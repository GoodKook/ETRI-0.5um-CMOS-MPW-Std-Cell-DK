magic
tech scmos
magscale 1 2
timestamp 0
<< metal1 >>
<< metal1 >>
rect 437 0 438 1
rect 436 0 437 1
rect 395 0 396 1
rect 394 0 395 1
rect 393 0 394 1
rect 437 1 438 2
rect 436 1 437 2
rect 435 1 436 2
rect 395 1 396 2
rect 394 1 395 2
rect 393 1 394 2
rect 437 2 438 3
rect 436 2 437 3
rect 435 2 436 3
rect 395 2 396 3
rect 394 2 395 3
rect 393 2 394 3
rect 437 3 438 4
rect 436 3 437 4
rect 435 3 436 4
rect 395 3 396 4
rect 394 3 395 4
rect 393 3 394 4
rect 437 4 438 5
rect 436 4 437 5
rect 435 4 436 5
rect 396 4 397 5
rect 395 4 396 5
rect 394 4 395 5
rect 393 4 394 5
rect 437 5 438 6
rect 436 5 437 6
rect 435 5 436 6
rect 434 5 435 6
rect 433 5 434 6
rect 397 5 398 6
rect 396 5 397 6
rect 395 5 396 6
rect 394 5 395 6
rect 393 5 394 6
rect 437 6 438 7
rect 436 6 437 7
rect 435 6 436 7
rect 434 6 435 7
rect 433 6 434 7
rect 432 6 433 7
rect 431 6 432 7
rect 430 6 431 7
rect 429 6 430 7
rect 428 6 429 7
rect 427 6 428 7
rect 426 6 427 7
rect 425 6 426 7
rect 424 6 425 7
rect 423 6 424 7
rect 422 6 423 7
rect 421 6 422 7
rect 420 6 421 7
rect 419 6 420 7
rect 418 6 419 7
rect 417 6 418 7
rect 416 6 417 7
rect 415 6 416 7
rect 414 6 415 7
rect 413 6 414 7
rect 412 6 413 7
rect 411 6 412 7
rect 410 6 411 7
rect 409 6 410 7
rect 408 6 409 7
rect 407 6 408 7
rect 406 6 407 7
rect 405 6 406 7
rect 404 6 405 7
rect 403 6 404 7
rect 402 6 403 7
rect 401 6 402 7
rect 400 6 401 7
rect 399 6 400 7
rect 398 6 399 7
rect 397 6 398 7
rect 396 6 397 7
rect 395 6 396 7
rect 394 6 395 7
rect 393 6 394 7
rect 437 7 438 8
rect 436 7 437 8
rect 435 7 436 8
rect 434 7 435 8
rect 433 7 434 8
rect 432 7 433 8
rect 431 7 432 8
rect 430 7 431 8
rect 429 7 430 8
rect 428 7 429 8
rect 427 7 428 8
rect 426 7 427 8
rect 425 7 426 8
rect 424 7 425 8
rect 423 7 424 8
rect 422 7 423 8
rect 421 7 422 8
rect 420 7 421 8
rect 419 7 420 8
rect 418 7 419 8
rect 417 7 418 8
rect 416 7 417 8
rect 415 7 416 8
rect 414 7 415 8
rect 413 7 414 8
rect 412 7 413 8
rect 411 7 412 8
rect 410 7 411 8
rect 409 7 410 8
rect 408 7 409 8
rect 407 7 408 8
rect 406 7 407 8
rect 405 7 406 8
rect 404 7 405 8
rect 403 7 404 8
rect 402 7 403 8
rect 401 7 402 8
rect 400 7 401 8
rect 399 7 400 8
rect 398 7 399 8
rect 397 7 398 8
rect 396 7 397 8
rect 395 7 396 8
rect 394 7 395 8
rect 393 7 394 8
rect 437 8 438 9
rect 436 8 437 9
rect 435 8 436 9
rect 434 8 435 9
rect 433 8 434 9
rect 432 8 433 9
rect 431 8 432 9
rect 430 8 431 9
rect 429 8 430 9
rect 428 8 429 9
rect 427 8 428 9
rect 426 8 427 9
rect 425 8 426 9
rect 424 8 425 9
rect 423 8 424 9
rect 422 8 423 9
rect 421 8 422 9
rect 420 8 421 9
rect 419 8 420 9
rect 418 8 419 9
rect 417 8 418 9
rect 416 8 417 9
rect 415 8 416 9
rect 414 8 415 9
rect 413 8 414 9
rect 412 8 413 9
rect 411 8 412 9
rect 410 8 411 9
rect 409 8 410 9
rect 408 8 409 9
rect 407 8 408 9
rect 406 8 407 9
rect 405 8 406 9
rect 404 8 405 9
rect 403 8 404 9
rect 402 8 403 9
rect 401 8 402 9
rect 400 8 401 9
rect 399 8 400 9
rect 398 8 399 9
rect 397 8 398 9
rect 396 8 397 9
rect 395 8 396 9
rect 394 8 395 9
rect 393 8 394 9
rect 437 9 438 10
rect 436 9 437 10
rect 435 9 436 10
rect 434 9 435 10
rect 433 9 434 10
rect 432 9 433 10
rect 431 9 432 10
rect 430 9 431 10
rect 429 9 430 10
rect 428 9 429 10
rect 427 9 428 10
rect 426 9 427 10
rect 425 9 426 10
rect 424 9 425 10
rect 423 9 424 10
rect 422 9 423 10
rect 421 9 422 10
rect 420 9 421 10
rect 419 9 420 10
rect 418 9 419 10
rect 417 9 418 10
rect 416 9 417 10
rect 415 9 416 10
rect 414 9 415 10
rect 413 9 414 10
rect 412 9 413 10
rect 411 9 412 10
rect 410 9 411 10
rect 409 9 410 10
rect 408 9 409 10
rect 407 9 408 10
rect 406 9 407 10
rect 405 9 406 10
rect 404 9 405 10
rect 403 9 404 10
rect 402 9 403 10
rect 401 9 402 10
rect 400 9 401 10
rect 399 9 400 10
rect 398 9 399 10
rect 397 9 398 10
rect 396 9 397 10
rect 395 9 396 10
rect 394 9 395 10
rect 393 9 394 10
rect 437 10 438 11
rect 436 10 437 11
rect 435 10 436 11
rect 434 10 435 11
rect 433 10 434 11
rect 432 10 433 11
rect 431 10 432 11
rect 430 10 431 11
rect 429 10 430 11
rect 428 10 429 11
rect 427 10 428 11
rect 426 10 427 11
rect 425 10 426 11
rect 424 10 425 11
rect 423 10 424 11
rect 422 10 423 11
rect 421 10 422 11
rect 420 10 421 11
rect 419 10 420 11
rect 418 10 419 11
rect 417 10 418 11
rect 416 10 417 11
rect 415 10 416 11
rect 414 10 415 11
rect 413 10 414 11
rect 412 10 413 11
rect 411 10 412 11
rect 410 10 411 11
rect 409 10 410 11
rect 408 10 409 11
rect 407 10 408 11
rect 406 10 407 11
rect 405 10 406 11
rect 404 10 405 11
rect 403 10 404 11
rect 402 10 403 11
rect 401 10 402 11
rect 400 10 401 11
rect 399 10 400 11
rect 398 10 399 11
rect 397 10 398 11
rect 396 10 397 11
rect 395 10 396 11
rect 394 10 395 11
rect 393 10 394 11
rect 437 11 438 12
rect 436 11 437 12
rect 435 11 436 12
rect 434 11 435 12
rect 433 11 434 12
rect 432 11 433 12
rect 431 11 432 12
rect 430 11 431 12
rect 429 11 430 12
rect 428 11 429 12
rect 427 11 428 12
rect 426 11 427 12
rect 425 11 426 12
rect 424 11 425 12
rect 423 11 424 12
rect 422 11 423 12
rect 421 11 422 12
rect 420 11 421 12
rect 419 11 420 12
rect 418 11 419 12
rect 417 11 418 12
rect 416 11 417 12
rect 415 11 416 12
rect 414 11 415 12
rect 413 11 414 12
rect 412 11 413 12
rect 411 11 412 12
rect 410 11 411 12
rect 409 11 410 12
rect 408 11 409 12
rect 407 11 408 12
rect 406 11 407 12
rect 405 11 406 12
rect 404 11 405 12
rect 403 11 404 12
rect 402 11 403 12
rect 401 11 402 12
rect 400 11 401 12
rect 399 11 400 12
rect 398 11 399 12
rect 397 11 398 12
rect 396 11 397 12
rect 395 11 396 12
rect 394 11 395 12
rect 393 11 394 12
rect 437 12 438 13
rect 436 12 437 13
rect 435 12 436 13
rect 434 12 435 13
rect 433 12 434 13
rect 432 12 433 13
rect 431 12 432 13
rect 430 12 431 13
rect 429 12 430 13
rect 428 12 429 13
rect 427 12 428 13
rect 426 12 427 13
rect 425 12 426 13
rect 424 12 425 13
rect 423 12 424 13
rect 422 12 423 13
rect 421 12 422 13
rect 420 12 421 13
rect 419 12 420 13
rect 418 12 419 13
rect 417 12 418 13
rect 416 12 417 13
rect 415 12 416 13
rect 414 12 415 13
rect 413 12 414 13
rect 412 12 413 13
rect 411 12 412 13
rect 410 12 411 13
rect 409 12 410 13
rect 408 12 409 13
rect 407 12 408 13
rect 406 12 407 13
rect 405 12 406 13
rect 404 12 405 13
rect 403 12 404 13
rect 402 12 403 13
rect 401 12 402 13
rect 400 12 401 13
rect 399 12 400 13
rect 398 12 399 13
rect 397 12 398 13
rect 396 12 397 13
rect 395 12 396 13
rect 394 12 395 13
rect 393 12 394 13
rect 437 13 438 14
rect 436 13 437 14
rect 435 13 436 14
rect 434 13 435 14
rect 433 13 434 14
rect 432 13 433 14
rect 431 13 432 14
rect 430 13 431 14
rect 429 13 430 14
rect 428 13 429 14
rect 427 13 428 14
rect 426 13 427 14
rect 425 13 426 14
rect 424 13 425 14
rect 423 13 424 14
rect 422 13 423 14
rect 421 13 422 14
rect 420 13 421 14
rect 419 13 420 14
rect 418 13 419 14
rect 417 13 418 14
rect 416 13 417 14
rect 415 13 416 14
rect 414 13 415 14
rect 413 13 414 14
rect 412 13 413 14
rect 411 13 412 14
rect 410 13 411 14
rect 409 13 410 14
rect 408 13 409 14
rect 407 13 408 14
rect 406 13 407 14
rect 405 13 406 14
rect 404 13 405 14
rect 403 13 404 14
rect 402 13 403 14
rect 401 13 402 14
rect 400 13 401 14
rect 399 13 400 14
rect 398 13 399 14
rect 397 13 398 14
rect 396 13 397 14
rect 395 13 396 14
rect 394 13 395 14
rect 393 13 394 14
rect 437 14 438 15
rect 436 14 437 15
rect 435 14 436 15
rect 434 14 435 15
rect 433 14 434 15
rect 432 14 433 15
rect 431 14 432 15
rect 430 14 431 15
rect 429 14 430 15
rect 428 14 429 15
rect 427 14 428 15
rect 426 14 427 15
rect 425 14 426 15
rect 424 14 425 15
rect 423 14 424 15
rect 422 14 423 15
rect 421 14 422 15
rect 420 14 421 15
rect 419 14 420 15
rect 418 14 419 15
rect 417 14 418 15
rect 416 14 417 15
rect 415 14 416 15
rect 414 14 415 15
rect 413 14 414 15
rect 412 14 413 15
rect 411 14 412 15
rect 410 14 411 15
rect 409 14 410 15
rect 408 14 409 15
rect 407 14 408 15
rect 406 14 407 15
rect 405 14 406 15
rect 404 14 405 15
rect 403 14 404 15
rect 402 14 403 15
rect 401 14 402 15
rect 400 14 401 15
rect 399 14 400 15
rect 398 14 399 15
rect 397 14 398 15
rect 396 14 397 15
rect 395 14 396 15
rect 394 14 395 15
rect 393 14 394 15
rect 437 15 438 16
rect 436 15 437 16
rect 435 15 436 16
rect 434 15 435 16
rect 433 15 434 16
rect 416 15 417 16
rect 415 15 416 16
rect 414 15 415 16
rect 397 15 398 16
rect 396 15 397 16
rect 395 15 396 16
rect 394 15 395 16
rect 393 15 394 16
rect 437 16 438 17
rect 436 16 437 17
rect 435 16 436 17
rect 434 16 435 17
rect 416 16 417 17
rect 415 16 416 17
rect 414 16 415 17
rect 413 16 414 17
rect 396 16 397 17
rect 395 16 396 17
rect 394 16 395 17
rect 393 16 394 17
rect 437 17 438 18
rect 436 17 437 18
rect 435 17 436 18
rect 417 17 418 18
rect 416 17 417 18
rect 415 17 416 18
rect 414 17 415 18
rect 413 17 414 18
rect 395 17 396 18
rect 394 17 395 18
rect 393 17 394 18
rect 437 18 438 19
rect 436 18 437 19
rect 435 18 436 19
rect 418 18 419 19
rect 417 18 418 19
rect 416 18 417 19
rect 415 18 416 19
rect 414 18 415 19
rect 413 18 414 19
rect 412 18 413 19
rect 395 18 396 19
rect 394 18 395 19
rect 393 18 394 19
rect 437 19 438 20
rect 436 19 437 20
rect 435 19 436 20
rect 419 19 420 20
rect 418 19 419 20
rect 417 19 418 20
rect 416 19 417 20
rect 415 19 416 20
rect 414 19 415 20
rect 413 19 414 20
rect 412 19 413 20
rect 411 19 412 20
rect 395 19 396 20
rect 394 19 395 20
rect 393 19 394 20
rect 437 20 438 21
rect 436 20 437 21
rect 435 20 436 21
rect 421 20 422 21
rect 420 20 421 21
rect 419 20 420 21
rect 418 20 419 21
rect 417 20 418 21
rect 416 20 417 21
rect 415 20 416 21
rect 414 20 415 21
rect 413 20 414 21
rect 412 20 413 21
rect 411 20 412 21
rect 410 20 411 21
rect 395 20 396 21
rect 394 20 395 21
rect 393 20 394 21
rect 422 21 423 22
rect 421 21 422 22
rect 420 21 421 22
rect 419 21 420 22
rect 418 21 419 22
rect 417 21 418 22
rect 416 21 417 22
rect 415 21 416 22
rect 414 21 415 22
rect 413 21 414 22
rect 412 21 413 22
rect 411 21 412 22
rect 410 21 411 22
rect 409 21 410 22
rect 424 22 425 23
rect 423 22 424 23
rect 422 22 423 23
rect 421 22 422 23
rect 420 22 421 23
rect 419 22 420 23
rect 418 22 419 23
rect 417 22 418 23
rect 416 22 417 23
rect 415 22 416 23
rect 414 22 415 23
rect 413 22 414 23
rect 412 22 413 23
rect 411 22 412 23
rect 410 22 411 23
rect 409 22 410 23
rect 408 22 409 23
rect 425 23 426 24
rect 424 23 425 24
rect 423 23 424 24
rect 422 23 423 24
rect 421 23 422 24
rect 420 23 421 24
rect 419 23 420 24
rect 418 23 419 24
rect 417 23 418 24
rect 416 23 417 24
rect 415 23 416 24
rect 414 23 415 24
rect 413 23 414 24
rect 412 23 413 24
rect 411 23 412 24
rect 410 23 411 24
rect 409 23 410 24
rect 408 23 409 24
rect 407 23 408 24
rect 427 24 428 25
rect 426 24 427 25
rect 425 24 426 25
rect 424 24 425 25
rect 423 24 424 25
rect 422 24 423 25
rect 421 24 422 25
rect 420 24 421 25
rect 419 24 420 25
rect 418 24 419 25
rect 417 24 418 25
rect 416 24 417 25
rect 415 24 416 25
rect 414 24 415 25
rect 413 24 414 25
rect 412 24 413 25
rect 411 24 412 25
rect 409 24 410 25
rect 408 24 409 25
rect 407 24 408 25
rect 406 24 407 25
rect 428 25 429 26
rect 427 25 428 26
rect 426 25 427 26
rect 425 25 426 26
rect 424 25 425 26
rect 423 25 424 26
rect 422 25 423 26
rect 421 25 422 26
rect 420 25 421 26
rect 419 25 420 26
rect 418 25 419 26
rect 417 25 418 26
rect 416 25 417 26
rect 415 25 416 26
rect 414 25 415 26
rect 413 25 414 26
rect 408 25 409 26
rect 407 25 408 26
rect 406 25 407 26
rect 405 25 406 26
rect 429 26 430 27
rect 428 26 429 27
rect 427 26 428 27
rect 426 26 427 27
rect 425 26 426 27
rect 424 26 425 27
rect 423 26 424 27
rect 422 26 423 27
rect 421 26 422 27
rect 420 26 421 27
rect 419 26 420 27
rect 418 26 419 27
rect 417 26 418 27
rect 416 26 417 27
rect 415 26 416 27
rect 414 26 415 27
rect 407 26 408 27
rect 406 26 407 27
rect 405 26 406 27
rect 404 26 405 27
rect 431 27 432 28
rect 430 27 431 28
rect 429 27 430 28
rect 428 27 429 28
rect 427 27 428 28
rect 426 27 427 28
rect 425 27 426 28
rect 424 27 425 28
rect 423 27 424 28
rect 422 27 423 28
rect 421 27 422 28
rect 420 27 421 28
rect 419 27 420 28
rect 418 27 419 28
rect 417 27 418 28
rect 416 27 417 28
rect 415 27 416 28
rect 406 27 407 28
rect 405 27 406 28
rect 404 27 405 28
rect 403 27 404 28
rect 402 27 403 28
rect 395 27 396 28
rect 394 27 395 28
rect 393 27 394 28
rect 432 28 433 29
rect 431 28 432 29
rect 430 28 431 29
rect 429 28 430 29
rect 428 28 429 29
rect 427 28 428 29
rect 426 28 427 29
rect 425 28 426 29
rect 424 28 425 29
rect 423 28 424 29
rect 422 28 423 29
rect 421 28 422 29
rect 420 28 421 29
rect 419 28 420 29
rect 418 28 419 29
rect 417 28 418 29
rect 405 28 406 29
rect 404 28 405 29
rect 403 28 404 29
rect 402 28 403 29
rect 401 28 402 29
rect 395 28 396 29
rect 394 28 395 29
rect 393 28 394 29
rect 434 29 435 30
rect 433 29 434 30
rect 432 29 433 30
rect 431 29 432 30
rect 430 29 431 30
rect 429 29 430 30
rect 428 29 429 30
rect 427 29 428 30
rect 426 29 427 30
rect 425 29 426 30
rect 424 29 425 30
rect 423 29 424 30
rect 422 29 423 30
rect 421 29 422 30
rect 420 29 421 30
rect 419 29 420 30
rect 418 29 419 30
rect 404 29 405 30
rect 403 29 404 30
rect 402 29 403 30
rect 401 29 402 30
rect 400 29 401 30
rect 395 29 396 30
rect 394 29 395 30
rect 393 29 394 30
rect 435 30 436 31
rect 434 30 435 31
rect 433 30 434 31
rect 432 30 433 31
rect 431 30 432 31
rect 430 30 431 31
rect 429 30 430 31
rect 428 30 429 31
rect 427 30 428 31
rect 426 30 427 31
rect 425 30 426 31
rect 424 30 425 31
rect 423 30 424 31
rect 422 30 423 31
rect 421 30 422 31
rect 420 30 421 31
rect 403 30 404 31
rect 402 30 403 31
rect 401 30 402 31
rect 400 30 401 31
rect 399 30 400 31
rect 398 30 399 31
rect 395 30 396 31
rect 394 30 395 31
rect 393 30 394 31
rect 437 31 438 32
rect 436 31 437 32
rect 435 31 436 32
rect 434 31 435 32
rect 433 31 434 32
rect 432 31 433 32
rect 431 31 432 32
rect 430 31 431 32
rect 429 31 430 32
rect 428 31 429 32
rect 427 31 428 32
rect 426 31 427 32
rect 425 31 426 32
rect 424 31 425 32
rect 423 31 424 32
rect 422 31 423 32
rect 421 31 422 32
rect 402 31 403 32
rect 401 31 402 32
rect 400 31 401 32
rect 399 31 400 32
rect 398 31 399 32
rect 397 31 398 32
rect 396 31 397 32
rect 395 31 396 32
rect 394 31 395 32
rect 393 31 394 32
rect 437 32 438 33
rect 436 32 437 33
rect 435 32 436 33
rect 434 32 435 33
rect 433 32 434 33
rect 432 32 433 33
rect 431 32 432 33
rect 430 32 431 33
rect 429 32 430 33
rect 428 32 429 33
rect 427 32 428 33
rect 426 32 427 33
rect 425 32 426 33
rect 424 32 425 33
rect 423 32 424 33
rect 422 32 423 33
rect 401 32 402 33
rect 400 32 401 33
rect 399 32 400 33
rect 398 32 399 33
rect 397 32 398 33
rect 396 32 397 33
rect 395 32 396 33
rect 394 32 395 33
rect 393 32 394 33
rect 437 33 438 34
rect 436 33 437 34
rect 435 33 436 34
rect 434 33 435 34
rect 433 33 434 34
rect 432 33 433 34
rect 431 33 432 34
rect 430 33 431 34
rect 429 33 430 34
rect 428 33 429 34
rect 427 33 428 34
rect 426 33 427 34
rect 425 33 426 34
rect 424 33 425 34
rect 400 33 401 34
rect 399 33 400 34
rect 398 33 399 34
rect 397 33 398 34
rect 396 33 397 34
rect 395 33 396 34
rect 394 33 395 34
rect 393 33 394 34
rect 437 34 438 35
rect 436 34 437 35
rect 435 34 436 35
rect 434 34 435 35
rect 433 34 434 35
rect 432 34 433 35
rect 431 34 432 35
rect 430 34 431 35
rect 429 34 430 35
rect 428 34 429 35
rect 427 34 428 35
rect 426 34 427 35
rect 425 34 426 35
rect 399 34 400 35
rect 398 34 399 35
rect 397 34 398 35
rect 396 34 397 35
rect 395 34 396 35
rect 394 34 395 35
rect 393 34 394 35
rect 437 35 438 36
rect 436 35 437 36
rect 435 35 436 36
rect 434 35 435 36
rect 433 35 434 36
rect 432 35 433 36
rect 431 35 432 36
rect 430 35 431 36
rect 429 35 430 36
rect 428 35 429 36
rect 427 35 428 36
rect 426 35 427 36
rect 398 35 399 36
rect 397 35 398 36
rect 396 35 397 36
rect 395 35 396 36
rect 394 35 395 36
rect 393 35 394 36
rect 437 36 438 37
rect 436 36 437 37
rect 435 36 436 37
rect 434 36 435 37
rect 433 36 434 37
rect 432 36 433 37
rect 431 36 432 37
rect 430 36 431 37
rect 429 36 430 37
rect 428 36 429 37
rect 398 36 399 37
rect 397 36 398 37
rect 396 36 397 37
rect 395 36 396 37
rect 394 36 395 37
rect 393 36 394 37
rect 437 37 438 38
rect 436 37 437 38
rect 435 37 436 38
rect 434 37 435 38
rect 433 37 434 38
rect 432 37 433 38
rect 431 37 432 38
rect 430 37 431 38
rect 429 37 430 38
rect 397 37 398 38
rect 396 37 397 38
rect 395 37 396 38
rect 394 37 395 38
rect 393 37 394 38
rect 437 38 438 39
rect 436 38 437 39
rect 435 38 436 39
rect 434 38 435 39
rect 433 38 434 39
rect 432 38 433 39
rect 431 38 432 39
rect 430 38 431 39
rect 396 38 397 39
rect 395 38 396 39
rect 394 38 395 39
rect 393 38 394 39
rect 437 39 438 40
rect 436 39 437 40
rect 435 39 436 40
rect 434 39 435 40
rect 433 39 434 40
rect 432 39 433 40
rect 431 39 432 40
rect 396 39 397 40
rect 395 39 396 40
rect 394 39 395 40
rect 393 39 394 40
rect 437 40 438 41
rect 436 40 437 41
rect 435 40 436 41
rect 434 40 435 41
rect 433 40 434 41
rect 396 40 397 41
rect 395 40 396 41
rect 394 40 395 41
rect 393 40 394 41
rect 437 41 438 42
rect 436 41 437 42
rect 435 41 436 42
rect 434 41 435 42
rect 433 41 434 42
rect 395 41 396 42
rect 394 41 395 42
rect 393 41 394 42
rect 437 42 438 43
rect 436 42 437 43
rect 435 42 436 43
rect 434 42 435 43
rect 395 42 396 43
rect 394 42 395 43
rect 393 42 394 43
rect 437 43 438 44
rect 436 43 437 44
rect 435 43 436 44
rect 395 43 396 44
rect 394 43 395 44
rect 393 43 394 44
rect 437 44 438 45
rect 436 44 437 45
rect 435 44 436 45
rect 395 44 396 45
rect 394 44 395 45
rect 393 44 394 45
rect 437 45 438 46
rect 436 45 437 46
rect 435 45 436 46
rect 89 47 90 48
rect 88 47 89 48
rect 87 47 88 48
rect 86 47 87 48
rect 85 47 86 48
rect 84 47 85 48
rect 91 48 92 49
rect 90 48 91 49
rect 89 48 90 49
rect 88 48 89 49
rect 87 48 88 49
rect 86 48 87 49
rect 85 48 86 49
rect 84 48 85 49
rect 83 48 84 49
rect 82 48 83 49
rect 92 49 93 50
rect 91 49 92 50
rect 90 49 91 50
rect 89 49 90 50
rect 88 49 89 50
rect 87 49 88 50
rect 86 49 87 50
rect 85 49 86 50
rect 84 49 85 50
rect 83 49 84 50
rect 82 49 83 50
rect 81 49 82 50
rect 394 50 395 51
rect 393 50 394 51
rect 92 50 93 51
rect 91 50 92 51
rect 90 50 91 51
rect 89 50 90 51
rect 88 50 89 51
rect 87 50 88 51
rect 86 50 87 51
rect 85 50 86 51
rect 84 50 85 51
rect 83 50 84 51
rect 82 50 83 51
rect 81 50 82 51
rect 80 50 81 51
rect 395 51 396 52
rect 394 51 395 52
rect 393 51 394 52
rect 93 51 94 52
rect 92 51 93 52
rect 91 51 92 52
rect 90 51 91 52
rect 89 51 90 52
rect 88 51 89 52
rect 87 51 88 52
rect 86 51 87 52
rect 85 51 86 52
rect 84 51 85 52
rect 83 51 84 52
rect 82 51 83 52
rect 81 51 82 52
rect 80 51 81 52
rect 79 51 80 52
rect 395 52 396 53
rect 394 52 395 53
rect 393 52 394 53
rect 93 52 94 53
rect 92 52 93 53
rect 91 52 92 53
rect 90 52 91 53
rect 89 52 90 53
rect 88 52 89 53
rect 87 52 88 53
rect 86 52 87 53
rect 85 52 86 53
rect 84 52 85 53
rect 83 52 84 53
rect 82 52 83 53
rect 81 52 82 53
rect 80 52 81 53
rect 79 52 80 53
rect 78 52 79 53
rect 395 53 396 54
rect 394 53 395 54
rect 393 53 394 54
rect 93 53 94 54
rect 92 53 93 54
rect 91 53 92 54
rect 90 53 91 54
rect 89 53 90 54
rect 88 53 89 54
rect 87 53 88 54
rect 86 53 87 54
rect 85 53 86 54
rect 84 53 85 54
rect 83 53 84 54
rect 82 53 83 54
rect 81 53 82 54
rect 80 53 81 54
rect 79 53 80 54
rect 78 53 79 54
rect 77 53 78 54
rect 396 54 397 55
rect 395 54 396 55
rect 394 54 395 55
rect 393 54 394 55
rect 105 54 106 55
rect 92 54 93 55
rect 91 54 92 55
rect 90 54 91 55
rect 89 54 90 55
rect 88 54 89 55
rect 87 54 88 55
rect 86 54 87 55
rect 85 54 86 55
rect 84 54 85 55
rect 83 54 84 55
rect 82 54 83 55
rect 81 54 82 55
rect 80 54 81 55
rect 79 54 80 55
rect 78 54 79 55
rect 77 54 78 55
rect 76 54 77 55
rect 397 55 398 56
rect 396 55 397 56
rect 395 55 396 56
rect 394 55 395 56
rect 393 55 394 56
rect 108 55 109 56
rect 107 55 108 56
rect 106 55 107 56
rect 105 55 106 56
rect 104 55 105 56
rect 103 55 104 56
rect 102 55 103 56
rect 92 55 93 56
rect 91 55 92 56
rect 90 55 91 56
rect 89 55 90 56
rect 88 55 89 56
rect 87 55 88 56
rect 86 55 87 56
rect 85 55 86 56
rect 84 55 85 56
rect 83 55 84 56
rect 82 55 83 56
rect 81 55 82 56
rect 80 55 81 56
rect 79 55 80 56
rect 78 55 79 56
rect 77 55 78 56
rect 76 55 77 56
rect 398 56 399 57
rect 397 56 398 57
rect 396 56 397 57
rect 395 56 396 57
rect 394 56 395 57
rect 393 56 394 57
rect 110 56 111 57
rect 109 56 110 57
rect 108 56 109 57
rect 107 56 108 57
rect 106 56 107 57
rect 105 56 106 57
rect 104 56 105 57
rect 103 56 104 57
rect 102 56 103 57
rect 101 56 102 57
rect 100 56 101 57
rect 92 56 93 57
rect 91 56 92 57
rect 90 56 91 57
rect 89 56 90 57
rect 88 56 89 57
rect 87 56 88 57
rect 86 56 87 57
rect 85 56 86 57
rect 84 56 85 57
rect 83 56 84 57
rect 82 56 83 57
rect 81 56 82 57
rect 80 56 81 57
rect 79 56 80 57
rect 78 56 79 57
rect 77 56 78 57
rect 76 56 77 57
rect 75 56 76 57
rect 400 57 401 58
rect 399 57 400 58
rect 398 57 399 58
rect 397 57 398 58
rect 396 57 397 58
rect 395 57 396 58
rect 394 57 395 58
rect 393 57 394 58
rect 112 57 113 58
rect 111 57 112 58
rect 110 57 111 58
rect 109 57 110 58
rect 108 57 109 58
rect 107 57 108 58
rect 106 57 107 58
rect 105 57 106 58
rect 104 57 105 58
rect 103 57 104 58
rect 102 57 103 58
rect 101 57 102 58
rect 100 57 101 58
rect 99 57 100 58
rect 92 57 93 58
rect 91 57 92 58
rect 90 57 91 58
rect 89 57 90 58
rect 88 57 89 58
rect 87 57 88 58
rect 86 57 87 58
rect 85 57 86 58
rect 84 57 85 58
rect 83 57 84 58
rect 82 57 83 58
rect 81 57 82 58
rect 80 57 81 58
rect 79 57 80 58
rect 78 57 79 58
rect 77 57 78 58
rect 76 57 77 58
rect 75 57 76 58
rect 74 57 75 58
rect 402 58 403 59
rect 401 58 402 59
rect 400 58 401 59
rect 399 58 400 59
rect 398 58 399 59
rect 397 58 398 59
rect 396 58 397 59
rect 395 58 396 59
rect 394 58 395 59
rect 393 58 394 59
rect 114 58 115 59
rect 113 58 114 59
rect 112 58 113 59
rect 111 58 112 59
rect 110 58 111 59
rect 109 58 110 59
rect 108 58 109 59
rect 107 58 108 59
rect 106 58 107 59
rect 105 58 106 59
rect 104 58 105 59
rect 103 58 104 59
rect 102 58 103 59
rect 101 58 102 59
rect 100 58 101 59
rect 99 58 100 59
rect 98 58 99 59
rect 91 58 92 59
rect 90 58 91 59
rect 89 58 90 59
rect 88 58 89 59
rect 87 58 88 59
rect 86 58 87 59
rect 85 58 86 59
rect 84 58 85 59
rect 83 58 84 59
rect 82 58 83 59
rect 81 58 82 59
rect 80 58 81 59
rect 79 58 80 59
rect 78 58 79 59
rect 77 58 78 59
rect 76 58 77 59
rect 75 58 76 59
rect 74 58 75 59
rect 403 59 404 60
rect 402 59 403 60
rect 401 59 402 60
rect 400 59 401 60
rect 399 59 400 60
rect 398 59 399 60
rect 397 59 398 60
rect 396 59 397 60
rect 395 59 396 60
rect 394 59 395 60
rect 393 59 394 60
rect 115 59 116 60
rect 114 59 115 60
rect 113 59 114 60
rect 112 59 113 60
rect 111 59 112 60
rect 110 59 111 60
rect 109 59 110 60
rect 108 59 109 60
rect 107 59 108 60
rect 106 59 107 60
rect 105 59 106 60
rect 104 59 105 60
rect 103 59 104 60
rect 102 59 103 60
rect 101 59 102 60
rect 100 59 101 60
rect 99 59 100 60
rect 98 59 99 60
rect 97 59 98 60
rect 91 59 92 60
rect 90 59 91 60
rect 89 59 90 60
rect 88 59 89 60
rect 87 59 88 60
rect 86 59 87 60
rect 85 59 86 60
rect 84 59 85 60
rect 83 59 84 60
rect 82 59 83 60
rect 81 59 82 60
rect 80 59 81 60
rect 79 59 80 60
rect 78 59 79 60
rect 77 59 78 60
rect 76 59 77 60
rect 75 59 76 60
rect 74 59 75 60
rect 73 59 74 60
rect 405 60 406 61
rect 404 60 405 61
rect 403 60 404 61
rect 402 60 403 61
rect 401 60 402 61
rect 400 60 401 61
rect 399 60 400 61
rect 398 60 399 61
rect 397 60 398 61
rect 396 60 397 61
rect 395 60 396 61
rect 394 60 395 61
rect 393 60 394 61
rect 116 60 117 61
rect 115 60 116 61
rect 114 60 115 61
rect 113 60 114 61
rect 112 60 113 61
rect 111 60 112 61
rect 110 60 111 61
rect 109 60 110 61
rect 108 60 109 61
rect 107 60 108 61
rect 106 60 107 61
rect 105 60 106 61
rect 104 60 105 61
rect 103 60 104 61
rect 102 60 103 61
rect 101 60 102 61
rect 100 60 101 61
rect 99 60 100 61
rect 98 60 99 61
rect 97 60 98 61
rect 96 60 97 61
rect 91 60 92 61
rect 90 60 91 61
rect 89 60 90 61
rect 88 60 89 61
rect 87 60 88 61
rect 86 60 87 61
rect 85 60 86 61
rect 84 60 85 61
rect 83 60 84 61
rect 82 60 83 61
rect 81 60 82 61
rect 80 60 81 61
rect 79 60 80 61
rect 78 60 79 61
rect 77 60 78 61
rect 76 60 77 61
rect 75 60 76 61
rect 74 60 75 61
rect 73 60 74 61
rect 437 61 438 62
rect 436 61 437 62
rect 407 61 408 62
rect 406 61 407 62
rect 405 61 406 62
rect 404 61 405 62
rect 403 61 404 62
rect 402 61 403 62
rect 401 61 402 62
rect 400 61 401 62
rect 399 61 400 62
rect 398 61 399 62
rect 397 61 398 62
rect 396 61 397 62
rect 395 61 396 62
rect 394 61 395 62
rect 393 61 394 62
rect 117 61 118 62
rect 116 61 117 62
rect 115 61 116 62
rect 114 61 115 62
rect 113 61 114 62
rect 112 61 113 62
rect 111 61 112 62
rect 110 61 111 62
rect 109 61 110 62
rect 108 61 109 62
rect 107 61 108 62
rect 106 61 107 62
rect 105 61 106 62
rect 104 61 105 62
rect 103 61 104 62
rect 102 61 103 62
rect 101 61 102 62
rect 100 61 101 62
rect 99 61 100 62
rect 98 61 99 62
rect 97 61 98 62
rect 96 61 97 62
rect 95 61 96 62
rect 90 61 91 62
rect 89 61 90 62
rect 88 61 89 62
rect 87 61 88 62
rect 86 61 87 62
rect 85 61 86 62
rect 84 61 85 62
rect 83 61 84 62
rect 82 61 83 62
rect 81 61 82 62
rect 80 61 81 62
rect 79 61 80 62
rect 78 61 79 62
rect 77 61 78 62
rect 76 61 77 62
rect 75 61 76 62
rect 74 61 75 62
rect 73 61 74 62
rect 72 61 73 62
rect 437 62 438 63
rect 436 62 437 63
rect 435 62 436 63
rect 409 62 410 63
rect 408 62 409 63
rect 407 62 408 63
rect 406 62 407 63
rect 405 62 406 63
rect 404 62 405 63
rect 403 62 404 63
rect 402 62 403 63
rect 401 62 402 63
rect 400 62 401 63
rect 399 62 400 63
rect 398 62 399 63
rect 397 62 398 63
rect 396 62 397 63
rect 395 62 396 63
rect 394 62 395 63
rect 393 62 394 63
rect 118 62 119 63
rect 117 62 118 63
rect 116 62 117 63
rect 115 62 116 63
rect 114 62 115 63
rect 113 62 114 63
rect 112 62 113 63
rect 111 62 112 63
rect 110 62 111 63
rect 109 62 110 63
rect 108 62 109 63
rect 107 62 108 63
rect 106 62 107 63
rect 105 62 106 63
rect 104 62 105 63
rect 103 62 104 63
rect 102 62 103 63
rect 101 62 102 63
rect 100 62 101 63
rect 99 62 100 63
rect 98 62 99 63
rect 97 62 98 63
rect 96 62 97 63
rect 95 62 96 63
rect 94 62 95 63
rect 90 62 91 63
rect 89 62 90 63
rect 88 62 89 63
rect 87 62 88 63
rect 86 62 87 63
rect 85 62 86 63
rect 84 62 85 63
rect 83 62 84 63
rect 82 62 83 63
rect 81 62 82 63
rect 80 62 81 63
rect 79 62 80 63
rect 78 62 79 63
rect 77 62 78 63
rect 76 62 77 63
rect 75 62 76 63
rect 74 62 75 63
rect 73 62 74 63
rect 72 62 73 63
rect 71 62 72 63
rect 437 63 438 64
rect 436 63 437 64
rect 435 63 436 64
rect 410 63 411 64
rect 409 63 410 64
rect 408 63 409 64
rect 407 63 408 64
rect 406 63 407 64
rect 405 63 406 64
rect 404 63 405 64
rect 403 63 404 64
rect 402 63 403 64
rect 401 63 402 64
rect 400 63 401 64
rect 399 63 400 64
rect 398 63 399 64
rect 397 63 398 64
rect 396 63 397 64
rect 395 63 396 64
rect 394 63 395 64
rect 393 63 394 64
rect 119 63 120 64
rect 118 63 119 64
rect 117 63 118 64
rect 116 63 117 64
rect 115 63 116 64
rect 114 63 115 64
rect 113 63 114 64
rect 112 63 113 64
rect 111 63 112 64
rect 110 63 111 64
rect 109 63 110 64
rect 108 63 109 64
rect 107 63 108 64
rect 106 63 107 64
rect 105 63 106 64
rect 104 63 105 64
rect 103 63 104 64
rect 102 63 103 64
rect 101 63 102 64
rect 100 63 101 64
rect 99 63 100 64
rect 98 63 99 64
rect 97 63 98 64
rect 96 63 97 64
rect 95 63 96 64
rect 94 63 95 64
rect 93 63 94 64
rect 89 63 90 64
rect 88 63 89 64
rect 87 63 88 64
rect 86 63 87 64
rect 85 63 86 64
rect 84 63 85 64
rect 83 63 84 64
rect 82 63 83 64
rect 81 63 82 64
rect 80 63 81 64
rect 79 63 80 64
rect 78 63 79 64
rect 77 63 78 64
rect 76 63 77 64
rect 75 63 76 64
rect 74 63 75 64
rect 73 63 74 64
rect 72 63 73 64
rect 71 63 72 64
rect 437 64 438 65
rect 436 64 437 65
rect 435 64 436 65
rect 412 64 413 65
rect 411 64 412 65
rect 410 64 411 65
rect 409 64 410 65
rect 408 64 409 65
rect 407 64 408 65
rect 406 64 407 65
rect 405 64 406 65
rect 404 64 405 65
rect 403 64 404 65
rect 402 64 403 65
rect 401 64 402 65
rect 400 64 401 65
rect 399 64 400 65
rect 398 64 399 65
rect 397 64 398 65
rect 396 64 397 65
rect 395 64 396 65
rect 394 64 395 65
rect 393 64 394 65
rect 120 64 121 65
rect 119 64 120 65
rect 118 64 119 65
rect 117 64 118 65
rect 116 64 117 65
rect 115 64 116 65
rect 114 64 115 65
rect 113 64 114 65
rect 112 64 113 65
rect 111 64 112 65
rect 110 64 111 65
rect 109 64 110 65
rect 108 64 109 65
rect 107 64 108 65
rect 106 64 107 65
rect 105 64 106 65
rect 104 64 105 65
rect 103 64 104 65
rect 102 64 103 65
rect 101 64 102 65
rect 100 64 101 65
rect 99 64 100 65
rect 98 64 99 65
rect 97 64 98 65
rect 96 64 97 65
rect 95 64 96 65
rect 94 64 95 65
rect 93 64 94 65
rect 92 64 93 65
rect 89 64 90 65
rect 88 64 89 65
rect 87 64 88 65
rect 86 64 87 65
rect 85 64 86 65
rect 84 64 85 65
rect 83 64 84 65
rect 82 64 83 65
rect 81 64 82 65
rect 80 64 81 65
rect 79 64 80 65
rect 78 64 79 65
rect 77 64 78 65
rect 76 64 77 65
rect 75 64 76 65
rect 74 64 75 65
rect 73 64 74 65
rect 72 64 73 65
rect 71 64 72 65
rect 70 64 71 65
rect 437 65 438 66
rect 436 65 437 66
rect 435 65 436 66
rect 414 65 415 66
rect 413 65 414 66
rect 412 65 413 66
rect 411 65 412 66
rect 410 65 411 66
rect 409 65 410 66
rect 408 65 409 66
rect 407 65 408 66
rect 406 65 407 66
rect 405 65 406 66
rect 404 65 405 66
rect 403 65 404 66
rect 402 65 403 66
rect 401 65 402 66
rect 400 65 401 66
rect 399 65 400 66
rect 398 65 399 66
rect 397 65 398 66
rect 396 65 397 66
rect 395 65 396 66
rect 394 65 395 66
rect 393 65 394 66
rect 121 65 122 66
rect 120 65 121 66
rect 119 65 120 66
rect 118 65 119 66
rect 117 65 118 66
rect 116 65 117 66
rect 115 65 116 66
rect 114 65 115 66
rect 113 65 114 66
rect 112 65 113 66
rect 111 65 112 66
rect 110 65 111 66
rect 109 65 110 66
rect 108 65 109 66
rect 107 65 108 66
rect 106 65 107 66
rect 105 65 106 66
rect 104 65 105 66
rect 103 65 104 66
rect 102 65 103 66
rect 101 65 102 66
rect 100 65 101 66
rect 99 65 100 66
rect 98 65 99 66
rect 97 65 98 66
rect 96 65 97 66
rect 95 65 96 66
rect 94 65 95 66
rect 93 65 94 66
rect 92 65 93 66
rect 91 65 92 66
rect 88 65 89 66
rect 87 65 88 66
rect 86 65 87 66
rect 85 65 86 66
rect 84 65 85 66
rect 83 65 84 66
rect 82 65 83 66
rect 81 65 82 66
rect 80 65 81 66
rect 79 65 80 66
rect 78 65 79 66
rect 77 65 78 66
rect 76 65 77 66
rect 75 65 76 66
rect 74 65 75 66
rect 73 65 74 66
rect 72 65 73 66
rect 71 65 72 66
rect 70 65 71 66
rect 437 66 438 67
rect 436 66 437 67
rect 435 66 436 67
rect 434 66 435 67
rect 416 66 417 67
rect 415 66 416 67
rect 414 66 415 67
rect 413 66 414 67
rect 412 66 413 67
rect 411 66 412 67
rect 410 66 411 67
rect 409 66 410 67
rect 408 66 409 67
rect 407 66 408 67
rect 406 66 407 67
rect 405 66 406 67
rect 404 66 405 67
rect 403 66 404 67
rect 402 66 403 67
rect 401 66 402 67
rect 400 66 401 67
rect 399 66 400 67
rect 398 66 399 67
rect 396 66 397 67
rect 395 66 396 67
rect 394 66 395 67
rect 393 66 394 67
rect 121 66 122 67
rect 120 66 121 67
rect 119 66 120 67
rect 118 66 119 67
rect 117 66 118 67
rect 116 66 117 67
rect 115 66 116 67
rect 114 66 115 67
rect 113 66 114 67
rect 112 66 113 67
rect 111 66 112 67
rect 110 66 111 67
rect 109 66 110 67
rect 108 66 109 67
rect 107 66 108 67
rect 106 66 107 67
rect 105 66 106 67
rect 104 66 105 67
rect 103 66 104 67
rect 102 66 103 67
rect 101 66 102 67
rect 100 66 101 67
rect 99 66 100 67
rect 98 66 99 67
rect 97 66 98 67
rect 96 66 97 67
rect 95 66 96 67
rect 94 66 95 67
rect 93 66 94 67
rect 92 66 93 67
rect 91 66 92 67
rect 90 66 91 67
rect 88 66 89 67
rect 87 66 88 67
rect 86 66 87 67
rect 85 66 86 67
rect 84 66 85 67
rect 83 66 84 67
rect 82 66 83 67
rect 81 66 82 67
rect 80 66 81 67
rect 79 66 80 67
rect 78 66 79 67
rect 77 66 78 67
rect 76 66 77 67
rect 75 66 76 67
rect 74 66 75 67
rect 73 66 74 67
rect 72 66 73 67
rect 71 66 72 67
rect 70 66 71 67
rect 437 67 438 68
rect 436 67 437 68
rect 435 67 436 68
rect 434 67 435 68
rect 433 67 434 68
rect 432 67 433 68
rect 431 67 432 68
rect 430 67 431 68
rect 429 67 430 68
rect 428 67 429 68
rect 427 67 428 68
rect 426 67 427 68
rect 425 67 426 68
rect 424 67 425 68
rect 423 67 424 68
rect 422 67 423 68
rect 421 67 422 68
rect 420 67 421 68
rect 419 67 420 68
rect 418 67 419 68
rect 417 67 418 68
rect 416 67 417 68
rect 415 67 416 68
rect 414 67 415 68
rect 413 67 414 68
rect 412 67 413 68
rect 411 67 412 68
rect 410 67 411 68
rect 409 67 410 68
rect 408 67 409 68
rect 407 67 408 68
rect 406 67 407 68
rect 405 67 406 68
rect 404 67 405 68
rect 403 67 404 68
rect 402 67 403 68
rect 401 67 402 68
rect 400 67 401 68
rect 395 67 396 68
rect 394 67 395 68
rect 393 67 394 68
rect 122 67 123 68
rect 121 67 122 68
rect 120 67 121 68
rect 119 67 120 68
rect 118 67 119 68
rect 117 67 118 68
rect 116 67 117 68
rect 115 67 116 68
rect 114 67 115 68
rect 113 67 114 68
rect 112 67 113 68
rect 111 67 112 68
rect 110 67 111 68
rect 109 67 110 68
rect 108 67 109 68
rect 107 67 108 68
rect 106 67 107 68
rect 105 67 106 68
rect 104 67 105 68
rect 103 67 104 68
rect 102 67 103 68
rect 101 67 102 68
rect 100 67 101 68
rect 99 67 100 68
rect 98 67 99 68
rect 97 67 98 68
rect 96 67 97 68
rect 95 67 96 68
rect 94 67 95 68
rect 93 67 94 68
rect 92 67 93 68
rect 91 67 92 68
rect 90 67 91 68
rect 89 67 90 68
rect 87 67 88 68
rect 86 67 87 68
rect 85 67 86 68
rect 84 67 85 68
rect 83 67 84 68
rect 82 67 83 68
rect 81 67 82 68
rect 80 67 81 68
rect 79 67 80 68
rect 78 67 79 68
rect 77 67 78 68
rect 76 67 77 68
rect 75 67 76 68
rect 74 67 75 68
rect 73 67 74 68
rect 72 67 73 68
rect 71 67 72 68
rect 70 67 71 68
rect 69 67 70 68
rect 437 68 438 69
rect 436 68 437 69
rect 435 68 436 69
rect 434 68 435 69
rect 433 68 434 69
rect 432 68 433 69
rect 431 68 432 69
rect 430 68 431 69
rect 429 68 430 69
rect 428 68 429 69
rect 427 68 428 69
rect 426 68 427 69
rect 425 68 426 69
rect 424 68 425 69
rect 423 68 424 69
rect 422 68 423 69
rect 421 68 422 69
rect 420 68 421 69
rect 419 68 420 69
rect 418 68 419 69
rect 417 68 418 69
rect 416 68 417 69
rect 415 68 416 69
rect 414 68 415 69
rect 413 68 414 69
rect 412 68 413 69
rect 411 68 412 69
rect 410 68 411 69
rect 409 68 410 69
rect 408 68 409 69
rect 407 68 408 69
rect 406 68 407 69
rect 405 68 406 69
rect 404 68 405 69
rect 403 68 404 69
rect 402 68 403 69
rect 395 68 396 69
rect 394 68 395 69
rect 393 68 394 69
rect 122 68 123 69
rect 121 68 122 69
rect 120 68 121 69
rect 119 68 120 69
rect 118 68 119 69
rect 117 68 118 69
rect 116 68 117 69
rect 115 68 116 69
rect 114 68 115 69
rect 113 68 114 69
rect 112 68 113 69
rect 111 68 112 69
rect 110 68 111 69
rect 109 68 110 69
rect 108 68 109 69
rect 107 68 108 69
rect 106 68 107 69
rect 105 68 106 69
rect 104 68 105 69
rect 103 68 104 69
rect 102 68 103 69
rect 101 68 102 69
rect 100 68 101 69
rect 99 68 100 69
rect 98 68 99 69
rect 97 68 98 69
rect 96 68 97 69
rect 95 68 96 69
rect 94 68 95 69
rect 93 68 94 69
rect 92 68 93 69
rect 91 68 92 69
rect 90 68 91 69
rect 89 68 90 69
rect 88 68 89 69
rect 87 68 88 69
rect 86 68 87 69
rect 85 68 86 69
rect 84 68 85 69
rect 83 68 84 69
rect 82 68 83 69
rect 81 68 82 69
rect 80 68 81 69
rect 79 68 80 69
rect 78 68 79 69
rect 77 68 78 69
rect 76 68 77 69
rect 75 68 76 69
rect 74 68 75 69
rect 73 68 74 69
rect 72 68 73 69
rect 71 68 72 69
rect 70 68 71 69
rect 69 68 70 69
rect 437 69 438 70
rect 436 69 437 70
rect 435 69 436 70
rect 434 69 435 70
rect 433 69 434 70
rect 432 69 433 70
rect 431 69 432 70
rect 430 69 431 70
rect 429 69 430 70
rect 428 69 429 70
rect 427 69 428 70
rect 426 69 427 70
rect 425 69 426 70
rect 424 69 425 70
rect 423 69 424 70
rect 422 69 423 70
rect 421 69 422 70
rect 420 69 421 70
rect 419 69 420 70
rect 418 69 419 70
rect 417 69 418 70
rect 416 69 417 70
rect 415 69 416 70
rect 414 69 415 70
rect 413 69 414 70
rect 412 69 413 70
rect 411 69 412 70
rect 410 69 411 70
rect 409 69 410 70
rect 408 69 409 70
rect 407 69 408 70
rect 406 69 407 70
rect 405 69 406 70
rect 404 69 405 70
rect 395 69 396 70
rect 394 69 395 70
rect 393 69 394 70
rect 137 69 138 70
rect 136 69 137 70
rect 135 69 136 70
rect 134 69 135 70
rect 133 69 134 70
rect 132 69 133 70
rect 122 69 123 70
rect 121 69 122 70
rect 120 69 121 70
rect 119 69 120 70
rect 118 69 119 70
rect 117 69 118 70
rect 116 69 117 70
rect 115 69 116 70
rect 114 69 115 70
rect 113 69 114 70
rect 112 69 113 70
rect 111 69 112 70
rect 110 69 111 70
rect 109 69 110 70
rect 108 69 109 70
rect 107 69 108 70
rect 106 69 107 70
rect 105 69 106 70
rect 104 69 105 70
rect 103 69 104 70
rect 102 69 103 70
rect 101 69 102 70
rect 100 69 101 70
rect 99 69 100 70
rect 98 69 99 70
rect 97 69 98 70
rect 96 69 97 70
rect 95 69 96 70
rect 94 69 95 70
rect 93 69 94 70
rect 92 69 93 70
rect 91 69 92 70
rect 90 69 91 70
rect 89 69 90 70
rect 88 69 89 70
rect 87 69 88 70
rect 86 69 87 70
rect 85 69 86 70
rect 84 69 85 70
rect 83 69 84 70
rect 82 69 83 70
rect 81 69 82 70
rect 80 69 81 70
rect 79 69 80 70
rect 78 69 79 70
rect 77 69 78 70
rect 76 69 77 70
rect 75 69 76 70
rect 74 69 75 70
rect 73 69 74 70
rect 72 69 73 70
rect 71 69 72 70
rect 70 69 71 70
rect 69 69 70 70
rect 68 69 69 70
rect 437 70 438 71
rect 436 70 437 71
rect 435 70 436 71
rect 434 70 435 71
rect 433 70 434 71
rect 432 70 433 71
rect 431 70 432 71
rect 430 70 431 71
rect 429 70 430 71
rect 428 70 429 71
rect 427 70 428 71
rect 426 70 427 71
rect 425 70 426 71
rect 424 70 425 71
rect 423 70 424 71
rect 422 70 423 71
rect 421 70 422 71
rect 420 70 421 71
rect 419 70 420 71
rect 418 70 419 71
rect 417 70 418 71
rect 416 70 417 71
rect 415 70 416 71
rect 414 70 415 71
rect 413 70 414 71
rect 412 70 413 71
rect 411 70 412 71
rect 410 70 411 71
rect 409 70 410 71
rect 408 70 409 71
rect 407 70 408 71
rect 406 70 407 71
rect 140 70 141 71
rect 139 70 140 71
rect 138 70 139 71
rect 137 70 138 71
rect 136 70 137 71
rect 135 70 136 71
rect 134 70 135 71
rect 133 70 134 71
rect 132 70 133 71
rect 131 70 132 71
rect 130 70 131 71
rect 122 70 123 71
rect 121 70 122 71
rect 120 70 121 71
rect 119 70 120 71
rect 118 70 119 71
rect 117 70 118 71
rect 116 70 117 71
rect 115 70 116 71
rect 114 70 115 71
rect 113 70 114 71
rect 112 70 113 71
rect 111 70 112 71
rect 110 70 111 71
rect 109 70 110 71
rect 108 70 109 71
rect 107 70 108 71
rect 106 70 107 71
rect 105 70 106 71
rect 104 70 105 71
rect 103 70 104 71
rect 102 70 103 71
rect 101 70 102 71
rect 100 70 101 71
rect 99 70 100 71
rect 98 70 99 71
rect 97 70 98 71
rect 96 70 97 71
rect 95 70 96 71
rect 94 70 95 71
rect 93 70 94 71
rect 92 70 93 71
rect 91 70 92 71
rect 90 70 91 71
rect 89 70 90 71
rect 88 70 89 71
rect 87 70 88 71
rect 86 70 87 71
rect 85 70 86 71
rect 84 70 85 71
rect 83 70 84 71
rect 82 70 83 71
rect 81 70 82 71
rect 80 70 81 71
rect 79 70 80 71
rect 78 70 79 71
rect 77 70 78 71
rect 76 70 77 71
rect 75 70 76 71
rect 74 70 75 71
rect 73 70 74 71
rect 72 70 73 71
rect 71 70 72 71
rect 70 70 71 71
rect 69 70 70 71
rect 68 70 69 71
rect 437 71 438 72
rect 436 71 437 72
rect 435 71 436 72
rect 434 71 435 72
rect 433 71 434 72
rect 432 71 433 72
rect 431 71 432 72
rect 430 71 431 72
rect 429 71 430 72
rect 428 71 429 72
rect 427 71 428 72
rect 426 71 427 72
rect 425 71 426 72
rect 424 71 425 72
rect 423 71 424 72
rect 422 71 423 72
rect 421 71 422 72
rect 420 71 421 72
rect 419 71 420 72
rect 418 71 419 72
rect 417 71 418 72
rect 416 71 417 72
rect 415 71 416 72
rect 414 71 415 72
rect 413 71 414 72
rect 412 71 413 72
rect 411 71 412 72
rect 410 71 411 72
rect 409 71 410 72
rect 408 71 409 72
rect 142 71 143 72
rect 141 71 142 72
rect 140 71 141 72
rect 139 71 140 72
rect 138 71 139 72
rect 137 71 138 72
rect 136 71 137 72
rect 135 71 136 72
rect 134 71 135 72
rect 133 71 134 72
rect 132 71 133 72
rect 131 71 132 72
rect 130 71 131 72
rect 122 71 123 72
rect 121 71 122 72
rect 120 71 121 72
rect 119 71 120 72
rect 118 71 119 72
rect 117 71 118 72
rect 116 71 117 72
rect 115 71 116 72
rect 114 71 115 72
rect 113 71 114 72
rect 112 71 113 72
rect 111 71 112 72
rect 110 71 111 72
rect 109 71 110 72
rect 108 71 109 72
rect 107 71 108 72
rect 106 71 107 72
rect 105 71 106 72
rect 104 71 105 72
rect 103 71 104 72
rect 102 71 103 72
rect 101 71 102 72
rect 100 71 101 72
rect 99 71 100 72
rect 98 71 99 72
rect 97 71 98 72
rect 96 71 97 72
rect 95 71 96 72
rect 94 71 95 72
rect 93 71 94 72
rect 92 71 93 72
rect 91 71 92 72
rect 90 71 91 72
rect 89 71 90 72
rect 88 71 89 72
rect 87 71 88 72
rect 86 71 87 72
rect 85 71 86 72
rect 84 71 85 72
rect 83 71 84 72
rect 82 71 83 72
rect 81 71 82 72
rect 80 71 81 72
rect 79 71 80 72
rect 78 71 79 72
rect 77 71 78 72
rect 76 71 77 72
rect 75 71 76 72
rect 74 71 75 72
rect 73 71 74 72
rect 72 71 73 72
rect 71 71 72 72
rect 70 71 71 72
rect 69 71 70 72
rect 68 71 69 72
rect 67 71 68 72
rect 437 72 438 73
rect 436 72 437 73
rect 435 72 436 73
rect 434 72 435 73
rect 433 72 434 73
rect 432 72 433 73
rect 431 72 432 73
rect 430 72 431 73
rect 429 72 430 73
rect 428 72 429 73
rect 427 72 428 73
rect 426 72 427 73
rect 425 72 426 73
rect 424 72 425 73
rect 423 72 424 73
rect 422 72 423 73
rect 421 72 422 73
rect 420 72 421 73
rect 419 72 420 73
rect 418 72 419 73
rect 417 72 418 73
rect 416 72 417 73
rect 415 72 416 73
rect 414 72 415 73
rect 413 72 414 73
rect 412 72 413 73
rect 411 72 412 73
rect 410 72 411 73
rect 144 72 145 73
rect 143 72 144 73
rect 142 72 143 73
rect 141 72 142 73
rect 140 72 141 73
rect 139 72 140 73
rect 138 72 139 73
rect 137 72 138 73
rect 136 72 137 73
rect 135 72 136 73
rect 134 72 135 73
rect 133 72 134 73
rect 132 72 133 73
rect 131 72 132 73
rect 130 72 131 73
rect 129 72 130 73
rect 123 72 124 73
rect 122 72 123 73
rect 121 72 122 73
rect 120 72 121 73
rect 119 72 120 73
rect 118 72 119 73
rect 117 72 118 73
rect 116 72 117 73
rect 115 72 116 73
rect 114 72 115 73
rect 113 72 114 73
rect 112 72 113 73
rect 111 72 112 73
rect 110 72 111 73
rect 109 72 110 73
rect 108 72 109 73
rect 107 72 108 73
rect 106 72 107 73
rect 105 72 106 73
rect 104 72 105 73
rect 103 72 104 73
rect 102 72 103 73
rect 101 72 102 73
rect 100 72 101 73
rect 99 72 100 73
rect 98 72 99 73
rect 97 72 98 73
rect 96 72 97 73
rect 95 72 96 73
rect 94 72 95 73
rect 93 72 94 73
rect 92 72 93 73
rect 91 72 92 73
rect 90 72 91 73
rect 89 72 90 73
rect 88 72 89 73
rect 87 72 88 73
rect 86 72 87 73
rect 85 72 86 73
rect 84 72 85 73
rect 83 72 84 73
rect 82 72 83 73
rect 81 72 82 73
rect 80 72 81 73
rect 79 72 80 73
rect 78 72 79 73
rect 77 72 78 73
rect 76 72 77 73
rect 75 72 76 73
rect 74 72 75 73
rect 73 72 74 73
rect 72 72 73 73
rect 71 72 72 73
rect 70 72 71 73
rect 69 72 70 73
rect 68 72 69 73
rect 67 72 68 73
rect 437 73 438 74
rect 436 73 437 74
rect 435 73 436 74
rect 434 73 435 74
rect 433 73 434 74
rect 432 73 433 74
rect 431 73 432 74
rect 430 73 431 74
rect 429 73 430 74
rect 428 73 429 74
rect 427 73 428 74
rect 426 73 427 74
rect 425 73 426 74
rect 424 73 425 74
rect 423 73 424 74
rect 422 73 423 74
rect 421 73 422 74
rect 420 73 421 74
rect 419 73 420 74
rect 418 73 419 74
rect 417 73 418 74
rect 416 73 417 74
rect 415 73 416 74
rect 414 73 415 74
rect 413 73 414 74
rect 412 73 413 74
rect 145 73 146 74
rect 144 73 145 74
rect 143 73 144 74
rect 142 73 143 74
rect 141 73 142 74
rect 140 73 141 74
rect 139 73 140 74
rect 138 73 139 74
rect 137 73 138 74
rect 136 73 137 74
rect 135 73 136 74
rect 134 73 135 74
rect 133 73 134 74
rect 132 73 133 74
rect 131 73 132 74
rect 130 73 131 74
rect 129 73 130 74
rect 122 73 123 74
rect 121 73 122 74
rect 120 73 121 74
rect 119 73 120 74
rect 118 73 119 74
rect 117 73 118 74
rect 116 73 117 74
rect 115 73 116 74
rect 114 73 115 74
rect 113 73 114 74
rect 112 73 113 74
rect 111 73 112 74
rect 110 73 111 74
rect 109 73 110 74
rect 108 73 109 74
rect 107 73 108 74
rect 106 73 107 74
rect 105 73 106 74
rect 104 73 105 74
rect 103 73 104 74
rect 102 73 103 74
rect 101 73 102 74
rect 100 73 101 74
rect 99 73 100 74
rect 98 73 99 74
rect 97 73 98 74
rect 96 73 97 74
rect 95 73 96 74
rect 94 73 95 74
rect 93 73 94 74
rect 92 73 93 74
rect 91 73 92 74
rect 90 73 91 74
rect 89 73 90 74
rect 88 73 89 74
rect 87 73 88 74
rect 86 73 87 74
rect 85 73 86 74
rect 84 73 85 74
rect 83 73 84 74
rect 82 73 83 74
rect 81 73 82 74
rect 80 73 81 74
rect 79 73 80 74
rect 78 73 79 74
rect 77 73 78 74
rect 76 73 77 74
rect 75 73 76 74
rect 74 73 75 74
rect 73 73 74 74
rect 72 73 73 74
rect 71 73 72 74
rect 70 73 71 74
rect 69 73 70 74
rect 68 73 69 74
rect 67 73 68 74
rect 66 73 67 74
rect 437 74 438 75
rect 436 74 437 75
rect 435 74 436 75
rect 434 74 435 75
rect 433 74 434 75
rect 432 74 433 75
rect 431 74 432 75
rect 430 74 431 75
rect 429 74 430 75
rect 428 74 429 75
rect 427 74 428 75
rect 426 74 427 75
rect 425 74 426 75
rect 424 74 425 75
rect 423 74 424 75
rect 422 74 423 75
rect 421 74 422 75
rect 420 74 421 75
rect 419 74 420 75
rect 418 74 419 75
rect 417 74 418 75
rect 416 74 417 75
rect 415 74 416 75
rect 414 74 415 75
rect 147 74 148 75
rect 146 74 147 75
rect 145 74 146 75
rect 144 74 145 75
rect 143 74 144 75
rect 142 74 143 75
rect 141 74 142 75
rect 140 74 141 75
rect 139 74 140 75
rect 138 74 139 75
rect 137 74 138 75
rect 136 74 137 75
rect 135 74 136 75
rect 134 74 135 75
rect 133 74 134 75
rect 132 74 133 75
rect 131 74 132 75
rect 130 74 131 75
rect 129 74 130 75
rect 122 74 123 75
rect 121 74 122 75
rect 120 74 121 75
rect 119 74 120 75
rect 118 74 119 75
rect 117 74 118 75
rect 116 74 117 75
rect 115 74 116 75
rect 114 74 115 75
rect 113 74 114 75
rect 112 74 113 75
rect 111 74 112 75
rect 110 74 111 75
rect 109 74 110 75
rect 108 74 109 75
rect 107 74 108 75
rect 106 74 107 75
rect 105 74 106 75
rect 104 74 105 75
rect 103 74 104 75
rect 102 74 103 75
rect 101 74 102 75
rect 100 74 101 75
rect 99 74 100 75
rect 98 74 99 75
rect 97 74 98 75
rect 96 74 97 75
rect 95 74 96 75
rect 94 74 95 75
rect 93 74 94 75
rect 92 74 93 75
rect 91 74 92 75
rect 90 74 91 75
rect 89 74 90 75
rect 88 74 89 75
rect 87 74 88 75
rect 86 74 87 75
rect 85 74 86 75
rect 84 74 85 75
rect 83 74 84 75
rect 82 74 83 75
rect 81 74 82 75
rect 80 74 81 75
rect 79 74 80 75
rect 78 74 79 75
rect 77 74 78 75
rect 76 74 77 75
rect 75 74 76 75
rect 74 74 75 75
rect 73 74 74 75
rect 72 74 73 75
rect 71 74 72 75
rect 70 74 71 75
rect 69 74 70 75
rect 68 74 69 75
rect 67 74 68 75
rect 66 74 67 75
rect 437 75 438 76
rect 436 75 437 76
rect 435 75 436 76
rect 434 75 435 76
rect 433 75 434 76
rect 432 75 433 76
rect 431 75 432 76
rect 430 75 431 76
rect 429 75 430 76
rect 428 75 429 76
rect 427 75 428 76
rect 426 75 427 76
rect 425 75 426 76
rect 424 75 425 76
rect 423 75 424 76
rect 422 75 423 76
rect 421 75 422 76
rect 420 75 421 76
rect 419 75 420 76
rect 418 75 419 76
rect 417 75 418 76
rect 416 75 417 76
rect 415 75 416 76
rect 414 75 415 76
rect 413 75 414 76
rect 148 75 149 76
rect 147 75 148 76
rect 146 75 147 76
rect 145 75 146 76
rect 144 75 145 76
rect 143 75 144 76
rect 142 75 143 76
rect 141 75 142 76
rect 140 75 141 76
rect 139 75 140 76
rect 138 75 139 76
rect 137 75 138 76
rect 136 75 137 76
rect 135 75 136 76
rect 134 75 135 76
rect 133 75 134 76
rect 132 75 133 76
rect 131 75 132 76
rect 130 75 131 76
rect 129 75 130 76
rect 122 75 123 76
rect 121 75 122 76
rect 120 75 121 76
rect 119 75 120 76
rect 118 75 119 76
rect 117 75 118 76
rect 116 75 117 76
rect 115 75 116 76
rect 114 75 115 76
rect 113 75 114 76
rect 112 75 113 76
rect 111 75 112 76
rect 110 75 111 76
rect 109 75 110 76
rect 108 75 109 76
rect 107 75 108 76
rect 106 75 107 76
rect 105 75 106 76
rect 104 75 105 76
rect 103 75 104 76
rect 102 75 103 76
rect 101 75 102 76
rect 100 75 101 76
rect 99 75 100 76
rect 98 75 99 76
rect 97 75 98 76
rect 96 75 97 76
rect 95 75 96 76
rect 94 75 95 76
rect 93 75 94 76
rect 92 75 93 76
rect 91 75 92 76
rect 90 75 91 76
rect 89 75 90 76
rect 88 75 89 76
rect 87 75 88 76
rect 86 75 87 76
rect 85 75 86 76
rect 84 75 85 76
rect 83 75 84 76
rect 82 75 83 76
rect 81 75 82 76
rect 80 75 81 76
rect 79 75 80 76
rect 78 75 79 76
rect 77 75 78 76
rect 76 75 77 76
rect 75 75 76 76
rect 74 75 75 76
rect 73 75 74 76
rect 72 75 73 76
rect 71 75 72 76
rect 70 75 71 76
rect 69 75 70 76
rect 68 75 69 76
rect 67 75 68 76
rect 66 75 67 76
rect 65 75 66 76
rect 437 76 438 77
rect 436 76 437 77
rect 435 76 436 77
rect 434 76 435 77
rect 433 76 434 77
rect 432 76 433 77
rect 431 76 432 77
rect 430 76 431 77
rect 429 76 430 77
rect 428 76 429 77
rect 427 76 428 77
rect 426 76 427 77
rect 425 76 426 77
rect 424 76 425 77
rect 423 76 424 77
rect 422 76 423 77
rect 421 76 422 77
rect 420 76 421 77
rect 419 76 420 77
rect 418 76 419 77
rect 417 76 418 77
rect 416 76 417 77
rect 415 76 416 77
rect 414 76 415 77
rect 413 76 414 77
rect 412 76 413 77
rect 411 76 412 77
rect 150 76 151 77
rect 149 76 150 77
rect 148 76 149 77
rect 147 76 148 77
rect 146 76 147 77
rect 145 76 146 77
rect 144 76 145 77
rect 143 76 144 77
rect 142 76 143 77
rect 141 76 142 77
rect 140 76 141 77
rect 139 76 140 77
rect 138 76 139 77
rect 137 76 138 77
rect 136 76 137 77
rect 135 76 136 77
rect 134 76 135 77
rect 133 76 134 77
rect 132 76 133 77
rect 131 76 132 77
rect 130 76 131 77
rect 129 76 130 77
rect 122 76 123 77
rect 121 76 122 77
rect 120 76 121 77
rect 119 76 120 77
rect 118 76 119 77
rect 117 76 118 77
rect 116 76 117 77
rect 115 76 116 77
rect 114 76 115 77
rect 113 76 114 77
rect 112 76 113 77
rect 111 76 112 77
rect 110 76 111 77
rect 109 76 110 77
rect 108 76 109 77
rect 107 76 108 77
rect 106 76 107 77
rect 105 76 106 77
rect 104 76 105 77
rect 103 76 104 77
rect 102 76 103 77
rect 101 76 102 77
rect 100 76 101 77
rect 99 76 100 77
rect 98 76 99 77
rect 97 76 98 77
rect 96 76 97 77
rect 95 76 96 77
rect 94 76 95 77
rect 93 76 94 77
rect 92 76 93 77
rect 91 76 92 77
rect 90 76 91 77
rect 89 76 90 77
rect 88 76 89 77
rect 87 76 88 77
rect 86 76 87 77
rect 85 76 86 77
rect 84 76 85 77
rect 83 76 84 77
rect 82 76 83 77
rect 81 76 82 77
rect 80 76 81 77
rect 79 76 80 77
rect 78 76 79 77
rect 77 76 78 77
rect 76 76 77 77
rect 75 76 76 77
rect 74 76 75 77
rect 73 76 74 77
rect 72 76 73 77
rect 71 76 72 77
rect 70 76 71 77
rect 69 76 70 77
rect 68 76 69 77
rect 67 76 68 77
rect 66 76 67 77
rect 65 76 66 77
rect 437 77 438 78
rect 436 77 437 78
rect 435 77 436 78
rect 434 77 435 78
rect 415 77 416 78
rect 414 77 415 78
rect 413 77 414 78
rect 412 77 413 78
rect 411 77 412 78
rect 410 77 411 78
rect 409 77 410 78
rect 152 77 153 78
rect 151 77 152 78
rect 150 77 151 78
rect 149 77 150 78
rect 148 77 149 78
rect 147 77 148 78
rect 146 77 147 78
rect 145 77 146 78
rect 144 77 145 78
rect 143 77 144 78
rect 142 77 143 78
rect 141 77 142 78
rect 140 77 141 78
rect 139 77 140 78
rect 138 77 139 78
rect 137 77 138 78
rect 136 77 137 78
rect 135 77 136 78
rect 134 77 135 78
rect 133 77 134 78
rect 132 77 133 78
rect 131 77 132 78
rect 130 77 131 78
rect 129 77 130 78
rect 122 77 123 78
rect 121 77 122 78
rect 120 77 121 78
rect 119 77 120 78
rect 118 77 119 78
rect 117 77 118 78
rect 116 77 117 78
rect 115 77 116 78
rect 114 77 115 78
rect 113 77 114 78
rect 112 77 113 78
rect 111 77 112 78
rect 110 77 111 78
rect 109 77 110 78
rect 108 77 109 78
rect 107 77 108 78
rect 106 77 107 78
rect 105 77 106 78
rect 104 77 105 78
rect 103 77 104 78
rect 102 77 103 78
rect 101 77 102 78
rect 100 77 101 78
rect 99 77 100 78
rect 98 77 99 78
rect 97 77 98 78
rect 96 77 97 78
rect 95 77 96 78
rect 94 77 95 78
rect 93 77 94 78
rect 92 77 93 78
rect 91 77 92 78
rect 90 77 91 78
rect 89 77 90 78
rect 88 77 89 78
rect 87 77 88 78
rect 86 77 87 78
rect 85 77 86 78
rect 84 77 85 78
rect 83 77 84 78
rect 82 77 83 78
rect 81 77 82 78
rect 80 77 81 78
rect 79 77 80 78
rect 78 77 79 78
rect 77 77 78 78
rect 76 77 77 78
rect 75 77 76 78
rect 74 77 75 78
rect 73 77 74 78
rect 72 77 73 78
rect 71 77 72 78
rect 70 77 71 78
rect 69 77 70 78
rect 68 77 69 78
rect 67 77 68 78
rect 66 77 67 78
rect 65 77 66 78
rect 64 77 65 78
rect 437 78 438 79
rect 436 78 437 79
rect 435 78 436 79
rect 413 78 414 79
rect 412 78 413 79
rect 411 78 412 79
rect 410 78 411 79
rect 409 78 410 79
rect 408 78 409 79
rect 407 78 408 79
rect 395 78 396 79
rect 394 78 395 79
rect 393 78 394 79
rect 155 78 156 79
rect 154 78 155 79
rect 153 78 154 79
rect 152 78 153 79
rect 151 78 152 79
rect 150 78 151 79
rect 149 78 150 79
rect 148 78 149 79
rect 147 78 148 79
rect 146 78 147 79
rect 145 78 146 79
rect 144 78 145 79
rect 143 78 144 79
rect 142 78 143 79
rect 141 78 142 79
rect 140 78 141 79
rect 139 78 140 79
rect 138 78 139 79
rect 137 78 138 79
rect 136 78 137 79
rect 135 78 136 79
rect 134 78 135 79
rect 133 78 134 79
rect 132 78 133 79
rect 131 78 132 79
rect 130 78 131 79
rect 129 78 130 79
rect 122 78 123 79
rect 121 78 122 79
rect 120 78 121 79
rect 119 78 120 79
rect 118 78 119 79
rect 117 78 118 79
rect 116 78 117 79
rect 115 78 116 79
rect 114 78 115 79
rect 113 78 114 79
rect 112 78 113 79
rect 111 78 112 79
rect 110 78 111 79
rect 109 78 110 79
rect 108 78 109 79
rect 107 78 108 79
rect 106 78 107 79
rect 105 78 106 79
rect 104 78 105 79
rect 103 78 104 79
rect 102 78 103 79
rect 101 78 102 79
rect 100 78 101 79
rect 99 78 100 79
rect 98 78 99 79
rect 97 78 98 79
rect 96 78 97 79
rect 95 78 96 79
rect 94 78 95 79
rect 93 78 94 79
rect 92 78 93 79
rect 91 78 92 79
rect 90 78 91 79
rect 89 78 90 79
rect 88 78 89 79
rect 87 78 88 79
rect 86 78 87 79
rect 85 78 86 79
rect 84 78 85 79
rect 83 78 84 79
rect 82 78 83 79
rect 81 78 82 79
rect 80 78 81 79
rect 79 78 80 79
rect 78 78 79 79
rect 77 78 78 79
rect 76 78 77 79
rect 75 78 76 79
rect 74 78 75 79
rect 73 78 74 79
rect 72 78 73 79
rect 71 78 72 79
rect 70 78 71 79
rect 69 78 70 79
rect 68 78 69 79
rect 67 78 68 79
rect 66 78 67 79
rect 65 78 66 79
rect 64 78 65 79
rect 63 78 64 79
rect 458 79 459 80
rect 437 79 438 80
rect 436 79 437 80
rect 435 79 436 80
rect 411 79 412 80
rect 410 79 411 80
rect 409 79 410 80
rect 408 79 409 80
rect 407 79 408 80
rect 406 79 407 80
rect 405 79 406 80
rect 395 79 396 80
rect 394 79 395 80
rect 393 79 394 80
rect 157 79 158 80
rect 156 79 157 80
rect 155 79 156 80
rect 154 79 155 80
rect 153 79 154 80
rect 152 79 153 80
rect 151 79 152 80
rect 150 79 151 80
rect 149 79 150 80
rect 148 79 149 80
rect 147 79 148 80
rect 146 79 147 80
rect 145 79 146 80
rect 144 79 145 80
rect 143 79 144 80
rect 142 79 143 80
rect 141 79 142 80
rect 140 79 141 80
rect 139 79 140 80
rect 138 79 139 80
rect 137 79 138 80
rect 136 79 137 80
rect 135 79 136 80
rect 134 79 135 80
rect 133 79 134 80
rect 132 79 133 80
rect 131 79 132 80
rect 130 79 131 80
rect 129 79 130 80
rect 122 79 123 80
rect 121 79 122 80
rect 120 79 121 80
rect 119 79 120 80
rect 118 79 119 80
rect 117 79 118 80
rect 116 79 117 80
rect 115 79 116 80
rect 114 79 115 80
rect 113 79 114 80
rect 112 79 113 80
rect 111 79 112 80
rect 110 79 111 80
rect 109 79 110 80
rect 108 79 109 80
rect 107 79 108 80
rect 106 79 107 80
rect 105 79 106 80
rect 104 79 105 80
rect 103 79 104 80
rect 102 79 103 80
rect 101 79 102 80
rect 100 79 101 80
rect 99 79 100 80
rect 98 79 99 80
rect 97 79 98 80
rect 96 79 97 80
rect 95 79 96 80
rect 94 79 95 80
rect 93 79 94 80
rect 92 79 93 80
rect 91 79 92 80
rect 90 79 91 80
rect 89 79 90 80
rect 88 79 89 80
rect 87 79 88 80
rect 86 79 87 80
rect 85 79 86 80
rect 84 79 85 80
rect 83 79 84 80
rect 82 79 83 80
rect 81 79 82 80
rect 80 79 81 80
rect 79 79 80 80
rect 78 79 79 80
rect 77 79 78 80
rect 76 79 77 80
rect 75 79 76 80
rect 74 79 75 80
rect 73 79 74 80
rect 72 79 73 80
rect 71 79 72 80
rect 70 79 71 80
rect 69 79 70 80
rect 68 79 69 80
rect 67 79 68 80
rect 66 79 67 80
rect 65 79 66 80
rect 64 79 65 80
rect 63 79 64 80
rect 458 80 459 81
rect 437 80 438 81
rect 436 80 437 81
rect 435 80 436 81
rect 409 80 410 81
rect 408 80 409 81
rect 407 80 408 81
rect 406 80 407 81
rect 405 80 406 81
rect 404 80 405 81
rect 403 80 404 81
rect 395 80 396 81
rect 394 80 395 81
rect 393 80 394 81
rect 159 80 160 81
rect 158 80 159 81
rect 157 80 158 81
rect 156 80 157 81
rect 155 80 156 81
rect 154 80 155 81
rect 153 80 154 81
rect 152 80 153 81
rect 151 80 152 81
rect 150 80 151 81
rect 149 80 150 81
rect 148 80 149 81
rect 147 80 148 81
rect 146 80 147 81
rect 145 80 146 81
rect 144 80 145 81
rect 143 80 144 81
rect 142 80 143 81
rect 141 80 142 81
rect 140 80 141 81
rect 139 80 140 81
rect 138 80 139 81
rect 137 80 138 81
rect 136 80 137 81
rect 135 80 136 81
rect 134 80 135 81
rect 133 80 134 81
rect 132 80 133 81
rect 131 80 132 81
rect 130 80 131 81
rect 129 80 130 81
rect 122 80 123 81
rect 121 80 122 81
rect 120 80 121 81
rect 119 80 120 81
rect 118 80 119 81
rect 117 80 118 81
rect 116 80 117 81
rect 115 80 116 81
rect 114 80 115 81
rect 113 80 114 81
rect 112 80 113 81
rect 111 80 112 81
rect 110 80 111 81
rect 109 80 110 81
rect 108 80 109 81
rect 107 80 108 81
rect 106 80 107 81
rect 105 80 106 81
rect 104 80 105 81
rect 103 80 104 81
rect 102 80 103 81
rect 101 80 102 81
rect 100 80 101 81
rect 99 80 100 81
rect 98 80 99 81
rect 97 80 98 81
rect 96 80 97 81
rect 95 80 96 81
rect 94 80 95 81
rect 93 80 94 81
rect 92 80 93 81
rect 91 80 92 81
rect 90 80 91 81
rect 89 80 90 81
rect 88 80 89 81
rect 87 80 88 81
rect 86 80 87 81
rect 85 80 86 81
rect 84 80 85 81
rect 83 80 84 81
rect 82 80 83 81
rect 81 80 82 81
rect 80 80 81 81
rect 79 80 80 81
rect 78 80 79 81
rect 77 80 78 81
rect 76 80 77 81
rect 75 80 76 81
rect 74 80 75 81
rect 73 80 74 81
rect 72 80 73 81
rect 71 80 72 81
rect 70 80 71 81
rect 69 80 70 81
rect 68 80 69 81
rect 67 80 68 81
rect 66 80 67 81
rect 65 80 66 81
rect 64 80 65 81
rect 63 80 64 81
rect 62 80 63 81
rect 459 81 460 82
rect 458 81 459 82
rect 437 81 438 82
rect 436 81 437 82
rect 435 81 436 82
rect 408 81 409 82
rect 407 81 408 82
rect 406 81 407 82
rect 405 81 406 82
rect 404 81 405 82
rect 403 81 404 82
rect 402 81 403 82
rect 401 81 402 82
rect 395 81 396 82
rect 394 81 395 82
rect 393 81 394 82
rect 223 81 224 82
rect 222 81 223 82
rect 221 81 222 82
rect 220 81 221 82
rect 219 81 220 82
rect 218 81 219 82
rect 217 81 218 82
rect 216 81 217 82
rect 215 81 216 82
rect 214 81 215 82
rect 213 81 214 82
rect 212 81 213 82
rect 211 81 212 82
rect 210 81 211 82
rect 209 81 210 82
rect 208 81 209 82
rect 207 81 208 82
rect 160 81 161 82
rect 159 81 160 82
rect 158 81 159 82
rect 157 81 158 82
rect 156 81 157 82
rect 155 81 156 82
rect 154 81 155 82
rect 153 81 154 82
rect 152 81 153 82
rect 151 81 152 82
rect 150 81 151 82
rect 149 81 150 82
rect 148 81 149 82
rect 147 81 148 82
rect 146 81 147 82
rect 145 81 146 82
rect 144 81 145 82
rect 143 81 144 82
rect 142 81 143 82
rect 141 81 142 82
rect 140 81 141 82
rect 139 81 140 82
rect 138 81 139 82
rect 137 81 138 82
rect 136 81 137 82
rect 135 81 136 82
rect 134 81 135 82
rect 133 81 134 82
rect 132 81 133 82
rect 131 81 132 82
rect 130 81 131 82
rect 129 81 130 82
rect 122 81 123 82
rect 121 81 122 82
rect 120 81 121 82
rect 119 81 120 82
rect 118 81 119 82
rect 117 81 118 82
rect 116 81 117 82
rect 115 81 116 82
rect 114 81 115 82
rect 113 81 114 82
rect 112 81 113 82
rect 111 81 112 82
rect 110 81 111 82
rect 109 81 110 82
rect 108 81 109 82
rect 107 81 108 82
rect 106 81 107 82
rect 105 81 106 82
rect 104 81 105 82
rect 103 81 104 82
rect 102 81 103 82
rect 101 81 102 82
rect 100 81 101 82
rect 99 81 100 82
rect 98 81 99 82
rect 97 81 98 82
rect 96 81 97 82
rect 95 81 96 82
rect 94 81 95 82
rect 93 81 94 82
rect 92 81 93 82
rect 91 81 92 82
rect 90 81 91 82
rect 89 81 90 82
rect 88 81 89 82
rect 87 81 88 82
rect 86 81 87 82
rect 85 81 86 82
rect 84 81 85 82
rect 83 81 84 82
rect 82 81 83 82
rect 81 81 82 82
rect 80 81 81 82
rect 79 81 80 82
rect 78 81 79 82
rect 77 81 78 82
rect 76 81 77 82
rect 75 81 76 82
rect 74 81 75 82
rect 73 81 74 82
rect 72 81 73 82
rect 71 81 72 82
rect 70 81 71 82
rect 69 81 70 82
rect 68 81 69 82
rect 67 81 68 82
rect 66 81 67 82
rect 65 81 66 82
rect 64 81 65 82
rect 63 81 64 82
rect 62 81 63 82
rect 474 82 475 83
rect 473 82 474 83
rect 472 82 473 83
rect 471 82 472 83
rect 470 82 471 83
rect 469 82 470 83
rect 468 82 469 83
rect 467 82 468 83
rect 466 82 467 83
rect 465 82 466 83
rect 464 82 465 83
rect 463 82 464 83
rect 462 82 463 83
rect 461 82 462 83
rect 460 82 461 83
rect 459 82 460 83
rect 458 82 459 83
rect 437 82 438 83
rect 436 82 437 83
rect 406 82 407 83
rect 405 82 406 83
rect 404 82 405 83
rect 403 82 404 83
rect 402 82 403 83
rect 401 82 402 83
rect 400 82 401 83
rect 399 82 400 83
rect 398 82 399 83
rect 397 82 398 83
rect 396 82 397 83
rect 395 82 396 83
rect 394 82 395 83
rect 393 82 394 83
rect 229 82 230 83
rect 228 82 229 83
rect 227 82 228 83
rect 226 82 227 83
rect 225 82 226 83
rect 224 82 225 83
rect 223 82 224 83
rect 222 82 223 83
rect 221 82 222 83
rect 220 82 221 83
rect 219 82 220 83
rect 218 82 219 83
rect 217 82 218 83
rect 216 82 217 83
rect 215 82 216 83
rect 214 82 215 83
rect 213 82 214 83
rect 212 82 213 83
rect 211 82 212 83
rect 210 82 211 83
rect 209 82 210 83
rect 208 82 209 83
rect 207 82 208 83
rect 206 82 207 83
rect 205 82 206 83
rect 204 82 205 83
rect 203 82 204 83
rect 202 82 203 83
rect 160 82 161 83
rect 159 82 160 83
rect 158 82 159 83
rect 157 82 158 83
rect 156 82 157 83
rect 155 82 156 83
rect 154 82 155 83
rect 153 82 154 83
rect 152 82 153 83
rect 151 82 152 83
rect 150 82 151 83
rect 149 82 150 83
rect 148 82 149 83
rect 147 82 148 83
rect 146 82 147 83
rect 145 82 146 83
rect 144 82 145 83
rect 143 82 144 83
rect 142 82 143 83
rect 141 82 142 83
rect 140 82 141 83
rect 139 82 140 83
rect 138 82 139 83
rect 137 82 138 83
rect 136 82 137 83
rect 135 82 136 83
rect 134 82 135 83
rect 133 82 134 83
rect 132 82 133 83
rect 131 82 132 83
rect 130 82 131 83
rect 129 82 130 83
rect 128 82 129 83
rect 121 82 122 83
rect 120 82 121 83
rect 119 82 120 83
rect 118 82 119 83
rect 117 82 118 83
rect 116 82 117 83
rect 115 82 116 83
rect 114 82 115 83
rect 113 82 114 83
rect 112 82 113 83
rect 111 82 112 83
rect 110 82 111 83
rect 109 82 110 83
rect 108 82 109 83
rect 107 82 108 83
rect 106 82 107 83
rect 105 82 106 83
rect 104 82 105 83
rect 103 82 104 83
rect 102 82 103 83
rect 101 82 102 83
rect 100 82 101 83
rect 99 82 100 83
rect 98 82 99 83
rect 97 82 98 83
rect 96 82 97 83
rect 95 82 96 83
rect 94 82 95 83
rect 93 82 94 83
rect 92 82 93 83
rect 91 82 92 83
rect 90 82 91 83
rect 89 82 90 83
rect 88 82 89 83
rect 87 82 88 83
rect 86 82 87 83
rect 85 82 86 83
rect 84 82 85 83
rect 83 82 84 83
rect 82 82 83 83
rect 81 82 82 83
rect 80 82 81 83
rect 79 82 80 83
rect 78 82 79 83
rect 77 82 78 83
rect 76 82 77 83
rect 75 82 76 83
rect 74 82 75 83
rect 73 82 74 83
rect 72 82 73 83
rect 71 82 72 83
rect 70 82 71 83
rect 69 82 70 83
rect 68 82 69 83
rect 67 82 68 83
rect 66 82 67 83
rect 65 82 66 83
rect 64 82 65 83
rect 63 82 64 83
rect 62 82 63 83
rect 61 82 62 83
rect 476 83 477 84
rect 475 83 476 84
rect 474 83 475 84
rect 473 83 474 84
rect 472 83 473 84
rect 471 83 472 84
rect 470 83 471 84
rect 469 83 470 84
rect 468 83 469 84
rect 467 83 468 84
rect 466 83 467 84
rect 465 83 466 84
rect 464 83 465 84
rect 463 83 464 84
rect 462 83 463 84
rect 461 83 462 84
rect 460 83 461 84
rect 459 83 460 84
rect 458 83 459 84
rect 437 83 438 84
rect 436 83 437 84
rect 404 83 405 84
rect 403 83 404 84
rect 402 83 403 84
rect 401 83 402 84
rect 400 83 401 84
rect 399 83 400 84
rect 398 83 399 84
rect 397 83 398 84
rect 396 83 397 84
rect 395 83 396 84
rect 394 83 395 84
rect 393 83 394 84
rect 233 83 234 84
rect 232 83 233 84
rect 231 83 232 84
rect 230 83 231 84
rect 229 83 230 84
rect 228 83 229 84
rect 227 83 228 84
rect 226 83 227 84
rect 225 83 226 84
rect 224 83 225 84
rect 223 83 224 84
rect 222 83 223 84
rect 221 83 222 84
rect 220 83 221 84
rect 219 83 220 84
rect 218 83 219 84
rect 217 83 218 84
rect 216 83 217 84
rect 215 83 216 84
rect 214 83 215 84
rect 213 83 214 84
rect 212 83 213 84
rect 211 83 212 84
rect 210 83 211 84
rect 209 83 210 84
rect 208 83 209 84
rect 207 83 208 84
rect 206 83 207 84
rect 205 83 206 84
rect 204 83 205 84
rect 203 83 204 84
rect 202 83 203 84
rect 201 83 202 84
rect 200 83 201 84
rect 199 83 200 84
rect 198 83 199 84
rect 160 83 161 84
rect 159 83 160 84
rect 158 83 159 84
rect 157 83 158 84
rect 156 83 157 84
rect 155 83 156 84
rect 154 83 155 84
rect 153 83 154 84
rect 152 83 153 84
rect 151 83 152 84
rect 150 83 151 84
rect 149 83 150 84
rect 148 83 149 84
rect 147 83 148 84
rect 146 83 147 84
rect 145 83 146 84
rect 144 83 145 84
rect 143 83 144 84
rect 142 83 143 84
rect 141 83 142 84
rect 140 83 141 84
rect 139 83 140 84
rect 138 83 139 84
rect 137 83 138 84
rect 136 83 137 84
rect 135 83 136 84
rect 134 83 135 84
rect 133 83 134 84
rect 132 83 133 84
rect 131 83 132 84
rect 130 83 131 84
rect 129 83 130 84
rect 128 83 129 84
rect 121 83 122 84
rect 120 83 121 84
rect 119 83 120 84
rect 118 83 119 84
rect 117 83 118 84
rect 116 83 117 84
rect 115 83 116 84
rect 114 83 115 84
rect 113 83 114 84
rect 112 83 113 84
rect 111 83 112 84
rect 110 83 111 84
rect 109 83 110 84
rect 108 83 109 84
rect 107 83 108 84
rect 106 83 107 84
rect 105 83 106 84
rect 104 83 105 84
rect 103 83 104 84
rect 102 83 103 84
rect 101 83 102 84
rect 100 83 101 84
rect 99 83 100 84
rect 98 83 99 84
rect 97 83 98 84
rect 96 83 97 84
rect 95 83 96 84
rect 94 83 95 84
rect 93 83 94 84
rect 92 83 93 84
rect 91 83 92 84
rect 90 83 91 84
rect 89 83 90 84
rect 88 83 89 84
rect 87 83 88 84
rect 86 83 87 84
rect 85 83 86 84
rect 84 83 85 84
rect 83 83 84 84
rect 82 83 83 84
rect 81 83 82 84
rect 80 83 81 84
rect 79 83 80 84
rect 78 83 79 84
rect 77 83 78 84
rect 76 83 77 84
rect 75 83 76 84
rect 74 83 75 84
rect 73 83 74 84
rect 72 83 73 84
rect 71 83 72 84
rect 70 83 71 84
rect 69 83 70 84
rect 68 83 69 84
rect 67 83 68 84
rect 66 83 67 84
rect 65 83 66 84
rect 64 83 65 84
rect 63 83 64 84
rect 62 83 63 84
rect 61 83 62 84
rect 60 83 61 84
rect 477 84 478 85
rect 476 84 477 85
rect 475 84 476 85
rect 474 84 475 85
rect 473 84 474 85
rect 472 84 473 85
rect 471 84 472 85
rect 470 84 471 85
rect 469 84 470 85
rect 468 84 469 85
rect 467 84 468 85
rect 466 84 467 85
rect 465 84 466 85
rect 464 84 465 85
rect 463 84 464 85
rect 462 84 463 85
rect 461 84 462 85
rect 460 84 461 85
rect 459 84 460 85
rect 458 84 459 85
rect 403 84 404 85
rect 402 84 403 85
rect 401 84 402 85
rect 400 84 401 85
rect 399 84 400 85
rect 398 84 399 85
rect 397 84 398 85
rect 396 84 397 85
rect 395 84 396 85
rect 394 84 395 85
rect 393 84 394 85
rect 236 84 237 85
rect 235 84 236 85
rect 234 84 235 85
rect 233 84 234 85
rect 232 84 233 85
rect 231 84 232 85
rect 230 84 231 85
rect 229 84 230 85
rect 228 84 229 85
rect 227 84 228 85
rect 226 84 227 85
rect 225 84 226 85
rect 224 84 225 85
rect 223 84 224 85
rect 222 84 223 85
rect 221 84 222 85
rect 220 84 221 85
rect 219 84 220 85
rect 218 84 219 85
rect 217 84 218 85
rect 216 84 217 85
rect 215 84 216 85
rect 214 84 215 85
rect 213 84 214 85
rect 212 84 213 85
rect 211 84 212 85
rect 210 84 211 85
rect 209 84 210 85
rect 208 84 209 85
rect 207 84 208 85
rect 206 84 207 85
rect 205 84 206 85
rect 204 84 205 85
rect 203 84 204 85
rect 202 84 203 85
rect 201 84 202 85
rect 200 84 201 85
rect 199 84 200 85
rect 198 84 199 85
rect 197 84 198 85
rect 196 84 197 85
rect 160 84 161 85
rect 159 84 160 85
rect 158 84 159 85
rect 157 84 158 85
rect 156 84 157 85
rect 155 84 156 85
rect 154 84 155 85
rect 153 84 154 85
rect 152 84 153 85
rect 151 84 152 85
rect 150 84 151 85
rect 149 84 150 85
rect 148 84 149 85
rect 147 84 148 85
rect 146 84 147 85
rect 145 84 146 85
rect 144 84 145 85
rect 143 84 144 85
rect 142 84 143 85
rect 141 84 142 85
rect 140 84 141 85
rect 139 84 140 85
rect 138 84 139 85
rect 137 84 138 85
rect 136 84 137 85
rect 135 84 136 85
rect 134 84 135 85
rect 133 84 134 85
rect 132 84 133 85
rect 131 84 132 85
rect 130 84 131 85
rect 129 84 130 85
rect 128 84 129 85
rect 121 84 122 85
rect 120 84 121 85
rect 119 84 120 85
rect 118 84 119 85
rect 117 84 118 85
rect 116 84 117 85
rect 115 84 116 85
rect 114 84 115 85
rect 113 84 114 85
rect 112 84 113 85
rect 111 84 112 85
rect 110 84 111 85
rect 109 84 110 85
rect 108 84 109 85
rect 107 84 108 85
rect 106 84 107 85
rect 105 84 106 85
rect 104 84 105 85
rect 103 84 104 85
rect 102 84 103 85
rect 101 84 102 85
rect 100 84 101 85
rect 99 84 100 85
rect 98 84 99 85
rect 97 84 98 85
rect 96 84 97 85
rect 95 84 96 85
rect 94 84 95 85
rect 93 84 94 85
rect 92 84 93 85
rect 91 84 92 85
rect 90 84 91 85
rect 89 84 90 85
rect 88 84 89 85
rect 87 84 88 85
rect 86 84 87 85
rect 85 84 86 85
rect 84 84 85 85
rect 83 84 84 85
rect 82 84 83 85
rect 81 84 82 85
rect 80 84 81 85
rect 79 84 80 85
rect 78 84 79 85
rect 77 84 78 85
rect 76 84 77 85
rect 75 84 76 85
rect 74 84 75 85
rect 73 84 74 85
rect 72 84 73 85
rect 71 84 72 85
rect 70 84 71 85
rect 69 84 70 85
rect 68 84 69 85
rect 67 84 68 85
rect 66 84 67 85
rect 65 84 66 85
rect 64 84 65 85
rect 63 84 64 85
rect 62 84 63 85
rect 61 84 62 85
rect 60 84 61 85
rect 478 85 479 86
rect 477 85 478 86
rect 476 85 477 86
rect 475 85 476 86
rect 474 85 475 86
rect 473 85 474 86
rect 472 85 473 86
rect 471 85 472 86
rect 470 85 471 86
rect 469 85 470 86
rect 468 85 469 86
rect 467 85 468 86
rect 466 85 467 86
rect 465 85 466 86
rect 464 85 465 86
rect 463 85 464 86
rect 462 85 463 86
rect 461 85 462 86
rect 460 85 461 86
rect 459 85 460 86
rect 458 85 459 86
rect 401 85 402 86
rect 400 85 401 86
rect 399 85 400 86
rect 398 85 399 86
rect 397 85 398 86
rect 396 85 397 86
rect 395 85 396 86
rect 394 85 395 86
rect 393 85 394 86
rect 239 85 240 86
rect 238 85 239 86
rect 237 85 238 86
rect 236 85 237 86
rect 235 85 236 86
rect 234 85 235 86
rect 233 85 234 86
rect 232 85 233 86
rect 231 85 232 86
rect 230 85 231 86
rect 229 85 230 86
rect 228 85 229 86
rect 227 85 228 86
rect 226 85 227 86
rect 225 85 226 86
rect 224 85 225 86
rect 223 85 224 86
rect 222 85 223 86
rect 221 85 222 86
rect 220 85 221 86
rect 219 85 220 86
rect 218 85 219 86
rect 217 85 218 86
rect 216 85 217 86
rect 215 85 216 86
rect 214 85 215 86
rect 213 85 214 86
rect 212 85 213 86
rect 211 85 212 86
rect 210 85 211 86
rect 209 85 210 86
rect 208 85 209 86
rect 207 85 208 86
rect 206 85 207 86
rect 205 85 206 86
rect 204 85 205 86
rect 203 85 204 86
rect 202 85 203 86
rect 201 85 202 86
rect 200 85 201 86
rect 199 85 200 86
rect 198 85 199 86
rect 197 85 198 86
rect 196 85 197 86
rect 195 85 196 86
rect 194 85 195 86
rect 160 85 161 86
rect 159 85 160 86
rect 158 85 159 86
rect 157 85 158 86
rect 156 85 157 86
rect 155 85 156 86
rect 154 85 155 86
rect 153 85 154 86
rect 152 85 153 86
rect 151 85 152 86
rect 150 85 151 86
rect 149 85 150 86
rect 148 85 149 86
rect 147 85 148 86
rect 146 85 147 86
rect 145 85 146 86
rect 144 85 145 86
rect 143 85 144 86
rect 142 85 143 86
rect 141 85 142 86
rect 140 85 141 86
rect 139 85 140 86
rect 138 85 139 86
rect 137 85 138 86
rect 136 85 137 86
rect 135 85 136 86
rect 134 85 135 86
rect 133 85 134 86
rect 132 85 133 86
rect 131 85 132 86
rect 130 85 131 86
rect 129 85 130 86
rect 128 85 129 86
rect 121 85 122 86
rect 120 85 121 86
rect 119 85 120 86
rect 118 85 119 86
rect 117 85 118 86
rect 116 85 117 86
rect 115 85 116 86
rect 114 85 115 86
rect 113 85 114 86
rect 112 85 113 86
rect 111 85 112 86
rect 110 85 111 86
rect 109 85 110 86
rect 108 85 109 86
rect 107 85 108 86
rect 106 85 107 86
rect 105 85 106 86
rect 104 85 105 86
rect 103 85 104 86
rect 102 85 103 86
rect 101 85 102 86
rect 100 85 101 86
rect 99 85 100 86
rect 98 85 99 86
rect 97 85 98 86
rect 96 85 97 86
rect 95 85 96 86
rect 94 85 95 86
rect 93 85 94 86
rect 92 85 93 86
rect 91 85 92 86
rect 90 85 91 86
rect 89 85 90 86
rect 88 85 89 86
rect 87 85 88 86
rect 86 85 87 86
rect 85 85 86 86
rect 84 85 85 86
rect 83 85 84 86
rect 82 85 83 86
rect 81 85 82 86
rect 80 85 81 86
rect 79 85 80 86
rect 78 85 79 86
rect 77 85 78 86
rect 76 85 77 86
rect 75 85 76 86
rect 74 85 75 86
rect 73 85 74 86
rect 72 85 73 86
rect 71 85 72 86
rect 70 85 71 86
rect 69 85 70 86
rect 68 85 69 86
rect 67 85 68 86
rect 66 85 67 86
rect 65 85 66 86
rect 64 85 65 86
rect 63 85 64 86
rect 62 85 63 86
rect 61 85 62 86
rect 60 85 61 86
rect 59 85 60 86
rect 479 86 480 87
rect 478 86 479 87
rect 477 86 478 87
rect 476 86 477 87
rect 475 86 476 87
rect 474 86 475 87
rect 473 86 474 87
rect 472 86 473 87
rect 471 86 472 87
rect 460 86 461 87
rect 459 86 460 87
rect 458 86 459 87
rect 399 86 400 87
rect 398 86 399 87
rect 397 86 398 87
rect 396 86 397 87
rect 395 86 396 87
rect 394 86 395 87
rect 393 86 394 87
rect 241 86 242 87
rect 240 86 241 87
rect 239 86 240 87
rect 238 86 239 87
rect 237 86 238 87
rect 236 86 237 87
rect 235 86 236 87
rect 234 86 235 87
rect 233 86 234 87
rect 232 86 233 87
rect 231 86 232 87
rect 230 86 231 87
rect 229 86 230 87
rect 228 86 229 87
rect 227 86 228 87
rect 226 86 227 87
rect 225 86 226 87
rect 224 86 225 87
rect 223 86 224 87
rect 222 86 223 87
rect 221 86 222 87
rect 220 86 221 87
rect 219 86 220 87
rect 218 86 219 87
rect 217 86 218 87
rect 216 86 217 87
rect 215 86 216 87
rect 214 86 215 87
rect 213 86 214 87
rect 212 86 213 87
rect 211 86 212 87
rect 210 86 211 87
rect 209 86 210 87
rect 208 86 209 87
rect 207 86 208 87
rect 206 86 207 87
rect 205 86 206 87
rect 204 86 205 87
rect 203 86 204 87
rect 202 86 203 87
rect 201 86 202 87
rect 200 86 201 87
rect 199 86 200 87
rect 198 86 199 87
rect 197 86 198 87
rect 196 86 197 87
rect 195 86 196 87
rect 194 86 195 87
rect 193 86 194 87
rect 192 86 193 87
rect 160 86 161 87
rect 159 86 160 87
rect 158 86 159 87
rect 157 86 158 87
rect 156 86 157 87
rect 155 86 156 87
rect 154 86 155 87
rect 153 86 154 87
rect 152 86 153 87
rect 151 86 152 87
rect 150 86 151 87
rect 149 86 150 87
rect 148 86 149 87
rect 147 86 148 87
rect 146 86 147 87
rect 145 86 146 87
rect 144 86 145 87
rect 143 86 144 87
rect 142 86 143 87
rect 141 86 142 87
rect 140 86 141 87
rect 139 86 140 87
rect 138 86 139 87
rect 137 86 138 87
rect 136 86 137 87
rect 135 86 136 87
rect 134 86 135 87
rect 133 86 134 87
rect 132 86 133 87
rect 131 86 132 87
rect 130 86 131 87
rect 129 86 130 87
rect 128 86 129 87
rect 121 86 122 87
rect 120 86 121 87
rect 119 86 120 87
rect 118 86 119 87
rect 117 86 118 87
rect 116 86 117 87
rect 115 86 116 87
rect 114 86 115 87
rect 113 86 114 87
rect 112 86 113 87
rect 111 86 112 87
rect 110 86 111 87
rect 109 86 110 87
rect 108 86 109 87
rect 107 86 108 87
rect 106 86 107 87
rect 105 86 106 87
rect 104 86 105 87
rect 103 86 104 87
rect 102 86 103 87
rect 101 86 102 87
rect 100 86 101 87
rect 99 86 100 87
rect 98 86 99 87
rect 97 86 98 87
rect 96 86 97 87
rect 95 86 96 87
rect 94 86 95 87
rect 93 86 94 87
rect 92 86 93 87
rect 91 86 92 87
rect 90 86 91 87
rect 89 86 90 87
rect 88 86 89 87
rect 87 86 88 87
rect 86 86 87 87
rect 85 86 86 87
rect 84 86 85 87
rect 83 86 84 87
rect 82 86 83 87
rect 81 86 82 87
rect 80 86 81 87
rect 79 86 80 87
rect 78 86 79 87
rect 77 86 78 87
rect 76 86 77 87
rect 75 86 76 87
rect 74 86 75 87
rect 73 86 74 87
rect 72 86 73 87
rect 71 86 72 87
rect 70 86 71 87
rect 69 86 70 87
rect 68 86 69 87
rect 67 86 68 87
rect 66 86 67 87
rect 65 86 66 87
rect 64 86 65 87
rect 63 86 64 87
rect 62 86 63 87
rect 61 86 62 87
rect 60 86 61 87
rect 59 86 60 87
rect 58 86 59 87
rect 479 87 480 88
rect 478 87 479 88
rect 477 87 478 88
rect 476 87 477 88
rect 475 87 476 88
rect 458 87 459 88
rect 398 87 399 88
rect 397 87 398 88
rect 396 87 397 88
rect 395 87 396 88
rect 394 87 395 88
rect 393 87 394 88
rect 244 87 245 88
rect 243 87 244 88
rect 242 87 243 88
rect 241 87 242 88
rect 240 87 241 88
rect 239 87 240 88
rect 238 87 239 88
rect 237 87 238 88
rect 236 87 237 88
rect 235 87 236 88
rect 234 87 235 88
rect 233 87 234 88
rect 232 87 233 88
rect 231 87 232 88
rect 230 87 231 88
rect 229 87 230 88
rect 228 87 229 88
rect 227 87 228 88
rect 226 87 227 88
rect 225 87 226 88
rect 224 87 225 88
rect 223 87 224 88
rect 222 87 223 88
rect 221 87 222 88
rect 220 87 221 88
rect 219 87 220 88
rect 218 87 219 88
rect 217 87 218 88
rect 216 87 217 88
rect 215 87 216 88
rect 214 87 215 88
rect 213 87 214 88
rect 212 87 213 88
rect 211 87 212 88
rect 210 87 211 88
rect 209 87 210 88
rect 208 87 209 88
rect 207 87 208 88
rect 206 87 207 88
rect 205 87 206 88
rect 204 87 205 88
rect 203 87 204 88
rect 202 87 203 88
rect 201 87 202 88
rect 200 87 201 88
rect 199 87 200 88
rect 198 87 199 88
rect 197 87 198 88
rect 196 87 197 88
rect 195 87 196 88
rect 194 87 195 88
rect 193 87 194 88
rect 192 87 193 88
rect 191 87 192 88
rect 190 87 191 88
rect 160 87 161 88
rect 159 87 160 88
rect 158 87 159 88
rect 157 87 158 88
rect 156 87 157 88
rect 155 87 156 88
rect 154 87 155 88
rect 153 87 154 88
rect 152 87 153 88
rect 151 87 152 88
rect 150 87 151 88
rect 149 87 150 88
rect 148 87 149 88
rect 147 87 148 88
rect 146 87 147 88
rect 145 87 146 88
rect 144 87 145 88
rect 143 87 144 88
rect 142 87 143 88
rect 141 87 142 88
rect 140 87 141 88
rect 139 87 140 88
rect 138 87 139 88
rect 137 87 138 88
rect 136 87 137 88
rect 135 87 136 88
rect 134 87 135 88
rect 133 87 134 88
rect 132 87 133 88
rect 131 87 132 88
rect 130 87 131 88
rect 129 87 130 88
rect 128 87 129 88
rect 121 87 122 88
rect 120 87 121 88
rect 119 87 120 88
rect 118 87 119 88
rect 117 87 118 88
rect 116 87 117 88
rect 115 87 116 88
rect 114 87 115 88
rect 113 87 114 88
rect 112 87 113 88
rect 111 87 112 88
rect 110 87 111 88
rect 109 87 110 88
rect 108 87 109 88
rect 107 87 108 88
rect 106 87 107 88
rect 105 87 106 88
rect 104 87 105 88
rect 103 87 104 88
rect 102 87 103 88
rect 101 87 102 88
rect 100 87 101 88
rect 99 87 100 88
rect 98 87 99 88
rect 97 87 98 88
rect 96 87 97 88
rect 95 87 96 88
rect 94 87 95 88
rect 93 87 94 88
rect 92 87 93 88
rect 91 87 92 88
rect 90 87 91 88
rect 89 87 90 88
rect 88 87 89 88
rect 87 87 88 88
rect 86 87 87 88
rect 85 87 86 88
rect 84 87 85 88
rect 83 87 84 88
rect 82 87 83 88
rect 81 87 82 88
rect 80 87 81 88
rect 79 87 80 88
rect 78 87 79 88
rect 77 87 78 88
rect 76 87 77 88
rect 75 87 76 88
rect 74 87 75 88
rect 73 87 74 88
rect 72 87 73 88
rect 71 87 72 88
rect 70 87 71 88
rect 69 87 70 88
rect 68 87 69 88
rect 67 87 68 88
rect 66 87 67 88
rect 65 87 66 88
rect 64 87 65 88
rect 63 87 64 88
rect 62 87 63 88
rect 61 87 62 88
rect 60 87 61 88
rect 59 87 60 88
rect 58 87 59 88
rect 479 88 480 89
rect 478 88 479 89
rect 477 88 478 89
rect 476 88 477 89
rect 458 88 459 89
rect 397 88 398 89
rect 396 88 397 89
rect 395 88 396 89
rect 394 88 395 89
rect 393 88 394 89
rect 246 88 247 89
rect 245 88 246 89
rect 244 88 245 89
rect 243 88 244 89
rect 242 88 243 89
rect 241 88 242 89
rect 240 88 241 89
rect 239 88 240 89
rect 238 88 239 89
rect 237 88 238 89
rect 236 88 237 89
rect 235 88 236 89
rect 234 88 235 89
rect 233 88 234 89
rect 232 88 233 89
rect 231 88 232 89
rect 230 88 231 89
rect 229 88 230 89
rect 228 88 229 89
rect 227 88 228 89
rect 226 88 227 89
rect 225 88 226 89
rect 224 88 225 89
rect 223 88 224 89
rect 222 88 223 89
rect 221 88 222 89
rect 220 88 221 89
rect 219 88 220 89
rect 218 88 219 89
rect 217 88 218 89
rect 216 88 217 89
rect 215 88 216 89
rect 214 88 215 89
rect 213 88 214 89
rect 212 88 213 89
rect 211 88 212 89
rect 210 88 211 89
rect 209 88 210 89
rect 208 88 209 89
rect 207 88 208 89
rect 206 88 207 89
rect 205 88 206 89
rect 204 88 205 89
rect 203 88 204 89
rect 202 88 203 89
rect 201 88 202 89
rect 200 88 201 89
rect 199 88 200 89
rect 198 88 199 89
rect 197 88 198 89
rect 196 88 197 89
rect 195 88 196 89
rect 194 88 195 89
rect 193 88 194 89
rect 192 88 193 89
rect 191 88 192 89
rect 190 88 191 89
rect 189 88 190 89
rect 188 88 189 89
rect 159 88 160 89
rect 158 88 159 89
rect 157 88 158 89
rect 156 88 157 89
rect 155 88 156 89
rect 154 88 155 89
rect 153 88 154 89
rect 152 88 153 89
rect 151 88 152 89
rect 150 88 151 89
rect 149 88 150 89
rect 148 88 149 89
rect 147 88 148 89
rect 146 88 147 89
rect 145 88 146 89
rect 144 88 145 89
rect 143 88 144 89
rect 142 88 143 89
rect 141 88 142 89
rect 140 88 141 89
rect 139 88 140 89
rect 138 88 139 89
rect 137 88 138 89
rect 136 88 137 89
rect 135 88 136 89
rect 134 88 135 89
rect 133 88 134 89
rect 132 88 133 89
rect 131 88 132 89
rect 130 88 131 89
rect 129 88 130 89
rect 128 88 129 89
rect 121 88 122 89
rect 120 88 121 89
rect 119 88 120 89
rect 118 88 119 89
rect 117 88 118 89
rect 116 88 117 89
rect 115 88 116 89
rect 114 88 115 89
rect 113 88 114 89
rect 112 88 113 89
rect 111 88 112 89
rect 110 88 111 89
rect 109 88 110 89
rect 108 88 109 89
rect 107 88 108 89
rect 106 88 107 89
rect 105 88 106 89
rect 104 88 105 89
rect 103 88 104 89
rect 102 88 103 89
rect 101 88 102 89
rect 100 88 101 89
rect 99 88 100 89
rect 98 88 99 89
rect 97 88 98 89
rect 96 88 97 89
rect 95 88 96 89
rect 94 88 95 89
rect 93 88 94 89
rect 92 88 93 89
rect 91 88 92 89
rect 90 88 91 89
rect 89 88 90 89
rect 88 88 89 89
rect 87 88 88 89
rect 86 88 87 89
rect 85 88 86 89
rect 84 88 85 89
rect 83 88 84 89
rect 82 88 83 89
rect 81 88 82 89
rect 80 88 81 89
rect 79 88 80 89
rect 78 88 79 89
rect 77 88 78 89
rect 76 88 77 89
rect 75 88 76 89
rect 74 88 75 89
rect 73 88 74 89
rect 72 88 73 89
rect 71 88 72 89
rect 70 88 71 89
rect 69 88 70 89
rect 68 88 69 89
rect 67 88 68 89
rect 66 88 67 89
rect 65 88 66 89
rect 64 88 65 89
rect 63 88 64 89
rect 62 88 63 89
rect 61 88 62 89
rect 60 88 61 89
rect 59 88 60 89
rect 58 88 59 89
rect 57 88 58 89
rect 479 89 480 90
rect 478 89 479 90
rect 477 89 478 90
rect 396 89 397 90
rect 395 89 396 90
rect 394 89 395 90
rect 393 89 394 90
rect 248 89 249 90
rect 247 89 248 90
rect 246 89 247 90
rect 245 89 246 90
rect 244 89 245 90
rect 243 89 244 90
rect 242 89 243 90
rect 241 89 242 90
rect 240 89 241 90
rect 239 89 240 90
rect 238 89 239 90
rect 237 89 238 90
rect 236 89 237 90
rect 235 89 236 90
rect 234 89 235 90
rect 233 89 234 90
rect 232 89 233 90
rect 231 89 232 90
rect 230 89 231 90
rect 229 89 230 90
rect 228 89 229 90
rect 227 89 228 90
rect 226 89 227 90
rect 225 89 226 90
rect 224 89 225 90
rect 223 89 224 90
rect 222 89 223 90
rect 221 89 222 90
rect 220 89 221 90
rect 219 89 220 90
rect 218 89 219 90
rect 217 89 218 90
rect 216 89 217 90
rect 215 89 216 90
rect 214 89 215 90
rect 213 89 214 90
rect 212 89 213 90
rect 211 89 212 90
rect 210 89 211 90
rect 209 89 210 90
rect 208 89 209 90
rect 207 89 208 90
rect 206 89 207 90
rect 205 89 206 90
rect 204 89 205 90
rect 203 89 204 90
rect 202 89 203 90
rect 201 89 202 90
rect 200 89 201 90
rect 199 89 200 90
rect 198 89 199 90
rect 197 89 198 90
rect 196 89 197 90
rect 195 89 196 90
rect 194 89 195 90
rect 193 89 194 90
rect 192 89 193 90
rect 191 89 192 90
rect 190 89 191 90
rect 189 89 190 90
rect 188 89 189 90
rect 187 89 188 90
rect 159 89 160 90
rect 158 89 159 90
rect 157 89 158 90
rect 156 89 157 90
rect 155 89 156 90
rect 154 89 155 90
rect 153 89 154 90
rect 152 89 153 90
rect 151 89 152 90
rect 150 89 151 90
rect 149 89 150 90
rect 148 89 149 90
rect 147 89 148 90
rect 146 89 147 90
rect 145 89 146 90
rect 144 89 145 90
rect 143 89 144 90
rect 142 89 143 90
rect 141 89 142 90
rect 140 89 141 90
rect 139 89 140 90
rect 138 89 139 90
rect 137 89 138 90
rect 136 89 137 90
rect 135 89 136 90
rect 134 89 135 90
rect 133 89 134 90
rect 132 89 133 90
rect 131 89 132 90
rect 130 89 131 90
rect 129 89 130 90
rect 128 89 129 90
rect 121 89 122 90
rect 120 89 121 90
rect 119 89 120 90
rect 118 89 119 90
rect 117 89 118 90
rect 116 89 117 90
rect 115 89 116 90
rect 114 89 115 90
rect 113 89 114 90
rect 112 89 113 90
rect 111 89 112 90
rect 110 89 111 90
rect 109 89 110 90
rect 108 89 109 90
rect 107 89 108 90
rect 106 89 107 90
rect 105 89 106 90
rect 104 89 105 90
rect 103 89 104 90
rect 102 89 103 90
rect 101 89 102 90
rect 100 89 101 90
rect 99 89 100 90
rect 98 89 99 90
rect 97 89 98 90
rect 96 89 97 90
rect 95 89 96 90
rect 94 89 95 90
rect 93 89 94 90
rect 92 89 93 90
rect 91 89 92 90
rect 90 89 91 90
rect 89 89 90 90
rect 88 89 89 90
rect 87 89 88 90
rect 86 89 87 90
rect 85 89 86 90
rect 84 89 85 90
rect 83 89 84 90
rect 82 89 83 90
rect 81 89 82 90
rect 80 89 81 90
rect 79 89 80 90
rect 78 89 79 90
rect 77 89 78 90
rect 76 89 77 90
rect 75 89 76 90
rect 74 89 75 90
rect 73 89 74 90
rect 72 89 73 90
rect 71 89 72 90
rect 70 89 71 90
rect 69 89 70 90
rect 68 89 69 90
rect 67 89 68 90
rect 66 89 67 90
rect 65 89 66 90
rect 64 89 65 90
rect 63 89 64 90
rect 62 89 63 90
rect 61 89 62 90
rect 60 89 61 90
rect 59 89 60 90
rect 58 89 59 90
rect 57 89 58 90
rect 56 89 57 90
rect 479 90 480 91
rect 478 90 479 91
rect 477 90 478 91
rect 396 90 397 91
rect 395 90 396 91
rect 394 90 395 91
rect 393 90 394 91
rect 250 90 251 91
rect 249 90 250 91
rect 248 90 249 91
rect 247 90 248 91
rect 246 90 247 91
rect 245 90 246 91
rect 244 90 245 91
rect 243 90 244 91
rect 242 90 243 91
rect 241 90 242 91
rect 240 90 241 91
rect 239 90 240 91
rect 238 90 239 91
rect 237 90 238 91
rect 236 90 237 91
rect 235 90 236 91
rect 234 90 235 91
rect 233 90 234 91
rect 232 90 233 91
rect 231 90 232 91
rect 230 90 231 91
rect 229 90 230 91
rect 228 90 229 91
rect 227 90 228 91
rect 226 90 227 91
rect 225 90 226 91
rect 224 90 225 91
rect 223 90 224 91
rect 222 90 223 91
rect 221 90 222 91
rect 220 90 221 91
rect 219 90 220 91
rect 218 90 219 91
rect 217 90 218 91
rect 216 90 217 91
rect 215 90 216 91
rect 214 90 215 91
rect 213 90 214 91
rect 212 90 213 91
rect 211 90 212 91
rect 210 90 211 91
rect 209 90 210 91
rect 208 90 209 91
rect 207 90 208 91
rect 206 90 207 91
rect 205 90 206 91
rect 204 90 205 91
rect 203 90 204 91
rect 202 90 203 91
rect 201 90 202 91
rect 200 90 201 91
rect 199 90 200 91
rect 198 90 199 91
rect 197 90 198 91
rect 196 90 197 91
rect 195 90 196 91
rect 194 90 195 91
rect 193 90 194 91
rect 192 90 193 91
rect 191 90 192 91
rect 190 90 191 91
rect 189 90 190 91
rect 188 90 189 91
rect 187 90 188 91
rect 186 90 187 91
rect 185 90 186 91
rect 159 90 160 91
rect 158 90 159 91
rect 157 90 158 91
rect 156 90 157 91
rect 155 90 156 91
rect 154 90 155 91
rect 153 90 154 91
rect 152 90 153 91
rect 151 90 152 91
rect 150 90 151 91
rect 149 90 150 91
rect 148 90 149 91
rect 147 90 148 91
rect 146 90 147 91
rect 145 90 146 91
rect 144 90 145 91
rect 143 90 144 91
rect 142 90 143 91
rect 141 90 142 91
rect 140 90 141 91
rect 139 90 140 91
rect 138 90 139 91
rect 137 90 138 91
rect 136 90 137 91
rect 135 90 136 91
rect 134 90 135 91
rect 133 90 134 91
rect 132 90 133 91
rect 131 90 132 91
rect 130 90 131 91
rect 129 90 130 91
rect 128 90 129 91
rect 120 90 121 91
rect 119 90 120 91
rect 118 90 119 91
rect 117 90 118 91
rect 116 90 117 91
rect 115 90 116 91
rect 114 90 115 91
rect 113 90 114 91
rect 112 90 113 91
rect 111 90 112 91
rect 110 90 111 91
rect 109 90 110 91
rect 108 90 109 91
rect 107 90 108 91
rect 106 90 107 91
rect 105 90 106 91
rect 104 90 105 91
rect 103 90 104 91
rect 102 90 103 91
rect 101 90 102 91
rect 100 90 101 91
rect 99 90 100 91
rect 98 90 99 91
rect 97 90 98 91
rect 96 90 97 91
rect 95 90 96 91
rect 94 90 95 91
rect 93 90 94 91
rect 92 90 93 91
rect 91 90 92 91
rect 90 90 91 91
rect 89 90 90 91
rect 88 90 89 91
rect 87 90 88 91
rect 86 90 87 91
rect 85 90 86 91
rect 84 90 85 91
rect 83 90 84 91
rect 82 90 83 91
rect 81 90 82 91
rect 80 90 81 91
rect 79 90 80 91
rect 78 90 79 91
rect 77 90 78 91
rect 76 90 77 91
rect 75 90 76 91
rect 74 90 75 91
rect 73 90 74 91
rect 72 90 73 91
rect 71 90 72 91
rect 70 90 71 91
rect 69 90 70 91
rect 68 90 69 91
rect 67 90 68 91
rect 66 90 67 91
rect 65 90 66 91
rect 64 90 65 91
rect 63 90 64 91
rect 62 90 63 91
rect 61 90 62 91
rect 60 90 61 91
rect 59 90 60 91
rect 58 90 59 91
rect 57 90 58 91
rect 56 90 57 91
rect 479 91 480 92
rect 478 91 479 92
rect 395 91 396 92
rect 394 91 395 92
rect 393 91 394 92
rect 252 91 253 92
rect 251 91 252 92
rect 250 91 251 92
rect 249 91 250 92
rect 248 91 249 92
rect 247 91 248 92
rect 246 91 247 92
rect 245 91 246 92
rect 244 91 245 92
rect 243 91 244 92
rect 242 91 243 92
rect 241 91 242 92
rect 240 91 241 92
rect 239 91 240 92
rect 238 91 239 92
rect 237 91 238 92
rect 236 91 237 92
rect 235 91 236 92
rect 234 91 235 92
rect 233 91 234 92
rect 232 91 233 92
rect 231 91 232 92
rect 230 91 231 92
rect 229 91 230 92
rect 228 91 229 92
rect 227 91 228 92
rect 226 91 227 92
rect 225 91 226 92
rect 224 91 225 92
rect 223 91 224 92
rect 222 91 223 92
rect 221 91 222 92
rect 220 91 221 92
rect 219 91 220 92
rect 218 91 219 92
rect 217 91 218 92
rect 216 91 217 92
rect 215 91 216 92
rect 214 91 215 92
rect 213 91 214 92
rect 212 91 213 92
rect 211 91 212 92
rect 210 91 211 92
rect 209 91 210 92
rect 208 91 209 92
rect 207 91 208 92
rect 206 91 207 92
rect 205 91 206 92
rect 204 91 205 92
rect 203 91 204 92
rect 202 91 203 92
rect 201 91 202 92
rect 200 91 201 92
rect 199 91 200 92
rect 198 91 199 92
rect 197 91 198 92
rect 196 91 197 92
rect 195 91 196 92
rect 194 91 195 92
rect 193 91 194 92
rect 192 91 193 92
rect 191 91 192 92
rect 190 91 191 92
rect 189 91 190 92
rect 188 91 189 92
rect 187 91 188 92
rect 186 91 187 92
rect 185 91 186 92
rect 184 91 185 92
rect 158 91 159 92
rect 157 91 158 92
rect 156 91 157 92
rect 155 91 156 92
rect 154 91 155 92
rect 153 91 154 92
rect 152 91 153 92
rect 151 91 152 92
rect 150 91 151 92
rect 149 91 150 92
rect 148 91 149 92
rect 147 91 148 92
rect 146 91 147 92
rect 145 91 146 92
rect 144 91 145 92
rect 143 91 144 92
rect 142 91 143 92
rect 141 91 142 92
rect 140 91 141 92
rect 139 91 140 92
rect 138 91 139 92
rect 137 91 138 92
rect 136 91 137 92
rect 135 91 136 92
rect 134 91 135 92
rect 133 91 134 92
rect 132 91 133 92
rect 131 91 132 92
rect 130 91 131 92
rect 129 91 130 92
rect 128 91 129 92
rect 127 91 128 92
rect 120 91 121 92
rect 119 91 120 92
rect 118 91 119 92
rect 117 91 118 92
rect 116 91 117 92
rect 115 91 116 92
rect 114 91 115 92
rect 113 91 114 92
rect 112 91 113 92
rect 111 91 112 92
rect 110 91 111 92
rect 109 91 110 92
rect 108 91 109 92
rect 107 91 108 92
rect 106 91 107 92
rect 105 91 106 92
rect 104 91 105 92
rect 103 91 104 92
rect 102 91 103 92
rect 101 91 102 92
rect 100 91 101 92
rect 99 91 100 92
rect 98 91 99 92
rect 97 91 98 92
rect 96 91 97 92
rect 95 91 96 92
rect 94 91 95 92
rect 93 91 94 92
rect 92 91 93 92
rect 91 91 92 92
rect 90 91 91 92
rect 89 91 90 92
rect 88 91 89 92
rect 87 91 88 92
rect 86 91 87 92
rect 85 91 86 92
rect 84 91 85 92
rect 83 91 84 92
rect 82 91 83 92
rect 81 91 82 92
rect 80 91 81 92
rect 79 91 80 92
rect 78 91 79 92
rect 77 91 78 92
rect 76 91 77 92
rect 75 91 76 92
rect 74 91 75 92
rect 73 91 74 92
rect 72 91 73 92
rect 71 91 72 92
rect 70 91 71 92
rect 69 91 70 92
rect 68 91 69 92
rect 67 91 68 92
rect 66 91 67 92
rect 65 91 66 92
rect 64 91 65 92
rect 63 91 64 92
rect 62 91 63 92
rect 61 91 62 92
rect 60 91 61 92
rect 59 91 60 92
rect 58 91 59 92
rect 57 91 58 92
rect 56 91 57 92
rect 55 91 56 92
rect 479 92 480 93
rect 478 92 479 93
rect 395 92 396 93
rect 394 92 395 93
rect 393 92 394 93
rect 253 92 254 93
rect 252 92 253 93
rect 251 92 252 93
rect 250 92 251 93
rect 249 92 250 93
rect 248 92 249 93
rect 247 92 248 93
rect 246 92 247 93
rect 245 92 246 93
rect 244 92 245 93
rect 243 92 244 93
rect 242 92 243 93
rect 241 92 242 93
rect 240 92 241 93
rect 239 92 240 93
rect 238 92 239 93
rect 237 92 238 93
rect 236 92 237 93
rect 235 92 236 93
rect 234 92 235 93
rect 233 92 234 93
rect 232 92 233 93
rect 231 92 232 93
rect 230 92 231 93
rect 229 92 230 93
rect 228 92 229 93
rect 227 92 228 93
rect 226 92 227 93
rect 225 92 226 93
rect 224 92 225 93
rect 223 92 224 93
rect 222 92 223 93
rect 221 92 222 93
rect 220 92 221 93
rect 219 92 220 93
rect 218 92 219 93
rect 217 92 218 93
rect 216 92 217 93
rect 215 92 216 93
rect 214 92 215 93
rect 213 92 214 93
rect 212 92 213 93
rect 211 92 212 93
rect 210 92 211 93
rect 209 92 210 93
rect 208 92 209 93
rect 207 92 208 93
rect 206 92 207 93
rect 205 92 206 93
rect 204 92 205 93
rect 203 92 204 93
rect 202 92 203 93
rect 201 92 202 93
rect 200 92 201 93
rect 199 92 200 93
rect 198 92 199 93
rect 197 92 198 93
rect 196 92 197 93
rect 195 92 196 93
rect 194 92 195 93
rect 193 92 194 93
rect 192 92 193 93
rect 191 92 192 93
rect 190 92 191 93
rect 189 92 190 93
rect 188 92 189 93
rect 187 92 188 93
rect 186 92 187 93
rect 185 92 186 93
rect 184 92 185 93
rect 183 92 184 93
rect 158 92 159 93
rect 157 92 158 93
rect 156 92 157 93
rect 155 92 156 93
rect 154 92 155 93
rect 153 92 154 93
rect 152 92 153 93
rect 151 92 152 93
rect 150 92 151 93
rect 149 92 150 93
rect 148 92 149 93
rect 147 92 148 93
rect 146 92 147 93
rect 145 92 146 93
rect 144 92 145 93
rect 143 92 144 93
rect 142 92 143 93
rect 141 92 142 93
rect 140 92 141 93
rect 139 92 140 93
rect 138 92 139 93
rect 137 92 138 93
rect 136 92 137 93
rect 135 92 136 93
rect 134 92 135 93
rect 133 92 134 93
rect 132 92 133 93
rect 131 92 132 93
rect 130 92 131 93
rect 129 92 130 93
rect 128 92 129 93
rect 127 92 128 93
rect 120 92 121 93
rect 119 92 120 93
rect 118 92 119 93
rect 117 92 118 93
rect 116 92 117 93
rect 115 92 116 93
rect 114 92 115 93
rect 113 92 114 93
rect 112 92 113 93
rect 111 92 112 93
rect 110 92 111 93
rect 109 92 110 93
rect 108 92 109 93
rect 107 92 108 93
rect 106 92 107 93
rect 105 92 106 93
rect 104 92 105 93
rect 103 92 104 93
rect 102 92 103 93
rect 101 92 102 93
rect 100 92 101 93
rect 99 92 100 93
rect 98 92 99 93
rect 97 92 98 93
rect 96 92 97 93
rect 95 92 96 93
rect 94 92 95 93
rect 93 92 94 93
rect 92 92 93 93
rect 91 92 92 93
rect 90 92 91 93
rect 89 92 90 93
rect 88 92 89 93
rect 87 92 88 93
rect 86 92 87 93
rect 85 92 86 93
rect 84 92 85 93
rect 83 92 84 93
rect 82 92 83 93
rect 81 92 82 93
rect 80 92 81 93
rect 79 92 80 93
rect 78 92 79 93
rect 77 92 78 93
rect 76 92 77 93
rect 75 92 76 93
rect 74 92 75 93
rect 73 92 74 93
rect 72 92 73 93
rect 71 92 72 93
rect 70 92 71 93
rect 69 92 70 93
rect 68 92 69 93
rect 67 92 68 93
rect 66 92 67 93
rect 65 92 66 93
rect 64 92 65 93
rect 63 92 64 93
rect 62 92 63 93
rect 61 92 62 93
rect 60 92 61 93
rect 59 92 60 93
rect 58 92 59 93
rect 57 92 58 93
rect 56 92 57 93
rect 55 92 56 93
rect 54 92 55 93
rect 479 93 480 94
rect 478 93 479 94
rect 477 93 478 94
rect 395 93 396 94
rect 394 93 395 94
rect 393 93 394 94
rect 255 93 256 94
rect 254 93 255 94
rect 253 93 254 94
rect 252 93 253 94
rect 251 93 252 94
rect 250 93 251 94
rect 249 93 250 94
rect 248 93 249 94
rect 247 93 248 94
rect 246 93 247 94
rect 245 93 246 94
rect 244 93 245 94
rect 243 93 244 94
rect 242 93 243 94
rect 241 93 242 94
rect 240 93 241 94
rect 239 93 240 94
rect 238 93 239 94
rect 237 93 238 94
rect 236 93 237 94
rect 235 93 236 94
rect 234 93 235 94
rect 233 93 234 94
rect 232 93 233 94
rect 231 93 232 94
rect 230 93 231 94
rect 229 93 230 94
rect 228 93 229 94
rect 227 93 228 94
rect 226 93 227 94
rect 225 93 226 94
rect 224 93 225 94
rect 223 93 224 94
rect 222 93 223 94
rect 221 93 222 94
rect 220 93 221 94
rect 219 93 220 94
rect 218 93 219 94
rect 217 93 218 94
rect 216 93 217 94
rect 215 93 216 94
rect 214 93 215 94
rect 213 93 214 94
rect 212 93 213 94
rect 211 93 212 94
rect 210 93 211 94
rect 209 93 210 94
rect 208 93 209 94
rect 207 93 208 94
rect 206 93 207 94
rect 205 93 206 94
rect 204 93 205 94
rect 203 93 204 94
rect 202 93 203 94
rect 201 93 202 94
rect 200 93 201 94
rect 199 93 200 94
rect 198 93 199 94
rect 197 93 198 94
rect 196 93 197 94
rect 195 93 196 94
rect 194 93 195 94
rect 193 93 194 94
rect 192 93 193 94
rect 191 93 192 94
rect 190 93 191 94
rect 189 93 190 94
rect 188 93 189 94
rect 187 93 188 94
rect 186 93 187 94
rect 185 93 186 94
rect 184 93 185 94
rect 183 93 184 94
rect 182 93 183 94
rect 158 93 159 94
rect 157 93 158 94
rect 156 93 157 94
rect 155 93 156 94
rect 154 93 155 94
rect 153 93 154 94
rect 152 93 153 94
rect 151 93 152 94
rect 150 93 151 94
rect 149 93 150 94
rect 148 93 149 94
rect 147 93 148 94
rect 146 93 147 94
rect 145 93 146 94
rect 144 93 145 94
rect 143 93 144 94
rect 142 93 143 94
rect 141 93 142 94
rect 140 93 141 94
rect 139 93 140 94
rect 138 93 139 94
rect 137 93 138 94
rect 136 93 137 94
rect 135 93 136 94
rect 134 93 135 94
rect 133 93 134 94
rect 132 93 133 94
rect 131 93 132 94
rect 130 93 131 94
rect 129 93 130 94
rect 128 93 129 94
rect 127 93 128 94
rect 120 93 121 94
rect 119 93 120 94
rect 118 93 119 94
rect 117 93 118 94
rect 116 93 117 94
rect 115 93 116 94
rect 114 93 115 94
rect 113 93 114 94
rect 112 93 113 94
rect 111 93 112 94
rect 110 93 111 94
rect 109 93 110 94
rect 108 93 109 94
rect 107 93 108 94
rect 106 93 107 94
rect 105 93 106 94
rect 104 93 105 94
rect 103 93 104 94
rect 102 93 103 94
rect 101 93 102 94
rect 100 93 101 94
rect 99 93 100 94
rect 98 93 99 94
rect 97 93 98 94
rect 96 93 97 94
rect 95 93 96 94
rect 94 93 95 94
rect 93 93 94 94
rect 92 93 93 94
rect 91 93 92 94
rect 90 93 91 94
rect 89 93 90 94
rect 88 93 89 94
rect 87 93 88 94
rect 86 93 87 94
rect 85 93 86 94
rect 84 93 85 94
rect 83 93 84 94
rect 82 93 83 94
rect 81 93 82 94
rect 80 93 81 94
rect 79 93 80 94
rect 78 93 79 94
rect 77 93 78 94
rect 76 93 77 94
rect 75 93 76 94
rect 74 93 75 94
rect 73 93 74 94
rect 72 93 73 94
rect 71 93 72 94
rect 70 93 71 94
rect 69 93 70 94
rect 68 93 69 94
rect 67 93 68 94
rect 66 93 67 94
rect 65 93 66 94
rect 64 93 65 94
rect 63 93 64 94
rect 62 93 63 94
rect 61 93 62 94
rect 60 93 61 94
rect 59 93 60 94
rect 58 93 59 94
rect 57 93 58 94
rect 56 93 57 94
rect 55 93 56 94
rect 54 93 55 94
rect 53 93 54 94
rect 478 94 479 95
rect 477 94 478 95
rect 458 94 459 95
rect 257 94 258 95
rect 256 94 257 95
rect 255 94 256 95
rect 254 94 255 95
rect 253 94 254 95
rect 252 94 253 95
rect 251 94 252 95
rect 250 94 251 95
rect 249 94 250 95
rect 248 94 249 95
rect 247 94 248 95
rect 246 94 247 95
rect 245 94 246 95
rect 244 94 245 95
rect 243 94 244 95
rect 242 94 243 95
rect 241 94 242 95
rect 240 94 241 95
rect 239 94 240 95
rect 238 94 239 95
rect 237 94 238 95
rect 236 94 237 95
rect 235 94 236 95
rect 234 94 235 95
rect 233 94 234 95
rect 232 94 233 95
rect 231 94 232 95
rect 230 94 231 95
rect 229 94 230 95
rect 228 94 229 95
rect 227 94 228 95
rect 226 94 227 95
rect 225 94 226 95
rect 224 94 225 95
rect 223 94 224 95
rect 222 94 223 95
rect 221 94 222 95
rect 220 94 221 95
rect 219 94 220 95
rect 218 94 219 95
rect 217 94 218 95
rect 216 94 217 95
rect 215 94 216 95
rect 214 94 215 95
rect 213 94 214 95
rect 212 94 213 95
rect 211 94 212 95
rect 210 94 211 95
rect 209 94 210 95
rect 208 94 209 95
rect 207 94 208 95
rect 206 94 207 95
rect 205 94 206 95
rect 204 94 205 95
rect 203 94 204 95
rect 202 94 203 95
rect 201 94 202 95
rect 200 94 201 95
rect 199 94 200 95
rect 198 94 199 95
rect 197 94 198 95
rect 196 94 197 95
rect 195 94 196 95
rect 194 94 195 95
rect 193 94 194 95
rect 192 94 193 95
rect 191 94 192 95
rect 190 94 191 95
rect 189 94 190 95
rect 188 94 189 95
rect 187 94 188 95
rect 186 94 187 95
rect 185 94 186 95
rect 184 94 185 95
rect 183 94 184 95
rect 182 94 183 95
rect 181 94 182 95
rect 157 94 158 95
rect 156 94 157 95
rect 155 94 156 95
rect 154 94 155 95
rect 153 94 154 95
rect 152 94 153 95
rect 151 94 152 95
rect 150 94 151 95
rect 149 94 150 95
rect 148 94 149 95
rect 147 94 148 95
rect 146 94 147 95
rect 145 94 146 95
rect 144 94 145 95
rect 143 94 144 95
rect 142 94 143 95
rect 141 94 142 95
rect 140 94 141 95
rect 139 94 140 95
rect 138 94 139 95
rect 137 94 138 95
rect 136 94 137 95
rect 135 94 136 95
rect 134 94 135 95
rect 133 94 134 95
rect 132 94 133 95
rect 131 94 132 95
rect 130 94 131 95
rect 129 94 130 95
rect 128 94 129 95
rect 127 94 128 95
rect 119 94 120 95
rect 118 94 119 95
rect 117 94 118 95
rect 116 94 117 95
rect 115 94 116 95
rect 114 94 115 95
rect 113 94 114 95
rect 112 94 113 95
rect 111 94 112 95
rect 110 94 111 95
rect 109 94 110 95
rect 108 94 109 95
rect 107 94 108 95
rect 106 94 107 95
rect 105 94 106 95
rect 104 94 105 95
rect 103 94 104 95
rect 102 94 103 95
rect 101 94 102 95
rect 100 94 101 95
rect 99 94 100 95
rect 98 94 99 95
rect 97 94 98 95
rect 96 94 97 95
rect 95 94 96 95
rect 94 94 95 95
rect 93 94 94 95
rect 92 94 93 95
rect 91 94 92 95
rect 90 94 91 95
rect 89 94 90 95
rect 88 94 89 95
rect 87 94 88 95
rect 86 94 87 95
rect 85 94 86 95
rect 84 94 85 95
rect 83 94 84 95
rect 82 94 83 95
rect 81 94 82 95
rect 80 94 81 95
rect 79 94 80 95
rect 78 94 79 95
rect 77 94 78 95
rect 76 94 77 95
rect 75 94 76 95
rect 74 94 75 95
rect 73 94 74 95
rect 72 94 73 95
rect 71 94 72 95
rect 70 94 71 95
rect 69 94 70 95
rect 68 94 69 95
rect 67 94 68 95
rect 66 94 67 95
rect 65 94 66 95
rect 64 94 65 95
rect 63 94 64 95
rect 62 94 63 95
rect 61 94 62 95
rect 60 94 61 95
rect 59 94 60 95
rect 58 94 59 95
rect 57 94 58 95
rect 56 94 57 95
rect 55 94 56 95
rect 54 94 55 95
rect 53 94 54 95
rect 52 94 53 95
rect 478 95 479 96
rect 477 95 478 96
rect 476 95 477 96
rect 458 95 459 96
rect 258 95 259 96
rect 257 95 258 96
rect 256 95 257 96
rect 255 95 256 96
rect 254 95 255 96
rect 253 95 254 96
rect 252 95 253 96
rect 251 95 252 96
rect 250 95 251 96
rect 249 95 250 96
rect 248 95 249 96
rect 247 95 248 96
rect 246 95 247 96
rect 245 95 246 96
rect 244 95 245 96
rect 243 95 244 96
rect 242 95 243 96
rect 241 95 242 96
rect 240 95 241 96
rect 239 95 240 96
rect 238 95 239 96
rect 237 95 238 96
rect 236 95 237 96
rect 235 95 236 96
rect 234 95 235 96
rect 233 95 234 96
rect 232 95 233 96
rect 231 95 232 96
rect 230 95 231 96
rect 229 95 230 96
rect 228 95 229 96
rect 227 95 228 96
rect 226 95 227 96
rect 225 95 226 96
rect 224 95 225 96
rect 223 95 224 96
rect 222 95 223 96
rect 221 95 222 96
rect 220 95 221 96
rect 219 95 220 96
rect 218 95 219 96
rect 217 95 218 96
rect 216 95 217 96
rect 215 95 216 96
rect 214 95 215 96
rect 213 95 214 96
rect 212 95 213 96
rect 211 95 212 96
rect 210 95 211 96
rect 209 95 210 96
rect 208 95 209 96
rect 207 95 208 96
rect 206 95 207 96
rect 205 95 206 96
rect 204 95 205 96
rect 203 95 204 96
rect 202 95 203 96
rect 201 95 202 96
rect 200 95 201 96
rect 199 95 200 96
rect 198 95 199 96
rect 197 95 198 96
rect 196 95 197 96
rect 195 95 196 96
rect 194 95 195 96
rect 193 95 194 96
rect 192 95 193 96
rect 191 95 192 96
rect 190 95 191 96
rect 189 95 190 96
rect 188 95 189 96
rect 187 95 188 96
rect 186 95 187 96
rect 185 95 186 96
rect 184 95 185 96
rect 183 95 184 96
rect 182 95 183 96
rect 181 95 182 96
rect 180 95 181 96
rect 157 95 158 96
rect 156 95 157 96
rect 155 95 156 96
rect 154 95 155 96
rect 153 95 154 96
rect 152 95 153 96
rect 151 95 152 96
rect 150 95 151 96
rect 149 95 150 96
rect 148 95 149 96
rect 147 95 148 96
rect 146 95 147 96
rect 145 95 146 96
rect 144 95 145 96
rect 143 95 144 96
rect 142 95 143 96
rect 141 95 142 96
rect 140 95 141 96
rect 139 95 140 96
rect 138 95 139 96
rect 137 95 138 96
rect 136 95 137 96
rect 135 95 136 96
rect 134 95 135 96
rect 133 95 134 96
rect 132 95 133 96
rect 131 95 132 96
rect 130 95 131 96
rect 129 95 130 96
rect 128 95 129 96
rect 127 95 128 96
rect 119 95 120 96
rect 118 95 119 96
rect 117 95 118 96
rect 116 95 117 96
rect 115 95 116 96
rect 114 95 115 96
rect 113 95 114 96
rect 112 95 113 96
rect 111 95 112 96
rect 110 95 111 96
rect 109 95 110 96
rect 108 95 109 96
rect 107 95 108 96
rect 106 95 107 96
rect 105 95 106 96
rect 104 95 105 96
rect 103 95 104 96
rect 102 95 103 96
rect 101 95 102 96
rect 100 95 101 96
rect 99 95 100 96
rect 98 95 99 96
rect 97 95 98 96
rect 96 95 97 96
rect 95 95 96 96
rect 94 95 95 96
rect 93 95 94 96
rect 92 95 93 96
rect 91 95 92 96
rect 90 95 91 96
rect 89 95 90 96
rect 88 95 89 96
rect 87 95 88 96
rect 86 95 87 96
rect 85 95 86 96
rect 84 95 85 96
rect 83 95 84 96
rect 82 95 83 96
rect 81 95 82 96
rect 80 95 81 96
rect 79 95 80 96
rect 78 95 79 96
rect 77 95 78 96
rect 76 95 77 96
rect 75 95 76 96
rect 74 95 75 96
rect 73 95 74 96
rect 70 95 71 96
rect 69 95 70 96
rect 68 95 69 96
rect 67 95 68 96
rect 66 95 67 96
rect 65 95 66 96
rect 64 95 65 96
rect 63 95 64 96
rect 62 95 63 96
rect 61 95 62 96
rect 60 95 61 96
rect 59 95 60 96
rect 58 95 59 96
rect 57 95 58 96
rect 56 95 57 96
rect 55 95 56 96
rect 54 95 55 96
rect 53 95 54 96
rect 52 95 53 96
rect 51 95 52 96
rect 477 96 478 97
rect 476 96 477 97
rect 475 96 476 97
rect 459 96 460 97
rect 458 96 459 97
rect 260 96 261 97
rect 259 96 260 97
rect 258 96 259 97
rect 257 96 258 97
rect 256 96 257 97
rect 255 96 256 97
rect 254 96 255 97
rect 253 96 254 97
rect 252 96 253 97
rect 251 96 252 97
rect 250 96 251 97
rect 249 96 250 97
rect 248 96 249 97
rect 247 96 248 97
rect 246 96 247 97
rect 245 96 246 97
rect 244 96 245 97
rect 243 96 244 97
rect 242 96 243 97
rect 241 96 242 97
rect 240 96 241 97
rect 239 96 240 97
rect 238 96 239 97
rect 237 96 238 97
rect 236 96 237 97
rect 235 96 236 97
rect 234 96 235 97
rect 233 96 234 97
rect 232 96 233 97
rect 231 96 232 97
rect 230 96 231 97
rect 229 96 230 97
rect 228 96 229 97
rect 227 96 228 97
rect 226 96 227 97
rect 225 96 226 97
rect 224 96 225 97
rect 223 96 224 97
rect 222 96 223 97
rect 221 96 222 97
rect 220 96 221 97
rect 219 96 220 97
rect 218 96 219 97
rect 217 96 218 97
rect 216 96 217 97
rect 215 96 216 97
rect 214 96 215 97
rect 213 96 214 97
rect 212 96 213 97
rect 211 96 212 97
rect 210 96 211 97
rect 209 96 210 97
rect 208 96 209 97
rect 207 96 208 97
rect 206 96 207 97
rect 205 96 206 97
rect 204 96 205 97
rect 203 96 204 97
rect 202 96 203 97
rect 201 96 202 97
rect 200 96 201 97
rect 199 96 200 97
rect 198 96 199 97
rect 197 96 198 97
rect 196 96 197 97
rect 195 96 196 97
rect 194 96 195 97
rect 193 96 194 97
rect 192 96 193 97
rect 191 96 192 97
rect 190 96 191 97
rect 189 96 190 97
rect 188 96 189 97
rect 187 96 188 97
rect 186 96 187 97
rect 185 96 186 97
rect 184 96 185 97
rect 183 96 184 97
rect 182 96 183 97
rect 181 96 182 97
rect 180 96 181 97
rect 179 96 180 97
rect 157 96 158 97
rect 156 96 157 97
rect 155 96 156 97
rect 154 96 155 97
rect 153 96 154 97
rect 152 96 153 97
rect 151 96 152 97
rect 150 96 151 97
rect 149 96 150 97
rect 148 96 149 97
rect 147 96 148 97
rect 146 96 147 97
rect 145 96 146 97
rect 144 96 145 97
rect 143 96 144 97
rect 142 96 143 97
rect 141 96 142 97
rect 140 96 141 97
rect 139 96 140 97
rect 138 96 139 97
rect 137 96 138 97
rect 136 96 137 97
rect 135 96 136 97
rect 134 96 135 97
rect 133 96 134 97
rect 132 96 133 97
rect 131 96 132 97
rect 130 96 131 97
rect 129 96 130 97
rect 128 96 129 97
rect 127 96 128 97
rect 119 96 120 97
rect 118 96 119 97
rect 117 96 118 97
rect 116 96 117 97
rect 115 96 116 97
rect 114 96 115 97
rect 113 96 114 97
rect 112 96 113 97
rect 111 96 112 97
rect 110 96 111 97
rect 109 96 110 97
rect 108 96 109 97
rect 107 96 108 97
rect 106 96 107 97
rect 105 96 106 97
rect 104 96 105 97
rect 103 96 104 97
rect 102 96 103 97
rect 101 96 102 97
rect 100 96 101 97
rect 99 96 100 97
rect 98 96 99 97
rect 97 96 98 97
rect 96 96 97 97
rect 95 96 96 97
rect 94 96 95 97
rect 93 96 94 97
rect 92 96 93 97
rect 91 96 92 97
rect 90 96 91 97
rect 89 96 90 97
rect 88 96 89 97
rect 87 96 88 97
rect 86 96 87 97
rect 85 96 86 97
rect 84 96 85 97
rect 83 96 84 97
rect 82 96 83 97
rect 81 96 82 97
rect 80 96 81 97
rect 79 96 80 97
rect 78 96 79 97
rect 77 96 78 97
rect 76 96 77 97
rect 75 96 76 97
rect 74 96 75 97
rect 73 96 74 97
rect 69 96 70 97
rect 68 96 69 97
rect 67 96 68 97
rect 66 96 67 97
rect 65 96 66 97
rect 64 96 65 97
rect 63 96 64 97
rect 62 96 63 97
rect 61 96 62 97
rect 60 96 61 97
rect 59 96 60 97
rect 58 96 59 97
rect 57 96 58 97
rect 56 96 57 97
rect 55 96 56 97
rect 54 96 55 97
rect 53 96 54 97
rect 52 96 53 97
rect 51 96 52 97
rect 50 96 51 97
rect 476 97 477 98
rect 475 97 476 98
rect 474 97 475 98
rect 473 97 474 98
rect 472 97 473 98
rect 471 97 472 98
rect 470 97 471 98
rect 469 97 470 98
rect 468 97 469 98
rect 467 97 468 98
rect 466 97 467 98
rect 465 97 466 98
rect 464 97 465 98
rect 463 97 464 98
rect 462 97 463 98
rect 461 97 462 98
rect 460 97 461 98
rect 459 97 460 98
rect 458 97 459 98
rect 261 97 262 98
rect 260 97 261 98
rect 259 97 260 98
rect 258 97 259 98
rect 257 97 258 98
rect 256 97 257 98
rect 255 97 256 98
rect 254 97 255 98
rect 253 97 254 98
rect 252 97 253 98
rect 251 97 252 98
rect 250 97 251 98
rect 249 97 250 98
rect 248 97 249 98
rect 247 97 248 98
rect 246 97 247 98
rect 245 97 246 98
rect 244 97 245 98
rect 243 97 244 98
rect 242 97 243 98
rect 241 97 242 98
rect 240 97 241 98
rect 239 97 240 98
rect 238 97 239 98
rect 237 97 238 98
rect 236 97 237 98
rect 235 97 236 98
rect 234 97 235 98
rect 233 97 234 98
rect 232 97 233 98
rect 231 97 232 98
rect 230 97 231 98
rect 229 97 230 98
rect 228 97 229 98
rect 227 97 228 98
rect 226 97 227 98
rect 225 97 226 98
rect 224 97 225 98
rect 223 97 224 98
rect 222 97 223 98
rect 221 97 222 98
rect 220 97 221 98
rect 219 97 220 98
rect 218 97 219 98
rect 217 97 218 98
rect 216 97 217 98
rect 215 97 216 98
rect 214 97 215 98
rect 213 97 214 98
rect 212 97 213 98
rect 211 97 212 98
rect 210 97 211 98
rect 209 97 210 98
rect 208 97 209 98
rect 207 97 208 98
rect 206 97 207 98
rect 205 97 206 98
rect 204 97 205 98
rect 203 97 204 98
rect 202 97 203 98
rect 201 97 202 98
rect 200 97 201 98
rect 199 97 200 98
rect 198 97 199 98
rect 197 97 198 98
rect 196 97 197 98
rect 195 97 196 98
rect 194 97 195 98
rect 193 97 194 98
rect 192 97 193 98
rect 191 97 192 98
rect 190 97 191 98
rect 189 97 190 98
rect 188 97 189 98
rect 187 97 188 98
rect 186 97 187 98
rect 185 97 186 98
rect 184 97 185 98
rect 183 97 184 98
rect 182 97 183 98
rect 181 97 182 98
rect 180 97 181 98
rect 179 97 180 98
rect 178 97 179 98
rect 156 97 157 98
rect 155 97 156 98
rect 154 97 155 98
rect 153 97 154 98
rect 152 97 153 98
rect 151 97 152 98
rect 150 97 151 98
rect 149 97 150 98
rect 148 97 149 98
rect 147 97 148 98
rect 146 97 147 98
rect 145 97 146 98
rect 144 97 145 98
rect 143 97 144 98
rect 142 97 143 98
rect 141 97 142 98
rect 140 97 141 98
rect 139 97 140 98
rect 138 97 139 98
rect 137 97 138 98
rect 136 97 137 98
rect 135 97 136 98
rect 134 97 135 98
rect 133 97 134 98
rect 132 97 133 98
rect 131 97 132 98
rect 130 97 131 98
rect 129 97 130 98
rect 128 97 129 98
rect 127 97 128 98
rect 126 97 127 98
rect 118 97 119 98
rect 117 97 118 98
rect 116 97 117 98
rect 115 97 116 98
rect 114 97 115 98
rect 113 97 114 98
rect 112 97 113 98
rect 111 97 112 98
rect 110 97 111 98
rect 109 97 110 98
rect 108 97 109 98
rect 107 97 108 98
rect 106 97 107 98
rect 105 97 106 98
rect 104 97 105 98
rect 103 97 104 98
rect 102 97 103 98
rect 101 97 102 98
rect 100 97 101 98
rect 99 97 100 98
rect 98 97 99 98
rect 97 97 98 98
rect 96 97 97 98
rect 95 97 96 98
rect 94 97 95 98
rect 93 97 94 98
rect 92 97 93 98
rect 91 97 92 98
rect 90 97 91 98
rect 89 97 90 98
rect 88 97 89 98
rect 87 97 88 98
rect 86 97 87 98
rect 85 97 86 98
rect 84 97 85 98
rect 83 97 84 98
rect 82 97 83 98
rect 81 97 82 98
rect 80 97 81 98
rect 79 97 80 98
rect 78 97 79 98
rect 77 97 78 98
rect 76 97 77 98
rect 75 97 76 98
rect 74 97 75 98
rect 73 97 74 98
rect 72 97 73 98
rect 68 97 69 98
rect 67 97 68 98
rect 66 97 67 98
rect 65 97 66 98
rect 64 97 65 98
rect 63 97 64 98
rect 62 97 63 98
rect 61 97 62 98
rect 60 97 61 98
rect 59 97 60 98
rect 58 97 59 98
rect 57 97 58 98
rect 56 97 57 98
rect 55 97 56 98
rect 54 97 55 98
rect 53 97 54 98
rect 52 97 53 98
rect 51 97 52 98
rect 50 97 51 98
rect 49 97 50 98
rect 474 98 475 99
rect 473 98 474 99
rect 472 98 473 99
rect 471 98 472 99
rect 470 98 471 99
rect 469 98 470 99
rect 468 98 469 99
rect 467 98 468 99
rect 466 98 467 99
rect 465 98 466 99
rect 464 98 465 99
rect 463 98 464 99
rect 462 98 463 99
rect 461 98 462 99
rect 460 98 461 99
rect 459 98 460 99
rect 458 98 459 99
rect 262 98 263 99
rect 261 98 262 99
rect 260 98 261 99
rect 259 98 260 99
rect 258 98 259 99
rect 257 98 258 99
rect 256 98 257 99
rect 255 98 256 99
rect 254 98 255 99
rect 253 98 254 99
rect 252 98 253 99
rect 251 98 252 99
rect 250 98 251 99
rect 249 98 250 99
rect 248 98 249 99
rect 247 98 248 99
rect 246 98 247 99
rect 245 98 246 99
rect 244 98 245 99
rect 243 98 244 99
rect 242 98 243 99
rect 241 98 242 99
rect 240 98 241 99
rect 239 98 240 99
rect 238 98 239 99
rect 237 98 238 99
rect 236 98 237 99
rect 235 98 236 99
rect 234 98 235 99
rect 233 98 234 99
rect 232 98 233 99
rect 231 98 232 99
rect 230 98 231 99
rect 229 98 230 99
rect 228 98 229 99
rect 227 98 228 99
rect 226 98 227 99
rect 225 98 226 99
rect 224 98 225 99
rect 223 98 224 99
rect 222 98 223 99
rect 221 98 222 99
rect 220 98 221 99
rect 219 98 220 99
rect 218 98 219 99
rect 217 98 218 99
rect 216 98 217 99
rect 215 98 216 99
rect 214 98 215 99
rect 213 98 214 99
rect 212 98 213 99
rect 211 98 212 99
rect 210 98 211 99
rect 209 98 210 99
rect 208 98 209 99
rect 207 98 208 99
rect 206 98 207 99
rect 205 98 206 99
rect 204 98 205 99
rect 203 98 204 99
rect 202 98 203 99
rect 201 98 202 99
rect 200 98 201 99
rect 199 98 200 99
rect 198 98 199 99
rect 197 98 198 99
rect 196 98 197 99
rect 195 98 196 99
rect 194 98 195 99
rect 193 98 194 99
rect 192 98 193 99
rect 191 98 192 99
rect 190 98 191 99
rect 189 98 190 99
rect 188 98 189 99
rect 187 98 188 99
rect 186 98 187 99
rect 185 98 186 99
rect 184 98 185 99
rect 183 98 184 99
rect 182 98 183 99
rect 181 98 182 99
rect 180 98 181 99
rect 179 98 180 99
rect 178 98 179 99
rect 177 98 178 99
rect 156 98 157 99
rect 155 98 156 99
rect 154 98 155 99
rect 153 98 154 99
rect 152 98 153 99
rect 151 98 152 99
rect 150 98 151 99
rect 149 98 150 99
rect 148 98 149 99
rect 147 98 148 99
rect 146 98 147 99
rect 145 98 146 99
rect 144 98 145 99
rect 143 98 144 99
rect 142 98 143 99
rect 141 98 142 99
rect 140 98 141 99
rect 139 98 140 99
rect 138 98 139 99
rect 137 98 138 99
rect 136 98 137 99
rect 135 98 136 99
rect 134 98 135 99
rect 133 98 134 99
rect 132 98 133 99
rect 131 98 132 99
rect 130 98 131 99
rect 129 98 130 99
rect 128 98 129 99
rect 127 98 128 99
rect 126 98 127 99
rect 117 98 118 99
rect 116 98 117 99
rect 115 98 116 99
rect 114 98 115 99
rect 113 98 114 99
rect 112 98 113 99
rect 111 98 112 99
rect 110 98 111 99
rect 109 98 110 99
rect 108 98 109 99
rect 107 98 108 99
rect 106 98 107 99
rect 105 98 106 99
rect 104 98 105 99
rect 103 98 104 99
rect 102 98 103 99
rect 101 98 102 99
rect 100 98 101 99
rect 99 98 100 99
rect 98 98 99 99
rect 97 98 98 99
rect 96 98 97 99
rect 95 98 96 99
rect 94 98 95 99
rect 93 98 94 99
rect 92 98 93 99
rect 91 98 92 99
rect 90 98 91 99
rect 89 98 90 99
rect 88 98 89 99
rect 87 98 88 99
rect 86 98 87 99
rect 85 98 86 99
rect 84 98 85 99
rect 83 98 84 99
rect 82 98 83 99
rect 81 98 82 99
rect 80 98 81 99
rect 79 98 80 99
rect 78 98 79 99
rect 77 98 78 99
rect 76 98 77 99
rect 75 98 76 99
rect 74 98 75 99
rect 73 98 74 99
rect 72 98 73 99
rect 67 98 68 99
rect 66 98 67 99
rect 65 98 66 99
rect 64 98 65 99
rect 63 98 64 99
rect 62 98 63 99
rect 61 98 62 99
rect 60 98 61 99
rect 59 98 60 99
rect 58 98 59 99
rect 57 98 58 99
rect 56 98 57 99
rect 55 98 56 99
rect 54 98 55 99
rect 53 98 54 99
rect 52 98 53 99
rect 51 98 52 99
rect 50 98 51 99
rect 49 98 50 99
rect 48 98 49 99
rect 461 99 462 100
rect 460 99 461 100
rect 459 99 460 100
rect 458 99 459 100
rect 263 99 264 100
rect 262 99 263 100
rect 261 99 262 100
rect 260 99 261 100
rect 259 99 260 100
rect 258 99 259 100
rect 257 99 258 100
rect 256 99 257 100
rect 255 99 256 100
rect 254 99 255 100
rect 253 99 254 100
rect 252 99 253 100
rect 251 99 252 100
rect 250 99 251 100
rect 249 99 250 100
rect 248 99 249 100
rect 247 99 248 100
rect 246 99 247 100
rect 245 99 246 100
rect 244 99 245 100
rect 243 99 244 100
rect 242 99 243 100
rect 241 99 242 100
rect 240 99 241 100
rect 239 99 240 100
rect 238 99 239 100
rect 237 99 238 100
rect 236 99 237 100
rect 235 99 236 100
rect 234 99 235 100
rect 233 99 234 100
rect 232 99 233 100
rect 231 99 232 100
rect 230 99 231 100
rect 229 99 230 100
rect 228 99 229 100
rect 227 99 228 100
rect 226 99 227 100
rect 225 99 226 100
rect 224 99 225 100
rect 223 99 224 100
rect 222 99 223 100
rect 221 99 222 100
rect 220 99 221 100
rect 219 99 220 100
rect 218 99 219 100
rect 217 99 218 100
rect 216 99 217 100
rect 215 99 216 100
rect 214 99 215 100
rect 213 99 214 100
rect 212 99 213 100
rect 211 99 212 100
rect 210 99 211 100
rect 209 99 210 100
rect 208 99 209 100
rect 207 99 208 100
rect 206 99 207 100
rect 205 99 206 100
rect 204 99 205 100
rect 203 99 204 100
rect 202 99 203 100
rect 201 99 202 100
rect 200 99 201 100
rect 199 99 200 100
rect 198 99 199 100
rect 197 99 198 100
rect 196 99 197 100
rect 195 99 196 100
rect 194 99 195 100
rect 193 99 194 100
rect 192 99 193 100
rect 191 99 192 100
rect 190 99 191 100
rect 189 99 190 100
rect 188 99 189 100
rect 187 99 188 100
rect 186 99 187 100
rect 185 99 186 100
rect 184 99 185 100
rect 183 99 184 100
rect 182 99 183 100
rect 181 99 182 100
rect 180 99 181 100
rect 179 99 180 100
rect 178 99 179 100
rect 177 99 178 100
rect 156 99 157 100
rect 155 99 156 100
rect 154 99 155 100
rect 153 99 154 100
rect 152 99 153 100
rect 151 99 152 100
rect 150 99 151 100
rect 149 99 150 100
rect 148 99 149 100
rect 147 99 148 100
rect 146 99 147 100
rect 145 99 146 100
rect 144 99 145 100
rect 143 99 144 100
rect 142 99 143 100
rect 141 99 142 100
rect 140 99 141 100
rect 139 99 140 100
rect 138 99 139 100
rect 137 99 138 100
rect 136 99 137 100
rect 135 99 136 100
rect 134 99 135 100
rect 133 99 134 100
rect 132 99 133 100
rect 131 99 132 100
rect 130 99 131 100
rect 129 99 130 100
rect 128 99 129 100
rect 127 99 128 100
rect 126 99 127 100
rect 116 99 117 100
rect 115 99 116 100
rect 114 99 115 100
rect 113 99 114 100
rect 112 99 113 100
rect 111 99 112 100
rect 110 99 111 100
rect 109 99 110 100
rect 108 99 109 100
rect 107 99 108 100
rect 106 99 107 100
rect 105 99 106 100
rect 104 99 105 100
rect 103 99 104 100
rect 102 99 103 100
rect 101 99 102 100
rect 100 99 101 100
rect 99 99 100 100
rect 98 99 99 100
rect 97 99 98 100
rect 96 99 97 100
rect 95 99 96 100
rect 94 99 95 100
rect 93 99 94 100
rect 92 99 93 100
rect 91 99 92 100
rect 90 99 91 100
rect 89 99 90 100
rect 88 99 89 100
rect 87 99 88 100
rect 86 99 87 100
rect 85 99 86 100
rect 84 99 85 100
rect 83 99 84 100
rect 82 99 83 100
rect 81 99 82 100
rect 80 99 81 100
rect 79 99 80 100
rect 78 99 79 100
rect 77 99 78 100
rect 76 99 77 100
rect 75 99 76 100
rect 74 99 75 100
rect 73 99 74 100
rect 72 99 73 100
rect 67 99 68 100
rect 66 99 67 100
rect 65 99 66 100
rect 64 99 65 100
rect 63 99 64 100
rect 62 99 63 100
rect 61 99 62 100
rect 60 99 61 100
rect 59 99 60 100
rect 58 99 59 100
rect 57 99 58 100
rect 56 99 57 100
rect 55 99 56 100
rect 54 99 55 100
rect 53 99 54 100
rect 52 99 53 100
rect 51 99 52 100
rect 50 99 51 100
rect 49 99 50 100
rect 48 99 49 100
rect 47 99 48 100
rect 459 100 460 101
rect 458 100 459 101
rect 395 100 396 101
rect 394 100 395 101
rect 393 100 394 101
rect 265 100 266 101
rect 264 100 265 101
rect 263 100 264 101
rect 262 100 263 101
rect 261 100 262 101
rect 260 100 261 101
rect 259 100 260 101
rect 258 100 259 101
rect 257 100 258 101
rect 256 100 257 101
rect 255 100 256 101
rect 254 100 255 101
rect 253 100 254 101
rect 252 100 253 101
rect 251 100 252 101
rect 250 100 251 101
rect 249 100 250 101
rect 248 100 249 101
rect 247 100 248 101
rect 246 100 247 101
rect 245 100 246 101
rect 244 100 245 101
rect 243 100 244 101
rect 242 100 243 101
rect 241 100 242 101
rect 240 100 241 101
rect 239 100 240 101
rect 238 100 239 101
rect 237 100 238 101
rect 236 100 237 101
rect 235 100 236 101
rect 234 100 235 101
rect 233 100 234 101
rect 232 100 233 101
rect 231 100 232 101
rect 230 100 231 101
rect 229 100 230 101
rect 228 100 229 101
rect 227 100 228 101
rect 226 100 227 101
rect 225 100 226 101
rect 224 100 225 101
rect 223 100 224 101
rect 222 100 223 101
rect 221 100 222 101
rect 220 100 221 101
rect 219 100 220 101
rect 218 100 219 101
rect 217 100 218 101
rect 216 100 217 101
rect 215 100 216 101
rect 214 100 215 101
rect 213 100 214 101
rect 212 100 213 101
rect 211 100 212 101
rect 210 100 211 101
rect 209 100 210 101
rect 208 100 209 101
rect 207 100 208 101
rect 206 100 207 101
rect 205 100 206 101
rect 204 100 205 101
rect 203 100 204 101
rect 202 100 203 101
rect 201 100 202 101
rect 200 100 201 101
rect 199 100 200 101
rect 198 100 199 101
rect 197 100 198 101
rect 196 100 197 101
rect 195 100 196 101
rect 194 100 195 101
rect 193 100 194 101
rect 192 100 193 101
rect 191 100 192 101
rect 190 100 191 101
rect 189 100 190 101
rect 188 100 189 101
rect 187 100 188 101
rect 186 100 187 101
rect 185 100 186 101
rect 184 100 185 101
rect 183 100 184 101
rect 182 100 183 101
rect 181 100 182 101
rect 180 100 181 101
rect 179 100 180 101
rect 178 100 179 101
rect 177 100 178 101
rect 176 100 177 101
rect 155 100 156 101
rect 154 100 155 101
rect 153 100 154 101
rect 152 100 153 101
rect 151 100 152 101
rect 150 100 151 101
rect 149 100 150 101
rect 148 100 149 101
rect 147 100 148 101
rect 146 100 147 101
rect 145 100 146 101
rect 144 100 145 101
rect 143 100 144 101
rect 142 100 143 101
rect 141 100 142 101
rect 140 100 141 101
rect 139 100 140 101
rect 138 100 139 101
rect 137 100 138 101
rect 136 100 137 101
rect 135 100 136 101
rect 134 100 135 101
rect 133 100 134 101
rect 132 100 133 101
rect 131 100 132 101
rect 130 100 131 101
rect 129 100 130 101
rect 128 100 129 101
rect 127 100 128 101
rect 126 100 127 101
rect 115 100 116 101
rect 114 100 115 101
rect 113 100 114 101
rect 112 100 113 101
rect 111 100 112 101
rect 110 100 111 101
rect 109 100 110 101
rect 108 100 109 101
rect 107 100 108 101
rect 106 100 107 101
rect 105 100 106 101
rect 104 100 105 101
rect 103 100 104 101
rect 102 100 103 101
rect 101 100 102 101
rect 100 100 101 101
rect 99 100 100 101
rect 98 100 99 101
rect 97 100 98 101
rect 96 100 97 101
rect 95 100 96 101
rect 94 100 95 101
rect 93 100 94 101
rect 92 100 93 101
rect 91 100 92 101
rect 90 100 91 101
rect 89 100 90 101
rect 88 100 89 101
rect 87 100 88 101
rect 86 100 87 101
rect 85 100 86 101
rect 84 100 85 101
rect 83 100 84 101
rect 82 100 83 101
rect 81 100 82 101
rect 80 100 81 101
rect 79 100 80 101
rect 78 100 79 101
rect 77 100 78 101
rect 76 100 77 101
rect 75 100 76 101
rect 74 100 75 101
rect 73 100 74 101
rect 72 100 73 101
rect 66 100 67 101
rect 65 100 66 101
rect 64 100 65 101
rect 63 100 64 101
rect 62 100 63 101
rect 61 100 62 101
rect 60 100 61 101
rect 59 100 60 101
rect 58 100 59 101
rect 57 100 58 101
rect 56 100 57 101
rect 55 100 56 101
rect 54 100 55 101
rect 53 100 54 101
rect 52 100 53 101
rect 51 100 52 101
rect 50 100 51 101
rect 49 100 50 101
rect 48 100 49 101
rect 47 100 48 101
rect 46 100 47 101
rect 458 101 459 102
rect 395 101 396 102
rect 394 101 395 102
rect 393 101 394 102
rect 266 101 267 102
rect 265 101 266 102
rect 264 101 265 102
rect 263 101 264 102
rect 262 101 263 102
rect 261 101 262 102
rect 260 101 261 102
rect 259 101 260 102
rect 258 101 259 102
rect 257 101 258 102
rect 256 101 257 102
rect 255 101 256 102
rect 254 101 255 102
rect 253 101 254 102
rect 252 101 253 102
rect 251 101 252 102
rect 250 101 251 102
rect 249 101 250 102
rect 248 101 249 102
rect 247 101 248 102
rect 246 101 247 102
rect 245 101 246 102
rect 244 101 245 102
rect 243 101 244 102
rect 242 101 243 102
rect 241 101 242 102
rect 240 101 241 102
rect 239 101 240 102
rect 238 101 239 102
rect 237 101 238 102
rect 236 101 237 102
rect 235 101 236 102
rect 234 101 235 102
rect 233 101 234 102
rect 232 101 233 102
rect 231 101 232 102
rect 230 101 231 102
rect 229 101 230 102
rect 228 101 229 102
rect 227 101 228 102
rect 226 101 227 102
rect 225 101 226 102
rect 224 101 225 102
rect 223 101 224 102
rect 222 101 223 102
rect 221 101 222 102
rect 220 101 221 102
rect 219 101 220 102
rect 218 101 219 102
rect 217 101 218 102
rect 216 101 217 102
rect 215 101 216 102
rect 214 101 215 102
rect 213 101 214 102
rect 212 101 213 102
rect 211 101 212 102
rect 210 101 211 102
rect 209 101 210 102
rect 208 101 209 102
rect 207 101 208 102
rect 206 101 207 102
rect 205 101 206 102
rect 204 101 205 102
rect 203 101 204 102
rect 202 101 203 102
rect 201 101 202 102
rect 200 101 201 102
rect 199 101 200 102
rect 198 101 199 102
rect 197 101 198 102
rect 196 101 197 102
rect 195 101 196 102
rect 194 101 195 102
rect 193 101 194 102
rect 192 101 193 102
rect 191 101 192 102
rect 190 101 191 102
rect 189 101 190 102
rect 188 101 189 102
rect 187 101 188 102
rect 186 101 187 102
rect 185 101 186 102
rect 184 101 185 102
rect 183 101 184 102
rect 182 101 183 102
rect 181 101 182 102
rect 180 101 181 102
rect 179 101 180 102
rect 178 101 179 102
rect 177 101 178 102
rect 176 101 177 102
rect 175 101 176 102
rect 155 101 156 102
rect 154 101 155 102
rect 153 101 154 102
rect 152 101 153 102
rect 151 101 152 102
rect 150 101 151 102
rect 149 101 150 102
rect 148 101 149 102
rect 147 101 148 102
rect 146 101 147 102
rect 145 101 146 102
rect 144 101 145 102
rect 143 101 144 102
rect 142 101 143 102
rect 141 101 142 102
rect 140 101 141 102
rect 139 101 140 102
rect 138 101 139 102
rect 137 101 138 102
rect 136 101 137 102
rect 135 101 136 102
rect 134 101 135 102
rect 133 101 134 102
rect 132 101 133 102
rect 131 101 132 102
rect 130 101 131 102
rect 129 101 130 102
rect 128 101 129 102
rect 127 101 128 102
rect 126 101 127 102
rect 125 101 126 102
rect 114 101 115 102
rect 113 101 114 102
rect 112 101 113 102
rect 111 101 112 102
rect 110 101 111 102
rect 109 101 110 102
rect 108 101 109 102
rect 107 101 108 102
rect 106 101 107 102
rect 105 101 106 102
rect 104 101 105 102
rect 103 101 104 102
rect 102 101 103 102
rect 101 101 102 102
rect 100 101 101 102
rect 99 101 100 102
rect 98 101 99 102
rect 97 101 98 102
rect 96 101 97 102
rect 95 101 96 102
rect 94 101 95 102
rect 93 101 94 102
rect 92 101 93 102
rect 91 101 92 102
rect 90 101 91 102
rect 89 101 90 102
rect 88 101 89 102
rect 87 101 88 102
rect 86 101 87 102
rect 85 101 86 102
rect 84 101 85 102
rect 83 101 84 102
rect 82 101 83 102
rect 81 101 82 102
rect 80 101 81 102
rect 79 101 80 102
rect 78 101 79 102
rect 77 101 78 102
rect 76 101 77 102
rect 75 101 76 102
rect 74 101 75 102
rect 73 101 74 102
rect 72 101 73 102
rect 66 101 67 102
rect 65 101 66 102
rect 64 101 65 102
rect 63 101 64 102
rect 62 101 63 102
rect 61 101 62 102
rect 60 101 61 102
rect 59 101 60 102
rect 58 101 59 102
rect 57 101 58 102
rect 56 101 57 102
rect 55 101 56 102
rect 54 101 55 102
rect 53 101 54 102
rect 52 101 53 102
rect 51 101 52 102
rect 50 101 51 102
rect 49 101 50 102
rect 48 101 49 102
rect 47 101 48 102
rect 46 101 47 102
rect 45 101 46 102
rect 395 102 396 103
rect 394 102 395 103
rect 393 102 394 103
rect 267 102 268 103
rect 266 102 267 103
rect 265 102 266 103
rect 264 102 265 103
rect 263 102 264 103
rect 262 102 263 103
rect 261 102 262 103
rect 260 102 261 103
rect 259 102 260 103
rect 258 102 259 103
rect 257 102 258 103
rect 256 102 257 103
rect 255 102 256 103
rect 254 102 255 103
rect 253 102 254 103
rect 252 102 253 103
rect 251 102 252 103
rect 250 102 251 103
rect 249 102 250 103
rect 248 102 249 103
rect 247 102 248 103
rect 246 102 247 103
rect 245 102 246 103
rect 244 102 245 103
rect 243 102 244 103
rect 242 102 243 103
rect 241 102 242 103
rect 240 102 241 103
rect 239 102 240 103
rect 238 102 239 103
rect 237 102 238 103
rect 236 102 237 103
rect 235 102 236 103
rect 234 102 235 103
rect 233 102 234 103
rect 232 102 233 103
rect 231 102 232 103
rect 230 102 231 103
rect 229 102 230 103
rect 228 102 229 103
rect 227 102 228 103
rect 226 102 227 103
rect 225 102 226 103
rect 224 102 225 103
rect 223 102 224 103
rect 222 102 223 103
rect 221 102 222 103
rect 220 102 221 103
rect 219 102 220 103
rect 218 102 219 103
rect 217 102 218 103
rect 216 102 217 103
rect 215 102 216 103
rect 214 102 215 103
rect 213 102 214 103
rect 212 102 213 103
rect 211 102 212 103
rect 210 102 211 103
rect 209 102 210 103
rect 208 102 209 103
rect 207 102 208 103
rect 206 102 207 103
rect 205 102 206 103
rect 204 102 205 103
rect 203 102 204 103
rect 202 102 203 103
rect 201 102 202 103
rect 200 102 201 103
rect 199 102 200 103
rect 198 102 199 103
rect 197 102 198 103
rect 196 102 197 103
rect 195 102 196 103
rect 194 102 195 103
rect 193 102 194 103
rect 192 102 193 103
rect 191 102 192 103
rect 190 102 191 103
rect 189 102 190 103
rect 188 102 189 103
rect 187 102 188 103
rect 186 102 187 103
rect 185 102 186 103
rect 184 102 185 103
rect 183 102 184 103
rect 182 102 183 103
rect 181 102 182 103
rect 180 102 181 103
rect 179 102 180 103
rect 178 102 179 103
rect 177 102 178 103
rect 176 102 177 103
rect 175 102 176 103
rect 155 102 156 103
rect 154 102 155 103
rect 153 102 154 103
rect 152 102 153 103
rect 151 102 152 103
rect 150 102 151 103
rect 149 102 150 103
rect 148 102 149 103
rect 147 102 148 103
rect 146 102 147 103
rect 145 102 146 103
rect 144 102 145 103
rect 143 102 144 103
rect 142 102 143 103
rect 141 102 142 103
rect 140 102 141 103
rect 139 102 140 103
rect 138 102 139 103
rect 137 102 138 103
rect 136 102 137 103
rect 135 102 136 103
rect 134 102 135 103
rect 133 102 134 103
rect 132 102 133 103
rect 131 102 132 103
rect 130 102 131 103
rect 129 102 130 103
rect 128 102 129 103
rect 127 102 128 103
rect 126 102 127 103
rect 125 102 126 103
rect 114 102 115 103
rect 113 102 114 103
rect 112 102 113 103
rect 111 102 112 103
rect 110 102 111 103
rect 109 102 110 103
rect 108 102 109 103
rect 107 102 108 103
rect 106 102 107 103
rect 105 102 106 103
rect 104 102 105 103
rect 103 102 104 103
rect 102 102 103 103
rect 101 102 102 103
rect 100 102 101 103
rect 99 102 100 103
rect 98 102 99 103
rect 97 102 98 103
rect 96 102 97 103
rect 95 102 96 103
rect 94 102 95 103
rect 93 102 94 103
rect 92 102 93 103
rect 91 102 92 103
rect 90 102 91 103
rect 89 102 90 103
rect 88 102 89 103
rect 87 102 88 103
rect 86 102 87 103
rect 85 102 86 103
rect 84 102 85 103
rect 83 102 84 103
rect 82 102 83 103
rect 81 102 82 103
rect 80 102 81 103
rect 79 102 80 103
rect 78 102 79 103
rect 77 102 78 103
rect 76 102 77 103
rect 75 102 76 103
rect 74 102 75 103
rect 73 102 74 103
rect 72 102 73 103
rect 71 102 72 103
rect 65 102 66 103
rect 64 102 65 103
rect 63 102 64 103
rect 62 102 63 103
rect 61 102 62 103
rect 60 102 61 103
rect 59 102 60 103
rect 58 102 59 103
rect 57 102 58 103
rect 56 102 57 103
rect 55 102 56 103
rect 54 102 55 103
rect 53 102 54 103
rect 52 102 53 103
rect 51 102 52 103
rect 50 102 51 103
rect 49 102 50 103
rect 48 102 49 103
rect 47 102 48 103
rect 46 102 47 103
rect 45 102 46 103
rect 44 102 45 103
rect 395 103 396 104
rect 394 103 395 104
rect 393 103 394 104
rect 268 103 269 104
rect 267 103 268 104
rect 266 103 267 104
rect 265 103 266 104
rect 264 103 265 104
rect 263 103 264 104
rect 262 103 263 104
rect 261 103 262 104
rect 260 103 261 104
rect 259 103 260 104
rect 258 103 259 104
rect 257 103 258 104
rect 256 103 257 104
rect 255 103 256 104
rect 254 103 255 104
rect 253 103 254 104
rect 252 103 253 104
rect 251 103 252 104
rect 250 103 251 104
rect 249 103 250 104
rect 248 103 249 104
rect 247 103 248 104
rect 246 103 247 104
rect 245 103 246 104
rect 244 103 245 104
rect 243 103 244 104
rect 242 103 243 104
rect 241 103 242 104
rect 240 103 241 104
rect 239 103 240 104
rect 238 103 239 104
rect 237 103 238 104
rect 236 103 237 104
rect 235 103 236 104
rect 234 103 235 104
rect 233 103 234 104
rect 232 103 233 104
rect 231 103 232 104
rect 230 103 231 104
rect 229 103 230 104
rect 228 103 229 104
rect 227 103 228 104
rect 226 103 227 104
rect 225 103 226 104
rect 224 103 225 104
rect 223 103 224 104
rect 222 103 223 104
rect 221 103 222 104
rect 220 103 221 104
rect 219 103 220 104
rect 218 103 219 104
rect 217 103 218 104
rect 216 103 217 104
rect 215 103 216 104
rect 214 103 215 104
rect 213 103 214 104
rect 212 103 213 104
rect 211 103 212 104
rect 210 103 211 104
rect 209 103 210 104
rect 208 103 209 104
rect 207 103 208 104
rect 206 103 207 104
rect 205 103 206 104
rect 204 103 205 104
rect 203 103 204 104
rect 202 103 203 104
rect 201 103 202 104
rect 200 103 201 104
rect 199 103 200 104
rect 198 103 199 104
rect 197 103 198 104
rect 196 103 197 104
rect 195 103 196 104
rect 194 103 195 104
rect 193 103 194 104
rect 192 103 193 104
rect 191 103 192 104
rect 190 103 191 104
rect 189 103 190 104
rect 188 103 189 104
rect 187 103 188 104
rect 186 103 187 104
rect 185 103 186 104
rect 184 103 185 104
rect 183 103 184 104
rect 182 103 183 104
rect 181 103 182 104
rect 180 103 181 104
rect 179 103 180 104
rect 178 103 179 104
rect 177 103 178 104
rect 176 103 177 104
rect 175 103 176 104
rect 174 103 175 104
rect 154 103 155 104
rect 153 103 154 104
rect 152 103 153 104
rect 151 103 152 104
rect 150 103 151 104
rect 149 103 150 104
rect 148 103 149 104
rect 147 103 148 104
rect 146 103 147 104
rect 145 103 146 104
rect 144 103 145 104
rect 143 103 144 104
rect 142 103 143 104
rect 141 103 142 104
rect 140 103 141 104
rect 139 103 140 104
rect 138 103 139 104
rect 137 103 138 104
rect 136 103 137 104
rect 135 103 136 104
rect 134 103 135 104
rect 133 103 134 104
rect 132 103 133 104
rect 131 103 132 104
rect 130 103 131 104
rect 129 103 130 104
rect 128 103 129 104
rect 127 103 128 104
rect 126 103 127 104
rect 125 103 126 104
rect 113 103 114 104
rect 112 103 113 104
rect 111 103 112 104
rect 110 103 111 104
rect 109 103 110 104
rect 108 103 109 104
rect 107 103 108 104
rect 106 103 107 104
rect 105 103 106 104
rect 104 103 105 104
rect 103 103 104 104
rect 102 103 103 104
rect 101 103 102 104
rect 100 103 101 104
rect 99 103 100 104
rect 98 103 99 104
rect 97 103 98 104
rect 96 103 97 104
rect 95 103 96 104
rect 94 103 95 104
rect 93 103 94 104
rect 92 103 93 104
rect 91 103 92 104
rect 90 103 91 104
rect 89 103 90 104
rect 88 103 89 104
rect 87 103 88 104
rect 86 103 87 104
rect 85 103 86 104
rect 84 103 85 104
rect 83 103 84 104
rect 82 103 83 104
rect 81 103 82 104
rect 80 103 81 104
rect 79 103 80 104
rect 78 103 79 104
rect 77 103 78 104
rect 76 103 77 104
rect 75 103 76 104
rect 74 103 75 104
rect 73 103 74 104
rect 72 103 73 104
rect 71 103 72 104
rect 65 103 66 104
rect 64 103 65 104
rect 63 103 64 104
rect 62 103 63 104
rect 61 103 62 104
rect 60 103 61 104
rect 59 103 60 104
rect 58 103 59 104
rect 57 103 58 104
rect 56 103 57 104
rect 55 103 56 104
rect 54 103 55 104
rect 53 103 54 104
rect 52 103 53 104
rect 51 103 52 104
rect 50 103 51 104
rect 49 103 50 104
rect 48 103 49 104
rect 47 103 48 104
rect 46 103 47 104
rect 45 103 46 104
rect 44 103 45 104
rect 43 103 44 104
rect 42 103 43 104
rect 396 104 397 105
rect 395 104 396 105
rect 394 104 395 105
rect 393 104 394 105
rect 269 104 270 105
rect 268 104 269 105
rect 267 104 268 105
rect 266 104 267 105
rect 265 104 266 105
rect 264 104 265 105
rect 263 104 264 105
rect 262 104 263 105
rect 261 104 262 105
rect 260 104 261 105
rect 259 104 260 105
rect 258 104 259 105
rect 257 104 258 105
rect 256 104 257 105
rect 255 104 256 105
rect 254 104 255 105
rect 253 104 254 105
rect 252 104 253 105
rect 251 104 252 105
rect 250 104 251 105
rect 249 104 250 105
rect 248 104 249 105
rect 247 104 248 105
rect 246 104 247 105
rect 245 104 246 105
rect 244 104 245 105
rect 243 104 244 105
rect 242 104 243 105
rect 241 104 242 105
rect 240 104 241 105
rect 239 104 240 105
rect 238 104 239 105
rect 237 104 238 105
rect 236 104 237 105
rect 235 104 236 105
rect 234 104 235 105
rect 233 104 234 105
rect 232 104 233 105
rect 231 104 232 105
rect 230 104 231 105
rect 229 104 230 105
rect 228 104 229 105
rect 227 104 228 105
rect 226 104 227 105
rect 225 104 226 105
rect 224 104 225 105
rect 223 104 224 105
rect 222 104 223 105
rect 221 104 222 105
rect 220 104 221 105
rect 219 104 220 105
rect 218 104 219 105
rect 217 104 218 105
rect 216 104 217 105
rect 215 104 216 105
rect 214 104 215 105
rect 213 104 214 105
rect 212 104 213 105
rect 211 104 212 105
rect 210 104 211 105
rect 209 104 210 105
rect 208 104 209 105
rect 207 104 208 105
rect 206 104 207 105
rect 205 104 206 105
rect 204 104 205 105
rect 203 104 204 105
rect 202 104 203 105
rect 201 104 202 105
rect 200 104 201 105
rect 199 104 200 105
rect 198 104 199 105
rect 197 104 198 105
rect 196 104 197 105
rect 195 104 196 105
rect 194 104 195 105
rect 193 104 194 105
rect 192 104 193 105
rect 191 104 192 105
rect 190 104 191 105
rect 189 104 190 105
rect 188 104 189 105
rect 187 104 188 105
rect 186 104 187 105
rect 185 104 186 105
rect 184 104 185 105
rect 183 104 184 105
rect 182 104 183 105
rect 181 104 182 105
rect 180 104 181 105
rect 179 104 180 105
rect 178 104 179 105
rect 177 104 178 105
rect 176 104 177 105
rect 175 104 176 105
rect 174 104 175 105
rect 173 104 174 105
rect 154 104 155 105
rect 153 104 154 105
rect 152 104 153 105
rect 151 104 152 105
rect 150 104 151 105
rect 149 104 150 105
rect 148 104 149 105
rect 147 104 148 105
rect 146 104 147 105
rect 145 104 146 105
rect 144 104 145 105
rect 143 104 144 105
rect 142 104 143 105
rect 141 104 142 105
rect 140 104 141 105
rect 139 104 140 105
rect 138 104 139 105
rect 137 104 138 105
rect 136 104 137 105
rect 135 104 136 105
rect 134 104 135 105
rect 133 104 134 105
rect 132 104 133 105
rect 131 104 132 105
rect 130 104 131 105
rect 129 104 130 105
rect 128 104 129 105
rect 127 104 128 105
rect 126 104 127 105
rect 125 104 126 105
rect 124 104 125 105
rect 113 104 114 105
rect 112 104 113 105
rect 111 104 112 105
rect 110 104 111 105
rect 109 104 110 105
rect 108 104 109 105
rect 107 104 108 105
rect 106 104 107 105
rect 105 104 106 105
rect 104 104 105 105
rect 103 104 104 105
rect 102 104 103 105
rect 101 104 102 105
rect 100 104 101 105
rect 99 104 100 105
rect 98 104 99 105
rect 97 104 98 105
rect 96 104 97 105
rect 95 104 96 105
rect 94 104 95 105
rect 93 104 94 105
rect 92 104 93 105
rect 91 104 92 105
rect 90 104 91 105
rect 89 104 90 105
rect 88 104 89 105
rect 87 104 88 105
rect 86 104 87 105
rect 85 104 86 105
rect 84 104 85 105
rect 83 104 84 105
rect 82 104 83 105
rect 81 104 82 105
rect 80 104 81 105
rect 79 104 80 105
rect 78 104 79 105
rect 77 104 78 105
rect 76 104 77 105
rect 75 104 76 105
rect 64 104 65 105
rect 63 104 64 105
rect 62 104 63 105
rect 61 104 62 105
rect 60 104 61 105
rect 59 104 60 105
rect 58 104 59 105
rect 57 104 58 105
rect 56 104 57 105
rect 55 104 56 105
rect 54 104 55 105
rect 53 104 54 105
rect 52 104 53 105
rect 51 104 52 105
rect 50 104 51 105
rect 49 104 50 105
rect 48 104 49 105
rect 47 104 48 105
rect 46 104 47 105
rect 45 104 46 105
rect 44 104 45 105
rect 43 104 44 105
rect 42 104 43 105
rect 41 104 42 105
rect 421 105 422 106
rect 420 105 421 106
rect 419 105 420 106
rect 418 105 419 106
rect 417 105 418 106
rect 416 105 417 106
rect 415 105 416 106
rect 414 105 415 106
rect 413 105 414 106
rect 412 105 413 106
rect 411 105 412 106
rect 410 105 411 106
rect 409 105 410 106
rect 408 105 409 106
rect 407 105 408 106
rect 406 105 407 106
rect 405 105 406 106
rect 404 105 405 106
rect 403 105 404 106
rect 402 105 403 106
rect 401 105 402 106
rect 400 105 401 106
rect 399 105 400 106
rect 398 105 399 106
rect 397 105 398 106
rect 396 105 397 106
rect 395 105 396 106
rect 394 105 395 106
rect 393 105 394 106
rect 270 105 271 106
rect 269 105 270 106
rect 268 105 269 106
rect 267 105 268 106
rect 266 105 267 106
rect 265 105 266 106
rect 264 105 265 106
rect 263 105 264 106
rect 262 105 263 106
rect 261 105 262 106
rect 260 105 261 106
rect 259 105 260 106
rect 258 105 259 106
rect 257 105 258 106
rect 256 105 257 106
rect 255 105 256 106
rect 254 105 255 106
rect 253 105 254 106
rect 252 105 253 106
rect 251 105 252 106
rect 250 105 251 106
rect 249 105 250 106
rect 248 105 249 106
rect 247 105 248 106
rect 246 105 247 106
rect 245 105 246 106
rect 244 105 245 106
rect 243 105 244 106
rect 242 105 243 106
rect 241 105 242 106
rect 240 105 241 106
rect 239 105 240 106
rect 238 105 239 106
rect 237 105 238 106
rect 236 105 237 106
rect 235 105 236 106
rect 234 105 235 106
rect 233 105 234 106
rect 232 105 233 106
rect 231 105 232 106
rect 230 105 231 106
rect 229 105 230 106
rect 228 105 229 106
rect 227 105 228 106
rect 226 105 227 106
rect 225 105 226 106
rect 224 105 225 106
rect 223 105 224 106
rect 222 105 223 106
rect 221 105 222 106
rect 220 105 221 106
rect 219 105 220 106
rect 218 105 219 106
rect 217 105 218 106
rect 216 105 217 106
rect 215 105 216 106
rect 214 105 215 106
rect 213 105 214 106
rect 212 105 213 106
rect 211 105 212 106
rect 210 105 211 106
rect 209 105 210 106
rect 208 105 209 106
rect 207 105 208 106
rect 206 105 207 106
rect 205 105 206 106
rect 204 105 205 106
rect 203 105 204 106
rect 202 105 203 106
rect 201 105 202 106
rect 200 105 201 106
rect 199 105 200 106
rect 198 105 199 106
rect 197 105 198 106
rect 196 105 197 106
rect 195 105 196 106
rect 194 105 195 106
rect 193 105 194 106
rect 192 105 193 106
rect 191 105 192 106
rect 190 105 191 106
rect 189 105 190 106
rect 188 105 189 106
rect 187 105 188 106
rect 186 105 187 106
rect 185 105 186 106
rect 184 105 185 106
rect 183 105 184 106
rect 182 105 183 106
rect 181 105 182 106
rect 180 105 181 106
rect 179 105 180 106
rect 178 105 179 106
rect 177 105 178 106
rect 176 105 177 106
rect 175 105 176 106
rect 174 105 175 106
rect 173 105 174 106
rect 154 105 155 106
rect 153 105 154 106
rect 152 105 153 106
rect 151 105 152 106
rect 150 105 151 106
rect 149 105 150 106
rect 148 105 149 106
rect 147 105 148 106
rect 146 105 147 106
rect 145 105 146 106
rect 144 105 145 106
rect 143 105 144 106
rect 142 105 143 106
rect 141 105 142 106
rect 140 105 141 106
rect 139 105 140 106
rect 138 105 139 106
rect 137 105 138 106
rect 136 105 137 106
rect 135 105 136 106
rect 134 105 135 106
rect 133 105 134 106
rect 132 105 133 106
rect 131 105 132 106
rect 130 105 131 106
rect 129 105 130 106
rect 128 105 129 106
rect 127 105 128 106
rect 126 105 127 106
rect 125 105 126 106
rect 124 105 125 106
rect 114 105 115 106
rect 113 105 114 106
rect 112 105 113 106
rect 111 105 112 106
rect 110 105 111 106
rect 109 105 110 106
rect 108 105 109 106
rect 107 105 108 106
rect 106 105 107 106
rect 105 105 106 106
rect 104 105 105 106
rect 103 105 104 106
rect 102 105 103 106
rect 101 105 102 106
rect 100 105 101 106
rect 99 105 100 106
rect 98 105 99 106
rect 97 105 98 106
rect 96 105 97 106
rect 95 105 96 106
rect 94 105 95 106
rect 93 105 94 106
rect 92 105 93 106
rect 91 105 92 106
rect 90 105 91 106
rect 89 105 90 106
rect 88 105 89 106
rect 87 105 88 106
rect 86 105 87 106
rect 85 105 86 106
rect 84 105 85 106
rect 83 105 84 106
rect 82 105 83 106
rect 81 105 82 106
rect 80 105 81 106
rect 79 105 80 106
rect 78 105 79 106
rect 63 105 64 106
rect 62 105 63 106
rect 61 105 62 106
rect 60 105 61 106
rect 59 105 60 106
rect 58 105 59 106
rect 57 105 58 106
rect 56 105 57 106
rect 55 105 56 106
rect 54 105 55 106
rect 53 105 54 106
rect 52 105 53 106
rect 51 105 52 106
rect 50 105 51 106
rect 49 105 50 106
rect 48 105 49 106
rect 47 105 48 106
rect 46 105 47 106
rect 45 105 46 106
rect 44 105 45 106
rect 43 105 44 106
rect 42 105 43 106
rect 41 105 42 106
rect 40 105 41 106
rect 39 105 40 106
rect 427 106 428 107
rect 426 106 427 107
rect 425 106 426 107
rect 424 106 425 107
rect 423 106 424 107
rect 422 106 423 107
rect 421 106 422 107
rect 420 106 421 107
rect 419 106 420 107
rect 418 106 419 107
rect 417 106 418 107
rect 416 106 417 107
rect 415 106 416 107
rect 414 106 415 107
rect 413 106 414 107
rect 412 106 413 107
rect 411 106 412 107
rect 410 106 411 107
rect 409 106 410 107
rect 408 106 409 107
rect 407 106 408 107
rect 406 106 407 107
rect 405 106 406 107
rect 404 106 405 107
rect 403 106 404 107
rect 402 106 403 107
rect 401 106 402 107
rect 400 106 401 107
rect 399 106 400 107
rect 398 106 399 107
rect 397 106 398 107
rect 396 106 397 107
rect 395 106 396 107
rect 394 106 395 107
rect 393 106 394 107
rect 271 106 272 107
rect 270 106 271 107
rect 269 106 270 107
rect 268 106 269 107
rect 267 106 268 107
rect 266 106 267 107
rect 265 106 266 107
rect 264 106 265 107
rect 263 106 264 107
rect 262 106 263 107
rect 261 106 262 107
rect 260 106 261 107
rect 259 106 260 107
rect 258 106 259 107
rect 257 106 258 107
rect 256 106 257 107
rect 255 106 256 107
rect 254 106 255 107
rect 253 106 254 107
rect 252 106 253 107
rect 251 106 252 107
rect 250 106 251 107
rect 249 106 250 107
rect 248 106 249 107
rect 247 106 248 107
rect 246 106 247 107
rect 245 106 246 107
rect 244 106 245 107
rect 243 106 244 107
rect 242 106 243 107
rect 241 106 242 107
rect 240 106 241 107
rect 239 106 240 107
rect 238 106 239 107
rect 237 106 238 107
rect 236 106 237 107
rect 235 106 236 107
rect 234 106 235 107
rect 233 106 234 107
rect 232 106 233 107
rect 231 106 232 107
rect 230 106 231 107
rect 229 106 230 107
rect 228 106 229 107
rect 227 106 228 107
rect 226 106 227 107
rect 225 106 226 107
rect 224 106 225 107
rect 223 106 224 107
rect 222 106 223 107
rect 221 106 222 107
rect 220 106 221 107
rect 219 106 220 107
rect 218 106 219 107
rect 217 106 218 107
rect 216 106 217 107
rect 215 106 216 107
rect 214 106 215 107
rect 213 106 214 107
rect 212 106 213 107
rect 211 106 212 107
rect 210 106 211 107
rect 209 106 210 107
rect 208 106 209 107
rect 207 106 208 107
rect 206 106 207 107
rect 205 106 206 107
rect 204 106 205 107
rect 203 106 204 107
rect 202 106 203 107
rect 201 106 202 107
rect 200 106 201 107
rect 199 106 200 107
rect 198 106 199 107
rect 197 106 198 107
rect 196 106 197 107
rect 195 106 196 107
rect 194 106 195 107
rect 193 106 194 107
rect 192 106 193 107
rect 191 106 192 107
rect 190 106 191 107
rect 189 106 190 107
rect 188 106 189 107
rect 187 106 188 107
rect 186 106 187 107
rect 185 106 186 107
rect 184 106 185 107
rect 183 106 184 107
rect 182 106 183 107
rect 181 106 182 107
rect 180 106 181 107
rect 179 106 180 107
rect 178 106 179 107
rect 177 106 178 107
rect 176 106 177 107
rect 175 106 176 107
rect 174 106 175 107
rect 173 106 174 107
rect 172 106 173 107
rect 153 106 154 107
rect 152 106 153 107
rect 151 106 152 107
rect 150 106 151 107
rect 149 106 150 107
rect 148 106 149 107
rect 147 106 148 107
rect 146 106 147 107
rect 145 106 146 107
rect 144 106 145 107
rect 143 106 144 107
rect 142 106 143 107
rect 141 106 142 107
rect 140 106 141 107
rect 139 106 140 107
rect 138 106 139 107
rect 137 106 138 107
rect 136 106 137 107
rect 135 106 136 107
rect 134 106 135 107
rect 133 106 134 107
rect 132 106 133 107
rect 131 106 132 107
rect 130 106 131 107
rect 129 106 130 107
rect 128 106 129 107
rect 127 106 128 107
rect 126 106 127 107
rect 125 106 126 107
rect 124 106 125 107
rect 114 106 115 107
rect 113 106 114 107
rect 112 106 113 107
rect 111 106 112 107
rect 110 106 111 107
rect 109 106 110 107
rect 108 106 109 107
rect 107 106 108 107
rect 106 106 107 107
rect 105 106 106 107
rect 104 106 105 107
rect 103 106 104 107
rect 102 106 103 107
rect 101 106 102 107
rect 100 106 101 107
rect 99 106 100 107
rect 98 106 99 107
rect 97 106 98 107
rect 96 106 97 107
rect 95 106 96 107
rect 94 106 95 107
rect 93 106 94 107
rect 92 106 93 107
rect 91 106 92 107
rect 90 106 91 107
rect 89 106 90 107
rect 88 106 89 107
rect 87 106 88 107
rect 86 106 87 107
rect 85 106 86 107
rect 84 106 85 107
rect 83 106 84 107
rect 82 106 83 107
rect 81 106 82 107
rect 80 106 81 107
rect 79 106 80 107
rect 63 106 64 107
rect 62 106 63 107
rect 61 106 62 107
rect 60 106 61 107
rect 59 106 60 107
rect 58 106 59 107
rect 57 106 58 107
rect 56 106 57 107
rect 55 106 56 107
rect 54 106 55 107
rect 53 106 54 107
rect 52 106 53 107
rect 51 106 52 107
rect 50 106 51 107
rect 49 106 50 107
rect 48 106 49 107
rect 47 106 48 107
rect 46 106 47 107
rect 45 106 46 107
rect 44 106 45 107
rect 43 106 44 107
rect 42 106 43 107
rect 41 106 42 107
rect 40 106 41 107
rect 39 106 40 107
rect 38 106 39 107
rect 430 107 431 108
rect 429 107 430 108
rect 428 107 429 108
rect 427 107 428 108
rect 426 107 427 108
rect 425 107 426 108
rect 424 107 425 108
rect 423 107 424 108
rect 422 107 423 108
rect 421 107 422 108
rect 420 107 421 108
rect 419 107 420 108
rect 418 107 419 108
rect 417 107 418 108
rect 416 107 417 108
rect 415 107 416 108
rect 414 107 415 108
rect 413 107 414 108
rect 412 107 413 108
rect 411 107 412 108
rect 410 107 411 108
rect 409 107 410 108
rect 408 107 409 108
rect 407 107 408 108
rect 406 107 407 108
rect 405 107 406 108
rect 404 107 405 108
rect 403 107 404 108
rect 402 107 403 108
rect 401 107 402 108
rect 400 107 401 108
rect 399 107 400 108
rect 398 107 399 108
rect 397 107 398 108
rect 396 107 397 108
rect 395 107 396 108
rect 394 107 395 108
rect 393 107 394 108
rect 272 107 273 108
rect 271 107 272 108
rect 270 107 271 108
rect 269 107 270 108
rect 268 107 269 108
rect 267 107 268 108
rect 266 107 267 108
rect 265 107 266 108
rect 264 107 265 108
rect 263 107 264 108
rect 262 107 263 108
rect 261 107 262 108
rect 260 107 261 108
rect 259 107 260 108
rect 258 107 259 108
rect 257 107 258 108
rect 256 107 257 108
rect 255 107 256 108
rect 254 107 255 108
rect 253 107 254 108
rect 252 107 253 108
rect 251 107 252 108
rect 250 107 251 108
rect 249 107 250 108
rect 248 107 249 108
rect 247 107 248 108
rect 246 107 247 108
rect 245 107 246 108
rect 244 107 245 108
rect 243 107 244 108
rect 242 107 243 108
rect 241 107 242 108
rect 240 107 241 108
rect 239 107 240 108
rect 238 107 239 108
rect 237 107 238 108
rect 236 107 237 108
rect 235 107 236 108
rect 234 107 235 108
rect 233 107 234 108
rect 232 107 233 108
rect 231 107 232 108
rect 230 107 231 108
rect 229 107 230 108
rect 228 107 229 108
rect 227 107 228 108
rect 226 107 227 108
rect 225 107 226 108
rect 224 107 225 108
rect 223 107 224 108
rect 222 107 223 108
rect 221 107 222 108
rect 220 107 221 108
rect 219 107 220 108
rect 218 107 219 108
rect 217 107 218 108
rect 216 107 217 108
rect 215 107 216 108
rect 214 107 215 108
rect 213 107 214 108
rect 212 107 213 108
rect 211 107 212 108
rect 210 107 211 108
rect 209 107 210 108
rect 208 107 209 108
rect 207 107 208 108
rect 206 107 207 108
rect 205 107 206 108
rect 204 107 205 108
rect 203 107 204 108
rect 202 107 203 108
rect 201 107 202 108
rect 200 107 201 108
rect 199 107 200 108
rect 198 107 199 108
rect 197 107 198 108
rect 196 107 197 108
rect 195 107 196 108
rect 194 107 195 108
rect 193 107 194 108
rect 192 107 193 108
rect 191 107 192 108
rect 190 107 191 108
rect 189 107 190 108
rect 188 107 189 108
rect 187 107 188 108
rect 186 107 187 108
rect 185 107 186 108
rect 184 107 185 108
rect 183 107 184 108
rect 182 107 183 108
rect 181 107 182 108
rect 180 107 181 108
rect 179 107 180 108
rect 178 107 179 108
rect 177 107 178 108
rect 176 107 177 108
rect 175 107 176 108
rect 174 107 175 108
rect 173 107 174 108
rect 172 107 173 108
rect 153 107 154 108
rect 152 107 153 108
rect 151 107 152 108
rect 150 107 151 108
rect 149 107 150 108
rect 148 107 149 108
rect 147 107 148 108
rect 146 107 147 108
rect 145 107 146 108
rect 144 107 145 108
rect 143 107 144 108
rect 142 107 143 108
rect 141 107 142 108
rect 140 107 141 108
rect 139 107 140 108
rect 138 107 139 108
rect 137 107 138 108
rect 136 107 137 108
rect 135 107 136 108
rect 134 107 135 108
rect 133 107 134 108
rect 132 107 133 108
rect 131 107 132 108
rect 130 107 131 108
rect 129 107 130 108
rect 128 107 129 108
rect 127 107 128 108
rect 126 107 127 108
rect 125 107 126 108
rect 124 107 125 108
rect 123 107 124 108
rect 115 107 116 108
rect 114 107 115 108
rect 113 107 114 108
rect 112 107 113 108
rect 111 107 112 108
rect 110 107 111 108
rect 109 107 110 108
rect 108 107 109 108
rect 107 107 108 108
rect 106 107 107 108
rect 105 107 106 108
rect 104 107 105 108
rect 103 107 104 108
rect 102 107 103 108
rect 101 107 102 108
rect 100 107 101 108
rect 99 107 100 108
rect 98 107 99 108
rect 97 107 98 108
rect 96 107 97 108
rect 95 107 96 108
rect 94 107 95 108
rect 93 107 94 108
rect 92 107 93 108
rect 91 107 92 108
rect 90 107 91 108
rect 89 107 90 108
rect 88 107 89 108
rect 87 107 88 108
rect 86 107 87 108
rect 85 107 86 108
rect 84 107 85 108
rect 83 107 84 108
rect 82 107 83 108
rect 81 107 82 108
rect 80 107 81 108
rect 62 107 63 108
rect 61 107 62 108
rect 60 107 61 108
rect 59 107 60 108
rect 58 107 59 108
rect 57 107 58 108
rect 56 107 57 108
rect 55 107 56 108
rect 54 107 55 108
rect 53 107 54 108
rect 52 107 53 108
rect 51 107 52 108
rect 50 107 51 108
rect 49 107 50 108
rect 48 107 49 108
rect 47 107 48 108
rect 46 107 47 108
rect 45 107 46 108
rect 44 107 45 108
rect 43 107 44 108
rect 42 107 43 108
rect 41 107 42 108
rect 40 107 41 108
rect 39 107 40 108
rect 38 107 39 108
rect 37 107 38 108
rect 36 107 37 108
rect 432 108 433 109
rect 431 108 432 109
rect 430 108 431 109
rect 429 108 430 109
rect 428 108 429 109
rect 427 108 428 109
rect 426 108 427 109
rect 425 108 426 109
rect 424 108 425 109
rect 423 108 424 109
rect 422 108 423 109
rect 421 108 422 109
rect 420 108 421 109
rect 419 108 420 109
rect 418 108 419 109
rect 417 108 418 109
rect 416 108 417 109
rect 415 108 416 109
rect 414 108 415 109
rect 413 108 414 109
rect 412 108 413 109
rect 411 108 412 109
rect 410 108 411 109
rect 409 108 410 109
rect 408 108 409 109
rect 407 108 408 109
rect 406 108 407 109
rect 405 108 406 109
rect 404 108 405 109
rect 403 108 404 109
rect 402 108 403 109
rect 401 108 402 109
rect 400 108 401 109
rect 399 108 400 109
rect 398 108 399 109
rect 397 108 398 109
rect 396 108 397 109
rect 395 108 396 109
rect 394 108 395 109
rect 393 108 394 109
rect 273 108 274 109
rect 272 108 273 109
rect 271 108 272 109
rect 270 108 271 109
rect 269 108 270 109
rect 268 108 269 109
rect 267 108 268 109
rect 266 108 267 109
rect 265 108 266 109
rect 264 108 265 109
rect 263 108 264 109
rect 262 108 263 109
rect 261 108 262 109
rect 260 108 261 109
rect 259 108 260 109
rect 258 108 259 109
rect 257 108 258 109
rect 256 108 257 109
rect 255 108 256 109
rect 254 108 255 109
rect 253 108 254 109
rect 252 108 253 109
rect 251 108 252 109
rect 250 108 251 109
rect 249 108 250 109
rect 248 108 249 109
rect 247 108 248 109
rect 246 108 247 109
rect 245 108 246 109
rect 244 108 245 109
rect 243 108 244 109
rect 242 108 243 109
rect 241 108 242 109
rect 240 108 241 109
rect 239 108 240 109
rect 238 108 239 109
rect 237 108 238 109
rect 236 108 237 109
rect 235 108 236 109
rect 234 108 235 109
rect 233 108 234 109
rect 232 108 233 109
rect 231 108 232 109
rect 230 108 231 109
rect 229 108 230 109
rect 228 108 229 109
rect 227 108 228 109
rect 226 108 227 109
rect 225 108 226 109
rect 224 108 225 109
rect 223 108 224 109
rect 222 108 223 109
rect 221 108 222 109
rect 220 108 221 109
rect 219 108 220 109
rect 218 108 219 109
rect 217 108 218 109
rect 216 108 217 109
rect 215 108 216 109
rect 214 108 215 109
rect 213 108 214 109
rect 212 108 213 109
rect 211 108 212 109
rect 210 108 211 109
rect 209 108 210 109
rect 208 108 209 109
rect 207 108 208 109
rect 206 108 207 109
rect 205 108 206 109
rect 204 108 205 109
rect 203 108 204 109
rect 202 108 203 109
rect 201 108 202 109
rect 200 108 201 109
rect 199 108 200 109
rect 198 108 199 109
rect 197 108 198 109
rect 196 108 197 109
rect 195 108 196 109
rect 194 108 195 109
rect 193 108 194 109
rect 192 108 193 109
rect 191 108 192 109
rect 190 108 191 109
rect 189 108 190 109
rect 188 108 189 109
rect 187 108 188 109
rect 186 108 187 109
rect 185 108 186 109
rect 184 108 185 109
rect 183 108 184 109
rect 182 108 183 109
rect 181 108 182 109
rect 180 108 181 109
rect 179 108 180 109
rect 178 108 179 109
rect 177 108 178 109
rect 176 108 177 109
rect 175 108 176 109
rect 174 108 175 109
rect 173 108 174 109
rect 172 108 173 109
rect 171 108 172 109
rect 153 108 154 109
rect 152 108 153 109
rect 151 108 152 109
rect 150 108 151 109
rect 149 108 150 109
rect 148 108 149 109
rect 147 108 148 109
rect 146 108 147 109
rect 145 108 146 109
rect 144 108 145 109
rect 143 108 144 109
rect 142 108 143 109
rect 141 108 142 109
rect 140 108 141 109
rect 139 108 140 109
rect 138 108 139 109
rect 137 108 138 109
rect 136 108 137 109
rect 135 108 136 109
rect 134 108 135 109
rect 133 108 134 109
rect 132 108 133 109
rect 131 108 132 109
rect 130 108 131 109
rect 129 108 130 109
rect 128 108 129 109
rect 127 108 128 109
rect 126 108 127 109
rect 125 108 126 109
rect 124 108 125 109
rect 123 108 124 109
rect 116 108 117 109
rect 115 108 116 109
rect 114 108 115 109
rect 113 108 114 109
rect 112 108 113 109
rect 111 108 112 109
rect 110 108 111 109
rect 109 108 110 109
rect 108 108 109 109
rect 107 108 108 109
rect 106 108 107 109
rect 105 108 106 109
rect 104 108 105 109
rect 103 108 104 109
rect 102 108 103 109
rect 101 108 102 109
rect 100 108 101 109
rect 99 108 100 109
rect 98 108 99 109
rect 97 108 98 109
rect 96 108 97 109
rect 95 108 96 109
rect 94 108 95 109
rect 93 108 94 109
rect 92 108 93 109
rect 91 108 92 109
rect 90 108 91 109
rect 89 108 90 109
rect 88 108 89 109
rect 87 108 88 109
rect 86 108 87 109
rect 85 108 86 109
rect 84 108 85 109
rect 83 108 84 109
rect 82 108 83 109
rect 81 108 82 109
rect 80 108 81 109
rect 62 108 63 109
rect 61 108 62 109
rect 60 108 61 109
rect 59 108 60 109
rect 58 108 59 109
rect 57 108 58 109
rect 56 108 57 109
rect 55 108 56 109
rect 54 108 55 109
rect 53 108 54 109
rect 52 108 53 109
rect 51 108 52 109
rect 50 108 51 109
rect 49 108 50 109
rect 48 108 49 109
rect 47 108 48 109
rect 46 108 47 109
rect 45 108 46 109
rect 44 108 45 109
rect 43 108 44 109
rect 42 108 43 109
rect 41 108 42 109
rect 40 108 41 109
rect 39 108 40 109
rect 38 108 39 109
rect 37 108 38 109
rect 36 108 37 109
rect 35 108 36 109
rect 478 109 479 110
rect 458 109 459 110
rect 433 109 434 110
rect 432 109 433 110
rect 431 109 432 110
rect 430 109 431 110
rect 429 109 430 110
rect 428 109 429 110
rect 427 109 428 110
rect 426 109 427 110
rect 425 109 426 110
rect 424 109 425 110
rect 423 109 424 110
rect 422 109 423 110
rect 421 109 422 110
rect 420 109 421 110
rect 419 109 420 110
rect 418 109 419 110
rect 417 109 418 110
rect 416 109 417 110
rect 415 109 416 110
rect 414 109 415 110
rect 413 109 414 110
rect 412 109 413 110
rect 411 109 412 110
rect 410 109 411 110
rect 409 109 410 110
rect 408 109 409 110
rect 407 109 408 110
rect 406 109 407 110
rect 405 109 406 110
rect 404 109 405 110
rect 403 109 404 110
rect 402 109 403 110
rect 401 109 402 110
rect 400 109 401 110
rect 399 109 400 110
rect 398 109 399 110
rect 397 109 398 110
rect 396 109 397 110
rect 395 109 396 110
rect 394 109 395 110
rect 393 109 394 110
rect 274 109 275 110
rect 273 109 274 110
rect 272 109 273 110
rect 271 109 272 110
rect 270 109 271 110
rect 269 109 270 110
rect 268 109 269 110
rect 267 109 268 110
rect 266 109 267 110
rect 265 109 266 110
rect 264 109 265 110
rect 263 109 264 110
rect 262 109 263 110
rect 261 109 262 110
rect 260 109 261 110
rect 259 109 260 110
rect 258 109 259 110
rect 257 109 258 110
rect 256 109 257 110
rect 255 109 256 110
rect 254 109 255 110
rect 253 109 254 110
rect 252 109 253 110
rect 251 109 252 110
rect 250 109 251 110
rect 249 109 250 110
rect 248 109 249 110
rect 247 109 248 110
rect 246 109 247 110
rect 245 109 246 110
rect 244 109 245 110
rect 243 109 244 110
rect 242 109 243 110
rect 241 109 242 110
rect 240 109 241 110
rect 239 109 240 110
rect 238 109 239 110
rect 237 109 238 110
rect 236 109 237 110
rect 235 109 236 110
rect 234 109 235 110
rect 233 109 234 110
rect 232 109 233 110
rect 231 109 232 110
rect 230 109 231 110
rect 229 109 230 110
rect 228 109 229 110
rect 227 109 228 110
rect 226 109 227 110
rect 225 109 226 110
rect 224 109 225 110
rect 223 109 224 110
rect 222 109 223 110
rect 221 109 222 110
rect 220 109 221 110
rect 219 109 220 110
rect 218 109 219 110
rect 217 109 218 110
rect 216 109 217 110
rect 215 109 216 110
rect 214 109 215 110
rect 213 109 214 110
rect 212 109 213 110
rect 211 109 212 110
rect 210 109 211 110
rect 209 109 210 110
rect 208 109 209 110
rect 207 109 208 110
rect 206 109 207 110
rect 205 109 206 110
rect 204 109 205 110
rect 203 109 204 110
rect 202 109 203 110
rect 201 109 202 110
rect 200 109 201 110
rect 199 109 200 110
rect 198 109 199 110
rect 197 109 198 110
rect 196 109 197 110
rect 195 109 196 110
rect 194 109 195 110
rect 193 109 194 110
rect 192 109 193 110
rect 191 109 192 110
rect 190 109 191 110
rect 189 109 190 110
rect 188 109 189 110
rect 187 109 188 110
rect 186 109 187 110
rect 185 109 186 110
rect 184 109 185 110
rect 183 109 184 110
rect 182 109 183 110
rect 181 109 182 110
rect 180 109 181 110
rect 179 109 180 110
rect 178 109 179 110
rect 177 109 178 110
rect 176 109 177 110
rect 175 109 176 110
rect 174 109 175 110
rect 173 109 174 110
rect 172 109 173 110
rect 171 109 172 110
rect 153 109 154 110
rect 152 109 153 110
rect 151 109 152 110
rect 150 109 151 110
rect 149 109 150 110
rect 148 109 149 110
rect 147 109 148 110
rect 146 109 147 110
rect 145 109 146 110
rect 144 109 145 110
rect 143 109 144 110
rect 142 109 143 110
rect 141 109 142 110
rect 140 109 141 110
rect 139 109 140 110
rect 138 109 139 110
rect 137 109 138 110
rect 136 109 137 110
rect 135 109 136 110
rect 134 109 135 110
rect 133 109 134 110
rect 132 109 133 110
rect 131 109 132 110
rect 130 109 131 110
rect 129 109 130 110
rect 128 109 129 110
rect 127 109 128 110
rect 126 109 127 110
rect 125 109 126 110
rect 124 109 125 110
rect 123 109 124 110
rect 122 109 123 110
rect 121 109 122 110
rect 118 109 119 110
rect 117 109 118 110
rect 116 109 117 110
rect 115 109 116 110
rect 114 109 115 110
rect 113 109 114 110
rect 112 109 113 110
rect 111 109 112 110
rect 110 109 111 110
rect 109 109 110 110
rect 108 109 109 110
rect 107 109 108 110
rect 106 109 107 110
rect 105 109 106 110
rect 104 109 105 110
rect 103 109 104 110
rect 102 109 103 110
rect 101 109 102 110
rect 100 109 101 110
rect 99 109 100 110
rect 98 109 99 110
rect 97 109 98 110
rect 96 109 97 110
rect 95 109 96 110
rect 94 109 95 110
rect 93 109 94 110
rect 92 109 93 110
rect 91 109 92 110
rect 90 109 91 110
rect 89 109 90 110
rect 88 109 89 110
rect 87 109 88 110
rect 86 109 87 110
rect 85 109 86 110
rect 84 109 85 110
rect 83 109 84 110
rect 82 109 83 110
rect 81 109 82 110
rect 80 109 81 110
rect 79 109 80 110
rect 61 109 62 110
rect 60 109 61 110
rect 59 109 60 110
rect 58 109 59 110
rect 57 109 58 110
rect 56 109 57 110
rect 55 109 56 110
rect 54 109 55 110
rect 53 109 54 110
rect 52 109 53 110
rect 51 109 52 110
rect 50 109 51 110
rect 49 109 50 110
rect 48 109 49 110
rect 47 109 48 110
rect 46 109 47 110
rect 45 109 46 110
rect 44 109 45 110
rect 43 109 44 110
rect 42 109 43 110
rect 41 109 42 110
rect 40 109 41 110
rect 39 109 40 110
rect 38 109 39 110
rect 37 109 38 110
rect 36 109 37 110
rect 35 109 36 110
rect 34 109 35 110
rect 478 110 479 111
rect 458 110 459 111
rect 434 110 435 111
rect 433 110 434 111
rect 432 110 433 111
rect 431 110 432 111
rect 430 110 431 111
rect 429 110 430 111
rect 428 110 429 111
rect 427 110 428 111
rect 426 110 427 111
rect 425 110 426 111
rect 424 110 425 111
rect 423 110 424 111
rect 422 110 423 111
rect 421 110 422 111
rect 420 110 421 111
rect 419 110 420 111
rect 418 110 419 111
rect 417 110 418 111
rect 416 110 417 111
rect 415 110 416 111
rect 414 110 415 111
rect 413 110 414 111
rect 412 110 413 111
rect 411 110 412 111
rect 410 110 411 111
rect 409 110 410 111
rect 408 110 409 111
rect 407 110 408 111
rect 406 110 407 111
rect 405 110 406 111
rect 404 110 405 111
rect 403 110 404 111
rect 402 110 403 111
rect 401 110 402 111
rect 400 110 401 111
rect 399 110 400 111
rect 398 110 399 111
rect 397 110 398 111
rect 396 110 397 111
rect 395 110 396 111
rect 394 110 395 111
rect 393 110 394 111
rect 275 110 276 111
rect 274 110 275 111
rect 273 110 274 111
rect 272 110 273 111
rect 271 110 272 111
rect 270 110 271 111
rect 269 110 270 111
rect 268 110 269 111
rect 267 110 268 111
rect 266 110 267 111
rect 265 110 266 111
rect 264 110 265 111
rect 263 110 264 111
rect 262 110 263 111
rect 261 110 262 111
rect 260 110 261 111
rect 259 110 260 111
rect 258 110 259 111
rect 257 110 258 111
rect 256 110 257 111
rect 255 110 256 111
rect 254 110 255 111
rect 253 110 254 111
rect 252 110 253 111
rect 251 110 252 111
rect 250 110 251 111
rect 249 110 250 111
rect 248 110 249 111
rect 247 110 248 111
rect 246 110 247 111
rect 245 110 246 111
rect 244 110 245 111
rect 243 110 244 111
rect 242 110 243 111
rect 241 110 242 111
rect 240 110 241 111
rect 239 110 240 111
rect 238 110 239 111
rect 237 110 238 111
rect 236 110 237 111
rect 235 110 236 111
rect 234 110 235 111
rect 233 110 234 111
rect 232 110 233 111
rect 231 110 232 111
rect 230 110 231 111
rect 229 110 230 111
rect 228 110 229 111
rect 227 110 228 111
rect 226 110 227 111
rect 225 110 226 111
rect 224 110 225 111
rect 223 110 224 111
rect 222 110 223 111
rect 221 110 222 111
rect 220 110 221 111
rect 219 110 220 111
rect 218 110 219 111
rect 217 110 218 111
rect 216 110 217 111
rect 215 110 216 111
rect 214 110 215 111
rect 213 110 214 111
rect 212 110 213 111
rect 211 110 212 111
rect 210 110 211 111
rect 209 110 210 111
rect 208 110 209 111
rect 207 110 208 111
rect 206 110 207 111
rect 205 110 206 111
rect 204 110 205 111
rect 203 110 204 111
rect 202 110 203 111
rect 201 110 202 111
rect 200 110 201 111
rect 199 110 200 111
rect 198 110 199 111
rect 197 110 198 111
rect 196 110 197 111
rect 195 110 196 111
rect 194 110 195 111
rect 193 110 194 111
rect 192 110 193 111
rect 191 110 192 111
rect 190 110 191 111
rect 189 110 190 111
rect 188 110 189 111
rect 187 110 188 111
rect 186 110 187 111
rect 185 110 186 111
rect 184 110 185 111
rect 183 110 184 111
rect 182 110 183 111
rect 181 110 182 111
rect 180 110 181 111
rect 179 110 180 111
rect 178 110 179 111
rect 177 110 178 111
rect 176 110 177 111
rect 175 110 176 111
rect 174 110 175 111
rect 173 110 174 111
rect 172 110 173 111
rect 171 110 172 111
rect 170 110 171 111
rect 152 110 153 111
rect 151 110 152 111
rect 150 110 151 111
rect 149 110 150 111
rect 148 110 149 111
rect 147 110 148 111
rect 146 110 147 111
rect 145 110 146 111
rect 144 110 145 111
rect 143 110 144 111
rect 142 110 143 111
rect 141 110 142 111
rect 140 110 141 111
rect 139 110 140 111
rect 138 110 139 111
rect 137 110 138 111
rect 136 110 137 111
rect 135 110 136 111
rect 134 110 135 111
rect 133 110 134 111
rect 132 110 133 111
rect 131 110 132 111
rect 130 110 131 111
rect 129 110 130 111
rect 128 110 129 111
rect 127 110 128 111
rect 126 110 127 111
rect 125 110 126 111
rect 124 110 125 111
rect 123 110 124 111
rect 122 110 123 111
rect 121 110 122 111
rect 120 110 121 111
rect 119 110 120 111
rect 118 110 119 111
rect 117 110 118 111
rect 116 110 117 111
rect 115 110 116 111
rect 114 110 115 111
rect 113 110 114 111
rect 112 110 113 111
rect 111 110 112 111
rect 110 110 111 111
rect 109 110 110 111
rect 108 110 109 111
rect 107 110 108 111
rect 106 110 107 111
rect 105 110 106 111
rect 104 110 105 111
rect 103 110 104 111
rect 102 110 103 111
rect 101 110 102 111
rect 100 110 101 111
rect 99 110 100 111
rect 98 110 99 111
rect 97 110 98 111
rect 96 110 97 111
rect 95 110 96 111
rect 94 110 95 111
rect 93 110 94 111
rect 92 110 93 111
rect 91 110 92 111
rect 90 110 91 111
rect 89 110 90 111
rect 88 110 89 111
rect 87 110 88 111
rect 86 110 87 111
rect 85 110 86 111
rect 84 110 85 111
rect 83 110 84 111
rect 82 110 83 111
rect 81 110 82 111
rect 80 110 81 111
rect 79 110 80 111
rect 78 110 79 111
rect 77 110 78 111
rect 61 110 62 111
rect 60 110 61 111
rect 59 110 60 111
rect 58 110 59 111
rect 57 110 58 111
rect 56 110 57 111
rect 55 110 56 111
rect 54 110 55 111
rect 53 110 54 111
rect 52 110 53 111
rect 51 110 52 111
rect 50 110 51 111
rect 49 110 50 111
rect 48 110 49 111
rect 47 110 48 111
rect 46 110 47 111
rect 45 110 46 111
rect 44 110 45 111
rect 43 110 44 111
rect 42 110 43 111
rect 41 110 42 111
rect 40 110 41 111
rect 39 110 40 111
rect 38 110 39 111
rect 37 110 38 111
rect 36 110 37 111
rect 35 110 36 111
rect 34 110 35 111
rect 33 110 34 111
rect 478 111 479 112
rect 477 111 478 112
rect 459 111 460 112
rect 458 111 459 112
rect 435 111 436 112
rect 434 111 435 112
rect 433 111 434 112
rect 432 111 433 112
rect 431 111 432 112
rect 430 111 431 112
rect 429 111 430 112
rect 428 111 429 112
rect 427 111 428 112
rect 426 111 427 112
rect 425 111 426 112
rect 424 111 425 112
rect 423 111 424 112
rect 422 111 423 112
rect 421 111 422 112
rect 420 111 421 112
rect 419 111 420 112
rect 418 111 419 112
rect 417 111 418 112
rect 416 111 417 112
rect 415 111 416 112
rect 414 111 415 112
rect 413 111 414 112
rect 412 111 413 112
rect 411 111 412 112
rect 410 111 411 112
rect 409 111 410 112
rect 408 111 409 112
rect 407 111 408 112
rect 406 111 407 112
rect 405 111 406 112
rect 404 111 405 112
rect 403 111 404 112
rect 402 111 403 112
rect 401 111 402 112
rect 400 111 401 112
rect 399 111 400 112
rect 398 111 399 112
rect 397 111 398 112
rect 396 111 397 112
rect 395 111 396 112
rect 394 111 395 112
rect 393 111 394 112
rect 263 111 264 112
rect 262 111 263 112
rect 261 111 262 112
rect 260 111 261 112
rect 259 111 260 112
rect 258 111 259 112
rect 257 111 258 112
rect 256 111 257 112
rect 255 111 256 112
rect 254 111 255 112
rect 253 111 254 112
rect 252 111 253 112
rect 251 111 252 112
rect 250 111 251 112
rect 249 111 250 112
rect 248 111 249 112
rect 247 111 248 112
rect 246 111 247 112
rect 245 111 246 112
rect 244 111 245 112
rect 243 111 244 112
rect 242 111 243 112
rect 241 111 242 112
rect 240 111 241 112
rect 239 111 240 112
rect 238 111 239 112
rect 237 111 238 112
rect 236 111 237 112
rect 235 111 236 112
rect 234 111 235 112
rect 233 111 234 112
rect 232 111 233 112
rect 231 111 232 112
rect 230 111 231 112
rect 229 111 230 112
rect 228 111 229 112
rect 227 111 228 112
rect 226 111 227 112
rect 225 111 226 112
rect 224 111 225 112
rect 223 111 224 112
rect 222 111 223 112
rect 221 111 222 112
rect 220 111 221 112
rect 219 111 220 112
rect 218 111 219 112
rect 217 111 218 112
rect 216 111 217 112
rect 215 111 216 112
rect 214 111 215 112
rect 213 111 214 112
rect 212 111 213 112
rect 211 111 212 112
rect 210 111 211 112
rect 209 111 210 112
rect 208 111 209 112
rect 207 111 208 112
rect 206 111 207 112
rect 205 111 206 112
rect 204 111 205 112
rect 203 111 204 112
rect 202 111 203 112
rect 201 111 202 112
rect 200 111 201 112
rect 199 111 200 112
rect 198 111 199 112
rect 197 111 198 112
rect 196 111 197 112
rect 195 111 196 112
rect 194 111 195 112
rect 193 111 194 112
rect 192 111 193 112
rect 191 111 192 112
rect 190 111 191 112
rect 189 111 190 112
rect 188 111 189 112
rect 187 111 188 112
rect 186 111 187 112
rect 185 111 186 112
rect 184 111 185 112
rect 183 111 184 112
rect 182 111 183 112
rect 181 111 182 112
rect 180 111 181 112
rect 179 111 180 112
rect 178 111 179 112
rect 177 111 178 112
rect 176 111 177 112
rect 175 111 176 112
rect 174 111 175 112
rect 173 111 174 112
rect 172 111 173 112
rect 171 111 172 112
rect 170 111 171 112
rect 152 111 153 112
rect 151 111 152 112
rect 150 111 151 112
rect 149 111 150 112
rect 148 111 149 112
rect 147 111 148 112
rect 146 111 147 112
rect 145 111 146 112
rect 144 111 145 112
rect 143 111 144 112
rect 142 111 143 112
rect 141 111 142 112
rect 140 111 141 112
rect 139 111 140 112
rect 138 111 139 112
rect 137 111 138 112
rect 136 111 137 112
rect 135 111 136 112
rect 134 111 135 112
rect 133 111 134 112
rect 132 111 133 112
rect 131 111 132 112
rect 130 111 131 112
rect 129 111 130 112
rect 128 111 129 112
rect 127 111 128 112
rect 126 111 127 112
rect 125 111 126 112
rect 124 111 125 112
rect 123 111 124 112
rect 122 111 123 112
rect 121 111 122 112
rect 120 111 121 112
rect 119 111 120 112
rect 118 111 119 112
rect 117 111 118 112
rect 116 111 117 112
rect 115 111 116 112
rect 114 111 115 112
rect 113 111 114 112
rect 112 111 113 112
rect 111 111 112 112
rect 110 111 111 112
rect 109 111 110 112
rect 108 111 109 112
rect 107 111 108 112
rect 106 111 107 112
rect 105 111 106 112
rect 104 111 105 112
rect 103 111 104 112
rect 102 111 103 112
rect 101 111 102 112
rect 100 111 101 112
rect 99 111 100 112
rect 98 111 99 112
rect 97 111 98 112
rect 96 111 97 112
rect 95 111 96 112
rect 94 111 95 112
rect 93 111 94 112
rect 92 111 93 112
rect 91 111 92 112
rect 90 111 91 112
rect 89 111 90 112
rect 88 111 89 112
rect 87 111 88 112
rect 86 111 87 112
rect 85 111 86 112
rect 84 111 85 112
rect 83 111 84 112
rect 82 111 83 112
rect 81 111 82 112
rect 80 111 81 112
rect 79 111 80 112
rect 78 111 79 112
rect 77 111 78 112
rect 76 111 77 112
rect 75 111 76 112
rect 61 111 62 112
rect 60 111 61 112
rect 59 111 60 112
rect 58 111 59 112
rect 57 111 58 112
rect 56 111 57 112
rect 55 111 56 112
rect 54 111 55 112
rect 53 111 54 112
rect 52 111 53 112
rect 51 111 52 112
rect 50 111 51 112
rect 49 111 50 112
rect 48 111 49 112
rect 47 111 48 112
rect 46 111 47 112
rect 45 111 46 112
rect 44 111 45 112
rect 43 111 44 112
rect 42 111 43 112
rect 41 111 42 112
rect 40 111 41 112
rect 39 111 40 112
rect 38 111 39 112
rect 37 111 38 112
rect 36 111 37 112
rect 35 111 36 112
rect 34 111 35 112
rect 33 111 34 112
rect 32 111 33 112
rect 478 112 479 113
rect 477 112 478 113
rect 476 112 477 113
rect 475 112 476 113
rect 474 112 475 113
rect 473 112 474 113
rect 472 112 473 113
rect 471 112 472 113
rect 470 112 471 113
rect 469 112 470 113
rect 468 112 469 113
rect 467 112 468 113
rect 466 112 467 113
rect 465 112 466 113
rect 464 112 465 113
rect 463 112 464 113
rect 462 112 463 113
rect 461 112 462 113
rect 460 112 461 113
rect 459 112 460 113
rect 458 112 459 113
rect 436 112 437 113
rect 435 112 436 113
rect 434 112 435 113
rect 433 112 434 113
rect 432 112 433 113
rect 431 112 432 113
rect 430 112 431 113
rect 429 112 430 113
rect 428 112 429 113
rect 427 112 428 113
rect 426 112 427 113
rect 425 112 426 113
rect 424 112 425 113
rect 423 112 424 113
rect 422 112 423 113
rect 421 112 422 113
rect 420 112 421 113
rect 419 112 420 113
rect 418 112 419 113
rect 417 112 418 113
rect 416 112 417 113
rect 415 112 416 113
rect 414 112 415 113
rect 413 112 414 113
rect 412 112 413 113
rect 411 112 412 113
rect 410 112 411 113
rect 409 112 410 113
rect 408 112 409 113
rect 407 112 408 113
rect 406 112 407 113
rect 405 112 406 113
rect 404 112 405 113
rect 403 112 404 113
rect 402 112 403 113
rect 401 112 402 113
rect 400 112 401 113
rect 399 112 400 113
rect 398 112 399 113
rect 397 112 398 113
rect 396 112 397 113
rect 395 112 396 113
rect 394 112 395 113
rect 393 112 394 113
rect 255 112 256 113
rect 254 112 255 113
rect 253 112 254 113
rect 252 112 253 113
rect 251 112 252 113
rect 250 112 251 113
rect 249 112 250 113
rect 248 112 249 113
rect 247 112 248 113
rect 246 112 247 113
rect 245 112 246 113
rect 244 112 245 113
rect 243 112 244 113
rect 242 112 243 113
rect 241 112 242 113
rect 240 112 241 113
rect 239 112 240 113
rect 238 112 239 113
rect 237 112 238 113
rect 236 112 237 113
rect 235 112 236 113
rect 234 112 235 113
rect 233 112 234 113
rect 232 112 233 113
rect 231 112 232 113
rect 230 112 231 113
rect 229 112 230 113
rect 228 112 229 113
rect 227 112 228 113
rect 226 112 227 113
rect 225 112 226 113
rect 224 112 225 113
rect 223 112 224 113
rect 222 112 223 113
rect 221 112 222 113
rect 220 112 221 113
rect 219 112 220 113
rect 218 112 219 113
rect 217 112 218 113
rect 216 112 217 113
rect 215 112 216 113
rect 214 112 215 113
rect 213 112 214 113
rect 212 112 213 113
rect 211 112 212 113
rect 210 112 211 113
rect 209 112 210 113
rect 208 112 209 113
rect 207 112 208 113
rect 206 112 207 113
rect 205 112 206 113
rect 204 112 205 113
rect 203 112 204 113
rect 202 112 203 113
rect 201 112 202 113
rect 200 112 201 113
rect 199 112 200 113
rect 198 112 199 113
rect 197 112 198 113
rect 196 112 197 113
rect 195 112 196 113
rect 194 112 195 113
rect 193 112 194 113
rect 192 112 193 113
rect 191 112 192 113
rect 190 112 191 113
rect 189 112 190 113
rect 188 112 189 113
rect 187 112 188 113
rect 186 112 187 113
rect 185 112 186 113
rect 184 112 185 113
rect 183 112 184 113
rect 182 112 183 113
rect 181 112 182 113
rect 180 112 181 113
rect 179 112 180 113
rect 178 112 179 113
rect 177 112 178 113
rect 176 112 177 113
rect 175 112 176 113
rect 174 112 175 113
rect 173 112 174 113
rect 172 112 173 113
rect 171 112 172 113
rect 170 112 171 113
rect 169 112 170 113
rect 151 112 152 113
rect 150 112 151 113
rect 149 112 150 113
rect 148 112 149 113
rect 147 112 148 113
rect 146 112 147 113
rect 145 112 146 113
rect 144 112 145 113
rect 143 112 144 113
rect 142 112 143 113
rect 141 112 142 113
rect 140 112 141 113
rect 139 112 140 113
rect 138 112 139 113
rect 137 112 138 113
rect 136 112 137 113
rect 135 112 136 113
rect 134 112 135 113
rect 133 112 134 113
rect 132 112 133 113
rect 131 112 132 113
rect 130 112 131 113
rect 129 112 130 113
rect 128 112 129 113
rect 127 112 128 113
rect 126 112 127 113
rect 125 112 126 113
rect 124 112 125 113
rect 123 112 124 113
rect 122 112 123 113
rect 121 112 122 113
rect 120 112 121 113
rect 119 112 120 113
rect 118 112 119 113
rect 117 112 118 113
rect 116 112 117 113
rect 115 112 116 113
rect 114 112 115 113
rect 113 112 114 113
rect 112 112 113 113
rect 111 112 112 113
rect 110 112 111 113
rect 109 112 110 113
rect 108 112 109 113
rect 107 112 108 113
rect 106 112 107 113
rect 105 112 106 113
rect 104 112 105 113
rect 103 112 104 113
rect 102 112 103 113
rect 101 112 102 113
rect 100 112 101 113
rect 99 112 100 113
rect 98 112 99 113
rect 97 112 98 113
rect 96 112 97 113
rect 95 112 96 113
rect 94 112 95 113
rect 93 112 94 113
rect 92 112 93 113
rect 91 112 92 113
rect 90 112 91 113
rect 89 112 90 113
rect 88 112 89 113
rect 87 112 88 113
rect 86 112 87 113
rect 85 112 86 113
rect 84 112 85 113
rect 83 112 84 113
rect 82 112 83 113
rect 81 112 82 113
rect 80 112 81 113
rect 79 112 80 113
rect 78 112 79 113
rect 77 112 78 113
rect 76 112 77 113
rect 75 112 76 113
rect 74 112 75 113
rect 73 112 74 113
rect 60 112 61 113
rect 59 112 60 113
rect 58 112 59 113
rect 57 112 58 113
rect 56 112 57 113
rect 55 112 56 113
rect 54 112 55 113
rect 53 112 54 113
rect 52 112 53 113
rect 51 112 52 113
rect 50 112 51 113
rect 49 112 50 113
rect 48 112 49 113
rect 47 112 48 113
rect 46 112 47 113
rect 45 112 46 113
rect 44 112 45 113
rect 43 112 44 113
rect 42 112 43 113
rect 41 112 42 113
rect 40 112 41 113
rect 39 112 40 113
rect 38 112 39 113
rect 37 112 38 113
rect 36 112 37 113
rect 35 112 36 113
rect 34 112 35 113
rect 33 112 34 113
rect 32 112 33 113
rect 31 112 32 113
rect 478 113 479 114
rect 477 113 478 114
rect 476 113 477 114
rect 475 113 476 114
rect 474 113 475 114
rect 473 113 474 114
rect 472 113 473 114
rect 471 113 472 114
rect 470 113 471 114
rect 469 113 470 114
rect 468 113 469 114
rect 467 113 468 114
rect 466 113 467 114
rect 465 113 466 114
rect 464 113 465 114
rect 463 113 464 114
rect 462 113 463 114
rect 461 113 462 114
rect 460 113 461 114
rect 459 113 460 114
rect 458 113 459 114
rect 436 113 437 114
rect 435 113 436 114
rect 434 113 435 114
rect 433 113 434 114
rect 432 113 433 114
rect 431 113 432 114
rect 430 113 431 114
rect 429 113 430 114
rect 428 113 429 114
rect 427 113 428 114
rect 426 113 427 114
rect 425 113 426 114
rect 424 113 425 114
rect 423 113 424 114
rect 422 113 423 114
rect 421 113 422 114
rect 420 113 421 114
rect 419 113 420 114
rect 418 113 419 114
rect 417 113 418 114
rect 416 113 417 114
rect 415 113 416 114
rect 414 113 415 114
rect 413 113 414 114
rect 412 113 413 114
rect 411 113 412 114
rect 410 113 411 114
rect 409 113 410 114
rect 408 113 409 114
rect 407 113 408 114
rect 406 113 407 114
rect 405 113 406 114
rect 404 113 405 114
rect 403 113 404 114
rect 402 113 403 114
rect 401 113 402 114
rect 400 113 401 114
rect 399 113 400 114
rect 398 113 399 114
rect 397 113 398 114
rect 396 113 397 114
rect 395 113 396 114
rect 394 113 395 114
rect 393 113 394 114
rect 251 113 252 114
rect 250 113 251 114
rect 249 113 250 114
rect 248 113 249 114
rect 247 113 248 114
rect 246 113 247 114
rect 245 113 246 114
rect 244 113 245 114
rect 243 113 244 114
rect 242 113 243 114
rect 241 113 242 114
rect 240 113 241 114
rect 239 113 240 114
rect 238 113 239 114
rect 237 113 238 114
rect 236 113 237 114
rect 235 113 236 114
rect 234 113 235 114
rect 233 113 234 114
rect 232 113 233 114
rect 231 113 232 114
rect 230 113 231 114
rect 229 113 230 114
rect 228 113 229 114
rect 227 113 228 114
rect 226 113 227 114
rect 225 113 226 114
rect 224 113 225 114
rect 223 113 224 114
rect 222 113 223 114
rect 221 113 222 114
rect 220 113 221 114
rect 219 113 220 114
rect 218 113 219 114
rect 217 113 218 114
rect 216 113 217 114
rect 215 113 216 114
rect 214 113 215 114
rect 213 113 214 114
rect 212 113 213 114
rect 211 113 212 114
rect 210 113 211 114
rect 209 113 210 114
rect 208 113 209 114
rect 207 113 208 114
rect 206 113 207 114
rect 205 113 206 114
rect 204 113 205 114
rect 203 113 204 114
rect 202 113 203 114
rect 201 113 202 114
rect 200 113 201 114
rect 199 113 200 114
rect 198 113 199 114
rect 197 113 198 114
rect 196 113 197 114
rect 195 113 196 114
rect 194 113 195 114
rect 193 113 194 114
rect 192 113 193 114
rect 191 113 192 114
rect 190 113 191 114
rect 189 113 190 114
rect 188 113 189 114
rect 187 113 188 114
rect 186 113 187 114
rect 185 113 186 114
rect 184 113 185 114
rect 183 113 184 114
rect 182 113 183 114
rect 181 113 182 114
rect 180 113 181 114
rect 179 113 180 114
rect 178 113 179 114
rect 177 113 178 114
rect 176 113 177 114
rect 175 113 176 114
rect 174 113 175 114
rect 173 113 174 114
rect 172 113 173 114
rect 171 113 172 114
rect 170 113 171 114
rect 169 113 170 114
rect 151 113 152 114
rect 150 113 151 114
rect 149 113 150 114
rect 148 113 149 114
rect 147 113 148 114
rect 146 113 147 114
rect 145 113 146 114
rect 144 113 145 114
rect 143 113 144 114
rect 142 113 143 114
rect 141 113 142 114
rect 140 113 141 114
rect 139 113 140 114
rect 138 113 139 114
rect 137 113 138 114
rect 136 113 137 114
rect 135 113 136 114
rect 134 113 135 114
rect 133 113 134 114
rect 132 113 133 114
rect 131 113 132 114
rect 130 113 131 114
rect 129 113 130 114
rect 128 113 129 114
rect 127 113 128 114
rect 126 113 127 114
rect 125 113 126 114
rect 124 113 125 114
rect 123 113 124 114
rect 122 113 123 114
rect 121 113 122 114
rect 120 113 121 114
rect 119 113 120 114
rect 118 113 119 114
rect 117 113 118 114
rect 116 113 117 114
rect 115 113 116 114
rect 114 113 115 114
rect 113 113 114 114
rect 112 113 113 114
rect 111 113 112 114
rect 110 113 111 114
rect 109 113 110 114
rect 108 113 109 114
rect 107 113 108 114
rect 106 113 107 114
rect 105 113 106 114
rect 104 113 105 114
rect 103 113 104 114
rect 102 113 103 114
rect 101 113 102 114
rect 100 113 101 114
rect 99 113 100 114
rect 98 113 99 114
rect 97 113 98 114
rect 96 113 97 114
rect 95 113 96 114
rect 94 113 95 114
rect 93 113 94 114
rect 92 113 93 114
rect 91 113 92 114
rect 90 113 91 114
rect 89 113 90 114
rect 88 113 89 114
rect 87 113 88 114
rect 86 113 87 114
rect 85 113 86 114
rect 84 113 85 114
rect 83 113 84 114
rect 82 113 83 114
rect 81 113 82 114
rect 80 113 81 114
rect 79 113 80 114
rect 78 113 79 114
rect 77 113 78 114
rect 76 113 77 114
rect 75 113 76 114
rect 74 113 75 114
rect 73 113 74 114
rect 72 113 73 114
rect 60 113 61 114
rect 59 113 60 114
rect 58 113 59 114
rect 57 113 58 114
rect 56 113 57 114
rect 55 113 56 114
rect 54 113 55 114
rect 53 113 54 114
rect 52 113 53 114
rect 51 113 52 114
rect 50 113 51 114
rect 49 113 50 114
rect 48 113 49 114
rect 47 113 48 114
rect 46 113 47 114
rect 45 113 46 114
rect 44 113 45 114
rect 43 113 44 114
rect 42 113 43 114
rect 41 113 42 114
rect 40 113 41 114
rect 39 113 40 114
rect 38 113 39 114
rect 37 113 38 114
rect 36 113 37 114
rect 35 113 36 114
rect 34 113 35 114
rect 33 113 34 114
rect 32 113 33 114
rect 31 113 32 114
rect 30 113 31 114
rect 478 114 479 115
rect 477 114 478 115
rect 476 114 477 115
rect 463 114 464 115
rect 462 114 463 115
rect 461 114 462 115
rect 460 114 461 115
rect 459 114 460 115
rect 458 114 459 115
rect 437 114 438 115
rect 436 114 437 115
rect 435 114 436 115
rect 434 114 435 115
rect 433 114 434 115
rect 432 114 433 115
rect 431 114 432 115
rect 430 114 431 115
rect 429 114 430 115
rect 428 114 429 115
rect 427 114 428 115
rect 426 114 427 115
rect 425 114 426 115
rect 424 114 425 115
rect 423 114 424 115
rect 422 114 423 115
rect 421 114 422 115
rect 420 114 421 115
rect 419 114 420 115
rect 418 114 419 115
rect 417 114 418 115
rect 416 114 417 115
rect 415 114 416 115
rect 414 114 415 115
rect 413 114 414 115
rect 412 114 413 115
rect 411 114 412 115
rect 410 114 411 115
rect 409 114 410 115
rect 408 114 409 115
rect 407 114 408 115
rect 406 114 407 115
rect 405 114 406 115
rect 404 114 405 115
rect 403 114 404 115
rect 402 114 403 115
rect 401 114 402 115
rect 400 114 401 115
rect 399 114 400 115
rect 398 114 399 115
rect 397 114 398 115
rect 396 114 397 115
rect 395 114 396 115
rect 394 114 395 115
rect 393 114 394 115
rect 247 114 248 115
rect 246 114 247 115
rect 245 114 246 115
rect 244 114 245 115
rect 243 114 244 115
rect 242 114 243 115
rect 241 114 242 115
rect 240 114 241 115
rect 239 114 240 115
rect 238 114 239 115
rect 237 114 238 115
rect 236 114 237 115
rect 235 114 236 115
rect 234 114 235 115
rect 233 114 234 115
rect 232 114 233 115
rect 231 114 232 115
rect 230 114 231 115
rect 229 114 230 115
rect 228 114 229 115
rect 227 114 228 115
rect 226 114 227 115
rect 225 114 226 115
rect 224 114 225 115
rect 223 114 224 115
rect 222 114 223 115
rect 221 114 222 115
rect 220 114 221 115
rect 219 114 220 115
rect 218 114 219 115
rect 217 114 218 115
rect 216 114 217 115
rect 215 114 216 115
rect 214 114 215 115
rect 213 114 214 115
rect 212 114 213 115
rect 211 114 212 115
rect 210 114 211 115
rect 209 114 210 115
rect 208 114 209 115
rect 207 114 208 115
rect 206 114 207 115
rect 205 114 206 115
rect 204 114 205 115
rect 203 114 204 115
rect 202 114 203 115
rect 201 114 202 115
rect 200 114 201 115
rect 199 114 200 115
rect 198 114 199 115
rect 197 114 198 115
rect 196 114 197 115
rect 195 114 196 115
rect 194 114 195 115
rect 193 114 194 115
rect 192 114 193 115
rect 191 114 192 115
rect 190 114 191 115
rect 189 114 190 115
rect 188 114 189 115
rect 187 114 188 115
rect 186 114 187 115
rect 185 114 186 115
rect 184 114 185 115
rect 183 114 184 115
rect 182 114 183 115
rect 181 114 182 115
rect 180 114 181 115
rect 179 114 180 115
rect 178 114 179 115
rect 177 114 178 115
rect 176 114 177 115
rect 175 114 176 115
rect 174 114 175 115
rect 173 114 174 115
rect 172 114 173 115
rect 171 114 172 115
rect 170 114 171 115
rect 169 114 170 115
rect 168 114 169 115
rect 151 114 152 115
rect 150 114 151 115
rect 149 114 150 115
rect 148 114 149 115
rect 147 114 148 115
rect 146 114 147 115
rect 145 114 146 115
rect 144 114 145 115
rect 143 114 144 115
rect 142 114 143 115
rect 141 114 142 115
rect 140 114 141 115
rect 139 114 140 115
rect 138 114 139 115
rect 137 114 138 115
rect 136 114 137 115
rect 135 114 136 115
rect 134 114 135 115
rect 133 114 134 115
rect 132 114 133 115
rect 131 114 132 115
rect 130 114 131 115
rect 129 114 130 115
rect 128 114 129 115
rect 127 114 128 115
rect 126 114 127 115
rect 125 114 126 115
rect 124 114 125 115
rect 123 114 124 115
rect 122 114 123 115
rect 121 114 122 115
rect 120 114 121 115
rect 119 114 120 115
rect 118 114 119 115
rect 117 114 118 115
rect 116 114 117 115
rect 115 114 116 115
rect 114 114 115 115
rect 113 114 114 115
rect 112 114 113 115
rect 111 114 112 115
rect 110 114 111 115
rect 109 114 110 115
rect 108 114 109 115
rect 107 114 108 115
rect 106 114 107 115
rect 105 114 106 115
rect 104 114 105 115
rect 103 114 104 115
rect 102 114 103 115
rect 101 114 102 115
rect 100 114 101 115
rect 99 114 100 115
rect 98 114 99 115
rect 97 114 98 115
rect 96 114 97 115
rect 95 114 96 115
rect 94 114 95 115
rect 93 114 94 115
rect 92 114 93 115
rect 91 114 92 115
rect 90 114 91 115
rect 89 114 90 115
rect 88 114 89 115
rect 87 114 88 115
rect 86 114 87 115
rect 85 114 86 115
rect 84 114 85 115
rect 83 114 84 115
rect 82 114 83 115
rect 81 114 82 115
rect 80 114 81 115
rect 79 114 80 115
rect 78 114 79 115
rect 77 114 78 115
rect 76 114 77 115
rect 75 114 76 115
rect 74 114 75 115
rect 73 114 74 115
rect 72 114 73 115
rect 71 114 72 115
rect 60 114 61 115
rect 59 114 60 115
rect 58 114 59 115
rect 57 114 58 115
rect 56 114 57 115
rect 55 114 56 115
rect 54 114 55 115
rect 53 114 54 115
rect 52 114 53 115
rect 51 114 52 115
rect 50 114 51 115
rect 49 114 50 115
rect 48 114 49 115
rect 47 114 48 115
rect 46 114 47 115
rect 45 114 46 115
rect 44 114 45 115
rect 43 114 44 115
rect 42 114 43 115
rect 41 114 42 115
rect 40 114 41 115
rect 39 114 40 115
rect 38 114 39 115
rect 37 114 38 115
rect 36 114 37 115
rect 35 114 36 115
rect 34 114 35 115
rect 33 114 34 115
rect 32 114 33 115
rect 31 114 32 115
rect 30 114 31 115
rect 478 115 479 116
rect 464 115 465 116
rect 463 115 464 116
rect 462 115 463 116
rect 461 115 462 116
rect 460 115 461 116
rect 459 115 460 116
rect 458 115 459 116
rect 437 115 438 116
rect 436 115 437 116
rect 435 115 436 116
rect 434 115 435 116
rect 433 115 434 116
rect 432 115 433 116
rect 431 115 432 116
rect 430 115 431 116
rect 429 115 430 116
rect 428 115 429 116
rect 427 115 428 116
rect 426 115 427 116
rect 425 115 426 116
rect 424 115 425 116
rect 397 115 398 116
rect 396 115 397 116
rect 395 115 396 116
rect 394 115 395 116
rect 393 115 394 116
rect 244 115 245 116
rect 243 115 244 116
rect 242 115 243 116
rect 241 115 242 116
rect 240 115 241 116
rect 239 115 240 116
rect 238 115 239 116
rect 237 115 238 116
rect 236 115 237 116
rect 235 115 236 116
rect 234 115 235 116
rect 233 115 234 116
rect 232 115 233 116
rect 231 115 232 116
rect 230 115 231 116
rect 229 115 230 116
rect 228 115 229 116
rect 227 115 228 116
rect 226 115 227 116
rect 225 115 226 116
rect 224 115 225 116
rect 223 115 224 116
rect 222 115 223 116
rect 221 115 222 116
rect 220 115 221 116
rect 219 115 220 116
rect 218 115 219 116
rect 217 115 218 116
rect 216 115 217 116
rect 215 115 216 116
rect 214 115 215 116
rect 213 115 214 116
rect 212 115 213 116
rect 211 115 212 116
rect 210 115 211 116
rect 209 115 210 116
rect 208 115 209 116
rect 207 115 208 116
rect 206 115 207 116
rect 205 115 206 116
rect 204 115 205 116
rect 203 115 204 116
rect 202 115 203 116
rect 201 115 202 116
rect 200 115 201 116
rect 199 115 200 116
rect 198 115 199 116
rect 197 115 198 116
rect 196 115 197 116
rect 195 115 196 116
rect 194 115 195 116
rect 193 115 194 116
rect 192 115 193 116
rect 191 115 192 116
rect 190 115 191 116
rect 189 115 190 116
rect 188 115 189 116
rect 187 115 188 116
rect 186 115 187 116
rect 185 115 186 116
rect 184 115 185 116
rect 183 115 184 116
rect 182 115 183 116
rect 181 115 182 116
rect 180 115 181 116
rect 179 115 180 116
rect 178 115 179 116
rect 177 115 178 116
rect 176 115 177 116
rect 175 115 176 116
rect 174 115 175 116
rect 173 115 174 116
rect 172 115 173 116
rect 171 115 172 116
rect 170 115 171 116
rect 169 115 170 116
rect 168 115 169 116
rect 150 115 151 116
rect 149 115 150 116
rect 148 115 149 116
rect 147 115 148 116
rect 146 115 147 116
rect 145 115 146 116
rect 144 115 145 116
rect 143 115 144 116
rect 142 115 143 116
rect 141 115 142 116
rect 140 115 141 116
rect 139 115 140 116
rect 138 115 139 116
rect 137 115 138 116
rect 136 115 137 116
rect 135 115 136 116
rect 134 115 135 116
rect 133 115 134 116
rect 132 115 133 116
rect 131 115 132 116
rect 130 115 131 116
rect 129 115 130 116
rect 128 115 129 116
rect 127 115 128 116
rect 126 115 127 116
rect 125 115 126 116
rect 124 115 125 116
rect 123 115 124 116
rect 122 115 123 116
rect 121 115 122 116
rect 120 115 121 116
rect 119 115 120 116
rect 118 115 119 116
rect 117 115 118 116
rect 116 115 117 116
rect 115 115 116 116
rect 114 115 115 116
rect 113 115 114 116
rect 112 115 113 116
rect 111 115 112 116
rect 110 115 111 116
rect 109 115 110 116
rect 108 115 109 116
rect 107 115 108 116
rect 106 115 107 116
rect 105 115 106 116
rect 104 115 105 116
rect 103 115 104 116
rect 102 115 103 116
rect 101 115 102 116
rect 100 115 101 116
rect 99 115 100 116
rect 98 115 99 116
rect 97 115 98 116
rect 96 115 97 116
rect 95 115 96 116
rect 94 115 95 116
rect 93 115 94 116
rect 92 115 93 116
rect 91 115 92 116
rect 90 115 91 116
rect 89 115 90 116
rect 88 115 89 116
rect 87 115 88 116
rect 86 115 87 116
rect 85 115 86 116
rect 84 115 85 116
rect 83 115 84 116
rect 82 115 83 116
rect 81 115 82 116
rect 80 115 81 116
rect 79 115 80 116
rect 78 115 79 116
rect 77 115 78 116
rect 76 115 77 116
rect 75 115 76 116
rect 74 115 75 116
rect 73 115 74 116
rect 72 115 73 116
rect 71 115 72 116
rect 70 115 71 116
rect 69 115 70 116
rect 60 115 61 116
rect 59 115 60 116
rect 58 115 59 116
rect 57 115 58 116
rect 56 115 57 116
rect 55 115 56 116
rect 54 115 55 116
rect 53 115 54 116
rect 52 115 53 116
rect 51 115 52 116
rect 50 115 51 116
rect 49 115 50 116
rect 48 115 49 116
rect 47 115 48 116
rect 46 115 47 116
rect 45 115 46 116
rect 44 115 45 116
rect 43 115 44 116
rect 42 115 43 116
rect 41 115 42 116
rect 40 115 41 116
rect 39 115 40 116
rect 38 115 39 116
rect 37 115 38 116
rect 36 115 37 116
rect 35 115 36 116
rect 34 115 35 116
rect 33 115 34 116
rect 32 115 33 116
rect 31 115 32 116
rect 30 115 31 116
rect 29 115 30 116
rect 478 116 479 117
rect 465 116 466 117
rect 464 116 465 117
rect 463 116 464 117
rect 462 116 463 117
rect 461 116 462 117
rect 460 116 461 117
rect 459 116 460 117
rect 437 116 438 117
rect 436 116 437 117
rect 435 116 436 117
rect 434 116 435 117
rect 433 116 434 117
rect 432 116 433 117
rect 431 116 432 117
rect 430 116 431 117
rect 429 116 430 117
rect 428 116 429 117
rect 396 116 397 117
rect 395 116 396 117
rect 394 116 395 117
rect 393 116 394 117
rect 242 116 243 117
rect 241 116 242 117
rect 240 116 241 117
rect 239 116 240 117
rect 238 116 239 117
rect 237 116 238 117
rect 236 116 237 117
rect 235 116 236 117
rect 234 116 235 117
rect 233 116 234 117
rect 232 116 233 117
rect 231 116 232 117
rect 230 116 231 117
rect 229 116 230 117
rect 228 116 229 117
rect 227 116 228 117
rect 226 116 227 117
rect 225 116 226 117
rect 224 116 225 117
rect 223 116 224 117
rect 222 116 223 117
rect 221 116 222 117
rect 220 116 221 117
rect 219 116 220 117
rect 218 116 219 117
rect 217 116 218 117
rect 216 116 217 117
rect 215 116 216 117
rect 214 116 215 117
rect 213 116 214 117
rect 212 116 213 117
rect 211 116 212 117
rect 210 116 211 117
rect 209 116 210 117
rect 208 116 209 117
rect 207 116 208 117
rect 206 116 207 117
rect 205 116 206 117
rect 204 116 205 117
rect 203 116 204 117
rect 202 116 203 117
rect 201 116 202 117
rect 200 116 201 117
rect 199 116 200 117
rect 198 116 199 117
rect 197 116 198 117
rect 196 116 197 117
rect 195 116 196 117
rect 194 116 195 117
rect 193 116 194 117
rect 192 116 193 117
rect 191 116 192 117
rect 190 116 191 117
rect 189 116 190 117
rect 188 116 189 117
rect 187 116 188 117
rect 186 116 187 117
rect 185 116 186 117
rect 184 116 185 117
rect 183 116 184 117
rect 182 116 183 117
rect 181 116 182 117
rect 180 116 181 117
rect 179 116 180 117
rect 178 116 179 117
rect 177 116 178 117
rect 176 116 177 117
rect 175 116 176 117
rect 174 116 175 117
rect 173 116 174 117
rect 172 116 173 117
rect 171 116 172 117
rect 170 116 171 117
rect 169 116 170 117
rect 168 116 169 117
rect 150 116 151 117
rect 149 116 150 117
rect 148 116 149 117
rect 147 116 148 117
rect 146 116 147 117
rect 145 116 146 117
rect 144 116 145 117
rect 143 116 144 117
rect 142 116 143 117
rect 141 116 142 117
rect 140 116 141 117
rect 139 116 140 117
rect 138 116 139 117
rect 137 116 138 117
rect 136 116 137 117
rect 135 116 136 117
rect 134 116 135 117
rect 133 116 134 117
rect 132 116 133 117
rect 131 116 132 117
rect 130 116 131 117
rect 129 116 130 117
rect 128 116 129 117
rect 127 116 128 117
rect 126 116 127 117
rect 125 116 126 117
rect 124 116 125 117
rect 123 116 124 117
rect 122 116 123 117
rect 121 116 122 117
rect 120 116 121 117
rect 119 116 120 117
rect 118 116 119 117
rect 117 116 118 117
rect 116 116 117 117
rect 115 116 116 117
rect 114 116 115 117
rect 113 116 114 117
rect 112 116 113 117
rect 111 116 112 117
rect 110 116 111 117
rect 109 116 110 117
rect 108 116 109 117
rect 107 116 108 117
rect 106 116 107 117
rect 105 116 106 117
rect 104 116 105 117
rect 103 116 104 117
rect 102 116 103 117
rect 101 116 102 117
rect 100 116 101 117
rect 99 116 100 117
rect 98 116 99 117
rect 97 116 98 117
rect 96 116 97 117
rect 95 116 96 117
rect 94 116 95 117
rect 93 116 94 117
rect 92 116 93 117
rect 91 116 92 117
rect 90 116 91 117
rect 89 116 90 117
rect 88 116 89 117
rect 87 116 88 117
rect 86 116 87 117
rect 85 116 86 117
rect 84 116 85 117
rect 83 116 84 117
rect 82 116 83 117
rect 81 116 82 117
rect 80 116 81 117
rect 79 116 80 117
rect 78 116 79 117
rect 77 116 78 117
rect 76 116 77 117
rect 75 116 76 117
rect 74 116 75 117
rect 73 116 74 117
rect 72 116 73 117
rect 71 116 72 117
rect 70 116 71 117
rect 69 116 70 117
rect 68 116 69 117
rect 59 116 60 117
rect 58 116 59 117
rect 57 116 58 117
rect 56 116 57 117
rect 55 116 56 117
rect 54 116 55 117
rect 53 116 54 117
rect 52 116 53 117
rect 51 116 52 117
rect 50 116 51 117
rect 49 116 50 117
rect 48 116 49 117
rect 47 116 48 117
rect 46 116 47 117
rect 45 116 46 117
rect 44 116 45 117
rect 43 116 44 117
rect 42 116 43 117
rect 41 116 42 117
rect 40 116 41 117
rect 39 116 40 117
rect 38 116 39 117
rect 37 116 38 117
rect 36 116 37 117
rect 35 116 36 117
rect 34 116 35 117
rect 33 116 34 117
rect 32 116 33 117
rect 31 116 32 117
rect 30 116 31 117
rect 29 116 30 117
rect 478 117 479 118
rect 466 117 467 118
rect 465 117 466 118
rect 464 117 465 118
rect 463 117 464 118
rect 462 117 463 118
rect 461 117 462 118
rect 460 117 461 118
rect 438 117 439 118
rect 437 117 438 118
rect 436 117 437 118
rect 435 117 436 118
rect 434 117 435 118
rect 433 117 434 118
rect 432 117 433 118
rect 431 117 432 118
rect 430 117 431 118
rect 395 117 396 118
rect 394 117 395 118
rect 393 117 394 118
rect 240 117 241 118
rect 239 117 240 118
rect 238 117 239 118
rect 237 117 238 118
rect 236 117 237 118
rect 235 117 236 118
rect 234 117 235 118
rect 233 117 234 118
rect 232 117 233 118
rect 231 117 232 118
rect 230 117 231 118
rect 229 117 230 118
rect 228 117 229 118
rect 227 117 228 118
rect 226 117 227 118
rect 225 117 226 118
rect 224 117 225 118
rect 223 117 224 118
rect 222 117 223 118
rect 221 117 222 118
rect 220 117 221 118
rect 219 117 220 118
rect 218 117 219 118
rect 217 117 218 118
rect 216 117 217 118
rect 215 117 216 118
rect 214 117 215 118
rect 213 117 214 118
rect 212 117 213 118
rect 211 117 212 118
rect 210 117 211 118
rect 209 117 210 118
rect 208 117 209 118
rect 207 117 208 118
rect 206 117 207 118
rect 205 117 206 118
rect 204 117 205 118
rect 203 117 204 118
rect 202 117 203 118
rect 201 117 202 118
rect 200 117 201 118
rect 199 117 200 118
rect 198 117 199 118
rect 197 117 198 118
rect 196 117 197 118
rect 195 117 196 118
rect 194 117 195 118
rect 193 117 194 118
rect 192 117 193 118
rect 191 117 192 118
rect 190 117 191 118
rect 189 117 190 118
rect 188 117 189 118
rect 187 117 188 118
rect 186 117 187 118
rect 185 117 186 118
rect 184 117 185 118
rect 183 117 184 118
rect 182 117 183 118
rect 181 117 182 118
rect 180 117 181 118
rect 179 117 180 118
rect 178 117 179 118
rect 177 117 178 118
rect 176 117 177 118
rect 175 117 176 118
rect 174 117 175 118
rect 173 117 174 118
rect 172 117 173 118
rect 171 117 172 118
rect 170 117 171 118
rect 169 117 170 118
rect 168 117 169 118
rect 167 117 168 118
rect 150 117 151 118
rect 149 117 150 118
rect 148 117 149 118
rect 147 117 148 118
rect 146 117 147 118
rect 145 117 146 118
rect 144 117 145 118
rect 143 117 144 118
rect 142 117 143 118
rect 141 117 142 118
rect 140 117 141 118
rect 139 117 140 118
rect 138 117 139 118
rect 137 117 138 118
rect 136 117 137 118
rect 135 117 136 118
rect 134 117 135 118
rect 133 117 134 118
rect 132 117 133 118
rect 131 117 132 118
rect 130 117 131 118
rect 129 117 130 118
rect 128 117 129 118
rect 127 117 128 118
rect 126 117 127 118
rect 125 117 126 118
rect 124 117 125 118
rect 123 117 124 118
rect 122 117 123 118
rect 121 117 122 118
rect 120 117 121 118
rect 119 117 120 118
rect 118 117 119 118
rect 117 117 118 118
rect 116 117 117 118
rect 115 117 116 118
rect 114 117 115 118
rect 113 117 114 118
rect 112 117 113 118
rect 111 117 112 118
rect 110 117 111 118
rect 109 117 110 118
rect 108 117 109 118
rect 107 117 108 118
rect 106 117 107 118
rect 105 117 106 118
rect 104 117 105 118
rect 103 117 104 118
rect 102 117 103 118
rect 101 117 102 118
rect 100 117 101 118
rect 99 117 100 118
rect 98 117 99 118
rect 97 117 98 118
rect 96 117 97 118
rect 95 117 96 118
rect 94 117 95 118
rect 93 117 94 118
rect 92 117 93 118
rect 91 117 92 118
rect 90 117 91 118
rect 89 117 90 118
rect 88 117 89 118
rect 87 117 88 118
rect 86 117 87 118
rect 85 117 86 118
rect 84 117 85 118
rect 83 117 84 118
rect 82 117 83 118
rect 81 117 82 118
rect 80 117 81 118
rect 79 117 80 118
rect 78 117 79 118
rect 77 117 78 118
rect 76 117 77 118
rect 75 117 76 118
rect 74 117 75 118
rect 73 117 74 118
rect 72 117 73 118
rect 71 117 72 118
rect 70 117 71 118
rect 69 117 70 118
rect 68 117 69 118
rect 67 117 68 118
rect 59 117 60 118
rect 58 117 59 118
rect 57 117 58 118
rect 56 117 57 118
rect 55 117 56 118
rect 54 117 55 118
rect 53 117 54 118
rect 52 117 53 118
rect 51 117 52 118
rect 50 117 51 118
rect 49 117 50 118
rect 48 117 49 118
rect 47 117 48 118
rect 46 117 47 118
rect 45 117 46 118
rect 44 117 45 118
rect 43 117 44 118
rect 42 117 43 118
rect 41 117 42 118
rect 40 117 41 118
rect 39 117 40 118
rect 38 117 39 118
rect 37 117 38 118
rect 36 117 37 118
rect 35 117 36 118
rect 34 117 35 118
rect 33 117 34 118
rect 32 117 33 118
rect 31 117 32 118
rect 30 117 31 118
rect 29 117 30 118
rect 28 117 29 118
rect 467 118 468 119
rect 466 118 467 119
rect 465 118 466 119
rect 464 118 465 119
rect 463 118 464 119
rect 462 118 463 119
rect 461 118 462 119
rect 438 118 439 119
rect 437 118 438 119
rect 436 118 437 119
rect 435 118 436 119
rect 434 118 435 119
rect 433 118 434 119
rect 432 118 433 119
rect 431 118 432 119
rect 395 118 396 119
rect 394 118 395 119
rect 393 118 394 119
rect 238 118 239 119
rect 237 118 238 119
rect 236 118 237 119
rect 235 118 236 119
rect 234 118 235 119
rect 233 118 234 119
rect 232 118 233 119
rect 231 118 232 119
rect 230 118 231 119
rect 229 118 230 119
rect 228 118 229 119
rect 227 118 228 119
rect 226 118 227 119
rect 225 118 226 119
rect 224 118 225 119
rect 223 118 224 119
rect 222 118 223 119
rect 221 118 222 119
rect 220 118 221 119
rect 219 118 220 119
rect 218 118 219 119
rect 217 118 218 119
rect 216 118 217 119
rect 215 118 216 119
rect 214 118 215 119
rect 213 118 214 119
rect 212 118 213 119
rect 211 118 212 119
rect 210 118 211 119
rect 209 118 210 119
rect 208 118 209 119
rect 207 118 208 119
rect 206 118 207 119
rect 205 118 206 119
rect 204 118 205 119
rect 203 118 204 119
rect 202 118 203 119
rect 201 118 202 119
rect 200 118 201 119
rect 199 118 200 119
rect 198 118 199 119
rect 197 118 198 119
rect 196 118 197 119
rect 195 118 196 119
rect 194 118 195 119
rect 193 118 194 119
rect 192 118 193 119
rect 191 118 192 119
rect 190 118 191 119
rect 189 118 190 119
rect 188 118 189 119
rect 187 118 188 119
rect 186 118 187 119
rect 185 118 186 119
rect 184 118 185 119
rect 183 118 184 119
rect 182 118 183 119
rect 181 118 182 119
rect 180 118 181 119
rect 179 118 180 119
rect 178 118 179 119
rect 177 118 178 119
rect 176 118 177 119
rect 175 118 176 119
rect 174 118 175 119
rect 173 118 174 119
rect 172 118 173 119
rect 171 118 172 119
rect 170 118 171 119
rect 169 118 170 119
rect 168 118 169 119
rect 167 118 168 119
rect 149 118 150 119
rect 148 118 149 119
rect 147 118 148 119
rect 146 118 147 119
rect 145 118 146 119
rect 144 118 145 119
rect 143 118 144 119
rect 142 118 143 119
rect 141 118 142 119
rect 140 118 141 119
rect 139 118 140 119
rect 138 118 139 119
rect 137 118 138 119
rect 136 118 137 119
rect 135 118 136 119
rect 134 118 135 119
rect 133 118 134 119
rect 132 118 133 119
rect 131 118 132 119
rect 130 118 131 119
rect 129 118 130 119
rect 128 118 129 119
rect 127 118 128 119
rect 126 118 127 119
rect 125 118 126 119
rect 124 118 125 119
rect 123 118 124 119
rect 122 118 123 119
rect 121 118 122 119
rect 120 118 121 119
rect 119 118 120 119
rect 118 118 119 119
rect 117 118 118 119
rect 116 118 117 119
rect 115 118 116 119
rect 114 118 115 119
rect 113 118 114 119
rect 112 118 113 119
rect 111 118 112 119
rect 110 118 111 119
rect 109 118 110 119
rect 108 118 109 119
rect 107 118 108 119
rect 106 118 107 119
rect 105 118 106 119
rect 104 118 105 119
rect 103 118 104 119
rect 102 118 103 119
rect 101 118 102 119
rect 100 118 101 119
rect 99 118 100 119
rect 98 118 99 119
rect 97 118 98 119
rect 96 118 97 119
rect 95 118 96 119
rect 94 118 95 119
rect 93 118 94 119
rect 92 118 93 119
rect 91 118 92 119
rect 90 118 91 119
rect 89 118 90 119
rect 88 118 89 119
rect 87 118 88 119
rect 86 118 87 119
rect 85 118 86 119
rect 84 118 85 119
rect 83 118 84 119
rect 82 118 83 119
rect 81 118 82 119
rect 80 118 81 119
rect 79 118 80 119
rect 78 118 79 119
rect 77 118 78 119
rect 76 118 77 119
rect 75 118 76 119
rect 74 118 75 119
rect 73 118 74 119
rect 72 118 73 119
rect 71 118 72 119
rect 70 118 71 119
rect 69 118 70 119
rect 68 118 69 119
rect 67 118 68 119
rect 59 118 60 119
rect 58 118 59 119
rect 57 118 58 119
rect 56 118 57 119
rect 55 118 56 119
rect 54 118 55 119
rect 53 118 54 119
rect 52 118 53 119
rect 51 118 52 119
rect 50 118 51 119
rect 49 118 50 119
rect 48 118 49 119
rect 47 118 48 119
rect 46 118 47 119
rect 45 118 46 119
rect 44 118 45 119
rect 43 118 44 119
rect 42 118 43 119
rect 41 118 42 119
rect 40 118 41 119
rect 39 118 40 119
rect 38 118 39 119
rect 37 118 38 119
rect 36 118 37 119
rect 35 118 36 119
rect 34 118 35 119
rect 33 118 34 119
rect 32 118 33 119
rect 31 118 32 119
rect 30 118 31 119
rect 29 118 30 119
rect 28 118 29 119
rect 469 119 470 120
rect 468 119 469 120
rect 467 119 468 120
rect 466 119 467 120
rect 465 119 466 120
rect 464 119 465 120
rect 463 119 464 120
rect 462 119 463 120
rect 438 119 439 120
rect 437 119 438 120
rect 436 119 437 120
rect 435 119 436 120
rect 434 119 435 120
rect 433 119 434 120
rect 432 119 433 120
rect 395 119 396 120
rect 394 119 395 120
rect 393 119 394 120
rect 236 119 237 120
rect 235 119 236 120
rect 234 119 235 120
rect 233 119 234 120
rect 232 119 233 120
rect 231 119 232 120
rect 230 119 231 120
rect 229 119 230 120
rect 228 119 229 120
rect 227 119 228 120
rect 226 119 227 120
rect 225 119 226 120
rect 224 119 225 120
rect 223 119 224 120
rect 222 119 223 120
rect 221 119 222 120
rect 220 119 221 120
rect 219 119 220 120
rect 218 119 219 120
rect 217 119 218 120
rect 216 119 217 120
rect 215 119 216 120
rect 214 119 215 120
rect 213 119 214 120
rect 212 119 213 120
rect 211 119 212 120
rect 210 119 211 120
rect 209 119 210 120
rect 208 119 209 120
rect 207 119 208 120
rect 206 119 207 120
rect 205 119 206 120
rect 204 119 205 120
rect 203 119 204 120
rect 202 119 203 120
rect 201 119 202 120
rect 200 119 201 120
rect 199 119 200 120
rect 198 119 199 120
rect 197 119 198 120
rect 196 119 197 120
rect 195 119 196 120
rect 194 119 195 120
rect 193 119 194 120
rect 192 119 193 120
rect 191 119 192 120
rect 190 119 191 120
rect 189 119 190 120
rect 188 119 189 120
rect 187 119 188 120
rect 186 119 187 120
rect 185 119 186 120
rect 184 119 185 120
rect 183 119 184 120
rect 182 119 183 120
rect 181 119 182 120
rect 180 119 181 120
rect 179 119 180 120
rect 178 119 179 120
rect 177 119 178 120
rect 176 119 177 120
rect 175 119 176 120
rect 174 119 175 120
rect 173 119 174 120
rect 172 119 173 120
rect 171 119 172 120
rect 170 119 171 120
rect 169 119 170 120
rect 168 119 169 120
rect 167 119 168 120
rect 166 119 167 120
rect 149 119 150 120
rect 148 119 149 120
rect 147 119 148 120
rect 146 119 147 120
rect 145 119 146 120
rect 144 119 145 120
rect 143 119 144 120
rect 142 119 143 120
rect 141 119 142 120
rect 140 119 141 120
rect 139 119 140 120
rect 138 119 139 120
rect 137 119 138 120
rect 136 119 137 120
rect 135 119 136 120
rect 134 119 135 120
rect 133 119 134 120
rect 132 119 133 120
rect 131 119 132 120
rect 130 119 131 120
rect 129 119 130 120
rect 128 119 129 120
rect 127 119 128 120
rect 126 119 127 120
rect 125 119 126 120
rect 124 119 125 120
rect 123 119 124 120
rect 122 119 123 120
rect 121 119 122 120
rect 120 119 121 120
rect 119 119 120 120
rect 118 119 119 120
rect 117 119 118 120
rect 116 119 117 120
rect 115 119 116 120
rect 114 119 115 120
rect 113 119 114 120
rect 112 119 113 120
rect 111 119 112 120
rect 110 119 111 120
rect 109 119 110 120
rect 108 119 109 120
rect 107 119 108 120
rect 106 119 107 120
rect 105 119 106 120
rect 104 119 105 120
rect 103 119 104 120
rect 102 119 103 120
rect 101 119 102 120
rect 100 119 101 120
rect 99 119 100 120
rect 98 119 99 120
rect 97 119 98 120
rect 96 119 97 120
rect 95 119 96 120
rect 94 119 95 120
rect 93 119 94 120
rect 92 119 93 120
rect 91 119 92 120
rect 90 119 91 120
rect 89 119 90 120
rect 88 119 89 120
rect 87 119 88 120
rect 86 119 87 120
rect 85 119 86 120
rect 84 119 85 120
rect 83 119 84 120
rect 82 119 83 120
rect 81 119 82 120
rect 80 119 81 120
rect 79 119 80 120
rect 78 119 79 120
rect 77 119 78 120
rect 76 119 77 120
rect 75 119 76 120
rect 74 119 75 120
rect 73 119 74 120
rect 72 119 73 120
rect 71 119 72 120
rect 70 119 71 120
rect 69 119 70 120
rect 68 119 69 120
rect 67 119 68 120
rect 66 119 67 120
rect 58 119 59 120
rect 57 119 58 120
rect 56 119 57 120
rect 55 119 56 120
rect 54 119 55 120
rect 53 119 54 120
rect 52 119 53 120
rect 51 119 52 120
rect 50 119 51 120
rect 49 119 50 120
rect 48 119 49 120
rect 47 119 48 120
rect 46 119 47 120
rect 45 119 46 120
rect 44 119 45 120
rect 43 119 44 120
rect 42 119 43 120
rect 41 119 42 120
rect 40 119 41 120
rect 39 119 40 120
rect 38 119 39 120
rect 37 119 38 120
rect 36 119 37 120
rect 35 119 36 120
rect 34 119 35 120
rect 33 119 34 120
rect 32 119 33 120
rect 31 119 32 120
rect 30 119 31 120
rect 29 119 30 120
rect 28 119 29 120
rect 470 120 471 121
rect 469 120 470 121
rect 468 120 469 121
rect 467 120 468 121
rect 466 120 467 121
rect 465 120 466 121
rect 464 120 465 121
rect 438 120 439 121
rect 437 120 438 121
rect 436 120 437 121
rect 435 120 436 121
rect 434 120 435 121
rect 433 120 434 121
rect 394 120 395 121
rect 393 120 394 121
rect 235 120 236 121
rect 234 120 235 121
rect 233 120 234 121
rect 232 120 233 121
rect 231 120 232 121
rect 230 120 231 121
rect 229 120 230 121
rect 228 120 229 121
rect 227 120 228 121
rect 226 120 227 121
rect 225 120 226 121
rect 224 120 225 121
rect 223 120 224 121
rect 222 120 223 121
rect 221 120 222 121
rect 220 120 221 121
rect 219 120 220 121
rect 218 120 219 121
rect 217 120 218 121
rect 216 120 217 121
rect 215 120 216 121
rect 214 120 215 121
rect 213 120 214 121
rect 212 120 213 121
rect 211 120 212 121
rect 210 120 211 121
rect 209 120 210 121
rect 208 120 209 121
rect 207 120 208 121
rect 206 120 207 121
rect 205 120 206 121
rect 204 120 205 121
rect 203 120 204 121
rect 202 120 203 121
rect 201 120 202 121
rect 200 120 201 121
rect 199 120 200 121
rect 198 120 199 121
rect 197 120 198 121
rect 196 120 197 121
rect 195 120 196 121
rect 194 120 195 121
rect 193 120 194 121
rect 192 120 193 121
rect 191 120 192 121
rect 190 120 191 121
rect 189 120 190 121
rect 188 120 189 121
rect 187 120 188 121
rect 186 120 187 121
rect 185 120 186 121
rect 184 120 185 121
rect 183 120 184 121
rect 182 120 183 121
rect 181 120 182 121
rect 180 120 181 121
rect 179 120 180 121
rect 178 120 179 121
rect 177 120 178 121
rect 176 120 177 121
rect 175 120 176 121
rect 174 120 175 121
rect 173 120 174 121
rect 172 120 173 121
rect 171 120 172 121
rect 170 120 171 121
rect 169 120 170 121
rect 168 120 169 121
rect 167 120 168 121
rect 166 120 167 121
rect 149 120 150 121
rect 148 120 149 121
rect 147 120 148 121
rect 146 120 147 121
rect 145 120 146 121
rect 144 120 145 121
rect 143 120 144 121
rect 142 120 143 121
rect 141 120 142 121
rect 140 120 141 121
rect 139 120 140 121
rect 138 120 139 121
rect 137 120 138 121
rect 136 120 137 121
rect 135 120 136 121
rect 134 120 135 121
rect 133 120 134 121
rect 132 120 133 121
rect 131 120 132 121
rect 130 120 131 121
rect 129 120 130 121
rect 128 120 129 121
rect 127 120 128 121
rect 126 120 127 121
rect 125 120 126 121
rect 124 120 125 121
rect 123 120 124 121
rect 122 120 123 121
rect 121 120 122 121
rect 120 120 121 121
rect 119 120 120 121
rect 118 120 119 121
rect 117 120 118 121
rect 116 120 117 121
rect 115 120 116 121
rect 114 120 115 121
rect 113 120 114 121
rect 112 120 113 121
rect 111 120 112 121
rect 110 120 111 121
rect 109 120 110 121
rect 108 120 109 121
rect 107 120 108 121
rect 106 120 107 121
rect 105 120 106 121
rect 104 120 105 121
rect 103 120 104 121
rect 102 120 103 121
rect 101 120 102 121
rect 100 120 101 121
rect 99 120 100 121
rect 98 120 99 121
rect 97 120 98 121
rect 96 120 97 121
rect 95 120 96 121
rect 94 120 95 121
rect 93 120 94 121
rect 92 120 93 121
rect 91 120 92 121
rect 90 120 91 121
rect 89 120 90 121
rect 88 120 89 121
rect 87 120 88 121
rect 86 120 87 121
rect 85 120 86 121
rect 84 120 85 121
rect 83 120 84 121
rect 82 120 83 121
rect 81 120 82 121
rect 80 120 81 121
rect 79 120 80 121
rect 78 120 79 121
rect 77 120 78 121
rect 76 120 77 121
rect 75 120 76 121
rect 74 120 75 121
rect 73 120 74 121
rect 72 120 73 121
rect 71 120 72 121
rect 70 120 71 121
rect 69 120 70 121
rect 68 120 69 121
rect 67 120 68 121
rect 66 120 67 121
rect 65 120 66 121
rect 58 120 59 121
rect 57 120 58 121
rect 56 120 57 121
rect 55 120 56 121
rect 54 120 55 121
rect 53 120 54 121
rect 52 120 53 121
rect 51 120 52 121
rect 50 120 51 121
rect 49 120 50 121
rect 48 120 49 121
rect 47 120 48 121
rect 46 120 47 121
rect 45 120 46 121
rect 44 120 45 121
rect 43 120 44 121
rect 42 120 43 121
rect 41 120 42 121
rect 40 120 41 121
rect 39 120 40 121
rect 38 120 39 121
rect 37 120 38 121
rect 36 120 37 121
rect 35 120 36 121
rect 34 120 35 121
rect 33 120 34 121
rect 32 120 33 121
rect 31 120 32 121
rect 30 120 31 121
rect 29 120 30 121
rect 28 120 29 121
rect 27 120 28 121
rect 471 121 472 122
rect 470 121 471 122
rect 469 121 470 122
rect 468 121 469 122
rect 467 121 468 122
rect 466 121 467 122
rect 465 121 466 122
rect 438 121 439 122
rect 437 121 438 122
rect 436 121 437 122
rect 435 121 436 122
rect 434 121 435 122
rect 433 121 434 122
rect 288 121 289 122
rect 287 121 288 122
rect 286 121 287 122
rect 285 121 286 122
rect 284 121 285 122
rect 283 121 284 122
rect 282 121 283 122
rect 281 121 282 122
rect 280 121 281 122
rect 279 121 280 122
rect 233 121 234 122
rect 232 121 233 122
rect 231 121 232 122
rect 230 121 231 122
rect 229 121 230 122
rect 228 121 229 122
rect 227 121 228 122
rect 226 121 227 122
rect 225 121 226 122
rect 224 121 225 122
rect 223 121 224 122
rect 222 121 223 122
rect 221 121 222 122
rect 220 121 221 122
rect 219 121 220 122
rect 218 121 219 122
rect 217 121 218 122
rect 216 121 217 122
rect 215 121 216 122
rect 214 121 215 122
rect 213 121 214 122
rect 212 121 213 122
rect 211 121 212 122
rect 210 121 211 122
rect 209 121 210 122
rect 208 121 209 122
rect 207 121 208 122
rect 206 121 207 122
rect 205 121 206 122
rect 204 121 205 122
rect 203 121 204 122
rect 202 121 203 122
rect 201 121 202 122
rect 200 121 201 122
rect 199 121 200 122
rect 198 121 199 122
rect 197 121 198 122
rect 196 121 197 122
rect 195 121 196 122
rect 194 121 195 122
rect 193 121 194 122
rect 192 121 193 122
rect 191 121 192 122
rect 190 121 191 122
rect 189 121 190 122
rect 188 121 189 122
rect 187 121 188 122
rect 186 121 187 122
rect 185 121 186 122
rect 184 121 185 122
rect 183 121 184 122
rect 182 121 183 122
rect 181 121 182 122
rect 180 121 181 122
rect 179 121 180 122
rect 178 121 179 122
rect 177 121 178 122
rect 176 121 177 122
rect 175 121 176 122
rect 174 121 175 122
rect 173 121 174 122
rect 172 121 173 122
rect 171 121 172 122
rect 170 121 171 122
rect 169 121 170 122
rect 168 121 169 122
rect 167 121 168 122
rect 166 121 167 122
rect 165 121 166 122
rect 148 121 149 122
rect 147 121 148 122
rect 146 121 147 122
rect 145 121 146 122
rect 144 121 145 122
rect 143 121 144 122
rect 142 121 143 122
rect 141 121 142 122
rect 140 121 141 122
rect 139 121 140 122
rect 138 121 139 122
rect 137 121 138 122
rect 136 121 137 122
rect 135 121 136 122
rect 134 121 135 122
rect 133 121 134 122
rect 132 121 133 122
rect 131 121 132 122
rect 130 121 131 122
rect 129 121 130 122
rect 128 121 129 122
rect 127 121 128 122
rect 126 121 127 122
rect 125 121 126 122
rect 124 121 125 122
rect 123 121 124 122
rect 122 121 123 122
rect 121 121 122 122
rect 120 121 121 122
rect 119 121 120 122
rect 118 121 119 122
rect 117 121 118 122
rect 116 121 117 122
rect 115 121 116 122
rect 114 121 115 122
rect 113 121 114 122
rect 112 121 113 122
rect 111 121 112 122
rect 110 121 111 122
rect 109 121 110 122
rect 108 121 109 122
rect 107 121 108 122
rect 106 121 107 122
rect 105 121 106 122
rect 104 121 105 122
rect 103 121 104 122
rect 102 121 103 122
rect 101 121 102 122
rect 100 121 101 122
rect 99 121 100 122
rect 98 121 99 122
rect 97 121 98 122
rect 96 121 97 122
rect 95 121 96 122
rect 94 121 95 122
rect 93 121 94 122
rect 92 121 93 122
rect 91 121 92 122
rect 90 121 91 122
rect 89 121 90 122
rect 88 121 89 122
rect 87 121 88 122
rect 86 121 87 122
rect 85 121 86 122
rect 84 121 85 122
rect 83 121 84 122
rect 82 121 83 122
rect 81 121 82 122
rect 80 121 81 122
rect 79 121 80 122
rect 78 121 79 122
rect 77 121 78 122
rect 76 121 77 122
rect 75 121 76 122
rect 74 121 75 122
rect 73 121 74 122
rect 72 121 73 122
rect 71 121 72 122
rect 70 121 71 122
rect 69 121 70 122
rect 68 121 69 122
rect 67 121 68 122
rect 66 121 67 122
rect 65 121 66 122
rect 58 121 59 122
rect 57 121 58 122
rect 56 121 57 122
rect 55 121 56 122
rect 54 121 55 122
rect 53 121 54 122
rect 52 121 53 122
rect 51 121 52 122
rect 50 121 51 122
rect 49 121 50 122
rect 48 121 49 122
rect 47 121 48 122
rect 46 121 47 122
rect 45 121 46 122
rect 44 121 45 122
rect 43 121 44 122
rect 42 121 43 122
rect 41 121 42 122
rect 40 121 41 122
rect 39 121 40 122
rect 38 121 39 122
rect 37 121 38 122
rect 36 121 37 122
rect 35 121 36 122
rect 34 121 35 122
rect 33 121 34 122
rect 32 121 33 122
rect 31 121 32 122
rect 30 121 31 122
rect 29 121 30 122
rect 28 121 29 122
rect 27 121 28 122
rect 472 122 473 123
rect 471 122 472 123
rect 470 122 471 123
rect 469 122 470 123
rect 468 122 469 123
rect 467 122 468 123
rect 466 122 467 123
rect 438 122 439 123
rect 437 122 438 123
rect 436 122 437 123
rect 435 122 436 123
rect 434 122 435 123
rect 291 122 292 123
rect 290 122 291 123
rect 289 122 290 123
rect 288 122 289 123
rect 287 122 288 123
rect 286 122 287 123
rect 285 122 286 123
rect 284 122 285 123
rect 283 122 284 123
rect 282 122 283 123
rect 281 122 282 123
rect 280 122 281 123
rect 279 122 280 123
rect 278 122 279 123
rect 277 122 278 123
rect 276 122 277 123
rect 275 122 276 123
rect 274 122 275 123
rect 232 122 233 123
rect 231 122 232 123
rect 230 122 231 123
rect 229 122 230 123
rect 228 122 229 123
rect 227 122 228 123
rect 226 122 227 123
rect 225 122 226 123
rect 224 122 225 123
rect 223 122 224 123
rect 222 122 223 123
rect 221 122 222 123
rect 220 122 221 123
rect 219 122 220 123
rect 218 122 219 123
rect 217 122 218 123
rect 216 122 217 123
rect 215 122 216 123
rect 214 122 215 123
rect 213 122 214 123
rect 212 122 213 123
rect 211 122 212 123
rect 210 122 211 123
rect 209 122 210 123
rect 208 122 209 123
rect 207 122 208 123
rect 206 122 207 123
rect 205 122 206 123
rect 204 122 205 123
rect 203 122 204 123
rect 202 122 203 123
rect 201 122 202 123
rect 200 122 201 123
rect 199 122 200 123
rect 198 122 199 123
rect 197 122 198 123
rect 196 122 197 123
rect 195 122 196 123
rect 194 122 195 123
rect 193 122 194 123
rect 192 122 193 123
rect 191 122 192 123
rect 190 122 191 123
rect 189 122 190 123
rect 188 122 189 123
rect 187 122 188 123
rect 186 122 187 123
rect 185 122 186 123
rect 184 122 185 123
rect 183 122 184 123
rect 182 122 183 123
rect 181 122 182 123
rect 180 122 181 123
rect 179 122 180 123
rect 178 122 179 123
rect 177 122 178 123
rect 176 122 177 123
rect 175 122 176 123
rect 174 122 175 123
rect 173 122 174 123
rect 172 122 173 123
rect 171 122 172 123
rect 170 122 171 123
rect 169 122 170 123
rect 168 122 169 123
rect 167 122 168 123
rect 166 122 167 123
rect 165 122 166 123
rect 148 122 149 123
rect 147 122 148 123
rect 146 122 147 123
rect 145 122 146 123
rect 144 122 145 123
rect 143 122 144 123
rect 142 122 143 123
rect 141 122 142 123
rect 140 122 141 123
rect 139 122 140 123
rect 138 122 139 123
rect 137 122 138 123
rect 136 122 137 123
rect 135 122 136 123
rect 134 122 135 123
rect 133 122 134 123
rect 132 122 133 123
rect 131 122 132 123
rect 130 122 131 123
rect 129 122 130 123
rect 128 122 129 123
rect 127 122 128 123
rect 126 122 127 123
rect 125 122 126 123
rect 124 122 125 123
rect 123 122 124 123
rect 122 122 123 123
rect 121 122 122 123
rect 120 122 121 123
rect 119 122 120 123
rect 118 122 119 123
rect 117 122 118 123
rect 116 122 117 123
rect 115 122 116 123
rect 114 122 115 123
rect 113 122 114 123
rect 112 122 113 123
rect 111 122 112 123
rect 110 122 111 123
rect 109 122 110 123
rect 108 122 109 123
rect 107 122 108 123
rect 106 122 107 123
rect 105 122 106 123
rect 104 122 105 123
rect 103 122 104 123
rect 102 122 103 123
rect 101 122 102 123
rect 100 122 101 123
rect 99 122 100 123
rect 98 122 99 123
rect 97 122 98 123
rect 96 122 97 123
rect 95 122 96 123
rect 94 122 95 123
rect 93 122 94 123
rect 92 122 93 123
rect 91 122 92 123
rect 90 122 91 123
rect 89 122 90 123
rect 88 122 89 123
rect 87 122 88 123
rect 86 122 87 123
rect 85 122 86 123
rect 84 122 85 123
rect 83 122 84 123
rect 82 122 83 123
rect 81 122 82 123
rect 80 122 81 123
rect 79 122 80 123
rect 78 122 79 123
rect 77 122 78 123
rect 76 122 77 123
rect 75 122 76 123
rect 74 122 75 123
rect 73 122 74 123
rect 72 122 73 123
rect 71 122 72 123
rect 70 122 71 123
rect 69 122 70 123
rect 68 122 69 123
rect 67 122 68 123
rect 66 122 67 123
rect 65 122 66 123
rect 64 122 65 123
rect 58 122 59 123
rect 57 122 58 123
rect 56 122 57 123
rect 55 122 56 123
rect 54 122 55 123
rect 53 122 54 123
rect 52 122 53 123
rect 51 122 52 123
rect 50 122 51 123
rect 49 122 50 123
rect 48 122 49 123
rect 47 122 48 123
rect 46 122 47 123
rect 45 122 46 123
rect 44 122 45 123
rect 43 122 44 123
rect 42 122 43 123
rect 41 122 42 123
rect 40 122 41 123
rect 39 122 40 123
rect 38 122 39 123
rect 37 122 38 123
rect 36 122 37 123
rect 35 122 36 123
rect 34 122 35 123
rect 33 122 34 123
rect 32 122 33 123
rect 31 122 32 123
rect 30 122 31 123
rect 29 122 30 123
rect 28 122 29 123
rect 27 122 28 123
rect 473 123 474 124
rect 472 123 473 124
rect 471 123 472 124
rect 470 123 471 124
rect 469 123 470 124
rect 468 123 469 124
rect 467 123 468 124
rect 438 123 439 124
rect 437 123 438 124
rect 436 123 437 124
rect 435 123 436 124
rect 434 123 435 124
rect 293 123 294 124
rect 292 123 293 124
rect 291 123 292 124
rect 290 123 291 124
rect 289 123 290 124
rect 288 123 289 124
rect 287 123 288 124
rect 286 123 287 124
rect 285 123 286 124
rect 284 123 285 124
rect 283 123 284 124
rect 282 123 283 124
rect 281 123 282 124
rect 280 123 281 124
rect 279 123 280 124
rect 278 123 279 124
rect 277 123 278 124
rect 276 123 277 124
rect 275 123 276 124
rect 274 123 275 124
rect 273 123 274 124
rect 272 123 273 124
rect 271 123 272 124
rect 270 123 271 124
rect 231 123 232 124
rect 230 123 231 124
rect 229 123 230 124
rect 228 123 229 124
rect 227 123 228 124
rect 226 123 227 124
rect 225 123 226 124
rect 224 123 225 124
rect 223 123 224 124
rect 222 123 223 124
rect 221 123 222 124
rect 220 123 221 124
rect 219 123 220 124
rect 218 123 219 124
rect 217 123 218 124
rect 216 123 217 124
rect 215 123 216 124
rect 214 123 215 124
rect 213 123 214 124
rect 212 123 213 124
rect 211 123 212 124
rect 210 123 211 124
rect 209 123 210 124
rect 208 123 209 124
rect 207 123 208 124
rect 206 123 207 124
rect 205 123 206 124
rect 204 123 205 124
rect 203 123 204 124
rect 202 123 203 124
rect 201 123 202 124
rect 200 123 201 124
rect 199 123 200 124
rect 198 123 199 124
rect 197 123 198 124
rect 196 123 197 124
rect 195 123 196 124
rect 194 123 195 124
rect 193 123 194 124
rect 192 123 193 124
rect 191 123 192 124
rect 190 123 191 124
rect 189 123 190 124
rect 188 123 189 124
rect 187 123 188 124
rect 186 123 187 124
rect 185 123 186 124
rect 184 123 185 124
rect 183 123 184 124
rect 182 123 183 124
rect 181 123 182 124
rect 180 123 181 124
rect 179 123 180 124
rect 178 123 179 124
rect 177 123 178 124
rect 176 123 177 124
rect 175 123 176 124
rect 174 123 175 124
rect 173 123 174 124
rect 172 123 173 124
rect 171 123 172 124
rect 170 123 171 124
rect 169 123 170 124
rect 168 123 169 124
rect 167 123 168 124
rect 166 123 167 124
rect 165 123 166 124
rect 147 123 148 124
rect 146 123 147 124
rect 145 123 146 124
rect 144 123 145 124
rect 143 123 144 124
rect 142 123 143 124
rect 141 123 142 124
rect 140 123 141 124
rect 139 123 140 124
rect 138 123 139 124
rect 137 123 138 124
rect 136 123 137 124
rect 135 123 136 124
rect 134 123 135 124
rect 133 123 134 124
rect 132 123 133 124
rect 131 123 132 124
rect 130 123 131 124
rect 129 123 130 124
rect 128 123 129 124
rect 127 123 128 124
rect 126 123 127 124
rect 125 123 126 124
rect 124 123 125 124
rect 123 123 124 124
rect 122 123 123 124
rect 121 123 122 124
rect 120 123 121 124
rect 119 123 120 124
rect 118 123 119 124
rect 117 123 118 124
rect 116 123 117 124
rect 115 123 116 124
rect 114 123 115 124
rect 113 123 114 124
rect 112 123 113 124
rect 111 123 112 124
rect 110 123 111 124
rect 109 123 110 124
rect 108 123 109 124
rect 107 123 108 124
rect 106 123 107 124
rect 105 123 106 124
rect 104 123 105 124
rect 103 123 104 124
rect 102 123 103 124
rect 101 123 102 124
rect 100 123 101 124
rect 99 123 100 124
rect 98 123 99 124
rect 97 123 98 124
rect 96 123 97 124
rect 95 123 96 124
rect 94 123 95 124
rect 93 123 94 124
rect 92 123 93 124
rect 91 123 92 124
rect 90 123 91 124
rect 89 123 90 124
rect 88 123 89 124
rect 87 123 88 124
rect 86 123 87 124
rect 85 123 86 124
rect 84 123 85 124
rect 83 123 84 124
rect 82 123 83 124
rect 81 123 82 124
rect 80 123 81 124
rect 79 123 80 124
rect 78 123 79 124
rect 77 123 78 124
rect 76 123 77 124
rect 75 123 76 124
rect 74 123 75 124
rect 73 123 74 124
rect 72 123 73 124
rect 71 123 72 124
rect 70 123 71 124
rect 69 123 70 124
rect 68 123 69 124
rect 67 123 68 124
rect 66 123 67 124
rect 65 123 66 124
rect 64 123 65 124
rect 57 123 58 124
rect 56 123 57 124
rect 55 123 56 124
rect 54 123 55 124
rect 53 123 54 124
rect 52 123 53 124
rect 51 123 52 124
rect 50 123 51 124
rect 49 123 50 124
rect 48 123 49 124
rect 47 123 48 124
rect 46 123 47 124
rect 45 123 46 124
rect 44 123 45 124
rect 43 123 44 124
rect 42 123 43 124
rect 41 123 42 124
rect 40 123 41 124
rect 39 123 40 124
rect 38 123 39 124
rect 37 123 38 124
rect 36 123 37 124
rect 35 123 36 124
rect 34 123 35 124
rect 33 123 34 124
rect 32 123 33 124
rect 31 123 32 124
rect 30 123 31 124
rect 29 123 30 124
rect 28 123 29 124
rect 27 123 28 124
rect 475 124 476 125
rect 474 124 475 125
rect 473 124 474 125
rect 472 124 473 125
rect 471 124 472 125
rect 470 124 471 125
rect 469 124 470 125
rect 468 124 469 125
rect 458 124 459 125
rect 438 124 439 125
rect 437 124 438 125
rect 436 124 437 125
rect 435 124 436 125
rect 434 124 435 125
rect 295 124 296 125
rect 294 124 295 125
rect 293 124 294 125
rect 292 124 293 125
rect 291 124 292 125
rect 290 124 291 125
rect 289 124 290 125
rect 288 124 289 125
rect 287 124 288 125
rect 286 124 287 125
rect 285 124 286 125
rect 284 124 285 125
rect 283 124 284 125
rect 282 124 283 125
rect 281 124 282 125
rect 280 124 281 125
rect 279 124 280 125
rect 278 124 279 125
rect 277 124 278 125
rect 276 124 277 125
rect 275 124 276 125
rect 274 124 275 125
rect 273 124 274 125
rect 272 124 273 125
rect 271 124 272 125
rect 270 124 271 125
rect 269 124 270 125
rect 268 124 269 125
rect 267 124 268 125
rect 230 124 231 125
rect 229 124 230 125
rect 228 124 229 125
rect 227 124 228 125
rect 226 124 227 125
rect 225 124 226 125
rect 224 124 225 125
rect 223 124 224 125
rect 222 124 223 125
rect 221 124 222 125
rect 220 124 221 125
rect 219 124 220 125
rect 218 124 219 125
rect 217 124 218 125
rect 216 124 217 125
rect 215 124 216 125
rect 214 124 215 125
rect 213 124 214 125
rect 212 124 213 125
rect 211 124 212 125
rect 210 124 211 125
rect 209 124 210 125
rect 208 124 209 125
rect 207 124 208 125
rect 206 124 207 125
rect 205 124 206 125
rect 204 124 205 125
rect 203 124 204 125
rect 202 124 203 125
rect 201 124 202 125
rect 200 124 201 125
rect 199 124 200 125
rect 198 124 199 125
rect 197 124 198 125
rect 196 124 197 125
rect 195 124 196 125
rect 194 124 195 125
rect 193 124 194 125
rect 192 124 193 125
rect 191 124 192 125
rect 190 124 191 125
rect 189 124 190 125
rect 188 124 189 125
rect 187 124 188 125
rect 186 124 187 125
rect 185 124 186 125
rect 184 124 185 125
rect 183 124 184 125
rect 182 124 183 125
rect 181 124 182 125
rect 180 124 181 125
rect 179 124 180 125
rect 178 124 179 125
rect 177 124 178 125
rect 176 124 177 125
rect 175 124 176 125
rect 174 124 175 125
rect 173 124 174 125
rect 172 124 173 125
rect 171 124 172 125
rect 170 124 171 125
rect 169 124 170 125
rect 168 124 169 125
rect 167 124 168 125
rect 166 124 167 125
rect 165 124 166 125
rect 164 124 165 125
rect 147 124 148 125
rect 146 124 147 125
rect 145 124 146 125
rect 144 124 145 125
rect 143 124 144 125
rect 142 124 143 125
rect 141 124 142 125
rect 140 124 141 125
rect 139 124 140 125
rect 138 124 139 125
rect 137 124 138 125
rect 136 124 137 125
rect 135 124 136 125
rect 134 124 135 125
rect 133 124 134 125
rect 132 124 133 125
rect 131 124 132 125
rect 130 124 131 125
rect 129 124 130 125
rect 128 124 129 125
rect 127 124 128 125
rect 126 124 127 125
rect 125 124 126 125
rect 124 124 125 125
rect 123 124 124 125
rect 122 124 123 125
rect 121 124 122 125
rect 120 124 121 125
rect 119 124 120 125
rect 118 124 119 125
rect 117 124 118 125
rect 116 124 117 125
rect 115 124 116 125
rect 114 124 115 125
rect 113 124 114 125
rect 112 124 113 125
rect 111 124 112 125
rect 110 124 111 125
rect 109 124 110 125
rect 108 124 109 125
rect 107 124 108 125
rect 106 124 107 125
rect 105 124 106 125
rect 104 124 105 125
rect 103 124 104 125
rect 102 124 103 125
rect 101 124 102 125
rect 100 124 101 125
rect 99 124 100 125
rect 98 124 99 125
rect 97 124 98 125
rect 96 124 97 125
rect 95 124 96 125
rect 94 124 95 125
rect 93 124 94 125
rect 92 124 93 125
rect 91 124 92 125
rect 90 124 91 125
rect 89 124 90 125
rect 88 124 89 125
rect 87 124 88 125
rect 86 124 87 125
rect 85 124 86 125
rect 84 124 85 125
rect 83 124 84 125
rect 82 124 83 125
rect 81 124 82 125
rect 80 124 81 125
rect 79 124 80 125
rect 78 124 79 125
rect 77 124 78 125
rect 76 124 77 125
rect 75 124 76 125
rect 74 124 75 125
rect 73 124 74 125
rect 72 124 73 125
rect 71 124 72 125
rect 70 124 71 125
rect 69 124 70 125
rect 68 124 69 125
rect 67 124 68 125
rect 66 124 67 125
rect 65 124 66 125
rect 64 124 65 125
rect 63 124 64 125
rect 57 124 58 125
rect 56 124 57 125
rect 55 124 56 125
rect 54 124 55 125
rect 53 124 54 125
rect 52 124 53 125
rect 51 124 52 125
rect 50 124 51 125
rect 49 124 50 125
rect 48 124 49 125
rect 47 124 48 125
rect 46 124 47 125
rect 45 124 46 125
rect 44 124 45 125
rect 43 124 44 125
rect 42 124 43 125
rect 41 124 42 125
rect 40 124 41 125
rect 39 124 40 125
rect 38 124 39 125
rect 37 124 38 125
rect 36 124 37 125
rect 35 124 36 125
rect 34 124 35 125
rect 33 124 34 125
rect 32 124 33 125
rect 31 124 32 125
rect 30 124 31 125
rect 29 124 30 125
rect 28 124 29 125
rect 27 124 28 125
rect 476 125 477 126
rect 475 125 476 126
rect 474 125 475 126
rect 473 125 474 126
rect 472 125 473 126
rect 471 125 472 126
rect 470 125 471 126
rect 469 125 470 126
rect 458 125 459 126
rect 438 125 439 126
rect 437 125 438 126
rect 436 125 437 126
rect 435 125 436 126
rect 434 125 435 126
rect 297 125 298 126
rect 296 125 297 126
rect 295 125 296 126
rect 294 125 295 126
rect 293 125 294 126
rect 292 125 293 126
rect 291 125 292 126
rect 290 125 291 126
rect 289 125 290 126
rect 288 125 289 126
rect 287 125 288 126
rect 286 125 287 126
rect 285 125 286 126
rect 284 125 285 126
rect 283 125 284 126
rect 282 125 283 126
rect 281 125 282 126
rect 280 125 281 126
rect 279 125 280 126
rect 278 125 279 126
rect 277 125 278 126
rect 276 125 277 126
rect 275 125 276 126
rect 274 125 275 126
rect 273 125 274 126
rect 272 125 273 126
rect 271 125 272 126
rect 270 125 271 126
rect 269 125 270 126
rect 268 125 269 126
rect 267 125 268 126
rect 266 125 267 126
rect 265 125 266 126
rect 264 125 265 126
rect 229 125 230 126
rect 228 125 229 126
rect 227 125 228 126
rect 226 125 227 126
rect 225 125 226 126
rect 224 125 225 126
rect 223 125 224 126
rect 222 125 223 126
rect 221 125 222 126
rect 220 125 221 126
rect 219 125 220 126
rect 218 125 219 126
rect 217 125 218 126
rect 216 125 217 126
rect 215 125 216 126
rect 214 125 215 126
rect 213 125 214 126
rect 212 125 213 126
rect 211 125 212 126
rect 210 125 211 126
rect 209 125 210 126
rect 208 125 209 126
rect 207 125 208 126
rect 206 125 207 126
rect 205 125 206 126
rect 204 125 205 126
rect 203 125 204 126
rect 202 125 203 126
rect 201 125 202 126
rect 200 125 201 126
rect 199 125 200 126
rect 198 125 199 126
rect 197 125 198 126
rect 196 125 197 126
rect 195 125 196 126
rect 194 125 195 126
rect 193 125 194 126
rect 192 125 193 126
rect 191 125 192 126
rect 190 125 191 126
rect 189 125 190 126
rect 188 125 189 126
rect 187 125 188 126
rect 186 125 187 126
rect 185 125 186 126
rect 184 125 185 126
rect 183 125 184 126
rect 182 125 183 126
rect 181 125 182 126
rect 180 125 181 126
rect 179 125 180 126
rect 178 125 179 126
rect 177 125 178 126
rect 176 125 177 126
rect 175 125 176 126
rect 174 125 175 126
rect 173 125 174 126
rect 172 125 173 126
rect 171 125 172 126
rect 170 125 171 126
rect 169 125 170 126
rect 168 125 169 126
rect 167 125 168 126
rect 166 125 167 126
rect 165 125 166 126
rect 164 125 165 126
rect 146 125 147 126
rect 145 125 146 126
rect 144 125 145 126
rect 143 125 144 126
rect 142 125 143 126
rect 141 125 142 126
rect 140 125 141 126
rect 139 125 140 126
rect 138 125 139 126
rect 137 125 138 126
rect 136 125 137 126
rect 135 125 136 126
rect 134 125 135 126
rect 133 125 134 126
rect 132 125 133 126
rect 131 125 132 126
rect 130 125 131 126
rect 129 125 130 126
rect 128 125 129 126
rect 127 125 128 126
rect 126 125 127 126
rect 125 125 126 126
rect 124 125 125 126
rect 123 125 124 126
rect 122 125 123 126
rect 121 125 122 126
rect 120 125 121 126
rect 119 125 120 126
rect 118 125 119 126
rect 117 125 118 126
rect 116 125 117 126
rect 115 125 116 126
rect 114 125 115 126
rect 113 125 114 126
rect 112 125 113 126
rect 111 125 112 126
rect 110 125 111 126
rect 109 125 110 126
rect 108 125 109 126
rect 107 125 108 126
rect 106 125 107 126
rect 105 125 106 126
rect 104 125 105 126
rect 103 125 104 126
rect 102 125 103 126
rect 101 125 102 126
rect 100 125 101 126
rect 99 125 100 126
rect 98 125 99 126
rect 97 125 98 126
rect 96 125 97 126
rect 95 125 96 126
rect 94 125 95 126
rect 93 125 94 126
rect 92 125 93 126
rect 91 125 92 126
rect 90 125 91 126
rect 89 125 90 126
rect 88 125 89 126
rect 87 125 88 126
rect 86 125 87 126
rect 85 125 86 126
rect 84 125 85 126
rect 83 125 84 126
rect 82 125 83 126
rect 81 125 82 126
rect 80 125 81 126
rect 79 125 80 126
rect 78 125 79 126
rect 77 125 78 126
rect 76 125 77 126
rect 75 125 76 126
rect 74 125 75 126
rect 73 125 74 126
rect 72 125 73 126
rect 71 125 72 126
rect 70 125 71 126
rect 69 125 70 126
rect 68 125 69 126
rect 67 125 68 126
rect 66 125 67 126
rect 65 125 66 126
rect 64 125 65 126
rect 63 125 64 126
rect 57 125 58 126
rect 56 125 57 126
rect 55 125 56 126
rect 54 125 55 126
rect 53 125 54 126
rect 52 125 53 126
rect 51 125 52 126
rect 50 125 51 126
rect 49 125 50 126
rect 48 125 49 126
rect 47 125 48 126
rect 46 125 47 126
rect 45 125 46 126
rect 44 125 45 126
rect 43 125 44 126
rect 42 125 43 126
rect 41 125 42 126
rect 40 125 41 126
rect 39 125 40 126
rect 38 125 39 126
rect 37 125 38 126
rect 36 125 37 126
rect 35 125 36 126
rect 34 125 35 126
rect 33 125 34 126
rect 32 125 33 126
rect 31 125 32 126
rect 30 125 31 126
rect 29 125 30 126
rect 28 125 29 126
rect 477 126 478 127
rect 476 126 477 127
rect 475 126 476 127
rect 474 126 475 127
rect 473 126 474 127
rect 472 126 473 127
rect 471 126 472 127
rect 470 126 471 127
rect 458 126 459 127
rect 438 126 439 127
rect 437 126 438 127
rect 436 126 437 127
rect 435 126 436 127
rect 434 126 435 127
rect 298 126 299 127
rect 297 126 298 127
rect 296 126 297 127
rect 295 126 296 127
rect 294 126 295 127
rect 293 126 294 127
rect 292 126 293 127
rect 291 126 292 127
rect 290 126 291 127
rect 289 126 290 127
rect 288 126 289 127
rect 287 126 288 127
rect 286 126 287 127
rect 285 126 286 127
rect 284 126 285 127
rect 283 126 284 127
rect 282 126 283 127
rect 281 126 282 127
rect 280 126 281 127
rect 279 126 280 127
rect 278 126 279 127
rect 277 126 278 127
rect 276 126 277 127
rect 275 126 276 127
rect 274 126 275 127
rect 273 126 274 127
rect 272 126 273 127
rect 271 126 272 127
rect 270 126 271 127
rect 269 126 270 127
rect 268 126 269 127
rect 267 126 268 127
rect 266 126 267 127
rect 265 126 266 127
rect 264 126 265 127
rect 263 126 264 127
rect 262 126 263 127
rect 228 126 229 127
rect 227 126 228 127
rect 226 126 227 127
rect 225 126 226 127
rect 224 126 225 127
rect 223 126 224 127
rect 222 126 223 127
rect 221 126 222 127
rect 220 126 221 127
rect 219 126 220 127
rect 218 126 219 127
rect 217 126 218 127
rect 216 126 217 127
rect 215 126 216 127
rect 214 126 215 127
rect 213 126 214 127
rect 212 126 213 127
rect 211 126 212 127
rect 210 126 211 127
rect 209 126 210 127
rect 208 126 209 127
rect 207 126 208 127
rect 206 126 207 127
rect 205 126 206 127
rect 204 126 205 127
rect 203 126 204 127
rect 202 126 203 127
rect 201 126 202 127
rect 200 126 201 127
rect 199 126 200 127
rect 198 126 199 127
rect 197 126 198 127
rect 196 126 197 127
rect 195 126 196 127
rect 194 126 195 127
rect 193 126 194 127
rect 192 126 193 127
rect 191 126 192 127
rect 190 126 191 127
rect 189 126 190 127
rect 188 126 189 127
rect 187 126 188 127
rect 186 126 187 127
rect 185 126 186 127
rect 184 126 185 127
rect 183 126 184 127
rect 182 126 183 127
rect 181 126 182 127
rect 180 126 181 127
rect 179 126 180 127
rect 178 126 179 127
rect 177 126 178 127
rect 176 126 177 127
rect 175 126 176 127
rect 174 126 175 127
rect 173 126 174 127
rect 172 126 173 127
rect 171 126 172 127
rect 170 126 171 127
rect 169 126 170 127
rect 168 126 169 127
rect 167 126 168 127
rect 166 126 167 127
rect 165 126 166 127
rect 164 126 165 127
rect 163 126 164 127
rect 146 126 147 127
rect 145 126 146 127
rect 144 126 145 127
rect 143 126 144 127
rect 142 126 143 127
rect 141 126 142 127
rect 140 126 141 127
rect 139 126 140 127
rect 138 126 139 127
rect 137 126 138 127
rect 136 126 137 127
rect 135 126 136 127
rect 134 126 135 127
rect 133 126 134 127
rect 132 126 133 127
rect 131 126 132 127
rect 130 126 131 127
rect 129 126 130 127
rect 128 126 129 127
rect 127 126 128 127
rect 126 126 127 127
rect 125 126 126 127
rect 124 126 125 127
rect 123 126 124 127
rect 122 126 123 127
rect 121 126 122 127
rect 120 126 121 127
rect 119 126 120 127
rect 118 126 119 127
rect 117 126 118 127
rect 116 126 117 127
rect 115 126 116 127
rect 114 126 115 127
rect 113 126 114 127
rect 112 126 113 127
rect 111 126 112 127
rect 110 126 111 127
rect 109 126 110 127
rect 108 126 109 127
rect 107 126 108 127
rect 106 126 107 127
rect 105 126 106 127
rect 104 126 105 127
rect 103 126 104 127
rect 102 126 103 127
rect 101 126 102 127
rect 100 126 101 127
rect 99 126 100 127
rect 98 126 99 127
rect 97 126 98 127
rect 96 126 97 127
rect 95 126 96 127
rect 94 126 95 127
rect 93 126 94 127
rect 92 126 93 127
rect 91 126 92 127
rect 90 126 91 127
rect 89 126 90 127
rect 88 126 89 127
rect 87 126 88 127
rect 86 126 87 127
rect 85 126 86 127
rect 84 126 85 127
rect 83 126 84 127
rect 82 126 83 127
rect 81 126 82 127
rect 80 126 81 127
rect 79 126 80 127
rect 78 126 79 127
rect 77 126 78 127
rect 76 126 77 127
rect 75 126 76 127
rect 74 126 75 127
rect 73 126 74 127
rect 72 126 73 127
rect 71 126 72 127
rect 70 126 71 127
rect 69 126 70 127
rect 68 126 69 127
rect 67 126 68 127
rect 66 126 67 127
rect 65 126 66 127
rect 64 126 65 127
rect 63 126 64 127
rect 62 126 63 127
rect 57 126 58 127
rect 56 126 57 127
rect 55 126 56 127
rect 54 126 55 127
rect 53 126 54 127
rect 52 126 53 127
rect 51 126 52 127
rect 50 126 51 127
rect 49 126 50 127
rect 48 126 49 127
rect 47 126 48 127
rect 46 126 47 127
rect 45 126 46 127
rect 44 126 45 127
rect 43 126 44 127
rect 42 126 43 127
rect 41 126 42 127
rect 40 126 41 127
rect 39 126 40 127
rect 38 126 39 127
rect 37 126 38 127
rect 36 126 37 127
rect 35 126 36 127
rect 34 126 35 127
rect 33 126 34 127
rect 32 126 33 127
rect 31 126 32 127
rect 30 126 31 127
rect 29 126 30 127
rect 28 126 29 127
rect 478 127 479 128
rect 477 127 478 128
rect 476 127 477 128
rect 475 127 476 128
rect 474 127 475 128
rect 473 127 474 128
rect 472 127 473 128
rect 471 127 472 128
rect 460 127 461 128
rect 459 127 460 128
rect 458 127 459 128
rect 438 127 439 128
rect 437 127 438 128
rect 436 127 437 128
rect 435 127 436 128
rect 434 127 435 128
rect 300 127 301 128
rect 299 127 300 128
rect 298 127 299 128
rect 297 127 298 128
rect 296 127 297 128
rect 295 127 296 128
rect 294 127 295 128
rect 293 127 294 128
rect 292 127 293 128
rect 291 127 292 128
rect 290 127 291 128
rect 289 127 290 128
rect 288 127 289 128
rect 287 127 288 128
rect 286 127 287 128
rect 285 127 286 128
rect 284 127 285 128
rect 283 127 284 128
rect 282 127 283 128
rect 281 127 282 128
rect 280 127 281 128
rect 279 127 280 128
rect 278 127 279 128
rect 277 127 278 128
rect 276 127 277 128
rect 275 127 276 128
rect 274 127 275 128
rect 273 127 274 128
rect 272 127 273 128
rect 271 127 272 128
rect 270 127 271 128
rect 269 127 270 128
rect 268 127 269 128
rect 267 127 268 128
rect 266 127 267 128
rect 265 127 266 128
rect 264 127 265 128
rect 263 127 264 128
rect 262 127 263 128
rect 261 127 262 128
rect 260 127 261 128
rect 228 127 229 128
rect 227 127 228 128
rect 226 127 227 128
rect 225 127 226 128
rect 224 127 225 128
rect 223 127 224 128
rect 222 127 223 128
rect 221 127 222 128
rect 220 127 221 128
rect 219 127 220 128
rect 218 127 219 128
rect 217 127 218 128
rect 216 127 217 128
rect 215 127 216 128
rect 214 127 215 128
rect 213 127 214 128
rect 212 127 213 128
rect 211 127 212 128
rect 210 127 211 128
rect 209 127 210 128
rect 208 127 209 128
rect 207 127 208 128
rect 206 127 207 128
rect 205 127 206 128
rect 204 127 205 128
rect 203 127 204 128
rect 202 127 203 128
rect 201 127 202 128
rect 200 127 201 128
rect 199 127 200 128
rect 198 127 199 128
rect 197 127 198 128
rect 196 127 197 128
rect 195 127 196 128
rect 194 127 195 128
rect 193 127 194 128
rect 192 127 193 128
rect 191 127 192 128
rect 190 127 191 128
rect 189 127 190 128
rect 188 127 189 128
rect 187 127 188 128
rect 186 127 187 128
rect 185 127 186 128
rect 184 127 185 128
rect 183 127 184 128
rect 182 127 183 128
rect 181 127 182 128
rect 180 127 181 128
rect 179 127 180 128
rect 178 127 179 128
rect 177 127 178 128
rect 176 127 177 128
rect 175 127 176 128
rect 174 127 175 128
rect 173 127 174 128
rect 172 127 173 128
rect 171 127 172 128
rect 170 127 171 128
rect 169 127 170 128
rect 168 127 169 128
rect 167 127 168 128
rect 166 127 167 128
rect 165 127 166 128
rect 164 127 165 128
rect 163 127 164 128
rect 145 127 146 128
rect 144 127 145 128
rect 143 127 144 128
rect 142 127 143 128
rect 141 127 142 128
rect 140 127 141 128
rect 139 127 140 128
rect 138 127 139 128
rect 137 127 138 128
rect 136 127 137 128
rect 135 127 136 128
rect 134 127 135 128
rect 133 127 134 128
rect 132 127 133 128
rect 131 127 132 128
rect 130 127 131 128
rect 129 127 130 128
rect 128 127 129 128
rect 127 127 128 128
rect 126 127 127 128
rect 125 127 126 128
rect 124 127 125 128
rect 123 127 124 128
rect 122 127 123 128
rect 121 127 122 128
rect 120 127 121 128
rect 119 127 120 128
rect 118 127 119 128
rect 117 127 118 128
rect 116 127 117 128
rect 115 127 116 128
rect 114 127 115 128
rect 113 127 114 128
rect 112 127 113 128
rect 111 127 112 128
rect 110 127 111 128
rect 109 127 110 128
rect 108 127 109 128
rect 107 127 108 128
rect 106 127 107 128
rect 105 127 106 128
rect 104 127 105 128
rect 103 127 104 128
rect 102 127 103 128
rect 101 127 102 128
rect 100 127 101 128
rect 99 127 100 128
rect 98 127 99 128
rect 97 127 98 128
rect 96 127 97 128
rect 95 127 96 128
rect 94 127 95 128
rect 93 127 94 128
rect 92 127 93 128
rect 91 127 92 128
rect 90 127 91 128
rect 89 127 90 128
rect 88 127 89 128
rect 87 127 88 128
rect 86 127 87 128
rect 85 127 86 128
rect 84 127 85 128
rect 83 127 84 128
rect 82 127 83 128
rect 81 127 82 128
rect 80 127 81 128
rect 79 127 80 128
rect 78 127 79 128
rect 77 127 78 128
rect 76 127 77 128
rect 75 127 76 128
rect 74 127 75 128
rect 73 127 74 128
rect 72 127 73 128
rect 71 127 72 128
rect 70 127 71 128
rect 69 127 70 128
rect 68 127 69 128
rect 67 127 68 128
rect 66 127 67 128
rect 65 127 66 128
rect 64 127 65 128
rect 63 127 64 128
rect 62 127 63 128
rect 61 127 62 128
rect 57 127 58 128
rect 56 127 57 128
rect 55 127 56 128
rect 54 127 55 128
rect 53 127 54 128
rect 52 127 53 128
rect 51 127 52 128
rect 50 127 51 128
rect 49 127 50 128
rect 48 127 49 128
rect 47 127 48 128
rect 46 127 47 128
rect 45 127 46 128
rect 44 127 45 128
rect 43 127 44 128
rect 42 127 43 128
rect 41 127 42 128
rect 40 127 41 128
rect 39 127 40 128
rect 38 127 39 128
rect 37 127 38 128
rect 36 127 37 128
rect 35 127 36 128
rect 34 127 35 128
rect 33 127 34 128
rect 32 127 33 128
rect 31 127 32 128
rect 30 127 31 128
rect 29 127 30 128
rect 28 127 29 128
rect 479 128 480 129
rect 478 128 479 129
rect 477 128 478 129
rect 476 128 477 129
rect 475 128 476 129
rect 474 128 475 129
rect 473 128 474 129
rect 472 128 473 129
rect 471 128 472 129
rect 470 128 471 129
rect 469 128 470 129
rect 468 128 469 129
rect 467 128 468 129
rect 466 128 467 129
rect 465 128 466 129
rect 464 128 465 129
rect 463 128 464 129
rect 462 128 463 129
rect 461 128 462 129
rect 460 128 461 129
rect 459 128 460 129
rect 458 128 459 129
rect 438 128 439 129
rect 437 128 438 129
rect 436 128 437 129
rect 435 128 436 129
rect 434 128 435 129
rect 301 128 302 129
rect 300 128 301 129
rect 299 128 300 129
rect 298 128 299 129
rect 297 128 298 129
rect 296 128 297 129
rect 295 128 296 129
rect 294 128 295 129
rect 293 128 294 129
rect 292 128 293 129
rect 291 128 292 129
rect 290 128 291 129
rect 289 128 290 129
rect 288 128 289 129
rect 287 128 288 129
rect 286 128 287 129
rect 285 128 286 129
rect 284 128 285 129
rect 283 128 284 129
rect 282 128 283 129
rect 281 128 282 129
rect 280 128 281 129
rect 279 128 280 129
rect 278 128 279 129
rect 277 128 278 129
rect 276 128 277 129
rect 275 128 276 129
rect 274 128 275 129
rect 273 128 274 129
rect 272 128 273 129
rect 271 128 272 129
rect 270 128 271 129
rect 269 128 270 129
rect 268 128 269 129
rect 267 128 268 129
rect 266 128 267 129
rect 265 128 266 129
rect 264 128 265 129
rect 263 128 264 129
rect 262 128 263 129
rect 261 128 262 129
rect 260 128 261 129
rect 259 128 260 129
rect 258 128 259 129
rect 227 128 228 129
rect 226 128 227 129
rect 225 128 226 129
rect 224 128 225 129
rect 223 128 224 129
rect 222 128 223 129
rect 221 128 222 129
rect 220 128 221 129
rect 219 128 220 129
rect 218 128 219 129
rect 217 128 218 129
rect 216 128 217 129
rect 215 128 216 129
rect 214 128 215 129
rect 213 128 214 129
rect 212 128 213 129
rect 211 128 212 129
rect 210 128 211 129
rect 209 128 210 129
rect 208 128 209 129
rect 207 128 208 129
rect 206 128 207 129
rect 205 128 206 129
rect 204 128 205 129
rect 203 128 204 129
rect 202 128 203 129
rect 201 128 202 129
rect 200 128 201 129
rect 199 128 200 129
rect 198 128 199 129
rect 197 128 198 129
rect 196 128 197 129
rect 195 128 196 129
rect 194 128 195 129
rect 193 128 194 129
rect 192 128 193 129
rect 191 128 192 129
rect 190 128 191 129
rect 189 128 190 129
rect 188 128 189 129
rect 187 128 188 129
rect 186 128 187 129
rect 185 128 186 129
rect 184 128 185 129
rect 183 128 184 129
rect 182 128 183 129
rect 181 128 182 129
rect 180 128 181 129
rect 179 128 180 129
rect 178 128 179 129
rect 177 128 178 129
rect 176 128 177 129
rect 175 128 176 129
rect 174 128 175 129
rect 173 128 174 129
rect 172 128 173 129
rect 171 128 172 129
rect 170 128 171 129
rect 169 128 170 129
rect 168 128 169 129
rect 167 128 168 129
rect 166 128 167 129
rect 165 128 166 129
rect 164 128 165 129
rect 163 128 164 129
rect 162 128 163 129
rect 145 128 146 129
rect 144 128 145 129
rect 143 128 144 129
rect 142 128 143 129
rect 141 128 142 129
rect 140 128 141 129
rect 139 128 140 129
rect 138 128 139 129
rect 137 128 138 129
rect 136 128 137 129
rect 135 128 136 129
rect 134 128 135 129
rect 133 128 134 129
rect 132 128 133 129
rect 131 128 132 129
rect 130 128 131 129
rect 129 128 130 129
rect 128 128 129 129
rect 127 128 128 129
rect 126 128 127 129
rect 125 128 126 129
rect 124 128 125 129
rect 123 128 124 129
rect 122 128 123 129
rect 121 128 122 129
rect 120 128 121 129
rect 119 128 120 129
rect 118 128 119 129
rect 117 128 118 129
rect 116 128 117 129
rect 115 128 116 129
rect 114 128 115 129
rect 113 128 114 129
rect 112 128 113 129
rect 111 128 112 129
rect 110 128 111 129
rect 109 128 110 129
rect 108 128 109 129
rect 107 128 108 129
rect 106 128 107 129
rect 105 128 106 129
rect 104 128 105 129
rect 103 128 104 129
rect 102 128 103 129
rect 101 128 102 129
rect 100 128 101 129
rect 99 128 100 129
rect 98 128 99 129
rect 97 128 98 129
rect 96 128 97 129
rect 95 128 96 129
rect 94 128 95 129
rect 93 128 94 129
rect 92 128 93 129
rect 91 128 92 129
rect 90 128 91 129
rect 89 128 90 129
rect 88 128 89 129
rect 87 128 88 129
rect 86 128 87 129
rect 85 128 86 129
rect 84 128 85 129
rect 83 128 84 129
rect 82 128 83 129
rect 81 128 82 129
rect 80 128 81 129
rect 79 128 80 129
rect 78 128 79 129
rect 77 128 78 129
rect 76 128 77 129
rect 75 128 76 129
rect 74 128 75 129
rect 73 128 74 129
rect 72 128 73 129
rect 71 128 72 129
rect 70 128 71 129
rect 69 128 70 129
rect 68 128 69 129
rect 67 128 68 129
rect 66 128 67 129
rect 65 128 66 129
rect 64 128 65 129
rect 63 128 64 129
rect 62 128 63 129
rect 61 128 62 129
rect 56 128 57 129
rect 55 128 56 129
rect 54 128 55 129
rect 53 128 54 129
rect 52 128 53 129
rect 51 128 52 129
rect 50 128 51 129
rect 49 128 50 129
rect 48 128 49 129
rect 47 128 48 129
rect 46 128 47 129
rect 45 128 46 129
rect 44 128 45 129
rect 43 128 44 129
rect 42 128 43 129
rect 41 128 42 129
rect 40 128 41 129
rect 39 128 40 129
rect 38 128 39 129
rect 37 128 38 129
rect 36 128 37 129
rect 35 128 36 129
rect 34 128 35 129
rect 33 128 34 129
rect 32 128 33 129
rect 31 128 32 129
rect 30 128 31 129
rect 29 128 30 129
rect 479 129 480 130
rect 478 129 479 130
rect 477 129 478 130
rect 476 129 477 130
rect 475 129 476 130
rect 474 129 475 130
rect 473 129 474 130
rect 472 129 473 130
rect 471 129 472 130
rect 470 129 471 130
rect 469 129 470 130
rect 468 129 469 130
rect 467 129 468 130
rect 466 129 467 130
rect 465 129 466 130
rect 464 129 465 130
rect 463 129 464 130
rect 462 129 463 130
rect 461 129 462 130
rect 460 129 461 130
rect 459 129 460 130
rect 458 129 459 130
rect 438 129 439 130
rect 437 129 438 130
rect 436 129 437 130
rect 435 129 436 130
rect 434 129 435 130
rect 302 129 303 130
rect 301 129 302 130
rect 300 129 301 130
rect 299 129 300 130
rect 298 129 299 130
rect 297 129 298 130
rect 296 129 297 130
rect 295 129 296 130
rect 294 129 295 130
rect 293 129 294 130
rect 292 129 293 130
rect 291 129 292 130
rect 290 129 291 130
rect 289 129 290 130
rect 288 129 289 130
rect 287 129 288 130
rect 286 129 287 130
rect 285 129 286 130
rect 284 129 285 130
rect 283 129 284 130
rect 282 129 283 130
rect 281 129 282 130
rect 280 129 281 130
rect 279 129 280 130
rect 278 129 279 130
rect 277 129 278 130
rect 276 129 277 130
rect 275 129 276 130
rect 274 129 275 130
rect 273 129 274 130
rect 272 129 273 130
rect 271 129 272 130
rect 270 129 271 130
rect 269 129 270 130
rect 268 129 269 130
rect 267 129 268 130
rect 266 129 267 130
rect 265 129 266 130
rect 264 129 265 130
rect 263 129 264 130
rect 262 129 263 130
rect 261 129 262 130
rect 260 129 261 130
rect 259 129 260 130
rect 258 129 259 130
rect 257 129 258 130
rect 256 129 257 130
rect 226 129 227 130
rect 225 129 226 130
rect 224 129 225 130
rect 223 129 224 130
rect 222 129 223 130
rect 221 129 222 130
rect 220 129 221 130
rect 219 129 220 130
rect 218 129 219 130
rect 217 129 218 130
rect 216 129 217 130
rect 215 129 216 130
rect 214 129 215 130
rect 213 129 214 130
rect 212 129 213 130
rect 211 129 212 130
rect 210 129 211 130
rect 209 129 210 130
rect 208 129 209 130
rect 207 129 208 130
rect 206 129 207 130
rect 205 129 206 130
rect 204 129 205 130
rect 203 129 204 130
rect 202 129 203 130
rect 201 129 202 130
rect 200 129 201 130
rect 199 129 200 130
rect 198 129 199 130
rect 197 129 198 130
rect 196 129 197 130
rect 195 129 196 130
rect 194 129 195 130
rect 193 129 194 130
rect 192 129 193 130
rect 191 129 192 130
rect 190 129 191 130
rect 189 129 190 130
rect 188 129 189 130
rect 187 129 188 130
rect 186 129 187 130
rect 185 129 186 130
rect 184 129 185 130
rect 183 129 184 130
rect 182 129 183 130
rect 181 129 182 130
rect 180 129 181 130
rect 179 129 180 130
rect 178 129 179 130
rect 177 129 178 130
rect 176 129 177 130
rect 175 129 176 130
rect 174 129 175 130
rect 173 129 174 130
rect 172 129 173 130
rect 171 129 172 130
rect 170 129 171 130
rect 169 129 170 130
rect 168 129 169 130
rect 167 129 168 130
rect 166 129 167 130
rect 165 129 166 130
rect 164 129 165 130
rect 163 129 164 130
rect 162 129 163 130
rect 144 129 145 130
rect 143 129 144 130
rect 142 129 143 130
rect 141 129 142 130
rect 140 129 141 130
rect 139 129 140 130
rect 138 129 139 130
rect 137 129 138 130
rect 136 129 137 130
rect 135 129 136 130
rect 134 129 135 130
rect 133 129 134 130
rect 132 129 133 130
rect 131 129 132 130
rect 130 129 131 130
rect 129 129 130 130
rect 128 129 129 130
rect 127 129 128 130
rect 126 129 127 130
rect 125 129 126 130
rect 124 129 125 130
rect 123 129 124 130
rect 122 129 123 130
rect 121 129 122 130
rect 120 129 121 130
rect 119 129 120 130
rect 118 129 119 130
rect 117 129 118 130
rect 116 129 117 130
rect 115 129 116 130
rect 114 129 115 130
rect 113 129 114 130
rect 112 129 113 130
rect 111 129 112 130
rect 110 129 111 130
rect 109 129 110 130
rect 108 129 109 130
rect 107 129 108 130
rect 106 129 107 130
rect 105 129 106 130
rect 104 129 105 130
rect 103 129 104 130
rect 102 129 103 130
rect 101 129 102 130
rect 100 129 101 130
rect 99 129 100 130
rect 98 129 99 130
rect 97 129 98 130
rect 96 129 97 130
rect 95 129 96 130
rect 94 129 95 130
rect 93 129 94 130
rect 92 129 93 130
rect 91 129 92 130
rect 90 129 91 130
rect 89 129 90 130
rect 88 129 89 130
rect 87 129 88 130
rect 86 129 87 130
rect 85 129 86 130
rect 84 129 85 130
rect 83 129 84 130
rect 82 129 83 130
rect 81 129 82 130
rect 80 129 81 130
rect 79 129 80 130
rect 78 129 79 130
rect 77 129 78 130
rect 76 129 77 130
rect 75 129 76 130
rect 74 129 75 130
rect 73 129 74 130
rect 72 129 73 130
rect 71 129 72 130
rect 70 129 71 130
rect 69 129 70 130
rect 68 129 69 130
rect 67 129 68 130
rect 66 129 67 130
rect 65 129 66 130
rect 64 129 65 130
rect 63 129 64 130
rect 62 129 63 130
rect 61 129 62 130
rect 60 129 61 130
rect 56 129 57 130
rect 55 129 56 130
rect 54 129 55 130
rect 53 129 54 130
rect 52 129 53 130
rect 51 129 52 130
rect 50 129 51 130
rect 49 129 50 130
rect 48 129 49 130
rect 47 129 48 130
rect 46 129 47 130
rect 45 129 46 130
rect 44 129 45 130
rect 43 129 44 130
rect 42 129 43 130
rect 41 129 42 130
rect 40 129 41 130
rect 39 129 40 130
rect 38 129 39 130
rect 37 129 38 130
rect 36 129 37 130
rect 35 129 36 130
rect 34 129 35 130
rect 33 129 34 130
rect 32 129 33 130
rect 31 129 32 130
rect 30 129 31 130
rect 29 129 30 130
rect 459 130 460 131
rect 458 130 459 131
rect 438 130 439 131
rect 437 130 438 131
rect 436 130 437 131
rect 435 130 436 131
rect 434 130 435 131
rect 433 130 434 131
rect 394 130 395 131
rect 393 130 394 131
rect 304 130 305 131
rect 303 130 304 131
rect 302 130 303 131
rect 301 130 302 131
rect 300 130 301 131
rect 299 130 300 131
rect 298 130 299 131
rect 297 130 298 131
rect 296 130 297 131
rect 295 130 296 131
rect 294 130 295 131
rect 293 130 294 131
rect 292 130 293 131
rect 291 130 292 131
rect 290 130 291 131
rect 289 130 290 131
rect 288 130 289 131
rect 287 130 288 131
rect 286 130 287 131
rect 285 130 286 131
rect 284 130 285 131
rect 283 130 284 131
rect 282 130 283 131
rect 281 130 282 131
rect 280 130 281 131
rect 279 130 280 131
rect 278 130 279 131
rect 277 130 278 131
rect 276 130 277 131
rect 275 130 276 131
rect 274 130 275 131
rect 273 130 274 131
rect 272 130 273 131
rect 271 130 272 131
rect 270 130 271 131
rect 269 130 270 131
rect 268 130 269 131
rect 267 130 268 131
rect 266 130 267 131
rect 265 130 266 131
rect 264 130 265 131
rect 263 130 264 131
rect 262 130 263 131
rect 261 130 262 131
rect 260 130 261 131
rect 259 130 260 131
rect 258 130 259 131
rect 257 130 258 131
rect 256 130 257 131
rect 255 130 256 131
rect 225 130 226 131
rect 224 130 225 131
rect 223 130 224 131
rect 222 130 223 131
rect 221 130 222 131
rect 220 130 221 131
rect 219 130 220 131
rect 218 130 219 131
rect 217 130 218 131
rect 216 130 217 131
rect 215 130 216 131
rect 214 130 215 131
rect 213 130 214 131
rect 212 130 213 131
rect 211 130 212 131
rect 210 130 211 131
rect 209 130 210 131
rect 208 130 209 131
rect 207 130 208 131
rect 206 130 207 131
rect 205 130 206 131
rect 204 130 205 131
rect 203 130 204 131
rect 202 130 203 131
rect 201 130 202 131
rect 200 130 201 131
rect 199 130 200 131
rect 198 130 199 131
rect 197 130 198 131
rect 196 130 197 131
rect 195 130 196 131
rect 194 130 195 131
rect 193 130 194 131
rect 192 130 193 131
rect 191 130 192 131
rect 190 130 191 131
rect 189 130 190 131
rect 188 130 189 131
rect 187 130 188 131
rect 186 130 187 131
rect 185 130 186 131
rect 184 130 185 131
rect 183 130 184 131
rect 182 130 183 131
rect 181 130 182 131
rect 180 130 181 131
rect 179 130 180 131
rect 178 130 179 131
rect 177 130 178 131
rect 176 130 177 131
rect 175 130 176 131
rect 174 130 175 131
rect 173 130 174 131
rect 172 130 173 131
rect 171 130 172 131
rect 170 130 171 131
rect 169 130 170 131
rect 168 130 169 131
rect 167 130 168 131
rect 166 130 167 131
rect 165 130 166 131
rect 164 130 165 131
rect 163 130 164 131
rect 162 130 163 131
rect 144 130 145 131
rect 143 130 144 131
rect 142 130 143 131
rect 141 130 142 131
rect 140 130 141 131
rect 139 130 140 131
rect 138 130 139 131
rect 137 130 138 131
rect 136 130 137 131
rect 135 130 136 131
rect 134 130 135 131
rect 133 130 134 131
rect 132 130 133 131
rect 131 130 132 131
rect 130 130 131 131
rect 129 130 130 131
rect 128 130 129 131
rect 127 130 128 131
rect 126 130 127 131
rect 125 130 126 131
rect 124 130 125 131
rect 123 130 124 131
rect 122 130 123 131
rect 121 130 122 131
rect 120 130 121 131
rect 119 130 120 131
rect 118 130 119 131
rect 117 130 118 131
rect 116 130 117 131
rect 115 130 116 131
rect 114 130 115 131
rect 113 130 114 131
rect 112 130 113 131
rect 111 130 112 131
rect 110 130 111 131
rect 109 130 110 131
rect 108 130 109 131
rect 107 130 108 131
rect 106 130 107 131
rect 105 130 106 131
rect 104 130 105 131
rect 103 130 104 131
rect 102 130 103 131
rect 101 130 102 131
rect 100 130 101 131
rect 99 130 100 131
rect 98 130 99 131
rect 97 130 98 131
rect 96 130 97 131
rect 95 130 96 131
rect 94 130 95 131
rect 93 130 94 131
rect 92 130 93 131
rect 91 130 92 131
rect 90 130 91 131
rect 89 130 90 131
rect 88 130 89 131
rect 87 130 88 131
rect 86 130 87 131
rect 85 130 86 131
rect 84 130 85 131
rect 83 130 84 131
rect 82 130 83 131
rect 81 130 82 131
rect 80 130 81 131
rect 79 130 80 131
rect 78 130 79 131
rect 77 130 78 131
rect 76 130 77 131
rect 75 130 76 131
rect 74 130 75 131
rect 73 130 74 131
rect 72 130 73 131
rect 71 130 72 131
rect 70 130 71 131
rect 69 130 70 131
rect 68 130 69 131
rect 67 130 68 131
rect 66 130 67 131
rect 65 130 66 131
rect 64 130 65 131
rect 63 130 64 131
rect 62 130 63 131
rect 61 130 62 131
rect 60 130 61 131
rect 59 130 60 131
rect 56 130 57 131
rect 55 130 56 131
rect 54 130 55 131
rect 53 130 54 131
rect 52 130 53 131
rect 51 130 52 131
rect 50 130 51 131
rect 49 130 50 131
rect 48 130 49 131
rect 47 130 48 131
rect 46 130 47 131
rect 45 130 46 131
rect 44 130 45 131
rect 43 130 44 131
rect 42 130 43 131
rect 41 130 42 131
rect 40 130 41 131
rect 39 130 40 131
rect 38 130 39 131
rect 37 130 38 131
rect 36 130 37 131
rect 35 130 36 131
rect 34 130 35 131
rect 33 130 34 131
rect 32 130 33 131
rect 31 130 32 131
rect 30 130 31 131
rect 29 130 30 131
rect 458 131 459 132
rect 437 131 438 132
rect 436 131 437 132
rect 435 131 436 132
rect 434 131 435 132
rect 433 131 434 132
rect 395 131 396 132
rect 394 131 395 132
rect 393 131 394 132
rect 305 131 306 132
rect 304 131 305 132
rect 303 131 304 132
rect 302 131 303 132
rect 301 131 302 132
rect 300 131 301 132
rect 299 131 300 132
rect 298 131 299 132
rect 297 131 298 132
rect 296 131 297 132
rect 295 131 296 132
rect 294 131 295 132
rect 293 131 294 132
rect 292 131 293 132
rect 291 131 292 132
rect 290 131 291 132
rect 289 131 290 132
rect 288 131 289 132
rect 287 131 288 132
rect 286 131 287 132
rect 285 131 286 132
rect 284 131 285 132
rect 283 131 284 132
rect 282 131 283 132
rect 281 131 282 132
rect 280 131 281 132
rect 279 131 280 132
rect 278 131 279 132
rect 277 131 278 132
rect 276 131 277 132
rect 275 131 276 132
rect 274 131 275 132
rect 273 131 274 132
rect 272 131 273 132
rect 271 131 272 132
rect 270 131 271 132
rect 269 131 270 132
rect 268 131 269 132
rect 267 131 268 132
rect 266 131 267 132
rect 265 131 266 132
rect 264 131 265 132
rect 263 131 264 132
rect 262 131 263 132
rect 261 131 262 132
rect 260 131 261 132
rect 259 131 260 132
rect 258 131 259 132
rect 257 131 258 132
rect 256 131 257 132
rect 255 131 256 132
rect 254 131 255 132
rect 253 131 254 132
rect 225 131 226 132
rect 224 131 225 132
rect 223 131 224 132
rect 222 131 223 132
rect 221 131 222 132
rect 220 131 221 132
rect 219 131 220 132
rect 218 131 219 132
rect 217 131 218 132
rect 216 131 217 132
rect 215 131 216 132
rect 214 131 215 132
rect 213 131 214 132
rect 212 131 213 132
rect 211 131 212 132
rect 210 131 211 132
rect 209 131 210 132
rect 208 131 209 132
rect 207 131 208 132
rect 206 131 207 132
rect 205 131 206 132
rect 204 131 205 132
rect 203 131 204 132
rect 202 131 203 132
rect 201 131 202 132
rect 200 131 201 132
rect 199 131 200 132
rect 198 131 199 132
rect 197 131 198 132
rect 196 131 197 132
rect 195 131 196 132
rect 194 131 195 132
rect 193 131 194 132
rect 192 131 193 132
rect 191 131 192 132
rect 190 131 191 132
rect 189 131 190 132
rect 188 131 189 132
rect 187 131 188 132
rect 186 131 187 132
rect 185 131 186 132
rect 184 131 185 132
rect 183 131 184 132
rect 182 131 183 132
rect 181 131 182 132
rect 180 131 181 132
rect 179 131 180 132
rect 178 131 179 132
rect 177 131 178 132
rect 176 131 177 132
rect 175 131 176 132
rect 174 131 175 132
rect 173 131 174 132
rect 172 131 173 132
rect 171 131 172 132
rect 170 131 171 132
rect 169 131 170 132
rect 168 131 169 132
rect 167 131 168 132
rect 166 131 167 132
rect 165 131 166 132
rect 164 131 165 132
rect 163 131 164 132
rect 162 131 163 132
rect 161 131 162 132
rect 143 131 144 132
rect 142 131 143 132
rect 141 131 142 132
rect 140 131 141 132
rect 139 131 140 132
rect 138 131 139 132
rect 137 131 138 132
rect 136 131 137 132
rect 135 131 136 132
rect 134 131 135 132
rect 133 131 134 132
rect 132 131 133 132
rect 131 131 132 132
rect 130 131 131 132
rect 129 131 130 132
rect 128 131 129 132
rect 127 131 128 132
rect 126 131 127 132
rect 125 131 126 132
rect 124 131 125 132
rect 123 131 124 132
rect 122 131 123 132
rect 121 131 122 132
rect 120 131 121 132
rect 119 131 120 132
rect 118 131 119 132
rect 117 131 118 132
rect 116 131 117 132
rect 115 131 116 132
rect 114 131 115 132
rect 113 131 114 132
rect 112 131 113 132
rect 111 131 112 132
rect 110 131 111 132
rect 109 131 110 132
rect 108 131 109 132
rect 107 131 108 132
rect 106 131 107 132
rect 105 131 106 132
rect 104 131 105 132
rect 103 131 104 132
rect 102 131 103 132
rect 101 131 102 132
rect 100 131 101 132
rect 99 131 100 132
rect 98 131 99 132
rect 97 131 98 132
rect 96 131 97 132
rect 95 131 96 132
rect 94 131 95 132
rect 93 131 94 132
rect 92 131 93 132
rect 91 131 92 132
rect 90 131 91 132
rect 89 131 90 132
rect 88 131 89 132
rect 87 131 88 132
rect 86 131 87 132
rect 85 131 86 132
rect 84 131 85 132
rect 83 131 84 132
rect 82 131 83 132
rect 81 131 82 132
rect 80 131 81 132
rect 79 131 80 132
rect 78 131 79 132
rect 77 131 78 132
rect 76 131 77 132
rect 75 131 76 132
rect 74 131 75 132
rect 73 131 74 132
rect 72 131 73 132
rect 71 131 72 132
rect 70 131 71 132
rect 69 131 70 132
rect 68 131 69 132
rect 67 131 68 132
rect 66 131 67 132
rect 65 131 66 132
rect 64 131 65 132
rect 63 131 64 132
rect 62 131 63 132
rect 61 131 62 132
rect 60 131 61 132
rect 59 131 60 132
rect 56 131 57 132
rect 55 131 56 132
rect 54 131 55 132
rect 53 131 54 132
rect 52 131 53 132
rect 51 131 52 132
rect 50 131 51 132
rect 49 131 50 132
rect 48 131 49 132
rect 47 131 48 132
rect 46 131 47 132
rect 45 131 46 132
rect 44 131 45 132
rect 43 131 44 132
rect 42 131 43 132
rect 41 131 42 132
rect 40 131 41 132
rect 39 131 40 132
rect 38 131 39 132
rect 37 131 38 132
rect 36 131 37 132
rect 35 131 36 132
rect 34 131 35 132
rect 33 131 34 132
rect 32 131 33 132
rect 31 131 32 132
rect 30 131 31 132
rect 458 132 459 133
rect 437 132 438 133
rect 436 132 437 133
rect 435 132 436 133
rect 434 132 435 133
rect 433 132 434 133
rect 432 132 433 133
rect 395 132 396 133
rect 394 132 395 133
rect 393 132 394 133
rect 306 132 307 133
rect 305 132 306 133
rect 304 132 305 133
rect 303 132 304 133
rect 302 132 303 133
rect 301 132 302 133
rect 300 132 301 133
rect 299 132 300 133
rect 298 132 299 133
rect 297 132 298 133
rect 296 132 297 133
rect 295 132 296 133
rect 294 132 295 133
rect 293 132 294 133
rect 292 132 293 133
rect 291 132 292 133
rect 290 132 291 133
rect 289 132 290 133
rect 288 132 289 133
rect 287 132 288 133
rect 286 132 287 133
rect 285 132 286 133
rect 284 132 285 133
rect 283 132 284 133
rect 282 132 283 133
rect 281 132 282 133
rect 280 132 281 133
rect 279 132 280 133
rect 278 132 279 133
rect 277 132 278 133
rect 276 132 277 133
rect 275 132 276 133
rect 274 132 275 133
rect 273 132 274 133
rect 272 132 273 133
rect 271 132 272 133
rect 270 132 271 133
rect 269 132 270 133
rect 268 132 269 133
rect 267 132 268 133
rect 266 132 267 133
rect 265 132 266 133
rect 264 132 265 133
rect 263 132 264 133
rect 262 132 263 133
rect 261 132 262 133
rect 260 132 261 133
rect 259 132 260 133
rect 258 132 259 133
rect 257 132 258 133
rect 256 132 257 133
rect 255 132 256 133
rect 254 132 255 133
rect 253 132 254 133
rect 252 132 253 133
rect 224 132 225 133
rect 223 132 224 133
rect 222 132 223 133
rect 221 132 222 133
rect 220 132 221 133
rect 219 132 220 133
rect 218 132 219 133
rect 217 132 218 133
rect 216 132 217 133
rect 215 132 216 133
rect 214 132 215 133
rect 213 132 214 133
rect 212 132 213 133
rect 211 132 212 133
rect 210 132 211 133
rect 209 132 210 133
rect 208 132 209 133
rect 207 132 208 133
rect 206 132 207 133
rect 205 132 206 133
rect 204 132 205 133
rect 203 132 204 133
rect 202 132 203 133
rect 201 132 202 133
rect 200 132 201 133
rect 199 132 200 133
rect 198 132 199 133
rect 197 132 198 133
rect 196 132 197 133
rect 195 132 196 133
rect 194 132 195 133
rect 193 132 194 133
rect 192 132 193 133
rect 191 132 192 133
rect 190 132 191 133
rect 189 132 190 133
rect 188 132 189 133
rect 187 132 188 133
rect 186 132 187 133
rect 185 132 186 133
rect 184 132 185 133
rect 183 132 184 133
rect 182 132 183 133
rect 181 132 182 133
rect 180 132 181 133
rect 179 132 180 133
rect 178 132 179 133
rect 177 132 178 133
rect 176 132 177 133
rect 175 132 176 133
rect 174 132 175 133
rect 173 132 174 133
rect 172 132 173 133
rect 171 132 172 133
rect 170 132 171 133
rect 169 132 170 133
rect 168 132 169 133
rect 167 132 168 133
rect 166 132 167 133
rect 165 132 166 133
rect 164 132 165 133
rect 163 132 164 133
rect 162 132 163 133
rect 161 132 162 133
rect 143 132 144 133
rect 142 132 143 133
rect 141 132 142 133
rect 140 132 141 133
rect 139 132 140 133
rect 138 132 139 133
rect 137 132 138 133
rect 136 132 137 133
rect 135 132 136 133
rect 134 132 135 133
rect 133 132 134 133
rect 132 132 133 133
rect 131 132 132 133
rect 130 132 131 133
rect 129 132 130 133
rect 128 132 129 133
rect 127 132 128 133
rect 126 132 127 133
rect 125 132 126 133
rect 124 132 125 133
rect 123 132 124 133
rect 122 132 123 133
rect 121 132 122 133
rect 120 132 121 133
rect 119 132 120 133
rect 118 132 119 133
rect 117 132 118 133
rect 116 132 117 133
rect 115 132 116 133
rect 114 132 115 133
rect 113 132 114 133
rect 112 132 113 133
rect 111 132 112 133
rect 110 132 111 133
rect 109 132 110 133
rect 108 132 109 133
rect 107 132 108 133
rect 106 132 107 133
rect 105 132 106 133
rect 104 132 105 133
rect 103 132 104 133
rect 102 132 103 133
rect 101 132 102 133
rect 100 132 101 133
rect 99 132 100 133
rect 98 132 99 133
rect 97 132 98 133
rect 96 132 97 133
rect 95 132 96 133
rect 94 132 95 133
rect 93 132 94 133
rect 92 132 93 133
rect 91 132 92 133
rect 90 132 91 133
rect 89 132 90 133
rect 88 132 89 133
rect 87 132 88 133
rect 86 132 87 133
rect 85 132 86 133
rect 84 132 85 133
rect 83 132 84 133
rect 82 132 83 133
rect 81 132 82 133
rect 80 132 81 133
rect 79 132 80 133
rect 78 132 79 133
rect 77 132 78 133
rect 76 132 77 133
rect 75 132 76 133
rect 74 132 75 133
rect 73 132 74 133
rect 72 132 73 133
rect 71 132 72 133
rect 70 132 71 133
rect 69 132 70 133
rect 68 132 69 133
rect 67 132 68 133
rect 66 132 67 133
rect 65 132 66 133
rect 64 132 65 133
rect 63 132 64 133
rect 62 132 63 133
rect 61 132 62 133
rect 60 132 61 133
rect 59 132 60 133
rect 58 132 59 133
rect 56 132 57 133
rect 55 132 56 133
rect 54 132 55 133
rect 53 132 54 133
rect 52 132 53 133
rect 51 132 52 133
rect 50 132 51 133
rect 49 132 50 133
rect 48 132 49 133
rect 47 132 48 133
rect 46 132 47 133
rect 45 132 46 133
rect 44 132 45 133
rect 43 132 44 133
rect 42 132 43 133
rect 41 132 42 133
rect 40 132 41 133
rect 39 132 40 133
rect 38 132 39 133
rect 37 132 38 133
rect 36 132 37 133
rect 35 132 36 133
rect 34 132 35 133
rect 33 132 34 133
rect 32 132 33 133
rect 31 132 32 133
rect 437 133 438 134
rect 436 133 437 134
rect 435 133 436 134
rect 434 133 435 134
rect 433 133 434 134
rect 432 133 433 134
rect 431 133 432 134
rect 395 133 396 134
rect 394 133 395 134
rect 393 133 394 134
rect 307 133 308 134
rect 306 133 307 134
rect 305 133 306 134
rect 304 133 305 134
rect 303 133 304 134
rect 302 133 303 134
rect 301 133 302 134
rect 300 133 301 134
rect 299 133 300 134
rect 298 133 299 134
rect 297 133 298 134
rect 296 133 297 134
rect 295 133 296 134
rect 294 133 295 134
rect 293 133 294 134
rect 292 133 293 134
rect 291 133 292 134
rect 290 133 291 134
rect 289 133 290 134
rect 288 133 289 134
rect 287 133 288 134
rect 286 133 287 134
rect 285 133 286 134
rect 284 133 285 134
rect 283 133 284 134
rect 282 133 283 134
rect 281 133 282 134
rect 280 133 281 134
rect 279 133 280 134
rect 278 133 279 134
rect 277 133 278 134
rect 276 133 277 134
rect 275 133 276 134
rect 274 133 275 134
rect 273 133 274 134
rect 272 133 273 134
rect 271 133 272 134
rect 270 133 271 134
rect 269 133 270 134
rect 268 133 269 134
rect 267 133 268 134
rect 266 133 267 134
rect 265 133 266 134
rect 264 133 265 134
rect 263 133 264 134
rect 262 133 263 134
rect 261 133 262 134
rect 260 133 261 134
rect 259 133 260 134
rect 258 133 259 134
rect 257 133 258 134
rect 256 133 257 134
rect 255 133 256 134
rect 254 133 255 134
rect 253 133 254 134
rect 252 133 253 134
rect 251 133 252 134
rect 223 133 224 134
rect 222 133 223 134
rect 221 133 222 134
rect 220 133 221 134
rect 219 133 220 134
rect 218 133 219 134
rect 217 133 218 134
rect 216 133 217 134
rect 215 133 216 134
rect 214 133 215 134
rect 213 133 214 134
rect 212 133 213 134
rect 211 133 212 134
rect 210 133 211 134
rect 209 133 210 134
rect 208 133 209 134
rect 207 133 208 134
rect 206 133 207 134
rect 205 133 206 134
rect 204 133 205 134
rect 203 133 204 134
rect 202 133 203 134
rect 201 133 202 134
rect 200 133 201 134
rect 199 133 200 134
rect 198 133 199 134
rect 197 133 198 134
rect 196 133 197 134
rect 195 133 196 134
rect 194 133 195 134
rect 193 133 194 134
rect 192 133 193 134
rect 191 133 192 134
rect 190 133 191 134
rect 189 133 190 134
rect 188 133 189 134
rect 187 133 188 134
rect 186 133 187 134
rect 185 133 186 134
rect 184 133 185 134
rect 183 133 184 134
rect 182 133 183 134
rect 181 133 182 134
rect 180 133 181 134
rect 179 133 180 134
rect 178 133 179 134
rect 177 133 178 134
rect 176 133 177 134
rect 175 133 176 134
rect 174 133 175 134
rect 173 133 174 134
rect 172 133 173 134
rect 171 133 172 134
rect 170 133 171 134
rect 169 133 170 134
rect 168 133 169 134
rect 167 133 168 134
rect 166 133 167 134
rect 165 133 166 134
rect 164 133 165 134
rect 163 133 164 134
rect 162 133 163 134
rect 161 133 162 134
rect 160 133 161 134
rect 142 133 143 134
rect 141 133 142 134
rect 140 133 141 134
rect 139 133 140 134
rect 138 133 139 134
rect 137 133 138 134
rect 136 133 137 134
rect 135 133 136 134
rect 134 133 135 134
rect 133 133 134 134
rect 132 133 133 134
rect 131 133 132 134
rect 130 133 131 134
rect 129 133 130 134
rect 128 133 129 134
rect 127 133 128 134
rect 126 133 127 134
rect 125 133 126 134
rect 124 133 125 134
rect 123 133 124 134
rect 122 133 123 134
rect 121 133 122 134
rect 120 133 121 134
rect 119 133 120 134
rect 118 133 119 134
rect 117 133 118 134
rect 116 133 117 134
rect 115 133 116 134
rect 114 133 115 134
rect 113 133 114 134
rect 112 133 113 134
rect 111 133 112 134
rect 110 133 111 134
rect 109 133 110 134
rect 108 133 109 134
rect 107 133 108 134
rect 106 133 107 134
rect 105 133 106 134
rect 104 133 105 134
rect 103 133 104 134
rect 102 133 103 134
rect 101 133 102 134
rect 100 133 101 134
rect 99 133 100 134
rect 98 133 99 134
rect 97 133 98 134
rect 96 133 97 134
rect 95 133 96 134
rect 94 133 95 134
rect 93 133 94 134
rect 92 133 93 134
rect 91 133 92 134
rect 90 133 91 134
rect 89 133 90 134
rect 88 133 89 134
rect 87 133 88 134
rect 86 133 87 134
rect 85 133 86 134
rect 84 133 85 134
rect 83 133 84 134
rect 82 133 83 134
rect 81 133 82 134
rect 80 133 81 134
rect 79 133 80 134
rect 78 133 79 134
rect 77 133 78 134
rect 76 133 77 134
rect 75 133 76 134
rect 74 133 75 134
rect 73 133 74 134
rect 72 133 73 134
rect 71 133 72 134
rect 70 133 71 134
rect 69 133 70 134
rect 68 133 69 134
rect 67 133 68 134
rect 66 133 67 134
rect 65 133 66 134
rect 64 133 65 134
rect 63 133 64 134
rect 62 133 63 134
rect 61 133 62 134
rect 60 133 61 134
rect 59 133 60 134
rect 58 133 59 134
rect 57 133 58 134
rect 56 133 57 134
rect 55 133 56 134
rect 54 133 55 134
rect 53 133 54 134
rect 52 133 53 134
rect 51 133 52 134
rect 50 133 51 134
rect 49 133 50 134
rect 48 133 49 134
rect 47 133 48 134
rect 46 133 47 134
rect 45 133 46 134
rect 44 133 45 134
rect 43 133 44 134
rect 42 133 43 134
rect 41 133 42 134
rect 40 133 41 134
rect 39 133 40 134
rect 38 133 39 134
rect 37 133 38 134
rect 36 133 37 134
rect 35 133 36 134
rect 34 133 35 134
rect 33 133 34 134
rect 32 133 33 134
rect 31 133 32 134
rect 436 134 437 135
rect 435 134 436 135
rect 434 134 435 135
rect 433 134 434 135
rect 432 134 433 135
rect 431 134 432 135
rect 430 134 431 135
rect 396 134 397 135
rect 395 134 396 135
rect 394 134 395 135
rect 393 134 394 135
rect 308 134 309 135
rect 307 134 308 135
rect 306 134 307 135
rect 305 134 306 135
rect 304 134 305 135
rect 303 134 304 135
rect 302 134 303 135
rect 301 134 302 135
rect 300 134 301 135
rect 299 134 300 135
rect 298 134 299 135
rect 297 134 298 135
rect 296 134 297 135
rect 295 134 296 135
rect 294 134 295 135
rect 293 134 294 135
rect 292 134 293 135
rect 291 134 292 135
rect 290 134 291 135
rect 289 134 290 135
rect 288 134 289 135
rect 287 134 288 135
rect 286 134 287 135
rect 285 134 286 135
rect 284 134 285 135
rect 283 134 284 135
rect 282 134 283 135
rect 281 134 282 135
rect 280 134 281 135
rect 279 134 280 135
rect 278 134 279 135
rect 277 134 278 135
rect 276 134 277 135
rect 275 134 276 135
rect 274 134 275 135
rect 273 134 274 135
rect 272 134 273 135
rect 271 134 272 135
rect 270 134 271 135
rect 269 134 270 135
rect 268 134 269 135
rect 267 134 268 135
rect 266 134 267 135
rect 265 134 266 135
rect 264 134 265 135
rect 263 134 264 135
rect 262 134 263 135
rect 261 134 262 135
rect 260 134 261 135
rect 259 134 260 135
rect 258 134 259 135
rect 257 134 258 135
rect 256 134 257 135
rect 255 134 256 135
rect 254 134 255 135
rect 253 134 254 135
rect 252 134 253 135
rect 251 134 252 135
rect 250 134 251 135
rect 249 134 250 135
rect 223 134 224 135
rect 222 134 223 135
rect 221 134 222 135
rect 220 134 221 135
rect 219 134 220 135
rect 218 134 219 135
rect 217 134 218 135
rect 216 134 217 135
rect 215 134 216 135
rect 214 134 215 135
rect 213 134 214 135
rect 212 134 213 135
rect 211 134 212 135
rect 210 134 211 135
rect 209 134 210 135
rect 208 134 209 135
rect 207 134 208 135
rect 206 134 207 135
rect 205 134 206 135
rect 204 134 205 135
rect 203 134 204 135
rect 202 134 203 135
rect 201 134 202 135
rect 200 134 201 135
rect 199 134 200 135
rect 198 134 199 135
rect 197 134 198 135
rect 196 134 197 135
rect 195 134 196 135
rect 194 134 195 135
rect 193 134 194 135
rect 192 134 193 135
rect 191 134 192 135
rect 190 134 191 135
rect 189 134 190 135
rect 188 134 189 135
rect 187 134 188 135
rect 186 134 187 135
rect 185 134 186 135
rect 184 134 185 135
rect 183 134 184 135
rect 182 134 183 135
rect 181 134 182 135
rect 180 134 181 135
rect 179 134 180 135
rect 178 134 179 135
rect 177 134 178 135
rect 176 134 177 135
rect 175 134 176 135
rect 174 134 175 135
rect 173 134 174 135
rect 172 134 173 135
rect 171 134 172 135
rect 170 134 171 135
rect 169 134 170 135
rect 168 134 169 135
rect 167 134 168 135
rect 166 134 167 135
rect 165 134 166 135
rect 164 134 165 135
rect 163 134 164 135
rect 162 134 163 135
rect 161 134 162 135
rect 160 134 161 135
rect 141 134 142 135
rect 140 134 141 135
rect 139 134 140 135
rect 138 134 139 135
rect 137 134 138 135
rect 136 134 137 135
rect 135 134 136 135
rect 134 134 135 135
rect 133 134 134 135
rect 132 134 133 135
rect 131 134 132 135
rect 130 134 131 135
rect 129 134 130 135
rect 128 134 129 135
rect 127 134 128 135
rect 126 134 127 135
rect 125 134 126 135
rect 124 134 125 135
rect 123 134 124 135
rect 122 134 123 135
rect 121 134 122 135
rect 120 134 121 135
rect 119 134 120 135
rect 118 134 119 135
rect 117 134 118 135
rect 116 134 117 135
rect 115 134 116 135
rect 114 134 115 135
rect 113 134 114 135
rect 112 134 113 135
rect 111 134 112 135
rect 110 134 111 135
rect 109 134 110 135
rect 108 134 109 135
rect 107 134 108 135
rect 106 134 107 135
rect 105 134 106 135
rect 104 134 105 135
rect 103 134 104 135
rect 102 134 103 135
rect 101 134 102 135
rect 100 134 101 135
rect 99 134 100 135
rect 98 134 99 135
rect 97 134 98 135
rect 96 134 97 135
rect 95 134 96 135
rect 94 134 95 135
rect 93 134 94 135
rect 92 134 93 135
rect 91 134 92 135
rect 90 134 91 135
rect 89 134 90 135
rect 88 134 89 135
rect 87 134 88 135
rect 86 134 87 135
rect 85 134 86 135
rect 84 134 85 135
rect 83 134 84 135
rect 82 134 83 135
rect 81 134 82 135
rect 80 134 81 135
rect 79 134 80 135
rect 78 134 79 135
rect 77 134 78 135
rect 76 134 77 135
rect 75 134 76 135
rect 74 134 75 135
rect 73 134 74 135
rect 72 134 73 135
rect 71 134 72 135
rect 70 134 71 135
rect 69 134 70 135
rect 68 134 69 135
rect 67 134 68 135
rect 66 134 67 135
rect 65 134 66 135
rect 64 134 65 135
rect 63 134 64 135
rect 62 134 63 135
rect 61 134 62 135
rect 60 134 61 135
rect 59 134 60 135
rect 58 134 59 135
rect 57 134 58 135
rect 56 134 57 135
rect 55 134 56 135
rect 54 134 55 135
rect 53 134 54 135
rect 52 134 53 135
rect 51 134 52 135
rect 50 134 51 135
rect 49 134 50 135
rect 48 134 49 135
rect 47 134 48 135
rect 46 134 47 135
rect 45 134 46 135
rect 44 134 45 135
rect 43 134 44 135
rect 42 134 43 135
rect 41 134 42 135
rect 40 134 41 135
rect 39 134 40 135
rect 38 134 39 135
rect 37 134 38 135
rect 36 134 37 135
rect 35 134 36 135
rect 34 134 35 135
rect 33 134 34 135
rect 32 134 33 135
rect 436 135 437 136
rect 435 135 436 136
rect 434 135 435 136
rect 433 135 434 136
rect 432 135 433 136
rect 431 135 432 136
rect 430 135 431 136
rect 429 135 430 136
rect 428 135 429 136
rect 427 135 428 136
rect 397 135 398 136
rect 396 135 397 136
rect 395 135 396 136
rect 394 135 395 136
rect 393 135 394 136
rect 308 135 309 136
rect 307 135 308 136
rect 306 135 307 136
rect 305 135 306 136
rect 304 135 305 136
rect 303 135 304 136
rect 302 135 303 136
rect 301 135 302 136
rect 300 135 301 136
rect 299 135 300 136
rect 298 135 299 136
rect 297 135 298 136
rect 296 135 297 136
rect 295 135 296 136
rect 294 135 295 136
rect 293 135 294 136
rect 292 135 293 136
rect 291 135 292 136
rect 290 135 291 136
rect 289 135 290 136
rect 288 135 289 136
rect 287 135 288 136
rect 286 135 287 136
rect 285 135 286 136
rect 284 135 285 136
rect 283 135 284 136
rect 282 135 283 136
rect 281 135 282 136
rect 280 135 281 136
rect 279 135 280 136
rect 278 135 279 136
rect 277 135 278 136
rect 276 135 277 136
rect 275 135 276 136
rect 274 135 275 136
rect 273 135 274 136
rect 272 135 273 136
rect 271 135 272 136
rect 270 135 271 136
rect 269 135 270 136
rect 268 135 269 136
rect 267 135 268 136
rect 266 135 267 136
rect 265 135 266 136
rect 264 135 265 136
rect 263 135 264 136
rect 262 135 263 136
rect 261 135 262 136
rect 260 135 261 136
rect 259 135 260 136
rect 258 135 259 136
rect 257 135 258 136
rect 256 135 257 136
rect 255 135 256 136
rect 254 135 255 136
rect 253 135 254 136
rect 252 135 253 136
rect 251 135 252 136
rect 250 135 251 136
rect 249 135 250 136
rect 248 135 249 136
rect 222 135 223 136
rect 221 135 222 136
rect 220 135 221 136
rect 219 135 220 136
rect 218 135 219 136
rect 217 135 218 136
rect 216 135 217 136
rect 215 135 216 136
rect 214 135 215 136
rect 213 135 214 136
rect 212 135 213 136
rect 211 135 212 136
rect 210 135 211 136
rect 209 135 210 136
rect 208 135 209 136
rect 207 135 208 136
rect 206 135 207 136
rect 205 135 206 136
rect 204 135 205 136
rect 203 135 204 136
rect 202 135 203 136
rect 201 135 202 136
rect 200 135 201 136
rect 199 135 200 136
rect 198 135 199 136
rect 197 135 198 136
rect 196 135 197 136
rect 195 135 196 136
rect 194 135 195 136
rect 193 135 194 136
rect 192 135 193 136
rect 191 135 192 136
rect 190 135 191 136
rect 189 135 190 136
rect 188 135 189 136
rect 187 135 188 136
rect 186 135 187 136
rect 185 135 186 136
rect 184 135 185 136
rect 183 135 184 136
rect 182 135 183 136
rect 181 135 182 136
rect 180 135 181 136
rect 179 135 180 136
rect 178 135 179 136
rect 177 135 178 136
rect 176 135 177 136
rect 175 135 176 136
rect 174 135 175 136
rect 173 135 174 136
rect 172 135 173 136
rect 171 135 172 136
rect 170 135 171 136
rect 169 135 170 136
rect 168 135 169 136
rect 167 135 168 136
rect 166 135 167 136
rect 165 135 166 136
rect 164 135 165 136
rect 163 135 164 136
rect 162 135 163 136
rect 161 135 162 136
rect 160 135 161 136
rect 159 135 160 136
rect 141 135 142 136
rect 140 135 141 136
rect 139 135 140 136
rect 138 135 139 136
rect 137 135 138 136
rect 136 135 137 136
rect 135 135 136 136
rect 134 135 135 136
rect 133 135 134 136
rect 132 135 133 136
rect 131 135 132 136
rect 130 135 131 136
rect 129 135 130 136
rect 128 135 129 136
rect 127 135 128 136
rect 126 135 127 136
rect 125 135 126 136
rect 124 135 125 136
rect 123 135 124 136
rect 122 135 123 136
rect 121 135 122 136
rect 120 135 121 136
rect 119 135 120 136
rect 118 135 119 136
rect 117 135 118 136
rect 116 135 117 136
rect 115 135 116 136
rect 114 135 115 136
rect 113 135 114 136
rect 112 135 113 136
rect 111 135 112 136
rect 110 135 111 136
rect 109 135 110 136
rect 108 135 109 136
rect 107 135 108 136
rect 106 135 107 136
rect 105 135 106 136
rect 104 135 105 136
rect 103 135 104 136
rect 102 135 103 136
rect 101 135 102 136
rect 100 135 101 136
rect 99 135 100 136
rect 98 135 99 136
rect 97 135 98 136
rect 96 135 97 136
rect 95 135 96 136
rect 94 135 95 136
rect 93 135 94 136
rect 92 135 93 136
rect 91 135 92 136
rect 90 135 91 136
rect 89 135 90 136
rect 88 135 89 136
rect 87 135 88 136
rect 86 135 87 136
rect 85 135 86 136
rect 84 135 85 136
rect 83 135 84 136
rect 82 135 83 136
rect 81 135 82 136
rect 80 135 81 136
rect 79 135 80 136
rect 78 135 79 136
rect 77 135 78 136
rect 76 135 77 136
rect 75 135 76 136
rect 74 135 75 136
rect 73 135 74 136
rect 72 135 73 136
rect 71 135 72 136
rect 70 135 71 136
rect 69 135 70 136
rect 68 135 69 136
rect 67 135 68 136
rect 66 135 67 136
rect 65 135 66 136
rect 64 135 65 136
rect 63 135 64 136
rect 62 135 63 136
rect 61 135 62 136
rect 60 135 61 136
rect 59 135 60 136
rect 58 135 59 136
rect 57 135 58 136
rect 56 135 57 136
rect 55 135 56 136
rect 54 135 55 136
rect 53 135 54 136
rect 52 135 53 136
rect 51 135 52 136
rect 50 135 51 136
rect 49 135 50 136
rect 48 135 49 136
rect 47 135 48 136
rect 46 135 47 136
rect 45 135 46 136
rect 44 135 45 136
rect 43 135 44 136
rect 42 135 43 136
rect 41 135 42 136
rect 40 135 41 136
rect 39 135 40 136
rect 38 135 39 136
rect 37 135 38 136
rect 36 135 37 136
rect 35 135 36 136
rect 34 135 35 136
rect 33 135 34 136
rect 435 136 436 137
rect 434 136 435 137
rect 433 136 434 137
rect 432 136 433 137
rect 431 136 432 137
rect 430 136 431 137
rect 429 136 430 137
rect 428 136 429 137
rect 427 136 428 137
rect 426 136 427 137
rect 425 136 426 137
rect 424 136 425 137
rect 423 136 424 137
rect 422 136 423 137
rect 403 136 404 137
rect 402 136 403 137
rect 401 136 402 137
rect 400 136 401 137
rect 399 136 400 137
rect 398 136 399 137
rect 397 136 398 137
rect 396 136 397 137
rect 395 136 396 137
rect 394 136 395 137
rect 393 136 394 137
rect 309 136 310 137
rect 308 136 309 137
rect 307 136 308 137
rect 306 136 307 137
rect 305 136 306 137
rect 304 136 305 137
rect 303 136 304 137
rect 302 136 303 137
rect 301 136 302 137
rect 300 136 301 137
rect 299 136 300 137
rect 298 136 299 137
rect 297 136 298 137
rect 296 136 297 137
rect 295 136 296 137
rect 294 136 295 137
rect 293 136 294 137
rect 292 136 293 137
rect 291 136 292 137
rect 290 136 291 137
rect 289 136 290 137
rect 288 136 289 137
rect 287 136 288 137
rect 286 136 287 137
rect 285 136 286 137
rect 284 136 285 137
rect 283 136 284 137
rect 282 136 283 137
rect 281 136 282 137
rect 280 136 281 137
rect 279 136 280 137
rect 278 136 279 137
rect 277 136 278 137
rect 276 136 277 137
rect 275 136 276 137
rect 274 136 275 137
rect 273 136 274 137
rect 272 136 273 137
rect 271 136 272 137
rect 270 136 271 137
rect 269 136 270 137
rect 268 136 269 137
rect 267 136 268 137
rect 266 136 267 137
rect 265 136 266 137
rect 264 136 265 137
rect 263 136 264 137
rect 262 136 263 137
rect 261 136 262 137
rect 260 136 261 137
rect 259 136 260 137
rect 258 136 259 137
rect 257 136 258 137
rect 256 136 257 137
rect 255 136 256 137
rect 254 136 255 137
rect 253 136 254 137
rect 252 136 253 137
rect 251 136 252 137
rect 250 136 251 137
rect 249 136 250 137
rect 248 136 249 137
rect 247 136 248 137
rect 222 136 223 137
rect 221 136 222 137
rect 220 136 221 137
rect 219 136 220 137
rect 218 136 219 137
rect 217 136 218 137
rect 216 136 217 137
rect 215 136 216 137
rect 214 136 215 137
rect 213 136 214 137
rect 212 136 213 137
rect 211 136 212 137
rect 210 136 211 137
rect 209 136 210 137
rect 208 136 209 137
rect 207 136 208 137
rect 206 136 207 137
rect 205 136 206 137
rect 204 136 205 137
rect 203 136 204 137
rect 202 136 203 137
rect 201 136 202 137
rect 200 136 201 137
rect 199 136 200 137
rect 198 136 199 137
rect 197 136 198 137
rect 196 136 197 137
rect 195 136 196 137
rect 194 136 195 137
rect 193 136 194 137
rect 192 136 193 137
rect 191 136 192 137
rect 190 136 191 137
rect 189 136 190 137
rect 188 136 189 137
rect 187 136 188 137
rect 186 136 187 137
rect 185 136 186 137
rect 184 136 185 137
rect 183 136 184 137
rect 182 136 183 137
rect 181 136 182 137
rect 180 136 181 137
rect 179 136 180 137
rect 178 136 179 137
rect 177 136 178 137
rect 176 136 177 137
rect 175 136 176 137
rect 174 136 175 137
rect 173 136 174 137
rect 172 136 173 137
rect 171 136 172 137
rect 170 136 171 137
rect 169 136 170 137
rect 168 136 169 137
rect 167 136 168 137
rect 166 136 167 137
rect 165 136 166 137
rect 164 136 165 137
rect 163 136 164 137
rect 162 136 163 137
rect 161 136 162 137
rect 160 136 161 137
rect 159 136 160 137
rect 140 136 141 137
rect 139 136 140 137
rect 138 136 139 137
rect 137 136 138 137
rect 136 136 137 137
rect 135 136 136 137
rect 134 136 135 137
rect 133 136 134 137
rect 132 136 133 137
rect 131 136 132 137
rect 130 136 131 137
rect 129 136 130 137
rect 128 136 129 137
rect 127 136 128 137
rect 126 136 127 137
rect 125 136 126 137
rect 124 136 125 137
rect 123 136 124 137
rect 122 136 123 137
rect 121 136 122 137
rect 120 136 121 137
rect 119 136 120 137
rect 118 136 119 137
rect 117 136 118 137
rect 116 136 117 137
rect 115 136 116 137
rect 114 136 115 137
rect 113 136 114 137
rect 112 136 113 137
rect 111 136 112 137
rect 110 136 111 137
rect 109 136 110 137
rect 108 136 109 137
rect 107 136 108 137
rect 106 136 107 137
rect 105 136 106 137
rect 104 136 105 137
rect 103 136 104 137
rect 102 136 103 137
rect 101 136 102 137
rect 100 136 101 137
rect 99 136 100 137
rect 98 136 99 137
rect 97 136 98 137
rect 96 136 97 137
rect 95 136 96 137
rect 94 136 95 137
rect 93 136 94 137
rect 92 136 93 137
rect 91 136 92 137
rect 90 136 91 137
rect 89 136 90 137
rect 88 136 89 137
rect 87 136 88 137
rect 86 136 87 137
rect 85 136 86 137
rect 84 136 85 137
rect 83 136 84 137
rect 82 136 83 137
rect 81 136 82 137
rect 80 136 81 137
rect 79 136 80 137
rect 78 136 79 137
rect 77 136 78 137
rect 76 136 77 137
rect 75 136 76 137
rect 74 136 75 137
rect 73 136 74 137
rect 72 136 73 137
rect 71 136 72 137
rect 70 136 71 137
rect 69 136 70 137
rect 68 136 69 137
rect 67 136 68 137
rect 66 136 67 137
rect 65 136 66 137
rect 64 136 65 137
rect 63 136 64 137
rect 62 136 63 137
rect 61 136 62 137
rect 60 136 61 137
rect 59 136 60 137
rect 58 136 59 137
rect 57 136 58 137
rect 56 136 57 137
rect 55 136 56 137
rect 54 136 55 137
rect 53 136 54 137
rect 52 136 53 137
rect 51 136 52 137
rect 50 136 51 137
rect 49 136 50 137
rect 48 136 49 137
rect 47 136 48 137
rect 46 136 47 137
rect 45 136 46 137
rect 44 136 45 137
rect 43 136 44 137
rect 42 136 43 137
rect 41 136 42 137
rect 40 136 41 137
rect 39 136 40 137
rect 38 136 39 137
rect 37 136 38 137
rect 36 136 37 137
rect 35 136 36 137
rect 34 136 35 137
rect 434 137 435 138
rect 433 137 434 138
rect 432 137 433 138
rect 431 137 432 138
rect 430 137 431 138
rect 429 137 430 138
rect 428 137 429 138
rect 427 137 428 138
rect 426 137 427 138
rect 425 137 426 138
rect 424 137 425 138
rect 423 137 424 138
rect 422 137 423 138
rect 421 137 422 138
rect 420 137 421 138
rect 419 137 420 138
rect 418 137 419 138
rect 417 137 418 138
rect 416 137 417 138
rect 415 137 416 138
rect 414 137 415 138
rect 413 137 414 138
rect 412 137 413 138
rect 411 137 412 138
rect 410 137 411 138
rect 409 137 410 138
rect 408 137 409 138
rect 407 137 408 138
rect 406 137 407 138
rect 405 137 406 138
rect 404 137 405 138
rect 403 137 404 138
rect 402 137 403 138
rect 401 137 402 138
rect 400 137 401 138
rect 399 137 400 138
rect 398 137 399 138
rect 397 137 398 138
rect 396 137 397 138
rect 395 137 396 138
rect 394 137 395 138
rect 393 137 394 138
rect 310 137 311 138
rect 309 137 310 138
rect 308 137 309 138
rect 307 137 308 138
rect 306 137 307 138
rect 305 137 306 138
rect 304 137 305 138
rect 303 137 304 138
rect 302 137 303 138
rect 301 137 302 138
rect 300 137 301 138
rect 299 137 300 138
rect 298 137 299 138
rect 297 137 298 138
rect 296 137 297 138
rect 295 137 296 138
rect 294 137 295 138
rect 293 137 294 138
rect 292 137 293 138
rect 291 137 292 138
rect 290 137 291 138
rect 289 137 290 138
rect 288 137 289 138
rect 287 137 288 138
rect 286 137 287 138
rect 285 137 286 138
rect 284 137 285 138
rect 283 137 284 138
rect 282 137 283 138
rect 281 137 282 138
rect 280 137 281 138
rect 279 137 280 138
rect 278 137 279 138
rect 277 137 278 138
rect 276 137 277 138
rect 275 137 276 138
rect 274 137 275 138
rect 273 137 274 138
rect 272 137 273 138
rect 271 137 272 138
rect 270 137 271 138
rect 269 137 270 138
rect 268 137 269 138
rect 267 137 268 138
rect 266 137 267 138
rect 265 137 266 138
rect 264 137 265 138
rect 263 137 264 138
rect 262 137 263 138
rect 261 137 262 138
rect 260 137 261 138
rect 259 137 260 138
rect 258 137 259 138
rect 257 137 258 138
rect 256 137 257 138
rect 255 137 256 138
rect 254 137 255 138
rect 253 137 254 138
rect 252 137 253 138
rect 251 137 252 138
rect 250 137 251 138
rect 249 137 250 138
rect 248 137 249 138
rect 247 137 248 138
rect 246 137 247 138
rect 221 137 222 138
rect 220 137 221 138
rect 219 137 220 138
rect 218 137 219 138
rect 217 137 218 138
rect 216 137 217 138
rect 215 137 216 138
rect 214 137 215 138
rect 213 137 214 138
rect 212 137 213 138
rect 211 137 212 138
rect 210 137 211 138
rect 209 137 210 138
rect 208 137 209 138
rect 207 137 208 138
rect 206 137 207 138
rect 205 137 206 138
rect 204 137 205 138
rect 203 137 204 138
rect 202 137 203 138
rect 201 137 202 138
rect 200 137 201 138
rect 199 137 200 138
rect 198 137 199 138
rect 197 137 198 138
rect 196 137 197 138
rect 195 137 196 138
rect 194 137 195 138
rect 193 137 194 138
rect 192 137 193 138
rect 191 137 192 138
rect 190 137 191 138
rect 189 137 190 138
rect 188 137 189 138
rect 187 137 188 138
rect 186 137 187 138
rect 185 137 186 138
rect 184 137 185 138
rect 183 137 184 138
rect 182 137 183 138
rect 181 137 182 138
rect 180 137 181 138
rect 179 137 180 138
rect 178 137 179 138
rect 177 137 178 138
rect 176 137 177 138
rect 175 137 176 138
rect 174 137 175 138
rect 173 137 174 138
rect 172 137 173 138
rect 171 137 172 138
rect 170 137 171 138
rect 169 137 170 138
rect 168 137 169 138
rect 167 137 168 138
rect 166 137 167 138
rect 165 137 166 138
rect 164 137 165 138
rect 163 137 164 138
rect 162 137 163 138
rect 161 137 162 138
rect 160 137 161 138
rect 159 137 160 138
rect 158 137 159 138
rect 139 137 140 138
rect 138 137 139 138
rect 137 137 138 138
rect 136 137 137 138
rect 135 137 136 138
rect 134 137 135 138
rect 133 137 134 138
rect 132 137 133 138
rect 131 137 132 138
rect 130 137 131 138
rect 129 137 130 138
rect 128 137 129 138
rect 127 137 128 138
rect 126 137 127 138
rect 125 137 126 138
rect 124 137 125 138
rect 123 137 124 138
rect 122 137 123 138
rect 121 137 122 138
rect 120 137 121 138
rect 119 137 120 138
rect 118 137 119 138
rect 117 137 118 138
rect 116 137 117 138
rect 115 137 116 138
rect 114 137 115 138
rect 113 137 114 138
rect 112 137 113 138
rect 111 137 112 138
rect 110 137 111 138
rect 109 137 110 138
rect 108 137 109 138
rect 107 137 108 138
rect 106 137 107 138
rect 105 137 106 138
rect 104 137 105 138
rect 103 137 104 138
rect 102 137 103 138
rect 101 137 102 138
rect 100 137 101 138
rect 99 137 100 138
rect 98 137 99 138
rect 97 137 98 138
rect 96 137 97 138
rect 95 137 96 138
rect 94 137 95 138
rect 93 137 94 138
rect 92 137 93 138
rect 91 137 92 138
rect 90 137 91 138
rect 89 137 90 138
rect 88 137 89 138
rect 87 137 88 138
rect 86 137 87 138
rect 85 137 86 138
rect 84 137 85 138
rect 83 137 84 138
rect 82 137 83 138
rect 81 137 82 138
rect 80 137 81 138
rect 79 137 80 138
rect 78 137 79 138
rect 77 137 78 138
rect 76 137 77 138
rect 75 137 76 138
rect 74 137 75 138
rect 73 137 74 138
rect 72 137 73 138
rect 71 137 72 138
rect 70 137 71 138
rect 69 137 70 138
rect 68 137 69 138
rect 67 137 68 138
rect 66 137 67 138
rect 65 137 66 138
rect 64 137 65 138
rect 63 137 64 138
rect 62 137 63 138
rect 61 137 62 138
rect 60 137 61 138
rect 59 137 60 138
rect 58 137 59 138
rect 57 137 58 138
rect 56 137 57 138
rect 55 137 56 138
rect 54 137 55 138
rect 53 137 54 138
rect 52 137 53 138
rect 51 137 52 138
rect 50 137 51 138
rect 49 137 50 138
rect 48 137 49 138
rect 47 137 48 138
rect 46 137 47 138
rect 45 137 46 138
rect 44 137 45 138
rect 43 137 44 138
rect 42 137 43 138
rect 41 137 42 138
rect 40 137 41 138
rect 39 137 40 138
rect 38 137 39 138
rect 37 137 38 138
rect 36 137 37 138
rect 35 137 36 138
rect 433 138 434 139
rect 432 138 433 139
rect 431 138 432 139
rect 430 138 431 139
rect 429 138 430 139
rect 428 138 429 139
rect 427 138 428 139
rect 426 138 427 139
rect 425 138 426 139
rect 424 138 425 139
rect 423 138 424 139
rect 422 138 423 139
rect 421 138 422 139
rect 420 138 421 139
rect 419 138 420 139
rect 418 138 419 139
rect 417 138 418 139
rect 416 138 417 139
rect 415 138 416 139
rect 414 138 415 139
rect 413 138 414 139
rect 412 138 413 139
rect 411 138 412 139
rect 410 138 411 139
rect 409 138 410 139
rect 408 138 409 139
rect 407 138 408 139
rect 406 138 407 139
rect 405 138 406 139
rect 404 138 405 139
rect 403 138 404 139
rect 402 138 403 139
rect 401 138 402 139
rect 400 138 401 139
rect 399 138 400 139
rect 398 138 399 139
rect 397 138 398 139
rect 396 138 397 139
rect 395 138 396 139
rect 394 138 395 139
rect 393 138 394 139
rect 311 138 312 139
rect 310 138 311 139
rect 309 138 310 139
rect 308 138 309 139
rect 307 138 308 139
rect 306 138 307 139
rect 305 138 306 139
rect 304 138 305 139
rect 303 138 304 139
rect 302 138 303 139
rect 301 138 302 139
rect 300 138 301 139
rect 299 138 300 139
rect 298 138 299 139
rect 297 138 298 139
rect 296 138 297 139
rect 295 138 296 139
rect 294 138 295 139
rect 293 138 294 139
rect 292 138 293 139
rect 291 138 292 139
rect 290 138 291 139
rect 289 138 290 139
rect 288 138 289 139
rect 287 138 288 139
rect 286 138 287 139
rect 285 138 286 139
rect 284 138 285 139
rect 283 138 284 139
rect 282 138 283 139
rect 281 138 282 139
rect 280 138 281 139
rect 279 138 280 139
rect 278 138 279 139
rect 277 138 278 139
rect 276 138 277 139
rect 275 138 276 139
rect 274 138 275 139
rect 273 138 274 139
rect 272 138 273 139
rect 271 138 272 139
rect 270 138 271 139
rect 269 138 270 139
rect 268 138 269 139
rect 267 138 268 139
rect 266 138 267 139
rect 265 138 266 139
rect 264 138 265 139
rect 263 138 264 139
rect 262 138 263 139
rect 261 138 262 139
rect 260 138 261 139
rect 259 138 260 139
rect 258 138 259 139
rect 257 138 258 139
rect 256 138 257 139
rect 255 138 256 139
rect 254 138 255 139
rect 253 138 254 139
rect 252 138 253 139
rect 251 138 252 139
rect 250 138 251 139
rect 249 138 250 139
rect 248 138 249 139
rect 247 138 248 139
rect 246 138 247 139
rect 245 138 246 139
rect 221 138 222 139
rect 220 138 221 139
rect 219 138 220 139
rect 218 138 219 139
rect 217 138 218 139
rect 216 138 217 139
rect 215 138 216 139
rect 214 138 215 139
rect 213 138 214 139
rect 212 138 213 139
rect 211 138 212 139
rect 210 138 211 139
rect 209 138 210 139
rect 208 138 209 139
rect 207 138 208 139
rect 206 138 207 139
rect 205 138 206 139
rect 204 138 205 139
rect 203 138 204 139
rect 202 138 203 139
rect 201 138 202 139
rect 200 138 201 139
rect 199 138 200 139
rect 198 138 199 139
rect 197 138 198 139
rect 196 138 197 139
rect 195 138 196 139
rect 194 138 195 139
rect 193 138 194 139
rect 192 138 193 139
rect 191 138 192 139
rect 190 138 191 139
rect 189 138 190 139
rect 188 138 189 139
rect 187 138 188 139
rect 186 138 187 139
rect 185 138 186 139
rect 184 138 185 139
rect 183 138 184 139
rect 182 138 183 139
rect 181 138 182 139
rect 180 138 181 139
rect 179 138 180 139
rect 178 138 179 139
rect 177 138 178 139
rect 176 138 177 139
rect 175 138 176 139
rect 174 138 175 139
rect 173 138 174 139
rect 172 138 173 139
rect 171 138 172 139
rect 170 138 171 139
rect 169 138 170 139
rect 168 138 169 139
rect 167 138 168 139
rect 166 138 167 139
rect 165 138 166 139
rect 164 138 165 139
rect 163 138 164 139
rect 162 138 163 139
rect 161 138 162 139
rect 160 138 161 139
rect 159 138 160 139
rect 158 138 159 139
rect 138 138 139 139
rect 137 138 138 139
rect 136 138 137 139
rect 135 138 136 139
rect 134 138 135 139
rect 133 138 134 139
rect 132 138 133 139
rect 131 138 132 139
rect 130 138 131 139
rect 129 138 130 139
rect 128 138 129 139
rect 127 138 128 139
rect 126 138 127 139
rect 125 138 126 139
rect 124 138 125 139
rect 123 138 124 139
rect 122 138 123 139
rect 121 138 122 139
rect 120 138 121 139
rect 119 138 120 139
rect 118 138 119 139
rect 117 138 118 139
rect 116 138 117 139
rect 115 138 116 139
rect 114 138 115 139
rect 113 138 114 139
rect 112 138 113 139
rect 111 138 112 139
rect 110 138 111 139
rect 109 138 110 139
rect 108 138 109 139
rect 107 138 108 139
rect 106 138 107 139
rect 105 138 106 139
rect 104 138 105 139
rect 103 138 104 139
rect 102 138 103 139
rect 101 138 102 139
rect 100 138 101 139
rect 99 138 100 139
rect 98 138 99 139
rect 97 138 98 139
rect 96 138 97 139
rect 95 138 96 139
rect 94 138 95 139
rect 93 138 94 139
rect 92 138 93 139
rect 91 138 92 139
rect 90 138 91 139
rect 89 138 90 139
rect 88 138 89 139
rect 87 138 88 139
rect 86 138 87 139
rect 85 138 86 139
rect 84 138 85 139
rect 83 138 84 139
rect 82 138 83 139
rect 81 138 82 139
rect 80 138 81 139
rect 79 138 80 139
rect 78 138 79 139
rect 77 138 78 139
rect 76 138 77 139
rect 75 138 76 139
rect 74 138 75 139
rect 73 138 74 139
rect 72 138 73 139
rect 71 138 72 139
rect 70 138 71 139
rect 69 138 70 139
rect 68 138 69 139
rect 67 138 68 139
rect 66 138 67 139
rect 65 138 66 139
rect 64 138 65 139
rect 63 138 64 139
rect 62 138 63 139
rect 61 138 62 139
rect 60 138 61 139
rect 59 138 60 139
rect 58 138 59 139
rect 57 138 58 139
rect 56 138 57 139
rect 55 138 56 139
rect 54 138 55 139
rect 53 138 54 139
rect 52 138 53 139
rect 51 138 52 139
rect 50 138 51 139
rect 49 138 50 139
rect 48 138 49 139
rect 47 138 48 139
rect 46 138 47 139
rect 45 138 46 139
rect 44 138 45 139
rect 43 138 44 139
rect 42 138 43 139
rect 41 138 42 139
rect 40 138 41 139
rect 39 138 40 139
rect 38 138 39 139
rect 37 138 38 139
rect 36 138 37 139
rect 431 139 432 140
rect 430 139 431 140
rect 429 139 430 140
rect 428 139 429 140
rect 427 139 428 140
rect 426 139 427 140
rect 425 139 426 140
rect 424 139 425 140
rect 423 139 424 140
rect 422 139 423 140
rect 421 139 422 140
rect 420 139 421 140
rect 419 139 420 140
rect 418 139 419 140
rect 417 139 418 140
rect 416 139 417 140
rect 415 139 416 140
rect 414 139 415 140
rect 413 139 414 140
rect 412 139 413 140
rect 411 139 412 140
rect 410 139 411 140
rect 409 139 410 140
rect 408 139 409 140
rect 407 139 408 140
rect 406 139 407 140
rect 405 139 406 140
rect 404 139 405 140
rect 403 139 404 140
rect 402 139 403 140
rect 401 139 402 140
rect 400 139 401 140
rect 399 139 400 140
rect 398 139 399 140
rect 397 139 398 140
rect 396 139 397 140
rect 395 139 396 140
rect 394 139 395 140
rect 393 139 394 140
rect 311 139 312 140
rect 310 139 311 140
rect 309 139 310 140
rect 308 139 309 140
rect 307 139 308 140
rect 306 139 307 140
rect 305 139 306 140
rect 304 139 305 140
rect 303 139 304 140
rect 302 139 303 140
rect 301 139 302 140
rect 300 139 301 140
rect 299 139 300 140
rect 298 139 299 140
rect 297 139 298 140
rect 296 139 297 140
rect 295 139 296 140
rect 294 139 295 140
rect 293 139 294 140
rect 292 139 293 140
rect 291 139 292 140
rect 290 139 291 140
rect 289 139 290 140
rect 288 139 289 140
rect 287 139 288 140
rect 286 139 287 140
rect 285 139 286 140
rect 284 139 285 140
rect 283 139 284 140
rect 282 139 283 140
rect 281 139 282 140
rect 280 139 281 140
rect 279 139 280 140
rect 278 139 279 140
rect 277 139 278 140
rect 276 139 277 140
rect 275 139 276 140
rect 274 139 275 140
rect 273 139 274 140
rect 272 139 273 140
rect 271 139 272 140
rect 270 139 271 140
rect 269 139 270 140
rect 268 139 269 140
rect 267 139 268 140
rect 266 139 267 140
rect 265 139 266 140
rect 264 139 265 140
rect 263 139 264 140
rect 262 139 263 140
rect 261 139 262 140
rect 260 139 261 140
rect 259 139 260 140
rect 258 139 259 140
rect 257 139 258 140
rect 256 139 257 140
rect 255 139 256 140
rect 254 139 255 140
rect 253 139 254 140
rect 252 139 253 140
rect 251 139 252 140
rect 250 139 251 140
rect 249 139 250 140
rect 248 139 249 140
rect 247 139 248 140
rect 246 139 247 140
rect 245 139 246 140
rect 244 139 245 140
rect 220 139 221 140
rect 219 139 220 140
rect 218 139 219 140
rect 217 139 218 140
rect 216 139 217 140
rect 215 139 216 140
rect 214 139 215 140
rect 213 139 214 140
rect 212 139 213 140
rect 211 139 212 140
rect 210 139 211 140
rect 209 139 210 140
rect 208 139 209 140
rect 207 139 208 140
rect 206 139 207 140
rect 205 139 206 140
rect 204 139 205 140
rect 203 139 204 140
rect 202 139 203 140
rect 201 139 202 140
rect 200 139 201 140
rect 199 139 200 140
rect 198 139 199 140
rect 197 139 198 140
rect 196 139 197 140
rect 195 139 196 140
rect 194 139 195 140
rect 193 139 194 140
rect 192 139 193 140
rect 191 139 192 140
rect 190 139 191 140
rect 189 139 190 140
rect 188 139 189 140
rect 187 139 188 140
rect 186 139 187 140
rect 185 139 186 140
rect 184 139 185 140
rect 183 139 184 140
rect 182 139 183 140
rect 181 139 182 140
rect 180 139 181 140
rect 179 139 180 140
rect 178 139 179 140
rect 177 139 178 140
rect 176 139 177 140
rect 175 139 176 140
rect 174 139 175 140
rect 173 139 174 140
rect 172 139 173 140
rect 171 139 172 140
rect 170 139 171 140
rect 169 139 170 140
rect 168 139 169 140
rect 167 139 168 140
rect 166 139 167 140
rect 165 139 166 140
rect 164 139 165 140
rect 163 139 164 140
rect 162 139 163 140
rect 161 139 162 140
rect 160 139 161 140
rect 159 139 160 140
rect 158 139 159 140
rect 157 139 158 140
rect 137 139 138 140
rect 136 139 137 140
rect 135 139 136 140
rect 134 139 135 140
rect 133 139 134 140
rect 132 139 133 140
rect 131 139 132 140
rect 130 139 131 140
rect 129 139 130 140
rect 128 139 129 140
rect 127 139 128 140
rect 126 139 127 140
rect 125 139 126 140
rect 124 139 125 140
rect 123 139 124 140
rect 122 139 123 140
rect 121 139 122 140
rect 120 139 121 140
rect 119 139 120 140
rect 118 139 119 140
rect 117 139 118 140
rect 116 139 117 140
rect 115 139 116 140
rect 114 139 115 140
rect 113 139 114 140
rect 112 139 113 140
rect 111 139 112 140
rect 110 139 111 140
rect 109 139 110 140
rect 108 139 109 140
rect 107 139 108 140
rect 106 139 107 140
rect 105 139 106 140
rect 104 139 105 140
rect 103 139 104 140
rect 102 139 103 140
rect 101 139 102 140
rect 100 139 101 140
rect 99 139 100 140
rect 98 139 99 140
rect 97 139 98 140
rect 96 139 97 140
rect 95 139 96 140
rect 94 139 95 140
rect 93 139 94 140
rect 92 139 93 140
rect 91 139 92 140
rect 90 139 91 140
rect 89 139 90 140
rect 88 139 89 140
rect 87 139 88 140
rect 86 139 87 140
rect 85 139 86 140
rect 84 139 85 140
rect 83 139 84 140
rect 82 139 83 140
rect 81 139 82 140
rect 80 139 81 140
rect 79 139 80 140
rect 78 139 79 140
rect 77 139 78 140
rect 76 139 77 140
rect 75 139 76 140
rect 74 139 75 140
rect 73 139 74 140
rect 72 139 73 140
rect 71 139 72 140
rect 70 139 71 140
rect 69 139 70 140
rect 68 139 69 140
rect 67 139 68 140
rect 66 139 67 140
rect 65 139 66 140
rect 64 139 65 140
rect 63 139 64 140
rect 62 139 63 140
rect 61 139 62 140
rect 60 139 61 140
rect 59 139 60 140
rect 58 139 59 140
rect 57 139 58 140
rect 56 139 57 140
rect 55 139 56 140
rect 54 139 55 140
rect 53 139 54 140
rect 52 139 53 140
rect 51 139 52 140
rect 50 139 51 140
rect 49 139 50 140
rect 48 139 49 140
rect 47 139 48 140
rect 46 139 47 140
rect 45 139 46 140
rect 44 139 45 140
rect 43 139 44 140
rect 42 139 43 140
rect 41 139 42 140
rect 40 139 41 140
rect 39 139 40 140
rect 38 139 39 140
rect 37 139 38 140
rect 478 140 479 141
rect 458 140 459 141
rect 429 140 430 141
rect 428 140 429 141
rect 427 140 428 141
rect 426 140 427 141
rect 425 140 426 141
rect 424 140 425 141
rect 423 140 424 141
rect 422 140 423 141
rect 421 140 422 141
rect 420 140 421 141
rect 419 140 420 141
rect 418 140 419 141
rect 417 140 418 141
rect 416 140 417 141
rect 415 140 416 141
rect 414 140 415 141
rect 413 140 414 141
rect 412 140 413 141
rect 411 140 412 141
rect 410 140 411 141
rect 409 140 410 141
rect 408 140 409 141
rect 407 140 408 141
rect 406 140 407 141
rect 405 140 406 141
rect 404 140 405 141
rect 403 140 404 141
rect 402 140 403 141
rect 401 140 402 141
rect 400 140 401 141
rect 399 140 400 141
rect 398 140 399 141
rect 397 140 398 141
rect 396 140 397 141
rect 395 140 396 141
rect 394 140 395 141
rect 393 140 394 141
rect 312 140 313 141
rect 311 140 312 141
rect 310 140 311 141
rect 309 140 310 141
rect 308 140 309 141
rect 307 140 308 141
rect 306 140 307 141
rect 305 140 306 141
rect 304 140 305 141
rect 303 140 304 141
rect 302 140 303 141
rect 301 140 302 141
rect 300 140 301 141
rect 299 140 300 141
rect 298 140 299 141
rect 297 140 298 141
rect 296 140 297 141
rect 295 140 296 141
rect 294 140 295 141
rect 293 140 294 141
rect 292 140 293 141
rect 291 140 292 141
rect 290 140 291 141
rect 289 140 290 141
rect 288 140 289 141
rect 287 140 288 141
rect 286 140 287 141
rect 285 140 286 141
rect 284 140 285 141
rect 283 140 284 141
rect 282 140 283 141
rect 281 140 282 141
rect 280 140 281 141
rect 279 140 280 141
rect 278 140 279 141
rect 277 140 278 141
rect 276 140 277 141
rect 275 140 276 141
rect 274 140 275 141
rect 273 140 274 141
rect 272 140 273 141
rect 271 140 272 141
rect 270 140 271 141
rect 269 140 270 141
rect 268 140 269 141
rect 267 140 268 141
rect 266 140 267 141
rect 265 140 266 141
rect 264 140 265 141
rect 263 140 264 141
rect 262 140 263 141
rect 261 140 262 141
rect 260 140 261 141
rect 259 140 260 141
rect 258 140 259 141
rect 257 140 258 141
rect 256 140 257 141
rect 255 140 256 141
rect 254 140 255 141
rect 253 140 254 141
rect 252 140 253 141
rect 251 140 252 141
rect 250 140 251 141
rect 249 140 250 141
rect 248 140 249 141
rect 247 140 248 141
rect 246 140 247 141
rect 245 140 246 141
rect 244 140 245 141
rect 243 140 244 141
rect 220 140 221 141
rect 219 140 220 141
rect 218 140 219 141
rect 217 140 218 141
rect 216 140 217 141
rect 215 140 216 141
rect 214 140 215 141
rect 213 140 214 141
rect 212 140 213 141
rect 211 140 212 141
rect 210 140 211 141
rect 209 140 210 141
rect 208 140 209 141
rect 207 140 208 141
rect 206 140 207 141
rect 205 140 206 141
rect 204 140 205 141
rect 203 140 204 141
rect 202 140 203 141
rect 201 140 202 141
rect 200 140 201 141
rect 199 140 200 141
rect 198 140 199 141
rect 197 140 198 141
rect 196 140 197 141
rect 195 140 196 141
rect 194 140 195 141
rect 193 140 194 141
rect 192 140 193 141
rect 191 140 192 141
rect 190 140 191 141
rect 189 140 190 141
rect 188 140 189 141
rect 187 140 188 141
rect 186 140 187 141
rect 185 140 186 141
rect 184 140 185 141
rect 183 140 184 141
rect 182 140 183 141
rect 181 140 182 141
rect 180 140 181 141
rect 179 140 180 141
rect 178 140 179 141
rect 177 140 178 141
rect 176 140 177 141
rect 175 140 176 141
rect 174 140 175 141
rect 173 140 174 141
rect 172 140 173 141
rect 171 140 172 141
rect 170 140 171 141
rect 169 140 170 141
rect 168 140 169 141
rect 167 140 168 141
rect 166 140 167 141
rect 165 140 166 141
rect 164 140 165 141
rect 163 140 164 141
rect 162 140 163 141
rect 161 140 162 141
rect 160 140 161 141
rect 159 140 160 141
rect 158 140 159 141
rect 157 140 158 141
rect 136 140 137 141
rect 135 140 136 141
rect 134 140 135 141
rect 133 140 134 141
rect 132 140 133 141
rect 131 140 132 141
rect 130 140 131 141
rect 129 140 130 141
rect 128 140 129 141
rect 127 140 128 141
rect 126 140 127 141
rect 125 140 126 141
rect 124 140 125 141
rect 123 140 124 141
rect 122 140 123 141
rect 121 140 122 141
rect 120 140 121 141
rect 119 140 120 141
rect 118 140 119 141
rect 117 140 118 141
rect 116 140 117 141
rect 115 140 116 141
rect 114 140 115 141
rect 113 140 114 141
rect 112 140 113 141
rect 111 140 112 141
rect 110 140 111 141
rect 109 140 110 141
rect 108 140 109 141
rect 107 140 108 141
rect 106 140 107 141
rect 105 140 106 141
rect 104 140 105 141
rect 103 140 104 141
rect 102 140 103 141
rect 101 140 102 141
rect 100 140 101 141
rect 99 140 100 141
rect 98 140 99 141
rect 97 140 98 141
rect 96 140 97 141
rect 95 140 96 141
rect 94 140 95 141
rect 93 140 94 141
rect 92 140 93 141
rect 91 140 92 141
rect 90 140 91 141
rect 89 140 90 141
rect 88 140 89 141
rect 87 140 88 141
rect 86 140 87 141
rect 85 140 86 141
rect 84 140 85 141
rect 83 140 84 141
rect 82 140 83 141
rect 81 140 82 141
rect 80 140 81 141
rect 79 140 80 141
rect 78 140 79 141
rect 77 140 78 141
rect 76 140 77 141
rect 75 140 76 141
rect 74 140 75 141
rect 73 140 74 141
rect 72 140 73 141
rect 71 140 72 141
rect 70 140 71 141
rect 69 140 70 141
rect 68 140 69 141
rect 67 140 68 141
rect 66 140 67 141
rect 65 140 66 141
rect 64 140 65 141
rect 63 140 64 141
rect 62 140 63 141
rect 61 140 62 141
rect 60 140 61 141
rect 59 140 60 141
rect 58 140 59 141
rect 57 140 58 141
rect 56 140 57 141
rect 55 140 56 141
rect 54 140 55 141
rect 53 140 54 141
rect 52 140 53 141
rect 51 140 52 141
rect 50 140 51 141
rect 49 140 50 141
rect 48 140 49 141
rect 47 140 48 141
rect 46 140 47 141
rect 45 140 46 141
rect 44 140 45 141
rect 43 140 44 141
rect 42 140 43 141
rect 41 140 42 141
rect 40 140 41 141
rect 39 140 40 141
rect 38 140 39 141
rect 37 140 38 141
rect 22 140 23 141
rect 21 140 22 141
rect 20 140 21 141
rect 19 140 20 141
rect 18 140 19 141
rect 478 141 479 142
rect 458 141 459 142
rect 425 141 426 142
rect 424 141 425 142
rect 423 141 424 142
rect 422 141 423 142
rect 421 141 422 142
rect 420 141 421 142
rect 419 141 420 142
rect 418 141 419 142
rect 417 141 418 142
rect 416 141 417 142
rect 415 141 416 142
rect 414 141 415 142
rect 413 141 414 142
rect 412 141 413 142
rect 411 141 412 142
rect 410 141 411 142
rect 409 141 410 142
rect 408 141 409 142
rect 407 141 408 142
rect 406 141 407 142
rect 405 141 406 142
rect 404 141 405 142
rect 403 141 404 142
rect 402 141 403 142
rect 401 141 402 142
rect 400 141 401 142
rect 399 141 400 142
rect 398 141 399 142
rect 397 141 398 142
rect 396 141 397 142
rect 395 141 396 142
rect 394 141 395 142
rect 393 141 394 142
rect 313 141 314 142
rect 312 141 313 142
rect 311 141 312 142
rect 310 141 311 142
rect 309 141 310 142
rect 308 141 309 142
rect 307 141 308 142
rect 306 141 307 142
rect 305 141 306 142
rect 304 141 305 142
rect 303 141 304 142
rect 302 141 303 142
rect 301 141 302 142
rect 300 141 301 142
rect 299 141 300 142
rect 298 141 299 142
rect 297 141 298 142
rect 296 141 297 142
rect 295 141 296 142
rect 294 141 295 142
rect 293 141 294 142
rect 292 141 293 142
rect 291 141 292 142
rect 290 141 291 142
rect 289 141 290 142
rect 288 141 289 142
rect 287 141 288 142
rect 286 141 287 142
rect 285 141 286 142
rect 284 141 285 142
rect 283 141 284 142
rect 282 141 283 142
rect 281 141 282 142
rect 280 141 281 142
rect 279 141 280 142
rect 278 141 279 142
rect 277 141 278 142
rect 276 141 277 142
rect 275 141 276 142
rect 274 141 275 142
rect 273 141 274 142
rect 272 141 273 142
rect 271 141 272 142
rect 270 141 271 142
rect 269 141 270 142
rect 268 141 269 142
rect 267 141 268 142
rect 266 141 267 142
rect 265 141 266 142
rect 264 141 265 142
rect 263 141 264 142
rect 262 141 263 142
rect 261 141 262 142
rect 260 141 261 142
rect 259 141 260 142
rect 258 141 259 142
rect 257 141 258 142
rect 256 141 257 142
rect 255 141 256 142
rect 254 141 255 142
rect 253 141 254 142
rect 252 141 253 142
rect 251 141 252 142
rect 250 141 251 142
rect 249 141 250 142
rect 248 141 249 142
rect 247 141 248 142
rect 246 141 247 142
rect 245 141 246 142
rect 244 141 245 142
rect 243 141 244 142
rect 242 141 243 142
rect 219 141 220 142
rect 218 141 219 142
rect 217 141 218 142
rect 216 141 217 142
rect 215 141 216 142
rect 214 141 215 142
rect 213 141 214 142
rect 212 141 213 142
rect 211 141 212 142
rect 210 141 211 142
rect 209 141 210 142
rect 208 141 209 142
rect 207 141 208 142
rect 206 141 207 142
rect 205 141 206 142
rect 204 141 205 142
rect 203 141 204 142
rect 202 141 203 142
rect 201 141 202 142
rect 200 141 201 142
rect 199 141 200 142
rect 198 141 199 142
rect 197 141 198 142
rect 196 141 197 142
rect 195 141 196 142
rect 194 141 195 142
rect 193 141 194 142
rect 192 141 193 142
rect 191 141 192 142
rect 190 141 191 142
rect 189 141 190 142
rect 188 141 189 142
rect 187 141 188 142
rect 186 141 187 142
rect 185 141 186 142
rect 184 141 185 142
rect 183 141 184 142
rect 182 141 183 142
rect 181 141 182 142
rect 180 141 181 142
rect 179 141 180 142
rect 178 141 179 142
rect 177 141 178 142
rect 176 141 177 142
rect 175 141 176 142
rect 174 141 175 142
rect 173 141 174 142
rect 172 141 173 142
rect 171 141 172 142
rect 170 141 171 142
rect 169 141 170 142
rect 168 141 169 142
rect 167 141 168 142
rect 166 141 167 142
rect 165 141 166 142
rect 164 141 165 142
rect 163 141 164 142
rect 162 141 163 142
rect 161 141 162 142
rect 160 141 161 142
rect 159 141 160 142
rect 158 141 159 142
rect 157 141 158 142
rect 156 141 157 142
rect 135 141 136 142
rect 134 141 135 142
rect 133 141 134 142
rect 132 141 133 142
rect 131 141 132 142
rect 130 141 131 142
rect 129 141 130 142
rect 128 141 129 142
rect 127 141 128 142
rect 126 141 127 142
rect 125 141 126 142
rect 124 141 125 142
rect 123 141 124 142
rect 122 141 123 142
rect 121 141 122 142
rect 120 141 121 142
rect 119 141 120 142
rect 118 141 119 142
rect 117 141 118 142
rect 116 141 117 142
rect 115 141 116 142
rect 114 141 115 142
rect 113 141 114 142
rect 112 141 113 142
rect 111 141 112 142
rect 110 141 111 142
rect 109 141 110 142
rect 108 141 109 142
rect 107 141 108 142
rect 106 141 107 142
rect 105 141 106 142
rect 104 141 105 142
rect 103 141 104 142
rect 102 141 103 142
rect 101 141 102 142
rect 100 141 101 142
rect 99 141 100 142
rect 98 141 99 142
rect 97 141 98 142
rect 96 141 97 142
rect 95 141 96 142
rect 94 141 95 142
rect 93 141 94 142
rect 92 141 93 142
rect 91 141 92 142
rect 90 141 91 142
rect 89 141 90 142
rect 88 141 89 142
rect 87 141 88 142
rect 86 141 87 142
rect 85 141 86 142
rect 84 141 85 142
rect 83 141 84 142
rect 82 141 83 142
rect 81 141 82 142
rect 80 141 81 142
rect 79 141 80 142
rect 78 141 79 142
rect 77 141 78 142
rect 76 141 77 142
rect 75 141 76 142
rect 74 141 75 142
rect 73 141 74 142
rect 72 141 73 142
rect 71 141 72 142
rect 70 141 71 142
rect 69 141 70 142
rect 68 141 69 142
rect 67 141 68 142
rect 66 141 67 142
rect 65 141 66 142
rect 64 141 65 142
rect 63 141 64 142
rect 62 141 63 142
rect 61 141 62 142
rect 60 141 61 142
rect 59 141 60 142
rect 58 141 59 142
rect 57 141 58 142
rect 56 141 57 142
rect 55 141 56 142
rect 54 141 55 142
rect 53 141 54 142
rect 52 141 53 142
rect 51 141 52 142
rect 50 141 51 142
rect 49 141 50 142
rect 48 141 49 142
rect 47 141 48 142
rect 46 141 47 142
rect 45 141 46 142
rect 44 141 45 142
rect 43 141 44 142
rect 42 141 43 142
rect 41 141 42 142
rect 40 141 41 142
rect 39 141 40 142
rect 38 141 39 142
rect 24 141 25 142
rect 23 141 24 142
rect 22 141 23 142
rect 21 141 22 142
rect 20 141 21 142
rect 19 141 20 142
rect 18 141 19 142
rect 17 141 18 142
rect 16 141 17 142
rect 15 141 16 142
rect 478 142 479 143
rect 477 142 478 143
rect 459 142 460 143
rect 458 142 459 143
rect 402 142 403 143
rect 401 142 402 143
rect 400 142 401 143
rect 399 142 400 143
rect 398 142 399 143
rect 397 142 398 143
rect 396 142 397 143
rect 395 142 396 143
rect 394 142 395 143
rect 393 142 394 143
rect 314 142 315 143
rect 313 142 314 143
rect 312 142 313 143
rect 311 142 312 143
rect 310 142 311 143
rect 309 142 310 143
rect 308 142 309 143
rect 307 142 308 143
rect 306 142 307 143
rect 305 142 306 143
rect 304 142 305 143
rect 303 142 304 143
rect 302 142 303 143
rect 301 142 302 143
rect 300 142 301 143
rect 299 142 300 143
rect 298 142 299 143
rect 297 142 298 143
rect 296 142 297 143
rect 295 142 296 143
rect 294 142 295 143
rect 293 142 294 143
rect 292 142 293 143
rect 291 142 292 143
rect 290 142 291 143
rect 289 142 290 143
rect 288 142 289 143
rect 287 142 288 143
rect 286 142 287 143
rect 285 142 286 143
rect 284 142 285 143
rect 283 142 284 143
rect 282 142 283 143
rect 281 142 282 143
rect 280 142 281 143
rect 279 142 280 143
rect 278 142 279 143
rect 277 142 278 143
rect 276 142 277 143
rect 275 142 276 143
rect 274 142 275 143
rect 273 142 274 143
rect 272 142 273 143
rect 271 142 272 143
rect 270 142 271 143
rect 269 142 270 143
rect 268 142 269 143
rect 267 142 268 143
rect 266 142 267 143
rect 265 142 266 143
rect 264 142 265 143
rect 263 142 264 143
rect 262 142 263 143
rect 261 142 262 143
rect 260 142 261 143
rect 259 142 260 143
rect 258 142 259 143
rect 257 142 258 143
rect 256 142 257 143
rect 255 142 256 143
rect 254 142 255 143
rect 253 142 254 143
rect 252 142 253 143
rect 251 142 252 143
rect 250 142 251 143
rect 249 142 250 143
rect 248 142 249 143
rect 247 142 248 143
rect 246 142 247 143
rect 245 142 246 143
rect 244 142 245 143
rect 243 142 244 143
rect 242 142 243 143
rect 241 142 242 143
rect 219 142 220 143
rect 218 142 219 143
rect 217 142 218 143
rect 216 142 217 143
rect 215 142 216 143
rect 214 142 215 143
rect 213 142 214 143
rect 212 142 213 143
rect 211 142 212 143
rect 210 142 211 143
rect 209 142 210 143
rect 208 142 209 143
rect 207 142 208 143
rect 206 142 207 143
rect 205 142 206 143
rect 204 142 205 143
rect 203 142 204 143
rect 202 142 203 143
rect 201 142 202 143
rect 200 142 201 143
rect 199 142 200 143
rect 198 142 199 143
rect 197 142 198 143
rect 196 142 197 143
rect 195 142 196 143
rect 194 142 195 143
rect 193 142 194 143
rect 192 142 193 143
rect 191 142 192 143
rect 190 142 191 143
rect 189 142 190 143
rect 188 142 189 143
rect 187 142 188 143
rect 186 142 187 143
rect 185 142 186 143
rect 184 142 185 143
rect 183 142 184 143
rect 182 142 183 143
rect 181 142 182 143
rect 180 142 181 143
rect 179 142 180 143
rect 178 142 179 143
rect 177 142 178 143
rect 176 142 177 143
rect 175 142 176 143
rect 174 142 175 143
rect 173 142 174 143
rect 172 142 173 143
rect 171 142 172 143
rect 170 142 171 143
rect 169 142 170 143
rect 168 142 169 143
rect 167 142 168 143
rect 166 142 167 143
rect 165 142 166 143
rect 164 142 165 143
rect 163 142 164 143
rect 162 142 163 143
rect 161 142 162 143
rect 160 142 161 143
rect 159 142 160 143
rect 158 142 159 143
rect 157 142 158 143
rect 156 142 157 143
rect 134 142 135 143
rect 133 142 134 143
rect 132 142 133 143
rect 131 142 132 143
rect 130 142 131 143
rect 129 142 130 143
rect 128 142 129 143
rect 127 142 128 143
rect 126 142 127 143
rect 125 142 126 143
rect 124 142 125 143
rect 123 142 124 143
rect 122 142 123 143
rect 121 142 122 143
rect 120 142 121 143
rect 119 142 120 143
rect 118 142 119 143
rect 117 142 118 143
rect 116 142 117 143
rect 115 142 116 143
rect 114 142 115 143
rect 113 142 114 143
rect 112 142 113 143
rect 111 142 112 143
rect 110 142 111 143
rect 109 142 110 143
rect 108 142 109 143
rect 107 142 108 143
rect 106 142 107 143
rect 105 142 106 143
rect 104 142 105 143
rect 103 142 104 143
rect 102 142 103 143
rect 101 142 102 143
rect 100 142 101 143
rect 99 142 100 143
rect 98 142 99 143
rect 97 142 98 143
rect 96 142 97 143
rect 95 142 96 143
rect 94 142 95 143
rect 93 142 94 143
rect 92 142 93 143
rect 91 142 92 143
rect 90 142 91 143
rect 89 142 90 143
rect 88 142 89 143
rect 87 142 88 143
rect 86 142 87 143
rect 85 142 86 143
rect 84 142 85 143
rect 83 142 84 143
rect 82 142 83 143
rect 81 142 82 143
rect 80 142 81 143
rect 79 142 80 143
rect 78 142 79 143
rect 77 142 78 143
rect 76 142 77 143
rect 75 142 76 143
rect 74 142 75 143
rect 73 142 74 143
rect 72 142 73 143
rect 71 142 72 143
rect 70 142 71 143
rect 69 142 70 143
rect 68 142 69 143
rect 67 142 68 143
rect 66 142 67 143
rect 65 142 66 143
rect 64 142 65 143
rect 63 142 64 143
rect 62 142 63 143
rect 61 142 62 143
rect 60 142 61 143
rect 59 142 60 143
rect 58 142 59 143
rect 57 142 58 143
rect 56 142 57 143
rect 55 142 56 143
rect 54 142 55 143
rect 53 142 54 143
rect 52 142 53 143
rect 51 142 52 143
rect 50 142 51 143
rect 49 142 50 143
rect 48 142 49 143
rect 47 142 48 143
rect 46 142 47 143
rect 45 142 46 143
rect 44 142 45 143
rect 43 142 44 143
rect 42 142 43 143
rect 41 142 42 143
rect 40 142 41 143
rect 39 142 40 143
rect 38 142 39 143
rect 25 142 26 143
rect 24 142 25 143
rect 23 142 24 143
rect 22 142 23 143
rect 21 142 22 143
rect 20 142 21 143
rect 19 142 20 143
rect 18 142 19 143
rect 17 142 18 143
rect 16 142 17 143
rect 15 142 16 143
rect 14 142 15 143
rect 478 143 479 144
rect 477 143 478 144
rect 476 143 477 144
rect 475 143 476 144
rect 474 143 475 144
rect 473 143 474 144
rect 472 143 473 144
rect 471 143 472 144
rect 470 143 471 144
rect 469 143 470 144
rect 468 143 469 144
rect 467 143 468 144
rect 466 143 467 144
rect 465 143 466 144
rect 464 143 465 144
rect 463 143 464 144
rect 462 143 463 144
rect 461 143 462 144
rect 460 143 461 144
rect 459 143 460 144
rect 458 143 459 144
rect 397 143 398 144
rect 396 143 397 144
rect 395 143 396 144
rect 394 143 395 144
rect 393 143 394 144
rect 314 143 315 144
rect 313 143 314 144
rect 312 143 313 144
rect 311 143 312 144
rect 310 143 311 144
rect 309 143 310 144
rect 308 143 309 144
rect 307 143 308 144
rect 306 143 307 144
rect 305 143 306 144
rect 304 143 305 144
rect 303 143 304 144
rect 302 143 303 144
rect 301 143 302 144
rect 300 143 301 144
rect 299 143 300 144
rect 298 143 299 144
rect 297 143 298 144
rect 296 143 297 144
rect 295 143 296 144
rect 294 143 295 144
rect 293 143 294 144
rect 292 143 293 144
rect 291 143 292 144
rect 290 143 291 144
rect 289 143 290 144
rect 288 143 289 144
rect 287 143 288 144
rect 286 143 287 144
rect 285 143 286 144
rect 284 143 285 144
rect 283 143 284 144
rect 282 143 283 144
rect 281 143 282 144
rect 280 143 281 144
rect 279 143 280 144
rect 278 143 279 144
rect 277 143 278 144
rect 276 143 277 144
rect 275 143 276 144
rect 274 143 275 144
rect 273 143 274 144
rect 272 143 273 144
rect 271 143 272 144
rect 270 143 271 144
rect 269 143 270 144
rect 268 143 269 144
rect 267 143 268 144
rect 266 143 267 144
rect 265 143 266 144
rect 264 143 265 144
rect 263 143 264 144
rect 262 143 263 144
rect 261 143 262 144
rect 260 143 261 144
rect 259 143 260 144
rect 258 143 259 144
rect 257 143 258 144
rect 256 143 257 144
rect 255 143 256 144
rect 254 143 255 144
rect 253 143 254 144
rect 252 143 253 144
rect 251 143 252 144
rect 250 143 251 144
rect 249 143 250 144
rect 248 143 249 144
rect 247 143 248 144
rect 246 143 247 144
rect 245 143 246 144
rect 244 143 245 144
rect 243 143 244 144
rect 242 143 243 144
rect 241 143 242 144
rect 219 143 220 144
rect 218 143 219 144
rect 217 143 218 144
rect 216 143 217 144
rect 215 143 216 144
rect 214 143 215 144
rect 213 143 214 144
rect 212 143 213 144
rect 211 143 212 144
rect 210 143 211 144
rect 209 143 210 144
rect 208 143 209 144
rect 207 143 208 144
rect 206 143 207 144
rect 205 143 206 144
rect 204 143 205 144
rect 203 143 204 144
rect 202 143 203 144
rect 201 143 202 144
rect 200 143 201 144
rect 199 143 200 144
rect 198 143 199 144
rect 197 143 198 144
rect 196 143 197 144
rect 195 143 196 144
rect 194 143 195 144
rect 193 143 194 144
rect 192 143 193 144
rect 191 143 192 144
rect 190 143 191 144
rect 189 143 190 144
rect 188 143 189 144
rect 187 143 188 144
rect 186 143 187 144
rect 185 143 186 144
rect 184 143 185 144
rect 183 143 184 144
rect 182 143 183 144
rect 181 143 182 144
rect 180 143 181 144
rect 179 143 180 144
rect 178 143 179 144
rect 177 143 178 144
rect 176 143 177 144
rect 175 143 176 144
rect 174 143 175 144
rect 173 143 174 144
rect 172 143 173 144
rect 171 143 172 144
rect 170 143 171 144
rect 169 143 170 144
rect 168 143 169 144
rect 167 143 168 144
rect 166 143 167 144
rect 165 143 166 144
rect 164 143 165 144
rect 163 143 164 144
rect 162 143 163 144
rect 161 143 162 144
rect 160 143 161 144
rect 159 143 160 144
rect 158 143 159 144
rect 157 143 158 144
rect 156 143 157 144
rect 155 143 156 144
rect 133 143 134 144
rect 132 143 133 144
rect 131 143 132 144
rect 130 143 131 144
rect 129 143 130 144
rect 128 143 129 144
rect 127 143 128 144
rect 126 143 127 144
rect 125 143 126 144
rect 124 143 125 144
rect 123 143 124 144
rect 122 143 123 144
rect 121 143 122 144
rect 120 143 121 144
rect 119 143 120 144
rect 118 143 119 144
rect 117 143 118 144
rect 116 143 117 144
rect 115 143 116 144
rect 114 143 115 144
rect 113 143 114 144
rect 112 143 113 144
rect 111 143 112 144
rect 110 143 111 144
rect 109 143 110 144
rect 108 143 109 144
rect 107 143 108 144
rect 106 143 107 144
rect 105 143 106 144
rect 104 143 105 144
rect 103 143 104 144
rect 102 143 103 144
rect 101 143 102 144
rect 100 143 101 144
rect 99 143 100 144
rect 98 143 99 144
rect 97 143 98 144
rect 96 143 97 144
rect 95 143 96 144
rect 94 143 95 144
rect 93 143 94 144
rect 92 143 93 144
rect 91 143 92 144
rect 90 143 91 144
rect 89 143 90 144
rect 88 143 89 144
rect 87 143 88 144
rect 86 143 87 144
rect 85 143 86 144
rect 84 143 85 144
rect 83 143 84 144
rect 82 143 83 144
rect 81 143 82 144
rect 80 143 81 144
rect 79 143 80 144
rect 78 143 79 144
rect 77 143 78 144
rect 76 143 77 144
rect 75 143 76 144
rect 74 143 75 144
rect 73 143 74 144
rect 72 143 73 144
rect 71 143 72 144
rect 70 143 71 144
rect 69 143 70 144
rect 68 143 69 144
rect 67 143 68 144
rect 66 143 67 144
rect 65 143 66 144
rect 64 143 65 144
rect 63 143 64 144
rect 62 143 63 144
rect 61 143 62 144
rect 60 143 61 144
rect 59 143 60 144
rect 58 143 59 144
rect 57 143 58 144
rect 56 143 57 144
rect 55 143 56 144
rect 54 143 55 144
rect 53 143 54 144
rect 52 143 53 144
rect 51 143 52 144
rect 50 143 51 144
rect 49 143 50 144
rect 48 143 49 144
rect 47 143 48 144
rect 46 143 47 144
rect 45 143 46 144
rect 44 143 45 144
rect 43 143 44 144
rect 42 143 43 144
rect 41 143 42 144
rect 40 143 41 144
rect 39 143 40 144
rect 38 143 39 144
rect 26 143 27 144
rect 25 143 26 144
rect 24 143 25 144
rect 23 143 24 144
rect 22 143 23 144
rect 21 143 22 144
rect 20 143 21 144
rect 19 143 20 144
rect 18 143 19 144
rect 17 143 18 144
rect 16 143 17 144
rect 15 143 16 144
rect 14 143 15 144
rect 13 143 14 144
rect 12 143 13 144
rect 478 144 479 145
rect 477 144 478 145
rect 476 144 477 145
rect 475 144 476 145
rect 474 144 475 145
rect 473 144 474 145
rect 472 144 473 145
rect 471 144 472 145
rect 470 144 471 145
rect 469 144 470 145
rect 468 144 469 145
rect 467 144 468 145
rect 466 144 467 145
rect 465 144 466 145
rect 464 144 465 145
rect 463 144 464 145
rect 462 144 463 145
rect 461 144 462 145
rect 460 144 461 145
rect 459 144 460 145
rect 458 144 459 145
rect 396 144 397 145
rect 395 144 396 145
rect 394 144 395 145
rect 393 144 394 145
rect 315 144 316 145
rect 314 144 315 145
rect 313 144 314 145
rect 312 144 313 145
rect 311 144 312 145
rect 310 144 311 145
rect 309 144 310 145
rect 308 144 309 145
rect 307 144 308 145
rect 306 144 307 145
rect 305 144 306 145
rect 304 144 305 145
rect 303 144 304 145
rect 302 144 303 145
rect 301 144 302 145
rect 300 144 301 145
rect 299 144 300 145
rect 298 144 299 145
rect 297 144 298 145
rect 296 144 297 145
rect 295 144 296 145
rect 294 144 295 145
rect 293 144 294 145
rect 292 144 293 145
rect 291 144 292 145
rect 290 144 291 145
rect 289 144 290 145
rect 288 144 289 145
rect 287 144 288 145
rect 286 144 287 145
rect 285 144 286 145
rect 284 144 285 145
rect 283 144 284 145
rect 282 144 283 145
rect 281 144 282 145
rect 280 144 281 145
rect 279 144 280 145
rect 278 144 279 145
rect 277 144 278 145
rect 276 144 277 145
rect 275 144 276 145
rect 274 144 275 145
rect 273 144 274 145
rect 272 144 273 145
rect 271 144 272 145
rect 270 144 271 145
rect 269 144 270 145
rect 268 144 269 145
rect 267 144 268 145
rect 266 144 267 145
rect 265 144 266 145
rect 264 144 265 145
rect 263 144 264 145
rect 262 144 263 145
rect 261 144 262 145
rect 260 144 261 145
rect 259 144 260 145
rect 258 144 259 145
rect 257 144 258 145
rect 256 144 257 145
rect 255 144 256 145
rect 254 144 255 145
rect 253 144 254 145
rect 252 144 253 145
rect 251 144 252 145
rect 250 144 251 145
rect 249 144 250 145
rect 248 144 249 145
rect 247 144 248 145
rect 246 144 247 145
rect 245 144 246 145
rect 244 144 245 145
rect 243 144 244 145
rect 242 144 243 145
rect 241 144 242 145
rect 240 144 241 145
rect 218 144 219 145
rect 217 144 218 145
rect 216 144 217 145
rect 215 144 216 145
rect 214 144 215 145
rect 213 144 214 145
rect 212 144 213 145
rect 211 144 212 145
rect 210 144 211 145
rect 209 144 210 145
rect 208 144 209 145
rect 207 144 208 145
rect 206 144 207 145
rect 205 144 206 145
rect 204 144 205 145
rect 203 144 204 145
rect 202 144 203 145
rect 201 144 202 145
rect 200 144 201 145
rect 199 144 200 145
rect 198 144 199 145
rect 197 144 198 145
rect 196 144 197 145
rect 195 144 196 145
rect 194 144 195 145
rect 193 144 194 145
rect 192 144 193 145
rect 191 144 192 145
rect 190 144 191 145
rect 189 144 190 145
rect 188 144 189 145
rect 187 144 188 145
rect 186 144 187 145
rect 185 144 186 145
rect 184 144 185 145
rect 183 144 184 145
rect 182 144 183 145
rect 181 144 182 145
rect 180 144 181 145
rect 179 144 180 145
rect 178 144 179 145
rect 177 144 178 145
rect 176 144 177 145
rect 175 144 176 145
rect 174 144 175 145
rect 173 144 174 145
rect 172 144 173 145
rect 171 144 172 145
rect 170 144 171 145
rect 169 144 170 145
rect 168 144 169 145
rect 167 144 168 145
rect 166 144 167 145
rect 165 144 166 145
rect 164 144 165 145
rect 163 144 164 145
rect 162 144 163 145
rect 161 144 162 145
rect 160 144 161 145
rect 159 144 160 145
rect 158 144 159 145
rect 157 144 158 145
rect 156 144 157 145
rect 155 144 156 145
rect 154 144 155 145
rect 132 144 133 145
rect 131 144 132 145
rect 130 144 131 145
rect 129 144 130 145
rect 128 144 129 145
rect 127 144 128 145
rect 126 144 127 145
rect 125 144 126 145
rect 124 144 125 145
rect 123 144 124 145
rect 122 144 123 145
rect 121 144 122 145
rect 120 144 121 145
rect 119 144 120 145
rect 118 144 119 145
rect 117 144 118 145
rect 116 144 117 145
rect 115 144 116 145
rect 114 144 115 145
rect 113 144 114 145
rect 112 144 113 145
rect 111 144 112 145
rect 110 144 111 145
rect 109 144 110 145
rect 108 144 109 145
rect 107 144 108 145
rect 106 144 107 145
rect 105 144 106 145
rect 104 144 105 145
rect 103 144 104 145
rect 102 144 103 145
rect 101 144 102 145
rect 100 144 101 145
rect 99 144 100 145
rect 98 144 99 145
rect 97 144 98 145
rect 96 144 97 145
rect 95 144 96 145
rect 94 144 95 145
rect 93 144 94 145
rect 92 144 93 145
rect 91 144 92 145
rect 90 144 91 145
rect 89 144 90 145
rect 88 144 89 145
rect 87 144 88 145
rect 86 144 87 145
rect 85 144 86 145
rect 84 144 85 145
rect 83 144 84 145
rect 82 144 83 145
rect 81 144 82 145
rect 80 144 81 145
rect 79 144 80 145
rect 78 144 79 145
rect 77 144 78 145
rect 76 144 77 145
rect 75 144 76 145
rect 74 144 75 145
rect 73 144 74 145
rect 72 144 73 145
rect 71 144 72 145
rect 70 144 71 145
rect 69 144 70 145
rect 68 144 69 145
rect 67 144 68 145
rect 66 144 67 145
rect 65 144 66 145
rect 64 144 65 145
rect 63 144 64 145
rect 62 144 63 145
rect 61 144 62 145
rect 60 144 61 145
rect 59 144 60 145
rect 58 144 59 145
rect 57 144 58 145
rect 56 144 57 145
rect 55 144 56 145
rect 54 144 55 145
rect 53 144 54 145
rect 52 144 53 145
rect 51 144 52 145
rect 50 144 51 145
rect 49 144 50 145
rect 48 144 49 145
rect 47 144 48 145
rect 46 144 47 145
rect 45 144 46 145
rect 44 144 45 145
rect 43 144 44 145
rect 42 144 43 145
rect 41 144 42 145
rect 40 144 41 145
rect 39 144 40 145
rect 38 144 39 145
rect 26 144 27 145
rect 25 144 26 145
rect 24 144 25 145
rect 23 144 24 145
rect 22 144 23 145
rect 21 144 22 145
rect 20 144 21 145
rect 19 144 20 145
rect 18 144 19 145
rect 17 144 18 145
rect 16 144 17 145
rect 15 144 16 145
rect 14 144 15 145
rect 13 144 14 145
rect 12 144 13 145
rect 11 144 12 145
rect 478 145 479 146
rect 477 145 478 146
rect 476 145 477 146
rect 475 145 476 146
rect 474 145 475 146
rect 473 145 474 146
rect 472 145 473 146
rect 471 145 472 146
rect 470 145 471 146
rect 469 145 470 146
rect 468 145 469 146
rect 467 145 468 146
rect 466 145 467 146
rect 465 145 466 146
rect 464 145 465 146
rect 463 145 464 146
rect 462 145 463 146
rect 461 145 462 146
rect 460 145 461 146
rect 459 145 460 146
rect 458 145 459 146
rect 395 145 396 146
rect 394 145 395 146
rect 393 145 394 146
rect 316 145 317 146
rect 315 145 316 146
rect 314 145 315 146
rect 313 145 314 146
rect 312 145 313 146
rect 311 145 312 146
rect 310 145 311 146
rect 309 145 310 146
rect 308 145 309 146
rect 307 145 308 146
rect 306 145 307 146
rect 305 145 306 146
rect 304 145 305 146
rect 303 145 304 146
rect 302 145 303 146
rect 301 145 302 146
rect 300 145 301 146
rect 299 145 300 146
rect 298 145 299 146
rect 297 145 298 146
rect 296 145 297 146
rect 295 145 296 146
rect 294 145 295 146
rect 293 145 294 146
rect 292 145 293 146
rect 291 145 292 146
rect 290 145 291 146
rect 289 145 290 146
rect 288 145 289 146
rect 287 145 288 146
rect 286 145 287 146
rect 285 145 286 146
rect 284 145 285 146
rect 283 145 284 146
rect 282 145 283 146
rect 281 145 282 146
rect 280 145 281 146
rect 279 145 280 146
rect 278 145 279 146
rect 277 145 278 146
rect 276 145 277 146
rect 275 145 276 146
rect 274 145 275 146
rect 273 145 274 146
rect 272 145 273 146
rect 271 145 272 146
rect 270 145 271 146
rect 269 145 270 146
rect 268 145 269 146
rect 267 145 268 146
rect 266 145 267 146
rect 265 145 266 146
rect 264 145 265 146
rect 263 145 264 146
rect 262 145 263 146
rect 261 145 262 146
rect 260 145 261 146
rect 259 145 260 146
rect 258 145 259 146
rect 257 145 258 146
rect 256 145 257 146
rect 255 145 256 146
rect 254 145 255 146
rect 253 145 254 146
rect 252 145 253 146
rect 251 145 252 146
rect 250 145 251 146
rect 249 145 250 146
rect 248 145 249 146
rect 247 145 248 146
rect 246 145 247 146
rect 245 145 246 146
rect 244 145 245 146
rect 243 145 244 146
rect 242 145 243 146
rect 241 145 242 146
rect 240 145 241 146
rect 239 145 240 146
rect 218 145 219 146
rect 217 145 218 146
rect 216 145 217 146
rect 215 145 216 146
rect 214 145 215 146
rect 213 145 214 146
rect 212 145 213 146
rect 211 145 212 146
rect 210 145 211 146
rect 209 145 210 146
rect 208 145 209 146
rect 207 145 208 146
rect 206 145 207 146
rect 205 145 206 146
rect 204 145 205 146
rect 203 145 204 146
rect 202 145 203 146
rect 201 145 202 146
rect 200 145 201 146
rect 199 145 200 146
rect 198 145 199 146
rect 197 145 198 146
rect 196 145 197 146
rect 195 145 196 146
rect 194 145 195 146
rect 193 145 194 146
rect 192 145 193 146
rect 191 145 192 146
rect 190 145 191 146
rect 189 145 190 146
rect 188 145 189 146
rect 187 145 188 146
rect 186 145 187 146
rect 185 145 186 146
rect 184 145 185 146
rect 183 145 184 146
rect 182 145 183 146
rect 181 145 182 146
rect 180 145 181 146
rect 179 145 180 146
rect 178 145 179 146
rect 177 145 178 146
rect 176 145 177 146
rect 175 145 176 146
rect 174 145 175 146
rect 173 145 174 146
rect 172 145 173 146
rect 171 145 172 146
rect 170 145 171 146
rect 169 145 170 146
rect 168 145 169 146
rect 167 145 168 146
rect 166 145 167 146
rect 165 145 166 146
rect 164 145 165 146
rect 163 145 164 146
rect 162 145 163 146
rect 161 145 162 146
rect 160 145 161 146
rect 159 145 160 146
rect 158 145 159 146
rect 157 145 158 146
rect 156 145 157 146
rect 155 145 156 146
rect 154 145 155 146
rect 130 145 131 146
rect 129 145 130 146
rect 128 145 129 146
rect 127 145 128 146
rect 126 145 127 146
rect 125 145 126 146
rect 124 145 125 146
rect 123 145 124 146
rect 122 145 123 146
rect 121 145 122 146
rect 120 145 121 146
rect 119 145 120 146
rect 118 145 119 146
rect 117 145 118 146
rect 116 145 117 146
rect 115 145 116 146
rect 114 145 115 146
rect 113 145 114 146
rect 112 145 113 146
rect 111 145 112 146
rect 110 145 111 146
rect 109 145 110 146
rect 108 145 109 146
rect 107 145 108 146
rect 106 145 107 146
rect 105 145 106 146
rect 104 145 105 146
rect 103 145 104 146
rect 102 145 103 146
rect 101 145 102 146
rect 100 145 101 146
rect 99 145 100 146
rect 98 145 99 146
rect 97 145 98 146
rect 96 145 97 146
rect 95 145 96 146
rect 94 145 95 146
rect 93 145 94 146
rect 92 145 93 146
rect 91 145 92 146
rect 90 145 91 146
rect 89 145 90 146
rect 88 145 89 146
rect 87 145 88 146
rect 86 145 87 146
rect 85 145 86 146
rect 84 145 85 146
rect 83 145 84 146
rect 82 145 83 146
rect 81 145 82 146
rect 80 145 81 146
rect 79 145 80 146
rect 78 145 79 146
rect 77 145 78 146
rect 76 145 77 146
rect 75 145 76 146
rect 74 145 75 146
rect 73 145 74 146
rect 72 145 73 146
rect 71 145 72 146
rect 70 145 71 146
rect 69 145 70 146
rect 68 145 69 146
rect 67 145 68 146
rect 66 145 67 146
rect 65 145 66 146
rect 64 145 65 146
rect 63 145 64 146
rect 62 145 63 146
rect 61 145 62 146
rect 60 145 61 146
rect 59 145 60 146
rect 58 145 59 146
rect 57 145 58 146
rect 56 145 57 146
rect 55 145 56 146
rect 54 145 55 146
rect 53 145 54 146
rect 52 145 53 146
rect 51 145 52 146
rect 50 145 51 146
rect 49 145 50 146
rect 48 145 49 146
rect 47 145 48 146
rect 46 145 47 146
rect 45 145 46 146
rect 44 145 45 146
rect 43 145 44 146
rect 42 145 43 146
rect 41 145 42 146
rect 40 145 41 146
rect 39 145 40 146
rect 38 145 39 146
rect 27 145 28 146
rect 26 145 27 146
rect 25 145 26 146
rect 24 145 25 146
rect 23 145 24 146
rect 22 145 23 146
rect 21 145 22 146
rect 20 145 21 146
rect 19 145 20 146
rect 18 145 19 146
rect 17 145 18 146
rect 16 145 17 146
rect 15 145 16 146
rect 14 145 15 146
rect 13 145 14 146
rect 12 145 13 146
rect 11 145 12 146
rect 10 145 11 146
rect 478 146 479 147
rect 477 146 478 147
rect 476 146 477 147
rect 475 146 476 147
rect 474 146 475 147
rect 473 146 474 147
rect 472 146 473 147
rect 471 146 472 147
rect 470 146 471 147
rect 469 146 470 147
rect 468 146 469 147
rect 467 146 468 147
rect 466 146 467 147
rect 465 146 466 147
rect 464 146 465 147
rect 463 146 464 147
rect 462 146 463 147
rect 461 146 462 147
rect 460 146 461 147
rect 459 146 460 147
rect 458 146 459 147
rect 395 146 396 147
rect 394 146 395 147
rect 393 146 394 147
rect 317 146 318 147
rect 316 146 317 147
rect 315 146 316 147
rect 314 146 315 147
rect 313 146 314 147
rect 312 146 313 147
rect 311 146 312 147
rect 310 146 311 147
rect 309 146 310 147
rect 308 146 309 147
rect 307 146 308 147
rect 306 146 307 147
rect 305 146 306 147
rect 304 146 305 147
rect 303 146 304 147
rect 302 146 303 147
rect 301 146 302 147
rect 300 146 301 147
rect 299 146 300 147
rect 298 146 299 147
rect 297 146 298 147
rect 296 146 297 147
rect 295 146 296 147
rect 294 146 295 147
rect 293 146 294 147
rect 292 146 293 147
rect 291 146 292 147
rect 290 146 291 147
rect 289 146 290 147
rect 288 146 289 147
rect 287 146 288 147
rect 286 146 287 147
rect 285 146 286 147
rect 284 146 285 147
rect 283 146 284 147
rect 282 146 283 147
rect 281 146 282 147
rect 280 146 281 147
rect 279 146 280 147
rect 278 146 279 147
rect 277 146 278 147
rect 276 146 277 147
rect 275 146 276 147
rect 274 146 275 147
rect 273 146 274 147
rect 272 146 273 147
rect 271 146 272 147
rect 270 146 271 147
rect 269 146 270 147
rect 268 146 269 147
rect 267 146 268 147
rect 266 146 267 147
rect 265 146 266 147
rect 264 146 265 147
rect 263 146 264 147
rect 262 146 263 147
rect 261 146 262 147
rect 260 146 261 147
rect 259 146 260 147
rect 258 146 259 147
rect 257 146 258 147
rect 256 146 257 147
rect 255 146 256 147
rect 254 146 255 147
rect 253 146 254 147
rect 252 146 253 147
rect 251 146 252 147
rect 250 146 251 147
rect 249 146 250 147
rect 248 146 249 147
rect 247 146 248 147
rect 246 146 247 147
rect 245 146 246 147
rect 244 146 245 147
rect 243 146 244 147
rect 242 146 243 147
rect 241 146 242 147
rect 240 146 241 147
rect 239 146 240 147
rect 238 146 239 147
rect 217 146 218 147
rect 216 146 217 147
rect 215 146 216 147
rect 214 146 215 147
rect 213 146 214 147
rect 212 146 213 147
rect 211 146 212 147
rect 210 146 211 147
rect 209 146 210 147
rect 208 146 209 147
rect 207 146 208 147
rect 206 146 207 147
rect 205 146 206 147
rect 204 146 205 147
rect 203 146 204 147
rect 202 146 203 147
rect 201 146 202 147
rect 200 146 201 147
rect 199 146 200 147
rect 198 146 199 147
rect 197 146 198 147
rect 196 146 197 147
rect 195 146 196 147
rect 194 146 195 147
rect 193 146 194 147
rect 192 146 193 147
rect 191 146 192 147
rect 190 146 191 147
rect 189 146 190 147
rect 188 146 189 147
rect 187 146 188 147
rect 186 146 187 147
rect 185 146 186 147
rect 184 146 185 147
rect 183 146 184 147
rect 182 146 183 147
rect 181 146 182 147
rect 180 146 181 147
rect 179 146 180 147
rect 178 146 179 147
rect 177 146 178 147
rect 176 146 177 147
rect 175 146 176 147
rect 174 146 175 147
rect 173 146 174 147
rect 172 146 173 147
rect 171 146 172 147
rect 170 146 171 147
rect 169 146 170 147
rect 168 146 169 147
rect 167 146 168 147
rect 166 146 167 147
rect 165 146 166 147
rect 164 146 165 147
rect 163 146 164 147
rect 162 146 163 147
rect 161 146 162 147
rect 160 146 161 147
rect 159 146 160 147
rect 158 146 159 147
rect 157 146 158 147
rect 156 146 157 147
rect 155 146 156 147
rect 154 146 155 147
rect 153 146 154 147
rect 129 146 130 147
rect 128 146 129 147
rect 127 146 128 147
rect 126 146 127 147
rect 125 146 126 147
rect 124 146 125 147
rect 123 146 124 147
rect 122 146 123 147
rect 121 146 122 147
rect 120 146 121 147
rect 119 146 120 147
rect 118 146 119 147
rect 117 146 118 147
rect 116 146 117 147
rect 115 146 116 147
rect 114 146 115 147
rect 113 146 114 147
rect 112 146 113 147
rect 111 146 112 147
rect 110 146 111 147
rect 109 146 110 147
rect 108 146 109 147
rect 107 146 108 147
rect 106 146 107 147
rect 105 146 106 147
rect 104 146 105 147
rect 103 146 104 147
rect 102 146 103 147
rect 101 146 102 147
rect 100 146 101 147
rect 99 146 100 147
rect 98 146 99 147
rect 97 146 98 147
rect 96 146 97 147
rect 95 146 96 147
rect 94 146 95 147
rect 93 146 94 147
rect 92 146 93 147
rect 91 146 92 147
rect 90 146 91 147
rect 89 146 90 147
rect 88 146 89 147
rect 87 146 88 147
rect 86 146 87 147
rect 85 146 86 147
rect 84 146 85 147
rect 83 146 84 147
rect 82 146 83 147
rect 81 146 82 147
rect 80 146 81 147
rect 79 146 80 147
rect 78 146 79 147
rect 77 146 78 147
rect 76 146 77 147
rect 75 146 76 147
rect 74 146 75 147
rect 73 146 74 147
rect 72 146 73 147
rect 71 146 72 147
rect 70 146 71 147
rect 69 146 70 147
rect 68 146 69 147
rect 67 146 68 147
rect 66 146 67 147
rect 65 146 66 147
rect 64 146 65 147
rect 63 146 64 147
rect 62 146 63 147
rect 61 146 62 147
rect 60 146 61 147
rect 59 146 60 147
rect 58 146 59 147
rect 57 146 58 147
rect 56 146 57 147
rect 55 146 56 147
rect 54 146 55 147
rect 53 146 54 147
rect 52 146 53 147
rect 51 146 52 147
rect 50 146 51 147
rect 49 146 50 147
rect 48 146 49 147
rect 47 146 48 147
rect 46 146 47 147
rect 45 146 46 147
rect 44 146 45 147
rect 43 146 44 147
rect 42 146 43 147
rect 41 146 42 147
rect 40 146 41 147
rect 39 146 40 147
rect 38 146 39 147
rect 27 146 28 147
rect 26 146 27 147
rect 25 146 26 147
rect 24 146 25 147
rect 23 146 24 147
rect 22 146 23 147
rect 21 146 22 147
rect 20 146 21 147
rect 19 146 20 147
rect 18 146 19 147
rect 17 146 18 147
rect 16 146 17 147
rect 15 146 16 147
rect 14 146 15 147
rect 13 146 14 147
rect 12 146 13 147
rect 11 146 12 147
rect 10 146 11 147
rect 9 146 10 147
rect 478 147 479 148
rect 477 147 478 148
rect 476 147 477 148
rect 475 147 476 148
rect 474 147 475 148
rect 473 147 474 148
rect 472 147 473 148
rect 471 147 472 148
rect 470 147 471 148
rect 469 147 470 148
rect 468 147 469 148
rect 467 147 468 148
rect 466 147 467 148
rect 465 147 466 148
rect 464 147 465 148
rect 463 147 464 148
rect 462 147 463 148
rect 461 147 462 148
rect 460 147 461 148
rect 459 147 460 148
rect 458 147 459 148
rect 395 147 396 148
rect 394 147 395 148
rect 393 147 394 148
rect 317 147 318 148
rect 316 147 317 148
rect 315 147 316 148
rect 314 147 315 148
rect 313 147 314 148
rect 312 147 313 148
rect 311 147 312 148
rect 310 147 311 148
rect 309 147 310 148
rect 308 147 309 148
rect 307 147 308 148
rect 306 147 307 148
rect 305 147 306 148
rect 304 147 305 148
rect 303 147 304 148
rect 302 147 303 148
rect 301 147 302 148
rect 300 147 301 148
rect 299 147 300 148
rect 298 147 299 148
rect 297 147 298 148
rect 296 147 297 148
rect 295 147 296 148
rect 294 147 295 148
rect 293 147 294 148
rect 292 147 293 148
rect 291 147 292 148
rect 290 147 291 148
rect 289 147 290 148
rect 288 147 289 148
rect 287 147 288 148
rect 286 147 287 148
rect 285 147 286 148
rect 284 147 285 148
rect 283 147 284 148
rect 282 147 283 148
rect 281 147 282 148
rect 280 147 281 148
rect 279 147 280 148
rect 278 147 279 148
rect 277 147 278 148
rect 276 147 277 148
rect 275 147 276 148
rect 274 147 275 148
rect 273 147 274 148
rect 272 147 273 148
rect 271 147 272 148
rect 270 147 271 148
rect 269 147 270 148
rect 268 147 269 148
rect 267 147 268 148
rect 266 147 267 148
rect 265 147 266 148
rect 264 147 265 148
rect 263 147 264 148
rect 262 147 263 148
rect 261 147 262 148
rect 260 147 261 148
rect 259 147 260 148
rect 258 147 259 148
rect 257 147 258 148
rect 256 147 257 148
rect 255 147 256 148
rect 254 147 255 148
rect 253 147 254 148
rect 252 147 253 148
rect 251 147 252 148
rect 250 147 251 148
rect 249 147 250 148
rect 248 147 249 148
rect 247 147 248 148
rect 246 147 247 148
rect 245 147 246 148
rect 244 147 245 148
rect 243 147 244 148
rect 242 147 243 148
rect 241 147 242 148
rect 240 147 241 148
rect 239 147 240 148
rect 238 147 239 148
rect 217 147 218 148
rect 216 147 217 148
rect 215 147 216 148
rect 214 147 215 148
rect 213 147 214 148
rect 212 147 213 148
rect 211 147 212 148
rect 210 147 211 148
rect 209 147 210 148
rect 208 147 209 148
rect 207 147 208 148
rect 206 147 207 148
rect 205 147 206 148
rect 204 147 205 148
rect 203 147 204 148
rect 202 147 203 148
rect 201 147 202 148
rect 200 147 201 148
rect 199 147 200 148
rect 198 147 199 148
rect 197 147 198 148
rect 196 147 197 148
rect 195 147 196 148
rect 194 147 195 148
rect 193 147 194 148
rect 192 147 193 148
rect 191 147 192 148
rect 190 147 191 148
rect 189 147 190 148
rect 188 147 189 148
rect 187 147 188 148
rect 186 147 187 148
rect 185 147 186 148
rect 184 147 185 148
rect 183 147 184 148
rect 182 147 183 148
rect 181 147 182 148
rect 180 147 181 148
rect 179 147 180 148
rect 178 147 179 148
rect 177 147 178 148
rect 176 147 177 148
rect 175 147 176 148
rect 174 147 175 148
rect 173 147 174 148
rect 172 147 173 148
rect 171 147 172 148
rect 170 147 171 148
rect 169 147 170 148
rect 168 147 169 148
rect 167 147 168 148
rect 166 147 167 148
rect 165 147 166 148
rect 164 147 165 148
rect 163 147 164 148
rect 162 147 163 148
rect 161 147 162 148
rect 160 147 161 148
rect 159 147 160 148
rect 158 147 159 148
rect 157 147 158 148
rect 156 147 157 148
rect 155 147 156 148
rect 154 147 155 148
rect 153 147 154 148
rect 127 147 128 148
rect 126 147 127 148
rect 125 147 126 148
rect 124 147 125 148
rect 123 147 124 148
rect 122 147 123 148
rect 121 147 122 148
rect 120 147 121 148
rect 119 147 120 148
rect 118 147 119 148
rect 117 147 118 148
rect 116 147 117 148
rect 115 147 116 148
rect 114 147 115 148
rect 113 147 114 148
rect 112 147 113 148
rect 111 147 112 148
rect 110 147 111 148
rect 109 147 110 148
rect 108 147 109 148
rect 107 147 108 148
rect 106 147 107 148
rect 105 147 106 148
rect 104 147 105 148
rect 103 147 104 148
rect 102 147 103 148
rect 101 147 102 148
rect 100 147 101 148
rect 99 147 100 148
rect 98 147 99 148
rect 97 147 98 148
rect 96 147 97 148
rect 95 147 96 148
rect 94 147 95 148
rect 93 147 94 148
rect 92 147 93 148
rect 91 147 92 148
rect 90 147 91 148
rect 89 147 90 148
rect 88 147 89 148
rect 87 147 88 148
rect 86 147 87 148
rect 85 147 86 148
rect 84 147 85 148
rect 83 147 84 148
rect 82 147 83 148
rect 81 147 82 148
rect 80 147 81 148
rect 79 147 80 148
rect 78 147 79 148
rect 77 147 78 148
rect 76 147 77 148
rect 75 147 76 148
rect 74 147 75 148
rect 73 147 74 148
rect 72 147 73 148
rect 71 147 72 148
rect 70 147 71 148
rect 69 147 70 148
rect 68 147 69 148
rect 67 147 68 148
rect 66 147 67 148
rect 65 147 66 148
rect 64 147 65 148
rect 63 147 64 148
rect 62 147 63 148
rect 61 147 62 148
rect 60 147 61 148
rect 59 147 60 148
rect 58 147 59 148
rect 57 147 58 148
rect 56 147 57 148
rect 55 147 56 148
rect 54 147 55 148
rect 53 147 54 148
rect 52 147 53 148
rect 51 147 52 148
rect 50 147 51 148
rect 49 147 50 148
rect 48 147 49 148
rect 47 147 48 148
rect 46 147 47 148
rect 45 147 46 148
rect 44 147 45 148
rect 43 147 44 148
rect 42 147 43 148
rect 41 147 42 148
rect 40 147 41 148
rect 39 147 40 148
rect 38 147 39 148
rect 37 147 38 148
rect 27 147 28 148
rect 26 147 27 148
rect 25 147 26 148
rect 24 147 25 148
rect 23 147 24 148
rect 22 147 23 148
rect 21 147 22 148
rect 20 147 21 148
rect 19 147 20 148
rect 18 147 19 148
rect 17 147 18 148
rect 16 147 17 148
rect 15 147 16 148
rect 14 147 15 148
rect 13 147 14 148
rect 12 147 13 148
rect 11 147 12 148
rect 10 147 11 148
rect 9 147 10 148
rect 478 148 479 149
rect 458 148 459 149
rect 318 148 319 149
rect 317 148 318 149
rect 316 148 317 149
rect 315 148 316 149
rect 314 148 315 149
rect 313 148 314 149
rect 312 148 313 149
rect 311 148 312 149
rect 310 148 311 149
rect 309 148 310 149
rect 308 148 309 149
rect 307 148 308 149
rect 306 148 307 149
rect 305 148 306 149
rect 304 148 305 149
rect 303 148 304 149
rect 302 148 303 149
rect 301 148 302 149
rect 300 148 301 149
rect 299 148 300 149
rect 298 148 299 149
rect 297 148 298 149
rect 296 148 297 149
rect 295 148 296 149
rect 294 148 295 149
rect 293 148 294 149
rect 292 148 293 149
rect 291 148 292 149
rect 290 148 291 149
rect 289 148 290 149
rect 288 148 289 149
rect 287 148 288 149
rect 286 148 287 149
rect 285 148 286 149
rect 284 148 285 149
rect 283 148 284 149
rect 282 148 283 149
rect 281 148 282 149
rect 280 148 281 149
rect 279 148 280 149
rect 278 148 279 149
rect 277 148 278 149
rect 276 148 277 149
rect 275 148 276 149
rect 274 148 275 149
rect 273 148 274 149
rect 272 148 273 149
rect 271 148 272 149
rect 270 148 271 149
rect 269 148 270 149
rect 268 148 269 149
rect 267 148 268 149
rect 266 148 267 149
rect 265 148 266 149
rect 264 148 265 149
rect 263 148 264 149
rect 262 148 263 149
rect 261 148 262 149
rect 260 148 261 149
rect 259 148 260 149
rect 258 148 259 149
rect 257 148 258 149
rect 256 148 257 149
rect 255 148 256 149
rect 254 148 255 149
rect 253 148 254 149
rect 252 148 253 149
rect 251 148 252 149
rect 250 148 251 149
rect 249 148 250 149
rect 248 148 249 149
rect 247 148 248 149
rect 246 148 247 149
rect 245 148 246 149
rect 244 148 245 149
rect 243 148 244 149
rect 242 148 243 149
rect 241 148 242 149
rect 240 148 241 149
rect 239 148 240 149
rect 238 148 239 149
rect 237 148 238 149
rect 216 148 217 149
rect 215 148 216 149
rect 214 148 215 149
rect 213 148 214 149
rect 212 148 213 149
rect 211 148 212 149
rect 210 148 211 149
rect 209 148 210 149
rect 208 148 209 149
rect 207 148 208 149
rect 206 148 207 149
rect 205 148 206 149
rect 204 148 205 149
rect 203 148 204 149
rect 202 148 203 149
rect 201 148 202 149
rect 200 148 201 149
rect 199 148 200 149
rect 198 148 199 149
rect 197 148 198 149
rect 196 148 197 149
rect 195 148 196 149
rect 194 148 195 149
rect 193 148 194 149
rect 192 148 193 149
rect 191 148 192 149
rect 190 148 191 149
rect 189 148 190 149
rect 188 148 189 149
rect 187 148 188 149
rect 186 148 187 149
rect 185 148 186 149
rect 184 148 185 149
rect 183 148 184 149
rect 182 148 183 149
rect 181 148 182 149
rect 180 148 181 149
rect 179 148 180 149
rect 178 148 179 149
rect 177 148 178 149
rect 176 148 177 149
rect 175 148 176 149
rect 174 148 175 149
rect 173 148 174 149
rect 172 148 173 149
rect 171 148 172 149
rect 170 148 171 149
rect 169 148 170 149
rect 168 148 169 149
rect 167 148 168 149
rect 166 148 167 149
rect 165 148 166 149
rect 164 148 165 149
rect 163 148 164 149
rect 162 148 163 149
rect 161 148 162 149
rect 160 148 161 149
rect 159 148 160 149
rect 158 148 159 149
rect 157 148 158 149
rect 156 148 157 149
rect 155 148 156 149
rect 154 148 155 149
rect 153 148 154 149
rect 152 148 153 149
rect 126 148 127 149
rect 125 148 126 149
rect 124 148 125 149
rect 123 148 124 149
rect 122 148 123 149
rect 121 148 122 149
rect 120 148 121 149
rect 119 148 120 149
rect 118 148 119 149
rect 117 148 118 149
rect 116 148 117 149
rect 115 148 116 149
rect 114 148 115 149
rect 113 148 114 149
rect 112 148 113 149
rect 111 148 112 149
rect 110 148 111 149
rect 109 148 110 149
rect 108 148 109 149
rect 107 148 108 149
rect 106 148 107 149
rect 105 148 106 149
rect 104 148 105 149
rect 103 148 104 149
rect 102 148 103 149
rect 101 148 102 149
rect 100 148 101 149
rect 99 148 100 149
rect 98 148 99 149
rect 97 148 98 149
rect 96 148 97 149
rect 95 148 96 149
rect 94 148 95 149
rect 93 148 94 149
rect 92 148 93 149
rect 91 148 92 149
rect 90 148 91 149
rect 89 148 90 149
rect 88 148 89 149
rect 87 148 88 149
rect 86 148 87 149
rect 85 148 86 149
rect 84 148 85 149
rect 83 148 84 149
rect 82 148 83 149
rect 81 148 82 149
rect 80 148 81 149
rect 79 148 80 149
rect 78 148 79 149
rect 77 148 78 149
rect 76 148 77 149
rect 75 148 76 149
rect 74 148 75 149
rect 73 148 74 149
rect 72 148 73 149
rect 71 148 72 149
rect 70 148 71 149
rect 69 148 70 149
rect 68 148 69 149
rect 67 148 68 149
rect 66 148 67 149
rect 65 148 66 149
rect 64 148 65 149
rect 63 148 64 149
rect 62 148 63 149
rect 61 148 62 149
rect 60 148 61 149
rect 59 148 60 149
rect 58 148 59 149
rect 57 148 58 149
rect 56 148 57 149
rect 55 148 56 149
rect 54 148 55 149
rect 53 148 54 149
rect 52 148 53 149
rect 51 148 52 149
rect 50 148 51 149
rect 49 148 50 149
rect 48 148 49 149
rect 47 148 48 149
rect 46 148 47 149
rect 45 148 46 149
rect 44 148 45 149
rect 43 148 44 149
rect 42 148 43 149
rect 41 148 42 149
rect 40 148 41 149
rect 39 148 40 149
rect 38 148 39 149
rect 37 148 38 149
rect 27 148 28 149
rect 26 148 27 149
rect 25 148 26 149
rect 24 148 25 149
rect 23 148 24 149
rect 22 148 23 149
rect 21 148 22 149
rect 20 148 21 149
rect 19 148 20 149
rect 18 148 19 149
rect 17 148 18 149
rect 16 148 17 149
rect 15 148 16 149
rect 14 148 15 149
rect 13 148 14 149
rect 12 148 13 149
rect 11 148 12 149
rect 10 148 11 149
rect 9 148 10 149
rect 8 148 9 149
rect 478 149 479 150
rect 458 149 459 150
rect 319 149 320 150
rect 318 149 319 150
rect 317 149 318 150
rect 316 149 317 150
rect 315 149 316 150
rect 314 149 315 150
rect 313 149 314 150
rect 312 149 313 150
rect 311 149 312 150
rect 310 149 311 150
rect 309 149 310 150
rect 308 149 309 150
rect 307 149 308 150
rect 306 149 307 150
rect 305 149 306 150
rect 304 149 305 150
rect 303 149 304 150
rect 302 149 303 150
rect 301 149 302 150
rect 300 149 301 150
rect 299 149 300 150
rect 298 149 299 150
rect 297 149 298 150
rect 296 149 297 150
rect 295 149 296 150
rect 294 149 295 150
rect 293 149 294 150
rect 292 149 293 150
rect 291 149 292 150
rect 290 149 291 150
rect 289 149 290 150
rect 288 149 289 150
rect 287 149 288 150
rect 286 149 287 150
rect 285 149 286 150
rect 284 149 285 150
rect 283 149 284 150
rect 282 149 283 150
rect 281 149 282 150
rect 280 149 281 150
rect 279 149 280 150
rect 278 149 279 150
rect 277 149 278 150
rect 276 149 277 150
rect 275 149 276 150
rect 274 149 275 150
rect 273 149 274 150
rect 272 149 273 150
rect 271 149 272 150
rect 270 149 271 150
rect 269 149 270 150
rect 268 149 269 150
rect 267 149 268 150
rect 266 149 267 150
rect 265 149 266 150
rect 264 149 265 150
rect 263 149 264 150
rect 262 149 263 150
rect 261 149 262 150
rect 260 149 261 150
rect 259 149 260 150
rect 258 149 259 150
rect 257 149 258 150
rect 256 149 257 150
rect 255 149 256 150
rect 254 149 255 150
rect 253 149 254 150
rect 252 149 253 150
rect 251 149 252 150
rect 250 149 251 150
rect 249 149 250 150
rect 248 149 249 150
rect 247 149 248 150
rect 246 149 247 150
rect 245 149 246 150
rect 244 149 245 150
rect 243 149 244 150
rect 242 149 243 150
rect 241 149 242 150
rect 240 149 241 150
rect 239 149 240 150
rect 238 149 239 150
rect 237 149 238 150
rect 236 149 237 150
rect 216 149 217 150
rect 215 149 216 150
rect 214 149 215 150
rect 213 149 214 150
rect 212 149 213 150
rect 211 149 212 150
rect 210 149 211 150
rect 209 149 210 150
rect 208 149 209 150
rect 207 149 208 150
rect 206 149 207 150
rect 205 149 206 150
rect 204 149 205 150
rect 203 149 204 150
rect 202 149 203 150
rect 201 149 202 150
rect 200 149 201 150
rect 199 149 200 150
rect 198 149 199 150
rect 197 149 198 150
rect 196 149 197 150
rect 195 149 196 150
rect 194 149 195 150
rect 193 149 194 150
rect 192 149 193 150
rect 191 149 192 150
rect 190 149 191 150
rect 189 149 190 150
rect 188 149 189 150
rect 187 149 188 150
rect 186 149 187 150
rect 185 149 186 150
rect 184 149 185 150
rect 183 149 184 150
rect 182 149 183 150
rect 181 149 182 150
rect 180 149 181 150
rect 179 149 180 150
rect 178 149 179 150
rect 177 149 178 150
rect 176 149 177 150
rect 175 149 176 150
rect 174 149 175 150
rect 173 149 174 150
rect 172 149 173 150
rect 171 149 172 150
rect 170 149 171 150
rect 169 149 170 150
rect 168 149 169 150
rect 167 149 168 150
rect 166 149 167 150
rect 165 149 166 150
rect 164 149 165 150
rect 163 149 164 150
rect 162 149 163 150
rect 161 149 162 150
rect 160 149 161 150
rect 159 149 160 150
rect 158 149 159 150
rect 157 149 158 150
rect 156 149 157 150
rect 155 149 156 150
rect 154 149 155 150
rect 153 149 154 150
rect 152 149 153 150
rect 151 149 152 150
rect 124 149 125 150
rect 123 149 124 150
rect 122 149 123 150
rect 121 149 122 150
rect 120 149 121 150
rect 119 149 120 150
rect 118 149 119 150
rect 117 149 118 150
rect 116 149 117 150
rect 115 149 116 150
rect 114 149 115 150
rect 113 149 114 150
rect 112 149 113 150
rect 111 149 112 150
rect 110 149 111 150
rect 109 149 110 150
rect 108 149 109 150
rect 107 149 108 150
rect 106 149 107 150
rect 105 149 106 150
rect 104 149 105 150
rect 103 149 104 150
rect 102 149 103 150
rect 101 149 102 150
rect 100 149 101 150
rect 99 149 100 150
rect 98 149 99 150
rect 97 149 98 150
rect 96 149 97 150
rect 95 149 96 150
rect 94 149 95 150
rect 93 149 94 150
rect 92 149 93 150
rect 91 149 92 150
rect 90 149 91 150
rect 89 149 90 150
rect 88 149 89 150
rect 87 149 88 150
rect 86 149 87 150
rect 85 149 86 150
rect 84 149 85 150
rect 83 149 84 150
rect 82 149 83 150
rect 81 149 82 150
rect 80 149 81 150
rect 79 149 80 150
rect 78 149 79 150
rect 77 149 78 150
rect 76 149 77 150
rect 75 149 76 150
rect 74 149 75 150
rect 73 149 74 150
rect 72 149 73 150
rect 71 149 72 150
rect 70 149 71 150
rect 69 149 70 150
rect 68 149 69 150
rect 67 149 68 150
rect 66 149 67 150
rect 65 149 66 150
rect 64 149 65 150
rect 63 149 64 150
rect 62 149 63 150
rect 61 149 62 150
rect 60 149 61 150
rect 59 149 60 150
rect 58 149 59 150
rect 57 149 58 150
rect 56 149 57 150
rect 55 149 56 150
rect 54 149 55 150
rect 53 149 54 150
rect 52 149 53 150
rect 51 149 52 150
rect 50 149 51 150
rect 49 149 50 150
rect 48 149 49 150
rect 47 149 48 150
rect 46 149 47 150
rect 45 149 46 150
rect 44 149 45 150
rect 43 149 44 150
rect 42 149 43 150
rect 41 149 42 150
rect 40 149 41 150
rect 39 149 40 150
rect 38 149 39 150
rect 37 149 38 150
rect 36 149 37 150
rect 27 149 28 150
rect 26 149 27 150
rect 25 149 26 150
rect 24 149 25 150
rect 23 149 24 150
rect 22 149 23 150
rect 21 149 22 150
rect 20 149 21 150
rect 19 149 20 150
rect 18 149 19 150
rect 17 149 18 150
rect 16 149 17 150
rect 15 149 16 150
rect 14 149 15 150
rect 13 149 14 150
rect 12 149 13 150
rect 11 149 12 150
rect 10 149 11 150
rect 9 149 10 150
rect 8 149 9 150
rect 7 149 8 150
rect 320 150 321 151
rect 319 150 320 151
rect 318 150 319 151
rect 317 150 318 151
rect 316 150 317 151
rect 315 150 316 151
rect 314 150 315 151
rect 313 150 314 151
rect 312 150 313 151
rect 311 150 312 151
rect 310 150 311 151
rect 309 150 310 151
rect 308 150 309 151
rect 307 150 308 151
rect 306 150 307 151
rect 305 150 306 151
rect 304 150 305 151
rect 303 150 304 151
rect 302 150 303 151
rect 301 150 302 151
rect 300 150 301 151
rect 299 150 300 151
rect 298 150 299 151
rect 297 150 298 151
rect 296 150 297 151
rect 295 150 296 151
rect 294 150 295 151
rect 293 150 294 151
rect 292 150 293 151
rect 291 150 292 151
rect 290 150 291 151
rect 289 150 290 151
rect 288 150 289 151
rect 287 150 288 151
rect 286 150 287 151
rect 285 150 286 151
rect 284 150 285 151
rect 283 150 284 151
rect 282 150 283 151
rect 281 150 282 151
rect 280 150 281 151
rect 279 150 280 151
rect 278 150 279 151
rect 277 150 278 151
rect 276 150 277 151
rect 275 150 276 151
rect 274 150 275 151
rect 273 150 274 151
rect 272 150 273 151
rect 271 150 272 151
rect 270 150 271 151
rect 269 150 270 151
rect 268 150 269 151
rect 267 150 268 151
rect 266 150 267 151
rect 265 150 266 151
rect 264 150 265 151
rect 263 150 264 151
rect 262 150 263 151
rect 261 150 262 151
rect 260 150 261 151
rect 259 150 260 151
rect 258 150 259 151
rect 257 150 258 151
rect 256 150 257 151
rect 255 150 256 151
rect 254 150 255 151
rect 253 150 254 151
rect 252 150 253 151
rect 251 150 252 151
rect 250 150 251 151
rect 249 150 250 151
rect 248 150 249 151
rect 247 150 248 151
rect 246 150 247 151
rect 245 150 246 151
rect 244 150 245 151
rect 243 150 244 151
rect 242 150 243 151
rect 241 150 242 151
rect 240 150 241 151
rect 239 150 240 151
rect 238 150 239 151
rect 237 150 238 151
rect 236 150 237 151
rect 216 150 217 151
rect 215 150 216 151
rect 214 150 215 151
rect 213 150 214 151
rect 212 150 213 151
rect 211 150 212 151
rect 210 150 211 151
rect 209 150 210 151
rect 208 150 209 151
rect 207 150 208 151
rect 206 150 207 151
rect 205 150 206 151
rect 204 150 205 151
rect 203 150 204 151
rect 202 150 203 151
rect 201 150 202 151
rect 200 150 201 151
rect 199 150 200 151
rect 198 150 199 151
rect 197 150 198 151
rect 196 150 197 151
rect 195 150 196 151
rect 194 150 195 151
rect 193 150 194 151
rect 192 150 193 151
rect 191 150 192 151
rect 190 150 191 151
rect 189 150 190 151
rect 188 150 189 151
rect 187 150 188 151
rect 186 150 187 151
rect 185 150 186 151
rect 184 150 185 151
rect 183 150 184 151
rect 182 150 183 151
rect 181 150 182 151
rect 180 150 181 151
rect 179 150 180 151
rect 178 150 179 151
rect 177 150 178 151
rect 176 150 177 151
rect 175 150 176 151
rect 174 150 175 151
rect 173 150 174 151
rect 172 150 173 151
rect 171 150 172 151
rect 170 150 171 151
rect 169 150 170 151
rect 168 150 169 151
rect 167 150 168 151
rect 166 150 167 151
rect 165 150 166 151
rect 164 150 165 151
rect 163 150 164 151
rect 162 150 163 151
rect 161 150 162 151
rect 160 150 161 151
rect 159 150 160 151
rect 158 150 159 151
rect 157 150 158 151
rect 156 150 157 151
rect 155 150 156 151
rect 154 150 155 151
rect 153 150 154 151
rect 152 150 153 151
rect 151 150 152 151
rect 150 150 151 151
rect 122 150 123 151
rect 121 150 122 151
rect 120 150 121 151
rect 119 150 120 151
rect 118 150 119 151
rect 117 150 118 151
rect 116 150 117 151
rect 115 150 116 151
rect 114 150 115 151
rect 113 150 114 151
rect 112 150 113 151
rect 111 150 112 151
rect 110 150 111 151
rect 109 150 110 151
rect 108 150 109 151
rect 107 150 108 151
rect 106 150 107 151
rect 105 150 106 151
rect 104 150 105 151
rect 103 150 104 151
rect 102 150 103 151
rect 101 150 102 151
rect 100 150 101 151
rect 99 150 100 151
rect 98 150 99 151
rect 97 150 98 151
rect 96 150 97 151
rect 95 150 96 151
rect 94 150 95 151
rect 93 150 94 151
rect 92 150 93 151
rect 91 150 92 151
rect 90 150 91 151
rect 89 150 90 151
rect 88 150 89 151
rect 87 150 88 151
rect 86 150 87 151
rect 85 150 86 151
rect 84 150 85 151
rect 83 150 84 151
rect 82 150 83 151
rect 81 150 82 151
rect 80 150 81 151
rect 79 150 80 151
rect 78 150 79 151
rect 77 150 78 151
rect 76 150 77 151
rect 75 150 76 151
rect 74 150 75 151
rect 73 150 74 151
rect 72 150 73 151
rect 71 150 72 151
rect 70 150 71 151
rect 69 150 70 151
rect 68 150 69 151
rect 67 150 68 151
rect 66 150 67 151
rect 65 150 66 151
rect 64 150 65 151
rect 63 150 64 151
rect 62 150 63 151
rect 61 150 62 151
rect 60 150 61 151
rect 59 150 60 151
rect 58 150 59 151
rect 57 150 58 151
rect 56 150 57 151
rect 55 150 56 151
rect 54 150 55 151
rect 53 150 54 151
rect 52 150 53 151
rect 51 150 52 151
rect 50 150 51 151
rect 49 150 50 151
rect 48 150 49 151
rect 47 150 48 151
rect 46 150 47 151
rect 45 150 46 151
rect 44 150 45 151
rect 43 150 44 151
rect 42 150 43 151
rect 41 150 42 151
rect 40 150 41 151
rect 39 150 40 151
rect 38 150 39 151
rect 37 150 38 151
rect 36 150 37 151
rect 26 150 27 151
rect 25 150 26 151
rect 24 150 25 151
rect 23 150 24 151
rect 22 150 23 151
rect 21 150 22 151
rect 20 150 21 151
rect 19 150 20 151
rect 18 150 19 151
rect 17 150 18 151
rect 16 150 17 151
rect 15 150 16 151
rect 14 150 15 151
rect 13 150 14 151
rect 12 150 13 151
rect 11 150 12 151
rect 10 150 11 151
rect 9 150 10 151
rect 8 150 9 151
rect 7 150 8 151
rect 321 151 322 152
rect 320 151 321 152
rect 319 151 320 152
rect 318 151 319 152
rect 317 151 318 152
rect 316 151 317 152
rect 315 151 316 152
rect 314 151 315 152
rect 313 151 314 152
rect 312 151 313 152
rect 311 151 312 152
rect 310 151 311 152
rect 309 151 310 152
rect 308 151 309 152
rect 307 151 308 152
rect 306 151 307 152
rect 305 151 306 152
rect 304 151 305 152
rect 303 151 304 152
rect 302 151 303 152
rect 301 151 302 152
rect 300 151 301 152
rect 299 151 300 152
rect 298 151 299 152
rect 297 151 298 152
rect 296 151 297 152
rect 295 151 296 152
rect 294 151 295 152
rect 293 151 294 152
rect 292 151 293 152
rect 291 151 292 152
rect 290 151 291 152
rect 289 151 290 152
rect 288 151 289 152
rect 287 151 288 152
rect 286 151 287 152
rect 285 151 286 152
rect 284 151 285 152
rect 283 151 284 152
rect 282 151 283 152
rect 281 151 282 152
rect 280 151 281 152
rect 279 151 280 152
rect 278 151 279 152
rect 277 151 278 152
rect 276 151 277 152
rect 275 151 276 152
rect 274 151 275 152
rect 273 151 274 152
rect 272 151 273 152
rect 271 151 272 152
rect 270 151 271 152
rect 269 151 270 152
rect 268 151 269 152
rect 267 151 268 152
rect 266 151 267 152
rect 265 151 266 152
rect 264 151 265 152
rect 263 151 264 152
rect 262 151 263 152
rect 261 151 262 152
rect 260 151 261 152
rect 259 151 260 152
rect 258 151 259 152
rect 257 151 258 152
rect 256 151 257 152
rect 255 151 256 152
rect 254 151 255 152
rect 253 151 254 152
rect 252 151 253 152
rect 251 151 252 152
rect 250 151 251 152
rect 249 151 250 152
rect 248 151 249 152
rect 247 151 248 152
rect 246 151 247 152
rect 245 151 246 152
rect 244 151 245 152
rect 243 151 244 152
rect 242 151 243 152
rect 241 151 242 152
rect 240 151 241 152
rect 239 151 240 152
rect 238 151 239 152
rect 237 151 238 152
rect 236 151 237 152
rect 235 151 236 152
rect 215 151 216 152
rect 214 151 215 152
rect 213 151 214 152
rect 212 151 213 152
rect 211 151 212 152
rect 210 151 211 152
rect 209 151 210 152
rect 208 151 209 152
rect 207 151 208 152
rect 206 151 207 152
rect 205 151 206 152
rect 204 151 205 152
rect 203 151 204 152
rect 202 151 203 152
rect 201 151 202 152
rect 200 151 201 152
rect 199 151 200 152
rect 198 151 199 152
rect 197 151 198 152
rect 196 151 197 152
rect 195 151 196 152
rect 194 151 195 152
rect 193 151 194 152
rect 192 151 193 152
rect 191 151 192 152
rect 190 151 191 152
rect 189 151 190 152
rect 188 151 189 152
rect 187 151 188 152
rect 186 151 187 152
rect 185 151 186 152
rect 184 151 185 152
rect 183 151 184 152
rect 182 151 183 152
rect 181 151 182 152
rect 180 151 181 152
rect 179 151 180 152
rect 178 151 179 152
rect 177 151 178 152
rect 176 151 177 152
rect 175 151 176 152
rect 174 151 175 152
rect 173 151 174 152
rect 172 151 173 152
rect 171 151 172 152
rect 170 151 171 152
rect 169 151 170 152
rect 168 151 169 152
rect 167 151 168 152
rect 166 151 167 152
rect 165 151 166 152
rect 164 151 165 152
rect 163 151 164 152
rect 162 151 163 152
rect 161 151 162 152
rect 160 151 161 152
rect 159 151 160 152
rect 158 151 159 152
rect 157 151 158 152
rect 156 151 157 152
rect 155 151 156 152
rect 154 151 155 152
rect 153 151 154 152
rect 152 151 153 152
rect 151 151 152 152
rect 150 151 151 152
rect 121 151 122 152
rect 120 151 121 152
rect 119 151 120 152
rect 118 151 119 152
rect 117 151 118 152
rect 116 151 117 152
rect 115 151 116 152
rect 114 151 115 152
rect 113 151 114 152
rect 112 151 113 152
rect 111 151 112 152
rect 110 151 111 152
rect 109 151 110 152
rect 108 151 109 152
rect 107 151 108 152
rect 106 151 107 152
rect 105 151 106 152
rect 104 151 105 152
rect 103 151 104 152
rect 102 151 103 152
rect 101 151 102 152
rect 100 151 101 152
rect 99 151 100 152
rect 98 151 99 152
rect 97 151 98 152
rect 96 151 97 152
rect 95 151 96 152
rect 94 151 95 152
rect 93 151 94 152
rect 92 151 93 152
rect 91 151 92 152
rect 90 151 91 152
rect 89 151 90 152
rect 88 151 89 152
rect 87 151 88 152
rect 86 151 87 152
rect 85 151 86 152
rect 84 151 85 152
rect 83 151 84 152
rect 82 151 83 152
rect 81 151 82 152
rect 80 151 81 152
rect 79 151 80 152
rect 78 151 79 152
rect 77 151 78 152
rect 76 151 77 152
rect 75 151 76 152
rect 74 151 75 152
rect 73 151 74 152
rect 72 151 73 152
rect 71 151 72 152
rect 70 151 71 152
rect 69 151 70 152
rect 68 151 69 152
rect 67 151 68 152
rect 66 151 67 152
rect 65 151 66 152
rect 64 151 65 152
rect 63 151 64 152
rect 62 151 63 152
rect 61 151 62 152
rect 60 151 61 152
rect 59 151 60 152
rect 58 151 59 152
rect 57 151 58 152
rect 56 151 57 152
rect 55 151 56 152
rect 54 151 55 152
rect 53 151 54 152
rect 52 151 53 152
rect 51 151 52 152
rect 50 151 51 152
rect 49 151 50 152
rect 48 151 49 152
rect 47 151 48 152
rect 46 151 47 152
rect 45 151 46 152
rect 44 151 45 152
rect 43 151 44 152
rect 42 151 43 152
rect 41 151 42 152
rect 40 151 41 152
rect 39 151 40 152
rect 38 151 39 152
rect 37 151 38 152
rect 36 151 37 152
rect 35 151 36 152
rect 26 151 27 152
rect 25 151 26 152
rect 24 151 25 152
rect 23 151 24 152
rect 22 151 23 152
rect 21 151 22 152
rect 20 151 21 152
rect 19 151 20 152
rect 18 151 19 152
rect 17 151 18 152
rect 16 151 17 152
rect 15 151 16 152
rect 14 151 15 152
rect 13 151 14 152
rect 12 151 13 152
rect 11 151 12 152
rect 10 151 11 152
rect 9 151 10 152
rect 8 151 9 152
rect 7 151 8 152
rect 6 151 7 152
rect 394 152 395 153
rect 393 152 394 153
rect 321 152 322 153
rect 320 152 321 153
rect 319 152 320 153
rect 318 152 319 153
rect 317 152 318 153
rect 316 152 317 153
rect 315 152 316 153
rect 314 152 315 153
rect 313 152 314 153
rect 312 152 313 153
rect 311 152 312 153
rect 310 152 311 153
rect 309 152 310 153
rect 308 152 309 153
rect 307 152 308 153
rect 306 152 307 153
rect 305 152 306 153
rect 304 152 305 153
rect 303 152 304 153
rect 302 152 303 153
rect 301 152 302 153
rect 300 152 301 153
rect 299 152 300 153
rect 298 152 299 153
rect 297 152 298 153
rect 296 152 297 153
rect 295 152 296 153
rect 294 152 295 153
rect 293 152 294 153
rect 292 152 293 153
rect 291 152 292 153
rect 290 152 291 153
rect 289 152 290 153
rect 288 152 289 153
rect 287 152 288 153
rect 286 152 287 153
rect 285 152 286 153
rect 284 152 285 153
rect 283 152 284 153
rect 282 152 283 153
rect 281 152 282 153
rect 280 152 281 153
rect 279 152 280 153
rect 278 152 279 153
rect 277 152 278 153
rect 276 152 277 153
rect 275 152 276 153
rect 274 152 275 153
rect 273 152 274 153
rect 272 152 273 153
rect 271 152 272 153
rect 270 152 271 153
rect 269 152 270 153
rect 268 152 269 153
rect 267 152 268 153
rect 266 152 267 153
rect 265 152 266 153
rect 264 152 265 153
rect 263 152 264 153
rect 262 152 263 153
rect 261 152 262 153
rect 260 152 261 153
rect 259 152 260 153
rect 258 152 259 153
rect 257 152 258 153
rect 256 152 257 153
rect 255 152 256 153
rect 254 152 255 153
rect 253 152 254 153
rect 252 152 253 153
rect 251 152 252 153
rect 250 152 251 153
rect 249 152 250 153
rect 248 152 249 153
rect 247 152 248 153
rect 246 152 247 153
rect 245 152 246 153
rect 244 152 245 153
rect 243 152 244 153
rect 242 152 243 153
rect 241 152 242 153
rect 240 152 241 153
rect 239 152 240 153
rect 238 152 239 153
rect 237 152 238 153
rect 236 152 237 153
rect 235 152 236 153
rect 234 152 235 153
rect 215 152 216 153
rect 214 152 215 153
rect 213 152 214 153
rect 212 152 213 153
rect 211 152 212 153
rect 210 152 211 153
rect 209 152 210 153
rect 208 152 209 153
rect 207 152 208 153
rect 206 152 207 153
rect 205 152 206 153
rect 204 152 205 153
rect 203 152 204 153
rect 202 152 203 153
rect 201 152 202 153
rect 200 152 201 153
rect 199 152 200 153
rect 198 152 199 153
rect 197 152 198 153
rect 196 152 197 153
rect 195 152 196 153
rect 194 152 195 153
rect 193 152 194 153
rect 192 152 193 153
rect 191 152 192 153
rect 190 152 191 153
rect 189 152 190 153
rect 188 152 189 153
rect 187 152 188 153
rect 186 152 187 153
rect 185 152 186 153
rect 184 152 185 153
rect 183 152 184 153
rect 182 152 183 153
rect 181 152 182 153
rect 180 152 181 153
rect 179 152 180 153
rect 178 152 179 153
rect 177 152 178 153
rect 176 152 177 153
rect 175 152 176 153
rect 174 152 175 153
rect 173 152 174 153
rect 172 152 173 153
rect 171 152 172 153
rect 170 152 171 153
rect 169 152 170 153
rect 168 152 169 153
rect 167 152 168 153
rect 166 152 167 153
rect 165 152 166 153
rect 164 152 165 153
rect 163 152 164 153
rect 162 152 163 153
rect 161 152 162 153
rect 160 152 161 153
rect 159 152 160 153
rect 158 152 159 153
rect 157 152 158 153
rect 156 152 157 153
rect 155 152 156 153
rect 154 152 155 153
rect 153 152 154 153
rect 152 152 153 153
rect 151 152 152 153
rect 150 152 151 153
rect 149 152 150 153
rect 119 152 120 153
rect 118 152 119 153
rect 117 152 118 153
rect 116 152 117 153
rect 115 152 116 153
rect 114 152 115 153
rect 113 152 114 153
rect 112 152 113 153
rect 111 152 112 153
rect 110 152 111 153
rect 109 152 110 153
rect 108 152 109 153
rect 107 152 108 153
rect 106 152 107 153
rect 105 152 106 153
rect 104 152 105 153
rect 103 152 104 153
rect 102 152 103 153
rect 101 152 102 153
rect 100 152 101 153
rect 99 152 100 153
rect 98 152 99 153
rect 97 152 98 153
rect 96 152 97 153
rect 95 152 96 153
rect 94 152 95 153
rect 93 152 94 153
rect 92 152 93 153
rect 91 152 92 153
rect 90 152 91 153
rect 89 152 90 153
rect 88 152 89 153
rect 87 152 88 153
rect 86 152 87 153
rect 85 152 86 153
rect 84 152 85 153
rect 83 152 84 153
rect 82 152 83 153
rect 81 152 82 153
rect 80 152 81 153
rect 79 152 80 153
rect 78 152 79 153
rect 77 152 78 153
rect 76 152 77 153
rect 75 152 76 153
rect 74 152 75 153
rect 73 152 74 153
rect 72 152 73 153
rect 71 152 72 153
rect 70 152 71 153
rect 69 152 70 153
rect 68 152 69 153
rect 67 152 68 153
rect 66 152 67 153
rect 65 152 66 153
rect 64 152 65 153
rect 63 152 64 153
rect 62 152 63 153
rect 61 152 62 153
rect 60 152 61 153
rect 59 152 60 153
rect 58 152 59 153
rect 57 152 58 153
rect 56 152 57 153
rect 55 152 56 153
rect 54 152 55 153
rect 53 152 54 153
rect 52 152 53 153
rect 51 152 52 153
rect 50 152 51 153
rect 49 152 50 153
rect 48 152 49 153
rect 47 152 48 153
rect 46 152 47 153
rect 45 152 46 153
rect 44 152 45 153
rect 43 152 44 153
rect 42 152 43 153
rect 41 152 42 153
rect 40 152 41 153
rect 39 152 40 153
rect 38 152 39 153
rect 37 152 38 153
rect 36 152 37 153
rect 35 152 36 153
rect 26 152 27 153
rect 25 152 26 153
rect 24 152 25 153
rect 23 152 24 153
rect 22 152 23 153
rect 21 152 22 153
rect 20 152 21 153
rect 19 152 20 153
rect 18 152 19 153
rect 17 152 18 153
rect 16 152 17 153
rect 15 152 16 153
rect 14 152 15 153
rect 13 152 14 153
rect 12 152 13 153
rect 11 152 12 153
rect 10 152 11 153
rect 9 152 10 153
rect 8 152 9 153
rect 7 152 8 153
rect 6 152 7 153
rect 437 153 438 154
rect 436 153 437 154
rect 395 153 396 154
rect 394 153 395 154
rect 393 153 394 154
rect 322 153 323 154
rect 321 153 322 154
rect 320 153 321 154
rect 319 153 320 154
rect 318 153 319 154
rect 317 153 318 154
rect 316 153 317 154
rect 315 153 316 154
rect 314 153 315 154
rect 313 153 314 154
rect 312 153 313 154
rect 311 153 312 154
rect 310 153 311 154
rect 309 153 310 154
rect 308 153 309 154
rect 307 153 308 154
rect 306 153 307 154
rect 305 153 306 154
rect 304 153 305 154
rect 303 153 304 154
rect 302 153 303 154
rect 301 153 302 154
rect 300 153 301 154
rect 299 153 300 154
rect 298 153 299 154
rect 297 153 298 154
rect 296 153 297 154
rect 295 153 296 154
rect 294 153 295 154
rect 293 153 294 154
rect 292 153 293 154
rect 291 153 292 154
rect 290 153 291 154
rect 289 153 290 154
rect 288 153 289 154
rect 287 153 288 154
rect 286 153 287 154
rect 285 153 286 154
rect 284 153 285 154
rect 283 153 284 154
rect 282 153 283 154
rect 281 153 282 154
rect 280 153 281 154
rect 279 153 280 154
rect 278 153 279 154
rect 277 153 278 154
rect 276 153 277 154
rect 275 153 276 154
rect 274 153 275 154
rect 273 153 274 154
rect 272 153 273 154
rect 271 153 272 154
rect 270 153 271 154
rect 269 153 270 154
rect 268 153 269 154
rect 267 153 268 154
rect 266 153 267 154
rect 265 153 266 154
rect 264 153 265 154
rect 263 153 264 154
rect 262 153 263 154
rect 261 153 262 154
rect 260 153 261 154
rect 259 153 260 154
rect 258 153 259 154
rect 257 153 258 154
rect 256 153 257 154
rect 255 153 256 154
rect 254 153 255 154
rect 253 153 254 154
rect 252 153 253 154
rect 251 153 252 154
rect 250 153 251 154
rect 249 153 250 154
rect 248 153 249 154
rect 247 153 248 154
rect 246 153 247 154
rect 245 153 246 154
rect 244 153 245 154
rect 243 153 244 154
rect 242 153 243 154
rect 241 153 242 154
rect 240 153 241 154
rect 239 153 240 154
rect 238 153 239 154
rect 237 153 238 154
rect 236 153 237 154
rect 235 153 236 154
rect 234 153 235 154
rect 214 153 215 154
rect 213 153 214 154
rect 212 153 213 154
rect 211 153 212 154
rect 210 153 211 154
rect 209 153 210 154
rect 208 153 209 154
rect 207 153 208 154
rect 206 153 207 154
rect 205 153 206 154
rect 204 153 205 154
rect 203 153 204 154
rect 202 153 203 154
rect 201 153 202 154
rect 200 153 201 154
rect 199 153 200 154
rect 198 153 199 154
rect 197 153 198 154
rect 196 153 197 154
rect 195 153 196 154
rect 194 153 195 154
rect 193 153 194 154
rect 192 153 193 154
rect 191 153 192 154
rect 190 153 191 154
rect 189 153 190 154
rect 188 153 189 154
rect 187 153 188 154
rect 186 153 187 154
rect 185 153 186 154
rect 184 153 185 154
rect 183 153 184 154
rect 182 153 183 154
rect 181 153 182 154
rect 180 153 181 154
rect 179 153 180 154
rect 178 153 179 154
rect 177 153 178 154
rect 176 153 177 154
rect 175 153 176 154
rect 174 153 175 154
rect 173 153 174 154
rect 172 153 173 154
rect 171 153 172 154
rect 170 153 171 154
rect 169 153 170 154
rect 168 153 169 154
rect 167 153 168 154
rect 166 153 167 154
rect 165 153 166 154
rect 164 153 165 154
rect 163 153 164 154
rect 162 153 163 154
rect 161 153 162 154
rect 160 153 161 154
rect 159 153 160 154
rect 158 153 159 154
rect 157 153 158 154
rect 156 153 157 154
rect 155 153 156 154
rect 154 153 155 154
rect 153 153 154 154
rect 152 153 153 154
rect 151 153 152 154
rect 150 153 151 154
rect 149 153 150 154
rect 148 153 149 154
rect 117 153 118 154
rect 116 153 117 154
rect 115 153 116 154
rect 114 153 115 154
rect 113 153 114 154
rect 112 153 113 154
rect 111 153 112 154
rect 110 153 111 154
rect 109 153 110 154
rect 108 153 109 154
rect 107 153 108 154
rect 106 153 107 154
rect 105 153 106 154
rect 104 153 105 154
rect 103 153 104 154
rect 102 153 103 154
rect 101 153 102 154
rect 100 153 101 154
rect 99 153 100 154
rect 98 153 99 154
rect 97 153 98 154
rect 96 153 97 154
rect 95 153 96 154
rect 94 153 95 154
rect 93 153 94 154
rect 92 153 93 154
rect 91 153 92 154
rect 90 153 91 154
rect 89 153 90 154
rect 88 153 89 154
rect 87 153 88 154
rect 86 153 87 154
rect 85 153 86 154
rect 84 153 85 154
rect 83 153 84 154
rect 82 153 83 154
rect 81 153 82 154
rect 80 153 81 154
rect 79 153 80 154
rect 78 153 79 154
rect 77 153 78 154
rect 76 153 77 154
rect 75 153 76 154
rect 74 153 75 154
rect 73 153 74 154
rect 72 153 73 154
rect 71 153 72 154
rect 70 153 71 154
rect 69 153 70 154
rect 68 153 69 154
rect 67 153 68 154
rect 66 153 67 154
rect 65 153 66 154
rect 64 153 65 154
rect 63 153 64 154
rect 62 153 63 154
rect 61 153 62 154
rect 60 153 61 154
rect 59 153 60 154
rect 58 153 59 154
rect 57 153 58 154
rect 56 153 57 154
rect 55 153 56 154
rect 54 153 55 154
rect 53 153 54 154
rect 52 153 53 154
rect 51 153 52 154
rect 50 153 51 154
rect 49 153 50 154
rect 48 153 49 154
rect 47 153 48 154
rect 46 153 47 154
rect 45 153 46 154
rect 44 153 45 154
rect 43 153 44 154
rect 42 153 43 154
rect 41 153 42 154
rect 40 153 41 154
rect 39 153 40 154
rect 38 153 39 154
rect 37 153 38 154
rect 36 153 37 154
rect 35 153 36 154
rect 34 153 35 154
rect 26 153 27 154
rect 25 153 26 154
rect 24 153 25 154
rect 23 153 24 154
rect 22 153 23 154
rect 21 153 22 154
rect 20 153 21 154
rect 19 153 20 154
rect 18 153 19 154
rect 17 153 18 154
rect 16 153 17 154
rect 15 153 16 154
rect 14 153 15 154
rect 13 153 14 154
rect 12 153 13 154
rect 11 153 12 154
rect 10 153 11 154
rect 9 153 10 154
rect 8 153 9 154
rect 7 153 8 154
rect 6 153 7 154
rect 437 154 438 155
rect 436 154 437 155
rect 435 154 436 155
rect 395 154 396 155
rect 394 154 395 155
rect 393 154 394 155
rect 323 154 324 155
rect 322 154 323 155
rect 321 154 322 155
rect 320 154 321 155
rect 319 154 320 155
rect 318 154 319 155
rect 317 154 318 155
rect 316 154 317 155
rect 315 154 316 155
rect 314 154 315 155
rect 313 154 314 155
rect 312 154 313 155
rect 311 154 312 155
rect 310 154 311 155
rect 309 154 310 155
rect 308 154 309 155
rect 307 154 308 155
rect 306 154 307 155
rect 305 154 306 155
rect 304 154 305 155
rect 303 154 304 155
rect 302 154 303 155
rect 301 154 302 155
rect 300 154 301 155
rect 299 154 300 155
rect 298 154 299 155
rect 297 154 298 155
rect 296 154 297 155
rect 295 154 296 155
rect 294 154 295 155
rect 293 154 294 155
rect 292 154 293 155
rect 291 154 292 155
rect 290 154 291 155
rect 289 154 290 155
rect 288 154 289 155
rect 287 154 288 155
rect 286 154 287 155
rect 285 154 286 155
rect 284 154 285 155
rect 283 154 284 155
rect 282 154 283 155
rect 281 154 282 155
rect 280 154 281 155
rect 279 154 280 155
rect 278 154 279 155
rect 277 154 278 155
rect 276 154 277 155
rect 275 154 276 155
rect 274 154 275 155
rect 273 154 274 155
rect 272 154 273 155
rect 271 154 272 155
rect 270 154 271 155
rect 269 154 270 155
rect 268 154 269 155
rect 267 154 268 155
rect 266 154 267 155
rect 265 154 266 155
rect 264 154 265 155
rect 263 154 264 155
rect 262 154 263 155
rect 261 154 262 155
rect 260 154 261 155
rect 259 154 260 155
rect 258 154 259 155
rect 257 154 258 155
rect 256 154 257 155
rect 255 154 256 155
rect 254 154 255 155
rect 253 154 254 155
rect 252 154 253 155
rect 251 154 252 155
rect 250 154 251 155
rect 249 154 250 155
rect 248 154 249 155
rect 247 154 248 155
rect 246 154 247 155
rect 245 154 246 155
rect 244 154 245 155
rect 243 154 244 155
rect 242 154 243 155
rect 241 154 242 155
rect 240 154 241 155
rect 239 154 240 155
rect 238 154 239 155
rect 237 154 238 155
rect 236 154 237 155
rect 235 154 236 155
rect 234 154 235 155
rect 233 154 234 155
rect 214 154 215 155
rect 213 154 214 155
rect 212 154 213 155
rect 211 154 212 155
rect 210 154 211 155
rect 209 154 210 155
rect 208 154 209 155
rect 207 154 208 155
rect 206 154 207 155
rect 205 154 206 155
rect 204 154 205 155
rect 203 154 204 155
rect 202 154 203 155
rect 201 154 202 155
rect 200 154 201 155
rect 199 154 200 155
rect 198 154 199 155
rect 197 154 198 155
rect 196 154 197 155
rect 195 154 196 155
rect 194 154 195 155
rect 193 154 194 155
rect 192 154 193 155
rect 191 154 192 155
rect 190 154 191 155
rect 189 154 190 155
rect 188 154 189 155
rect 187 154 188 155
rect 186 154 187 155
rect 185 154 186 155
rect 184 154 185 155
rect 183 154 184 155
rect 182 154 183 155
rect 181 154 182 155
rect 180 154 181 155
rect 179 154 180 155
rect 178 154 179 155
rect 177 154 178 155
rect 176 154 177 155
rect 175 154 176 155
rect 174 154 175 155
rect 173 154 174 155
rect 172 154 173 155
rect 171 154 172 155
rect 170 154 171 155
rect 169 154 170 155
rect 168 154 169 155
rect 167 154 168 155
rect 166 154 167 155
rect 165 154 166 155
rect 164 154 165 155
rect 163 154 164 155
rect 162 154 163 155
rect 161 154 162 155
rect 160 154 161 155
rect 159 154 160 155
rect 158 154 159 155
rect 157 154 158 155
rect 156 154 157 155
rect 155 154 156 155
rect 154 154 155 155
rect 153 154 154 155
rect 152 154 153 155
rect 151 154 152 155
rect 150 154 151 155
rect 149 154 150 155
rect 148 154 149 155
rect 147 154 148 155
rect 116 154 117 155
rect 115 154 116 155
rect 114 154 115 155
rect 113 154 114 155
rect 112 154 113 155
rect 111 154 112 155
rect 110 154 111 155
rect 109 154 110 155
rect 108 154 109 155
rect 107 154 108 155
rect 106 154 107 155
rect 105 154 106 155
rect 104 154 105 155
rect 103 154 104 155
rect 102 154 103 155
rect 101 154 102 155
rect 100 154 101 155
rect 99 154 100 155
rect 98 154 99 155
rect 97 154 98 155
rect 96 154 97 155
rect 95 154 96 155
rect 94 154 95 155
rect 93 154 94 155
rect 92 154 93 155
rect 91 154 92 155
rect 90 154 91 155
rect 89 154 90 155
rect 88 154 89 155
rect 87 154 88 155
rect 86 154 87 155
rect 85 154 86 155
rect 84 154 85 155
rect 83 154 84 155
rect 82 154 83 155
rect 81 154 82 155
rect 80 154 81 155
rect 79 154 80 155
rect 78 154 79 155
rect 77 154 78 155
rect 76 154 77 155
rect 75 154 76 155
rect 74 154 75 155
rect 73 154 74 155
rect 72 154 73 155
rect 71 154 72 155
rect 70 154 71 155
rect 69 154 70 155
rect 68 154 69 155
rect 67 154 68 155
rect 66 154 67 155
rect 65 154 66 155
rect 64 154 65 155
rect 63 154 64 155
rect 62 154 63 155
rect 61 154 62 155
rect 60 154 61 155
rect 59 154 60 155
rect 58 154 59 155
rect 57 154 58 155
rect 56 154 57 155
rect 55 154 56 155
rect 54 154 55 155
rect 53 154 54 155
rect 52 154 53 155
rect 51 154 52 155
rect 50 154 51 155
rect 49 154 50 155
rect 48 154 49 155
rect 47 154 48 155
rect 46 154 47 155
rect 45 154 46 155
rect 44 154 45 155
rect 43 154 44 155
rect 42 154 43 155
rect 41 154 42 155
rect 40 154 41 155
rect 39 154 40 155
rect 38 154 39 155
rect 37 154 38 155
rect 36 154 37 155
rect 35 154 36 155
rect 34 154 35 155
rect 25 154 26 155
rect 24 154 25 155
rect 23 154 24 155
rect 22 154 23 155
rect 21 154 22 155
rect 20 154 21 155
rect 19 154 20 155
rect 18 154 19 155
rect 17 154 18 155
rect 16 154 17 155
rect 15 154 16 155
rect 14 154 15 155
rect 13 154 14 155
rect 12 154 13 155
rect 11 154 12 155
rect 10 154 11 155
rect 9 154 10 155
rect 8 154 9 155
rect 7 154 8 155
rect 6 154 7 155
rect 437 155 438 156
rect 436 155 437 156
rect 435 155 436 156
rect 395 155 396 156
rect 394 155 395 156
rect 393 155 394 156
rect 324 155 325 156
rect 323 155 324 156
rect 322 155 323 156
rect 321 155 322 156
rect 320 155 321 156
rect 319 155 320 156
rect 318 155 319 156
rect 317 155 318 156
rect 316 155 317 156
rect 315 155 316 156
rect 314 155 315 156
rect 313 155 314 156
rect 312 155 313 156
rect 311 155 312 156
rect 310 155 311 156
rect 309 155 310 156
rect 308 155 309 156
rect 307 155 308 156
rect 306 155 307 156
rect 305 155 306 156
rect 304 155 305 156
rect 303 155 304 156
rect 302 155 303 156
rect 301 155 302 156
rect 300 155 301 156
rect 299 155 300 156
rect 298 155 299 156
rect 297 155 298 156
rect 296 155 297 156
rect 295 155 296 156
rect 294 155 295 156
rect 293 155 294 156
rect 292 155 293 156
rect 291 155 292 156
rect 290 155 291 156
rect 289 155 290 156
rect 288 155 289 156
rect 287 155 288 156
rect 286 155 287 156
rect 285 155 286 156
rect 284 155 285 156
rect 283 155 284 156
rect 282 155 283 156
rect 281 155 282 156
rect 280 155 281 156
rect 279 155 280 156
rect 278 155 279 156
rect 277 155 278 156
rect 276 155 277 156
rect 275 155 276 156
rect 274 155 275 156
rect 273 155 274 156
rect 272 155 273 156
rect 271 155 272 156
rect 270 155 271 156
rect 269 155 270 156
rect 268 155 269 156
rect 267 155 268 156
rect 266 155 267 156
rect 265 155 266 156
rect 264 155 265 156
rect 263 155 264 156
rect 262 155 263 156
rect 261 155 262 156
rect 260 155 261 156
rect 259 155 260 156
rect 258 155 259 156
rect 257 155 258 156
rect 256 155 257 156
rect 255 155 256 156
rect 254 155 255 156
rect 253 155 254 156
rect 252 155 253 156
rect 251 155 252 156
rect 250 155 251 156
rect 249 155 250 156
rect 248 155 249 156
rect 247 155 248 156
rect 246 155 247 156
rect 245 155 246 156
rect 244 155 245 156
rect 243 155 244 156
rect 242 155 243 156
rect 241 155 242 156
rect 240 155 241 156
rect 239 155 240 156
rect 238 155 239 156
rect 237 155 238 156
rect 236 155 237 156
rect 235 155 236 156
rect 234 155 235 156
rect 233 155 234 156
rect 213 155 214 156
rect 212 155 213 156
rect 211 155 212 156
rect 210 155 211 156
rect 209 155 210 156
rect 208 155 209 156
rect 207 155 208 156
rect 206 155 207 156
rect 205 155 206 156
rect 204 155 205 156
rect 203 155 204 156
rect 202 155 203 156
rect 201 155 202 156
rect 200 155 201 156
rect 199 155 200 156
rect 198 155 199 156
rect 197 155 198 156
rect 196 155 197 156
rect 195 155 196 156
rect 194 155 195 156
rect 193 155 194 156
rect 192 155 193 156
rect 191 155 192 156
rect 190 155 191 156
rect 189 155 190 156
rect 188 155 189 156
rect 187 155 188 156
rect 186 155 187 156
rect 185 155 186 156
rect 184 155 185 156
rect 183 155 184 156
rect 182 155 183 156
rect 181 155 182 156
rect 180 155 181 156
rect 179 155 180 156
rect 178 155 179 156
rect 177 155 178 156
rect 176 155 177 156
rect 175 155 176 156
rect 174 155 175 156
rect 173 155 174 156
rect 172 155 173 156
rect 171 155 172 156
rect 170 155 171 156
rect 169 155 170 156
rect 168 155 169 156
rect 167 155 168 156
rect 166 155 167 156
rect 165 155 166 156
rect 164 155 165 156
rect 163 155 164 156
rect 162 155 163 156
rect 161 155 162 156
rect 160 155 161 156
rect 159 155 160 156
rect 158 155 159 156
rect 157 155 158 156
rect 156 155 157 156
rect 155 155 156 156
rect 154 155 155 156
rect 153 155 154 156
rect 152 155 153 156
rect 151 155 152 156
rect 150 155 151 156
rect 149 155 150 156
rect 148 155 149 156
rect 147 155 148 156
rect 146 155 147 156
rect 115 155 116 156
rect 114 155 115 156
rect 113 155 114 156
rect 112 155 113 156
rect 111 155 112 156
rect 110 155 111 156
rect 109 155 110 156
rect 108 155 109 156
rect 107 155 108 156
rect 106 155 107 156
rect 105 155 106 156
rect 104 155 105 156
rect 103 155 104 156
rect 102 155 103 156
rect 101 155 102 156
rect 100 155 101 156
rect 99 155 100 156
rect 98 155 99 156
rect 97 155 98 156
rect 96 155 97 156
rect 95 155 96 156
rect 94 155 95 156
rect 93 155 94 156
rect 92 155 93 156
rect 91 155 92 156
rect 90 155 91 156
rect 89 155 90 156
rect 88 155 89 156
rect 87 155 88 156
rect 86 155 87 156
rect 85 155 86 156
rect 84 155 85 156
rect 83 155 84 156
rect 82 155 83 156
rect 81 155 82 156
rect 80 155 81 156
rect 79 155 80 156
rect 78 155 79 156
rect 77 155 78 156
rect 76 155 77 156
rect 75 155 76 156
rect 74 155 75 156
rect 73 155 74 156
rect 72 155 73 156
rect 71 155 72 156
rect 70 155 71 156
rect 69 155 70 156
rect 68 155 69 156
rect 67 155 68 156
rect 66 155 67 156
rect 65 155 66 156
rect 64 155 65 156
rect 63 155 64 156
rect 62 155 63 156
rect 61 155 62 156
rect 60 155 61 156
rect 59 155 60 156
rect 58 155 59 156
rect 57 155 58 156
rect 56 155 57 156
rect 55 155 56 156
rect 54 155 55 156
rect 53 155 54 156
rect 52 155 53 156
rect 51 155 52 156
rect 50 155 51 156
rect 49 155 50 156
rect 48 155 49 156
rect 47 155 48 156
rect 46 155 47 156
rect 45 155 46 156
rect 44 155 45 156
rect 43 155 44 156
rect 42 155 43 156
rect 41 155 42 156
rect 40 155 41 156
rect 39 155 40 156
rect 38 155 39 156
rect 37 155 38 156
rect 36 155 37 156
rect 35 155 36 156
rect 34 155 35 156
rect 33 155 34 156
rect 25 155 26 156
rect 24 155 25 156
rect 23 155 24 156
rect 22 155 23 156
rect 21 155 22 156
rect 20 155 21 156
rect 19 155 20 156
rect 18 155 19 156
rect 17 155 18 156
rect 16 155 17 156
rect 15 155 16 156
rect 14 155 15 156
rect 13 155 14 156
rect 12 155 13 156
rect 11 155 12 156
rect 10 155 11 156
rect 9 155 10 156
rect 8 155 9 156
rect 7 155 8 156
rect 6 155 7 156
rect 5 155 6 156
rect 437 156 438 157
rect 436 156 437 157
rect 435 156 436 157
rect 396 156 397 157
rect 395 156 396 157
rect 394 156 395 157
rect 393 156 394 157
rect 324 156 325 157
rect 323 156 324 157
rect 322 156 323 157
rect 321 156 322 157
rect 320 156 321 157
rect 319 156 320 157
rect 318 156 319 157
rect 317 156 318 157
rect 316 156 317 157
rect 315 156 316 157
rect 314 156 315 157
rect 313 156 314 157
rect 294 156 295 157
rect 293 156 294 157
rect 292 156 293 157
rect 291 156 292 157
rect 290 156 291 157
rect 289 156 290 157
rect 288 156 289 157
rect 287 156 288 157
rect 286 156 287 157
rect 285 156 286 157
rect 284 156 285 157
rect 283 156 284 157
rect 282 156 283 157
rect 281 156 282 157
rect 280 156 281 157
rect 279 156 280 157
rect 278 156 279 157
rect 277 156 278 157
rect 276 156 277 157
rect 275 156 276 157
rect 274 156 275 157
rect 273 156 274 157
rect 272 156 273 157
rect 271 156 272 157
rect 270 156 271 157
rect 269 156 270 157
rect 268 156 269 157
rect 267 156 268 157
rect 266 156 267 157
rect 265 156 266 157
rect 264 156 265 157
rect 263 156 264 157
rect 262 156 263 157
rect 261 156 262 157
rect 260 156 261 157
rect 259 156 260 157
rect 258 156 259 157
rect 257 156 258 157
rect 256 156 257 157
rect 255 156 256 157
rect 254 156 255 157
rect 253 156 254 157
rect 252 156 253 157
rect 251 156 252 157
rect 250 156 251 157
rect 249 156 250 157
rect 248 156 249 157
rect 247 156 248 157
rect 246 156 247 157
rect 245 156 246 157
rect 244 156 245 157
rect 243 156 244 157
rect 242 156 243 157
rect 241 156 242 157
rect 240 156 241 157
rect 239 156 240 157
rect 238 156 239 157
rect 237 156 238 157
rect 236 156 237 157
rect 235 156 236 157
rect 234 156 235 157
rect 233 156 234 157
rect 232 156 233 157
rect 213 156 214 157
rect 212 156 213 157
rect 211 156 212 157
rect 210 156 211 157
rect 209 156 210 157
rect 208 156 209 157
rect 207 156 208 157
rect 206 156 207 157
rect 205 156 206 157
rect 204 156 205 157
rect 203 156 204 157
rect 202 156 203 157
rect 201 156 202 157
rect 200 156 201 157
rect 199 156 200 157
rect 198 156 199 157
rect 197 156 198 157
rect 196 156 197 157
rect 195 156 196 157
rect 194 156 195 157
rect 193 156 194 157
rect 192 156 193 157
rect 191 156 192 157
rect 190 156 191 157
rect 189 156 190 157
rect 188 156 189 157
rect 187 156 188 157
rect 186 156 187 157
rect 185 156 186 157
rect 184 156 185 157
rect 183 156 184 157
rect 182 156 183 157
rect 181 156 182 157
rect 180 156 181 157
rect 179 156 180 157
rect 178 156 179 157
rect 177 156 178 157
rect 176 156 177 157
rect 175 156 176 157
rect 174 156 175 157
rect 173 156 174 157
rect 172 156 173 157
rect 171 156 172 157
rect 170 156 171 157
rect 169 156 170 157
rect 168 156 169 157
rect 167 156 168 157
rect 166 156 167 157
rect 165 156 166 157
rect 164 156 165 157
rect 163 156 164 157
rect 162 156 163 157
rect 161 156 162 157
rect 160 156 161 157
rect 159 156 160 157
rect 158 156 159 157
rect 157 156 158 157
rect 156 156 157 157
rect 155 156 156 157
rect 154 156 155 157
rect 153 156 154 157
rect 152 156 153 157
rect 151 156 152 157
rect 150 156 151 157
rect 149 156 150 157
rect 148 156 149 157
rect 147 156 148 157
rect 146 156 147 157
rect 145 156 146 157
rect 113 156 114 157
rect 112 156 113 157
rect 111 156 112 157
rect 110 156 111 157
rect 109 156 110 157
rect 108 156 109 157
rect 107 156 108 157
rect 106 156 107 157
rect 105 156 106 157
rect 104 156 105 157
rect 103 156 104 157
rect 102 156 103 157
rect 101 156 102 157
rect 100 156 101 157
rect 99 156 100 157
rect 98 156 99 157
rect 97 156 98 157
rect 96 156 97 157
rect 95 156 96 157
rect 94 156 95 157
rect 93 156 94 157
rect 92 156 93 157
rect 91 156 92 157
rect 90 156 91 157
rect 89 156 90 157
rect 88 156 89 157
rect 87 156 88 157
rect 86 156 87 157
rect 85 156 86 157
rect 84 156 85 157
rect 83 156 84 157
rect 82 156 83 157
rect 81 156 82 157
rect 80 156 81 157
rect 79 156 80 157
rect 78 156 79 157
rect 77 156 78 157
rect 76 156 77 157
rect 75 156 76 157
rect 74 156 75 157
rect 73 156 74 157
rect 72 156 73 157
rect 71 156 72 157
rect 70 156 71 157
rect 69 156 70 157
rect 68 156 69 157
rect 67 156 68 157
rect 66 156 67 157
rect 65 156 66 157
rect 64 156 65 157
rect 63 156 64 157
rect 62 156 63 157
rect 61 156 62 157
rect 60 156 61 157
rect 59 156 60 157
rect 58 156 59 157
rect 57 156 58 157
rect 56 156 57 157
rect 55 156 56 157
rect 54 156 55 157
rect 53 156 54 157
rect 52 156 53 157
rect 51 156 52 157
rect 50 156 51 157
rect 49 156 50 157
rect 48 156 49 157
rect 47 156 48 157
rect 46 156 47 157
rect 45 156 46 157
rect 44 156 45 157
rect 43 156 44 157
rect 42 156 43 157
rect 41 156 42 157
rect 40 156 41 157
rect 39 156 40 157
rect 38 156 39 157
rect 37 156 38 157
rect 36 156 37 157
rect 35 156 36 157
rect 34 156 35 157
rect 33 156 34 157
rect 24 156 25 157
rect 23 156 24 157
rect 22 156 23 157
rect 21 156 22 157
rect 20 156 21 157
rect 19 156 20 157
rect 18 156 19 157
rect 17 156 18 157
rect 16 156 17 157
rect 15 156 16 157
rect 14 156 15 157
rect 13 156 14 157
rect 12 156 13 157
rect 11 156 12 157
rect 10 156 11 157
rect 9 156 10 157
rect 8 156 9 157
rect 7 156 8 157
rect 6 156 7 157
rect 5 156 6 157
rect 437 157 438 158
rect 436 157 437 158
rect 435 157 436 158
rect 434 157 435 158
rect 396 157 397 158
rect 395 157 396 158
rect 394 157 395 158
rect 393 157 394 158
rect 325 157 326 158
rect 324 157 325 158
rect 323 157 324 158
rect 322 157 323 158
rect 321 157 322 158
rect 320 157 321 158
rect 319 157 320 158
rect 290 157 291 158
rect 289 157 290 158
rect 288 157 289 158
rect 287 157 288 158
rect 286 157 287 158
rect 285 157 286 158
rect 284 157 285 158
rect 283 157 284 158
rect 282 157 283 158
rect 281 157 282 158
rect 280 157 281 158
rect 279 157 280 158
rect 278 157 279 158
rect 277 157 278 158
rect 276 157 277 158
rect 275 157 276 158
rect 274 157 275 158
rect 273 157 274 158
rect 272 157 273 158
rect 271 157 272 158
rect 270 157 271 158
rect 269 157 270 158
rect 268 157 269 158
rect 267 157 268 158
rect 266 157 267 158
rect 265 157 266 158
rect 264 157 265 158
rect 263 157 264 158
rect 262 157 263 158
rect 261 157 262 158
rect 260 157 261 158
rect 259 157 260 158
rect 258 157 259 158
rect 257 157 258 158
rect 256 157 257 158
rect 255 157 256 158
rect 254 157 255 158
rect 253 157 254 158
rect 252 157 253 158
rect 251 157 252 158
rect 250 157 251 158
rect 249 157 250 158
rect 248 157 249 158
rect 247 157 248 158
rect 246 157 247 158
rect 245 157 246 158
rect 244 157 245 158
rect 243 157 244 158
rect 242 157 243 158
rect 241 157 242 158
rect 240 157 241 158
rect 239 157 240 158
rect 238 157 239 158
rect 237 157 238 158
rect 236 157 237 158
rect 235 157 236 158
rect 234 157 235 158
rect 233 157 234 158
rect 232 157 233 158
rect 231 157 232 158
rect 212 157 213 158
rect 211 157 212 158
rect 210 157 211 158
rect 209 157 210 158
rect 208 157 209 158
rect 207 157 208 158
rect 206 157 207 158
rect 205 157 206 158
rect 204 157 205 158
rect 203 157 204 158
rect 202 157 203 158
rect 201 157 202 158
rect 200 157 201 158
rect 199 157 200 158
rect 198 157 199 158
rect 197 157 198 158
rect 196 157 197 158
rect 195 157 196 158
rect 194 157 195 158
rect 193 157 194 158
rect 192 157 193 158
rect 191 157 192 158
rect 190 157 191 158
rect 189 157 190 158
rect 188 157 189 158
rect 187 157 188 158
rect 186 157 187 158
rect 185 157 186 158
rect 184 157 185 158
rect 183 157 184 158
rect 182 157 183 158
rect 181 157 182 158
rect 180 157 181 158
rect 179 157 180 158
rect 178 157 179 158
rect 177 157 178 158
rect 176 157 177 158
rect 175 157 176 158
rect 174 157 175 158
rect 173 157 174 158
rect 172 157 173 158
rect 171 157 172 158
rect 170 157 171 158
rect 169 157 170 158
rect 168 157 169 158
rect 167 157 168 158
rect 166 157 167 158
rect 165 157 166 158
rect 164 157 165 158
rect 163 157 164 158
rect 162 157 163 158
rect 161 157 162 158
rect 160 157 161 158
rect 159 157 160 158
rect 158 157 159 158
rect 157 157 158 158
rect 156 157 157 158
rect 155 157 156 158
rect 154 157 155 158
rect 153 157 154 158
rect 152 157 153 158
rect 151 157 152 158
rect 150 157 151 158
rect 149 157 150 158
rect 148 157 149 158
rect 147 157 148 158
rect 146 157 147 158
rect 145 157 146 158
rect 112 157 113 158
rect 111 157 112 158
rect 110 157 111 158
rect 109 157 110 158
rect 108 157 109 158
rect 107 157 108 158
rect 106 157 107 158
rect 105 157 106 158
rect 104 157 105 158
rect 103 157 104 158
rect 102 157 103 158
rect 101 157 102 158
rect 100 157 101 158
rect 99 157 100 158
rect 98 157 99 158
rect 97 157 98 158
rect 96 157 97 158
rect 95 157 96 158
rect 94 157 95 158
rect 93 157 94 158
rect 92 157 93 158
rect 91 157 92 158
rect 90 157 91 158
rect 89 157 90 158
rect 88 157 89 158
rect 87 157 88 158
rect 86 157 87 158
rect 85 157 86 158
rect 84 157 85 158
rect 83 157 84 158
rect 82 157 83 158
rect 81 157 82 158
rect 80 157 81 158
rect 79 157 80 158
rect 78 157 79 158
rect 77 157 78 158
rect 76 157 77 158
rect 75 157 76 158
rect 74 157 75 158
rect 73 157 74 158
rect 72 157 73 158
rect 71 157 72 158
rect 70 157 71 158
rect 69 157 70 158
rect 68 157 69 158
rect 67 157 68 158
rect 66 157 67 158
rect 65 157 66 158
rect 64 157 65 158
rect 63 157 64 158
rect 62 157 63 158
rect 61 157 62 158
rect 60 157 61 158
rect 59 157 60 158
rect 58 157 59 158
rect 57 157 58 158
rect 56 157 57 158
rect 55 157 56 158
rect 54 157 55 158
rect 53 157 54 158
rect 52 157 53 158
rect 51 157 52 158
rect 50 157 51 158
rect 49 157 50 158
rect 48 157 49 158
rect 47 157 48 158
rect 46 157 47 158
rect 45 157 46 158
rect 44 157 45 158
rect 43 157 44 158
rect 42 157 43 158
rect 41 157 42 158
rect 40 157 41 158
rect 39 157 40 158
rect 38 157 39 158
rect 37 157 38 158
rect 36 157 37 158
rect 35 157 36 158
rect 34 157 35 158
rect 33 157 34 158
rect 32 157 33 158
rect 23 157 24 158
rect 22 157 23 158
rect 21 157 22 158
rect 20 157 21 158
rect 19 157 20 158
rect 18 157 19 158
rect 17 157 18 158
rect 16 157 17 158
rect 15 157 16 158
rect 14 157 15 158
rect 13 157 14 158
rect 12 157 13 158
rect 11 157 12 158
rect 10 157 11 158
rect 9 157 10 158
rect 8 157 9 158
rect 7 157 8 158
rect 6 157 7 158
rect 5 157 6 158
rect 458 158 459 159
rect 437 158 438 159
rect 436 158 437 159
rect 435 158 436 159
rect 434 158 435 159
rect 433 158 434 159
rect 432 158 433 159
rect 398 158 399 159
rect 397 158 398 159
rect 396 158 397 159
rect 395 158 396 159
rect 394 158 395 159
rect 393 158 394 159
rect 326 158 327 159
rect 325 158 326 159
rect 324 158 325 159
rect 323 158 324 159
rect 287 158 288 159
rect 286 158 287 159
rect 285 158 286 159
rect 284 158 285 159
rect 283 158 284 159
rect 282 158 283 159
rect 281 158 282 159
rect 280 158 281 159
rect 279 158 280 159
rect 278 158 279 159
rect 277 158 278 159
rect 276 158 277 159
rect 275 158 276 159
rect 274 158 275 159
rect 273 158 274 159
rect 272 158 273 159
rect 271 158 272 159
rect 270 158 271 159
rect 269 158 270 159
rect 268 158 269 159
rect 267 158 268 159
rect 266 158 267 159
rect 265 158 266 159
rect 264 158 265 159
rect 263 158 264 159
rect 262 158 263 159
rect 261 158 262 159
rect 260 158 261 159
rect 259 158 260 159
rect 258 158 259 159
rect 257 158 258 159
rect 256 158 257 159
rect 255 158 256 159
rect 254 158 255 159
rect 253 158 254 159
rect 252 158 253 159
rect 251 158 252 159
rect 250 158 251 159
rect 249 158 250 159
rect 248 158 249 159
rect 247 158 248 159
rect 246 158 247 159
rect 245 158 246 159
rect 244 158 245 159
rect 243 158 244 159
rect 242 158 243 159
rect 241 158 242 159
rect 240 158 241 159
rect 239 158 240 159
rect 238 158 239 159
rect 237 158 238 159
rect 236 158 237 159
rect 235 158 236 159
rect 234 158 235 159
rect 233 158 234 159
rect 232 158 233 159
rect 231 158 232 159
rect 212 158 213 159
rect 211 158 212 159
rect 210 158 211 159
rect 209 158 210 159
rect 208 158 209 159
rect 207 158 208 159
rect 206 158 207 159
rect 205 158 206 159
rect 204 158 205 159
rect 203 158 204 159
rect 202 158 203 159
rect 201 158 202 159
rect 200 158 201 159
rect 199 158 200 159
rect 198 158 199 159
rect 197 158 198 159
rect 196 158 197 159
rect 195 158 196 159
rect 194 158 195 159
rect 193 158 194 159
rect 192 158 193 159
rect 191 158 192 159
rect 190 158 191 159
rect 189 158 190 159
rect 188 158 189 159
rect 187 158 188 159
rect 186 158 187 159
rect 185 158 186 159
rect 184 158 185 159
rect 183 158 184 159
rect 182 158 183 159
rect 181 158 182 159
rect 180 158 181 159
rect 179 158 180 159
rect 178 158 179 159
rect 177 158 178 159
rect 176 158 177 159
rect 175 158 176 159
rect 174 158 175 159
rect 173 158 174 159
rect 172 158 173 159
rect 171 158 172 159
rect 170 158 171 159
rect 169 158 170 159
rect 168 158 169 159
rect 167 158 168 159
rect 166 158 167 159
rect 165 158 166 159
rect 164 158 165 159
rect 163 158 164 159
rect 162 158 163 159
rect 161 158 162 159
rect 160 158 161 159
rect 159 158 160 159
rect 158 158 159 159
rect 157 158 158 159
rect 156 158 157 159
rect 155 158 156 159
rect 154 158 155 159
rect 153 158 154 159
rect 152 158 153 159
rect 151 158 152 159
rect 150 158 151 159
rect 149 158 150 159
rect 148 158 149 159
rect 147 158 148 159
rect 146 158 147 159
rect 145 158 146 159
rect 144 158 145 159
rect 110 158 111 159
rect 109 158 110 159
rect 108 158 109 159
rect 107 158 108 159
rect 106 158 107 159
rect 105 158 106 159
rect 104 158 105 159
rect 103 158 104 159
rect 102 158 103 159
rect 101 158 102 159
rect 100 158 101 159
rect 99 158 100 159
rect 98 158 99 159
rect 97 158 98 159
rect 96 158 97 159
rect 95 158 96 159
rect 94 158 95 159
rect 93 158 94 159
rect 92 158 93 159
rect 91 158 92 159
rect 90 158 91 159
rect 89 158 90 159
rect 88 158 89 159
rect 87 158 88 159
rect 86 158 87 159
rect 85 158 86 159
rect 84 158 85 159
rect 83 158 84 159
rect 82 158 83 159
rect 81 158 82 159
rect 80 158 81 159
rect 79 158 80 159
rect 78 158 79 159
rect 77 158 78 159
rect 76 158 77 159
rect 75 158 76 159
rect 74 158 75 159
rect 73 158 74 159
rect 72 158 73 159
rect 71 158 72 159
rect 70 158 71 159
rect 69 158 70 159
rect 68 158 69 159
rect 67 158 68 159
rect 66 158 67 159
rect 65 158 66 159
rect 64 158 65 159
rect 63 158 64 159
rect 62 158 63 159
rect 61 158 62 159
rect 60 158 61 159
rect 59 158 60 159
rect 58 158 59 159
rect 57 158 58 159
rect 56 158 57 159
rect 55 158 56 159
rect 54 158 55 159
rect 53 158 54 159
rect 52 158 53 159
rect 51 158 52 159
rect 50 158 51 159
rect 49 158 50 159
rect 48 158 49 159
rect 47 158 48 159
rect 46 158 47 159
rect 45 158 46 159
rect 44 158 45 159
rect 43 158 44 159
rect 42 158 43 159
rect 41 158 42 159
rect 40 158 41 159
rect 39 158 40 159
rect 38 158 39 159
rect 37 158 38 159
rect 36 158 37 159
rect 35 158 36 159
rect 34 158 35 159
rect 33 158 34 159
rect 32 158 33 159
rect 23 158 24 159
rect 22 158 23 159
rect 21 158 22 159
rect 20 158 21 159
rect 19 158 20 159
rect 18 158 19 159
rect 17 158 18 159
rect 16 158 17 159
rect 15 158 16 159
rect 14 158 15 159
rect 13 158 14 159
rect 12 158 13 159
rect 11 158 12 159
rect 10 158 11 159
rect 9 158 10 159
rect 8 158 9 159
rect 7 158 8 159
rect 6 158 7 159
rect 5 158 6 159
rect 458 159 459 160
rect 437 159 438 160
rect 436 159 437 160
rect 435 159 436 160
rect 434 159 435 160
rect 433 159 434 160
rect 432 159 433 160
rect 431 159 432 160
rect 430 159 431 160
rect 429 159 430 160
rect 428 159 429 160
rect 427 159 428 160
rect 426 159 427 160
rect 425 159 426 160
rect 424 159 425 160
rect 423 159 424 160
rect 422 159 423 160
rect 421 159 422 160
rect 420 159 421 160
rect 419 159 420 160
rect 418 159 419 160
rect 417 159 418 160
rect 416 159 417 160
rect 415 159 416 160
rect 414 159 415 160
rect 413 159 414 160
rect 412 159 413 160
rect 411 159 412 160
rect 410 159 411 160
rect 409 159 410 160
rect 408 159 409 160
rect 407 159 408 160
rect 406 159 407 160
rect 405 159 406 160
rect 404 159 405 160
rect 403 159 404 160
rect 402 159 403 160
rect 401 159 402 160
rect 400 159 401 160
rect 399 159 400 160
rect 398 159 399 160
rect 397 159 398 160
rect 396 159 397 160
rect 395 159 396 160
rect 394 159 395 160
rect 393 159 394 160
rect 284 159 285 160
rect 283 159 284 160
rect 282 159 283 160
rect 281 159 282 160
rect 280 159 281 160
rect 279 159 280 160
rect 278 159 279 160
rect 277 159 278 160
rect 276 159 277 160
rect 275 159 276 160
rect 274 159 275 160
rect 273 159 274 160
rect 272 159 273 160
rect 271 159 272 160
rect 270 159 271 160
rect 269 159 270 160
rect 268 159 269 160
rect 267 159 268 160
rect 266 159 267 160
rect 265 159 266 160
rect 264 159 265 160
rect 263 159 264 160
rect 262 159 263 160
rect 261 159 262 160
rect 260 159 261 160
rect 259 159 260 160
rect 258 159 259 160
rect 257 159 258 160
rect 256 159 257 160
rect 255 159 256 160
rect 254 159 255 160
rect 253 159 254 160
rect 252 159 253 160
rect 251 159 252 160
rect 250 159 251 160
rect 249 159 250 160
rect 248 159 249 160
rect 247 159 248 160
rect 246 159 247 160
rect 245 159 246 160
rect 244 159 245 160
rect 243 159 244 160
rect 242 159 243 160
rect 241 159 242 160
rect 240 159 241 160
rect 239 159 240 160
rect 238 159 239 160
rect 237 159 238 160
rect 236 159 237 160
rect 235 159 236 160
rect 234 159 235 160
rect 233 159 234 160
rect 232 159 233 160
rect 231 159 232 160
rect 230 159 231 160
rect 211 159 212 160
rect 210 159 211 160
rect 209 159 210 160
rect 208 159 209 160
rect 207 159 208 160
rect 206 159 207 160
rect 205 159 206 160
rect 204 159 205 160
rect 203 159 204 160
rect 202 159 203 160
rect 201 159 202 160
rect 200 159 201 160
rect 199 159 200 160
rect 198 159 199 160
rect 197 159 198 160
rect 196 159 197 160
rect 195 159 196 160
rect 194 159 195 160
rect 193 159 194 160
rect 192 159 193 160
rect 191 159 192 160
rect 190 159 191 160
rect 189 159 190 160
rect 188 159 189 160
rect 187 159 188 160
rect 186 159 187 160
rect 185 159 186 160
rect 184 159 185 160
rect 183 159 184 160
rect 182 159 183 160
rect 181 159 182 160
rect 180 159 181 160
rect 179 159 180 160
rect 178 159 179 160
rect 177 159 178 160
rect 176 159 177 160
rect 175 159 176 160
rect 174 159 175 160
rect 173 159 174 160
rect 172 159 173 160
rect 171 159 172 160
rect 170 159 171 160
rect 169 159 170 160
rect 168 159 169 160
rect 167 159 168 160
rect 166 159 167 160
rect 165 159 166 160
rect 164 159 165 160
rect 163 159 164 160
rect 162 159 163 160
rect 161 159 162 160
rect 160 159 161 160
rect 159 159 160 160
rect 158 159 159 160
rect 157 159 158 160
rect 156 159 157 160
rect 155 159 156 160
rect 154 159 155 160
rect 153 159 154 160
rect 152 159 153 160
rect 151 159 152 160
rect 150 159 151 160
rect 149 159 150 160
rect 148 159 149 160
rect 147 159 148 160
rect 146 159 147 160
rect 145 159 146 160
rect 144 159 145 160
rect 143 159 144 160
rect 109 159 110 160
rect 108 159 109 160
rect 107 159 108 160
rect 106 159 107 160
rect 105 159 106 160
rect 104 159 105 160
rect 103 159 104 160
rect 102 159 103 160
rect 101 159 102 160
rect 100 159 101 160
rect 99 159 100 160
rect 98 159 99 160
rect 97 159 98 160
rect 96 159 97 160
rect 95 159 96 160
rect 94 159 95 160
rect 93 159 94 160
rect 92 159 93 160
rect 91 159 92 160
rect 90 159 91 160
rect 89 159 90 160
rect 88 159 89 160
rect 87 159 88 160
rect 86 159 87 160
rect 85 159 86 160
rect 84 159 85 160
rect 83 159 84 160
rect 82 159 83 160
rect 81 159 82 160
rect 80 159 81 160
rect 79 159 80 160
rect 78 159 79 160
rect 77 159 78 160
rect 76 159 77 160
rect 75 159 76 160
rect 74 159 75 160
rect 73 159 74 160
rect 72 159 73 160
rect 71 159 72 160
rect 70 159 71 160
rect 69 159 70 160
rect 68 159 69 160
rect 67 159 68 160
rect 66 159 67 160
rect 65 159 66 160
rect 64 159 65 160
rect 63 159 64 160
rect 62 159 63 160
rect 61 159 62 160
rect 60 159 61 160
rect 59 159 60 160
rect 58 159 59 160
rect 57 159 58 160
rect 56 159 57 160
rect 55 159 56 160
rect 54 159 55 160
rect 53 159 54 160
rect 52 159 53 160
rect 51 159 52 160
rect 50 159 51 160
rect 49 159 50 160
rect 48 159 49 160
rect 47 159 48 160
rect 46 159 47 160
rect 45 159 46 160
rect 44 159 45 160
rect 43 159 44 160
rect 42 159 43 160
rect 41 159 42 160
rect 40 159 41 160
rect 39 159 40 160
rect 38 159 39 160
rect 37 159 38 160
rect 36 159 37 160
rect 35 159 36 160
rect 34 159 35 160
rect 33 159 34 160
rect 32 159 33 160
rect 22 159 23 160
rect 21 159 22 160
rect 20 159 21 160
rect 19 159 20 160
rect 18 159 19 160
rect 17 159 18 160
rect 16 159 17 160
rect 15 159 16 160
rect 14 159 15 160
rect 13 159 14 160
rect 12 159 13 160
rect 11 159 12 160
rect 10 159 11 160
rect 9 159 10 160
rect 8 159 9 160
rect 7 159 8 160
rect 6 159 7 160
rect 459 160 460 161
rect 458 160 459 161
rect 437 160 438 161
rect 436 160 437 161
rect 435 160 436 161
rect 434 160 435 161
rect 433 160 434 161
rect 432 160 433 161
rect 431 160 432 161
rect 430 160 431 161
rect 429 160 430 161
rect 428 160 429 161
rect 427 160 428 161
rect 426 160 427 161
rect 425 160 426 161
rect 424 160 425 161
rect 423 160 424 161
rect 422 160 423 161
rect 421 160 422 161
rect 420 160 421 161
rect 419 160 420 161
rect 418 160 419 161
rect 417 160 418 161
rect 416 160 417 161
rect 415 160 416 161
rect 414 160 415 161
rect 413 160 414 161
rect 412 160 413 161
rect 411 160 412 161
rect 410 160 411 161
rect 409 160 410 161
rect 408 160 409 161
rect 407 160 408 161
rect 406 160 407 161
rect 405 160 406 161
rect 404 160 405 161
rect 403 160 404 161
rect 402 160 403 161
rect 401 160 402 161
rect 400 160 401 161
rect 399 160 400 161
rect 398 160 399 161
rect 397 160 398 161
rect 396 160 397 161
rect 395 160 396 161
rect 394 160 395 161
rect 393 160 394 161
rect 282 160 283 161
rect 281 160 282 161
rect 280 160 281 161
rect 279 160 280 161
rect 278 160 279 161
rect 277 160 278 161
rect 276 160 277 161
rect 275 160 276 161
rect 274 160 275 161
rect 273 160 274 161
rect 272 160 273 161
rect 271 160 272 161
rect 270 160 271 161
rect 269 160 270 161
rect 268 160 269 161
rect 267 160 268 161
rect 266 160 267 161
rect 265 160 266 161
rect 264 160 265 161
rect 263 160 264 161
rect 262 160 263 161
rect 261 160 262 161
rect 260 160 261 161
rect 259 160 260 161
rect 258 160 259 161
rect 257 160 258 161
rect 256 160 257 161
rect 255 160 256 161
rect 254 160 255 161
rect 253 160 254 161
rect 252 160 253 161
rect 251 160 252 161
rect 250 160 251 161
rect 249 160 250 161
rect 248 160 249 161
rect 247 160 248 161
rect 246 160 247 161
rect 245 160 246 161
rect 244 160 245 161
rect 243 160 244 161
rect 242 160 243 161
rect 241 160 242 161
rect 240 160 241 161
rect 239 160 240 161
rect 238 160 239 161
rect 237 160 238 161
rect 236 160 237 161
rect 235 160 236 161
rect 234 160 235 161
rect 233 160 234 161
rect 232 160 233 161
rect 231 160 232 161
rect 230 160 231 161
rect 211 160 212 161
rect 210 160 211 161
rect 209 160 210 161
rect 208 160 209 161
rect 207 160 208 161
rect 206 160 207 161
rect 205 160 206 161
rect 204 160 205 161
rect 203 160 204 161
rect 202 160 203 161
rect 201 160 202 161
rect 200 160 201 161
rect 199 160 200 161
rect 198 160 199 161
rect 197 160 198 161
rect 196 160 197 161
rect 195 160 196 161
rect 194 160 195 161
rect 193 160 194 161
rect 192 160 193 161
rect 191 160 192 161
rect 190 160 191 161
rect 189 160 190 161
rect 188 160 189 161
rect 187 160 188 161
rect 186 160 187 161
rect 185 160 186 161
rect 184 160 185 161
rect 183 160 184 161
rect 182 160 183 161
rect 181 160 182 161
rect 180 160 181 161
rect 179 160 180 161
rect 178 160 179 161
rect 177 160 178 161
rect 176 160 177 161
rect 175 160 176 161
rect 174 160 175 161
rect 173 160 174 161
rect 172 160 173 161
rect 171 160 172 161
rect 170 160 171 161
rect 169 160 170 161
rect 168 160 169 161
rect 167 160 168 161
rect 166 160 167 161
rect 165 160 166 161
rect 164 160 165 161
rect 163 160 164 161
rect 162 160 163 161
rect 161 160 162 161
rect 160 160 161 161
rect 159 160 160 161
rect 158 160 159 161
rect 157 160 158 161
rect 156 160 157 161
rect 155 160 156 161
rect 154 160 155 161
rect 153 160 154 161
rect 152 160 153 161
rect 151 160 152 161
rect 150 160 151 161
rect 149 160 150 161
rect 148 160 149 161
rect 147 160 148 161
rect 146 160 147 161
rect 145 160 146 161
rect 144 160 145 161
rect 143 160 144 161
rect 142 160 143 161
rect 141 160 142 161
rect 107 160 108 161
rect 106 160 107 161
rect 105 160 106 161
rect 104 160 105 161
rect 103 160 104 161
rect 102 160 103 161
rect 101 160 102 161
rect 100 160 101 161
rect 99 160 100 161
rect 98 160 99 161
rect 97 160 98 161
rect 96 160 97 161
rect 95 160 96 161
rect 94 160 95 161
rect 93 160 94 161
rect 92 160 93 161
rect 91 160 92 161
rect 90 160 91 161
rect 89 160 90 161
rect 88 160 89 161
rect 87 160 88 161
rect 86 160 87 161
rect 85 160 86 161
rect 84 160 85 161
rect 83 160 84 161
rect 82 160 83 161
rect 81 160 82 161
rect 80 160 81 161
rect 79 160 80 161
rect 78 160 79 161
rect 77 160 78 161
rect 76 160 77 161
rect 75 160 76 161
rect 74 160 75 161
rect 73 160 74 161
rect 72 160 73 161
rect 71 160 72 161
rect 70 160 71 161
rect 69 160 70 161
rect 68 160 69 161
rect 67 160 68 161
rect 66 160 67 161
rect 65 160 66 161
rect 64 160 65 161
rect 63 160 64 161
rect 62 160 63 161
rect 61 160 62 161
rect 60 160 61 161
rect 59 160 60 161
rect 58 160 59 161
rect 57 160 58 161
rect 56 160 57 161
rect 55 160 56 161
rect 54 160 55 161
rect 53 160 54 161
rect 52 160 53 161
rect 51 160 52 161
rect 50 160 51 161
rect 49 160 50 161
rect 48 160 49 161
rect 47 160 48 161
rect 46 160 47 161
rect 45 160 46 161
rect 44 160 45 161
rect 43 160 44 161
rect 42 160 43 161
rect 41 160 42 161
rect 40 160 41 161
rect 39 160 40 161
rect 38 160 39 161
rect 37 160 38 161
rect 36 160 37 161
rect 35 160 36 161
rect 34 160 35 161
rect 33 160 34 161
rect 32 160 33 161
rect 22 160 23 161
rect 21 160 22 161
rect 20 160 21 161
rect 19 160 20 161
rect 18 160 19 161
rect 17 160 18 161
rect 16 160 17 161
rect 15 160 16 161
rect 14 160 15 161
rect 13 160 14 161
rect 12 160 13 161
rect 11 160 12 161
rect 10 160 11 161
rect 9 160 10 161
rect 8 160 9 161
rect 7 160 8 161
rect 6 160 7 161
rect 461 161 462 162
rect 460 161 461 162
rect 459 161 460 162
rect 458 161 459 162
rect 437 161 438 162
rect 436 161 437 162
rect 435 161 436 162
rect 434 161 435 162
rect 433 161 434 162
rect 432 161 433 162
rect 431 161 432 162
rect 430 161 431 162
rect 429 161 430 162
rect 428 161 429 162
rect 427 161 428 162
rect 426 161 427 162
rect 425 161 426 162
rect 424 161 425 162
rect 423 161 424 162
rect 422 161 423 162
rect 421 161 422 162
rect 420 161 421 162
rect 419 161 420 162
rect 418 161 419 162
rect 417 161 418 162
rect 416 161 417 162
rect 415 161 416 162
rect 414 161 415 162
rect 413 161 414 162
rect 412 161 413 162
rect 411 161 412 162
rect 410 161 411 162
rect 409 161 410 162
rect 408 161 409 162
rect 407 161 408 162
rect 406 161 407 162
rect 405 161 406 162
rect 404 161 405 162
rect 403 161 404 162
rect 402 161 403 162
rect 401 161 402 162
rect 400 161 401 162
rect 399 161 400 162
rect 398 161 399 162
rect 397 161 398 162
rect 396 161 397 162
rect 395 161 396 162
rect 394 161 395 162
rect 393 161 394 162
rect 280 161 281 162
rect 279 161 280 162
rect 278 161 279 162
rect 277 161 278 162
rect 276 161 277 162
rect 275 161 276 162
rect 274 161 275 162
rect 273 161 274 162
rect 272 161 273 162
rect 271 161 272 162
rect 270 161 271 162
rect 269 161 270 162
rect 268 161 269 162
rect 267 161 268 162
rect 266 161 267 162
rect 265 161 266 162
rect 264 161 265 162
rect 263 161 264 162
rect 262 161 263 162
rect 261 161 262 162
rect 260 161 261 162
rect 259 161 260 162
rect 258 161 259 162
rect 257 161 258 162
rect 256 161 257 162
rect 255 161 256 162
rect 254 161 255 162
rect 253 161 254 162
rect 252 161 253 162
rect 251 161 252 162
rect 250 161 251 162
rect 249 161 250 162
rect 248 161 249 162
rect 247 161 248 162
rect 246 161 247 162
rect 245 161 246 162
rect 244 161 245 162
rect 243 161 244 162
rect 242 161 243 162
rect 241 161 242 162
rect 240 161 241 162
rect 239 161 240 162
rect 238 161 239 162
rect 237 161 238 162
rect 236 161 237 162
rect 235 161 236 162
rect 234 161 235 162
rect 233 161 234 162
rect 232 161 233 162
rect 231 161 232 162
rect 230 161 231 162
rect 229 161 230 162
rect 211 161 212 162
rect 210 161 211 162
rect 209 161 210 162
rect 208 161 209 162
rect 207 161 208 162
rect 206 161 207 162
rect 205 161 206 162
rect 204 161 205 162
rect 203 161 204 162
rect 202 161 203 162
rect 201 161 202 162
rect 200 161 201 162
rect 199 161 200 162
rect 198 161 199 162
rect 197 161 198 162
rect 196 161 197 162
rect 195 161 196 162
rect 194 161 195 162
rect 193 161 194 162
rect 192 161 193 162
rect 191 161 192 162
rect 190 161 191 162
rect 189 161 190 162
rect 188 161 189 162
rect 187 161 188 162
rect 186 161 187 162
rect 185 161 186 162
rect 184 161 185 162
rect 183 161 184 162
rect 182 161 183 162
rect 181 161 182 162
rect 180 161 181 162
rect 179 161 180 162
rect 178 161 179 162
rect 177 161 178 162
rect 176 161 177 162
rect 175 161 176 162
rect 174 161 175 162
rect 173 161 174 162
rect 172 161 173 162
rect 171 161 172 162
rect 170 161 171 162
rect 169 161 170 162
rect 168 161 169 162
rect 167 161 168 162
rect 166 161 167 162
rect 165 161 166 162
rect 164 161 165 162
rect 163 161 164 162
rect 162 161 163 162
rect 161 161 162 162
rect 160 161 161 162
rect 159 161 160 162
rect 158 161 159 162
rect 157 161 158 162
rect 156 161 157 162
rect 155 161 156 162
rect 154 161 155 162
rect 153 161 154 162
rect 152 161 153 162
rect 151 161 152 162
rect 150 161 151 162
rect 149 161 150 162
rect 148 161 149 162
rect 147 161 148 162
rect 146 161 147 162
rect 145 161 146 162
rect 144 161 145 162
rect 143 161 144 162
rect 142 161 143 162
rect 141 161 142 162
rect 140 161 141 162
rect 106 161 107 162
rect 105 161 106 162
rect 104 161 105 162
rect 103 161 104 162
rect 102 161 103 162
rect 101 161 102 162
rect 100 161 101 162
rect 99 161 100 162
rect 98 161 99 162
rect 97 161 98 162
rect 96 161 97 162
rect 95 161 96 162
rect 94 161 95 162
rect 93 161 94 162
rect 92 161 93 162
rect 91 161 92 162
rect 90 161 91 162
rect 89 161 90 162
rect 88 161 89 162
rect 87 161 88 162
rect 86 161 87 162
rect 85 161 86 162
rect 84 161 85 162
rect 83 161 84 162
rect 82 161 83 162
rect 81 161 82 162
rect 80 161 81 162
rect 79 161 80 162
rect 78 161 79 162
rect 77 161 78 162
rect 76 161 77 162
rect 75 161 76 162
rect 74 161 75 162
rect 73 161 74 162
rect 72 161 73 162
rect 71 161 72 162
rect 70 161 71 162
rect 69 161 70 162
rect 68 161 69 162
rect 67 161 68 162
rect 66 161 67 162
rect 65 161 66 162
rect 64 161 65 162
rect 63 161 64 162
rect 62 161 63 162
rect 61 161 62 162
rect 60 161 61 162
rect 59 161 60 162
rect 58 161 59 162
rect 57 161 58 162
rect 56 161 57 162
rect 55 161 56 162
rect 54 161 55 162
rect 53 161 54 162
rect 52 161 53 162
rect 51 161 52 162
rect 50 161 51 162
rect 49 161 50 162
rect 48 161 49 162
rect 47 161 48 162
rect 46 161 47 162
rect 45 161 46 162
rect 44 161 45 162
rect 43 161 44 162
rect 42 161 43 162
rect 41 161 42 162
rect 40 161 41 162
rect 39 161 40 162
rect 38 161 39 162
rect 37 161 38 162
rect 36 161 37 162
rect 35 161 36 162
rect 34 161 35 162
rect 33 161 34 162
rect 32 161 33 162
rect 31 161 32 162
rect 22 161 23 162
rect 21 161 22 162
rect 20 161 21 162
rect 19 161 20 162
rect 18 161 19 162
rect 17 161 18 162
rect 16 161 17 162
rect 15 161 16 162
rect 14 161 15 162
rect 13 161 14 162
rect 12 161 13 162
rect 11 161 12 162
rect 10 161 11 162
rect 9 161 10 162
rect 8 161 9 162
rect 7 161 8 162
rect 6 161 7 162
rect 463 162 464 163
rect 462 162 463 163
rect 461 162 462 163
rect 460 162 461 163
rect 459 162 460 163
rect 458 162 459 163
rect 437 162 438 163
rect 436 162 437 163
rect 435 162 436 163
rect 434 162 435 163
rect 433 162 434 163
rect 432 162 433 163
rect 431 162 432 163
rect 430 162 431 163
rect 429 162 430 163
rect 428 162 429 163
rect 427 162 428 163
rect 426 162 427 163
rect 425 162 426 163
rect 424 162 425 163
rect 423 162 424 163
rect 422 162 423 163
rect 421 162 422 163
rect 420 162 421 163
rect 419 162 420 163
rect 418 162 419 163
rect 417 162 418 163
rect 416 162 417 163
rect 415 162 416 163
rect 414 162 415 163
rect 413 162 414 163
rect 412 162 413 163
rect 411 162 412 163
rect 410 162 411 163
rect 409 162 410 163
rect 408 162 409 163
rect 407 162 408 163
rect 406 162 407 163
rect 405 162 406 163
rect 404 162 405 163
rect 403 162 404 163
rect 402 162 403 163
rect 401 162 402 163
rect 400 162 401 163
rect 399 162 400 163
rect 398 162 399 163
rect 397 162 398 163
rect 396 162 397 163
rect 395 162 396 163
rect 394 162 395 163
rect 393 162 394 163
rect 278 162 279 163
rect 277 162 278 163
rect 276 162 277 163
rect 275 162 276 163
rect 274 162 275 163
rect 273 162 274 163
rect 272 162 273 163
rect 271 162 272 163
rect 270 162 271 163
rect 269 162 270 163
rect 268 162 269 163
rect 267 162 268 163
rect 266 162 267 163
rect 265 162 266 163
rect 264 162 265 163
rect 263 162 264 163
rect 262 162 263 163
rect 261 162 262 163
rect 260 162 261 163
rect 259 162 260 163
rect 258 162 259 163
rect 257 162 258 163
rect 256 162 257 163
rect 255 162 256 163
rect 254 162 255 163
rect 253 162 254 163
rect 252 162 253 163
rect 251 162 252 163
rect 250 162 251 163
rect 249 162 250 163
rect 248 162 249 163
rect 247 162 248 163
rect 246 162 247 163
rect 245 162 246 163
rect 244 162 245 163
rect 243 162 244 163
rect 242 162 243 163
rect 241 162 242 163
rect 240 162 241 163
rect 239 162 240 163
rect 238 162 239 163
rect 237 162 238 163
rect 236 162 237 163
rect 235 162 236 163
rect 234 162 235 163
rect 233 162 234 163
rect 232 162 233 163
rect 231 162 232 163
rect 230 162 231 163
rect 229 162 230 163
rect 210 162 211 163
rect 209 162 210 163
rect 208 162 209 163
rect 207 162 208 163
rect 206 162 207 163
rect 205 162 206 163
rect 204 162 205 163
rect 203 162 204 163
rect 202 162 203 163
rect 201 162 202 163
rect 200 162 201 163
rect 199 162 200 163
rect 198 162 199 163
rect 197 162 198 163
rect 196 162 197 163
rect 195 162 196 163
rect 194 162 195 163
rect 193 162 194 163
rect 192 162 193 163
rect 191 162 192 163
rect 190 162 191 163
rect 189 162 190 163
rect 188 162 189 163
rect 187 162 188 163
rect 186 162 187 163
rect 185 162 186 163
rect 184 162 185 163
rect 183 162 184 163
rect 182 162 183 163
rect 181 162 182 163
rect 180 162 181 163
rect 179 162 180 163
rect 178 162 179 163
rect 177 162 178 163
rect 176 162 177 163
rect 175 162 176 163
rect 174 162 175 163
rect 173 162 174 163
rect 172 162 173 163
rect 171 162 172 163
rect 170 162 171 163
rect 169 162 170 163
rect 168 162 169 163
rect 167 162 168 163
rect 166 162 167 163
rect 165 162 166 163
rect 164 162 165 163
rect 163 162 164 163
rect 162 162 163 163
rect 161 162 162 163
rect 160 162 161 163
rect 159 162 160 163
rect 158 162 159 163
rect 157 162 158 163
rect 156 162 157 163
rect 155 162 156 163
rect 154 162 155 163
rect 153 162 154 163
rect 152 162 153 163
rect 151 162 152 163
rect 150 162 151 163
rect 149 162 150 163
rect 148 162 149 163
rect 147 162 148 163
rect 146 162 147 163
rect 145 162 146 163
rect 144 162 145 163
rect 143 162 144 163
rect 142 162 143 163
rect 141 162 142 163
rect 140 162 141 163
rect 139 162 140 163
rect 104 162 105 163
rect 103 162 104 163
rect 102 162 103 163
rect 101 162 102 163
rect 100 162 101 163
rect 99 162 100 163
rect 98 162 99 163
rect 97 162 98 163
rect 96 162 97 163
rect 95 162 96 163
rect 94 162 95 163
rect 93 162 94 163
rect 92 162 93 163
rect 91 162 92 163
rect 90 162 91 163
rect 89 162 90 163
rect 88 162 89 163
rect 87 162 88 163
rect 86 162 87 163
rect 85 162 86 163
rect 84 162 85 163
rect 83 162 84 163
rect 82 162 83 163
rect 81 162 82 163
rect 80 162 81 163
rect 79 162 80 163
rect 78 162 79 163
rect 77 162 78 163
rect 76 162 77 163
rect 75 162 76 163
rect 74 162 75 163
rect 73 162 74 163
rect 72 162 73 163
rect 71 162 72 163
rect 66 162 67 163
rect 65 162 66 163
rect 64 162 65 163
rect 63 162 64 163
rect 62 162 63 163
rect 61 162 62 163
rect 60 162 61 163
rect 59 162 60 163
rect 58 162 59 163
rect 57 162 58 163
rect 56 162 57 163
rect 55 162 56 163
rect 54 162 55 163
rect 53 162 54 163
rect 52 162 53 163
rect 51 162 52 163
rect 50 162 51 163
rect 49 162 50 163
rect 48 162 49 163
rect 47 162 48 163
rect 46 162 47 163
rect 45 162 46 163
rect 44 162 45 163
rect 43 162 44 163
rect 42 162 43 163
rect 41 162 42 163
rect 40 162 41 163
rect 39 162 40 163
rect 38 162 39 163
rect 37 162 38 163
rect 36 162 37 163
rect 35 162 36 163
rect 34 162 35 163
rect 33 162 34 163
rect 32 162 33 163
rect 31 162 32 163
rect 21 162 22 163
rect 20 162 21 163
rect 19 162 20 163
rect 18 162 19 163
rect 17 162 18 163
rect 16 162 17 163
rect 15 162 16 163
rect 14 162 15 163
rect 13 162 14 163
rect 12 162 13 163
rect 11 162 12 163
rect 10 162 11 163
rect 9 162 10 163
rect 8 162 9 163
rect 7 162 8 163
rect 6 162 7 163
rect 466 163 467 164
rect 465 163 466 164
rect 464 163 465 164
rect 463 163 464 164
rect 462 163 463 164
rect 461 163 462 164
rect 460 163 461 164
rect 459 163 460 164
rect 458 163 459 164
rect 437 163 438 164
rect 436 163 437 164
rect 435 163 436 164
rect 434 163 435 164
rect 433 163 434 164
rect 432 163 433 164
rect 431 163 432 164
rect 404 163 405 164
rect 403 163 404 164
rect 402 163 403 164
rect 401 163 402 164
rect 400 163 401 164
rect 399 163 400 164
rect 398 163 399 164
rect 397 163 398 164
rect 396 163 397 164
rect 395 163 396 164
rect 394 163 395 164
rect 393 163 394 164
rect 277 163 278 164
rect 276 163 277 164
rect 275 163 276 164
rect 274 163 275 164
rect 273 163 274 164
rect 272 163 273 164
rect 271 163 272 164
rect 270 163 271 164
rect 269 163 270 164
rect 268 163 269 164
rect 267 163 268 164
rect 266 163 267 164
rect 265 163 266 164
rect 264 163 265 164
rect 263 163 264 164
rect 262 163 263 164
rect 261 163 262 164
rect 260 163 261 164
rect 259 163 260 164
rect 258 163 259 164
rect 257 163 258 164
rect 256 163 257 164
rect 255 163 256 164
rect 254 163 255 164
rect 253 163 254 164
rect 252 163 253 164
rect 251 163 252 164
rect 250 163 251 164
rect 249 163 250 164
rect 248 163 249 164
rect 247 163 248 164
rect 246 163 247 164
rect 245 163 246 164
rect 244 163 245 164
rect 243 163 244 164
rect 242 163 243 164
rect 241 163 242 164
rect 240 163 241 164
rect 239 163 240 164
rect 238 163 239 164
rect 237 163 238 164
rect 236 163 237 164
rect 235 163 236 164
rect 234 163 235 164
rect 233 163 234 164
rect 232 163 233 164
rect 231 163 232 164
rect 230 163 231 164
rect 229 163 230 164
rect 228 163 229 164
rect 209 163 210 164
rect 208 163 209 164
rect 207 163 208 164
rect 206 163 207 164
rect 205 163 206 164
rect 204 163 205 164
rect 203 163 204 164
rect 202 163 203 164
rect 201 163 202 164
rect 200 163 201 164
rect 199 163 200 164
rect 198 163 199 164
rect 197 163 198 164
rect 196 163 197 164
rect 195 163 196 164
rect 194 163 195 164
rect 193 163 194 164
rect 192 163 193 164
rect 191 163 192 164
rect 190 163 191 164
rect 189 163 190 164
rect 188 163 189 164
rect 187 163 188 164
rect 186 163 187 164
rect 185 163 186 164
rect 184 163 185 164
rect 183 163 184 164
rect 182 163 183 164
rect 181 163 182 164
rect 180 163 181 164
rect 179 163 180 164
rect 178 163 179 164
rect 177 163 178 164
rect 176 163 177 164
rect 175 163 176 164
rect 174 163 175 164
rect 173 163 174 164
rect 172 163 173 164
rect 171 163 172 164
rect 170 163 171 164
rect 169 163 170 164
rect 168 163 169 164
rect 167 163 168 164
rect 166 163 167 164
rect 165 163 166 164
rect 164 163 165 164
rect 163 163 164 164
rect 162 163 163 164
rect 161 163 162 164
rect 160 163 161 164
rect 159 163 160 164
rect 158 163 159 164
rect 157 163 158 164
rect 156 163 157 164
rect 155 163 156 164
rect 154 163 155 164
rect 153 163 154 164
rect 152 163 153 164
rect 151 163 152 164
rect 150 163 151 164
rect 149 163 150 164
rect 148 163 149 164
rect 147 163 148 164
rect 146 163 147 164
rect 145 163 146 164
rect 144 163 145 164
rect 143 163 144 164
rect 142 163 143 164
rect 141 163 142 164
rect 140 163 141 164
rect 139 163 140 164
rect 138 163 139 164
rect 102 163 103 164
rect 101 163 102 164
rect 100 163 101 164
rect 99 163 100 164
rect 98 163 99 164
rect 97 163 98 164
rect 96 163 97 164
rect 95 163 96 164
rect 94 163 95 164
rect 93 163 94 164
rect 92 163 93 164
rect 91 163 92 164
rect 90 163 91 164
rect 89 163 90 164
rect 88 163 89 164
rect 87 163 88 164
rect 86 163 87 164
rect 85 163 86 164
rect 84 163 85 164
rect 83 163 84 164
rect 82 163 83 164
rect 81 163 82 164
rect 80 163 81 164
rect 79 163 80 164
rect 78 163 79 164
rect 77 163 78 164
rect 76 163 77 164
rect 64 163 65 164
rect 63 163 64 164
rect 62 163 63 164
rect 61 163 62 164
rect 60 163 61 164
rect 59 163 60 164
rect 58 163 59 164
rect 57 163 58 164
rect 56 163 57 164
rect 55 163 56 164
rect 54 163 55 164
rect 53 163 54 164
rect 52 163 53 164
rect 51 163 52 164
rect 50 163 51 164
rect 49 163 50 164
rect 48 163 49 164
rect 47 163 48 164
rect 46 163 47 164
rect 45 163 46 164
rect 44 163 45 164
rect 43 163 44 164
rect 42 163 43 164
rect 41 163 42 164
rect 40 163 41 164
rect 39 163 40 164
rect 38 163 39 164
rect 37 163 38 164
rect 36 163 37 164
rect 35 163 36 164
rect 34 163 35 164
rect 33 163 34 164
rect 32 163 33 164
rect 31 163 32 164
rect 21 163 22 164
rect 20 163 21 164
rect 19 163 20 164
rect 18 163 19 164
rect 17 163 18 164
rect 16 163 17 164
rect 15 163 16 164
rect 14 163 15 164
rect 13 163 14 164
rect 12 163 13 164
rect 11 163 12 164
rect 10 163 11 164
rect 9 163 10 164
rect 8 163 9 164
rect 7 163 8 164
rect 6 163 7 164
rect 468 164 469 165
rect 467 164 468 165
rect 466 164 467 165
rect 465 164 466 165
rect 464 164 465 165
rect 463 164 464 165
rect 462 164 463 165
rect 461 164 462 165
rect 460 164 461 165
rect 459 164 460 165
rect 458 164 459 165
rect 437 164 438 165
rect 436 164 437 165
rect 435 164 436 165
rect 434 164 435 165
rect 405 164 406 165
rect 404 164 405 165
rect 403 164 404 165
rect 402 164 403 165
rect 401 164 402 165
rect 400 164 401 165
rect 399 164 400 165
rect 398 164 399 165
rect 397 164 398 165
rect 396 164 397 165
rect 395 164 396 165
rect 394 164 395 165
rect 393 164 394 165
rect 275 164 276 165
rect 274 164 275 165
rect 273 164 274 165
rect 272 164 273 165
rect 271 164 272 165
rect 270 164 271 165
rect 269 164 270 165
rect 268 164 269 165
rect 267 164 268 165
rect 266 164 267 165
rect 265 164 266 165
rect 264 164 265 165
rect 263 164 264 165
rect 262 164 263 165
rect 261 164 262 165
rect 260 164 261 165
rect 259 164 260 165
rect 258 164 259 165
rect 257 164 258 165
rect 256 164 257 165
rect 255 164 256 165
rect 254 164 255 165
rect 253 164 254 165
rect 252 164 253 165
rect 251 164 252 165
rect 250 164 251 165
rect 249 164 250 165
rect 248 164 249 165
rect 247 164 248 165
rect 246 164 247 165
rect 245 164 246 165
rect 244 164 245 165
rect 243 164 244 165
rect 242 164 243 165
rect 241 164 242 165
rect 240 164 241 165
rect 239 164 240 165
rect 238 164 239 165
rect 237 164 238 165
rect 236 164 237 165
rect 235 164 236 165
rect 234 164 235 165
rect 233 164 234 165
rect 232 164 233 165
rect 231 164 232 165
rect 230 164 231 165
rect 229 164 230 165
rect 228 164 229 165
rect 209 164 210 165
rect 208 164 209 165
rect 207 164 208 165
rect 206 164 207 165
rect 205 164 206 165
rect 204 164 205 165
rect 203 164 204 165
rect 202 164 203 165
rect 201 164 202 165
rect 200 164 201 165
rect 199 164 200 165
rect 198 164 199 165
rect 197 164 198 165
rect 196 164 197 165
rect 195 164 196 165
rect 194 164 195 165
rect 193 164 194 165
rect 192 164 193 165
rect 191 164 192 165
rect 190 164 191 165
rect 189 164 190 165
rect 188 164 189 165
rect 187 164 188 165
rect 186 164 187 165
rect 185 164 186 165
rect 184 164 185 165
rect 183 164 184 165
rect 182 164 183 165
rect 181 164 182 165
rect 180 164 181 165
rect 179 164 180 165
rect 178 164 179 165
rect 177 164 178 165
rect 176 164 177 165
rect 175 164 176 165
rect 174 164 175 165
rect 173 164 174 165
rect 172 164 173 165
rect 171 164 172 165
rect 170 164 171 165
rect 169 164 170 165
rect 168 164 169 165
rect 167 164 168 165
rect 166 164 167 165
rect 165 164 166 165
rect 164 164 165 165
rect 163 164 164 165
rect 162 164 163 165
rect 161 164 162 165
rect 160 164 161 165
rect 159 164 160 165
rect 158 164 159 165
rect 157 164 158 165
rect 156 164 157 165
rect 155 164 156 165
rect 154 164 155 165
rect 153 164 154 165
rect 152 164 153 165
rect 151 164 152 165
rect 150 164 151 165
rect 149 164 150 165
rect 148 164 149 165
rect 147 164 148 165
rect 146 164 147 165
rect 145 164 146 165
rect 144 164 145 165
rect 143 164 144 165
rect 142 164 143 165
rect 141 164 142 165
rect 140 164 141 165
rect 139 164 140 165
rect 138 164 139 165
rect 137 164 138 165
rect 99 164 100 165
rect 98 164 99 165
rect 97 164 98 165
rect 96 164 97 165
rect 95 164 96 165
rect 94 164 95 165
rect 93 164 94 165
rect 92 164 93 165
rect 91 164 92 165
rect 90 164 91 165
rect 89 164 90 165
rect 88 164 89 165
rect 87 164 88 165
rect 86 164 87 165
rect 85 164 86 165
rect 84 164 85 165
rect 83 164 84 165
rect 82 164 83 165
rect 81 164 82 165
rect 80 164 81 165
rect 62 164 63 165
rect 61 164 62 165
rect 60 164 61 165
rect 59 164 60 165
rect 58 164 59 165
rect 57 164 58 165
rect 56 164 57 165
rect 55 164 56 165
rect 54 164 55 165
rect 53 164 54 165
rect 52 164 53 165
rect 51 164 52 165
rect 50 164 51 165
rect 49 164 50 165
rect 48 164 49 165
rect 47 164 48 165
rect 46 164 47 165
rect 45 164 46 165
rect 44 164 45 165
rect 43 164 44 165
rect 42 164 43 165
rect 41 164 42 165
rect 40 164 41 165
rect 39 164 40 165
rect 38 164 39 165
rect 37 164 38 165
rect 36 164 37 165
rect 35 164 36 165
rect 34 164 35 165
rect 33 164 34 165
rect 32 164 33 165
rect 31 164 32 165
rect 21 164 22 165
rect 20 164 21 165
rect 19 164 20 165
rect 18 164 19 165
rect 17 164 18 165
rect 16 164 17 165
rect 15 164 16 165
rect 14 164 15 165
rect 13 164 14 165
rect 12 164 13 165
rect 11 164 12 165
rect 10 164 11 165
rect 9 164 10 165
rect 8 164 9 165
rect 7 164 8 165
rect 6 164 7 165
rect 471 165 472 166
rect 470 165 471 166
rect 469 165 470 166
rect 468 165 469 166
rect 467 165 468 166
rect 466 165 467 166
rect 465 165 466 166
rect 464 165 465 166
rect 463 165 464 166
rect 462 165 463 166
rect 461 165 462 166
rect 460 165 461 166
rect 459 165 460 166
rect 458 165 459 166
rect 437 165 438 166
rect 436 165 437 166
rect 435 165 436 166
rect 407 165 408 166
rect 406 165 407 166
rect 405 165 406 166
rect 404 165 405 166
rect 403 165 404 166
rect 402 165 403 166
rect 401 165 402 166
rect 400 165 401 166
rect 399 165 400 166
rect 398 165 399 166
rect 397 165 398 166
rect 396 165 397 166
rect 395 165 396 166
rect 394 165 395 166
rect 393 165 394 166
rect 274 165 275 166
rect 273 165 274 166
rect 272 165 273 166
rect 271 165 272 166
rect 270 165 271 166
rect 269 165 270 166
rect 268 165 269 166
rect 267 165 268 166
rect 266 165 267 166
rect 265 165 266 166
rect 264 165 265 166
rect 263 165 264 166
rect 262 165 263 166
rect 261 165 262 166
rect 260 165 261 166
rect 259 165 260 166
rect 258 165 259 166
rect 257 165 258 166
rect 256 165 257 166
rect 255 165 256 166
rect 254 165 255 166
rect 253 165 254 166
rect 252 165 253 166
rect 251 165 252 166
rect 250 165 251 166
rect 249 165 250 166
rect 248 165 249 166
rect 247 165 248 166
rect 246 165 247 166
rect 245 165 246 166
rect 244 165 245 166
rect 243 165 244 166
rect 242 165 243 166
rect 241 165 242 166
rect 240 165 241 166
rect 239 165 240 166
rect 238 165 239 166
rect 237 165 238 166
rect 236 165 237 166
rect 235 165 236 166
rect 234 165 235 166
rect 233 165 234 166
rect 232 165 233 166
rect 231 165 232 166
rect 230 165 231 166
rect 229 165 230 166
rect 228 165 229 166
rect 227 165 228 166
rect 208 165 209 166
rect 207 165 208 166
rect 206 165 207 166
rect 205 165 206 166
rect 204 165 205 166
rect 203 165 204 166
rect 202 165 203 166
rect 201 165 202 166
rect 200 165 201 166
rect 199 165 200 166
rect 198 165 199 166
rect 197 165 198 166
rect 196 165 197 166
rect 195 165 196 166
rect 194 165 195 166
rect 193 165 194 166
rect 192 165 193 166
rect 191 165 192 166
rect 190 165 191 166
rect 189 165 190 166
rect 188 165 189 166
rect 187 165 188 166
rect 186 165 187 166
rect 185 165 186 166
rect 184 165 185 166
rect 183 165 184 166
rect 182 165 183 166
rect 181 165 182 166
rect 180 165 181 166
rect 179 165 180 166
rect 178 165 179 166
rect 177 165 178 166
rect 176 165 177 166
rect 175 165 176 166
rect 174 165 175 166
rect 173 165 174 166
rect 172 165 173 166
rect 171 165 172 166
rect 170 165 171 166
rect 169 165 170 166
rect 168 165 169 166
rect 167 165 168 166
rect 166 165 167 166
rect 165 165 166 166
rect 164 165 165 166
rect 163 165 164 166
rect 162 165 163 166
rect 161 165 162 166
rect 160 165 161 166
rect 159 165 160 166
rect 158 165 159 166
rect 157 165 158 166
rect 156 165 157 166
rect 155 165 156 166
rect 154 165 155 166
rect 153 165 154 166
rect 152 165 153 166
rect 151 165 152 166
rect 150 165 151 166
rect 149 165 150 166
rect 148 165 149 166
rect 147 165 148 166
rect 146 165 147 166
rect 145 165 146 166
rect 144 165 145 166
rect 143 165 144 166
rect 142 165 143 166
rect 141 165 142 166
rect 140 165 141 166
rect 139 165 140 166
rect 138 165 139 166
rect 137 165 138 166
rect 136 165 137 166
rect 135 165 136 166
rect 95 165 96 166
rect 94 165 95 166
rect 93 165 94 166
rect 92 165 93 166
rect 91 165 92 166
rect 90 165 91 166
rect 89 165 90 166
rect 88 165 89 166
rect 87 165 88 166
rect 86 165 87 166
rect 61 165 62 166
rect 60 165 61 166
rect 59 165 60 166
rect 58 165 59 166
rect 57 165 58 166
rect 56 165 57 166
rect 55 165 56 166
rect 54 165 55 166
rect 53 165 54 166
rect 52 165 53 166
rect 51 165 52 166
rect 50 165 51 166
rect 49 165 50 166
rect 48 165 49 166
rect 47 165 48 166
rect 46 165 47 166
rect 45 165 46 166
rect 44 165 45 166
rect 43 165 44 166
rect 42 165 43 166
rect 41 165 42 166
rect 40 165 41 166
rect 39 165 40 166
rect 38 165 39 166
rect 37 165 38 166
rect 36 165 37 166
rect 35 165 36 166
rect 34 165 35 166
rect 33 165 34 166
rect 32 165 33 166
rect 31 165 32 166
rect 21 165 22 166
rect 20 165 21 166
rect 19 165 20 166
rect 18 165 19 166
rect 17 165 18 166
rect 16 165 17 166
rect 15 165 16 166
rect 14 165 15 166
rect 13 165 14 166
rect 12 165 13 166
rect 11 165 12 166
rect 10 165 11 166
rect 9 165 10 166
rect 8 165 9 166
rect 7 165 8 166
rect 473 166 474 167
rect 472 166 473 167
rect 471 166 472 167
rect 470 166 471 167
rect 469 166 470 167
rect 468 166 469 167
rect 467 166 468 167
rect 466 166 467 167
rect 465 166 466 167
rect 464 166 465 167
rect 463 166 464 167
rect 462 166 463 167
rect 461 166 462 167
rect 459 166 460 167
rect 458 166 459 167
rect 437 166 438 167
rect 436 166 437 167
rect 435 166 436 167
rect 408 166 409 167
rect 407 166 408 167
rect 406 166 407 167
rect 405 166 406 167
rect 404 166 405 167
rect 403 166 404 167
rect 402 166 403 167
rect 401 166 402 167
rect 400 166 401 167
rect 399 166 400 167
rect 398 166 399 167
rect 397 166 398 167
rect 396 166 397 167
rect 395 166 396 167
rect 394 166 395 167
rect 273 166 274 167
rect 272 166 273 167
rect 271 166 272 167
rect 270 166 271 167
rect 269 166 270 167
rect 268 166 269 167
rect 267 166 268 167
rect 266 166 267 167
rect 265 166 266 167
rect 264 166 265 167
rect 263 166 264 167
rect 262 166 263 167
rect 261 166 262 167
rect 260 166 261 167
rect 259 166 260 167
rect 258 166 259 167
rect 257 166 258 167
rect 256 166 257 167
rect 255 166 256 167
rect 254 166 255 167
rect 253 166 254 167
rect 252 166 253 167
rect 251 166 252 167
rect 250 166 251 167
rect 249 166 250 167
rect 248 166 249 167
rect 247 166 248 167
rect 246 166 247 167
rect 245 166 246 167
rect 244 166 245 167
rect 243 166 244 167
rect 242 166 243 167
rect 241 166 242 167
rect 240 166 241 167
rect 239 166 240 167
rect 238 166 239 167
rect 237 166 238 167
rect 236 166 237 167
rect 235 166 236 167
rect 234 166 235 167
rect 233 166 234 167
rect 232 166 233 167
rect 231 166 232 167
rect 230 166 231 167
rect 229 166 230 167
rect 228 166 229 167
rect 227 166 228 167
rect 208 166 209 167
rect 207 166 208 167
rect 206 166 207 167
rect 205 166 206 167
rect 204 166 205 167
rect 203 166 204 167
rect 202 166 203 167
rect 201 166 202 167
rect 200 166 201 167
rect 199 166 200 167
rect 198 166 199 167
rect 197 166 198 167
rect 196 166 197 167
rect 195 166 196 167
rect 194 166 195 167
rect 193 166 194 167
rect 192 166 193 167
rect 191 166 192 167
rect 190 166 191 167
rect 189 166 190 167
rect 188 166 189 167
rect 187 166 188 167
rect 186 166 187 167
rect 185 166 186 167
rect 184 166 185 167
rect 183 166 184 167
rect 182 166 183 167
rect 181 166 182 167
rect 180 166 181 167
rect 179 166 180 167
rect 178 166 179 167
rect 177 166 178 167
rect 176 166 177 167
rect 175 166 176 167
rect 174 166 175 167
rect 173 166 174 167
rect 172 166 173 167
rect 171 166 172 167
rect 170 166 171 167
rect 169 166 170 167
rect 168 166 169 167
rect 167 166 168 167
rect 166 166 167 167
rect 165 166 166 167
rect 164 166 165 167
rect 163 166 164 167
rect 162 166 163 167
rect 161 166 162 167
rect 160 166 161 167
rect 159 166 160 167
rect 158 166 159 167
rect 157 166 158 167
rect 156 166 157 167
rect 155 166 156 167
rect 154 166 155 167
rect 153 166 154 167
rect 152 166 153 167
rect 151 166 152 167
rect 150 166 151 167
rect 149 166 150 167
rect 148 166 149 167
rect 147 166 148 167
rect 146 166 147 167
rect 145 166 146 167
rect 144 166 145 167
rect 143 166 144 167
rect 142 166 143 167
rect 141 166 142 167
rect 140 166 141 167
rect 139 166 140 167
rect 138 166 139 167
rect 137 166 138 167
rect 136 166 137 167
rect 135 166 136 167
rect 134 166 135 167
rect 60 166 61 167
rect 59 166 60 167
rect 58 166 59 167
rect 57 166 58 167
rect 56 166 57 167
rect 55 166 56 167
rect 54 166 55 167
rect 53 166 54 167
rect 52 166 53 167
rect 51 166 52 167
rect 50 166 51 167
rect 49 166 50 167
rect 48 166 49 167
rect 47 166 48 167
rect 46 166 47 167
rect 45 166 46 167
rect 44 166 45 167
rect 43 166 44 167
rect 42 166 43 167
rect 41 166 42 167
rect 40 166 41 167
rect 39 166 40 167
rect 38 166 39 167
rect 37 166 38 167
rect 36 166 37 167
rect 35 166 36 167
rect 34 166 35 167
rect 33 166 34 167
rect 32 166 33 167
rect 31 166 32 167
rect 21 166 22 167
rect 20 166 21 167
rect 19 166 20 167
rect 18 166 19 167
rect 17 166 18 167
rect 16 166 17 167
rect 15 166 16 167
rect 14 166 15 167
rect 13 166 14 167
rect 12 166 13 167
rect 11 166 12 167
rect 10 166 11 167
rect 9 166 10 167
rect 8 166 9 167
rect 7 166 8 167
rect 476 167 477 168
rect 475 167 476 168
rect 474 167 475 168
rect 473 167 474 168
rect 472 167 473 168
rect 471 167 472 168
rect 470 167 471 168
rect 469 167 470 168
rect 468 167 469 168
rect 467 167 468 168
rect 466 167 467 168
rect 465 167 466 168
rect 464 167 465 168
rect 458 167 459 168
rect 437 167 438 168
rect 436 167 437 168
rect 435 167 436 168
rect 409 167 410 168
rect 408 167 409 168
rect 407 167 408 168
rect 406 167 407 168
rect 405 167 406 168
rect 404 167 405 168
rect 403 167 404 168
rect 402 167 403 168
rect 401 167 402 168
rect 400 167 401 168
rect 399 167 400 168
rect 398 167 399 168
rect 397 167 398 168
rect 396 167 397 168
rect 272 167 273 168
rect 271 167 272 168
rect 270 167 271 168
rect 269 167 270 168
rect 268 167 269 168
rect 267 167 268 168
rect 266 167 267 168
rect 265 167 266 168
rect 264 167 265 168
rect 263 167 264 168
rect 262 167 263 168
rect 261 167 262 168
rect 260 167 261 168
rect 259 167 260 168
rect 258 167 259 168
rect 257 167 258 168
rect 256 167 257 168
rect 255 167 256 168
rect 254 167 255 168
rect 253 167 254 168
rect 252 167 253 168
rect 251 167 252 168
rect 250 167 251 168
rect 249 167 250 168
rect 248 167 249 168
rect 247 167 248 168
rect 246 167 247 168
rect 245 167 246 168
rect 244 167 245 168
rect 243 167 244 168
rect 242 167 243 168
rect 241 167 242 168
rect 240 167 241 168
rect 239 167 240 168
rect 238 167 239 168
rect 237 167 238 168
rect 236 167 237 168
rect 235 167 236 168
rect 234 167 235 168
rect 233 167 234 168
rect 232 167 233 168
rect 231 167 232 168
rect 230 167 231 168
rect 229 167 230 168
rect 228 167 229 168
rect 227 167 228 168
rect 226 167 227 168
rect 207 167 208 168
rect 206 167 207 168
rect 205 167 206 168
rect 204 167 205 168
rect 203 167 204 168
rect 202 167 203 168
rect 201 167 202 168
rect 200 167 201 168
rect 199 167 200 168
rect 198 167 199 168
rect 197 167 198 168
rect 196 167 197 168
rect 195 167 196 168
rect 194 167 195 168
rect 193 167 194 168
rect 192 167 193 168
rect 191 167 192 168
rect 190 167 191 168
rect 189 167 190 168
rect 188 167 189 168
rect 187 167 188 168
rect 186 167 187 168
rect 185 167 186 168
rect 184 167 185 168
rect 183 167 184 168
rect 182 167 183 168
rect 181 167 182 168
rect 180 167 181 168
rect 179 167 180 168
rect 178 167 179 168
rect 177 167 178 168
rect 176 167 177 168
rect 175 167 176 168
rect 174 167 175 168
rect 173 167 174 168
rect 172 167 173 168
rect 171 167 172 168
rect 170 167 171 168
rect 169 167 170 168
rect 168 167 169 168
rect 167 167 168 168
rect 166 167 167 168
rect 165 167 166 168
rect 164 167 165 168
rect 163 167 164 168
rect 162 167 163 168
rect 161 167 162 168
rect 160 167 161 168
rect 159 167 160 168
rect 158 167 159 168
rect 157 167 158 168
rect 156 167 157 168
rect 155 167 156 168
rect 154 167 155 168
rect 153 167 154 168
rect 152 167 153 168
rect 151 167 152 168
rect 150 167 151 168
rect 149 167 150 168
rect 148 167 149 168
rect 147 167 148 168
rect 146 167 147 168
rect 145 167 146 168
rect 144 167 145 168
rect 143 167 144 168
rect 142 167 143 168
rect 141 167 142 168
rect 140 167 141 168
rect 139 167 140 168
rect 138 167 139 168
rect 137 167 138 168
rect 136 167 137 168
rect 135 167 136 168
rect 134 167 135 168
rect 133 167 134 168
rect 59 167 60 168
rect 58 167 59 168
rect 57 167 58 168
rect 56 167 57 168
rect 55 167 56 168
rect 54 167 55 168
rect 53 167 54 168
rect 52 167 53 168
rect 51 167 52 168
rect 50 167 51 168
rect 49 167 50 168
rect 48 167 49 168
rect 47 167 48 168
rect 46 167 47 168
rect 45 167 46 168
rect 44 167 45 168
rect 43 167 44 168
rect 42 167 43 168
rect 41 167 42 168
rect 40 167 41 168
rect 39 167 40 168
rect 38 167 39 168
rect 37 167 38 168
rect 36 167 37 168
rect 35 167 36 168
rect 34 167 35 168
rect 33 167 34 168
rect 32 167 33 168
rect 31 167 32 168
rect 21 167 22 168
rect 20 167 21 168
rect 19 167 20 168
rect 18 167 19 168
rect 17 167 18 168
rect 16 167 17 168
rect 15 167 16 168
rect 14 167 15 168
rect 13 167 14 168
rect 12 167 13 168
rect 11 167 12 168
rect 10 167 11 168
rect 9 167 10 168
rect 8 167 9 168
rect 7 167 8 168
rect 479 168 480 169
rect 478 168 479 169
rect 477 168 478 169
rect 476 168 477 169
rect 475 168 476 169
rect 474 168 475 169
rect 473 168 474 169
rect 472 168 473 169
rect 471 168 472 169
rect 470 168 471 169
rect 469 168 470 169
rect 468 168 469 169
rect 467 168 468 169
rect 437 168 438 169
rect 436 168 437 169
rect 435 168 436 169
rect 410 168 411 169
rect 409 168 410 169
rect 408 168 409 169
rect 407 168 408 169
rect 406 168 407 169
rect 405 168 406 169
rect 404 168 405 169
rect 403 168 404 169
rect 402 168 403 169
rect 401 168 402 169
rect 400 168 401 169
rect 399 168 400 169
rect 398 168 399 169
rect 397 168 398 169
rect 270 168 271 169
rect 269 168 270 169
rect 268 168 269 169
rect 267 168 268 169
rect 266 168 267 169
rect 265 168 266 169
rect 264 168 265 169
rect 263 168 264 169
rect 262 168 263 169
rect 261 168 262 169
rect 260 168 261 169
rect 259 168 260 169
rect 258 168 259 169
rect 257 168 258 169
rect 256 168 257 169
rect 255 168 256 169
rect 254 168 255 169
rect 253 168 254 169
rect 252 168 253 169
rect 251 168 252 169
rect 250 168 251 169
rect 249 168 250 169
rect 248 168 249 169
rect 247 168 248 169
rect 246 168 247 169
rect 245 168 246 169
rect 244 168 245 169
rect 243 168 244 169
rect 242 168 243 169
rect 241 168 242 169
rect 240 168 241 169
rect 239 168 240 169
rect 238 168 239 169
rect 237 168 238 169
rect 236 168 237 169
rect 235 168 236 169
rect 234 168 235 169
rect 233 168 234 169
rect 232 168 233 169
rect 231 168 232 169
rect 230 168 231 169
rect 229 168 230 169
rect 228 168 229 169
rect 227 168 228 169
rect 226 168 227 169
rect 207 168 208 169
rect 206 168 207 169
rect 205 168 206 169
rect 204 168 205 169
rect 203 168 204 169
rect 202 168 203 169
rect 201 168 202 169
rect 200 168 201 169
rect 199 168 200 169
rect 198 168 199 169
rect 197 168 198 169
rect 196 168 197 169
rect 195 168 196 169
rect 194 168 195 169
rect 193 168 194 169
rect 192 168 193 169
rect 191 168 192 169
rect 190 168 191 169
rect 189 168 190 169
rect 188 168 189 169
rect 187 168 188 169
rect 186 168 187 169
rect 185 168 186 169
rect 184 168 185 169
rect 183 168 184 169
rect 182 168 183 169
rect 181 168 182 169
rect 180 168 181 169
rect 179 168 180 169
rect 178 168 179 169
rect 177 168 178 169
rect 176 168 177 169
rect 175 168 176 169
rect 174 168 175 169
rect 173 168 174 169
rect 172 168 173 169
rect 171 168 172 169
rect 170 168 171 169
rect 169 168 170 169
rect 168 168 169 169
rect 167 168 168 169
rect 166 168 167 169
rect 165 168 166 169
rect 164 168 165 169
rect 163 168 164 169
rect 162 168 163 169
rect 161 168 162 169
rect 160 168 161 169
rect 159 168 160 169
rect 158 168 159 169
rect 157 168 158 169
rect 156 168 157 169
rect 155 168 156 169
rect 154 168 155 169
rect 153 168 154 169
rect 152 168 153 169
rect 151 168 152 169
rect 150 168 151 169
rect 149 168 150 169
rect 148 168 149 169
rect 147 168 148 169
rect 146 168 147 169
rect 145 168 146 169
rect 144 168 145 169
rect 143 168 144 169
rect 142 168 143 169
rect 141 168 142 169
rect 140 168 141 169
rect 139 168 140 169
rect 138 168 139 169
rect 137 168 138 169
rect 136 168 137 169
rect 135 168 136 169
rect 134 168 135 169
rect 133 168 134 169
rect 132 168 133 169
rect 131 168 132 169
rect 58 168 59 169
rect 57 168 58 169
rect 56 168 57 169
rect 55 168 56 169
rect 54 168 55 169
rect 53 168 54 169
rect 52 168 53 169
rect 51 168 52 169
rect 50 168 51 169
rect 49 168 50 169
rect 48 168 49 169
rect 47 168 48 169
rect 46 168 47 169
rect 45 168 46 169
rect 44 168 45 169
rect 43 168 44 169
rect 42 168 43 169
rect 41 168 42 169
rect 40 168 41 169
rect 39 168 40 169
rect 38 168 39 169
rect 37 168 38 169
rect 36 168 37 169
rect 35 168 36 169
rect 34 168 35 169
rect 33 168 34 169
rect 32 168 33 169
rect 31 168 32 169
rect 21 168 22 169
rect 20 168 21 169
rect 19 168 20 169
rect 18 168 19 169
rect 17 168 18 169
rect 16 168 17 169
rect 15 168 16 169
rect 14 168 15 169
rect 13 168 14 169
rect 12 168 13 169
rect 11 168 12 169
rect 10 168 11 169
rect 9 168 10 169
rect 8 168 9 169
rect 7 168 8 169
rect 479 169 480 170
rect 478 169 479 170
rect 477 169 478 170
rect 476 169 477 170
rect 475 169 476 170
rect 474 169 475 170
rect 473 169 474 170
rect 472 169 473 170
rect 471 169 472 170
rect 470 169 471 170
rect 469 169 470 170
rect 437 169 438 170
rect 436 169 437 170
rect 411 169 412 170
rect 410 169 411 170
rect 409 169 410 170
rect 408 169 409 170
rect 407 169 408 170
rect 406 169 407 170
rect 405 169 406 170
rect 404 169 405 170
rect 403 169 404 170
rect 402 169 403 170
rect 401 169 402 170
rect 400 169 401 170
rect 399 169 400 170
rect 398 169 399 170
rect 269 169 270 170
rect 268 169 269 170
rect 267 169 268 170
rect 266 169 267 170
rect 265 169 266 170
rect 264 169 265 170
rect 263 169 264 170
rect 262 169 263 170
rect 261 169 262 170
rect 260 169 261 170
rect 259 169 260 170
rect 258 169 259 170
rect 257 169 258 170
rect 256 169 257 170
rect 255 169 256 170
rect 254 169 255 170
rect 253 169 254 170
rect 252 169 253 170
rect 251 169 252 170
rect 250 169 251 170
rect 249 169 250 170
rect 248 169 249 170
rect 247 169 248 170
rect 246 169 247 170
rect 245 169 246 170
rect 244 169 245 170
rect 243 169 244 170
rect 242 169 243 170
rect 241 169 242 170
rect 240 169 241 170
rect 239 169 240 170
rect 238 169 239 170
rect 237 169 238 170
rect 236 169 237 170
rect 235 169 236 170
rect 234 169 235 170
rect 233 169 234 170
rect 232 169 233 170
rect 231 169 232 170
rect 230 169 231 170
rect 229 169 230 170
rect 228 169 229 170
rect 227 169 228 170
rect 226 169 227 170
rect 225 169 226 170
rect 206 169 207 170
rect 205 169 206 170
rect 204 169 205 170
rect 203 169 204 170
rect 202 169 203 170
rect 201 169 202 170
rect 200 169 201 170
rect 199 169 200 170
rect 198 169 199 170
rect 197 169 198 170
rect 196 169 197 170
rect 195 169 196 170
rect 194 169 195 170
rect 193 169 194 170
rect 192 169 193 170
rect 191 169 192 170
rect 190 169 191 170
rect 189 169 190 170
rect 188 169 189 170
rect 187 169 188 170
rect 186 169 187 170
rect 185 169 186 170
rect 184 169 185 170
rect 183 169 184 170
rect 182 169 183 170
rect 181 169 182 170
rect 180 169 181 170
rect 179 169 180 170
rect 178 169 179 170
rect 177 169 178 170
rect 176 169 177 170
rect 175 169 176 170
rect 174 169 175 170
rect 173 169 174 170
rect 172 169 173 170
rect 171 169 172 170
rect 170 169 171 170
rect 169 169 170 170
rect 168 169 169 170
rect 167 169 168 170
rect 166 169 167 170
rect 165 169 166 170
rect 164 169 165 170
rect 163 169 164 170
rect 162 169 163 170
rect 161 169 162 170
rect 160 169 161 170
rect 159 169 160 170
rect 158 169 159 170
rect 157 169 158 170
rect 156 169 157 170
rect 155 169 156 170
rect 154 169 155 170
rect 153 169 154 170
rect 152 169 153 170
rect 151 169 152 170
rect 150 169 151 170
rect 149 169 150 170
rect 148 169 149 170
rect 147 169 148 170
rect 146 169 147 170
rect 145 169 146 170
rect 144 169 145 170
rect 143 169 144 170
rect 142 169 143 170
rect 141 169 142 170
rect 140 169 141 170
rect 139 169 140 170
rect 138 169 139 170
rect 137 169 138 170
rect 136 169 137 170
rect 135 169 136 170
rect 134 169 135 170
rect 133 169 134 170
rect 132 169 133 170
rect 131 169 132 170
rect 130 169 131 170
rect 57 169 58 170
rect 56 169 57 170
rect 55 169 56 170
rect 54 169 55 170
rect 53 169 54 170
rect 52 169 53 170
rect 51 169 52 170
rect 50 169 51 170
rect 49 169 50 170
rect 48 169 49 170
rect 47 169 48 170
rect 46 169 47 170
rect 45 169 46 170
rect 44 169 45 170
rect 43 169 44 170
rect 42 169 43 170
rect 41 169 42 170
rect 40 169 41 170
rect 39 169 40 170
rect 38 169 39 170
rect 37 169 38 170
rect 36 169 37 170
rect 35 169 36 170
rect 34 169 35 170
rect 33 169 34 170
rect 32 169 33 170
rect 20 169 21 170
rect 19 169 20 170
rect 18 169 19 170
rect 17 169 18 170
rect 16 169 17 170
rect 15 169 16 170
rect 14 169 15 170
rect 13 169 14 170
rect 12 169 13 170
rect 11 169 12 170
rect 10 169 11 170
rect 9 169 10 170
rect 8 169 9 170
rect 478 170 479 171
rect 477 170 478 171
rect 476 170 477 171
rect 475 170 476 171
rect 474 170 475 171
rect 473 170 474 171
rect 472 170 473 171
rect 412 170 413 171
rect 411 170 412 171
rect 410 170 411 171
rect 409 170 410 171
rect 408 170 409 171
rect 407 170 408 171
rect 406 170 407 171
rect 405 170 406 171
rect 404 170 405 171
rect 403 170 404 171
rect 402 170 403 171
rect 401 170 402 171
rect 400 170 401 171
rect 399 170 400 171
rect 268 170 269 171
rect 267 170 268 171
rect 266 170 267 171
rect 265 170 266 171
rect 264 170 265 171
rect 263 170 264 171
rect 262 170 263 171
rect 261 170 262 171
rect 260 170 261 171
rect 259 170 260 171
rect 258 170 259 171
rect 257 170 258 171
rect 256 170 257 171
rect 255 170 256 171
rect 254 170 255 171
rect 253 170 254 171
rect 252 170 253 171
rect 251 170 252 171
rect 250 170 251 171
rect 249 170 250 171
rect 248 170 249 171
rect 247 170 248 171
rect 246 170 247 171
rect 245 170 246 171
rect 244 170 245 171
rect 243 170 244 171
rect 242 170 243 171
rect 241 170 242 171
rect 240 170 241 171
rect 239 170 240 171
rect 238 170 239 171
rect 237 170 238 171
rect 236 170 237 171
rect 235 170 236 171
rect 234 170 235 171
rect 233 170 234 171
rect 232 170 233 171
rect 231 170 232 171
rect 230 170 231 171
rect 229 170 230 171
rect 228 170 229 171
rect 227 170 228 171
rect 226 170 227 171
rect 225 170 226 171
rect 224 170 225 171
rect 206 170 207 171
rect 205 170 206 171
rect 204 170 205 171
rect 203 170 204 171
rect 202 170 203 171
rect 201 170 202 171
rect 200 170 201 171
rect 199 170 200 171
rect 198 170 199 171
rect 197 170 198 171
rect 196 170 197 171
rect 195 170 196 171
rect 194 170 195 171
rect 193 170 194 171
rect 192 170 193 171
rect 191 170 192 171
rect 190 170 191 171
rect 189 170 190 171
rect 188 170 189 171
rect 187 170 188 171
rect 186 170 187 171
rect 185 170 186 171
rect 184 170 185 171
rect 183 170 184 171
rect 182 170 183 171
rect 181 170 182 171
rect 180 170 181 171
rect 179 170 180 171
rect 178 170 179 171
rect 177 170 178 171
rect 176 170 177 171
rect 175 170 176 171
rect 174 170 175 171
rect 173 170 174 171
rect 172 170 173 171
rect 171 170 172 171
rect 170 170 171 171
rect 169 170 170 171
rect 168 170 169 171
rect 167 170 168 171
rect 166 170 167 171
rect 165 170 166 171
rect 164 170 165 171
rect 163 170 164 171
rect 162 170 163 171
rect 161 170 162 171
rect 160 170 161 171
rect 159 170 160 171
rect 158 170 159 171
rect 157 170 158 171
rect 156 170 157 171
rect 155 170 156 171
rect 154 170 155 171
rect 153 170 154 171
rect 152 170 153 171
rect 151 170 152 171
rect 150 170 151 171
rect 149 170 150 171
rect 148 170 149 171
rect 147 170 148 171
rect 146 170 147 171
rect 145 170 146 171
rect 144 170 145 171
rect 143 170 144 171
rect 142 170 143 171
rect 141 170 142 171
rect 140 170 141 171
rect 139 170 140 171
rect 138 170 139 171
rect 137 170 138 171
rect 136 170 137 171
rect 135 170 136 171
rect 134 170 135 171
rect 133 170 134 171
rect 132 170 133 171
rect 131 170 132 171
rect 130 170 131 171
rect 129 170 130 171
rect 128 170 129 171
rect 56 170 57 171
rect 55 170 56 171
rect 54 170 55 171
rect 53 170 54 171
rect 52 170 53 171
rect 51 170 52 171
rect 50 170 51 171
rect 49 170 50 171
rect 48 170 49 171
rect 47 170 48 171
rect 46 170 47 171
rect 45 170 46 171
rect 44 170 45 171
rect 43 170 44 171
rect 42 170 43 171
rect 41 170 42 171
rect 40 170 41 171
rect 39 170 40 171
rect 38 170 39 171
rect 37 170 38 171
rect 36 170 37 171
rect 35 170 36 171
rect 34 170 35 171
rect 33 170 34 171
rect 32 170 33 171
rect 20 170 21 171
rect 19 170 20 171
rect 18 170 19 171
rect 17 170 18 171
rect 16 170 17 171
rect 15 170 16 171
rect 14 170 15 171
rect 13 170 14 171
rect 12 170 13 171
rect 11 170 12 171
rect 10 170 11 171
rect 9 170 10 171
rect 8 170 9 171
rect 476 171 477 172
rect 475 171 476 172
rect 474 171 475 172
rect 473 171 474 172
rect 472 171 473 172
rect 414 171 415 172
rect 413 171 414 172
rect 412 171 413 172
rect 411 171 412 172
rect 410 171 411 172
rect 409 171 410 172
rect 408 171 409 172
rect 407 171 408 172
rect 406 171 407 172
rect 405 171 406 172
rect 404 171 405 172
rect 403 171 404 172
rect 402 171 403 172
rect 401 171 402 172
rect 400 171 401 172
rect 267 171 268 172
rect 266 171 267 172
rect 265 171 266 172
rect 264 171 265 172
rect 263 171 264 172
rect 262 171 263 172
rect 261 171 262 172
rect 260 171 261 172
rect 259 171 260 172
rect 258 171 259 172
rect 257 171 258 172
rect 256 171 257 172
rect 255 171 256 172
rect 254 171 255 172
rect 253 171 254 172
rect 252 171 253 172
rect 251 171 252 172
rect 250 171 251 172
rect 249 171 250 172
rect 248 171 249 172
rect 247 171 248 172
rect 246 171 247 172
rect 245 171 246 172
rect 244 171 245 172
rect 243 171 244 172
rect 242 171 243 172
rect 241 171 242 172
rect 240 171 241 172
rect 239 171 240 172
rect 238 171 239 172
rect 237 171 238 172
rect 236 171 237 172
rect 235 171 236 172
rect 234 171 235 172
rect 233 171 234 172
rect 232 171 233 172
rect 231 171 232 172
rect 230 171 231 172
rect 229 171 230 172
rect 228 171 229 172
rect 227 171 228 172
rect 226 171 227 172
rect 225 171 226 172
rect 224 171 225 172
rect 205 171 206 172
rect 204 171 205 172
rect 203 171 204 172
rect 202 171 203 172
rect 201 171 202 172
rect 200 171 201 172
rect 199 171 200 172
rect 198 171 199 172
rect 197 171 198 172
rect 196 171 197 172
rect 195 171 196 172
rect 194 171 195 172
rect 193 171 194 172
rect 192 171 193 172
rect 191 171 192 172
rect 190 171 191 172
rect 189 171 190 172
rect 188 171 189 172
rect 187 171 188 172
rect 186 171 187 172
rect 185 171 186 172
rect 184 171 185 172
rect 183 171 184 172
rect 182 171 183 172
rect 181 171 182 172
rect 180 171 181 172
rect 179 171 180 172
rect 178 171 179 172
rect 177 171 178 172
rect 176 171 177 172
rect 175 171 176 172
rect 174 171 175 172
rect 173 171 174 172
rect 172 171 173 172
rect 171 171 172 172
rect 170 171 171 172
rect 169 171 170 172
rect 168 171 169 172
rect 167 171 168 172
rect 166 171 167 172
rect 165 171 166 172
rect 164 171 165 172
rect 163 171 164 172
rect 162 171 163 172
rect 161 171 162 172
rect 160 171 161 172
rect 159 171 160 172
rect 158 171 159 172
rect 157 171 158 172
rect 156 171 157 172
rect 155 171 156 172
rect 154 171 155 172
rect 153 171 154 172
rect 152 171 153 172
rect 151 171 152 172
rect 150 171 151 172
rect 149 171 150 172
rect 148 171 149 172
rect 147 171 148 172
rect 146 171 147 172
rect 145 171 146 172
rect 144 171 145 172
rect 143 171 144 172
rect 142 171 143 172
rect 141 171 142 172
rect 140 171 141 172
rect 139 171 140 172
rect 138 171 139 172
rect 137 171 138 172
rect 136 171 137 172
rect 135 171 136 172
rect 134 171 135 172
rect 133 171 134 172
rect 132 171 133 172
rect 131 171 132 172
rect 130 171 131 172
rect 129 171 130 172
rect 128 171 129 172
rect 127 171 128 172
rect 126 171 127 172
rect 55 171 56 172
rect 54 171 55 172
rect 53 171 54 172
rect 52 171 53 172
rect 51 171 52 172
rect 50 171 51 172
rect 49 171 50 172
rect 48 171 49 172
rect 47 171 48 172
rect 46 171 47 172
rect 45 171 46 172
rect 44 171 45 172
rect 43 171 44 172
rect 42 171 43 172
rect 41 171 42 172
rect 40 171 41 172
rect 39 171 40 172
rect 38 171 39 172
rect 37 171 38 172
rect 36 171 37 172
rect 35 171 36 172
rect 34 171 35 172
rect 33 171 34 172
rect 32 171 33 172
rect 20 171 21 172
rect 19 171 20 172
rect 18 171 19 172
rect 17 171 18 172
rect 16 171 17 172
rect 15 171 16 172
rect 14 171 15 172
rect 13 171 14 172
rect 12 171 13 172
rect 11 171 12 172
rect 10 171 11 172
rect 9 171 10 172
rect 8 171 9 172
rect 473 172 474 173
rect 472 172 473 173
rect 471 172 472 173
rect 470 172 471 173
rect 469 172 470 173
rect 415 172 416 173
rect 414 172 415 173
rect 413 172 414 173
rect 412 172 413 173
rect 411 172 412 173
rect 410 172 411 173
rect 409 172 410 173
rect 408 172 409 173
rect 407 172 408 173
rect 406 172 407 173
rect 405 172 406 173
rect 404 172 405 173
rect 403 172 404 173
rect 402 172 403 173
rect 401 172 402 173
rect 266 172 267 173
rect 265 172 266 173
rect 264 172 265 173
rect 263 172 264 173
rect 262 172 263 173
rect 261 172 262 173
rect 260 172 261 173
rect 259 172 260 173
rect 258 172 259 173
rect 257 172 258 173
rect 256 172 257 173
rect 255 172 256 173
rect 254 172 255 173
rect 253 172 254 173
rect 252 172 253 173
rect 251 172 252 173
rect 250 172 251 173
rect 249 172 250 173
rect 248 172 249 173
rect 247 172 248 173
rect 246 172 247 173
rect 245 172 246 173
rect 244 172 245 173
rect 243 172 244 173
rect 242 172 243 173
rect 241 172 242 173
rect 240 172 241 173
rect 239 172 240 173
rect 238 172 239 173
rect 237 172 238 173
rect 236 172 237 173
rect 235 172 236 173
rect 234 172 235 173
rect 233 172 234 173
rect 232 172 233 173
rect 231 172 232 173
rect 230 172 231 173
rect 229 172 230 173
rect 228 172 229 173
rect 227 172 228 173
rect 226 172 227 173
rect 225 172 226 173
rect 224 172 225 173
rect 223 172 224 173
rect 204 172 205 173
rect 203 172 204 173
rect 202 172 203 173
rect 201 172 202 173
rect 200 172 201 173
rect 199 172 200 173
rect 198 172 199 173
rect 197 172 198 173
rect 196 172 197 173
rect 195 172 196 173
rect 194 172 195 173
rect 193 172 194 173
rect 192 172 193 173
rect 191 172 192 173
rect 190 172 191 173
rect 189 172 190 173
rect 188 172 189 173
rect 187 172 188 173
rect 186 172 187 173
rect 185 172 186 173
rect 184 172 185 173
rect 183 172 184 173
rect 182 172 183 173
rect 181 172 182 173
rect 180 172 181 173
rect 179 172 180 173
rect 178 172 179 173
rect 177 172 178 173
rect 176 172 177 173
rect 175 172 176 173
rect 174 172 175 173
rect 173 172 174 173
rect 172 172 173 173
rect 171 172 172 173
rect 170 172 171 173
rect 169 172 170 173
rect 168 172 169 173
rect 167 172 168 173
rect 166 172 167 173
rect 165 172 166 173
rect 164 172 165 173
rect 163 172 164 173
rect 162 172 163 173
rect 161 172 162 173
rect 160 172 161 173
rect 159 172 160 173
rect 158 172 159 173
rect 157 172 158 173
rect 156 172 157 173
rect 155 172 156 173
rect 154 172 155 173
rect 153 172 154 173
rect 152 172 153 173
rect 151 172 152 173
rect 150 172 151 173
rect 149 172 150 173
rect 148 172 149 173
rect 147 172 148 173
rect 146 172 147 173
rect 145 172 146 173
rect 144 172 145 173
rect 143 172 144 173
rect 142 172 143 173
rect 141 172 142 173
rect 140 172 141 173
rect 139 172 140 173
rect 138 172 139 173
rect 137 172 138 173
rect 136 172 137 173
rect 135 172 136 173
rect 134 172 135 173
rect 133 172 134 173
rect 132 172 133 173
rect 131 172 132 173
rect 130 172 131 173
rect 129 172 130 173
rect 128 172 129 173
rect 127 172 128 173
rect 126 172 127 173
rect 125 172 126 173
rect 55 172 56 173
rect 54 172 55 173
rect 53 172 54 173
rect 52 172 53 173
rect 51 172 52 173
rect 50 172 51 173
rect 49 172 50 173
rect 48 172 49 173
rect 47 172 48 173
rect 46 172 47 173
rect 45 172 46 173
rect 44 172 45 173
rect 43 172 44 173
rect 42 172 43 173
rect 41 172 42 173
rect 40 172 41 173
rect 39 172 40 173
rect 38 172 39 173
rect 37 172 38 173
rect 36 172 37 173
rect 35 172 36 173
rect 34 172 35 173
rect 33 172 34 173
rect 20 172 21 173
rect 19 172 20 173
rect 18 172 19 173
rect 17 172 18 173
rect 16 172 17 173
rect 15 172 16 173
rect 14 172 15 173
rect 13 172 14 173
rect 12 172 13 173
rect 11 172 12 173
rect 10 172 11 173
rect 9 172 10 173
rect 471 173 472 174
rect 470 173 471 174
rect 469 173 470 174
rect 468 173 469 174
rect 467 173 468 174
rect 458 173 459 174
rect 416 173 417 174
rect 415 173 416 174
rect 414 173 415 174
rect 413 173 414 174
rect 412 173 413 174
rect 411 173 412 174
rect 410 173 411 174
rect 409 173 410 174
rect 408 173 409 174
rect 407 173 408 174
rect 406 173 407 174
rect 405 173 406 174
rect 404 173 405 174
rect 403 173 404 174
rect 265 173 266 174
rect 264 173 265 174
rect 263 173 264 174
rect 262 173 263 174
rect 261 173 262 174
rect 260 173 261 174
rect 259 173 260 174
rect 258 173 259 174
rect 257 173 258 174
rect 256 173 257 174
rect 255 173 256 174
rect 254 173 255 174
rect 253 173 254 174
rect 252 173 253 174
rect 251 173 252 174
rect 250 173 251 174
rect 249 173 250 174
rect 248 173 249 174
rect 247 173 248 174
rect 246 173 247 174
rect 245 173 246 174
rect 244 173 245 174
rect 243 173 244 174
rect 242 173 243 174
rect 241 173 242 174
rect 240 173 241 174
rect 239 173 240 174
rect 238 173 239 174
rect 237 173 238 174
rect 236 173 237 174
rect 235 173 236 174
rect 234 173 235 174
rect 233 173 234 174
rect 232 173 233 174
rect 231 173 232 174
rect 230 173 231 174
rect 229 173 230 174
rect 228 173 229 174
rect 227 173 228 174
rect 226 173 227 174
rect 225 173 226 174
rect 224 173 225 174
rect 223 173 224 174
rect 204 173 205 174
rect 203 173 204 174
rect 202 173 203 174
rect 201 173 202 174
rect 200 173 201 174
rect 199 173 200 174
rect 198 173 199 174
rect 197 173 198 174
rect 196 173 197 174
rect 195 173 196 174
rect 194 173 195 174
rect 193 173 194 174
rect 192 173 193 174
rect 191 173 192 174
rect 190 173 191 174
rect 189 173 190 174
rect 188 173 189 174
rect 187 173 188 174
rect 186 173 187 174
rect 185 173 186 174
rect 184 173 185 174
rect 183 173 184 174
rect 182 173 183 174
rect 181 173 182 174
rect 180 173 181 174
rect 179 173 180 174
rect 178 173 179 174
rect 177 173 178 174
rect 176 173 177 174
rect 175 173 176 174
rect 174 173 175 174
rect 173 173 174 174
rect 172 173 173 174
rect 171 173 172 174
rect 170 173 171 174
rect 169 173 170 174
rect 168 173 169 174
rect 167 173 168 174
rect 166 173 167 174
rect 165 173 166 174
rect 164 173 165 174
rect 163 173 164 174
rect 162 173 163 174
rect 161 173 162 174
rect 160 173 161 174
rect 159 173 160 174
rect 158 173 159 174
rect 157 173 158 174
rect 156 173 157 174
rect 155 173 156 174
rect 154 173 155 174
rect 153 173 154 174
rect 152 173 153 174
rect 151 173 152 174
rect 150 173 151 174
rect 149 173 150 174
rect 148 173 149 174
rect 147 173 148 174
rect 146 173 147 174
rect 145 173 146 174
rect 144 173 145 174
rect 143 173 144 174
rect 142 173 143 174
rect 141 173 142 174
rect 140 173 141 174
rect 139 173 140 174
rect 138 173 139 174
rect 137 173 138 174
rect 136 173 137 174
rect 135 173 136 174
rect 134 173 135 174
rect 133 173 134 174
rect 132 173 133 174
rect 131 173 132 174
rect 130 173 131 174
rect 129 173 130 174
rect 128 173 129 174
rect 127 173 128 174
rect 126 173 127 174
rect 125 173 126 174
rect 124 173 125 174
rect 123 173 124 174
rect 54 173 55 174
rect 53 173 54 174
rect 52 173 53 174
rect 51 173 52 174
rect 50 173 51 174
rect 49 173 50 174
rect 48 173 49 174
rect 47 173 48 174
rect 46 173 47 174
rect 45 173 46 174
rect 44 173 45 174
rect 43 173 44 174
rect 42 173 43 174
rect 41 173 42 174
rect 40 173 41 174
rect 39 173 40 174
rect 38 173 39 174
rect 37 173 38 174
rect 36 173 37 174
rect 35 173 36 174
rect 34 173 35 174
rect 33 173 34 174
rect 21 173 22 174
rect 20 173 21 174
rect 19 173 20 174
rect 18 173 19 174
rect 17 173 18 174
rect 16 173 17 174
rect 15 173 16 174
rect 14 173 15 174
rect 13 173 14 174
rect 12 173 13 174
rect 11 173 12 174
rect 10 173 11 174
rect 9 173 10 174
rect 468 174 469 175
rect 467 174 468 175
rect 466 174 467 175
rect 465 174 466 175
rect 464 174 465 175
rect 458 174 459 175
rect 417 174 418 175
rect 416 174 417 175
rect 415 174 416 175
rect 414 174 415 175
rect 413 174 414 175
rect 412 174 413 175
rect 411 174 412 175
rect 410 174 411 175
rect 409 174 410 175
rect 408 174 409 175
rect 407 174 408 175
rect 406 174 407 175
rect 405 174 406 175
rect 404 174 405 175
rect 264 174 265 175
rect 263 174 264 175
rect 262 174 263 175
rect 261 174 262 175
rect 260 174 261 175
rect 259 174 260 175
rect 258 174 259 175
rect 257 174 258 175
rect 256 174 257 175
rect 255 174 256 175
rect 254 174 255 175
rect 253 174 254 175
rect 252 174 253 175
rect 251 174 252 175
rect 250 174 251 175
rect 249 174 250 175
rect 248 174 249 175
rect 247 174 248 175
rect 246 174 247 175
rect 245 174 246 175
rect 244 174 245 175
rect 243 174 244 175
rect 242 174 243 175
rect 241 174 242 175
rect 240 174 241 175
rect 239 174 240 175
rect 238 174 239 175
rect 237 174 238 175
rect 236 174 237 175
rect 235 174 236 175
rect 234 174 235 175
rect 233 174 234 175
rect 232 174 233 175
rect 231 174 232 175
rect 230 174 231 175
rect 229 174 230 175
rect 228 174 229 175
rect 227 174 228 175
rect 226 174 227 175
rect 225 174 226 175
rect 224 174 225 175
rect 223 174 224 175
rect 222 174 223 175
rect 203 174 204 175
rect 202 174 203 175
rect 201 174 202 175
rect 200 174 201 175
rect 199 174 200 175
rect 198 174 199 175
rect 197 174 198 175
rect 196 174 197 175
rect 195 174 196 175
rect 194 174 195 175
rect 193 174 194 175
rect 192 174 193 175
rect 191 174 192 175
rect 190 174 191 175
rect 189 174 190 175
rect 188 174 189 175
rect 187 174 188 175
rect 186 174 187 175
rect 185 174 186 175
rect 184 174 185 175
rect 183 174 184 175
rect 182 174 183 175
rect 181 174 182 175
rect 180 174 181 175
rect 179 174 180 175
rect 178 174 179 175
rect 177 174 178 175
rect 176 174 177 175
rect 175 174 176 175
rect 174 174 175 175
rect 173 174 174 175
rect 172 174 173 175
rect 171 174 172 175
rect 170 174 171 175
rect 169 174 170 175
rect 168 174 169 175
rect 167 174 168 175
rect 166 174 167 175
rect 165 174 166 175
rect 164 174 165 175
rect 163 174 164 175
rect 162 174 163 175
rect 161 174 162 175
rect 160 174 161 175
rect 159 174 160 175
rect 158 174 159 175
rect 157 174 158 175
rect 156 174 157 175
rect 155 174 156 175
rect 154 174 155 175
rect 153 174 154 175
rect 152 174 153 175
rect 151 174 152 175
rect 150 174 151 175
rect 149 174 150 175
rect 148 174 149 175
rect 147 174 148 175
rect 146 174 147 175
rect 145 174 146 175
rect 144 174 145 175
rect 143 174 144 175
rect 142 174 143 175
rect 141 174 142 175
rect 140 174 141 175
rect 139 174 140 175
rect 138 174 139 175
rect 137 174 138 175
rect 136 174 137 175
rect 135 174 136 175
rect 134 174 135 175
rect 133 174 134 175
rect 132 174 133 175
rect 131 174 132 175
rect 130 174 131 175
rect 129 174 130 175
rect 128 174 129 175
rect 127 174 128 175
rect 126 174 127 175
rect 125 174 126 175
rect 124 174 125 175
rect 123 174 124 175
rect 122 174 123 175
rect 121 174 122 175
rect 53 174 54 175
rect 52 174 53 175
rect 51 174 52 175
rect 50 174 51 175
rect 49 174 50 175
rect 48 174 49 175
rect 47 174 48 175
rect 46 174 47 175
rect 45 174 46 175
rect 44 174 45 175
rect 43 174 44 175
rect 42 174 43 175
rect 41 174 42 175
rect 40 174 41 175
rect 39 174 40 175
rect 38 174 39 175
rect 37 174 38 175
rect 36 174 37 175
rect 35 174 36 175
rect 34 174 35 175
rect 21 174 22 175
rect 20 174 21 175
rect 19 174 20 175
rect 18 174 19 175
rect 17 174 18 175
rect 16 174 17 175
rect 15 174 16 175
rect 14 174 15 175
rect 13 174 14 175
rect 12 174 13 175
rect 11 174 12 175
rect 10 174 11 175
rect 9 174 10 175
rect 465 175 466 176
rect 464 175 465 176
rect 463 175 464 176
rect 462 175 463 176
rect 461 175 462 176
rect 460 175 461 176
rect 459 175 460 176
rect 458 175 459 176
rect 418 175 419 176
rect 417 175 418 176
rect 416 175 417 176
rect 415 175 416 176
rect 414 175 415 176
rect 413 175 414 176
rect 412 175 413 176
rect 411 175 412 176
rect 410 175 411 176
rect 409 175 410 176
rect 408 175 409 176
rect 407 175 408 176
rect 406 175 407 176
rect 405 175 406 176
rect 263 175 264 176
rect 262 175 263 176
rect 261 175 262 176
rect 260 175 261 176
rect 259 175 260 176
rect 258 175 259 176
rect 257 175 258 176
rect 256 175 257 176
rect 255 175 256 176
rect 254 175 255 176
rect 253 175 254 176
rect 252 175 253 176
rect 251 175 252 176
rect 250 175 251 176
rect 249 175 250 176
rect 248 175 249 176
rect 247 175 248 176
rect 246 175 247 176
rect 245 175 246 176
rect 244 175 245 176
rect 243 175 244 176
rect 242 175 243 176
rect 241 175 242 176
rect 240 175 241 176
rect 239 175 240 176
rect 238 175 239 176
rect 237 175 238 176
rect 236 175 237 176
rect 235 175 236 176
rect 234 175 235 176
rect 233 175 234 176
rect 232 175 233 176
rect 231 175 232 176
rect 230 175 231 176
rect 229 175 230 176
rect 228 175 229 176
rect 227 175 228 176
rect 226 175 227 176
rect 225 175 226 176
rect 224 175 225 176
rect 223 175 224 176
rect 222 175 223 176
rect 202 175 203 176
rect 201 175 202 176
rect 200 175 201 176
rect 199 175 200 176
rect 198 175 199 176
rect 197 175 198 176
rect 196 175 197 176
rect 195 175 196 176
rect 194 175 195 176
rect 193 175 194 176
rect 192 175 193 176
rect 191 175 192 176
rect 190 175 191 176
rect 189 175 190 176
rect 188 175 189 176
rect 187 175 188 176
rect 186 175 187 176
rect 185 175 186 176
rect 184 175 185 176
rect 183 175 184 176
rect 182 175 183 176
rect 181 175 182 176
rect 180 175 181 176
rect 179 175 180 176
rect 178 175 179 176
rect 177 175 178 176
rect 176 175 177 176
rect 175 175 176 176
rect 174 175 175 176
rect 173 175 174 176
rect 172 175 173 176
rect 171 175 172 176
rect 170 175 171 176
rect 169 175 170 176
rect 168 175 169 176
rect 167 175 168 176
rect 166 175 167 176
rect 165 175 166 176
rect 164 175 165 176
rect 163 175 164 176
rect 162 175 163 176
rect 161 175 162 176
rect 160 175 161 176
rect 159 175 160 176
rect 158 175 159 176
rect 157 175 158 176
rect 156 175 157 176
rect 155 175 156 176
rect 154 175 155 176
rect 153 175 154 176
rect 152 175 153 176
rect 151 175 152 176
rect 150 175 151 176
rect 149 175 150 176
rect 148 175 149 176
rect 147 175 148 176
rect 146 175 147 176
rect 145 175 146 176
rect 144 175 145 176
rect 143 175 144 176
rect 142 175 143 176
rect 141 175 142 176
rect 140 175 141 176
rect 139 175 140 176
rect 138 175 139 176
rect 137 175 138 176
rect 136 175 137 176
rect 135 175 136 176
rect 134 175 135 176
rect 133 175 134 176
rect 132 175 133 176
rect 131 175 132 176
rect 130 175 131 176
rect 129 175 130 176
rect 128 175 129 176
rect 127 175 128 176
rect 126 175 127 176
rect 125 175 126 176
rect 124 175 125 176
rect 123 175 124 176
rect 122 175 123 176
rect 121 175 122 176
rect 120 175 121 176
rect 119 175 120 176
rect 52 175 53 176
rect 51 175 52 176
rect 50 175 51 176
rect 49 175 50 176
rect 48 175 49 176
rect 47 175 48 176
rect 46 175 47 176
rect 45 175 46 176
rect 44 175 45 176
rect 43 175 44 176
rect 42 175 43 176
rect 41 175 42 176
rect 40 175 41 176
rect 39 175 40 176
rect 38 175 39 176
rect 37 175 38 176
rect 36 175 37 176
rect 35 175 36 176
rect 34 175 35 176
rect 21 175 22 176
rect 20 175 21 176
rect 19 175 20 176
rect 18 175 19 176
rect 17 175 18 176
rect 16 175 17 176
rect 15 175 16 176
rect 14 175 15 176
rect 13 175 14 176
rect 12 175 13 176
rect 11 175 12 176
rect 10 175 11 176
rect 9 175 10 176
rect 463 176 464 177
rect 462 176 463 177
rect 461 176 462 177
rect 460 176 461 177
rect 459 176 460 177
rect 458 176 459 177
rect 420 176 421 177
rect 419 176 420 177
rect 418 176 419 177
rect 417 176 418 177
rect 416 176 417 177
rect 415 176 416 177
rect 414 176 415 177
rect 413 176 414 177
rect 412 176 413 177
rect 411 176 412 177
rect 410 176 411 177
rect 409 176 410 177
rect 408 176 409 177
rect 407 176 408 177
rect 406 176 407 177
rect 263 176 264 177
rect 262 176 263 177
rect 261 176 262 177
rect 260 176 261 177
rect 259 176 260 177
rect 258 176 259 177
rect 257 176 258 177
rect 256 176 257 177
rect 255 176 256 177
rect 254 176 255 177
rect 253 176 254 177
rect 252 176 253 177
rect 251 176 252 177
rect 250 176 251 177
rect 249 176 250 177
rect 248 176 249 177
rect 247 176 248 177
rect 246 176 247 177
rect 245 176 246 177
rect 244 176 245 177
rect 243 176 244 177
rect 242 176 243 177
rect 241 176 242 177
rect 240 176 241 177
rect 239 176 240 177
rect 238 176 239 177
rect 237 176 238 177
rect 236 176 237 177
rect 235 176 236 177
rect 234 176 235 177
rect 233 176 234 177
rect 232 176 233 177
rect 231 176 232 177
rect 230 176 231 177
rect 229 176 230 177
rect 228 176 229 177
rect 227 176 228 177
rect 226 176 227 177
rect 225 176 226 177
rect 224 176 225 177
rect 223 176 224 177
rect 222 176 223 177
rect 221 176 222 177
rect 202 176 203 177
rect 201 176 202 177
rect 200 176 201 177
rect 199 176 200 177
rect 198 176 199 177
rect 197 176 198 177
rect 196 176 197 177
rect 195 176 196 177
rect 194 176 195 177
rect 193 176 194 177
rect 192 176 193 177
rect 191 176 192 177
rect 190 176 191 177
rect 189 176 190 177
rect 188 176 189 177
rect 187 176 188 177
rect 186 176 187 177
rect 185 176 186 177
rect 184 176 185 177
rect 183 176 184 177
rect 182 176 183 177
rect 181 176 182 177
rect 180 176 181 177
rect 179 176 180 177
rect 178 176 179 177
rect 177 176 178 177
rect 176 176 177 177
rect 175 176 176 177
rect 174 176 175 177
rect 173 176 174 177
rect 172 176 173 177
rect 171 176 172 177
rect 170 176 171 177
rect 169 176 170 177
rect 168 176 169 177
rect 167 176 168 177
rect 166 176 167 177
rect 165 176 166 177
rect 164 176 165 177
rect 163 176 164 177
rect 162 176 163 177
rect 161 176 162 177
rect 160 176 161 177
rect 159 176 160 177
rect 158 176 159 177
rect 157 176 158 177
rect 156 176 157 177
rect 155 176 156 177
rect 154 176 155 177
rect 153 176 154 177
rect 152 176 153 177
rect 151 176 152 177
rect 150 176 151 177
rect 149 176 150 177
rect 148 176 149 177
rect 147 176 148 177
rect 146 176 147 177
rect 145 176 146 177
rect 144 176 145 177
rect 143 176 144 177
rect 142 176 143 177
rect 141 176 142 177
rect 140 176 141 177
rect 139 176 140 177
rect 138 176 139 177
rect 137 176 138 177
rect 136 176 137 177
rect 135 176 136 177
rect 134 176 135 177
rect 133 176 134 177
rect 132 176 133 177
rect 131 176 132 177
rect 130 176 131 177
rect 129 176 130 177
rect 128 176 129 177
rect 127 176 128 177
rect 126 176 127 177
rect 125 176 126 177
rect 124 176 125 177
rect 123 176 124 177
rect 122 176 123 177
rect 121 176 122 177
rect 120 176 121 177
rect 119 176 120 177
rect 118 176 119 177
rect 117 176 118 177
rect 116 176 117 177
rect 51 176 52 177
rect 50 176 51 177
rect 49 176 50 177
rect 48 176 49 177
rect 47 176 48 177
rect 46 176 47 177
rect 45 176 46 177
rect 44 176 45 177
rect 43 176 44 177
rect 42 176 43 177
rect 41 176 42 177
rect 40 176 41 177
rect 39 176 40 177
rect 38 176 39 177
rect 37 176 38 177
rect 36 176 37 177
rect 35 176 36 177
rect 21 176 22 177
rect 20 176 21 177
rect 19 176 20 177
rect 18 176 19 177
rect 17 176 18 177
rect 16 176 17 177
rect 15 176 16 177
rect 14 176 15 177
rect 13 176 14 177
rect 12 176 13 177
rect 11 176 12 177
rect 10 176 11 177
rect 9 176 10 177
rect 461 177 462 178
rect 460 177 461 178
rect 459 177 460 178
rect 458 177 459 178
rect 421 177 422 178
rect 420 177 421 178
rect 419 177 420 178
rect 418 177 419 178
rect 417 177 418 178
rect 416 177 417 178
rect 415 177 416 178
rect 414 177 415 178
rect 413 177 414 178
rect 412 177 413 178
rect 411 177 412 178
rect 410 177 411 178
rect 409 177 410 178
rect 408 177 409 178
rect 407 177 408 178
rect 262 177 263 178
rect 261 177 262 178
rect 260 177 261 178
rect 259 177 260 178
rect 258 177 259 178
rect 257 177 258 178
rect 256 177 257 178
rect 255 177 256 178
rect 254 177 255 178
rect 253 177 254 178
rect 252 177 253 178
rect 251 177 252 178
rect 250 177 251 178
rect 249 177 250 178
rect 248 177 249 178
rect 247 177 248 178
rect 246 177 247 178
rect 245 177 246 178
rect 244 177 245 178
rect 243 177 244 178
rect 242 177 243 178
rect 241 177 242 178
rect 240 177 241 178
rect 239 177 240 178
rect 238 177 239 178
rect 237 177 238 178
rect 236 177 237 178
rect 235 177 236 178
rect 234 177 235 178
rect 233 177 234 178
rect 232 177 233 178
rect 231 177 232 178
rect 230 177 231 178
rect 229 177 230 178
rect 228 177 229 178
rect 227 177 228 178
rect 226 177 227 178
rect 225 177 226 178
rect 224 177 225 178
rect 223 177 224 178
rect 222 177 223 178
rect 221 177 222 178
rect 201 177 202 178
rect 200 177 201 178
rect 199 177 200 178
rect 198 177 199 178
rect 197 177 198 178
rect 196 177 197 178
rect 195 177 196 178
rect 194 177 195 178
rect 193 177 194 178
rect 192 177 193 178
rect 191 177 192 178
rect 190 177 191 178
rect 189 177 190 178
rect 188 177 189 178
rect 187 177 188 178
rect 186 177 187 178
rect 185 177 186 178
rect 184 177 185 178
rect 183 177 184 178
rect 182 177 183 178
rect 181 177 182 178
rect 180 177 181 178
rect 179 177 180 178
rect 178 177 179 178
rect 177 177 178 178
rect 176 177 177 178
rect 175 177 176 178
rect 174 177 175 178
rect 173 177 174 178
rect 172 177 173 178
rect 171 177 172 178
rect 170 177 171 178
rect 169 177 170 178
rect 168 177 169 178
rect 167 177 168 178
rect 166 177 167 178
rect 165 177 166 178
rect 164 177 165 178
rect 163 177 164 178
rect 162 177 163 178
rect 161 177 162 178
rect 160 177 161 178
rect 159 177 160 178
rect 158 177 159 178
rect 157 177 158 178
rect 156 177 157 178
rect 155 177 156 178
rect 154 177 155 178
rect 153 177 154 178
rect 152 177 153 178
rect 151 177 152 178
rect 150 177 151 178
rect 149 177 150 178
rect 148 177 149 178
rect 147 177 148 178
rect 146 177 147 178
rect 145 177 146 178
rect 144 177 145 178
rect 143 177 144 178
rect 142 177 143 178
rect 141 177 142 178
rect 140 177 141 178
rect 139 177 140 178
rect 138 177 139 178
rect 137 177 138 178
rect 136 177 137 178
rect 135 177 136 178
rect 134 177 135 178
rect 133 177 134 178
rect 132 177 133 178
rect 131 177 132 178
rect 130 177 131 178
rect 129 177 130 178
rect 128 177 129 178
rect 127 177 128 178
rect 126 177 127 178
rect 125 177 126 178
rect 124 177 125 178
rect 123 177 124 178
rect 122 177 123 178
rect 121 177 122 178
rect 120 177 121 178
rect 119 177 120 178
rect 118 177 119 178
rect 117 177 118 178
rect 116 177 117 178
rect 115 177 116 178
rect 114 177 115 178
rect 50 177 51 178
rect 49 177 50 178
rect 48 177 49 178
rect 47 177 48 178
rect 46 177 47 178
rect 45 177 46 178
rect 44 177 45 178
rect 43 177 44 178
rect 42 177 43 178
rect 41 177 42 178
rect 40 177 41 178
rect 39 177 40 178
rect 38 177 39 178
rect 37 177 38 178
rect 36 177 37 178
rect 21 177 22 178
rect 20 177 21 178
rect 19 177 20 178
rect 18 177 19 178
rect 17 177 18 178
rect 16 177 17 178
rect 15 177 16 178
rect 14 177 15 178
rect 13 177 14 178
rect 12 177 13 178
rect 11 177 12 178
rect 10 177 11 178
rect 459 178 460 179
rect 458 178 459 179
rect 422 178 423 179
rect 421 178 422 179
rect 420 178 421 179
rect 419 178 420 179
rect 418 178 419 179
rect 417 178 418 179
rect 416 178 417 179
rect 415 178 416 179
rect 414 178 415 179
rect 413 178 414 179
rect 412 178 413 179
rect 411 178 412 179
rect 410 178 411 179
rect 409 178 410 179
rect 408 178 409 179
rect 315 178 316 179
rect 314 178 315 179
rect 313 178 314 179
rect 312 178 313 179
rect 311 178 312 179
rect 310 178 311 179
rect 309 178 310 179
rect 308 178 309 179
rect 307 178 308 179
rect 306 178 307 179
rect 305 178 306 179
rect 304 178 305 179
rect 303 178 304 179
rect 302 178 303 179
rect 301 178 302 179
rect 300 178 301 179
rect 299 178 300 179
rect 261 178 262 179
rect 260 178 261 179
rect 259 178 260 179
rect 258 178 259 179
rect 257 178 258 179
rect 256 178 257 179
rect 255 178 256 179
rect 254 178 255 179
rect 253 178 254 179
rect 252 178 253 179
rect 251 178 252 179
rect 250 178 251 179
rect 249 178 250 179
rect 248 178 249 179
rect 247 178 248 179
rect 246 178 247 179
rect 245 178 246 179
rect 244 178 245 179
rect 243 178 244 179
rect 242 178 243 179
rect 241 178 242 179
rect 240 178 241 179
rect 239 178 240 179
rect 238 178 239 179
rect 237 178 238 179
rect 236 178 237 179
rect 235 178 236 179
rect 234 178 235 179
rect 233 178 234 179
rect 232 178 233 179
rect 231 178 232 179
rect 230 178 231 179
rect 229 178 230 179
rect 228 178 229 179
rect 227 178 228 179
rect 226 178 227 179
rect 225 178 226 179
rect 224 178 225 179
rect 223 178 224 179
rect 222 178 223 179
rect 221 178 222 179
rect 220 178 221 179
rect 200 178 201 179
rect 199 178 200 179
rect 198 178 199 179
rect 197 178 198 179
rect 196 178 197 179
rect 195 178 196 179
rect 194 178 195 179
rect 193 178 194 179
rect 192 178 193 179
rect 191 178 192 179
rect 190 178 191 179
rect 189 178 190 179
rect 188 178 189 179
rect 187 178 188 179
rect 186 178 187 179
rect 185 178 186 179
rect 184 178 185 179
rect 183 178 184 179
rect 182 178 183 179
rect 181 178 182 179
rect 180 178 181 179
rect 179 178 180 179
rect 178 178 179 179
rect 177 178 178 179
rect 176 178 177 179
rect 175 178 176 179
rect 174 178 175 179
rect 173 178 174 179
rect 172 178 173 179
rect 171 178 172 179
rect 170 178 171 179
rect 169 178 170 179
rect 168 178 169 179
rect 167 178 168 179
rect 166 178 167 179
rect 165 178 166 179
rect 164 178 165 179
rect 163 178 164 179
rect 162 178 163 179
rect 161 178 162 179
rect 160 178 161 179
rect 159 178 160 179
rect 158 178 159 179
rect 157 178 158 179
rect 156 178 157 179
rect 155 178 156 179
rect 154 178 155 179
rect 153 178 154 179
rect 152 178 153 179
rect 151 178 152 179
rect 150 178 151 179
rect 149 178 150 179
rect 148 178 149 179
rect 147 178 148 179
rect 146 178 147 179
rect 145 178 146 179
rect 144 178 145 179
rect 143 178 144 179
rect 142 178 143 179
rect 141 178 142 179
rect 140 178 141 179
rect 139 178 140 179
rect 138 178 139 179
rect 137 178 138 179
rect 136 178 137 179
rect 135 178 136 179
rect 134 178 135 179
rect 133 178 134 179
rect 132 178 133 179
rect 131 178 132 179
rect 130 178 131 179
rect 129 178 130 179
rect 128 178 129 179
rect 127 178 128 179
rect 126 178 127 179
rect 125 178 126 179
rect 124 178 125 179
rect 123 178 124 179
rect 122 178 123 179
rect 121 178 122 179
rect 120 178 121 179
rect 119 178 120 179
rect 118 178 119 179
rect 117 178 118 179
rect 116 178 117 179
rect 115 178 116 179
rect 114 178 115 179
rect 113 178 114 179
rect 112 178 113 179
rect 111 178 112 179
rect 68 178 69 179
rect 67 178 68 179
rect 48 178 49 179
rect 47 178 48 179
rect 46 178 47 179
rect 45 178 46 179
rect 44 178 45 179
rect 43 178 44 179
rect 42 178 43 179
rect 41 178 42 179
rect 40 178 41 179
rect 39 178 40 179
rect 38 178 39 179
rect 37 178 38 179
rect 21 178 22 179
rect 20 178 21 179
rect 19 178 20 179
rect 18 178 19 179
rect 17 178 18 179
rect 16 178 17 179
rect 15 178 16 179
rect 14 178 15 179
rect 13 178 14 179
rect 12 178 13 179
rect 11 178 12 179
rect 10 178 11 179
rect 458 179 459 180
rect 423 179 424 180
rect 422 179 423 180
rect 421 179 422 180
rect 420 179 421 180
rect 419 179 420 180
rect 418 179 419 180
rect 417 179 418 180
rect 416 179 417 180
rect 415 179 416 180
rect 414 179 415 180
rect 413 179 414 180
rect 412 179 413 180
rect 411 179 412 180
rect 410 179 411 180
rect 409 179 410 180
rect 320 179 321 180
rect 319 179 320 180
rect 318 179 319 180
rect 317 179 318 180
rect 316 179 317 180
rect 315 179 316 180
rect 314 179 315 180
rect 313 179 314 180
rect 312 179 313 180
rect 311 179 312 180
rect 310 179 311 180
rect 309 179 310 180
rect 308 179 309 180
rect 307 179 308 180
rect 306 179 307 180
rect 305 179 306 180
rect 304 179 305 180
rect 303 179 304 180
rect 302 179 303 180
rect 301 179 302 180
rect 300 179 301 180
rect 299 179 300 180
rect 298 179 299 180
rect 297 179 298 180
rect 296 179 297 180
rect 295 179 296 180
rect 294 179 295 180
rect 260 179 261 180
rect 259 179 260 180
rect 258 179 259 180
rect 257 179 258 180
rect 256 179 257 180
rect 255 179 256 180
rect 254 179 255 180
rect 253 179 254 180
rect 252 179 253 180
rect 251 179 252 180
rect 250 179 251 180
rect 249 179 250 180
rect 248 179 249 180
rect 247 179 248 180
rect 246 179 247 180
rect 245 179 246 180
rect 244 179 245 180
rect 243 179 244 180
rect 242 179 243 180
rect 241 179 242 180
rect 240 179 241 180
rect 239 179 240 180
rect 238 179 239 180
rect 237 179 238 180
rect 236 179 237 180
rect 235 179 236 180
rect 234 179 235 180
rect 233 179 234 180
rect 232 179 233 180
rect 231 179 232 180
rect 230 179 231 180
rect 229 179 230 180
rect 228 179 229 180
rect 227 179 228 180
rect 226 179 227 180
rect 225 179 226 180
rect 224 179 225 180
rect 223 179 224 180
rect 222 179 223 180
rect 221 179 222 180
rect 220 179 221 180
rect 199 179 200 180
rect 198 179 199 180
rect 197 179 198 180
rect 196 179 197 180
rect 195 179 196 180
rect 194 179 195 180
rect 193 179 194 180
rect 192 179 193 180
rect 191 179 192 180
rect 190 179 191 180
rect 189 179 190 180
rect 188 179 189 180
rect 187 179 188 180
rect 186 179 187 180
rect 185 179 186 180
rect 184 179 185 180
rect 183 179 184 180
rect 182 179 183 180
rect 181 179 182 180
rect 180 179 181 180
rect 179 179 180 180
rect 178 179 179 180
rect 177 179 178 180
rect 176 179 177 180
rect 175 179 176 180
rect 174 179 175 180
rect 173 179 174 180
rect 172 179 173 180
rect 171 179 172 180
rect 170 179 171 180
rect 169 179 170 180
rect 168 179 169 180
rect 167 179 168 180
rect 166 179 167 180
rect 165 179 166 180
rect 164 179 165 180
rect 163 179 164 180
rect 162 179 163 180
rect 161 179 162 180
rect 160 179 161 180
rect 159 179 160 180
rect 158 179 159 180
rect 157 179 158 180
rect 156 179 157 180
rect 155 179 156 180
rect 154 179 155 180
rect 153 179 154 180
rect 152 179 153 180
rect 151 179 152 180
rect 150 179 151 180
rect 149 179 150 180
rect 148 179 149 180
rect 147 179 148 180
rect 146 179 147 180
rect 145 179 146 180
rect 144 179 145 180
rect 143 179 144 180
rect 142 179 143 180
rect 141 179 142 180
rect 140 179 141 180
rect 139 179 140 180
rect 138 179 139 180
rect 137 179 138 180
rect 136 179 137 180
rect 135 179 136 180
rect 134 179 135 180
rect 133 179 134 180
rect 132 179 133 180
rect 131 179 132 180
rect 130 179 131 180
rect 129 179 130 180
rect 128 179 129 180
rect 127 179 128 180
rect 126 179 127 180
rect 125 179 126 180
rect 124 179 125 180
rect 123 179 124 180
rect 122 179 123 180
rect 121 179 122 180
rect 120 179 121 180
rect 119 179 120 180
rect 118 179 119 180
rect 117 179 118 180
rect 116 179 117 180
rect 115 179 116 180
rect 114 179 115 180
rect 113 179 114 180
rect 112 179 113 180
rect 111 179 112 180
rect 110 179 111 180
rect 109 179 110 180
rect 70 179 71 180
rect 69 179 70 180
rect 68 179 69 180
rect 67 179 68 180
rect 46 179 47 180
rect 45 179 46 180
rect 44 179 45 180
rect 43 179 44 180
rect 42 179 43 180
rect 41 179 42 180
rect 40 179 41 180
rect 39 179 40 180
rect 21 179 22 180
rect 20 179 21 180
rect 19 179 20 180
rect 18 179 19 180
rect 17 179 18 180
rect 16 179 17 180
rect 15 179 16 180
rect 14 179 15 180
rect 13 179 14 180
rect 12 179 13 180
rect 11 179 12 180
rect 10 179 11 180
rect 458 180 459 181
rect 424 180 425 181
rect 423 180 424 181
rect 422 180 423 181
rect 421 180 422 181
rect 420 180 421 181
rect 419 180 420 181
rect 418 180 419 181
rect 417 180 418 181
rect 416 180 417 181
rect 415 180 416 181
rect 414 180 415 181
rect 413 180 414 181
rect 412 180 413 181
rect 411 180 412 181
rect 323 180 324 181
rect 322 180 323 181
rect 321 180 322 181
rect 320 180 321 181
rect 319 180 320 181
rect 318 180 319 181
rect 317 180 318 181
rect 316 180 317 181
rect 315 180 316 181
rect 314 180 315 181
rect 313 180 314 181
rect 312 180 313 181
rect 311 180 312 181
rect 310 180 311 181
rect 309 180 310 181
rect 308 180 309 181
rect 307 180 308 181
rect 306 180 307 181
rect 305 180 306 181
rect 304 180 305 181
rect 303 180 304 181
rect 302 180 303 181
rect 301 180 302 181
rect 300 180 301 181
rect 299 180 300 181
rect 298 180 299 181
rect 297 180 298 181
rect 296 180 297 181
rect 295 180 296 181
rect 294 180 295 181
rect 293 180 294 181
rect 292 180 293 181
rect 291 180 292 181
rect 290 180 291 181
rect 259 180 260 181
rect 258 180 259 181
rect 257 180 258 181
rect 256 180 257 181
rect 255 180 256 181
rect 254 180 255 181
rect 253 180 254 181
rect 252 180 253 181
rect 251 180 252 181
rect 250 180 251 181
rect 249 180 250 181
rect 248 180 249 181
rect 247 180 248 181
rect 246 180 247 181
rect 245 180 246 181
rect 244 180 245 181
rect 243 180 244 181
rect 242 180 243 181
rect 241 180 242 181
rect 240 180 241 181
rect 239 180 240 181
rect 238 180 239 181
rect 237 180 238 181
rect 236 180 237 181
rect 235 180 236 181
rect 234 180 235 181
rect 233 180 234 181
rect 232 180 233 181
rect 231 180 232 181
rect 230 180 231 181
rect 229 180 230 181
rect 228 180 229 181
rect 227 180 228 181
rect 226 180 227 181
rect 225 180 226 181
rect 224 180 225 181
rect 223 180 224 181
rect 222 180 223 181
rect 221 180 222 181
rect 220 180 221 181
rect 219 180 220 181
rect 199 180 200 181
rect 198 180 199 181
rect 197 180 198 181
rect 196 180 197 181
rect 195 180 196 181
rect 194 180 195 181
rect 193 180 194 181
rect 192 180 193 181
rect 191 180 192 181
rect 190 180 191 181
rect 189 180 190 181
rect 188 180 189 181
rect 187 180 188 181
rect 186 180 187 181
rect 185 180 186 181
rect 184 180 185 181
rect 183 180 184 181
rect 182 180 183 181
rect 181 180 182 181
rect 180 180 181 181
rect 179 180 180 181
rect 178 180 179 181
rect 177 180 178 181
rect 176 180 177 181
rect 175 180 176 181
rect 174 180 175 181
rect 173 180 174 181
rect 172 180 173 181
rect 171 180 172 181
rect 170 180 171 181
rect 169 180 170 181
rect 168 180 169 181
rect 167 180 168 181
rect 166 180 167 181
rect 165 180 166 181
rect 164 180 165 181
rect 163 180 164 181
rect 162 180 163 181
rect 161 180 162 181
rect 160 180 161 181
rect 159 180 160 181
rect 158 180 159 181
rect 157 180 158 181
rect 156 180 157 181
rect 155 180 156 181
rect 154 180 155 181
rect 153 180 154 181
rect 152 180 153 181
rect 151 180 152 181
rect 150 180 151 181
rect 149 180 150 181
rect 148 180 149 181
rect 147 180 148 181
rect 146 180 147 181
rect 145 180 146 181
rect 144 180 145 181
rect 143 180 144 181
rect 142 180 143 181
rect 141 180 142 181
rect 140 180 141 181
rect 139 180 140 181
rect 138 180 139 181
rect 137 180 138 181
rect 136 180 137 181
rect 135 180 136 181
rect 134 180 135 181
rect 133 180 134 181
rect 132 180 133 181
rect 131 180 132 181
rect 130 180 131 181
rect 129 180 130 181
rect 128 180 129 181
rect 127 180 128 181
rect 126 180 127 181
rect 125 180 126 181
rect 124 180 125 181
rect 123 180 124 181
rect 122 180 123 181
rect 121 180 122 181
rect 120 180 121 181
rect 119 180 120 181
rect 118 180 119 181
rect 117 180 118 181
rect 116 180 117 181
rect 115 180 116 181
rect 114 180 115 181
rect 113 180 114 181
rect 112 180 113 181
rect 111 180 112 181
rect 110 180 111 181
rect 109 180 110 181
rect 108 180 109 181
rect 107 180 108 181
rect 106 180 107 181
rect 105 180 106 181
rect 73 180 74 181
rect 72 180 73 181
rect 71 180 72 181
rect 70 180 71 181
rect 69 180 70 181
rect 68 180 69 181
rect 67 180 68 181
rect 22 180 23 181
rect 21 180 22 181
rect 20 180 21 181
rect 19 180 20 181
rect 18 180 19 181
rect 17 180 18 181
rect 16 180 17 181
rect 15 180 16 181
rect 14 180 15 181
rect 13 180 14 181
rect 12 180 13 181
rect 11 180 12 181
rect 10 180 11 181
rect 426 181 427 182
rect 425 181 426 182
rect 424 181 425 182
rect 423 181 424 182
rect 422 181 423 182
rect 421 181 422 182
rect 420 181 421 182
rect 419 181 420 182
rect 418 181 419 182
rect 417 181 418 182
rect 416 181 417 182
rect 415 181 416 182
rect 414 181 415 182
rect 413 181 414 182
rect 412 181 413 182
rect 325 181 326 182
rect 324 181 325 182
rect 323 181 324 182
rect 322 181 323 182
rect 321 181 322 182
rect 320 181 321 182
rect 319 181 320 182
rect 318 181 319 182
rect 317 181 318 182
rect 316 181 317 182
rect 315 181 316 182
rect 314 181 315 182
rect 313 181 314 182
rect 312 181 313 182
rect 311 181 312 182
rect 310 181 311 182
rect 309 181 310 182
rect 308 181 309 182
rect 307 181 308 182
rect 306 181 307 182
rect 305 181 306 182
rect 304 181 305 182
rect 303 181 304 182
rect 302 181 303 182
rect 301 181 302 182
rect 300 181 301 182
rect 299 181 300 182
rect 298 181 299 182
rect 297 181 298 182
rect 296 181 297 182
rect 295 181 296 182
rect 294 181 295 182
rect 293 181 294 182
rect 292 181 293 182
rect 291 181 292 182
rect 290 181 291 182
rect 289 181 290 182
rect 288 181 289 182
rect 287 181 288 182
rect 259 181 260 182
rect 258 181 259 182
rect 257 181 258 182
rect 256 181 257 182
rect 255 181 256 182
rect 254 181 255 182
rect 253 181 254 182
rect 252 181 253 182
rect 251 181 252 182
rect 250 181 251 182
rect 249 181 250 182
rect 248 181 249 182
rect 247 181 248 182
rect 246 181 247 182
rect 245 181 246 182
rect 244 181 245 182
rect 243 181 244 182
rect 242 181 243 182
rect 241 181 242 182
rect 240 181 241 182
rect 239 181 240 182
rect 238 181 239 182
rect 237 181 238 182
rect 236 181 237 182
rect 235 181 236 182
rect 234 181 235 182
rect 233 181 234 182
rect 232 181 233 182
rect 231 181 232 182
rect 230 181 231 182
rect 229 181 230 182
rect 228 181 229 182
rect 227 181 228 182
rect 226 181 227 182
rect 225 181 226 182
rect 224 181 225 182
rect 223 181 224 182
rect 222 181 223 182
rect 221 181 222 182
rect 220 181 221 182
rect 219 181 220 182
rect 198 181 199 182
rect 197 181 198 182
rect 196 181 197 182
rect 195 181 196 182
rect 194 181 195 182
rect 193 181 194 182
rect 192 181 193 182
rect 191 181 192 182
rect 190 181 191 182
rect 189 181 190 182
rect 188 181 189 182
rect 187 181 188 182
rect 186 181 187 182
rect 185 181 186 182
rect 184 181 185 182
rect 183 181 184 182
rect 182 181 183 182
rect 181 181 182 182
rect 180 181 181 182
rect 179 181 180 182
rect 178 181 179 182
rect 177 181 178 182
rect 176 181 177 182
rect 175 181 176 182
rect 174 181 175 182
rect 173 181 174 182
rect 172 181 173 182
rect 171 181 172 182
rect 170 181 171 182
rect 169 181 170 182
rect 168 181 169 182
rect 167 181 168 182
rect 166 181 167 182
rect 165 181 166 182
rect 164 181 165 182
rect 163 181 164 182
rect 162 181 163 182
rect 161 181 162 182
rect 160 181 161 182
rect 159 181 160 182
rect 158 181 159 182
rect 157 181 158 182
rect 156 181 157 182
rect 155 181 156 182
rect 154 181 155 182
rect 153 181 154 182
rect 152 181 153 182
rect 151 181 152 182
rect 150 181 151 182
rect 149 181 150 182
rect 148 181 149 182
rect 147 181 148 182
rect 146 181 147 182
rect 145 181 146 182
rect 144 181 145 182
rect 143 181 144 182
rect 142 181 143 182
rect 141 181 142 182
rect 140 181 141 182
rect 139 181 140 182
rect 138 181 139 182
rect 137 181 138 182
rect 136 181 137 182
rect 135 181 136 182
rect 134 181 135 182
rect 133 181 134 182
rect 132 181 133 182
rect 131 181 132 182
rect 130 181 131 182
rect 129 181 130 182
rect 128 181 129 182
rect 127 181 128 182
rect 126 181 127 182
rect 125 181 126 182
rect 124 181 125 182
rect 123 181 124 182
rect 122 181 123 182
rect 121 181 122 182
rect 120 181 121 182
rect 119 181 120 182
rect 118 181 119 182
rect 117 181 118 182
rect 116 181 117 182
rect 115 181 116 182
rect 114 181 115 182
rect 113 181 114 182
rect 112 181 113 182
rect 111 181 112 182
rect 110 181 111 182
rect 109 181 110 182
rect 108 181 109 182
rect 107 181 108 182
rect 106 181 107 182
rect 105 181 106 182
rect 104 181 105 182
rect 103 181 104 182
rect 102 181 103 182
rect 75 181 76 182
rect 74 181 75 182
rect 73 181 74 182
rect 72 181 73 182
rect 71 181 72 182
rect 70 181 71 182
rect 69 181 70 182
rect 68 181 69 182
rect 22 181 23 182
rect 21 181 22 182
rect 20 181 21 182
rect 19 181 20 182
rect 18 181 19 182
rect 17 181 18 182
rect 16 181 17 182
rect 15 181 16 182
rect 14 181 15 182
rect 13 181 14 182
rect 12 181 13 182
rect 11 181 12 182
rect 10 181 11 182
rect 427 182 428 183
rect 426 182 427 183
rect 425 182 426 183
rect 424 182 425 183
rect 423 182 424 183
rect 422 182 423 183
rect 421 182 422 183
rect 420 182 421 183
rect 419 182 420 183
rect 418 182 419 183
rect 417 182 418 183
rect 416 182 417 183
rect 415 182 416 183
rect 414 182 415 183
rect 413 182 414 183
rect 327 182 328 183
rect 326 182 327 183
rect 325 182 326 183
rect 324 182 325 183
rect 323 182 324 183
rect 322 182 323 183
rect 321 182 322 183
rect 320 182 321 183
rect 319 182 320 183
rect 318 182 319 183
rect 317 182 318 183
rect 316 182 317 183
rect 315 182 316 183
rect 314 182 315 183
rect 313 182 314 183
rect 312 182 313 183
rect 311 182 312 183
rect 310 182 311 183
rect 309 182 310 183
rect 308 182 309 183
rect 307 182 308 183
rect 306 182 307 183
rect 305 182 306 183
rect 304 182 305 183
rect 303 182 304 183
rect 302 182 303 183
rect 301 182 302 183
rect 300 182 301 183
rect 299 182 300 183
rect 298 182 299 183
rect 297 182 298 183
rect 296 182 297 183
rect 295 182 296 183
rect 294 182 295 183
rect 293 182 294 183
rect 292 182 293 183
rect 291 182 292 183
rect 290 182 291 183
rect 289 182 290 183
rect 288 182 289 183
rect 287 182 288 183
rect 286 182 287 183
rect 285 182 286 183
rect 258 182 259 183
rect 257 182 258 183
rect 256 182 257 183
rect 255 182 256 183
rect 254 182 255 183
rect 253 182 254 183
rect 252 182 253 183
rect 251 182 252 183
rect 250 182 251 183
rect 249 182 250 183
rect 248 182 249 183
rect 247 182 248 183
rect 246 182 247 183
rect 245 182 246 183
rect 244 182 245 183
rect 243 182 244 183
rect 242 182 243 183
rect 241 182 242 183
rect 240 182 241 183
rect 239 182 240 183
rect 238 182 239 183
rect 237 182 238 183
rect 236 182 237 183
rect 235 182 236 183
rect 234 182 235 183
rect 233 182 234 183
rect 232 182 233 183
rect 231 182 232 183
rect 230 182 231 183
rect 229 182 230 183
rect 228 182 229 183
rect 227 182 228 183
rect 226 182 227 183
rect 225 182 226 183
rect 224 182 225 183
rect 223 182 224 183
rect 222 182 223 183
rect 221 182 222 183
rect 220 182 221 183
rect 219 182 220 183
rect 218 182 219 183
rect 197 182 198 183
rect 196 182 197 183
rect 195 182 196 183
rect 194 182 195 183
rect 193 182 194 183
rect 192 182 193 183
rect 191 182 192 183
rect 190 182 191 183
rect 189 182 190 183
rect 188 182 189 183
rect 187 182 188 183
rect 186 182 187 183
rect 185 182 186 183
rect 184 182 185 183
rect 183 182 184 183
rect 182 182 183 183
rect 181 182 182 183
rect 180 182 181 183
rect 179 182 180 183
rect 178 182 179 183
rect 177 182 178 183
rect 176 182 177 183
rect 175 182 176 183
rect 174 182 175 183
rect 173 182 174 183
rect 172 182 173 183
rect 171 182 172 183
rect 170 182 171 183
rect 169 182 170 183
rect 168 182 169 183
rect 167 182 168 183
rect 166 182 167 183
rect 165 182 166 183
rect 164 182 165 183
rect 163 182 164 183
rect 162 182 163 183
rect 161 182 162 183
rect 160 182 161 183
rect 159 182 160 183
rect 158 182 159 183
rect 157 182 158 183
rect 156 182 157 183
rect 155 182 156 183
rect 154 182 155 183
rect 153 182 154 183
rect 152 182 153 183
rect 151 182 152 183
rect 150 182 151 183
rect 149 182 150 183
rect 148 182 149 183
rect 147 182 148 183
rect 146 182 147 183
rect 145 182 146 183
rect 144 182 145 183
rect 143 182 144 183
rect 142 182 143 183
rect 141 182 142 183
rect 140 182 141 183
rect 139 182 140 183
rect 138 182 139 183
rect 137 182 138 183
rect 136 182 137 183
rect 135 182 136 183
rect 134 182 135 183
rect 133 182 134 183
rect 132 182 133 183
rect 131 182 132 183
rect 130 182 131 183
rect 129 182 130 183
rect 128 182 129 183
rect 127 182 128 183
rect 126 182 127 183
rect 125 182 126 183
rect 124 182 125 183
rect 123 182 124 183
rect 122 182 123 183
rect 121 182 122 183
rect 120 182 121 183
rect 119 182 120 183
rect 118 182 119 183
rect 117 182 118 183
rect 116 182 117 183
rect 115 182 116 183
rect 114 182 115 183
rect 113 182 114 183
rect 112 182 113 183
rect 111 182 112 183
rect 110 182 111 183
rect 109 182 110 183
rect 108 182 109 183
rect 107 182 108 183
rect 106 182 107 183
rect 105 182 106 183
rect 104 182 105 183
rect 103 182 104 183
rect 102 182 103 183
rect 101 182 102 183
rect 100 182 101 183
rect 99 182 100 183
rect 98 182 99 183
rect 97 182 98 183
rect 79 182 80 183
rect 78 182 79 183
rect 77 182 78 183
rect 76 182 77 183
rect 75 182 76 183
rect 74 182 75 183
rect 73 182 74 183
rect 72 182 73 183
rect 71 182 72 183
rect 70 182 71 183
rect 69 182 70 183
rect 68 182 69 183
rect 22 182 23 183
rect 21 182 22 183
rect 20 182 21 183
rect 19 182 20 183
rect 18 182 19 183
rect 17 182 18 183
rect 16 182 17 183
rect 15 182 16 183
rect 14 182 15 183
rect 13 182 14 183
rect 12 182 13 183
rect 11 182 12 183
rect 10 182 11 183
rect 428 183 429 184
rect 427 183 428 184
rect 426 183 427 184
rect 425 183 426 184
rect 424 183 425 184
rect 423 183 424 184
rect 422 183 423 184
rect 421 183 422 184
rect 420 183 421 184
rect 419 183 420 184
rect 418 183 419 184
rect 417 183 418 184
rect 416 183 417 184
rect 415 183 416 184
rect 414 183 415 184
rect 329 183 330 184
rect 328 183 329 184
rect 327 183 328 184
rect 326 183 327 184
rect 325 183 326 184
rect 324 183 325 184
rect 323 183 324 184
rect 322 183 323 184
rect 321 183 322 184
rect 320 183 321 184
rect 319 183 320 184
rect 318 183 319 184
rect 317 183 318 184
rect 316 183 317 184
rect 315 183 316 184
rect 314 183 315 184
rect 313 183 314 184
rect 312 183 313 184
rect 311 183 312 184
rect 310 183 311 184
rect 309 183 310 184
rect 308 183 309 184
rect 307 183 308 184
rect 306 183 307 184
rect 305 183 306 184
rect 304 183 305 184
rect 303 183 304 184
rect 302 183 303 184
rect 301 183 302 184
rect 300 183 301 184
rect 299 183 300 184
rect 298 183 299 184
rect 297 183 298 184
rect 296 183 297 184
rect 295 183 296 184
rect 294 183 295 184
rect 293 183 294 184
rect 292 183 293 184
rect 291 183 292 184
rect 290 183 291 184
rect 289 183 290 184
rect 288 183 289 184
rect 287 183 288 184
rect 286 183 287 184
rect 285 183 286 184
rect 284 183 285 184
rect 283 183 284 184
rect 282 183 283 184
rect 257 183 258 184
rect 256 183 257 184
rect 255 183 256 184
rect 254 183 255 184
rect 253 183 254 184
rect 252 183 253 184
rect 251 183 252 184
rect 250 183 251 184
rect 249 183 250 184
rect 248 183 249 184
rect 247 183 248 184
rect 246 183 247 184
rect 245 183 246 184
rect 244 183 245 184
rect 243 183 244 184
rect 242 183 243 184
rect 241 183 242 184
rect 240 183 241 184
rect 239 183 240 184
rect 238 183 239 184
rect 237 183 238 184
rect 236 183 237 184
rect 235 183 236 184
rect 234 183 235 184
rect 233 183 234 184
rect 232 183 233 184
rect 231 183 232 184
rect 230 183 231 184
rect 229 183 230 184
rect 228 183 229 184
rect 227 183 228 184
rect 226 183 227 184
rect 225 183 226 184
rect 224 183 225 184
rect 223 183 224 184
rect 222 183 223 184
rect 221 183 222 184
rect 220 183 221 184
rect 219 183 220 184
rect 218 183 219 184
rect 217 183 218 184
rect 196 183 197 184
rect 195 183 196 184
rect 194 183 195 184
rect 193 183 194 184
rect 192 183 193 184
rect 191 183 192 184
rect 190 183 191 184
rect 189 183 190 184
rect 188 183 189 184
rect 187 183 188 184
rect 186 183 187 184
rect 185 183 186 184
rect 184 183 185 184
rect 183 183 184 184
rect 182 183 183 184
rect 181 183 182 184
rect 180 183 181 184
rect 179 183 180 184
rect 178 183 179 184
rect 177 183 178 184
rect 176 183 177 184
rect 175 183 176 184
rect 174 183 175 184
rect 173 183 174 184
rect 172 183 173 184
rect 171 183 172 184
rect 170 183 171 184
rect 169 183 170 184
rect 168 183 169 184
rect 167 183 168 184
rect 166 183 167 184
rect 165 183 166 184
rect 164 183 165 184
rect 163 183 164 184
rect 162 183 163 184
rect 161 183 162 184
rect 160 183 161 184
rect 159 183 160 184
rect 158 183 159 184
rect 157 183 158 184
rect 156 183 157 184
rect 155 183 156 184
rect 154 183 155 184
rect 153 183 154 184
rect 152 183 153 184
rect 151 183 152 184
rect 150 183 151 184
rect 149 183 150 184
rect 148 183 149 184
rect 147 183 148 184
rect 146 183 147 184
rect 145 183 146 184
rect 144 183 145 184
rect 143 183 144 184
rect 142 183 143 184
rect 141 183 142 184
rect 140 183 141 184
rect 139 183 140 184
rect 138 183 139 184
rect 137 183 138 184
rect 136 183 137 184
rect 135 183 136 184
rect 134 183 135 184
rect 133 183 134 184
rect 132 183 133 184
rect 131 183 132 184
rect 130 183 131 184
rect 129 183 130 184
rect 128 183 129 184
rect 127 183 128 184
rect 126 183 127 184
rect 125 183 126 184
rect 124 183 125 184
rect 123 183 124 184
rect 122 183 123 184
rect 121 183 122 184
rect 120 183 121 184
rect 119 183 120 184
rect 118 183 119 184
rect 117 183 118 184
rect 116 183 117 184
rect 115 183 116 184
rect 114 183 115 184
rect 113 183 114 184
rect 112 183 113 184
rect 111 183 112 184
rect 110 183 111 184
rect 109 183 110 184
rect 108 183 109 184
rect 107 183 108 184
rect 106 183 107 184
rect 105 183 106 184
rect 104 183 105 184
rect 103 183 104 184
rect 102 183 103 184
rect 101 183 102 184
rect 100 183 101 184
rect 99 183 100 184
rect 98 183 99 184
rect 97 183 98 184
rect 96 183 97 184
rect 95 183 96 184
rect 94 183 95 184
rect 93 183 94 184
rect 92 183 93 184
rect 91 183 92 184
rect 90 183 91 184
rect 89 183 90 184
rect 88 183 89 184
rect 87 183 88 184
rect 86 183 87 184
rect 85 183 86 184
rect 84 183 85 184
rect 83 183 84 184
rect 82 183 83 184
rect 81 183 82 184
rect 80 183 81 184
rect 79 183 80 184
rect 78 183 79 184
rect 77 183 78 184
rect 76 183 77 184
rect 75 183 76 184
rect 74 183 75 184
rect 73 183 74 184
rect 72 183 73 184
rect 71 183 72 184
rect 70 183 71 184
rect 69 183 70 184
rect 68 183 69 184
rect 22 183 23 184
rect 21 183 22 184
rect 20 183 21 184
rect 19 183 20 184
rect 18 183 19 184
rect 17 183 18 184
rect 16 183 17 184
rect 15 183 16 184
rect 14 183 15 184
rect 13 183 14 184
rect 12 183 13 184
rect 11 183 12 184
rect 10 183 11 184
rect 429 184 430 185
rect 428 184 429 185
rect 427 184 428 185
rect 426 184 427 185
rect 425 184 426 185
rect 424 184 425 185
rect 423 184 424 185
rect 422 184 423 185
rect 421 184 422 185
rect 420 184 421 185
rect 419 184 420 185
rect 418 184 419 185
rect 417 184 418 185
rect 416 184 417 185
rect 415 184 416 185
rect 394 184 395 185
rect 393 184 394 185
rect 331 184 332 185
rect 330 184 331 185
rect 329 184 330 185
rect 328 184 329 185
rect 327 184 328 185
rect 326 184 327 185
rect 325 184 326 185
rect 324 184 325 185
rect 323 184 324 185
rect 322 184 323 185
rect 321 184 322 185
rect 320 184 321 185
rect 319 184 320 185
rect 318 184 319 185
rect 317 184 318 185
rect 316 184 317 185
rect 315 184 316 185
rect 314 184 315 185
rect 313 184 314 185
rect 312 184 313 185
rect 311 184 312 185
rect 310 184 311 185
rect 309 184 310 185
rect 308 184 309 185
rect 307 184 308 185
rect 306 184 307 185
rect 305 184 306 185
rect 304 184 305 185
rect 303 184 304 185
rect 302 184 303 185
rect 301 184 302 185
rect 300 184 301 185
rect 299 184 300 185
rect 298 184 299 185
rect 297 184 298 185
rect 296 184 297 185
rect 295 184 296 185
rect 294 184 295 185
rect 293 184 294 185
rect 292 184 293 185
rect 291 184 292 185
rect 290 184 291 185
rect 289 184 290 185
rect 288 184 289 185
rect 287 184 288 185
rect 286 184 287 185
rect 285 184 286 185
rect 284 184 285 185
rect 283 184 284 185
rect 282 184 283 185
rect 281 184 282 185
rect 280 184 281 185
rect 257 184 258 185
rect 256 184 257 185
rect 255 184 256 185
rect 254 184 255 185
rect 253 184 254 185
rect 252 184 253 185
rect 251 184 252 185
rect 250 184 251 185
rect 249 184 250 185
rect 248 184 249 185
rect 247 184 248 185
rect 246 184 247 185
rect 245 184 246 185
rect 244 184 245 185
rect 243 184 244 185
rect 242 184 243 185
rect 241 184 242 185
rect 240 184 241 185
rect 239 184 240 185
rect 238 184 239 185
rect 237 184 238 185
rect 236 184 237 185
rect 235 184 236 185
rect 234 184 235 185
rect 233 184 234 185
rect 232 184 233 185
rect 231 184 232 185
rect 230 184 231 185
rect 229 184 230 185
rect 228 184 229 185
rect 227 184 228 185
rect 226 184 227 185
rect 225 184 226 185
rect 224 184 225 185
rect 223 184 224 185
rect 222 184 223 185
rect 221 184 222 185
rect 220 184 221 185
rect 219 184 220 185
rect 218 184 219 185
rect 217 184 218 185
rect 195 184 196 185
rect 194 184 195 185
rect 193 184 194 185
rect 192 184 193 185
rect 191 184 192 185
rect 190 184 191 185
rect 189 184 190 185
rect 188 184 189 185
rect 187 184 188 185
rect 186 184 187 185
rect 185 184 186 185
rect 184 184 185 185
rect 183 184 184 185
rect 182 184 183 185
rect 181 184 182 185
rect 180 184 181 185
rect 179 184 180 185
rect 178 184 179 185
rect 177 184 178 185
rect 176 184 177 185
rect 175 184 176 185
rect 174 184 175 185
rect 173 184 174 185
rect 172 184 173 185
rect 171 184 172 185
rect 170 184 171 185
rect 169 184 170 185
rect 168 184 169 185
rect 167 184 168 185
rect 166 184 167 185
rect 165 184 166 185
rect 164 184 165 185
rect 163 184 164 185
rect 162 184 163 185
rect 161 184 162 185
rect 160 184 161 185
rect 159 184 160 185
rect 158 184 159 185
rect 157 184 158 185
rect 156 184 157 185
rect 155 184 156 185
rect 154 184 155 185
rect 153 184 154 185
rect 152 184 153 185
rect 151 184 152 185
rect 150 184 151 185
rect 149 184 150 185
rect 148 184 149 185
rect 147 184 148 185
rect 146 184 147 185
rect 145 184 146 185
rect 144 184 145 185
rect 143 184 144 185
rect 142 184 143 185
rect 141 184 142 185
rect 140 184 141 185
rect 139 184 140 185
rect 138 184 139 185
rect 137 184 138 185
rect 136 184 137 185
rect 135 184 136 185
rect 134 184 135 185
rect 133 184 134 185
rect 132 184 133 185
rect 131 184 132 185
rect 130 184 131 185
rect 129 184 130 185
rect 128 184 129 185
rect 127 184 128 185
rect 126 184 127 185
rect 125 184 126 185
rect 124 184 125 185
rect 123 184 124 185
rect 122 184 123 185
rect 121 184 122 185
rect 120 184 121 185
rect 119 184 120 185
rect 118 184 119 185
rect 117 184 118 185
rect 116 184 117 185
rect 115 184 116 185
rect 114 184 115 185
rect 113 184 114 185
rect 112 184 113 185
rect 111 184 112 185
rect 110 184 111 185
rect 109 184 110 185
rect 108 184 109 185
rect 107 184 108 185
rect 106 184 107 185
rect 105 184 106 185
rect 104 184 105 185
rect 103 184 104 185
rect 102 184 103 185
rect 101 184 102 185
rect 100 184 101 185
rect 99 184 100 185
rect 98 184 99 185
rect 97 184 98 185
rect 96 184 97 185
rect 95 184 96 185
rect 94 184 95 185
rect 93 184 94 185
rect 92 184 93 185
rect 91 184 92 185
rect 90 184 91 185
rect 89 184 90 185
rect 88 184 89 185
rect 87 184 88 185
rect 86 184 87 185
rect 85 184 86 185
rect 84 184 85 185
rect 83 184 84 185
rect 82 184 83 185
rect 81 184 82 185
rect 80 184 81 185
rect 79 184 80 185
rect 78 184 79 185
rect 77 184 78 185
rect 76 184 77 185
rect 75 184 76 185
rect 74 184 75 185
rect 73 184 74 185
rect 72 184 73 185
rect 71 184 72 185
rect 70 184 71 185
rect 69 184 70 185
rect 68 184 69 185
rect 23 184 24 185
rect 22 184 23 185
rect 21 184 22 185
rect 20 184 21 185
rect 19 184 20 185
rect 18 184 19 185
rect 17 184 18 185
rect 16 184 17 185
rect 15 184 16 185
rect 14 184 15 185
rect 13 184 14 185
rect 12 184 13 185
rect 11 184 12 185
rect 10 184 11 185
rect 430 185 431 186
rect 429 185 430 186
rect 428 185 429 186
rect 427 185 428 186
rect 426 185 427 186
rect 425 185 426 186
rect 424 185 425 186
rect 423 185 424 186
rect 422 185 423 186
rect 421 185 422 186
rect 420 185 421 186
rect 419 185 420 186
rect 418 185 419 186
rect 417 185 418 186
rect 416 185 417 186
rect 395 185 396 186
rect 394 185 395 186
rect 393 185 394 186
rect 333 185 334 186
rect 332 185 333 186
rect 331 185 332 186
rect 330 185 331 186
rect 329 185 330 186
rect 328 185 329 186
rect 327 185 328 186
rect 326 185 327 186
rect 325 185 326 186
rect 324 185 325 186
rect 323 185 324 186
rect 322 185 323 186
rect 321 185 322 186
rect 320 185 321 186
rect 319 185 320 186
rect 318 185 319 186
rect 317 185 318 186
rect 316 185 317 186
rect 315 185 316 186
rect 314 185 315 186
rect 313 185 314 186
rect 312 185 313 186
rect 311 185 312 186
rect 310 185 311 186
rect 309 185 310 186
rect 308 185 309 186
rect 307 185 308 186
rect 306 185 307 186
rect 305 185 306 186
rect 304 185 305 186
rect 303 185 304 186
rect 302 185 303 186
rect 301 185 302 186
rect 300 185 301 186
rect 299 185 300 186
rect 298 185 299 186
rect 297 185 298 186
rect 296 185 297 186
rect 295 185 296 186
rect 294 185 295 186
rect 293 185 294 186
rect 292 185 293 186
rect 291 185 292 186
rect 290 185 291 186
rect 289 185 290 186
rect 288 185 289 186
rect 287 185 288 186
rect 286 185 287 186
rect 285 185 286 186
rect 284 185 285 186
rect 283 185 284 186
rect 282 185 283 186
rect 281 185 282 186
rect 280 185 281 186
rect 279 185 280 186
rect 278 185 279 186
rect 256 185 257 186
rect 255 185 256 186
rect 254 185 255 186
rect 253 185 254 186
rect 252 185 253 186
rect 251 185 252 186
rect 250 185 251 186
rect 249 185 250 186
rect 248 185 249 186
rect 247 185 248 186
rect 246 185 247 186
rect 245 185 246 186
rect 244 185 245 186
rect 243 185 244 186
rect 242 185 243 186
rect 241 185 242 186
rect 240 185 241 186
rect 239 185 240 186
rect 238 185 239 186
rect 237 185 238 186
rect 236 185 237 186
rect 235 185 236 186
rect 234 185 235 186
rect 233 185 234 186
rect 232 185 233 186
rect 231 185 232 186
rect 230 185 231 186
rect 229 185 230 186
rect 228 185 229 186
rect 227 185 228 186
rect 226 185 227 186
rect 225 185 226 186
rect 224 185 225 186
rect 223 185 224 186
rect 222 185 223 186
rect 221 185 222 186
rect 220 185 221 186
rect 219 185 220 186
rect 218 185 219 186
rect 217 185 218 186
rect 216 185 217 186
rect 194 185 195 186
rect 193 185 194 186
rect 192 185 193 186
rect 191 185 192 186
rect 190 185 191 186
rect 189 185 190 186
rect 188 185 189 186
rect 187 185 188 186
rect 186 185 187 186
rect 185 185 186 186
rect 184 185 185 186
rect 183 185 184 186
rect 182 185 183 186
rect 181 185 182 186
rect 180 185 181 186
rect 179 185 180 186
rect 178 185 179 186
rect 177 185 178 186
rect 176 185 177 186
rect 175 185 176 186
rect 174 185 175 186
rect 173 185 174 186
rect 172 185 173 186
rect 171 185 172 186
rect 170 185 171 186
rect 169 185 170 186
rect 168 185 169 186
rect 167 185 168 186
rect 166 185 167 186
rect 165 185 166 186
rect 164 185 165 186
rect 163 185 164 186
rect 162 185 163 186
rect 161 185 162 186
rect 160 185 161 186
rect 159 185 160 186
rect 158 185 159 186
rect 157 185 158 186
rect 156 185 157 186
rect 155 185 156 186
rect 154 185 155 186
rect 153 185 154 186
rect 152 185 153 186
rect 151 185 152 186
rect 150 185 151 186
rect 149 185 150 186
rect 148 185 149 186
rect 147 185 148 186
rect 146 185 147 186
rect 145 185 146 186
rect 144 185 145 186
rect 143 185 144 186
rect 142 185 143 186
rect 141 185 142 186
rect 140 185 141 186
rect 139 185 140 186
rect 138 185 139 186
rect 137 185 138 186
rect 136 185 137 186
rect 135 185 136 186
rect 134 185 135 186
rect 133 185 134 186
rect 132 185 133 186
rect 131 185 132 186
rect 130 185 131 186
rect 129 185 130 186
rect 128 185 129 186
rect 127 185 128 186
rect 126 185 127 186
rect 125 185 126 186
rect 124 185 125 186
rect 123 185 124 186
rect 122 185 123 186
rect 121 185 122 186
rect 120 185 121 186
rect 119 185 120 186
rect 118 185 119 186
rect 117 185 118 186
rect 116 185 117 186
rect 115 185 116 186
rect 114 185 115 186
rect 113 185 114 186
rect 112 185 113 186
rect 111 185 112 186
rect 110 185 111 186
rect 109 185 110 186
rect 108 185 109 186
rect 107 185 108 186
rect 106 185 107 186
rect 105 185 106 186
rect 104 185 105 186
rect 103 185 104 186
rect 102 185 103 186
rect 101 185 102 186
rect 100 185 101 186
rect 99 185 100 186
rect 98 185 99 186
rect 97 185 98 186
rect 96 185 97 186
rect 95 185 96 186
rect 94 185 95 186
rect 93 185 94 186
rect 92 185 93 186
rect 91 185 92 186
rect 90 185 91 186
rect 89 185 90 186
rect 88 185 89 186
rect 87 185 88 186
rect 86 185 87 186
rect 85 185 86 186
rect 84 185 85 186
rect 83 185 84 186
rect 82 185 83 186
rect 81 185 82 186
rect 80 185 81 186
rect 79 185 80 186
rect 78 185 79 186
rect 77 185 78 186
rect 76 185 77 186
rect 75 185 76 186
rect 74 185 75 186
rect 73 185 74 186
rect 72 185 73 186
rect 71 185 72 186
rect 70 185 71 186
rect 69 185 70 186
rect 68 185 69 186
rect 23 185 24 186
rect 22 185 23 186
rect 21 185 22 186
rect 20 185 21 186
rect 19 185 20 186
rect 18 185 19 186
rect 17 185 18 186
rect 16 185 17 186
rect 15 185 16 186
rect 14 185 15 186
rect 13 185 14 186
rect 12 185 13 186
rect 11 185 12 186
rect 10 185 11 186
rect 432 186 433 187
rect 431 186 432 187
rect 430 186 431 187
rect 429 186 430 187
rect 428 186 429 187
rect 427 186 428 187
rect 426 186 427 187
rect 425 186 426 187
rect 424 186 425 187
rect 423 186 424 187
rect 422 186 423 187
rect 421 186 422 187
rect 420 186 421 187
rect 419 186 420 187
rect 418 186 419 187
rect 417 186 418 187
rect 395 186 396 187
rect 394 186 395 187
rect 393 186 394 187
rect 334 186 335 187
rect 333 186 334 187
rect 332 186 333 187
rect 331 186 332 187
rect 330 186 331 187
rect 329 186 330 187
rect 328 186 329 187
rect 327 186 328 187
rect 326 186 327 187
rect 325 186 326 187
rect 324 186 325 187
rect 323 186 324 187
rect 322 186 323 187
rect 321 186 322 187
rect 320 186 321 187
rect 319 186 320 187
rect 318 186 319 187
rect 317 186 318 187
rect 316 186 317 187
rect 315 186 316 187
rect 314 186 315 187
rect 313 186 314 187
rect 312 186 313 187
rect 311 186 312 187
rect 310 186 311 187
rect 309 186 310 187
rect 308 186 309 187
rect 307 186 308 187
rect 306 186 307 187
rect 305 186 306 187
rect 304 186 305 187
rect 303 186 304 187
rect 302 186 303 187
rect 301 186 302 187
rect 300 186 301 187
rect 299 186 300 187
rect 298 186 299 187
rect 297 186 298 187
rect 296 186 297 187
rect 295 186 296 187
rect 294 186 295 187
rect 293 186 294 187
rect 292 186 293 187
rect 291 186 292 187
rect 290 186 291 187
rect 289 186 290 187
rect 288 186 289 187
rect 287 186 288 187
rect 286 186 287 187
rect 285 186 286 187
rect 284 186 285 187
rect 283 186 284 187
rect 282 186 283 187
rect 281 186 282 187
rect 280 186 281 187
rect 279 186 280 187
rect 278 186 279 187
rect 277 186 278 187
rect 276 186 277 187
rect 255 186 256 187
rect 254 186 255 187
rect 253 186 254 187
rect 252 186 253 187
rect 251 186 252 187
rect 250 186 251 187
rect 249 186 250 187
rect 248 186 249 187
rect 247 186 248 187
rect 246 186 247 187
rect 245 186 246 187
rect 244 186 245 187
rect 243 186 244 187
rect 242 186 243 187
rect 241 186 242 187
rect 240 186 241 187
rect 239 186 240 187
rect 238 186 239 187
rect 237 186 238 187
rect 236 186 237 187
rect 235 186 236 187
rect 234 186 235 187
rect 233 186 234 187
rect 232 186 233 187
rect 231 186 232 187
rect 230 186 231 187
rect 229 186 230 187
rect 228 186 229 187
rect 227 186 228 187
rect 226 186 227 187
rect 225 186 226 187
rect 224 186 225 187
rect 223 186 224 187
rect 222 186 223 187
rect 221 186 222 187
rect 220 186 221 187
rect 219 186 220 187
rect 218 186 219 187
rect 217 186 218 187
rect 216 186 217 187
rect 193 186 194 187
rect 192 186 193 187
rect 191 186 192 187
rect 190 186 191 187
rect 189 186 190 187
rect 188 186 189 187
rect 187 186 188 187
rect 186 186 187 187
rect 185 186 186 187
rect 184 186 185 187
rect 183 186 184 187
rect 182 186 183 187
rect 181 186 182 187
rect 180 186 181 187
rect 179 186 180 187
rect 178 186 179 187
rect 177 186 178 187
rect 176 186 177 187
rect 175 186 176 187
rect 174 186 175 187
rect 173 186 174 187
rect 172 186 173 187
rect 171 186 172 187
rect 170 186 171 187
rect 169 186 170 187
rect 168 186 169 187
rect 167 186 168 187
rect 166 186 167 187
rect 165 186 166 187
rect 164 186 165 187
rect 163 186 164 187
rect 162 186 163 187
rect 161 186 162 187
rect 160 186 161 187
rect 159 186 160 187
rect 158 186 159 187
rect 157 186 158 187
rect 156 186 157 187
rect 155 186 156 187
rect 154 186 155 187
rect 153 186 154 187
rect 152 186 153 187
rect 151 186 152 187
rect 150 186 151 187
rect 149 186 150 187
rect 148 186 149 187
rect 147 186 148 187
rect 146 186 147 187
rect 145 186 146 187
rect 144 186 145 187
rect 143 186 144 187
rect 142 186 143 187
rect 141 186 142 187
rect 140 186 141 187
rect 139 186 140 187
rect 138 186 139 187
rect 137 186 138 187
rect 136 186 137 187
rect 135 186 136 187
rect 134 186 135 187
rect 133 186 134 187
rect 132 186 133 187
rect 131 186 132 187
rect 130 186 131 187
rect 129 186 130 187
rect 128 186 129 187
rect 127 186 128 187
rect 126 186 127 187
rect 125 186 126 187
rect 124 186 125 187
rect 123 186 124 187
rect 122 186 123 187
rect 121 186 122 187
rect 120 186 121 187
rect 119 186 120 187
rect 118 186 119 187
rect 117 186 118 187
rect 116 186 117 187
rect 115 186 116 187
rect 114 186 115 187
rect 113 186 114 187
rect 112 186 113 187
rect 111 186 112 187
rect 110 186 111 187
rect 109 186 110 187
rect 108 186 109 187
rect 107 186 108 187
rect 106 186 107 187
rect 105 186 106 187
rect 104 186 105 187
rect 103 186 104 187
rect 102 186 103 187
rect 101 186 102 187
rect 100 186 101 187
rect 99 186 100 187
rect 98 186 99 187
rect 97 186 98 187
rect 96 186 97 187
rect 95 186 96 187
rect 94 186 95 187
rect 93 186 94 187
rect 92 186 93 187
rect 91 186 92 187
rect 90 186 91 187
rect 89 186 90 187
rect 88 186 89 187
rect 87 186 88 187
rect 86 186 87 187
rect 85 186 86 187
rect 84 186 85 187
rect 83 186 84 187
rect 82 186 83 187
rect 81 186 82 187
rect 80 186 81 187
rect 79 186 80 187
rect 78 186 79 187
rect 77 186 78 187
rect 76 186 77 187
rect 75 186 76 187
rect 74 186 75 187
rect 73 186 74 187
rect 72 186 73 187
rect 71 186 72 187
rect 70 186 71 187
rect 69 186 70 187
rect 68 186 69 187
rect 24 186 25 187
rect 23 186 24 187
rect 22 186 23 187
rect 21 186 22 187
rect 20 186 21 187
rect 19 186 20 187
rect 18 186 19 187
rect 17 186 18 187
rect 16 186 17 187
rect 15 186 16 187
rect 14 186 15 187
rect 13 186 14 187
rect 12 186 13 187
rect 11 186 12 187
rect 10 186 11 187
rect 433 187 434 188
rect 432 187 433 188
rect 431 187 432 188
rect 430 187 431 188
rect 429 187 430 188
rect 428 187 429 188
rect 427 187 428 188
rect 426 187 427 188
rect 425 187 426 188
rect 424 187 425 188
rect 423 187 424 188
rect 422 187 423 188
rect 421 187 422 188
rect 420 187 421 188
rect 419 187 420 188
rect 395 187 396 188
rect 394 187 395 188
rect 393 187 394 188
rect 336 187 337 188
rect 335 187 336 188
rect 334 187 335 188
rect 333 187 334 188
rect 332 187 333 188
rect 331 187 332 188
rect 330 187 331 188
rect 329 187 330 188
rect 328 187 329 188
rect 327 187 328 188
rect 326 187 327 188
rect 325 187 326 188
rect 324 187 325 188
rect 323 187 324 188
rect 322 187 323 188
rect 321 187 322 188
rect 320 187 321 188
rect 319 187 320 188
rect 318 187 319 188
rect 317 187 318 188
rect 316 187 317 188
rect 315 187 316 188
rect 314 187 315 188
rect 313 187 314 188
rect 312 187 313 188
rect 311 187 312 188
rect 310 187 311 188
rect 309 187 310 188
rect 308 187 309 188
rect 307 187 308 188
rect 306 187 307 188
rect 305 187 306 188
rect 304 187 305 188
rect 303 187 304 188
rect 302 187 303 188
rect 301 187 302 188
rect 300 187 301 188
rect 299 187 300 188
rect 298 187 299 188
rect 297 187 298 188
rect 296 187 297 188
rect 295 187 296 188
rect 294 187 295 188
rect 293 187 294 188
rect 292 187 293 188
rect 291 187 292 188
rect 290 187 291 188
rect 289 187 290 188
rect 288 187 289 188
rect 287 187 288 188
rect 286 187 287 188
rect 285 187 286 188
rect 284 187 285 188
rect 283 187 284 188
rect 282 187 283 188
rect 281 187 282 188
rect 280 187 281 188
rect 279 187 280 188
rect 278 187 279 188
rect 277 187 278 188
rect 276 187 277 188
rect 275 187 276 188
rect 274 187 275 188
rect 255 187 256 188
rect 254 187 255 188
rect 253 187 254 188
rect 252 187 253 188
rect 251 187 252 188
rect 250 187 251 188
rect 249 187 250 188
rect 248 187 249 188
rect 247 187 248 188
rect 246 187 247 188
rect 245 187 246 188
rect 244 187 245 188
rect 243 187 244 188
rect 242 187 243 188
rect 241 187 242 188
rect 240 187 241 188
rect 239 187 240 188
rect 238 187 239 188
rect 237 187 238 188
rect 236 187 237 188
rect 235 187 236 188
rect 234 187 235 188
rect 233 187 234 188
rect 232 187 233 188
rect 231 187 232 188
rect 230 187 231 188
rect 229 187 230 188
rect 228 187 229 188
rect 227 187 228 188
rect 226 187 227 188
rect 225 187 226 188
rect 224 187 225 188
rect 223 187 224 188
rect 222 187 223 188
rect 221 187 222 188
rect 220 187 221 188
rect 219 187 220 188
rect 218 187 219 188
rect 217 187 218 188
rect 216 187 217 188
rect 215 187 216 188
rect 192 187 193 188
rect 191 187 192 188
rect 190 187 191 188
rect 189 187 190 188
rect 188 187 189 188
rect 187 187 188 188
rect 186 187 187 188
rect 185 187 186 188
rect 184 187 185 188
rect 183 187 184 188
rect 182 187 183 188
rect 181 187 182 188
rect 180 187 181 188
rect 179 187 180 188
rect 178 187 179 188
rect 177 187 178 188
rect 176 187 177 188
rect 175 187 176 188
rect 174 187 175 188
rect 173 187 174 188
rect 172 187 173 188
rect 171 187 172 188
rect 170 187 171 188
rect 169 187 170 188
rect 168 187 169 188
rect 167 187 168 188
rect 166 187 167 188
rect 165 187 166 188
rect 164 187 165 188
rect 163 187 164 188
rect 162 187 163 188
rect 161 187 162 188
rect 160 187 161 188
rect 159 187 160 188
rect 158 187 159 188
rect 157 187 158 188
rect 156 187 157 188
rect 155 187 156 188
rect 154 187 155 188
rect 153 187 154 188
rect 152 187 153 188
rect 151 187 152 188
rect 150 187 151 188
rect 149 187 150 188
rect 148 187 149 188
rect 147 187 148 188
rect 146 187 147 188
rect 145 187 146 188
rect 144 187 145 188
rect 143 187 144 188
rect 142 187 143 188
rect 141 187 142 188
rect 140 187 141 188
rect 139 187 140 188
rect 138 187 139 188
rect 137 187 138 188
rect 136 187 137 188
rect 135 187 136 188
rect 134 187 135 188
rect 133 187 134 188
rect 132 187 133 188
rect 131 187 132 188
rect 130 187 131 188
rect 129 187 130 188
rect 128 187 129 188
rect 127 187 128 188
rect 126 187 127 188
rect 125 187 126 188
rect 124 187 125 188
rect 123 187 124 188
rect 122 187 123 188
rect 121 187 122 188
rect 120 187 121 188
rect 119 187 120 188
rect 118 187 119 188
rect 117 187 118 188
rect 116 187 117 188
rect 115 187 116 188
rect 114 187 115 188
rect 113 187 114 188
rect 112 187 113 188
rect 111 187 112 188
rect 110 187 111 188
rect 109 187 110 188
rect 108 187 109 188
rect 107 187 108 188
rect 106 187 107 188
rect 105 187 106 188
rect 104 187 105 188
rect 103 187 104 188
rect 102 187 103 188
rect 101 187 102 188
rect 100 187 101 188
rect 99 187 100 188
rect 98 187 99 188
rect 97 187 98 188
rect 96 187 97 188
rect 95 187 96 188
rect 94 187 95 188
rect 93 187 94 188
rect 92 187 93 188
rect 91 187 92 188
rect 90 187 91 188
rect 89 187 90 188
rect 88 187 89 188
rect 87 187 88 188
rect 86 187 87 188
rect 85 187 86 188
rect 84 187 85 188
rect 83 187 84 188
rect 82 187 83 188
rect 81 187 82 188
rect 80 187 81 188
rect 79 187 80 188
rect 78 187 79 188
rect 77 187 78 188
rect 76 187 77 188
rect 75 187 76 188
rect 74 187 75 188
rect 73 187 74 188
rect 72 187 73 188
rect 71 187 72 188
rect 70 187 71 188
rect 69 187 70 188
rect 68 187 69 188
rect 24 187 25 188
rect 23 187 24 188
rect 22 187 23 188
rect 21 187 22 188
rect 20 187 21 188
rect 19 187 20 188
rect 18 187 19 188
rect 17 187 18 188
rect 16 187 17 188
rect 15 187 16 188
rect 14 187 15 188
rect 13 187 14 188
rect 12 187 13 188
rect 11 187 12 188
rect 10 187 11 188
rect 478 188 479 189
rect 434 188 435 189
rect 433 188 434 189
rect 432 188 433 189
rect 431 188 432 189
rect 430 188 431 189
rect 429 188 430 189
rect 428 188 429 189
rect 427 188 428 189
rect 426 188 427 189
rect 425 188 426 189
rect 424 188 425 189
rect 423 188 424 189
rect 422 188 423 189
rect 421 188 422 189
rect 420 188 421 189
rect 395 188 396 189
rect 394 188 395 189
rect 393 188 394 189
rect 337 188 338 189
rect 336 188 337 189
rect 335 188 336 189
rect 334 188 335 189
rect 333 188 334 189
rect 332 188 333 189
rect 331 188 332 189
rect 330 188 331 189
rect 329 188 330 189
rect 328 188 329 189
rect 327 188 328 189
rect 326 188 327 189
rect 325 188 326 189
rect 324 188 325 189
rect 323 188 324 189
rect 322 188 323 189
rect 321 188 322 189
rect 320 188 321 189
rect 319 188 320 189
rect 318 188 319 189
rect 317 188 318 189
rect 316 188 317 189
rect 315 188 316 189
rect 314 188 315 189
rect 313 188 314 189
rect 312 188 313 189
rect 311 188 312 189
rect 310 188 311 189
rect 309 188 310 189
rect 308 188 309 189
rect 307 188 308 189
rect 306 188 307 189
rect 305 188 306 189
rect 304 188 305 189
rect 303 188 304 189
rect 302 188 303 189
rect 301 188 302 189
rect 300 188 301 189
rect 299 188 300 189
rect 298 188 299 189
rect 297 188 298 189
rect 296 188 297 189
rect 295 188 296 189
rect 294 188 295 189
rect 293 188 294 189
rect 292 188 293 189
rect 291 188 292 189
rect 290 188 291 189
rect 289 188 290 189
rect 288 188 289 189
rect 287 188 288 189
rect 286 188 287 189
rect 285 188 286 189
rect 284 188 285 189
rect 283 188 284 189
rect 282 188 283 189
rect 281 188 282 189
rect 280 188 281 189
rect 279 188 280 189
rect 278 188 279 189
rect 277 188 278 189
rect 276 188 277 189
rect 275 188 276 189
rect 274 188 275 189
rect 273 188 274 189
rect 254 188 255 189
rect 253 188 254 189
rect 252 188 253 189
rect 251 188 252 189
rect 250 188 251 189
rect 249 188 250 189
rect 248 188 249 189
rect 247 188 248 189
rect 246 188 247 189
rect 245 188 246 189
rect 244 188 245 189
rect 243 188 244 189
rect 242 188 243 189
rect 241 188 242 189
rect 240 188 241 189
rect 239 188 240 189
rect 238 188 239 189
rect 237 188 238 189
rect 236 188 237 189
rect 235 188 236 189
rect 234 188 235 189
rect 233 188 234 189
rect 232 188 233 189
rect 231 188 232 189
rect 230 188 231 189
rect 229 188 230 189
rect 228 188 229 189
rect 227 188 228 189
rect 226 188 227 189
rect 225 188 226 189
rect 224 188 225 189
rect 223 188 224 189
rect 222 188 223 189
rect 221 188 222 189
rect 220 188 221 189
rect 219 188 220 189
rect 218 188 219 189
rect 217 188 218 189
rect 216 188 217 189
rect 215 188 216 189
rect 214 188 215 189
rect 191 188 192 189
rect 190 188 191 189
rect 189 188 190 189
rect 188 188 189 189
rect 187 188 188 189
rect 186 188 187 189
rect 185 188 186 189
rect 184 188 185 189
rect 183 188 184 189
rect 182 188 183 189
rect 181 188 182 189
rect 180 188 181 189
rect 179 188 180 189
rect 178 188 179 189
rect 177 188 178 189
rect 176 188 177 189
rect 175 188 176 189
rect 174 188 175 189
rect 173 188 174 189
rect 172 188 173 189
rect 171 188 172 189
rect 170 188 171 189
rect 169 188 170 189
rect 168 188 169 189
rect 167 188 168 189
rect 166 188 167 189
rect 165 188 166 189
rect 164 188 165 189
rect 163 188 164 189
rect 162 188 163 189
rect 161 188 162 189
rect 160 188 161 189
rect 159 188 160 189
rect 158 188 159 189
rect 157 188 158 189
rect 156 188 157 189
rect 155 188 156 189
rect 154 188 155 189
rect 153 188 154 189
rect 152 188 153 189
rect 151 188 152 189
rect 150 188 151 189
rect 149 188 150 189
rect 148 188 149 189
rect 147 188 148 189
rect 146 188 147 189
rect 145 188 146 189
rect 144 188 145 189
rect 143 188 144 189
rect 142 188 143 189
rect 141 188 142 189
rect 140 188 141 189
rect 139 188 140 189
rect 138 188 139 189
rect 137 188 138 189
rect 136 188 137 189
rect 135 188 136 189
rect 134 188 135 189
rect 133 188 134 189
rect 132 188 133 189
rect 131 188 132 189
rect 130 188 131 189
rect 129 188 130 189
rect 128 188 129 189
rect 127 188 128 189
rect 126 188 127 189
rect 125 188 126 189
rect 124 188 125 189
rect 123 188 124 189
rect 122 188 123 189
rect 121 188 122 189
rect 120 188 121 189
rect 119 188 120 189
rect 118 188 119 189
rect 117 188 118 189
rect 116 188 117 189
rect 115 188 116 189
rect 114 188 115 189
rect 113 188 114 189
rect 112 188 113 189
rect 111 188 112 189
rect 110 188 111 189
rect 109 188 110 189
rect 108 188 109 189
rect 107 188 108 189
rect 106 188 107 189
rect 105 188 106 189
rect 104 188 105 189
rect 103 188 104 189
rect 102 188 103 189
rect 101 188 102 189
rect 100 188 101 189
rect 99 188 100 189
rect 98 188 99 189
rect 97 188 98 189
rect 96 188 97 189
rect 95 188 96 189
rect 94 188 95 189
rect 93 188 94 189
rect 92 188 93 189
rect 91 188 92 189
rect 90 188 91 189
rect 89 188 90 189
rect 88 188 89 189
rect 87 188 88 189
rect 86 188 87 189
rect 85 188 86 189
rect 84 188 85 189
rect 83 188 84 189
rect 82 188 83 189
rect 81 188 82 189
rect 80 188 81 189
rect 79 188 80 189
rect 78 188 79 189
rect 77 188 78 189
rect 76 188 77 189
rect 75 188 76 189
rect 74 188 75 189
rect 73 188 74 189
rect 72 188 73 189
rect 71 188 72 189
rect 70 188 71 189
rect 69 188 70 189
rect 68 188 69 189
rect 67 188 68 189
rect 25 188 26 189
rect 24 188 25 189
rect 23 188 24 189
rect 22 188 23 189
rect 21 188 22 189
rect 20 188 21 189
rect 19 188 20 189
rect 18 188 19 189
rect 17 188 18 189
rect 16 188 17 189
rect 15 188 16 189
rect 14 188 15 189
rect 13 188 14 189
rect 12 188 13 189
rect 11 188 12 189
rect 10 188 11 189
rect 478 189 479 190
rect 458 189 459 190
rect 435 189 436 190
rect 434 189 435 190
rect 433 189 434 190
rect 432 189 433 190
rect 431 189 432 190
rect 430 189 431 190
rect 429 189 430 190
rect 428 189 429 190
rect 427 189 428 190
rect 426 189 427 190
rect 425 189 426 190
rect 424 189 425 190
rect 423 189 424 190
rect 422 189 423 190
rect 421 189 422 190
rect 396 189 397 190
rect 395 189 396 190
rect 394 189 395 190
rect 393 189 394 190
rect 338 189 339 190
rect 337 189 338 190
rect 336 189 337 190
rect 335 189 336 190
rect 334 189 335 190
rect 333 189 334 190
rect 332 189 333 190
rect 331 189 332 190
rect 330 189 331 190
rect 329 189 330 190
rect 328 189 329 190
rect 327 189 328 190
rect 326 189 327 190
rect 325 189 326 190
rect 324 189 325 190
rect 323 189 324 190
rect 322 189 323 190
rect 321 189 322 190
rect 320 189 321 190
rect 319 189 320 190
rect 318 189 319 190
rect 317 189 318 190
rect 316 189 317 190
rect 315 189 316 190
rect 314 189 315 190
rect 313 189 314 190
rect 312 189 313 190
rect 311 189 312 190
rect 310 189 311 190
rect 309 189 310 190
rect 308 189 309 190
rect 307 189 308 190
rect 306 189 307 190
rect 305 189 306 190
rect 304 189 305 190
rect 303 189 304 190
rect 302 189 303 190
rect 301 189 302 190
rect 300 189 301 190
rect 299 189 300 190
rect 298 189 299 190
rect 297 189 298 190
rect 296 189 297 190
rect 295 189 296 190
rect 294 189 295 190
rect 293 189 294 190
rect 292 189 293 190
rect 291 189 292 190
rect 290 189 291 190
rect 289 189 290 190
rect 288 189 289 190
rect 287 189 288 190
rect 286 189 287 190
rect 285 189 286 190
rect 284 189 285 190
rect 283 189 284 190
rect 282 189 283 190
rect 281 189 282 190
rect 280 189 281 190
rect 279 189 280 190
rect 278 189 279 190
rect 277 189 278 190
rect 276 189 277 190
rect 275 189 276 190
rect 274 189 275 190
rect 273 189 274 190
rect 272 189 273 190
rect 271 189 272 190
rect 253 189 254 190
rect 252 189 253 190
rect 251 189 252 190
rect 250 189 251 190
rect 249 189 250 190
rect 248 189 249 190
rect 247 189 248 190
rect 246 189 247 190
rect 245 189 246 190
rect 244 189 245 190
rect 243 189 244 190
rect 242 189 243 190
rect 241 189 242 190
rect 240 189 241 190
rect 239 189 240 190
rect 238 189 239 190
rect 237 189 238 190
rect 236 189 237 190
rect 235 189 236 190
rect 234 189 235 190
rect 233 189 234 190
rect 232 189 233 190
rect 231 189 232 190
rect 230 189 231 190
rect 229 189 230 190
rect 228 189 229 190
rect 227 189 228 190
rect 226 189 227 190
rect 225 189 226 190
rect 224 189 225 190
rect 223 189 224 190
rect 222 189 223 190
rect 221 189 222 190
rect 220 189 221 190
rect 219 189 220 190
rect 218 189 219 190
rect 217 189 218 190
rect 216 189 217 190
rect 215 189 216 190
rect 214 189 215 190
rect 190 189 191 190
rect 189 189 190 190
rect 188 189 189 190
rect 187 189 188 190
rect 186 189 187 190
rect 185 189 186 190
rect 184 189 185 190
rect 183 189 184 190
rect 182 189 183 190
rect 181 189 182 190
rect 180 189 181 190
rect 179 189 180 190
rect 178 189 179 190
rect 177 189 178 190
rect 176 189 177 190
rect 175 189 176 190
rect 174 189 175 190
rect 173 189 174 190
rect 172 189 173 190
rect 171 189 172 190
rect 170 189 171 190
rect 169 189 170 190
rect 168 189 169 190
rect 167 189 168 190
rect 166 189 167 190
rect 165 189 166 190
rect 164 189 165 190
rect 163 189 164 190
rect 162 189 163 190
rect 161 189 162 190
rect 160 189 161 190
rect 159 189 160 190
rect 158 189 159 190
rect 157 189 158 190
rect 156 189 157 190
rect 155 189 156 190
rect 154 189 155 190
rect 153 189 154 190
rect 152 189 153 190
rect 151 189 152 190
rect 150 189 151 190
rect 149 189 150 190
rect 148 189 149 190
rect 147 189 148 190
rect 146 189 147 190
rect 145 189 146 190
rect 144 189 145 190
rect 143 189 144 190
rect 142 189 143 190
rect 141 189 142 190
rect 140 189 141 190
rect 139 189 140 190
rect 138 189 139 190
rect 137 189 138 190
rect 136 189 137 190
rect 135 189 136 190
rect 134 189 135 190
rect 133 189 134 190
rect 132 189 133 190
rect 131 189 132 190
rect 130 189 131 190
rect 129 189 130 190
rect 128 189 129 190
rect 127 189 128 190
rect 126 189 127 190
rect 125 189 126 190
rect 124 189 125 190
rect 123 189 124 190
rect 122 189 123 190
rect 121 189 122 190
rect 120 189 121 190
rect 119 189 120 190
rect 118 189 119 190
rect 117 189 118 190
rect 116 189 117 190
rect 115 189 116 190
rect 114 189 115 190
rect 113 189 114 190
rect 112 189 113 190
rect 111 189 112 190
rect 110 189 111 190
rect 109 189 110 190
rect 108 189 109 190
rect 107 189 108 190
rect 106 189 107 190
rect 105 189 106 190
rect 104 189 105 190
rect 103 189 104 190
rect 102 189 103 190
rect 101 189 102 190
rect 100 189 101 190
rect 99 189 100 190
rect 98 189 99 190
rect 97 189 98 190
rect 96 189 97 190
rect 95 189 96 190
rect 94 189 95 190
rect 93 189 94 190
rect 92 189 93 190
rect 91 189 92 190
rect 90 189 91 190
rect 89 189 90 190
rect 88 189 89 190
rect 87 189 88 190
rect 86 189 87 190
rect 85 189 86 190
rect 84 189 85 190
rect 83 189 84 190
rect 82 189 83 190
rect 81 189 82 190
rect 80 189 81 190
rect 79 189 80 190
rect 78 189 79 190
rect 77 189 78 190
rect 76 189 77 190
rect 75 189 76 190
rect 74 189 75 190
rect 73 189 74 190
rect 72 189 73 190
rect 71 189 72 190
rect 70 189 71 190
rect 69 189 70 190
rect 68 189 69 190
rect 67 189 68 190
rect 26 189 27 190
rect 25 189 26 190
rect 24 189 25 190
rect 23 189 24 190
rect 22 189 23 190
rect 21 189 22 190
rect 20 189 21 190
rect 19 189 20 190
rect 18 189 19 190
rect 17 189 18 190
rect 16 189 17 190
rect 15 189 16 190
rect 14 189 15 190
rect 13 189 14 190
rect 12 189 13 190
rect 11 189 12 190
rect 10 189 11 190
rect 478 190 479 191
rect 477 190 478 191
rect 458 190 459 191
rect 436 190 437 191
rect 435 190 436 191
rect 434 190 435 191
rect 433 190 434 191
rect 432 190 433 191
rect 431 190 432 191
rect 430 190 431 191
rect 429 190 430 191
rect 428 190 429 191
rect 427 190 428 191
rect 426 190 427 191
rect 425 190 426 191
rect 424 190 425 191
rect 423 190 424 191
rect 422 190 423 191
rect 397 190 398 191
rect 396 190 397 191
rect 395 190 396 191
rect 394 190 395 191
rect 393 190 394 191
rect 339 190 340 191
rect 338 190 339 191
rect 337 190 338 191
rect 336 190 337 191
rect 335 190 336 191
rect 334 190 335 191
rect 333 190 334 191
rect 332 190 333 191
rect 331 190 332 191
rect 330 190 331 191
rect 329 190 330 191
rect 328 190 329 191
rect 327 190 328 191
rect 326 190 327 191
rect 325 190 326 191
rect 324 190 325 191
rect 323 190 324 191
rect 322 190 323 191
rect 321 190 322 191
rect 320 190 321 191
rect 319 190 320 191
rect 318 190 319 191
rect 317 190 318 191
rect 316 190 317 191
rect 315 190 316 191
rect 314 190 315 191
rect 313 190 314 191
rect 312 190 313 191
rect 311 190 312 191
rect 310 190 311 191
rect 309 190 310 191
rect 308 190 309 191
rect 307 190 308 191
rect 306 190 307 191
rect 305 190 306 191
rect 304 190 305 191
rect 303 190 304 191
rect 302 190 303 191
rect 301 190 302 191
rect 300 190 301 191
rect 299 190 300 191
rect 298 190 299 191
rect 297 190 298 191
rect 296 190 297 191
rect 295 190 296 191
rect 294 190 295 191
rect 293 190 294 191
rect 292 190 293 191
rect 291 190 292 191
rect 290 190 291 191
rect 289 190 290 191
rect 288 190 289 191
rect 287 190 288 191
rect 286 190 287 191
rect 285 190 286 191
rect 284 190 285 191
rect 283 190 284 191
rect 282 190 283 191
rect 281 190 282 191
rect 280 190 281 191
rect 279 190 280 191
rect 278 190 279 191
rect 277 190 278 191
rect 276 190 277 191
rect 275 190 276 191
rect 274 190 275 191
rect 273 190 274 191
rect 272 190 273 191
rect 271 190 272 191
rect 270 190 271 191
rect 253 190 254 191
rect 252 190 253 191
rect 251 190 252 191
rect 250 190 251 191
rect 249 190 250 191
rect 248 190 249 191
rect 247 190 248 191
rect 246 190 247 191
rect 245 190 246 191
rect 244 190 245 191
rect 243 190 244 191
rect 242 190 243 191
rect 241 190 242 191
rect 240 190 241 191
rect 239 190 240 191
rect 238 190 239 191
rect 237 190 238 191
rect 236 190 237 191
rect 235 190 236 191
rect 234 190 235 191
rect 233 190 234 191
rect 232 190 233 191
rect 231 190 232 191
rect 230 190 231 191
rect 229 190 230 191
rect 228 190 229 191
rect 227 190 228 191
rect 226 190 227 191
rect 225 190 226 191
rect 224 190 225 191
rect 223 190 224 191
rect 222 190 223 191
rect 221 190 222 191
rect 220 190 221 191
rect 219 190 220 191
rect 218 190 219 191
rect 217 190 218 191
rect 216 190 217 191
rect 215 190 216 191
rect 214 190 215 191
rect 213 190 214 191
rect 189 190 190 191
rect 188 190 189 191
rect 187 190 188 191
rect 186 190 187 191
rect 185 190 186 191
rect 184 190 185 191
rect 183 190 184 191
rect 182 190 183 191
rect 181 190 182 191
rect 180 190 181 191
rect 179 190 180 191
rect 178 190 179 191
rect 177 190 178 191
rect 176 190 177 191
rect 175 190 176 191
rect 174 190 175 191
rect 173 190 174 191
rect 172 190 173 191
rect 171 190 172 191
rect 170 190 171 191
rect 169 190 170 191
rect 168 190 169 191
rect 167 190 168 191
rect 166 190 167 191
rect 165 190 166 191
rect 164 190 165 191
rect 163 190 164 191
rect 162 190 163 191
rect 161 190 162 191
rect 160 190 161 191
rect 159 190 160 191
rect 158 190 159 191
rect 157 190 158 191
rect 156 190 157 191
rect 155 190 156 191
rect 154 190 155 191
rect 153 190 154 191
rect 152 190 153 191
rect 151 190 152 191
rect 150 190 151 191
rect 149 190 150 191
rect 148 190 149 191
rect 147 190 148 191
rect 146 190 147 191
rect 145 190 146 191
rect 144 190 145 191
rect 143 190 144 191
rect 142 190 143 191
rect 141 190 142 191
rect 140 190 141 191
rect 139 190 140 191
rect 138 190 139 191
rect 137 190 138 191
rect 136 190 137 191
rect 135 190 136 191
rect 134 190 135 191
rect 133 190 134 191
rect 132 190 133 191
rect 131 190 132 191
rect 130 190 131 191
rect 129 190 130 191
rect 128 190 129 191
rect 127 190 128 191
rect 126 190 127 191
rect 125 190 126 191
rect 124 190 125 191
rect 123 190 124 191
rect 122 190 123 191
rect 121 190 122 191
rect 120 190 121 191
rect 119 190 120 191
rect 118 190 119 191
rect 117 190 118 191
rect 116 190 117 191
rect 115 190 116 191
rect 114 190 115 191
rect 113 190 114 191
rect 112 190 113 191
rect 111 190 112 191
rect 110 190 111 191
rect 109 190 110 191
rect 108 190 109 191
rect 107 190 108 191
rect 106 190 107 191
rect 105 190 106 191
rect 104 190 105 191
rect 103 190 104 191
rect 102 190 103 191
rect 101 190 102 191
rect 100 190 101 191
rect 99 190 100 191
rect 98 190 99 191
rect 97 190 98 191
rect 96 190 97 191
rect 95 190 96 191
rect 94 190 95 191
rect 93 190 94 191
rect 92 190 93 191
rect 91 190 92 191
rect 90 190 91 191
rect 89 190 90 191
rect 88 190 89 191
rect 87 190 88 191
rect 86 190 87 191
rect 85 190 86 191
rect 84 190 85 191
rect 83 190 84 191
rect 82 190 83 191
rect 81 190 82 191
rect 80 190 81 191
rect 79 190 80 191
rect 78 190 79 191
rect 77 190 78 191
rect 76 190 77 191
rect 75 190 76 191
rect 74 190 75 191
rect 73 190 74 191
rect 72 190 73 191
rect 71 190 72 191
rect 70 190 71 191
rect 69 190 70 191
rect 68 190 69 191
rect 67 190 68 191
rect 26 190 27 191
rect 25 190 26 191
rect 24 190 25 191
rect 23 190 24 191
rect 22 190 23 191
rect 21 190 22 191
rect 20 190 21 191
rect 19 190 20 191
rect 18 190 19 191
rect 17 190 18 191
rect 16 190 17 191
rect 15 190 16 191
rect 14 190 15 191
rect 13 190 14 191
rect 12 190 13 191
rect 11 190 12 191
rect 10 190 11 191
rect 478 191 479 192
rect 477 191 478 192
rect 476 191 477 192
rect 475 191 476 192
rect 474 191 475 192
rect 473 191 474 192
rect 472 191 473 192
rect 471 191 472 192
rect 470 191 471 192
rect 469 191 470 192
rect 468 191 469 192
rect 467 191 468 192
rect 466 191 467 192
rect 465 191 466 192
rect 464 191 465 192
rect 463 191 464 192
rect 462 191 463 192
rect 461 191 462 192
rect 460 191 461 192
rect 459 191 460 192
rect 458 191 459 192
rect 438 191 439 192
rect 437 191 438 192
rect 436 191 437 192
rect 435 191 436 192
rect 434 191 435 192
rect 433 191 434 192
rect 432 191 433 192
rect 431 191 432 192
rect 430 191 431 192
rect 429 191 430 192
rect 428 191 429 192
rect 427 191 428 192
rect 426 191 427 192
rect 425 191 426 192
rect 424 191 425 192
rect 423 191 424 192
rect 403 191 404 192
rect 402 191 403 192
rect 401 191 402 192
rect 400 191 401 192
rect 399 191 400 192
rect 398 191 399 192
rect 397 191 398 192
rect 396 191 397 192
rect 395 191 396 192
rect 394 191 395 192
rect 393 191 394 192
rect 340 191 341 192
rect 339 191 340 192
rect 338 191 339 192
rect 337 191 338 192
rect 336 191 337 192
rect 335 191 336 192
rect 334 191 335 192
rect 333 191 334 192
rect 332 191 333 192
rect 331 191 332 192
rect 330 191 331 192
rect 329 191 330 192
rect 328 191 329 192
rect 327 191 328 192
rect 326 191 327 192
rect 325 191 326 192
rect 324 191 325 192
rect 323 191 324 192
rect 322 191 323 192
rect 321 191 322 192
rect 320 191 321 192
rect 319 191 320 192
rect 318 191 319 192
rect 317 191 318 192
rect 316 191 317 192
rect 315 191 316 192
rect 314 191 315 192
rect 313 191 314 192
rect 312 191 313 192
rect 311 191 312 192
rect 310 191 311 192
rect 309 191 310 192
rect 308 191 309 192
rect 307 191 308 192
rect 306 191 307 192
rect 305 191 306 192
rect 304 191 305 192
rect 303 191 304 192
rect 302 191 303 192
rect 301 191 302 192
rect 300 191 301 192
rect 299 191 300 192
rect 298 191 299 192
rect 297 191 298 192
rect 296 191 297 192
rect 295 191 296 192
rect 294 191 295 192
rect 293 191 294 192
rect 292 191 293 192
rect 291 191 292 192
rect 290 191 291 192
rect 289 191 290 192
rect 288 191 289 192
rect 287 191 288 192
rect 286 191 287 192
rect 285 191 286 192
rect 284 191 285 192
rect 283 191 284 192
rect 282 191 283 192
rect 281 191 282 192
rect 280 191 281 192
rect 279 191 280 192
rect 278 191 279 192
rect 277 191 278 192
rect 276 191 277 192
rect 275 191 276 192
rect 274 191 275 192
rect 273 191 274 192
rect 272 191 273 192
rect 271 191 272 192
rect 270 191 271 192
rect 269 191 270 192
rect 252 191 253 192
rect 251 191 252 192
rect 250 191 251 192
rect 249 191 250 192
rect 248 191 249 192
rect 247 191 248 192
rect 246 191 247 192
rect 245 191 246 192
rect 244 191 245 192
rect 243 191 244 192
rect 242 191 243 192
rect 241 191 242 192
rect 240 191 241 192
rect 239 191 240 192
rect 238 191 239 192
rect 237 191 238 192
rect 236 191 237 192
rect 235 191 236 192
rect 234 191 235 192
rect 233 191 234 192
rect 232 191 233 192
rect 231 191 232 192
rect 230 191 231 192
rect 229 191 230 192
rect 228 191 229 192
rect 227 191 228 192
rect 226 191 227 192
rect 225 191 226 192
rect 224 191 225 192
rect 223 191 224 192
rect 222 191 223 192
rect 221 191 222 192
rect 220 191 221 192
rect 219 191 220 192
rect 218 191 219 192
rect 217 191 218 192
rect 216 191 217 192
rect 215 191 216 192
rect 214 191 215 192
rect 213 191 214 192
rect 212 191 213 192
rect 188 191 189 192
rect 187 191 188 192
rect 186 191 187 192
rect 185 191 186 192
rect 184 191 185 192
rect 183 191 184 192
rect 182 191 183 192
rect 181 191 182 192
rect 180 191 181 192
rect 179 191 180 192
rect 178 191 179 192
rect 177 191 178 192
rect 176 191 177 192
rect 175 191 176 192
rect 174 191 175 192
rect 173 191 174 192
rect 172 191 173 192
rect 171 191 172 192
rect 170 191 171 192
rect 169 191 170 192
rect 168 191 169 192
rect 167 191 168 192
rect 166 191 167 192
rect 165 191 166 192
rect 164 191 165 192
rect 163 191 164 192
rect 162 191 163 192
rect 161 191 162 192
rect 160 191 161 192
rect 159 191 160 192
rect 158 191 159 192
rect 157 191 158 192
rect 156 191 157 192
rect 155 191 156 192
rect 154 191 155 192
rect 153 191 154 192
rect 152 191 153 192
rect 151 191 152 192
rect 150 191 151 192
rect 149 191 150 192
rect 148 191 149 192
rect 147 191 148 192
rect 146 191 147 192
rect 145 191 146 192
rect 144 191 145 192
rect 143 191 144 192
rect 142 191 143 192
rect 141 191 142 192
rect 140 191 141 192
rect 139 191 140 192
rect 138 191 139 192
rect 137 191 138 192
rect 136 191 137 192
rect 135 191 136 192
rect 134 191 135 192
rect 133 191 134 192
rect 132 191 133 192
rect 131 191 132 192
rect 130 191 131 192
rect 129 191 130 192
rect 128 191 129 192
rect 127 191 128 192
rect 126 191 127 192
rect 125 191 126 192
rect 124 191 125 192
rect 123 191 124 192
rect 122 191 123 192
rect 121 191 122 192
rect 120 191 121 192
rect 119 191 120 192
rect 118 191 119 192
rect 117 191 118 192
rect 116 191 117 192
rect 115 191 116 192
rect 114 191 115 192
rect 113 191 114 192
rect 112 191 113 192
rect 111 191 112 192
rect 110 191 111 192
rect 109 191 110 192
rect 108 191 109 192
rect 107 191 108 192
rect 106 191 107 192
rect 105 191 106 192
rect 104 191 105 192
rect 103 191 104 192
rect 102 191 103 192
rect 101 191 102 192
rect 100 191 101 192
rect 99 191 100 192
rect 98 191 99 192
rect 97 191 98 192
rect 96 191 97 192
rect 95 191 96 192
rect 94 191 95 192
rect 93 191 94 192
rect 92 191 93 192
rect 91 191 92 192
rect 90 191 91 192
rect 89 191 90 192
rect 88 191 89 192
rect 87 191 88 192
rect 86 191 87 192
rect 85 191 86 192
rect 84 191 85 192
rect 83 191 84 192
rect 82 191 83 192
rect 81 191 82 192
rect 80 191 81 192
rect 79 191 80 192
rect 78 191 79 192
rect 77 191 78 192
rect 76 191 77 192
rect 75 191 76 192
rect 74 191 75 192
rect 73 191 74 192
rect 72 191 73 192
rect 71 191 72 192
rect 70 191 71 192
rect 69 191 70 192
rect 68 191 69 192
rect 48 191 49 192
rect 47 191 48 192
rect 46 191 47 192
rect 27 191 28 192
rect 26 191 27 192
rect 25 191 26 192
rect 24 191 25 192
rect 23 191 24 192
rect 22 191 23 192
rect 21 191 22 192
rect 20 191 21 192
rect 19 191 20 192
rect 18 191 19 192
rect 17 191 18 192
rect 16 191 17 192
rect 15 191 16 192
rect 14 191 15 192
rect 13 191 14 192
rect 12 191 13 192
rect 11 191 12 192
rect 10 191 11 192
rect 478 192 479 193
rect 477 192 478 193
rect 476 192 477 193
rect 475 192 476 193
rect 474 192 475 193
rect 473 192 474 193
rect 472 192 473 193
rect 471 192 472 193
rect 470 192 471 193
rect 469 192 470 193
rect 468 192 469 193
rect 467 192 468 193
rect 466 192 467 193
rect 465 192 466 193
rect 464 192 465 193
rect 463 192 464 193
rect 462 192 463 193
rect 461 192 462 193
rect 460 192 461 193
rect 459 192 460 193
rect 458 192 459 193
rect 438 192 439 193
rect 437 192 438 193
rect 436 192 437 193
rect 435 192 436 193
rect 434 192 435 193
rect 433 192 434 193
rect 432 192 433 193
rect 431 192 432 193
rect 430 192 431 193
rect 429 192 430 193
rect 428 192 429 193
rect 427 192 428 193
rect 426 192 427 193
rect 425 192 426 193
rect 424 192 425 193
rect 423 192 424 193
rect 422 192 423 193
rect 421 192 422 193
rect 420 192 421 193
rect 419 192 420 193
rect 418 192 419 193
rect 417 192 418 193
rect 416 192 417 193
rect 415 192 416 193
rect 414 192 415 193
rect 413 192 414 193
rect 412 192 413 193
rect 411 192 412 193
rect 410 192 411 193
rect 409 192 410 193
rect 408 192 409 193
rect 407 192 408 193
rect 406 192 407 193
rect 405 192 406 193
rect 404 192 405 193
rect 403 192 404 193
rect 402 192 403 193
rect 401 192 402 193
rect 400 192 401 193
rect 399 192 400 193
rect 398 192 399 193
rect 397 192 398 193
rect 396 192 397 193
rect 395 192 396 193
rect 394 192 395 193
rect 393 192 394 193
rect 341 192 342 193
rect 340 192 341 193
rect 339 192 340 193
rect 338 192 339 193
rect 337 192 338 193
rect 336 192 337 193
rect 335 192 336 193
rect 334 192 335 193
rect 333 192 334 193
rect 332 192 333 193
rect 331 192 332 193
rect 330 192 331 193
rect 329 192 330 193
rect 328 192 329 193
rect 327 192 328 193
rect 326 192 327 193
rect 325 192 326 193
rect 324 192 325 193
rect 323 192 324 193
rect 322 192 323 193
rect 321 192 322 193
rect 320 192 321 193
rect 319 192 320 193
rect 318 192 319 193
rect 317 192 318 193
rect 316 192 317 193
rect 315 192 316 193
rect 314 192 315 193
rect 313 192 314 193
rect 312 192 313 193
rect 311 192 312 193
rect 310 192 311 193
rect 309 192 310 193
rect 308 192 309 193
rect 307 192 308 193
rect 306 192 307 193
rect 305 192 306 193
rect 304 192 305 193
rect 303 192 304 193
rect 302 192 303 193
rect 301 192 302 193
rect 300 192 301 193
rect 299 192 300 193
rect 298 192 299 193
rect 297 192 298 193
rect 296 192 297 193
rect 295 192 296 193
rect 294 192 295 193
rect 293 192 294 193
rect 292 192 293 193
rect 291 192 292 193
rect 290 192 291 193
rect 289 192 290 193
rect 288 192 289 193
rect 287 192 288 193
rect 286 192 287 193
rect 285 192 286 193
rect 284 192 285 193
rect 283 192 284 193
rect 282 192 283 193
rect 281 192 282 193
rect 280 192 281 193
rect 279 192 280 193
rect 278 192 279 193
rect 277 192 278 193
rect 276 192 277 193
rect 275 192 276 193
rect 274 192 275 193
rect 273 192 274 193
rect 272 192 273 193
rect 271 192 272 193
rect 270 192 271 193
rect 269 192 270 193
rect 268 192 269 193
rect 267 192 268 193
rect 252 192 253 193
rect 251 192 252 193
rect 250 192 251 193
rect 249 192 250 193
rect 248 192 249 193
rect 247 192 248 193
rect 246 192 247 193
rect 245 192 246 193
rect 244 192 245 193
rect 243 192 244 193
rect 242 192 243 193
rect 241 192 242 193
rect 240 192 241 193
rect 239 192 240 193
rect 238 192 239 193
rect 237 192 238 193
rect 236 192 237 193
rect 235 192 236 193
rect 234 192 235 193
rect 233 192 234 193
rect 232 192 233 193
rect 231 192 232 193
rect 230 192 231 193
rect 229 192 230 193
rect 228 192 229 193
rect 227 192 228 193
rect 226 192 227 193
rect 225 192 226 193
rect 224 192 225 193
rect 223 192 224 193
rect 222 192 223 193
rect 221 192 222 193
rect 220 192 221 193
rect 219 192 220 193
rect 218 192 219 193
rect 217 192 218 193
rect 216 192 217 193
rect 215 192 216 193
rect 214 192 215 193
rect 213 192 214 193
rect 212 192 213 193
rect 187 192 188 193
rect 186 192 187 193
rect 185 192 186 193
rect 184 192 185 193
rect 183 192 184 193
rect 182 192 183 193
rect 181 192 182 193
rect 180 192 181 193
rect 179 192 180 193
rect 178 192 179 193
rect 177 192 178 193
rect 176 192 177 193
rect 175 192 176 193
rect 174 192 175 193
rect 173 192 174 193
rect 172 192 173 193
rect 171 192 172 193
rect 170 192 171 193
rect 169 192 170 193
rect 168 192 169 193
rect 167 192 168 193
rect 166 192 167 193
rect 165 192 166 193
rect 164 192 165 193
rect 163 192 164 193
rect 162 192 163 193
rect 161 192 162 193
rect 160 192 161 193
rect 159 192 160 193
rect 158 192 159 193
rect 157 192 158 193
rect 156 192 157 193
rect 155 192 156 193
rect 154 192 155 193
rect 153 192 154 193
rect 152 192 153 193
rect 151 192 152 193
rect 150 192 151 193
rect 149 192 150 193
rect 148 192 149 193
rect 147 192 148 193
rect 146 192 147 193
rect 145 192 146 193
rect 144 192 145 193
rect 143 192 144 193
rect 142 192 143 193
rect 141 192 142 193
rect 140 192 141 193
rect 139 192 140 193
rect 138 192 139 193
rect 137 192 138 193
rect 136 192 137 193
rect 135 192 136 193
rect 134 192 135 193
rect 133 192 134 193
rect 132 192 133 193
rect 131 192 132 193
rect 130 192 131 193
rect 129 192 130 193
rect 128 192 129 193
rect 127 192 128 193
rect 126 192 127 193
rect 125 192 126 193
rect 124 192 125 193
rect 123 192 124 193
rect 122 192 123 193
rect 121 192 122 193
rect 120 192 121 193
rect 119 192 120 193
rect 118 192 119 193
rect 117 192 118 193
rect 116 192 117 193
rect 115 192 116 193
rect 114 192 115 193
rect 113 192 114 193
rect 112 192 113 193
rect 111 192 112 193
rect 110 192 111 193
rect 109 192 110 193
rect 108 192 109 193
rect 107 192 108 193
rect 106 192 107 193
rect 105 192 106 193
rect 104 192 105 193
rect 103 192 104 193
rect 102 192 103 193
rect 101 192 102 193
rect 100 192 101 193
rect 99 192 100 193
rect 98 192 99 193
rect 97 192 98 193
rect 96 192 97 193
rect 95 192 96 193
rect 94 192 95 193
rect 93 192 94 193
rect 92 192 93 193
rect 91 192 92 193
rect 90 192 91 193
rect 89 192 90 193
rect 88 192 89 193
rect 87 192 88 193
rect 86 192 87 193
rect 85 192 86 193
rect 84 192 85 193
rect 83 192 84 193
rect 82 192 83 193
rect 81 192 82 193
rect 80 192 81 193
rect 79 192 80 193
rect 78 192 79 193
rect 77 192 78 193
rect 76 192 77 193
rect 75 192 76 193
rect 74 192 75 193
rect 73 192 74 193
rect 72 192 73 193
rect 71 192 72 193
rect 70 192 71 193
rect 69 192 70 193
rect 68 192 69 193
rect 49 192 50 193
rect 48 192 49 193
rect 47 192 48 193
rect 46 192 47 193
rect 45 192 46 193
rect 44 192 45 193
rect 29 192 30 193
rect 28 192 29 193
rect 27 192 28 193
rect 26 192 27 193
rect 25 192 26 193
rect 24 192 25 193
rect 23 192 24 193
rect 22 192 23 193
rect 21 192 22 193
rect 20 192 21 193
rect 19 192 20 193
rect 18 192 19 193
rect 17 192 18 193
rect 16 192 17 193
rect 15 192 16 193
rect 14 192 15 193
rect 13 192 14 193
rect 12 192 13 193
rect 11 192 12 193
rect 10 192 11 193
rect 478 193 479 194
rect 477 193 478 194
rect 476 193 477 194
rect 475 193 476 194
rect 474 193 475 194
rect 473 193 474 194
rect 472 193 473 194
rect 471 193 472 194
rect 470 193 471 194
rect 469 193 470 194
rect 468 193 469 194
rect 467 193 468 194
rect 466 193 467 194
rect 465 193 466 194
rect 464 193 465 194
rect 463 193 464 194
rect 462 193 463 194
rect 461 193 462 194
rect 460 193 461 194
rect 459 193 460 194
rect 458 193 459 194
rect 438 193 439 194
rect 437 193 438 194
rect 436 193 437 194
rect 435 193 436 194
rect 434 193 435 194
rect 433 193 434 194
rect 432 193 433 194
rect 431 193 432 194
rect 430 193 431 194
rect 429 193 430 194
rect 428 193 429 194
rect 427 193 428 194
rect 426 193 427 194
rect 425 193 426 194
rect 424 193 425 194
rect 423 193 424 194
rect 422 193 423 194
rect 421 193 422 194
rect 420 193 421 194
rect 419 193 420 194
rect 418 193 419 194
rect 417 193 418 194
rect 416 193 417 194
rect 415 193 416 194
rect 414 193 415 194
rect 413 193 414 194
rect 412 193 413 194
rect 411 193 412 194
rect 410 193 411 194
rect 409 193 410 194
rect 408 193 409 194
rect 407 193 408 194
rect 406 193 407 194
rect 405 193 406 194
rect 404 193 405 194
rect 403 193 404 194
rect 402 193 403 194
rect 401 193 402 194
rect 400 193 401 194
rect 399 193 400 194
rect 398 193 399 194
rect 397 193 398 194
rect 396 193 397 194
rect 395 193 396 194
rect 394 193 395 194
rect 393 193 394 194
rect 342 193 343 194
rect 341 193 342 194
rect 340 193 341 194
rect 339 193 340 194
rect 338 193 339 194
rect 337 193 338 194
rect 336 193 337 194
rect 335 193 336 194
rect 334 193 335 194
rect 333 193 334 194
rect 332 193 333 194
rect 331 193 332 194
rect 330 193 331 194
rect 329 193 330 194
rect 328 193 329 194
rect 327 193 328 194
rect 326 193 327 194
rect 325 193 326 194
rect 324 193 325 194
rect 323 193 324 194
rect 322 193 323 194
rect 321 193 322 194
rect 320 193 321 194
rect 319 193 320 194
rect 318 193 319 194
rect 317 193 318 194
rect 316 193 317 194
rect 315 193 316 194
rect 314 193 315 194
rect 313 193 314 194
rect 312 193 313 194
rect 311 193 312 194
rect 310 193 311 194
rect 309 193 310 194
rect 308 193 309 194
rect 307 193 308 194
rect 306 193 307 194
rect 305 193 306 194
rect 304 193 305 194
rect 303 193 304 194
rect 302 193 303 194
rect 301 193 302 194
rect 300 193 301 194
rect 299 193 300 194
rect 298 193 299 194
rect 297 193 298 194
rect 296 193 297 194
rect 295 193 296 194
rect 294 193 295 194
rect 293 193 294 194
rect 292 193 293 194
rect 291 193 292 194
rect 290 193 291 194
rect 289 193 290 194
rect 288 193 289 194
rect 287 193 288 194
rect 286 193 287 194
rect 285 193 286 194
rect 284 193 285 194
rect 283 193 284 194
rect 282 193 283 194
rect 281 193 282 194
rect 280 193 281 194
rect 279 193 280 194
rect 278 193 279 194
rect 277 193 278 194
rect 276 193 277 194
rect 275 193 276 194
rect 274 193 275 194
rect 273 193 274 194
rect 272 193 273 194
rect 271 193 272 194
rect 270 193 271 194
rect 269 193 270 194
rect 268 193 269 194
rect 267 193 268 194
rect 266 193 267 194
rect 251 193 252 194
rect 250 193 251 194
rect 249 193 250 194
rect 248 193 249 194
rect 247 193 248 194
rect 246 193 247 194
rect 245 193 246 194
rect 244 193 245 194
rect 243 193 244 194
rect 242 193 243 194
rect 241 193 242 194
rect 240 193 241 194
rect 239 193 240 194
rect 238 193 239 194
rect 237 193 238 194
rect 236 193 237 194
rect 235 193 236 194
rect 234 193 235 194
rect 233 193 234 194
rect 232 193 233 194
rect 231 193 232 194
rect 230 193 231 194
rect 229 193 230 194
rect 228 193 229 194
rect 227 193 228 194
rect 226 193 227 194
rect 225 193 226 194
rect 224 193 225 194
rect 223 193 224 194
rect 222 193 223 194
rect 221 193 222 194
rect 220 193 221 194
rect 219 193 220 194
rect 218 193 219 194
rect 217 193 218 194
rect 216 193 217 194
rect 215 193 216 194
rect 214 193 215 194
rect 213 193 214 194
rect 212 193 213 194
rect 211 193 212 194
rect 186 193 187 194
rect 185 193 186 194
rect 184 193 185 194
rect 183 193 184 194
rect 182 193 183 194
rect 181 193 182 194
rect 180 193 181 194
rect 179 193 180 194
rect 178 193 179 194
rect 177 193 178 194
rect 176 193 177 194
rect 175 193 176 194
rect 174 193 175 194
rect 173 193 174 194
rect 172 193 173 194
rect 171 193 172 194
rect 170 193 171 194
rect 169 193 170 194
rect 168 193 169 194
rect 167 193 168 194
rect 166 193 167 194
rect 165 193 166 194
rect 164 193 165 194
rect 163 193 164 194
rect 162 193 163 194
rect 161 193 162 194
rect 160 193 161 194
rect 159 193 160 194
rect 158 193 159 194
rect 157 193 158 194
rect 156 193 157 194
rect 155 193 156 194
rect 154 193 155 194
rect 153 193 154 194
rect 152 193 153 194
rect 151 193 152 194
rect 150 193 151 194
rect 149 193 150 194
rect 148 193 149 194
rect 147 193 148 194
rect 146 193 147 194
rect 145 193 146 194
rect 144 193 145 194
rect 143 193 144 194
rect 142 193 143 194
rect 141 193 142 194
rect 140 193 141 194
rect 139 193 140 194
rect 138 193 139 194
rect 137 193 138 194
rect 136 193 137 194
rect 135 193 136 194
rect 134 193 135 194
rect 133 193 134 194
rect 132 193 133 194
rect 131 193 132 194
rect 130 193 131 194
rect 129 193 130 194
rect 128 193 129 194
rect 127 193 128 194
rect 126 193 127 194
rect 125 193 126 194
rect 124 193 125 194
rect 123 193 124 194
rect 122 193 123 194
rect 121 193 122 194
rect 120 193 121 194
rect 119 193 120 194
rect 118 193 119 194
rect 117 193 118 194
rect 116 193 117 194
rect 115 193 116 194
rect 114 193 115 194
rect 113 193 114 194
rect 112 193 113 194
rect 111 193 112 194
rect 110 193 111 194
rect 109 193 110 194
rect 108 193 109 194
rect 107 193 108 194
rect 106 193 107 194
rect 105 193 106 194
rect 104 193 105 194
rect 103 193 104 194
rect 102 193 103 194
rect 101 193 102 194
rect 100 193 101 194
rect 99 193 100 194
rect 98 193 99 194
rect 97 193 98 194
rect 96 193 97 194
rect 95 193 96 194
rect 94 193 95 194
rect 93 193 94 194
rect 92 193 93 194
rect 91 193 92 194
rect 90 193 91 194
rect 89 193 90 194
rect 88 193 89 194
rect 87 193 88 194
rect 86 193 87 194
rect 85 193 86 194
rect 84 193 85 194
rect 83 193 84 194
rect 82 193 83 194
rect 81 193 82 194
rect 80 193 81 194
rect 79 193 80 194
rect 78 193 79 194
rect 77 193 78 194
rect 76 193 77 194
rect 75 193 76 194
rect 74 193 75 194
rect 73 193 74 194
rect 72 193 73 194
rect 71 193 72 194
rect 70 193 71 194
rect 69 193 70 194
rect 68 193 69 194
rect 49 193 50 194
rect 48 193 49 194
rect 47 193 48 194
rect 46 193 47 194
rect 45 193 46 194
rect 44 193 45 194
rect 43 193 44 194
rect 42 193 43 194
rect 30 193 31 194
rect 29 193 30 194
rect 28 193 29 194
rect 27 193 28 194
rect 26 193 27 194
rect 25 193 26 194
rect 24 193 25 194
rect 23 193 24 194
rect 22 193 23 194
rect 21 193 22 194
rect 20 193 21 194
rect 19 193 20 194
rect 18 193 19 194
rect 17 193 18 194
rect 16 193 17 194
rect 15 193 16 194
rect 14 193 15 194
rect 13 193 14 194
rect 12 193 13 194
rect 11 193 12 194
rect 10 193 11 194
rect 478 194 479 195
rect 477 194 478 195
rect 476 194 477 195
rect 475 194 476 195
rect 474 194 475 195
rect 473 194 474 195
rect 472 194 473 195
rect 471 194 472 195
rect 470 194 471 195
rect 469 194 470 195
rect 468 194 469 195
rect 467 194 468 195
rect 466 194 467 195
rect 465 194 466 195
rect 464 194 465 195
rect 463 194 464 195
rect 462 194 463 195
rect 461 194 462 195
rect 460 194 461 195
rect 459 194 460 195
rect 458 194 459 195
rect 438 194 439 195
rect 437 194 438 195
rect 436 194 437 195
rect 435 194 436 195
rect 434 194 435 195
rect 433 194 434 195
rect 432 194 433 195
rect 431 194 432 195
rect 430 194 431 195
rect 429 194 430 195
rect 428 194 429 195
rect 427 194 428 195
rect 426 194 427 195
rect 425 194 426 195
rect 424 194 425 195
rect 423 194 424 195
rect 422 194 423 195
rect 421 194 422 195
rect 420 194 421 195
rect 419 194 420 195
rect 418 194 419 195
rect 417 194 418 195
rect 416 194 417 195
rect 415 194 416 195
rect 414 194 415 195
rect 413 194 414 195
rect 412 194 413 195
rect 411 194 412 195
rect 410 194 411 195
rect 409 194 410 195
rect 408 194 409 195
rect 407 194 408 195
rect 406 194 407 195
rect 405 194 406 195
rect 404 194 405 195
rect 403 194 404 195
rect 402 194 403 195
rect 401 194 402 195
rect 400 194 401 195
rect 399 194 400 195
rect 398 194 399 195
rect 397 194 398 195
rect 396 194 397 195
rect 395 194 396 195
rect 394 194 395 195
rect 393 194 394 195
rect 343 194 344 195
rect 342 194 343 195
rect 341 194 342 195
rect 340 194 341 195
rect 339 194 340 195
rect 338 194 339 195
rect 337 194 338 195
rect 336 194 337 195
rect 335 194 336 195
rect 334 194 335 195
rect 333 194 334 195
rect 332 194 333 195
rect 331 194 332 195
rect 330 194 331 195
rect 329 194 330 195
rect 328 194 329 195
rect 327 194 328 195
rect 326 194 327 195
rect 325 194 326 195
rect 324 194 325 195
rect 323 194 324 195
rect 322 194 323 195
rect 321 194 322 195
rect 320 194 321 195
rect 319 194 320 195
rect 318 194 319 195
rect 317 194 318 195
rect 316 194 317 195
rect 315 194 316 195
rect 314 194 315 195
rect 313 194 314 195
rect 312 194 313 195
rect 311 194 312 195
rect 310 194 311 195
rect 309 194 310 195
rect 308 194 309 195
rect 307 194 308 195
rect 306 194 307 195
rect 305 194 306 195
rect 304 194 305 195
rect 303 194 304 195
rect 302 194 303 195
rect 301 194 302 195
rect 300 194 301 195
rect 299 194 300 195
rect 298 194 299 195
rect 297 194 298 195
rect 296 194 297 195
rect 295 194 296 195
rect 294 194 295 195
rect 293 194 294 195
rect 292 194 293 195
rect 291 194 292 195
rect 290 194 291 195
rect 289 194 290 195
rect 288 194 289 195
rect 287 194 288 195
rect 286 194 287 195
rect 285 194 286 195
rect 284 194 285 195
rect 283 194 284 195
rect 282 194 283 195
rect 281 194 282 195
rect 280 194 281 195
rect 279 194 280 195
rect 278 194 279 195
rect 277 194 278 195
rect 276 194 277 195
rect 275 194 276 195
rect 274 194 275 195
rect 273 194 274 195
rect 272 194 273 195
rect 271 194 272 195
rect 270 194 271 195
rect 269 194 270 195
rect 268 194 269 195
rect 267 194 268 195
rect 266 194 267 195
rect 265 194 266 195
rect 250 194 251 195
rect 249 194 250 195
rect 248 194 249 195
rect 247 194 248 195
rect 246 194 247 195
rect 245 194 246 195
rect 244 194 245 195
rect 243 194 244 195
rect 242 194 243 195
rect 241 194 242 195
rect 240 194 241 195
rect 239 194 240 195
rect 238 194 239 195
rect 237 194 238 195
rect 236 194 237 195
rect 235 194 236 195
rect 234 194 235 195
rect 233 194 234 195
rect 232 194 233 195
rect 231 194 232 195
rect 230 194 231 195
rect 229 194 230 195
rect 228 194 229 195
rect 227 194 228 195
rect 226 194 227 195
rect 225 194 226 195
rect 224 194 225 195
rect 223 194 224 195
rect 222 194 223 195
rect 221 194 222 195
rect 220 194 221 195
rect 219 194 220 195
rect 218 194 219 195
rect 217 194 218 195
rect 216 194 217 195
rect 215 194 216 195
rect 214 194 215 195
rect 213 194 214 195
rect 212 194 213 195
rect 211 194 212 195
rect 210 194 211 195
rect 185 194 186 195
rect 184 194 185 195
rect 183 194 184 195
rect 182 194 183 195
rect 181 194 182 195
rect 180 194 181 195
rect 179 194 180 195
rect 178 194 179 195
rect 177 194 178 195
rect 176 194 177 195
rect 175 194 176 195
rect 174 194 175 195
rect 173 194 174 195
rect 172 194 173 195
rect 171 194 172 195
rect 170 194 171 195
rect 169 194 170 195
rect 168 194 169 195
rect 167 194 168 195
rect 166 194 167 195
rect 165 194 166 195
rect 164 194 165 195
rect 163 194 164 195
rect 162 194 163 195
rect 161 194 162 195
rect 160 194 161 195
rect 159 194 160 195
rect 158 194 159 195
rect 157 194 158 195
rect 156 194 157 195
rect 155 194 156 195
rect 154 194 155 195
rect 153 194 154 195
rect 152 194 153 195
rect 151 194 152 195
rect 150 194 151 195
rect 149 194 150 195
rect 148 194 149 195
rect 147 194 148 195
rect 146 194 147 195
rect 145 194 146 195
rect 144 194 145 195
rect 143 194 144 195
rect 142 194 143 195
rect 141 194 142 195
rect 140 194 141 195
rect 139 194 140 195
rect 138 194 139 195
rect 137 194 138 195
rect 136 194 137 195
rect 135 194 136 195
rect 134 194 135 195
rect 133 194 134 195
rect 132 194 133 195
rect 131 194 132 195
rect 130 194 131 195
rect 129 194 130 195
rect 128 194 129 195
rect 127 194 128 195
rect 126 194 127 195
rect 125 194 126 195
rect 124 194 125 195
rect 123 194 124 195
rect 122 194 123 195
rect 121 194 122 195
rect 120 194 121 195
rect 119 194 120 195
rect 118 194 119 195
rect 117 194 118 195
rect 116 194 117 195
rect 115 194 116 195
rect 114 194 115 195
rect 113 194 114 195
rect 112 194 113 195
rect 111 194 112 195
rect 110 194 111 195
rect 109 194 110 195
rect 108 194 109 195
rect 107 194 108 195
rect 106 194 107 195
rect 105 194 106 195
rect 104 194 105 195
rect 103 194 104 195
rect 102 194 103 195
rect 101 194 102 195
rect 100 194 101 195
rect 99 194 100 195
rect 98 194 99 195
rect 97 194 98 195
rect 96 194 97 195
rect 95 194 96 195
rect 94 194 95 195
rect 93 194 94 195
rect 92 194 93 195
rect 91 194 92 195
rect 90 194 91 195
rect 89 194 90 195
rect 88 194 89 195
rect 87 194 88 195
rect 86 194 87 195
rect 85 194 86 195
rect 84 194 85 195
rect 83 194 84 195
rect 82 194 83 195
rect 81 194 82 195
rect 80 194 81 195
rect 79 194 80 195
rect 78 194 79 195
rect 77 194 78 195
rect 76 194 77 195
rect 75 194 76 195
rect 74 194 75 195
rect 73 194 74 195
rect 72 194 73 195
rect 71 194 72 195
rect 70 194 71 195
rect 69 194 70 195
rect 68 194 69 195
rect 50 194 51 195
rect 49 194 50 195
rect 48 194 49 195
rect 47 194 48 195
rect 46 194 47 195
rect 45 194 46 195
rect 44 194 45 195
rect 43 194 44 195
rect 42 194 43 195
rect 41 194 42 195
rect 40 194 41 195
rect 39 194 40 195
rect 38 194 39 195
rect 33 194 34 195
rect 32 194 33 195
rect 31 194 32 195
rect 30 194 31 195
rect 29 194 30 195
rect 28 194 29 195
rect 27 194 28 195
rect 26 194 27 195
rect 25 194 26 195
rect 24 194 25 195
rect 23 194 24 195
rect 22 194 23 195
rect 21 194 22 195
rect 20 194 21 195
rect 19 194 20 195
rect 18 194 19 195
rect 17 194 18 195
rect 16 194 17 195
rect 15 194 16 195
rect 14 194 15 195
rect 13 194 14 195
rect 12 194 13 195
rect 11 194 12 195
rect 10 194 11 195
rect 478 195 479 196
rect 477 195 478 196
rect 476 195 477 196
rect 475 195 476 196
rect 474 195 475 196
rect 473 195 474 196
rect 472 195 473 196
rect 471 195 472 196
rect 470 195 471 196
rect 469 195 470 196
rect 468 195 469 196
rect 467 195 468 196
rect 466 195 467 196
rect 465 195 466 196
rect 464 195 465 196
rect 463 195 464 196
rect 462 195 463 196
rect 461 195 462 196
rect 460 195 461 196
rect 459 195 460 196
rect 458 195 459 196
rect 403 195 404 196
rect 402 195 403 196
rect 401 195 402 196
rect 400 195 401 196
rect 399 195 400 196
rect 398 195 399 196
rect 397 195 398 196
rect 396 195 397 196
rect 395 195 396 196
rect 394 195 395 196
rect 393 195 394 196
rect 344 195 345 196
rect 343 195 344 196
rect 342 195 343 196
rect 341 195 342 196
rect 340 195 341 196
rect 339 195 340 196
rect 338 195 339 196
rect 337 195 338 196
rect 336 195 337 196
rect 335 195 336 196
rect 334 195 335 196
rect 333 195 334 196
rect 332 195 333 196
rect 331 195 332 196
rect 330 195 331 196
rect 329 195 330 196
rect 328 195 329 196
rect 327 195 328 196
rect 326 195 327 196
rect 325 195 326 196
rect 324 195 325 196
rect 323 195 324 196
rect 322 195 323 196
rect 321 195 322 196
rect 320 195 321 196
rect 319 195 320 196
rect 318 195 319 196
rect 317 195 318 196
rect 316 195 317 196
rect 315 195 316 196
rect 314 195 315 196
rect 313 195 314 196
rect 312 195 313 196
rect 311 195 312 196
rect 310 195 311 196
rect 309 195 310 196
rect 308 195 309 196
rect 307 195 308 196
rect 306 195 307 196
rect 305 195 306 196
rect 304 195 305 196
rect 303 195 304 196
rect 302 195 303 196
rect 301 195 302 196
rect 300 195 301 196
rect 299 195 300 196
rect 298 195 299 196
rect 297 195 298 196
rect 296 195 297 196
rect 295 195 296 196
rect 294 195 295 196
rect 293 195 294 196
rect 292 195 293 196
rect 291 195 292 196
rect 290 195 291 196
rect 289 195 290 196
rect 288 195 289 196
rect 287 195 288 196
rect 286 195 287 196
rect 285 195 286 196
rect 284 195 285 196
rect 283 195 284 196
rect 282 195 283 196
rect 281 195 282 196
rect 280 195 281 196
rect 279 195 280 196
rect 278 195 279 196
rect 277 195 278 196
rect 276 195 277 196
rect 275 195 276 196
rect 274 195 275 196
rect 273 195 274 196
rect 272 195 273 196
rect 271 195 272 196
rect 270 195 271 196
rect 269 195 270 196
rect 268 195 269 196
rect 267 195 268 196
rect 266 195 267 196
rect 265 195 266 196
rect 264 195 265 196
rect 263 195 264 196
rect 250 195 251 196
rect 249 195 250 196
rect 248 195 249 196
rect 247 195 248 196
rect 246 195 247 196
rect 245 195 246 196
rect 244 195 245 196
rect 243 195 244 196
rect 242 195 243 196
rect 241 195 242 196
rect 240 195 241 196
rect 239 195 240 196
rect 238 195 239 196
rect 237 195 238 196
rect 236 195 237 196
rect 235 195 236 196
rect 234 195 235 196
rect 233 195 234 196
rect 232 195 233 196
rect 231 195 232 196
rect 230 195 231 196
rect 229 195 230 196
rect 228 195 229 196
rect 227 195 228 196
rect 226 195 227 196
rect 225 195 226 196
rect 224 195 225 196
rect 223 195 224 196
rect 222 195 223 196
rect 221 195 222 196
rect 220 195 221 196
rect 219 195 220 196
rect 218 195 219 196
rect 217 195 218 196
rect 216 195 217 196
rect 215 195 216 196
rect 214 195 215 196
rect 213 195 214 196
rect 212 195 213 196
rect 211 195 212 196
rect 210 195 211 196
rect 209 195 210 196
rect 183 195 184 196
rect 182 195 183 196
rect 181 195 182 196
rect 180 195 181 196
rect 179 195 180 196
rect 178 195 179 196
rect 177 195 178 196
rect 176 195 177 196
rect 175 195 176 196
rect 174 195 175 196
rect 173 195 174 196
rect 172 195 173 196
rect 171 195 172 196
rect 170 195 171 196
rect 169 195 170 196
rect 168 195 169 196
rect 167 195 168 196
rect 166 195 167 196
rect 165 195 166 196
rect 164 195 165 196
rect 163 195 164 196
rect 162 195 163 196
rect 161 195 162 196
rect 160 195 161 196
rect 159 195 160 196
rect 158 195 159 196
rect 157 195 158 196
rect 156 195 157 196
rect 155 195 156 196
rect 154 195 155 196
rect 153 195 154 196
rect 152 195 153 196
rect 151 195 152 196
rect 150 195 151 196
rect 149 195 150 196
rect 148 195 149 196
rect 147 195 148 196
rect 146 195 147 196
rect 145 195 146 196
rect 144 195 145 196
rect 143 195 144 196
rect 142 195 143 196
rect 141 195 142 196
rect 140 195 141 196
rect 139 195 140 196
rect 138 195 139 196
rect 137 195 138 196
rect 136 195 137 196
rect 135 195 136 196
rect 134 195 135 196
rect 133 195 134 196
rect 132 195 133 196
rect 131 195 132 196
rect 130 195 131 196
rect 129 195 130 196
rect 128 195 129 196
rect 127 195 128 196
rect 126 195 127 196
rect 125 195 126 196
rect 124 195 125 196
rect 123 195 124 196
rect 122 195 123 196
rect 121 195 122 196
rect 120 195 121 196
rect 119 195 120 196
rect 118 195 119 196
rect 117 195 118 196
rect 116 195 117 196
rect 115 195 116 196
rect 114 195 115 196
rect 113 195 114 196
rect 112 195 113 196
rect 111 195 112 196
rect 110 195 111 196
rect 109 195 110 196
rect 108 195 109 196
rect 107 195 108 196
rect 106 195 107 196
rect 105 195 106 196
rect 104 195 105 196
rect 103 195 104 196
rect 102 195 103 196
rect 101 195 102 196
rect 100 195 101 196
rect 99 195 100 196
rect 98 195 99 196
rect 97 195 98 196
rect 96 195 97 196
rect 95 195 96 196
rect 94 195 95 196
rect 93 195 94 196
rect 92 195 93 196
rect 91 195 92 196
rect 90 195 91 196
rect 89 195 90 196
rect 88 195 89 196
rect 87 195 88 196
rect 86 195 87 196
rect 85 195 86 196
rect 84 195 85 196
rect 83 195 84 196
rect 82 195 83 196
rect 81 195 82 196
rect 80 195 81 196
rect 79 195 80 196
rect 78 195 79 196
rect 77 195 78 196
rect 76 195 77 196
rect 75 195 76 196
rect 74 195 75 196
rect 73 195 74 196
rect 72 195 73 196
rect 71 195 72 196
rect 70 195 71 196
rect 69 195 70 196
rect 68 195 69 196
rect 50 195 51 196
rect 49 195 50 196
rect 48 195 49 196
rect 47 195 48 196
rect 46 195 47 196
rect 45 195 46 196
rect 44 195 45 196
rect 43 195 44 196
rect 42 195 43 196
rect 41 195 42 196
rect 40 195 41 196
rect 39 195 40 196
rect 38 195 39 196
rect 37 195 38 196
rect 36 195 37 196
rect 35 195 36 196
rect 34 195 35 196
rect 33 195 34 196
rect 32 195 33 196
rect 31 195 32 196
rect 30 195 31 196
rect 29 195 30 196
rect 28 195 29 196
rect 27 195 28 196
rect 26 195 27 196
rect 25 195 26 196
rect 24 195 25 196
rect 23 195 24 196
rect 22 195 23 196
rect 21 195 22 196
rect 20 195 21 196
rect 19 195 20 196
rect 18 195 19 196
rect 17 195 18 196
rect 16 195 17 196
rect 15 195 16 196
rect 14 195 15 196
rect 13 195 14 196
rect 12 195 13 196
rect 11 195 12 196
rect 10 195 11 196
rect 478 196 479 197
rect 477 196 478 197
rect 468 196 469 197
rect 467 196 468 197
rect 458 196 459 197
rect 397 196 398 197
rect 396 196 397 197
rect 395 196 396 197
rect 394 196 395 197
rect 393 196 394 197
rect 345 196 346 197
rect 344 196 345 197
rect 343 196 344 197
rect 342 196 343 197
rect 341 196 342 197
rect 340 196 341 197
rect 339 196 340 197
rect 338 196 339 197
rect 337 196 338 197
rect 336 196 337 197
rect 335 196 336 197
rect 334 196 335 197
rect 333 196 334 197
rect 332 196 333 197
rect 331 196 332 197
rect 330 196 331 197
rect 329 196 330 197
rect 328 196 329 197
rect 327 196 328 197
rect 326 196 327 197
rect 325 196 326 197
rect 324 196 325 197
rect 323 196 324 197
rect 322 196 323 197
rect 321 196 322 197
rect 320 196 321 197
rect 319 196 320 197
rect 318 196 319 197
rect 317 196 318 197
rect 316 196 317 197
rect 315 196 316 197
rect 314 196 315 197
rect 313 196 314 197
rect 312 196 313 197
rect 311 196 312 197
rect 310 196 311 197
rect 309 196 310 197
rect 308 196 309 197
rect 307 196 308 197
rect 306 196 307 197
rect 305 196 306 197
rect 304 196 305 197
rect 303 196 304 197
rect 302 196 303 197
rect 301 196 302 197
rect 300 196 301 197
rect 299 196 300 197
rect 298 196 299 197
rect 297 196 298 197
rect 296 196 297 197
rect 295 196 296 197
rect 294 196 295 197
rect 293 196 294 197
rect 292 196 293 197
rect 291 196 292 197
rect 290 196 291 197
rect 289 196 290 197
rect 288 196 289 197
rect 287 196 288 197
rect 286 196 287 197
rect 285 196 286 197
rect 284 196 285 197
rect 283 196 284 197
rect 282 196 283 197
rect 281 196 282 197
rect 280 196 281 197
rect 279 196 280 197
rect 278 196 279 197
rect 277 196 278 197
rect 276 196 277 197
rect 275 196 276 197
rect 274 196 275 197
rect 273 196 274 197
rect 272 196 273 197
rect 271 196 272 197
rect 270 196 271 197
rect 269 196 270 197
rect 268 196 269 197
rect 267 196 268 197
rect 266 196 267 197
rect 265 196 266 197
rect 264 196 265 197
rect 263 196 264 197
rect 262 196 263 197
rect 249 196 250 197
rect 248 196 249 197
rect 247 196 248 197
rect 246 196 247 197
rect 245 196 246 197
rect 244 196 245 197
rect 243 196 244 197
rect 242 196 243 197
rect 241 196 242 197
rect 240 196 241 197
rect 239 196 240 197
rect 238 196 239 197
rect 237 196 238 197
rect 236 196 237 197
rect 235 196 236 197
rect 234 196 235 197
rect 233 196 234 197
rect 232 196 233 197
rect 231 196 232 197
rect 230 196 231 197
rect 229 196 230 197
rect 228 196 229 197
rect 227 196 228 197
rect 226 196 227 197
rect 225 196 226 197
rect 224 196 225 197
rect 223 196 224 197
rect 222 196 223 197
rect 221 196 222 197
rect 220 196 221 197
rect 219 196 220 197
rect 218 196 219 197
rect 217 196 218 197
rect 216 196 217 197
rect 215 196 216 197
rect 214 196 215 197
rect 213 196 214 197
rect 212 196 213 197
rect 211 196 212 197
rect 210 196 211 197
rect 209 196 210 197
rect 208 196 209 197
rect 182 196 183 197
rect 181 196 182 197
rect 180 196 181 197
rect 179 196 180 197
rect 178 196 179 197
rect 177 196 178 197
rect 176 196 177 197
rect 175 196 176 197
rect 174 196 175 197
rect 173 196 174 197
rect 172 196 173 197
rect 171 196 172 197
rect 170 196 171 197
rect 169 196 170 197
rect 168 196 169 197
rect 167 196 168 197
rect 166 196 167 197
rect 165 196 166 197
rect 164 196 165 197
rect 163 196 164 197
rect 162 196 163 197
rect 161 196 162 197
rect 160 196 161 197
rect 159 196 160 197
rect 158 196 159 197
rect 157 196 158 197
rect 156 196 157 197
rect 155 196 156 197
rect 154 196 155 197
rect 153 196 154 197
rect 152 196 153 197
rect 151 196 152 197
rect 150 196 151 197
rect 149 196 150 197
rect 148 196 149 197
rect 147 196 148 197
rect 146 196 147 197
rect 145 196 146 197
rect 144 196 145 197
rect 143 196 144 197
rect 142 196 143 197
rect 141 196 142 197
rect 140 196 141 197
rect 139 196 140 197
rect 138 196 139 197
rect 137 196 138 197
rect 136 196 137 197
rect 135 196 136 197
rect 134 196 135 197
rect 133 196 134 197
rect 132 196 133 197
rect 131 196 132 197
rect 130 196 131 197
rect 129 196 130 197
rect 128 196 129 197
rect 127 196 128 197
rect 126 196 127 197
rect 125 196 126 197
rect 124 196 125 197
rect 123 196 124 197
rect 122 196 123 197
rect 121 196 122 197
rect 120 196 121 197
rect 119 196 120 197
rect 118 196 119 197
rect 117 196 118 197
rect 116 196 117 197
rect 115 196 116 197
rect 114 196 115 197
rect 113 196 114 197
rect 112 196 113 197
rect 111 196 112 197
rect 110 196 111 197
rect 109 196 110 197
rect 108 196 109 197
rect 107 196 108 197
rect 106 196 107 197
rect 105 196 106 197
rect 104 196 105 197
rect 103 196 104 197
rect 102 196 103 197
rect 101 196 102 197
rect 100 196 101 197
rect 99 196 100 197
rect 98 196 99 197
rect 97 196 98 197
rect 96 196 97 197
rect 95 196 96 197
rect 94 196 95 197
rect 93 196 94 197
rect 92 196 93 197
rect 91 196 92 197
rect 90 196 91 197
rect 89 196 90 197
rect 88 196 89 197
rect 87 196 88 197
rect 86 196 87 197
rect 85 196 86 197
rect 84 196 85 197
rect 83 196 84 197
rect 82 196 83 197
rect 81 196 82 197
rect 80 196 81 197
rect 79 196 80 197
rect 78 196 79 197
rect 77 196 78 197
rect 76 196 77 197
rect 75 196 76 197
rect 74 196 75 197
rect 73 196 74 197
rect 72 196 73 197
rect 71 196 72 197
rect 70 196 71 197
rect 69 196 70 197
rect 51 196 52 197
rect 50 196 51 197
rect 49 196 50 197
rect 48 196 49 197
rect 47 196 48 197
rect 46 196 47 197
rect 45 196 46 197
rect 44 196 45 197
rect 43 196 44 197
rect 42 196 43 197
rect 41 196 42 197
rect 40 196 41 197
rect 39 196 40 197
rect 38 196 39 197
rect 37 196 38 197
rect 36 196 37 197
rect 35 196 36 197
rect 34 196 35 197
rect 33 196 34 197
rect 32 196 33 197
rect 31 196 32 197
rect 30 196 31 197
rect 29 196 30 197
rect 28 196 29 197
rect 27 196 28 197
rect 26 196 27 197
rect 25 196 26 197
rect 24 196 25 197
rect 23 196 24 197
rect 22 196 23 197
rect 21 196 22 197
rect 20 196 21 197
rect 19 196 20 197
rect 18 196 19 197
rect 17 196 18 197
rect 16 196 17 197
rect 15 196 16 197
rect 14 196 15 197
rect 13 196 14 197
rect 12 196 13 197
rect 11 196 12 197
rect 10 196 11 197
rect 9 196 10 197
rect 478 197 479 198
rect 468 197 469 198
rect 467 197 468 198
rect 458 197 459 198
rect 396 197 397 198
rect 395 197 396 198
rect 394 197 395 198
rect 393 197 394 198
rect 346 197 347 198
rect 345 197 346 198
rect 344 197 345 198
rect 343 197 344 198
rect 342 197 343 198
rect 341 197 342 198
rect 340 197 341 198
rect 339 197 340 198
rect 338 197 339 198
rect 337 197 338 198
rect 336 197 337 198
rect 335 197 336 198
rect 334 197 335 198
rect 333 197 334 198
rect 332 197 333 198
rect 331 197 332 198
rect 330 197 331 198
rect 329 197 330 198
rect 328 197 329 198
rect 327 197 328 198
rect 326 197 327 198
rect 325 197 326 198
rect 324 197 325 198
rect 323 197 324 198
rect 322 197 323 198
rect 321 197 322 198
rect 320 197 321 198
rect 319 197 320 198
rect 318 197 319 198
rect 317 197 318 198
rect 316 197 317 198
rect 315 197 316 198
rect 314 197 315 198
rect 313 197 314 198
rect 312 197 313 198
rect 311 197 312 198
rect 310 197 311 198
rect 309 197 310 198
rect 308 197 309 198
rect 307 197 308 198
rect 306 197 307 198
rect 305 197 306 198
rect 304 197 305 198
rect 303 197 304 198
rect 302 197 303 198
rect 301 197 302 198
rect 300 197 301 198
rect 299 197 300 198
rect 298 197 299 198
rect 297 197 298 198
rect 296 197 297 198
rect 295 197 296 198
rect 294 197 295 198
rect 293 197 294 198
rect 292 197 293 198
rect 291 197 292 198
rect 290 197 291 198
rect 289 197 290 198
rect 288 197 289 198
rect 287 197 288 198
rect 286 197 287 198
rect 285 197 286 198
rect 284 197 285 198
rect 283 197 284 198
rect 282 197 283 198
rect 281 197 282 198
rect 280 197 281 198
rect 279 197 280 198
rect 278 197 279 198
rect 277 197 278 198
rect 276 197 277 198
rect 275 197 276 198
rect 274 197 275 198
rect 273 197 274 198
rect 272 197 273 198
rect 271 197 272 198
rect 270 197 271 198
rect 269 197 270 198
rect 268 197 269 198
rect 267 197 268 198
rect 266 197 267 198
rect 265 197 266 198
rect 264 197 265 198
rect 263 197 264 198
rect 262 197 263 198
rect 261 197 262 198
rect 248 197 249 198
rect 247 197 248 198
rect 246 197 247 198
rect 245 197 246 198
rect 244 197 245 198
rect 243 197 244 198
rect 242 197 243 198
rect 241 197 242 198
rect 240 197 241 198
rect 239 197 240 198
rect 238 197 239 198
rect 237 197 238 198
rect 236 197 237 198
rect 235 197 236 198
rect 234 197 235 198
rect 233 197 234 198
rect 232 197 233 198
rect 231 197 232 198
rect 230 197 231 198
rect 229 197 230 198
rect 228 197 229 198
rect 227 197 228 198
rect 226 197 227 198
rect 225 197 226 198
rect 224 197 225 198
rect 223 197 224 198
rect 222 197 223 198
rect 221 197 222 198
rect 220 197 221 198
rect 219 197 220 198
rect 218 197 219 198
rect 217 197 218 198
rect 216 197 217 198
rect 215 197 216 198
rect 214 197 215 198
rect 213 197 214 198
rect 212 197 213 198
rect 211 197 212 198
rect 210 197 211 198
rect 209 197 210 198
rect 208 197 209 198
rect 181 197 182 198
rect 180 197 181 198
rect 179 197 180 198
rect 178 197 179 198
rect 177 197 178 198
rect 176 197 177 198
rect 175 197 176 198
rect 174 197 175 198
rect 173 197 174 198
rect 172 197 173 198
rect 171 197 172 198
rect 170 197 171 198
rect 169 197 170 198
rect 168 197 169 198
rect 167 197 168 198
rect 166 197 167 198
rect 165 197 166 198
rect 164 197 165 198
rect 163 197 164 198
rect 162 197 163 198
rect 161 197 162 198
rect 160 197 161 198
rect 159 197 160 198
rect 158 197 159 198
rect 157 197 158 198
rect 156 197 157 198
rect 155 197 156 198
rect 154 197 155 198
rect 153 197 154 198
rect 152 197 153 198
rect 151 197 152 198
rect 150 197 151 198
rect 149 197 150 198
rect 148 197 149 198
rect 147 197 148 198
rect 146 197 147 198
rect 145 197 146 198
rect 144 197 145 198
rect 143 197 144 198
rect 142 197 143 198
rect 141 197 142 198
rect 140 197 141 198
rect 139 197 140 198
rect 138 197 139 198
rect 137 197 138 198
rect 136 197 137 198
rect 135 197 136 198
rect 134 197 135 198
rect 133 197 134 198
rect 132 197 133 198
rect 131 197 132 198
rect 130 197 131 198
rect 129 197 130 198
rect 128 197 129 198
rect 127 197 128 198
rect 126 197 127 198
rect 125 197 126 198
rect 124 197 125 198
rect 123 197 124 198
rect 122 197 123 198
rect 121 197 122 198
rect 120 197 121 198
rect 119 197 120 198
rect 118 197 119 198
rect 117 197 118 198
rect 116 197 117 198
rect 115 197 116 198
rect 114 197 115 198
rect 113 197 114 198
rect 112 197 113 198
rect 111 197 112 198
rect 110 197 111 198
rect 109 197 110 198
rect 108 197 109 198
rect 107 197 108 198
rect 106 197 107 198
rect 105 197 106 198
rect 104 197 105 198
rect 103 197 104 198
rect 102 197 103 198
rect 101 197 102 198
rect 100 197 101 198
rect 99 197 100 198
rect 98 197 99 198
rect 97 197 98 198
rect 96 197 97 198
rect 95 197 96 198
rect 94 197 95 198
rect 93 197 94 198
rect 92 197 93 198
rect 91 197 92 198
rect 90 197 91 198
rect 89 197 90 198
rect 88 197 89 198
rect 87 197 88 198
rect 86 197 87 198
rect 85 197 86 198
rect 84 197 85 198
rect 83 197 84 198
rect 82 197 83 198
rect 81 197 82 198
rect 80 197 81 198
rect 79 197 80 198
rect 78 197 79 198
rect 77 197 78 198
rect 76 197 77 198
rect 75 197 76 198
rect 74 197 75 198
rect 73 197 74 198
rect 72 197 73 198
rect 71 197 72 198
rect 70 197 71 198
rect 69 197 70 198
rect 52 197 53 198
rect 51 197 52 198
rect 50 197 51 198
rect 49 197 50 198
rect 48 197 49 198
rect 47 197 48 198
rect 46 197 47 198
rect 45 197 46 198
rect 44 197 45 198
rect 43 197 44 198
rect 42 197 43 198
rect 41 197 42 198
rect 40 197 41 198
rect 39 197 40 198
rect 38 197 39 198
rect 37 197 38 198
rect 36 197 37 198
rect 35 197 36 198
rect 34 197 35 198
rect 33 197 34 198
rect 32 197 33 198
rect 31 197 32 198
rect 30 197 31 198
rect 29 197 30 198
rect 28 197 29 198
rect 27 197 28 198
rect 26 197 27 198
rect 25 197 26 198
rect 24 197 25 198
rect 23 197 24 198
rect 22 197 23 198
rect 21 197 22 198
rect 20 197 21 198
rect 19 197 20 198
rect 18 197 19 198
rect 17 197 18 198
rect 16 197 17 198
rect 15 197 16 198
rect 14 197 15 198
rect 13 197 14 198
rect 12 197 13 198
rect 11 197 12 198
rect 10 197 11 198
rect 9 197 10 198
rect 478 198 479 199
rect 468 198 469 199
rect 467 198 468 199
rect 458 198 459 199
rect 395 198 396 199
rect 394 198 395 199
rect 393 198 394 199
rect 347 198 348 199
rect 346 198 347 199
rect 345 198 346 199
rect 344 198 345 199
rect 343 198 344 199
rect 342 198 343 199
rect 341 198 342 199
rect 340 198 341 199
rect 339 198 340 199
rect 338 198 339 199
rect 337 198 338 199
rect 336 198 337 199
rect 335 198 336 199
rect 334 198 335 199
rect 333 198 334 199
rect 332 198 333 199
rect 331 198 332 199
rect 330 198 331 199
rect 329 198 330 199
rect 328 198 329 199
rect 327 198 328 199
rect 326 198 327 199
rect 325 198 326 199
rect 324 198 325 199
rect 323 198 324 199
rect 322 198 323 199
rect 321 198 322 199
rect 320 198 321 199
rect 319 198 320 199
rect 318 198 319 199
rect 317 198 318 199
rect 316 198 317 199
rect 315 198 316 199
rect 314 198 315 199
rect 313 198 314 199
rect 312 198 313 199
rect 311 198 312 199
rect 310 198 311 199
rect 309 198 310 199
rect 308 198 309 199
rect 307 198 308 199
rect 306 198 307 199
rect 305 198 306 199
rect 304 198 305 199
rect 303 198 304 199
rect 302 198 303 199
rect 301 198 302 199
rect 300 198 301 199
rect 299 198 300 199
rect 298 198 299 199
rect 297 198 298 199
rect 296 198 297 199
rect 295 198 296 199
rect 294 198 295 199
rect 293 198 294 199
rect 292 198 293 199
rect 291 198 292 199
rect 290 198 291 199
rect 289 198 290 199
rect 288 198 289 199
rect 287 198 288 199
rect 286 198 287 199
rect 285 198 286 199
rect 284 198 285 199
rect 283 198 284 199
rect 282 198 283 199
rect 281 198 282 199
rect 280 198 281 199
rect 279 198 280 199
rect 278 198 279 199
rect 277 198 278 199
rect 276 198 277 199
rect 275 198 276 199
rect 274 198 275 199
rect 273 198 274 199
rect 272 198 273 199
rect 271 198 272 199
rect 270 198 271 199
rect 269 198 270 199
rect 268 198 269 199
rect 267 198 268 199
rect 266 198 267 199
rect 265 198 266 199
rect 264 198 265 199
rect 263 198 264 199
rect 262 198 263 199
rect 261 198 262 199
rect 260 198 261 199
rect 259 198 260 199
rect 248 198 249 199
rect 247 198 248 199
rect 246 198 247 199
rect 245 198 246 199
rect 244 198 245 199
rect 243 198 244 199
rect 242 198 243 199
rect 241 198 242 199
rect 240 198 241 199
rect 239 198 240 199
rect 238 198 239 199
rect 237 198 238 199
rect 236 198 237 199
rect 235 198 236 199
rect 234 198 235 199
rect 233 198 234 199
rect 232 198 233 199
rect 231 198 232 199
rect 230 198 231 199
rect 229 198 230 199
rect 228 198 229 199
rect 227 198 228 199
rect 226 198 227 199
rect 225 198 226 199
rect 224 198 225 199
rect 223 198 224 199
rect 222 198 223 199
rect 221 198 222 199
rect 220 198 221 199
rect 219 198 220 199
rect 218 198 219 199
rect 217 198 218 199
rect 216 198 217 199
rect 215 198 216 199
rect 214 198 215 199
rect 213 198 214 199
rect 212 198 213 199
rect 211 198 212 199
rect 210 198 211 199
rect 209 198 210 199
rect 208 198 209 199
rect 207 198 208 199
rect 180 198 181 199
rect 179 198 180 199
rect 178 198 179 199
rect 177 198 178 199
rect 176 198 177 199
rect 175 198 176 199
rect 174 198 175 199
rect 173 198 174 199
rect 172 198 173 199
rect 171 198 172 199
rect 170 198 171 199
rect 169 198 170 199
rect 168 198 169 199
rect 167 198 168 199
rect 166 198 167 199
rect 165 198 166 199
rect 164 198 165 199
rect 163 198 164 199
rect 162 198 163 199
rect 161 198 162 199
rect 160 198 161 199
rect 159 198 160 199
rect 158 198 159 199
rect 157 198 158 199
rect 156 198 157 199
rect 155 198 156 199
rect 154 198 155 199
rect 153 198 154 199
rect 152 198 153 199
rect 151 198 152 199
rect 150 198 151 199
rect 149 198 150 199
rect 148 198 149 199
rect 147 198 148 199
rect 146 198 147 199
rect 145 198 146 199
rect 144 198 145 199
rect 143 198 144 199
rect 142 198 143 199
rect 141 198 142 199
rect 140 198 141 199
rect 139 198 140 199
rect 138 198 139 199
rect 137 198 138 199
rect 136 198 137 199
rect 135 198 136 199
rect 134 198 135 199
rect 133 198 134 199
rect 132 198 133 199
rect 131 198 132 199
rect 130 198 131 199
rect 129 198 130 199
rect 128 198 129 199
rect 127 198 128 199
rect 126 198 127 199
rect 125 198 126 199
rect 124 198 125 199
rect 123 198 124 199
rect 122 198 123 199
rect 121 198 122 199
rect 120 198 121 199
rect 119 198 120 199
rect 118 198 119 199
rect 117 198 118 199
rect 116 198 117 199
rect 115 198 116 199
rect 114 198 115 199
rect 113 198 114 199
rect 112 198 113 199
rect 111 198 112 199
rect 110 198 111 199
rect 109 198 110 199
rect 108 198 109 199
rect 107 198 108 199
rect 106 198 107 199
rect 105 198 106 199
rect 104 198 105 199
rect 103 198 104 199
rect 102 198 103 199
rect 101 198 102 199
rect 100 198 101 199
rect 99 198 100 199
rect 98 198 99 199
rect 97 198 98 199
rect 96 198 97 199
rect 95 198 96 199
rect 94 198 95 199
rect 93 198 94 199
rect 92 198 93 199
rect 91 198 92 199
rect 90 198 91 199
rect 89 198 90 199
rect 88 198 89 199
rect 87 198 88 199
rect 86 198 87 199
rect 85 198 86 199
rect 84 198 85 199
rect 83 198 84 199
rect 82 198 83 199
rect 81 198 82 199
rect 80 198 81 199
rect 79 198 80 199
rect 78 198 79 199
rect 77 198 78 199
rect 76 198 77 199
rect 75 198 76 199
rect 74 198 75 199
rect 73 198 74 199
rect 72 198 73 199
rect 71 198 72 199
rect 70 198 71 199
rect 69 198 70 199
rect 52 198 53 199
rect 51 198 52 199
rect 50 198 51 199
rect 49 198 50 199
rect 48 198 49 199
rect 47 198 48 199
rect 46 198 47 199
rect 45 198 46 199
rect 44 198 45 199
rect 43 198 44 199
rect 42 198 43 199
rect 41 198 42 199
rect 40 198 41 199
rect 39 198 40 199
rect 38 198 39 199
rect 37 198 38 199
rect 36 198 37 199
rect 35 198 36 199
rect 34 198 35 199
rect 33 198 34 199
rect 32 198 33 199
rect 31 198 32 199
rect 30 198 31 199
rect 29 198 30 199
rect 28 198 29 199
rect 27 198 28 199
rect 26 198 27 199
rect 25 198 26 199
rect 24 198 25 199
rect 23 198 24 199
rect 22 198 23 199
rect 21 198 22 199
rect 20 198 21 199
rect 19 198 20 199
rect 18 198 19 199
rect 17 198 18 199
rect 16 198 17 199
rect 15 198 16 199
rect 14 198 15 199
rect 13 198 14 199
rect 12 198 13 199
rect 11 198 12 199
rect 10 198 11 199
rect 9 198 10 199
rect 478 199 479 200
rect 468 199 469 200
rect 467 199 468 200
rect 458 199 459 200
rect 395 199 396 200
rect 394 199 395 200
rect 393 199 394 200
rect 348 199 349 200
rect 347 199 348 200
rect 346 199 347 200
rect 345 199 346 200
rect 344 199 345 200
rect 343 199 344 200
rect 342 199 343 200
rect 341 199 342 200
rect 340 199 341 200
rect 339 199 340 200
rect 338 199 339 200
rect 337 199 338 200
rect 336 199 337 200
rect 335 199 336 200
rect 334 199 335 200
rect 333 199 334 200
rect 332 199 333 200
rect 331 199 332 200
rect 330 199 331 200
rect 329 199 330 200
rect 328 199 329 200
rect 327 199 328 200
rect 326 199 327 200
rect 325 199 326 200
rect 324 199 325 200
rect 323 199 324 200
rect 322 199 323 200
rect 321 199 322 200
rect 320 199 321 200
rect 319 199 320 200
rect 318 199 319 200
rect 317 199 318 200
rect 316 199 317 200
rect 315 199 316 200
rect 314 199 315 200
rect 313 199 314 200
rect 312 199 313 200
rect 311 199 312 200
rect 310 199 311 200
rect 309 199 310 200
rect 308 199 309 200
rect 307 199 308 200
rect 306 199 307 200
rect 305 199 306 200
rect 304 199 305 200
rect 303 199 304 200
rect 302 199 303 200
rect 301 199 302 200
rect 300 199 301 200
rect 299 199 300 200
rect 298 199 299 200
rect 297 199 298 200
rect 296 199 297 200
rect 295 199 296 200
rect 294 199 295 200
rect 293 199 294 200
rect 292 199 293 200
rect 291 199 292 200
rect 290 199 291 200
rect 289 199 290 200
rect 288 199 289 200
rect 287 199 288 200
rect 286 199 287 200
rect 285 199 286 200
rect 284 199 285 200
rect 283 199 284 200
rect 282 199 283 200
rect 281 199 282 200
rect 280 199 281 200
rect 279 199 280 200
rect 278 199 279 200
rect 277 199 278 200
rect 276 199 277 200
rect 275 199 276 200
rect 274 199 275 200
rect 273 199 274 200
rect 272 199 273 200
rect 271 199 272 200
rect 270 199 271 200
rect 269 199 270 200
rect 268 199 269 200
rect 267 199 268 200
rect 266 199 267 200
rect 265 199 266 200
rect 264 199 265 200
rect 263 199 264 200
rect 262 199 263 200
rect 261 199 262 200
rect 260 199 261 200
rect 259 199 260 200
rect 258 199 259 200
rect 247 199 248 200
rect 246 199 247 200
rect 245 199 246 200
rect 244 199 245 200
rect 243 199 244 200
rect 242 199 243 200
rect 241 199 242 200
rect 240 199 241 200
rect 239 199 240 200
rect 238 199 239 200
rect 237 199 238 200
rect 236 199 237 200
rect 235 199 236 200
rect 234 199 235 200
rect 233 199 234 200
rect 232 199 233 200
rect 231 199 232 200
rect 230 199 231 200
rect 229 199 230 200
rect 228 199 229 200
rect 227 199 228 200
rect 226 199 227 200
rect 225 199 226 200
rect 224 199 225 200
rect 223 199 224 200
rect 222 199 223 200
rect 221 199 222 200
rect 220 199 221 200
rect 219 199 220 200
rect 218 199 219 200
rect 217 199 218 200
rect 216 199 217 200
rect 215 199 216 200
rect 214 199 215 200
rect 213 199 214 200
rect 212 199 213 200
rect 211 199 212 200
rect 210 199 211 200
rect 209 199 210 200
rect 208 199 209 200
rect 207 199 208 200
rect 206 199 207 200
rect 178 199 179 200
rect 177 199 178 200
rect 176 199 177 200
rect 175 199 176 200
rect 174 199 175 200
rect 173 199 174 200
rect 172 199 173 200
rect 171 199 172 200
rect 170 199 171 200
rect 169 199 170 200
rect 168 199 169 200
rect 167 199 168 200
rect 166 199 167 200
rect 165 199 166 200
rect 164 199 165 200
rect 163 199 164 200
rect 162 199 163 200
rect 161 199 162 200
rect 160 199 161 200
rect 159 199 160 200
rect 158 199 159 200
rect 157 199 158 200
rect 156 199 157 200
rect 155 199 156 200
rect 154 199 155 200
rect 153 199 154 200
rect 152 199 153 200
rect 151 199 152 200
rect 150 199 151 200
rect 149 199 150 200
rect 148 199 149 200
rect 147 199 148 200
rect 146 199 147 200
rect 145 199 146 200
rect 144 199 145 200
rect 143 199 144 200
rect 142 199 143 200
rect 141 199 142 200
rect 140 199 141 200
rect 139 199 140 200
rect 138 199 139 200
rect 137 199 138 200
rect 136 199 137 200
rect 135 199 136 200
rect 134 199 135 200
rect 133 199 134 200
rect 132 199 133 200
rect 131 199 132 200
rect 130 199 131 200
rect 129 199 130 200
rect 128 199 129 200
rect 127 199 128 200
rect 126 199 127 200
rect 125 199 126 200
rect 124 199 125 200
rect 123 199 124 200
rect 122 199 123 200
rect 121 199 122 200
rect 120 199 121 200
rect 119 199 120 200
rect 118 199 119 200
rect 117 199 118 200
rect 116 199 117 200
rect 115 199 116 200
rect 114 199 115 200
rect 113 199 114 200
rect 112 199 113 200
rect 111 199 112 200
rect 110 199 111 200
rect 109 199 110 200
rect 108 199 109 200
rect 107 199 108 200
rect 106 199 107 200
rect 105 199 106 200
rect 104 199 105 200
rect 103 199 104 200
rect 102 199 103 200
rect 101 199 102 200
rect 100 199 101 200
rect 99 199 100 200
rect 98 199 99 200
rect 97 199 98 200
rect 96 199 97 200
rect 95 199 96 200
rect 94 199 95 200
rect 93 199 94 200
rect 92 199 93 200
rect 91 199 92 200
rect 90 199 91 200
rect 89 199 90 200
rect 88 199 89 200
rect 87 199 88 200
rect 86 199 87 200
rect 85 199 86 200
rect 84 199 85 200
rect 83 199 84 200
rect 82 199 83 200
rect 81 199 82 200
rect 80 199 81 200
rect 79 199 80 200
rect 78 199 79 200
rect 77 199 78 200
rect 76 199 77 200
rect 75 199 76 200
rect 74 199 75 200
rect 73 199 74 200
rect 72 199 73 200
rect 71 199 72 200
rect 70 199 71 200
rect 53 199 54 200
rect 52 199 53 200
rect 51 199 52 200
rect 50 199 51 200
rect 49 199 50 200
rect 48 199 49 200
rect 47 199 48 200
rect 46 199 47 200
rect 45 199 46 200
rect 44 199 45 200
rect 43 199 44 200
rect 42 199 43 200
rect 41 199 42 200
rect 40 199 41 200
rect 39 199 40 200
rect 38 199 39 200
rect 37 199 38 200
rect 36 199 37 200
rect 35 199 36 200
rect 34 199 35 200
rect 33 199 34 200
rect 32 199 33 200
rect 31 199 32 200
rect 30 199 31 200
rect 29 199 30 200
rect 28 199 29 200
rect 27 199 28 200
rect 26 199 27 200
rect 25 199 26 200
rect 24 199 25 200
rect 23 199 24 200
rect 22 199 23 200
rect 21 199 22 200
rect 20 199 21 200
rect 19 199 20 200
rect 18 199 19 200
rect 17 199 18 200
rect 16 199 17 200
rect 15 199 16 200
rect 14 199 15 200
rect 13 199 14 200
rect 12 199 13 200
rect 11 199 12 200
rect 10 199 11 200
rect 9 199 10 200
rect 478 200 479 201
rect 468 200 469 201
rect 467 200 468 201
rect 458 200 459 201
rect 395 200 396 201
rect 394 200 395 201
rect 393 200 394 201
rect 348 200 349 201
rect 347 200 348 201
rect 346 200 347 201
rect 345 200 346 201
rect 344 200 345 201
rect 343 200 344 201
rect 342 200 343 201
rect 341 200 342 201
rect 340 200 341 201
rect 339 200 340 201
rect 338 200 339 201
rect 337 200 338 201
rect 336 200 337 201
rect 335 200 336 201
rect 334 200 335 201
rect 333 200 334 201
rect 332 200 333 201
rect 331 200 332 201
rect 330 200 331 201
rect 329 200 330 201
rect 328 200 329 201
rect 327 200 328 201
rect 326 200 327 201
rect 325 200 326 201
rect 324 200 325 201
rect 323 200 324 201
rect 322 200 323 201
rect 321 200 322 201
rect 320 200 321 201
rect 319 200 320 201
rect 318 200 319 201
rect 317 200 318 201
rect 316 200 317 201
rect 315 200 316 201
rect 314 200 315 201
rect 313 200 314 201
rect 312 200 313 201
rect 311 200 312 201
rect 310 200 311 201
rect 309 200 310 201
rect 308 200 309 201
rect 307 200 308 201
rect 306 200 307 201
rect 305 200 306 201
rect 304 200 305 201
rect 303 200 304 201
rect 302 200 303 201
rect 301 200 302 201
rect 300 200 301 201
rect 299 200 300 201
rect 298 200 299 201
rect 297 200 298 201
rect 296 200 297 201
rect 295 200 296 201
rect 294 200 295 201
rect 293 200 294 201
rect 292 200 293 201
rect 291 200 292 201
rect 290 200 291 201
rect 289 200 290 201
rect 288 200 289 201
rect 287 200 288 201
rect 286 200 287 201
rect 285 200 286 201
rect 284 200 285 201
rect 283 200 284 201
rect 282 200 283 201
rect 281 200 282 201
rect 280 200 281 201
rect 279 200 280 201
rect 278 200 279 201
rect 277 200 278 201
rect 276 200 277 201
rect 275 200 276 201
rect 274 200 275 201
rect 273 200 274 201
rect 272 200 273 201
rect 271 200 272 201
rect 270 200 271 201
rect 269 200 270 201
rect 268 200 269 201
rect 267 200 268 201
rect 266 200 267 201
rect 265 200 266 201
rect 264 200 265 201
rect 263 200 264 201
rect 262 200 263 201
rect 261 200 262 201
rect 260 200 261 201
rect 259 200 260 201
rect 258 200 259 201
rect 257 200 258 201
rect 256 200 257 201
rect 247 200 248 201
rect 246 200 247 201
rect 245 200 246 201
rect 244 200 245 201
rect 243 200 244 201
rect 242 200 243 201
rect 241 200 242 201
rect 240 200 241 201
rect 239 200 240 201
rect 238 200 239 201
rect 237 200 238 201
rect 236 200 237 201
rect 235 200 236 201
rect 234 200 235 201
rect 233 200 234 201
rect 232 200 233 201
rect 231 200 232 201
rect 230 200 231 201
rect 229 200 230 201
rect 228 200 229 201
rect 227 200 228 201
rect 226 200 227 201
rect 225 200 226 201
rect 224 200 225 201
rect 223 200 224 201
rect 222 200 223 201
rect 221 200 222 201
rect 220 200 221 201
rect 219 200 220 201
rect 218 200 219 201
rect 217 200 218 201
rect 216 200 217 201
rect 215 200 216 201
rect 214 200 215 201
rect 213 200 214 201
rect 212 200 213 201
rect 211 200 212 201
rect 210 200 211 201
rect 209 200 210 201
rect 208 200 209 201
rect 207 200 208 201
rect 206 200 207 201
rect 205 200 206 201
rect 177 200 178 201
rect 176 200 177 201
rect 175 200 176 201
rect 174 200 175 201
rect 173 200 174 201
rect 172 200 173 201
rect 171 200 172 201
rect 170 200 171 201
rect 169 200 170 201
rect 168 200 169 201
rect 167 200 168 201
rect 166 200 167 201
rect 165 200 166 201
rect 164 200 165 201
rect 163 200 164 201
rect 162 200 163 201
rect 161 200 162 201
rect 160 200 161 201
rect 159 200 160 201
rect 158 200 159 201
rect 157 200 158 201
rect 156 200 157 201
rect 155 200 156 201
rect 154 200 155 201
rect 153 200 154 201
rect 152 200 153 201
rect 151 200 152 201
rect 150 200 151 201
rect 149 200 150 201
rect 148 200 149 201
rect 147 200 148 201
rect 146 200 147 201
rect 145 200 146 201
rect 144 200 145 201
rect 143 200 144 201
rect 142 200 143 201
rect 141 200 142 201
rect 140 200 141 201
rect 139 200 140 201
rect 138 200 139 201
rect 137 200 138 201
rect 136 200 137 201
rect 135 200 136 201
rect 134 200 135 201
rect 133 200 134 201
rect 132 200 133 201
rect 131 200 132 201
rect 130 200 131 201
rect 129 200 130 201
rect 128 200 129 201
rect 127 200 128 201
rect 126 200 127 201
rect 125 200 126 201
rect 124 200 125 201
rect 123 200 124 201
rect 122 200 123 201
rect 121 200 122 201
rect 120 200 121 201
rect 119 200 120 201
rect 118 200 119 201
rect 117 200 118 201
rect 116 200 117 201
rect 115 200 116 201
rect 114 200 115 201
rect 113 200 114 201
rect 112 200 113 201
rect 111 200 112 201
rect 110 200 111 201
rect 109 200 110 201
rect 108 200 109 201
rect 107 200 108 201
rect 106 200 107 201
rect 105 200 106 201
rect 104 200 105 201
rect 103 200 104 201
rect 102 200 103 201
rect 101 200 102 201
rect 100 200 101 201
rect 99 200 100 201
rect 98 200 99 201
rect 97 200 98 201
rect 96 200 97 201
rect 95 200 96 201
rect 94 200 95 201
rect 93 200 94 201
rect 92 200 93 201
rect 91 200 92 201
rect 90 200 91 201
rect 89 200 90 201
rect 88 200 89 201
rect 87 200 88 201
rect 86 200 87 201
rect 85 200 86 201
rect 84 200 85 201
rect 83 200 84 201
rect 82 200 83 201
rect 81 200 82 201
rect 80 200 81 201
rect 79 200 80 201
rect 78 200 79 201
rect 77 200 78 201
rect 76 200 77 201
rect 75 200 76 201
rect 74 200 75 201
rect 73 200 74 201
rect 72 200 73 201
rect 71 200 72 201
rect 54 200 55 201
rect 53 200 54 201
rect 52 200 53 201
rect 51 200 52 201
rect 50 200 51 201
rect 49 200 50 201
rect 48 200 49 201
rect 47 200 48 201
rect 46 200 47 201
rect 45 200 46 201
rect 44 200 45 201
rect 43 200 44 201
rect 42 200 43 201
rect 41 200 42 201
rect 40 200 41 201
rect 39 200 40 201
rect 38 200 39 201
rect 37 200 38 201
rect 36 200 37 201
rect 35 200 36 201
rect 34 200 35 201
rect 33 200 34 201
rect 32 200 33 201
rect 31 200 32 201
rect 30 200 31 201
rect 29 200 30 201
rect 28 200 29 201
rect 27 200 28 201
rect 26 200 27 201
rect 25 200 26 201
rect 24 200 25 201
rect 23 200 24 201
rect 22 200 23 201
rect 21 200 22 201
rect 20 200 21 201
rect 19 200 20 201
rect 18 200 19 201
rect 17 200 18 201
rect 16 200 17 201
rect 15 200 16 201
rect 14 200 15 201
rect 13 200 14 201
rect 12 200 13 201
rect 11 200 12 201
rect 10 200 11 201
rect 9 200 10 201
rect 478 201 479 202
rect 470 201 471 202
rect 469 201 470 202
rect 468 201 469 202
rect 467 201 468 202
rect 466 201 467 202
rect 465 201 466 202
rect 459 201 460 202
rect 458 201 459 202
rect 394 201 395 202
rect 349 201 350 202
rect 348 201 349 202
rect 347 201 348 202
rect 346 201 347 202
rect 345 201 346 202
rect 344 201 345 202
rect 343 201 344 202
rect 342 201 343 202
rect 341 201 342 202
rect 340 201 341 202
rect 339 201 340 202
rect 338 201 339 202
rect 337 201 338 202
rect 336 201 337 202
rect 335 201 336 202
rect 334 201 335 202
rect 333 201 334 202
rect 332 201 333 202
rect 331 201 332 202
rect 330 201 331 202
rect 329 201 330 202
rect 328 201 329 202
rect 327 201 328 202
rect 326 201 327 202
rect 325 201 326 202
rect 324 201 325 202
rect 323 201 324 202
rect 322 201 323 202
rect 321 201 322 202
rect 320 201 321 202
rect 319 201 320 202
rect 318 201 319 202
rect 317 201 318 202
rect 316 201 317 202
rect 315 201 316 202
rect 314 201 315 202
rect 313 201 314 202
rect 312 201 313 202
rect 311 201 312 202
rect 310 201 311 202
rect 309 201 310 202
rect 308 201 309 202
rect 307 201 308 202
rect 306 201 307 202
rect 305 201 306 202
rect 304 201 305 202
rect 303 201 304 202
rect 302 201 303 202
rect 301 201 302 202
rect 300 201 301 202
rect 299 201 300 202
rect 298 201 299 202
rect 297 201 298 202
rect 296 201 297 202
rect 295 201 296 202
rect 294 201 295 202
rect 293 201 294 202
rect 292 201 293 202
rect 291 201 292 202
rect 290 201 291 202
rect 289 201 290 202
rect 288 201 289 202
rect 287 201 288 202
rect 286 201 287 202
rect 285 201 286 202
rect 284 201 285 202
rect 283 201 284 202
rect 282 201 283 202
rect 281 201 282 202
rect 280 201 281 202
rect 279 201 280 202
rect 278 201 279 202
rect 277 201 278 202
rect 276 201 277 202
rect 275 201 276 202
rect 274 201 275 202
rect 273 201 274 202
rect 272 201 273 202
rect 271 201 272 202
rect 270 201 271 202
rect 269 201 270 202
rect 268 201 269 202
rect 267 201 268 202
rect 266 201 267 202
rect 265 201 266 202
rect 264 201 265 202
rect 263 201 264 202
rect 262 201 263 202
rect 261 201 262 202
rect 260 201 261 202
rect 259 201 260 202
rect 258 201 259 202
rect 257 201 258 202
rect 256 201 257 202
rect 255 201 256 202
rect 246 201 247 202
rect 245 201 246 202
rect 244 201 245 202
rect 243 201 244 202
rect 242 201 243 202
rect 241 201 242 202
rect 240 201 241 202
rect 239 201 240 202
rect 238 201 239 202
rect 237 201 238 202
rect 236 201 237 202
rect 235 201 236 202
rect 234 201 235 202
rect 233 201 234 202
rect 232 201 233 202
rect 231 201 232 202
rect 230 201 231 202
rect 229 201 230 202
rect 228 201 229 202
rect 227 201 228 202
rect 226 201 227 202
rect 225 201 226 202
rect 224 201 225 202
rect 223 201 224 202
rect 222 201 223 202
rect 221 201 222 202
rect 220 201 221 202
rect 219 201 220 202
rect 218 201 219 202
rect 217 201 218 202
rect 216 201 217 202
rect 215 201 216 202
rect 214 201 215 202
rect 213 201 214 202
rect 212 201 213 202
rect 211 201 212 202
rect 210 201 211 202
rect 209 201 210 202
rect 208 201 209 202
rect 207 201 208 202
rect 206 201 207 202
rect 205 201 206 202
rect 204 201 205 202
rect 175 201 176 202
rect 174 201 175 202
rect 173 201 174 202
rect 172 201 173 202
rect 171 201 172 202
rect 170 201 171 202
rect 169 201 170 202
rect 168 201 169 202
rect 167 201 168 202
rect 166 201 167 202
rect 165 201 166 202
rect 164 201 165 202
rect 163 201 164 202
rect 162 201 163 202
rect 161 201 162 202
rect 160 201 161 202
rect 159 201 160 202
rect 158 201 159 202
rect 157 201 158 202
rect 156 201 157 202
rect 155 201 156 202
rect 154 201 155 202
rect 153 201 154 202
rect 152 201 153 202
rect 151 201 152 202
rect 150 201 151 202
rect 149 201 150 202
rect 148 201 149 202
rect 147 201 148 202
rect 146 201 147 202
rect 145 201 146 202
rect 144 201 145 202
rect 143 201 144 202
rect 142 201 143 202
rect 141 201 142 202
rect 140 201 141 202
rect 139 201 140 202
rect 138 201 139 202
rect 137 201 138 202
rect 136 201 137 202
rect 135 201 136 202
rect 134 201 135 202
rect 133 201 134 202
rect 132 201 133 202
rect 131 201 132 202
rect 130 201 131 202
rect 129 201 130 202
rect 128 201 129 202
rect 127 201 128 202
rect 126 201 127 202
rect 125 201 126 202
rect 124 201 125 202
rect 123 201 124 202
rect 122 201 123 202
rect 121 201 122 202
rect 120 201 121 202
rect 119 201 120 202
rect 118 201 119 202
rect 117 201 118 202
rect 116 201 117 202
rect 115 201 116 202
rect 114 201 115 202
rect 113 201 114 202
rect 112 201 113 202
rect 111 201 112 202
rect 110 201 111 202
rect 109 201 110 202
rect 108 201 109 202
rect 107 201 108 202
rect 106 201 107 202
rect 105 201 106 202
rect 104 201 105 202
rect 103 201 104 202
rect 102 201 103 202
rect 101 201 102 202
rect 100 201 101 202
rect 99 201 100 202
rect 98 201 99 202
rect 97 201 98 202
rect 96 201 97 202
rect 95 201 96 202
rect 94 201 95 202
rect 93 201 94 202
rect 92 201 93 202
rect 91 201 92 202
rect 90 201 91 202
rect 89 201 90 202
rect 88 201 89 202
rect 87 201 88 202
rect 86 201 87 202
rect 85 201 86 202
rect 84 201 85 202
rect 83 201 84 202
rect 82 201 83 202
rect 81 201 82 202
rect 80 201 81 202
rect 79 201 80 202
rect 78 201 79 202
rect 77 201 78 202
rect 76 201 77 202
rect 75 201 76 202
rect 74 201 75 202
rect 73 201 74 202
rect 72 201 73 202
rect 71 201 72 202
rect 54 201 55 202
rect 53 201 54 202
rect 52 201 53 202
rect 51 201 52 202
rect 50 201 51 202
rect 49 201 50 202
rect 48 201 49 202
rect 47 201 48 202
rect 46 201 47 202
rect 45 201 46 202
rect 44 201 45 202
rect 43 201 44 202
rect 42 201 43 202
rect 41 201 42 202
rect 40 201 41 202
rect 39 201 40 202
rect 38 201 39 202
rect 37 201 38 202
rect 36 201 37 202
rect 35 201 36 202
rect 34 201 35 202
rect 33 201 34 202
rect 32 201 33 202
rect 31 201 32 202
rect 30 201 31 202
rect 29 201 30 202
rect 28 201 29 202
rect 27 201 28 202
rect 26 201 27 202
rect 25 201 26 202
rect 24 201 25 202
rect 23 201 24 202
rect 22 201 23 202
rect 21 201 22 202
rect 20 201 21 202
rect 19 201 20 202
rect 18 201 19 202
rect 17 201 18 202
rect 16 201 17 202
rect 15 201 16 202
rect 14 201 15 202
rect 13 201 14 202
rect 12 201 13 202
rect 11 201 12 202
rect 10 201 11 202
rect 9 201 10 202
rect 478 202 479 203
rect 477 202 478 203
rect 471 202 472 203
rect 470 202 471 203
rect 469 202 470 203
rect 468 202 469 203
rect 467 202 468 203
rect 466 202 467 203
rect 465 202 466 203
rect 460 202 461 203
rect 459 202 460 203
rect 458 202 459 203
rect 350 202 351 203
rect 349 202 350 203
rect 348 202 349 203
rect 347 202 348 203
rect 346 202 347 203
rect 345 202 346 203
rect 344 202 345 203
rect 343 202 344 203
rect 342 202 343 203
rect 341 202 342 203
rect 340 202 341 203
rect 339 202 340 203
rect 338 202 339 203
rect 337 202 338 203
rect 336 202 337 203
rect 335 202 336 203
rect 334 202 335 203
rect 333 202 334 203
rect 332 202 333 203
rect 331 202 332 203
rect 330 202 331 203
rect 329 202 330 203
rect 328 202 329 203
rect 327 202 328 203
rect 326 202 327 203
rect 325 202 326 203
rect 324 202 325 203
rect 323 202 324 203
rect 322 202 323 203
rect 321 202 322 203
rect 320 202 321 203
rect 319 202 320 203
rect 318 202 319 203
rect 317 202 318 203
rect 316 202 317 203
rect 315 202 316 203
rect 314 202 315 203
rect 313 202 314 203
rect 312 202 313 203
rect 311 202 312 203
rect 310 202 311 203
rect 309 202 310 203
rect 308 202 309 203
rect 307 202 308 203
rect 306 202 307 203
rect 305 202 306 203
rect 304 202 305 203
rect 303 202 304 203
rect 302 202 303 203
rect 301 202 302 203
rect 300 202 301 203
rect 299 202 300 203
rect 298 202 299 203
rect 297 202 298 203
rect 296 202 297 203
rect 295 202 296 203
rect 294 202 295 203
rect 293 202 294 203
rect 292 202 293 203
rect 291 202 292 203
rect 290 202 291 203
rect 289 202 290 203
rect 288 202 289 203
rect 287 202 288 203
rect 286 202 287 203
rect 285 202 286 203
rect 284 202 285 203
rect 283 202 284 203
rect 282 202 283 203
rect 281 202 282 203
rect 280 202 281 203
rect 279 202 280 203
rect 278 202 279 203
rect 277 202 278 203
rect 276 202 277 203
rect 275 202 276 203
rect 274 202 275 203
rect 273 202 274 203
rect 272 202 273 203
rect 271 202 272 203
rect 270 202 271 203
rect 269 202 270 203
rect 268 202 269 203
rect 267 202 268 203
rect 266 202 267 203
rect 265 202 266 203
rect 264 202 265 203
rect 263 202 264 203
rect 262 202 263 203
rect 261 202 262 203
rect 260 202 261 203
rect 259 202 260 203
rect 258 202 259 203
rect 257 202 258 203
rect 256 202 257 203
rect 255 202 256 203
rect 254 202 255 203
rect 253 202 254 203
rect 245 202 246 203
rect 244 202 245 203
rect 243 202 244 203
rect 242 202 243 203
rect 241 202 242 203
rect 240 202 241 203
rect 239 202 240 203
rect 238 202 239 203
rect 237 202 238 203
rect 236 202 237 203
rect 235 202 236 203
rect 234 202 235 203
rect 233 202 234 203
rect 232 202 233 203
rect 231 202 232 203
rect 230 202 231 203
rect 229 202 230 203
rect 228 202 229 203
rect 227 202 228 203
rect 226 202 227 203
rect 225 202 226 203
rect 224 202 225 203
rect 223 202 224 203
rect 222 202 223 203
rect 221 202 222 203
rect 220 202 221 203
rect 219 202 220 203
rect 218 202 219 203
rect 217 202 218 203
rect 216 202 217 203
rect 215 202 216 203
rect 214 202 215 203
rect 213 202 214 203
rect 212 202 213 203
rect 211 202 212 203
rect 210 202 211 203
rect 209 202 210 203
rect 208 202 209 203
rect 207 202 208 203
rect 206 202 207 203
rect 205 202 206 203
rect 204 202 205 203
rect 203 202 204 203
rect 173 202 174 203
rect 172 202 173 203
rect 171 202 172 203
rect 170 202 171 203
rect 169 202 170 203
rect 168 202 169 203
rect 167 202 168 203
rect 166 202 167 203
rect 165 202 166 203
rect 164 202 165 203
rect 163 202 164 203
rect 162 202 163 203
rect 161 202 162 203
rect 160 202 161 203
rect 159 202 160 203
rect 158 202 159 203
rect 157 202 158 203
rect 156 202 157 203
rect 155 202 156 203
rect 154 202 155 203
rect 153 202 154 203
rect 152 202 153 203
rect 151 202 152 203
rect 150 202 151 203
rect 149 202 150 203
rect 148 202 149 203
rect 147 202 148 203
rect 146 202 147 203
rect 145 202 146 203
rect 144 202 145 203
rect 143 202 144 203
rect 142 202 143 203
rect 141 202 142 203
rect 140 202 141 203
rect 139 202 140 203
rect 138 202 139 203
rect 137 202 138 203
rect 136 202 137 203
rect 135 202 136 203
rect 134 202 135 203
rect 133 202 134 203
rect 132 202 133 203
rect 131 202 132 203
rect 130 202 131 203
rect 129 202 130 203
rect 128 202 129 203
rect 127 202 128 203
rect 126 202 127 203
rect 125 202 126 203
rect 124 202 125 203
rect 123 202 124 203
rect 122 202 123 203
rect 121 202 122 203
rect 120 202 121 203
rect 119 202 120 203
rect 118 202 119 203
rect 117 202 118 203
rect 116 202 117 203
rect 115 202 116 203
rect 114 202 115 203
rect 113 202 114 203
rect 112 202 113 203
rect 111 202 112 203
rect 110 202 111 203
rect 109 202 110 203
rect 108 202 109 203
rect 107 202 108 203
rect 106 202 107 203
rect 105 202 106 203
rect 104 202 105 203
rect 103 202 104 203
rect 102 202 103 203
rect 101 202 102 203
rect 100 202 101 203
rect 99 202 100 203
rect 98 202 99 203
rect 97 202 98 203
rect 96 202 97 203
rect 95 202 96 203
rect 94 202 95 203
rect 93 202 94 203
rect 92 202 93 203
rect 91 202 92 203
rect 90 202 91 203
rect 89 202 90 203
rect 88 202 89 203
rect 87 202 88 203
rect 86 202 87 203
rect 85 202 86 203
rect 84 202 85 203
rect 83 202 84 203
rect 82 202 83 203
rect 81 202 82 203
rect 80 202 81 203
rect 79 202 80 203
rect 78 202 79 203
rect 77 202 78 203
rect 76 202 77 203
rect 75 202 76 203
rect 74 202 75 203
rect 73 202 74 203
rect 72 202 73 203
rect 55 202 56 203
rect 54 202 55 203
rect 53 202 54 203
rect 52 202 53 203
rect 51 202 52 203
rect 50 202 51 203
rect 49 202 50 203
rect 48 202 49 203
rect 47 202 48 203
rect 46 202 47 203
rect 45 202 46 203
rect 44 202 45 203
rect 43 202 44 203
rect 42 202 43 203
rect 41 202 42 203
rect 40 202 41 203
rect 39 202 40 203
rect 38 202 39 203
rect 37 202 38 203
rect 36 202 37 203
rect 35 202 36 203
rect 34 202 35 203
rect 33 202 34 203
rect 32 202 33 203
rect 31 202 32 203
rect 30 202 31 203
rect 29 202 30 203
rect 28 202 29 203
rect 27 202 28 203
rect 26 202 27 203
rect 25 202 26 203
rect 24 202 25 203
rect 23 202 24 203
rect 22 202 23 203
rect 21 202 22 203
rect 20 202 21 203
rect 19 202 20 203
rect 18 202 19 203
rect 17 202 18 203
rect 16 202 17 203
rect 15 202 16 203
rect 14 202 15 203
rect 13 202 14 203
rect 12 202 13 203
rect 11 202 12 203
rect 10 202 11 203
rect 9 202 10 203
rect 8 202 9 203
rect 478 203 479 204
rect 477 203 478 204
rect 476 203 477 204
rect 462 203 463 204
rect 461 203 462 204
rect 460 203 461 204
rect 459 203 460 204
rect 458 203 459 204
rect 351 203 352 204
rect 350 203 351 204
rect 349 203 350 204
rect 348 203 349 204
rect 347 203 348 204
rect 346 203 347 204
rect 345 203 346 204
rect 344 203 345 204
rect 343 203 344 204
rect 342 203 343 204
rect 341 203 342 204
rect 340 203 341 204
rect 339 203 340 204
rect 338 203 339 204
rect 337 203 338 204
rect 336 203 337 204
rect 335 203 336 204
rect 334 203 335 204
rect 333 203 334 204
rect 332 203 333 204
rect 331 203 332 204
rect 330 203 331 204
rect 329 203 330 204
rect 328 203 329 204
rect 327 203 328 204
rect 326 203 327 204
rect 325 203 326 204
rect 324 203 325 204
rect 323 203 324 204
rect 322 203 323 204
rect 321 203 322 204
rect 320 203 321 204
rect 319 203 320 204
rect 318 203 319 204
rect 317 203 318 204
rect 316 203 317 204
rect 315 203 316 204
rect 314 203 315 204
rect 313 203 314 204
rect 312 203 313 204
rect 311 203 312 204
rect 310 203 311 204
rect 309 203 310 204
rect 308 203 309 204
rect 307 203 308 204
rect 306 203 307 204
rect 305 203 306 204
rect 304 203 305 204
rect 303 203 304 204
rect 302 203 303 204
rect 301 203 302 204
rect 300 203 301 204
rect 299 203 300 204
rect 298 203 299 204
rect 297 203 298 204
rect 296 203 297 204
rect 295 203 296 204
rect 294 203 295 204
rect 293 203 294 204
rect 292 203 293 204
rect 291 203 292 204
rect 290 203 291 204
rect 289 203 290 204
rect 288 203 289 204
rect 287 203 288 204
rect 286 203 287 204
rect 285 203 286 204
rect 284 203 285 204
rect 283 203 284 204
rect 282 203 283 204
rect 281 203 282 204
rect 280 203 281 204
rect 279 203 280 204
rect 278 203 279 204
rect 277 203 278 204
rect 276 203 277 204
rect 275 203 276 204
rect 274 203 275 204
rect 273 203 274 204
rect 272 203 273 204
rect 271 203 272 204
rect 270 203 271 204
rect 269 203 270 204
rect 268 203 269 204
rect 267 203 268 204
rect 266 203 267 204
rect 265 203 266 204
rect 264 203 265 204
rect 263 203 264 204
rect 262 203 263 204
rect 261 203 262 204
rect 260 203 261 204
rect 259 203 260 204
rect 258 203 259 204
rect 257 203 258 204
rect 256 203 257 204
rect 255 203 256 204
rect 254 203 255 204
rect 253 203 254 204
rect 252 203 253 204
rect 251 203 252 204
rect 245 203 246 204
rect 244 203 245 204
rect 243 203 244 204
rect 242 203 243 204
rect 241 203 242 204
rect 240 203 241 204
rect 239 203 240 204
rect 238 203 239 204
rect 237 203 238 204
rect 236 203 237 204
rect 235 203 236 204
rect 234 203 235 204
rect 233 203 234 204
rect 232 203 233 204
rect 231 203 232 204
rect 230 203 231 204
rect 229 203 230 204
rect 228 203 229 204
rect 227 203 228 204
rect 226 203 227 204
rect 225 203 226 204
rect 224 203 225 204
rect 223 203 224 204
rect 222 203 223 204
rect 221 203 222 204
rect 220 203 221 204
rect 219 203 220 204
rect 218 203 219 204
rect 217 203 218 204
rect 216 203 217 204
rect 215 203 216 204
rect 214 203 215 204
rect 213 203 214 204
rect 212 203 213 204
rect 211 203 212 204
rect 210 203 211 204
rect 209 203 210 204
rect 208 203 209 204
rect 207 203 208 204
rect 206 203 207 204
rect 205 203 206 204
rect 204 203 205 204
rect 203 203 204 204
rect 202 203 203 204
rect 171 203 172 204
rect 170 203 171 204
rect 169 203 170 204
rect 168 203 169 204
rect 167 203 168 204
rect 166 203 167 204
rect 165 203 166 204
rect 164 203 165 204
rect 163 203 164 204
rect 162 203 163 204
rect 161 203 162 204
rect 160 203 161 204
rect 159 203 160 204
rect 158 203 159 204
rect 157 203 158 204
rect 156 203 157 204
rect 155 203 156 204
rect 154 203 155 204
rect 153 203 154 204
rect 152 203 153 204
rect 151 203 152 204
rect 150 203 151 204
rect 149 203 150 204
rect 148 203 149 204
rect 147 203 148 204
rect 146 203 147 204
rect 145 203 146 204
rect 144 203 145 204
rect 143 203 144 204
rect 142 203 143 204
rect 141 203 142 204
rect 140 203 141 204
rect 139 203 140 204
rect 138 203 139 204
rect 137 203 138 204
rect 136 203 137 204
rect 135 203 136 204
rect 134 203 135 204
rect 133 203 134 204
rect 132 203 133 204
rect 131 203 132 204
rect 130 203 131 204
rect 129 203 130 204
rect 128 203 129 204
rect 127 203 128 204
rect 126 203 127 204
rect 125 203 126 204
rect 124 203 125 204
rect 123 203 124 204
rect 122 203 123 204
rect 121 203 122 204
rect 120 203 121 204
rect 119 203 120 204
rect 118 203 119 204
rect 117 203 118 204
rect 116 203 117 204
rect 115 203 116 204
rect 114 203 115 204
rect 113 203 114 204
rect 112 203 113 204
rect 111 203 112 204
rect 110 203 111 204
rect 109 203 110 204
rect 108 203 109 204
rect 107 203 108 204
rect 106 203 107 204
rect 105 203 106 204
rect 104 203 105 204
rect 103 203 104 204
rect 102 203 103 204
rect 101 203 102 204
rect 100 203 101 204
rect 99 203 100 204
rect 98 203 99 204
rect 97 203 98 204
rect 96 203 97 204
rect 95 203 96 204
rect 94 203 95 204
rect 93 203 94 204
rect 92 203 93 204
rect 91 203 92 204
rect 90 203 91 204
rect 89 203 90 204
rect 88 203 89 204
rect 87 203 88 204
rect 86 203 87 204
rect 85 203 86 204
rect 84 203 85 204
rect 83 203 84 204
rect 82 203 83 204
rect 81 203 82 204
rect 80 203 81 204
rect 79 203 80 204
rect 78 203 79 204
rect 77 203 78 204
rect 76 203 77 204
rect 75 203 76 204
rect 74 203 75 204
rect 73 203 74 204
rect 56 203 57 204
rect 55 203 56 204
rect 54 203 55 204
rect 53 203 54 204
rect 52 203 53 204
rect 51 203 52 204
rect 50 203 51 204
rect 49 203 50 204
rect 48 203 49 204
rect 47 203 48 204
rect 46 203 47 204
rect 45 203 46 204
rect 44 203 45 204
rect 43 203 44 204
rect 42 203 43 204
rect 41 203 42 204
rect 40 203 41 204
rect 39 203 40 204
rect 38 203 39 204
rect 37 203 38 204
rect 36 203 37 204
rect 35 203 36 204
rect 34 203 35 204
rect 33 203 34 204
rect 32 203 33 204
rect 31 203 32 204
rect 30 203 31 204
rect 29 203 30 204
rect 28 203 29 204
rect 27 203 28 204
rect 26 203 27 204
rect 25 203 26 204
rect 24 203 25 204
rect 23 203 24 204
rect 22 203 23 204
rect 21 203 22 204
rect 20 203 21 204
rect 19 203 20 204
rect 18 203 19 204
rect 17 203 18 204
rect 16 203 17 204
rect 15 203 16 204
rect 14 203 15 204
rect 13 203 14 204
rect 12 203 13 204
rect 11 203 12 204
rect 10 203 11 204
rect 9 203 10 204
rect 8 203 9 204
rect 478 204 479 205
rect 477 204 478 205
rect 476 204 477 205
rect 475 204 476 205
rect 474 204 475 205
rect 462 204 463 205
rect 461 204 462 205
rect 460 204 461 205
rect 351 204 352 205
rect 350 204 351 205
rect 349 204 350 205
rect 348 204 349 205
rect 347 204 348 205
rect 346 204 347 205
rect 345 204 346 205
rect 344 204 345 205
rect 343 204 344 205
rect 342 204 343 205
rect 341 204 342 205
rect 340 204 341 205
rect 339 204 340 205
rect 338 204 339 205
rect 337 204 338 205
rect 336 204 337 205
rect 335 204 336 205
rect 334 204 335 205
rect 333 204 334 205
rect 332 204 333 205
rect 331 204 332 205
rect 330 204 331 205
rect 329 204 330 205
rect 328 204 329 205
rect 327 204 328 205
rect 326 204 327 205
rect 325 204 326 205
rect 324 204 325 205
rect 323 204 324 205
rect 322 204 323 205
rect 321 204 322 205
rect 320 204 321 205
rect 319 204 320 205
rect 318 204 319 205
rect 317 204 318 205
rect 316 204 317 205
rect 315 204 316 205
rect 314 204 315 205
rect 313 204 314 205
rect 312 204 313 205
rect 311 204 312 205
rect 310 204 311 205
rect 309 204 310 205
rect 308 204 309 205
rect 307 204 308 205
rect 306 204 307 205
rect 305 204 306 205
rect 304 204 305 205
rect 303 204 304 205
rect 302 204 303 205
rect 301 204 302 205
rect 300 204 301 205
rect 299 204 300 205
rect 298 204 299 205
rect 297 204 298 205
rect 296 204 297 205
rect 295 204 296 205
rect 294 204 295 205
rect 293 204 294 205
rect 292 204 293 205
rect 291 204 292 205
rect 290 204 291 205
rect 289 204 290 205
rect 288 204 289 205
rect 287 204 288 205
rect 286 204 287 205
rect 285 204 286 205
rect 284 204 285 205
rect 283 204 284 205
rect 282 204 283 205
rect 281 204 282 205
rect 280 204 281 205
rect 279 204 280 205
rect 278 204 279 205
rect 277 204 278 205
rect 276 204 277 205
rect 275 204 276 205
rect 274 204 275 205
rect 273 204 274 205
rect 272 204 273 205
rect 271 204 272 205
rect 270 204 271 205
rect 269 204 270 205
rect 268 204 269 205
rect 267 204 268 205
rect 266 204 267 205
rect 265 204 266 205
rect 264 204 265 205
rect 263 204 264 205
rect 262 204 263 205
rect 261 204 262 205
rect 260 204 261 205
rect 259 204 260 205
rect 258 204 259 205
rect 257 204 258 205
rect 256 204 257 205
rect 255 204 256 205
rect 254 204 255 205
rect 253 204 254 205
rect 252 204 253 205
rect 251 204 252 205
rect 250 204 251 205
rect 249 204 250 205
rect 244 204 245 205
rect 243 204 244 205
rect 242 204 243 205
rect 241 204 242 205
rect 240 204 241 205
rect 239 204 240 205
rect 238 204 239 205
rect 237 204 238 205
rect 236 204 237 205
rect 235 204 236 205
rect 234 204 235 205
rect 233 204 234 205
rect 232 204 233 205
rect 231 204 232 205
rect 230 204 231 205
rect 229 204 230 205
rect 228 204 229 205
rect 227 204 228 205
rect 226 204 227 205
rect 225 204 226 205
rect 224 204 225 205
rect 223 204 224 205
rect 222 204 223 205
rect 221 204 222 205
rect 220 204 221 205
rect 219 204 220 205
rect 218 204 219 205
rect 217 204 218 205
rect 216 204 217 205
rect 215 204 216 205
rect 214 204 215 205
rect 213 204 214 205
rect 212 204 213 205
rect 211 204 212 205
rect 210 204 211 205
rect 209 204 210 205
rect 208 204 209 205
rect 207 204 208 205
rect 206 204 207 205
rect 205 204 206 205
rect 204 204 205 205
rect 203 204 204 205
rect 202 204 203 205
rect 201 204 202 205
rect 169 204 170 205
rect 168 204 169 205
rect 167 204 168 205
rect 166 204 167 205
rect 165 204 166 205
rect 164 204 165 205
rect 163 204 164 205
rect 162 204 163 205
rect 161 204 162 205
rect 160 204 161 205
rect 159 204 160 205
rect 158 204 159 205
rect 157 204 158 205
rect 156 204 157 205
rect 155 204 156 205
rect 154 204 155 205
rect 153 204 154 205
rect 152 204 153 205
rect 151 204 152 205
rect 150 204 151 205
rect 149 204 150 205
rect 148 204 149 205
rect 147 204 148 205
rect 146 204 147 205
rect 145 204 146 205
rect 144 204 145 205
rect 143 204 144 205
rect 142 204 143 205
rect 141 204 142 205
rect 140 204 141 205
rect 139 204 140 205
rect 138 204 139 205
rect 137 204 138 205
rect 136 204 137 205
rect 135 204 136 205
rect 134 204 135 205
rect 133 204 134 205
rect 132 204 133 205
rect 131 204 132 205
rect 130 204 131 205
rect 129 204 130 205
rect 128 204 129 205
rect 127 204 128 205
rect 126 204 127 205
rect 125 204 126 205
rect 124 204 125 205
rect 123 204 124 205
rect 122 204 123 205
rect 121 204 122 205
rect 120 204 121 205
rect 119 204 120 205
rect 118 204 119 205
rect 117 204 118 205
rect 116 204 117 205
rect 115 204 116 205
rect 114 204 115 205
rect 113 204 114 205
rect 112 204 113 205
rect 111 204 112 205
rect 110 204 111 205
rect 109 204 110 205
rect 108 204 109 205
rect 107 204 108 205
rect 106 204 107 205
rect 105 204 106 205
rect 104 204 105 205
rect 103 204 104 205
rect 102 204 103 205
rect 101 204 102 205
rect 100 204 101 205
rect 99 204 100 205
rect 98 204 99 205
rect 97 204 98 205
rect 96 204 97 205
rect 95 204 96 205
rect 94 204 95 205
rect 93 204 94 205
rect 92 204 93 205
rect 91 204 92 205
rect 90 204 91 205
rect 89 204 90 205
rect 88 204 89 205
rect 87 204 88 205
rect 86 204 87 205
rect 85 204 86 205
rect 84 204 85 205
rect 83 204 84 205
rect 82 204 83 205
rect 81 204 82 205
rect 80 204 81 205
rect 79 204 80 205
rect 78 204 79 205
rect 77 204 78 205
rect 76 204 77 205
rect 75 204 76 205
rect 74 204 75 205
rect 56 204 57 205
rect 55 204 56 205
rect 54 204 55 205
rect 53 204 54 205
rect 52 204 53 205
rect 51 204 52 205
rect 50 204 51 205
rect 49 204 50 205
rect 48 204 49 205
rect 47 204 48 205
rect 46 204 47 205
rect 45 204 46 205
rect 44 204 45 205
rect 43 204 44 205
rect 42 204 43 205
rect 41 204 42 205
rect 40 204 41 205
rect 39 204 40 205
rect 38 204 39 205
rect 37 204 38 205
rect 36 204 37 205
rect 35 204 36 205
rect 34 204 35 205
rect 33 204 34 205
rect 32 204 33 205
rect 31 204 32 205
rect 30 204 31 205
rect 29 204 30 205
rect 28 204 29 205
rect 27 204 28 205
rect 26 204 27 205
rect 25 204 26 205
rect 24 204 25 205
rect 23 204 24 205
rect 22 204 23 205
rect 21 204 22 205
rect 20 204 21 205
rect 19 204 20 205
rect 18 204 19 205
rect 17 204 18 205
rect 16 204 17 205
rect 15 204 16 205
rect 14 204 15 205
rect 13 204 14 205
rect 12 204 13 205
rect 11 204 12 205
rect 10 204 11 205
rect 9 204 10 205
rect 8 204 9 205
rect 477 205 478 206
rect 476 205 477 206
rect 475 205 476 206
rect 474 205 475 206
rect 473 205 474 206
rect 420 205 421 206
rect 419 205 420 206
rect 418 205 419 206
rect 417 205 418 206
rect 416 205 417 206
rect 415 205 416 206
rect 414 205 415 206
rect 413 205 414 206
rect 412 205 413 206
rect 411 205 412 206
rect 352 205 353 206
rect 351 205 352 206
rect 350 205 351 206
rect 349 205 350 206
rect 348 205 349 206
rect 347 205 348 206
rect 346 205 347 206
rect 345 205 346 206
rect 344 205 345 206
rect 343 205 344 206
rect 342 205 343 206
rect 341 205 342 206
rect 340 205 341 206
rect 339 205 340 206
rect 338 205 339 206
rect 337 205 338 206
rect 336 205 337 206
rect 335 205 336 206
rect 334 205 335 206
rect 333 205 334 206
rect 332 205 333 206
rect 331 205 332 206
rect 330 205 331 206
rect 329 205 330 206
rect 328 205 329 206
rect 327 205 328 206
rect 326 205 327 206
rect 325 205 326 206
rect 324 205 325 206
rect 323 205 324 206
rect 322 205 323 206
rect 321 205 322 206
rect 320 205 321 206
rect 319 205 320 206
rect 318 205 319 206
rect 317 205 318 206
rect 316 205 317 206
rect 315 205 316 206
rect 314 205 315 206
rect 313 205 314 206
rect 312 205 313 206
rect 311 205 312 206
rect 310 205 311 206
rect 309 205 310 206
rect 308 205 309 206
rect 307 205 308 206
rect 306 205 307 206
rect 305 205 306 206
rect 304 205 305 206
rect 303 205 304 206
rect 302 205 303 206
rect 301 205 302 206
rect 300 205 301 206
rect 299 205 300 206
rect 298 205 299 206
rect 297 205 298 206
rect 296 205 297 206
rect 295 205 296 206
rect 294 205 295 206
rect 293 205 294 206
rect 292 205 293 206
rect 291 205 292 206
rect 290 205 291 206
rect 289 205 290 206
rect 288 205 289 206
rect 287 205 288 206
rect 286 205 287 206
rect 285 205 286 206
rect 284 205 285 206
rect 283 205 284 206
rect 282 205 283 206
rect 281 205 282 206
rect 280 205 281 206
rect 279 205 280 206
rect 278 205 279 206
rect 277 205 278 206
rect 276 205 277 206
rect 275 205 276 206
rect 274 205 275 206
rect 273 205 274 206
rect 272 205 273 206
rect 271 205 272 206
rect 270 205 271 206
rect 269 205 270 206
rect 268 205 269 206
rect 267 205 268 206
rect 266 205 267 206
rect 265 205 266 206
rect 264 205 265 206
rect 263 205 264 206
rect 262 205 263 206
rect 261 205 262 206
rect 260 205 261 206
rect 259 205 260 206
rect 258 205 259 206
rect 257 205 258 206
rect 256 205 257 206
rect 255 205 256 206
rect 254 205 255 206
rect 253 205 254 206
rect 252 205 253 206
rect 251 205 252 206
rect 250 205 251 206
rect 249 205 250 206
rect 248 205 249 206
rect 247 205 248 206
rect 246 205 247 206
rect 245 205 246 206
rect 244 205 245 206
rect 243 205 244 206
rect 242 205 243 206
rect 241 205 242 206
rect 240 205 241 206
rect 239 205 240 206
rect 238 205 239 206
rect 237 205 238 206
rect 236 205 237 206
rect 235 205 236 206
rect 234 205 235 206
rect 233 205 234 206
rect 232 205 233 206
rect 231 205 232 206
rect 230 205 231 206
rect 229 205 230 206
rect 228 205 229 206
rect 227 205 228 206
rect 226 205 227 206
rect 225 205 226 206
rect 224 205 225 206
rect 223 205 224 206
rect 222 205 223 206
rect 221 205 222 206
rect 220 205 221 206
rect 219 205 220 206
rect 218 205 219 206
rect 217 205 218 206
rect 216 205 217 206
rect 215 205 216 206
rect 214 205 215 206
rect 213 205 214 206
rect 212 205 213 206
rect 211 205 212 206
rect 210 205 211 206
rect 209 205 210 206
rect 208 205 209 206
rect 207 205 208 206
rect 206 205 207 206
rect 205 205 206 206
rect 204 205 205 206
rect 203 205 204 206
rect 202 205 203 206
rect 201 205 202 206
rect 200 205 201 206
rect 167 205 168 206
rect 166 205 167 206
rect 165 205 166 206
rect 164 205 165 206
rect 163 205 164 206
rect 162 205 163 206
rect 161 205 162 206
rect 160 205 161 206
rect 159 205 160 206
rect 158 205 159 206
rect 157 205 158 206
rect 156 205 157 206
rect 155 205 156 206
rect 154 205 155 206
rect 153 205 154 206
rect 152 205 153 206
rect 151 205 152 206
rect 150 205 151 206
rect 149 205 150 206
rect 148 205 149 206
rect 147 205 148 206
rect 146 205 147 206
rect 145 205 146 206
rect 144 205 145 206
rect 143 205 144 206
rect 142 205 143 206
rect 141 205 142 206
rect 140 205 141 206
rect 139 205 140 206
rect 138 205 139 206
rect 137 205 138 206
rect 136 205 137 206
rect 135 205 136 206
rect 134 205 135 206
rect 133 205 134 206
rect 132 205 133 206
rect 131 205 132 206
rect 130 205 131 206
rect 129 205 130 206
rect 128 205 129 206
rect 127 205 128 206
rect 126 205 127 206
rect 125 205 126 206
rect 124 205 125 206
rect 123 205 124 206
rect 122 205 123 206
rect 121 205 122 206
rect 120 205 121 206
rect 119 205 120 206
rect 118 205 119 206
rect 117 205 118 206
rect 116 205 117 206
rect 115 205 116 206
rect 114 205 115 206
rect 113 205 114 206
rect 112 205 113 206
rect 111 205 112 206
rect 110 205 111 206
rect 109 205 110 206
rect 108 205 109 206
rect 107 205 108 206
rect 106 205 107 206
rect 105 205 106 206
rect 104 205 105 206
rect 103 205 104 206
rect 102 205 103 206
rect 101 205 102 206
rect 100 205 101 206
rect 99 205 100 206
rect 98 205 99 206
rect 97 205 98 206
rect 96 205 97 206
rect 95 205 96 206
rect 94 205 95 206
rect 93 205 94 206
rect 92 205 93 206
rect 91 205 92 206
rect 90 205 91 206
rect 89 205 90 206
rect 88 205 89 206
rect 87 205 88 206
rect 86 205 87 206
rect 85 205 86 206
rect 84 205 85 206
rect 83 205 84 206
rect 82 205 83 206
rect 81 205 82 206
rect 80 205 81 206
rect 79 205 80 206
rect 78 205 79 206
rect 77 205 78 206
rect 76 205 77 206
rect 57 205 58 206
rect 56 205 57 206
rect 55 205 56 206
rect 54 205 55 206
rect 53 205 54 206
rect 52 205 53 206
rect 51 205 52 206
rect 50 205 51 206
rect 49 205 50 206
rect 48 205 49 206
rect 47 205 48 206
rect 46 205 47 206
rect 45 205 46 206
rect 44 205 45 206
rect 43 205 44 206
rect 42 205 43 206
rect 41 205 42 206
rect 40 205 41 206
rect 39 205 40 206
rect 38 205 39 206
rect 37 205 38 206
rect 36 205 37 206
rect 35 205 36 206
rect 34 205 35 206
rect 33 205 34 206
rect 32 205 33 206
rect 31 205 32 206
rect 30 205 31 206
rect 29 205 30 206
rect 28 205 29 206
rect 27 205 28 206
rect 26 205 27 206
rect 25 205 26 206
rect 24 205 25 206
rect 23 205 24 206
rect 22 205 23 206
rect 21 205 22 206
rect 20 205 21 206
rect 19 205 20 206
rect 18 205 19 206
rect 17 205 18 206
rect 16 205 17 206
rect 15 205 16 206
rect 14 205 15 206
rect 13 205 14 206
rect 12 205 13 206
rect 11 205 12 206
rect 10 205 11 206
rect 9 205 10 206
rect 8 205 9 206
rect 424 206 425 207
rect 423 206 424 207
rect 422 206 423 207
rect 421 206 422 207
rect 420 206 421 207
rect 419 206 420 207
rect 418 206 419 207
rect 417 206 418 207
rect 416 206 417 207
rect 415 206 416 207
rect 414 206 415 207
rect 413 206 414 207
rect 412 206 413 207
rect 411 206 412 207
rect 410 206 411 207
rect 409 206 410 207
rect 408 206 409 207
rect 353 206 354 207
rect 352 206 353 207
rect 351 206 352 207
rect 350 206 351 207
rect 349 206 350 207
rect 348 206 349 207
rect 347 206 348 207
rect 346 206 347 207
rect 345 206 346 207
rect 344 206 345 207
rect 343 206 344 207
rect 342 206 343 207
rect 341 206 342 207
rect 340 206 341 207
rect 339 206 340 207
rect 338 206 339 207
rect 337 206 338 207
rect 336 206 337 207
rect 335 206 336 207
rect 334 206 335 207
rect 333 206 334 207
rect 332 206 333 207
rect 331 206 332 207
rect 330 206 331 207
rect 329 206 330 207
rect 328 206 329 207
rect 327 206 328 207
rect 326 206 327 207
rect 325 206 326 207
rect 324 206 325 207
rect 323 206 324 207
rect 322 206 323 207
rect 321 206 322 207
rect 320 206 321 207
rect 319 206 320 207
rect 318 206 319 207
rect 317 206 318 207
rect 316 206 317 207
rect 315 206 316 207
rect 314 206 315 207
rect 313 206 314 207
rect 312 206 313 207
rect 311 206 312 207
rect 310 206 311 207
rect 309 206 310 207
rect 308 206 309 207
rect 307 206 308 207
rect 306 206 307 207
rect 305 206 306 207
rect 304 206 305 207
rect 303 206 304 207
rect 302 206 303 207
rect 301 206 302 207
rect 300 206 301 207
rect 299 206 300 207
rect 298 206 299 207
rect 297 206 298 207
rect 296 206 297 207
rect 295 206 296 207
rect 294 206 295 207
rect 293 206 294 207
rect 292 206 293 207
rect 291 206 292 207
rect 290 206 291 207
rect 289 206 290 207
rect 288 206 289 207
rect 287 206 288 207
rect 286 206 287 207
rect 285 206 286 207
rect 284 206 285 207
rect 283 206 284 207
rect 282 206 283 207
rect 281 206 282 207
rect 280 206 281 207
rect 279 206 280 207
rect 278 206 279 207
rect 277 206 278 207
rect 276 206 277 207
rect 275 206 276 207
rect 274 206 275 207
rect 273 206 274 207
rect 272 206 273 207
rect 271 206 272 207
rect 270 206 271 207
rect 269 206 270 207
rect 268 206 269 207
rect 267 206 268 207
rect 266 206 267 207
rect 265 206 266 207
rect 264 206 265 207
rect 263 206 264 207
rect 262 206 263 207
rect 261 206 262 207
rect 260 206 261 207
rect 259 206 260 207
rect 258 206 259 207
rect 257 206 258 207
rect 256 206 257 207
rect 255 206 256 207
rect 254 206 255 207
rect 253 206 254 207
rect 252 206 253 207
rect 251 206 252 207
rect 250 206 251 207
rect 249 206 250 207
rect 248 206 249 207
rect 247 206 248 207
rect 246 206 247 207
rect 245 206 246 207
rect 244 206 245 207
rect 243 206 244 207
rect 242 206 243 207
rect 241 206 242 207
rect 240 206 241 207
rect 239 206 240 207
rect 238 206 239 207
rect 237 206 238 207
rect 236 206 237 207
rect 235 206 236 207
rect 234 206 235 207
rect 233 206 234 207
rect 232 206 233 207
rect 231 206 232 207
rect 230 206 231 207
rect 229 206 230 207
rect 228 206 229 207
rect 227 206 228 207
rect 226 206 227 207
rect 225 206 226 207
rect 224 206 225 207
rect 223 206 224 207
rect 222 206 223 207
rect 221 206 222 207
rect 220 206 221 207
rect 219 206 220 207
rect 218 206 219 207
rect 217 206 218 207
rect 216 206 217 207
rect 215 206 216 207
rect 214 206 215 207
rect 213 206 214 207
rect 212 206 213 207
rect 211 206 212 207
rect 210 206 211 207
rect 209 206 210 207
rect 208 206 209 207
rect 207 206 208 207
rect 206 206 207 207
rect 205 206 206 207
rect 204 206 205 207
rect 203 206 204 207
rect 202 206 203 207
rect 201 206 202 207
rect 200 206 201 207
rect 199 206 200 207
rect 198 206 199 207
rect 165 206 166 207
rect 164 206 165 207
rect 163 206 164 207
rect 162 206 163 207
rect 161 206 162 207
rect 160 206 161 207
rect 159 206 160 207
rect 158 206 159 207
rect 157 206 158 207
rect 156 206 157 207
rect 155 206 156 207
rect 154 206 155 207
rect 153 206 154 207
rect 152 206 153 207
rect 151 206 152 207
rect 150 206 151 207
rect 149 206 150 207
rect 148 206 149 207
rect 147 206 148 207
rect 146 206 147 207
rect 145 206 146 207
rect 144 206 145 207
rect 143 206 144 207
rect 142 206 143 207
rect 141 206 142 207
rect 140 206 141 207
rect 139 206 140 207
rect 138 206 139 207
rect 137 206 138 207
rect 136 206 137 207
rect 135 206 136 207
rect 134 206 135 207
rect 133 206 134 207
rect 132 206 133 207
rect 131 206 132 207
rect 130 206 131 207
rect 129 206 130 207
rect 128 206 129 207
rect 127 206 128 207
rect 126 206 127 207
rect 125 206 126 207
rect 124 206 125 207
rect 123 206 124 207
rect 122 206 123 207
rect 121 206 122 207
rect 120 206 121 207
rect 119 206 120 207
rect 118 206 119 207
rect 117 206 118 207
rect 116 206 117 207
rect 115 206 116 207
rect 114 206 115 207
rect 113 206 114 207
rect 112 206 113 207
rect 111 206 112 207
rect 110 206 111 207
rect 109 206 110 207
rect 108 206 109 207
rect 107 206 108 207
rect 106 206 107 207
rect 105 206 106 207
rect 104 206 105 207
rect 103 206 104 207
rect 102 206 103 207
rect 101 206 102 207
rect 100 206 101 207
rect 99 206 100 207
rect 98 206 99 207
rect 97 206 98 207
rect 96 206 97 207
rect 95 206 96 207
rect 94 206 95 207
rect 93 206 94 207
rect 92 206 93 207
rect 91 206 92 207
rect 90 206 91 207
rect 89 206 90 207
rect 88 206 89 207
rect 87 206 88 207
rect 86 206 87 207
rect 85 206 86 207
rect 84 206 85 207
rect 83 206 84 207
rect 82 206 83 207
rect 81 206 82 207
rect 80 206 81 207
rect 79 206 80 207
rect 78 206 79 207
rect 77 206 78 207
rect 58 206 59 207
rect 57 206 58 207
rect 56 206 57 207
rect 55 206 56 207
rect 54 206 55 207
rect 53 206 54 207
rect 52 206 53 207
rect 51 206 52 207
rect 50 206 51 207
rect 49 206 50 207
rect 48 206 49 207
rect 47 206 48 207
rect 46 206 47 207
rect 45 206 46 207
rect 44 206 45 207
rect 43 206 44 207
rect 42 206 43 207
rect 41 206 42 207
rect 40 206 41 207
rect 39 206 40 207
rect 38 206 39 207
rect 37 206 38 207
rect 36 206 37 207
rect 35 206 36 207
rect 34 206 35 207
rect 33 206 34 207
rect 32 206 33 207
rect 31 206 32 207
rect 30 206 31 207
rect 29 206 30 207
rect 28 206 29 207
rect 27 206 28 207
rect 26 206 27 207
rect 25 206 26 207
rect 24 206 25 207
rect 23 206 24 207
rect 22 206 23 207
rect 21 206 22 207
rect 20 206 21 207
rect 19 206 20 207
rect 18 206 19 207
rect 17 206 18 207
rect 16 206 17 207
rect 15 206 16 207
rect 14 206 15 207
rect 13 206 14 207
rect 12 206 13 207
rect 11 206 12 207
rect 10 206 11 207
rect 9 206 10 207
rect 8 206 9 207
rect 426 207 427 208
rect 425 207 426 208
rect 424 207 425 208
rect 423 207 424 208
rect 422 207 423 208
rect 421 207 422 208
rect 420 207 421 208
rect 419 207 420 208
rect 418 207 419 208
rect 417 207 418 208
rect 416 207 417 208
rect 415 207 416 208
rect 414 207 415 208
rect 413 207 414 208
rect 412 207 413 208
rect 411 207 412 208
rect 410 207 411 208
rect 409 207 410 208
rect 408 207 409 208
rect 407 207 408 208
rect 406 207 407 208
rect 405 207 406 208
rect 353 207 354 208
rect 352 207 353 208
rect 351 207 352 208
rect 350 207 351 208
rect 349 207 350 208
rect 348 207 349 208
rect 347 207 348 208
rect 346 207 347 208
rect 345 207 346 208
rect 344 207 345 208
rect 343 207 344 208
rect 342 207 343 208
rect 341 207 342 208
rect 340 207 341 208
rect 339 207 340 208
rect 338 207 339 208
rect 337 207 338 208
rect 336 207 337 208
rect 335 207 336 208
rect 334 207 335 208
rect 333 207 334 208
rect 332 207 333 208
rect 331 207 332 208
rect 330 207 331 208
rect 329 207 330 208
rect 328 207 329 208
rect 327 207 328 208
rect 326 207 327 208
rect 325 207 326 208
rect 324 207 325 208
rect 323 207 324 208
rect 322 207 323 208
rect 321 207 322 208
rect 320 207 321 208
rect 319 207 320 208
rect 318 207 319 208
rect 317 207 318 208
rect 316 207 317 208
rect 315 207 316 208
rect 314 207 315 208
rect 313 207 314 208
rect 312 207 313 208
rect 311 207 312 208
rect 310 207 311 208
rect 309 207 310 208
rect 308 207 309 208
rect 307 207 308 208
rect 306 207 307 208
rect 305 207 306 208
rect 304 207 305 208
rect 303 207 304 208
rect 302 207 303 208
rect 301 207 302 208
rect 300 207 301 208
rect 299 207 300 208
rect 298 207 299 208
rect 297 207 298 208
rect 296 207 297 208
rect 295 207 296 208
rect 294 207 295 208
rect 293 207 294 208
rect 292 207 293 208
rect 291 207 292 208
rect 290 207 291 208
rect 289 207 290 208
rect 288 207 289 208
rect 287 207 288 208
rect 286 207 287 208
rect 285 207 286 208
rect 284 207 285 208
rect 283 207 284 208
rect 282 207 283 208
rect 281 207 282 208
rect 280 207 281 208
rect 279 207 280 208
rect 278 207 279 208
rect 277 207 278 208
rect 276 207 277 208
rect 275 207 276 208
rect 274 207 275 208
rect 273 207 274 208
rect 272 207 273 208
rect 271 207 272 208
rect 270 207 271 208
rect 269 207 270 208
rect 268 207 269 208
rect 267 207 268 208
rect 266 207 267 208
rect 265 207 266 208
rect 264 207 265 208
rect 263 207 264 208
rect 262 207 263 208
rect 261 207 262 208
rect 260 207 261 208
rect 259 207 260 208
rect 258 207 259 208
rect 257 207 258 208
rect 256 207 257 208
rect 255 207 256 208
rect 254 207 255 208
rect 253 207 254 208
rect 252 207 253 208
rect 251 207 252 208
rect 250 207 251 208
rect 249 207 250 208
rect 248 207 249 208
rect 247 207 248 208
rect 246 207 247 208
rect 245 207 246 208
rect 244 207 245 208
rect 243 207 244 208
rect 242 207 243 208
rect 241 207 242 208
rect 240 207 241 208
rect 239 207 240 208
rect 238 207 239 208
rect 237 207 238 208
rect 236 207 237 208
rect 235 207 236 208
rect 234 207 235 208
rect 233 207 234 208
rect 232 207 233 208
rect 231 207 232 208
rect 230 207 231 208
rect 229 207 230 208
rect 228 207 229 208
rect 227 207 228 208
rect 226 207 227 208
rect 225 207 226 208
rect 224 207 225 208
rect 223 207 224 208
rect 222 207 223 208
rect 221 207 222 208
rect 220 207 221 208
rect 219 207 220 208
rect 218 207 219 208
rect 217 207 218 208
rect 216 207 217 208
rect 215 207 216 208
rect 214 207 215 208
rect 213 207 214 208
rect 212 207 213 208
rect 211 207 212 208
rect 210 207 211 208
rect 209 207 210 208
rect 208 207 209 208
rect 207 207 208 208
rect 206 207 207 208
rect 205 207 206 208
rect 204 207 205 208
rect 203 207 204 208
rect 202 207 203 208
rect 201 207 202 208
rect 200 207 201 208
rect 199 207 200 208
rect 198 207 199 208
rect 197 207 198 208
rect 163 207 164 208
rect 162 207 163 208
rect 161 207 162 208
rect 160 207 161 208
rect 159 207 160 208
rect 158 207 159 208
rect 157 207 158 208
rect 156 207 157 208
rect 155 207 156 208
rect 154 207 155 208
rect 153 207 154 208
rect 152 207 153 208
rect 151 207 152 208
rect 150 207 151 208
rect 149 207 150 208
rect 148 207 149 208
rect 147 207 148 208
rect 146 207 147 208
rect 145 207 146 208
rect 144 207 145 208
rect 143 207 144 208
rect 142 207 143 208
rect 141 207 142 208
rect 140 207 141 208
rect 139 207 140 208
rect 138 207 139 208
rect 137 207 138 208
rect 136 207 137 208
rect 135 207 136 208
rect 134 207 135 208
rect 133 207 134 208
rect 132 207 133 208
rect 131 207 132 208
rect 130 207 131 208
rect 129 207 130 208
rect 128 207 129 208
rect 127 207 128 208
rect 126 207 127 208
rect 125 207 126 208
rect 124 207 125 208
rect 123 207 124 208
rect 122 207 123 208
rect 121 207 122 208
rect 120 207 121 208
rect 119 207 120 208
rect 118 207 119 208
rect 117 207 118 208
rect 116 207 117 208
rect 115 207 116 208
rect 114 207 115 208
rect 113 207 114 208
rect 112 207 113 208
rect 111 207 112 208
rect 110 207 111 208
rect 109 207 110 208
rect 108 207 109 208
rect 107 207 108 208
rect 106 207 107 208
rect 105 207 106 208
rect 104 207 105 208
rect 103 207 104 208
rect 102 207 103 208
rect 101 207 102 208
rect 100 207 101 208
rect 99 207 100 208
rect 98 207 99 208
rect 97 207 98 208
rect 96 207 97 208
rect 95 207 96 208
rect 94 207 95 208
rect 93 207 94 208
rect 92 207 93 208
rect 91 207 92 208
rect 90 207 91 208
rect 89 207 90 208
rect 88 207 89 208
rect 87 207 88 208
rect 86 207 87 208
rect 85 207 86 208
rect 84 207 85 208
rect 83 207 84 208
rect 82 207 83 208
rect 81 207 82 208
rect 80 207 81 208
rect 79 207 80 208
rect 59 207 60 208
rect 58 207 59 208
rect 57 207 58 208
rect 56 207 57 208
rect 55 207 56 208
rect 54 207 55 208
rect 53 207 54 208
rect 52 207 53 208
rect 51 207 52 208
rect 50 207 51 208
rect 49 207 50 208
rect 48 207 49 208
rect 47 207 48 208
rect 46 207 47 208
rect 45 207 46 208
rect 44 207 45 208
rect 43 207 44 208
rect 42 207 43 208
rect 41 207 42 208
rect 40 207 41 208
rect 39 207 40 208
rect 38 207 39 208
rect 37 207 38 208
rect 36 207 37 208
rect 35 207 36 208
rect 34 207 35 208
rect 33 207 34 208
rect 32 207 33 208
rect 31 207 32 208
rect 30 207 31 208
rect 29 207 30 208
rect 28 207 29 208
rect 27 207 28 208
rect 26 207 27 208
rect 25 207 26 208
rect 24 207 25 208
rect 23 207 24 208
rect 22 207 23 208
rect 21 207 22 208
rect 20 207 21 208
rect 19 207 20 208
rect 18 207 19 208
rect 17 207 18 208
rect 16 207 17 208
rect 15 207 16 208
rect 14 207 15 208
rect 13 207 14 208
rect 12 207 13 208
rect 11 207 12 208
rect 10 207 11 208
rect 9 207 10 208
rect 8 207 9 208
rect 7 207 8 208
rect 428 208 429 209
rect 427 208 428 209
rect 426 208 427 209
rect 425 208 426 209
rect 424 208 425 209
rect 423 208 424 209
rect 422 208 423 209
rect 421 208 422 209
rect 420 208 421 209
rect 419 208 420 209
rect 418 208 419 209
rect 417 208 418 209
rect 416 208 417 209
rect 415 208 416 209
rect 414 208 415 209
rect 413 208 414 209
rect 412 208 413 209
rect 411 208 412 209
rect 410 208 411 209
rect 409 208 410 209
rect 408 208 409 209
rect 407 208 408 209
rect 406 208 407 209
rect 405 208 406 209
rect 404 208 405 209
rect 403 208 404 209
rect 354 208 355 209
rect 353 208 354 209
rect 352 208 353 209
rect 351 208 352 209
rect 350 208 351 209
rect 349 208 350 209
rect 348 208 349 209
rect 347 208 348 209
rect 346 208 347 209
rect 345 208 346 209
rect 344 208 345 209
rect 343 208 344 209
rect 342 208 343 209
rect 341 208 342 209
rect 340 208 341 209
rect 339 208 340 209
rect 338 208 339 209
rect 337 208 338 209
rect 336 208 337 209
rect 335 208 336 209
rect 334 208 335 209
rect 333 208 334 209
rect 332 208 333 209
rect 331 208 332 209
rect 330 208 331 209
rect 329 208 330 209
rect 328 208 329 209
rect 327 208 328 209
rect 326 208 327 209
rect 325 208 326 209
rect 324 208 325 209
rect 323 208 324 209
rect 322 208 323 209
rect 321 208 322 209
rect 320 208 321 209
rect 319 208 320 209
rect 318 208 319 209
rect 317 208 318 209
rect 316 208 317 209
rect 315 208 316 209
rect 314 208 315 209
rect 313 208 314 209
rect 312 208 313 209
rect 311 208 312 209
rect 310 208 311 209
rect 309 208 310 209
rect 308 208 309 209
rect 307 208 308 209
rect 306 208 307 209
rect 305 208 306 209
rect 304 208 305 209
rect 303 208 304 209
rect 302 208 303 209
rect 301 208 302 209
rect 300 208 301 209
rect 299 208 300 209
rect 298 208 299 209
rect 297 208 298 209
rect 296 208 297 209
rect 295 208 296 209
rect 294 208 295 209
rect 293 208 294 209
rect 292 208 293 209
rect 291 208 292 209
rect 290 208 291 209
rect 289 208 290 209
rect 288 208 289 209
rect 287 208 288 209
rect 286 208 287 209
rect 285 208 286 209
rect 284 208 285 209
rect 283 208 284 209
rect 282 208 283 209
rect 281 208 282 209
rect 280 208 281 209
rect 279 208 280 209
rect 278 208 279 209
rect 277 208 278 209
rect 276 208 277 209
rect 275 208 276 209
rect 274 208 275 209
rect 273 208 274 209
rect 272 208 273 209
rect 271 208 272 209
rect 270 208 271 209
rect 269 208 270 209
rect 268 208 269 209
rect 267 208 268 209
rect 266 208 267 209
rect 265 208 266 209
rect 264 208 265 209
rect 263 208 264 209
rect 262 208 263 209
rect 261 208 262 209
rect 260 208 261 209
rect 259 208 260 209
rect 258 208 259 209
rect 257 208 258 209
rect 256 208 257 209
rect 255 208 256 209
rect 254 208 255 209
rect 253 208 254 209
rect 252 208 253 209
rect 251 208 252 209
rect 250 208 251 209
rect 249 208 250 209
rect 248 208 249 209
rect 247 208 248 209
rect 246 208 247 209
rect 245 208 246 209
rect 244 208 245 209
rect 243 208 244 209
rect 242 208 243 209
rect 241 208 242 209
rect 240 208 241 209
rect 239 208 240 209
rect 238 208 239 209
rect 237 208 238 209
rect 236 208 237 209
rect 235 208 236 209
rect 234 208 235 209
rect 233 208 234 209
rect 232 208 233 209
rect 231 208 232 209
rect 230 208 231 209
rect 229 208 230 209
rect 228 208 229 209
rect 227 208 228 209
rect 226 208 227 209
rect 225 208 226 209
rect 224 208 225 209
rect 223 208 224 209
rect 222 208 223 209
rect 221 208 222 209
rect 220 208 221 209
rect 219 208 220 209
rect 218 208 219 209
rect 217 208 218 209
rect 216 208 217 209
rect 215 208 216 209
rect 214 208 215 209
rect 213 208 214 209
rect 212 208 213 209
rect 211 208 212 209
rect 210 208 211 209
rect 209 208 210 209
rect 208 208 209 209
rect 207 208 208 209
rect 206 208 207 209
rect 205 208 206 209
rect 204 208 205 209
rect 203 208 204 209
rect 202 208 203 209
rect 201 208 202 209
rect 200 208 201 209
rect 199 208 200 209
rect 198 208 199 209
rect 197 208 198 209
rect 196 208 197 209
rect 160 208 161 209
rect 159 208 160 209
rect 158 208 159 209
rect 157 208 158 209
rect 156 208 157 209
rect 155 208 156 209
rect 154 208 155 209
rect 153 208 154 209
rect 152 208 153 209
rect 151 208 152 209
rect 150 208 151 209
rect 149 208 150 209
rect 148 208 149 209
rect 147 208 148 209
rect 146 208 147 209
rect 145 208 146 209
rect 144 208 145 209
rect 143 208 144 209
rect 142 208 143 209
rect 141 208 142 209
rect 140 208 141 209
rect 139 208 140 209
rect 138 208 139 209
rect 137 208 138 209
rect 136 208 137 209
rect 135 208 136 209
rect 134 208 135 209
rect 133 208 134 209
rect 132 208 133 209
rect 131 208 132 209
rect 130 208 131 209
rect 129 208 130 209
rect 128 208 129 209
rect 127 208 128 209
rect 126 208 127 209
rect 125 208 126 209
rect 124 208 125 209
rect 123 208 124 209
rect 122 208 123 209
rect 121 208 122 209
rect 120 208 121 209
rect 119 208 120 209
rect 118 208 119 209
rect 117 208 118 209
rect 116 208 117 209
rect 115 208 116 209
rect 114 208 115 209
rect 113 208 114 209
rect 112 208 113 209
rect 111 208 112 209
rect 110 208 111 209
rect 109 208 110 209
rect 108 208 109 209
rect 107 208 108 209
rect 106 208 107 209
rect 105 208 106 209
rect 104 208 105 209
rect 103 208 104 209
rect 102 208 103 209
rect 101 208 102 209
rect 100 208 101 209
rect 99 208 100 209
rect 98 208 99 209
rect 97 208 98 209
rect 96 208 97 209
rect 95 208 96 209
rect 94 208 95 209
rect 93 208 94 209
rect 92 208 93 209
rect 91 208 92 209
rect 90 208 91 209
rect 89 208 90 209
rect 88 208 89 209
rect 87 208 88 209
rect 86 208 87 209
rect 85 208 86 209
rect 84 208 85 209
rect 83 208 84 209
rect 82 208 83 209
rect 81 208 82 209
rect 80 208 81 209
rect 59 208 60 209
rect 58 208 59 209
rect 57 208 58 209
rect 56 208 57 209
rect 55 208 56 209
rect 54 208 55 209
rect 53 208 54 209
rect 52 208 53 209
rect 51 208 52 209
rect 50 208 51 209
rect 49 208 50 209
rect 48 208 49 209
rect 47 208 48 209
rect 46 208 47 209
rect 45 208 46 209
rect 44 208 45 209
rect 43 208 44 209
rect 42 208 43 209
rect 41 208 42 209
rect 40 208 41 209
rect 39 208 40 209
rect 38 208 39 209
rect 37 208 38 209
rect 36 208 37 209
rect 35 208 36 209
rect 34 208 35 209
rect 33 208 34 209
rect 32 208 33 209
rect 31 208 32 209
rect 30 208 31 209
rect 29 208 30 209
rect 28 208 29 209
rect 27 208 28 209
rect 26 208 27 209
rect 25 208 26 209
rect 24 208 25 209
rect 23 208 24 209
rect 22 208 23 209
rect 21 208 22 209
rect 20 208 21 209
rect 19 208 20 209
rect 18 208 19 209
rect 17 208 18 209
rect 16 208 17 209
rect 15 208 16 209
rect 14 208 15 209
rect 13 208 14 209
rect 12 208 13 209
rect 11 208 12 209
rect 10 208 11 209
rect 9 208 10 209
rect 8 208 9 209
rect 7 208 8 209
rect 429 209 430 210
rect 428 209 429 210
rect 427 209 428 210
rect 426 209 427 210
rect 425 209 426 210
rect 424 209 425 210
rect 423 209 424 210
rect 422 209 423 210
rect 421 209 422 210
rect 420 209 421 210
rect 419 209 420 210
rect 418 209 419 210
rect 417 209 418 210
rect 416 209 417 210
rect 415 209 416 210
rect 414 209 415 210
rect 413 209 414 210
rect 412 209 413 210
rect 411 209 412 210
rect 410 209 411 210
rect 409 209 410 210
rect 408 209 409 210
rect 407 209 408 210
rect 406 209 407 210
rect 405 209 406 210
rect 404 209 405 210
rect 403 209 404 210
rect 402 209 403 210
rect 354 209 355 210
rect 353 209 354 210
rect 352 209 353 210
rect 351 209 352 210
rect 350 209 351 210
rect 349 209 350 210
rect 348 209 349 210
rect 347 209 348 210
rect 346 209 347 210
rect 345 209 346 210
rect 344 209 345 210
rect 343 209 344 210
rect 342 209 343 210
rect 341 209 342 210
rect 340 209 341 210
rect 339 209 340 210
rect 338 209 339 210
rect 337 209 338 210
rect 336 209 337 210
rect 335 209 336 210
rect 334 209 335 210
rect 333 209 334 210
rect 332 209 333 210
rect 331 209 332 210
rect 330 209 331 210
rect 329 209 330 210
rect 328 209 329 210
rect 327 209 328 210
rect 326 209 327 210
rect 325 209 326 210
rect 324 209 325 210
rect 323 209 324 210
rect 322 209 323 210
rect 321 209 322 210
rect 320 209 321 210
rect 319 209 320 210
rect 318 209 319 210
rect 317 209 318 210
rect 316 209 317 210
rect 315 209 316 210
rect 314 209 315 210
rect 313 209 314 210
rect 312 209 313 210
rect 311 209 312 210
rect 310 209 311 210
rect 309 209 310 210
rect 308 209 309 210
rect 307 209 308 210
rect 306 209 307 210
rect 305 209 306 210
rect 304 209 305 210
rect 303 209 304 210
rect 302 209 303 210
rect 301 209 302 210
rect 300 209 301 210
rect 299 209 300 210
rect 298 209 299 210
rect 297 209 298 210
rect 296 209 297 210
rect 295 209 296 210
rect 294 209 295 210
rect 293 209 294 210
rect 292 209 293 210
rect 291 209 292 210
rect 290 209 291 210
rect 289 209 290 210
rect 288 209 289 210
rect 287 209 288 210
rect 286 209 287 210
rect 285 209 286 210
rect 284 209 285 210
rect 283 209 284 210
rect 282 209 283 210
rect 281 209 282 210
rect 280 209 281 210
rect 279 209 280 210
rect 278 209 279 210
rect 277 209 278 210
rect 276 209 277 210
rect 275 209 276 210
rect 274 209 275 210
rect 273 209 274 210
rect 272 209 273 210
rect 271 209 272 210
rect 270 209 271 210
rect 269 209 270 210
rect 268 209 269 210
rect 267 209 268 210
rect 266 209 267 210
rect 265 209 266 210
rect 264 209 265 210
rect 263 209 264 210
rect 262 209 263 210
rect 261 209 262 210
rect 260 209 261 210
rect 259 209 260 210
rect 258 209 259 210
rect 257 209 258 210
rect 256 209 257 210
rect 255 209 256 210
rect 254 209 255 210
rect 253 209 254 210
rect 252 209 253 210
rect 251 209 252 210
rect 250 209 251 210
rect 249 209 250 210
rect 248 209 249 210
rect 247 209 248 210
rect 246 209 247 210
rect 245 209 246 210
rect 244 209 245 210
rect 243 209 244 210
rect 242 209 243 210
rect 241 209 242 210
rect 240 209 241 210
rect 239 209 240 210
rect 238 209 239 210
rect 237 209 238 210
rect 236 209 237 210
rect 235 209 236 210
rect 234 209 235 210
rect 233 209 234 210
rect 232 209 233 210
rect 231 209 232 210
rect 230 209 231 210
rect 229 209 230 210
rect 228 209 229 210
rect 227 209 228 210
rect 226 209 227 210
rect 225 209 226 210
rect 224 209 225 210
rect 223 209 224 210
rect 222 209 223 210
rect 221 209 222 210
rect 220 209 221 210
rect 219 209 220 210
rect 218 209 219 210
rect 217 209 218 210
rect 216 209 217 210
rect 215 209 216 210
rect 214 209 215 210
rect 213 209 214 210
rect 212 209 213 210
rect 211 209 212 210
rect 210 209 211 210
rect 209 209 210 210
rect 208 209 209 210
rect 207 209 208 210
rect 206 209 207 210
rect 205 209 206 210
rect 204 209 205 210
rect 203 209 204 210
rect 202 209 203 210
rect 201 209 202 210
rect 200 209 201 210
rect 199 209 200 210
rect 198 209 199 210
rect 197 209 198 210
rect 196 209 197 210
rect 195 209 196 210
rect 194 209 195 210
rect 157 209 158 210
rect 156 209 157 210
rect 155 209 156 210
rect 154 209 155 210
rect 153 209 154 210
rect 152 209 153 210
rect 151 209 152 210
rect 150 209 151 210
rect 149 209 150 210
rect 148 209 149 210
rect 147 209 148 210
rect 146 209 147 210
rect 145 209 146 210
rect 144 209 145 210
rect 143 209 144 210
rect 142 209 143 210
rect 141 209 142 210
rect 140 209 141 210
rect 139 209 140 210
rect 138 209 139 210
rect 137 209 138 210
rect 136 209 137 210
rect 135 209 136 210
rect 134 209 135 210
rect 133 209 134 210
rect 132 209 133 210
rect 131 209 132 210
rect 130 209 131 210
rect 129 209 130 210
rect 128 209 129 210
rect 127 209 128 210
rect 126 209 127 210
rect 125 209 126 210
rect 124 209 125 210
rect 123 209 124 210
rect 122 209 123 210
rect 121 209 122 210
rect 120 209 121 210
rect 119 209 120 210
rect 118 209 119 210
rect 117 209 118 210
rect 116 209 117 210
rect 115 209 116 210
rect 114 209 115 210
rect 113 209 114 210
rect 112 209 113 210
rect 111 209 112 210
rect 110 209 111 210
rect 109 209 110 210
rect 108 209 109 210
rect 107 209 108 210
rect 106 209 107 210
rect 105 209 106 210
rect 104 209 105 210
rect 103 209 104 210
rect 102 209 103 210
rect 101 209 102 210
rect 100 209 101 210
rect 99 209 100 210
rect 98 209 99 210
rect 97 209 98 210
rect 96 209 97 210
rect 95 209 96 210
rect 94 209 95 210
rect 93 209 94 210
rect 92 209 93 210
rect 91 209 92 210
rect 90 209 91 210
rect 89 209 90 210
rect 88 209 89 210
rect 87 209 88 210
rect 86 209 87 210
rect 85 209 86 210
rect 84 209 85 210
rect 83 209 84 210
rect 82 209 83 210
rect 60 209 61 210
rect 59 209 60 210
rect 58 209 59 210
rect 57 209 58 210
rect 56 209 57 210
rect 55 209 56 210
rect 54 209 55 210
rect 53 209 54 210
rect 52 209 53 210
rect 51 209 52 210
rect 50 209 51 210
rect 49 209 50 210
rect 48 209 49 210
rect 47 209 48 210
rect 46 209 47 210
rect 45 209 46 210
rect 44 209 45 210
rect 43 209 44 210
rect 42 209 43 210
rect 41 209 42 210
rect 40 209 41 210
rect 39 209 40 210
rect 38 209 39 210
rect 37 209 38 210
rect 36 209 37 210
rect 35 209 36 210
rect 34 209 35 210
rect 33 209 34 210
rect 32 209 33 210
rect 31 209 32 210
rect 30 209 31 210
rect 29 209 30 210
rect 28 209 29 210
rect 27 209 28 210
rect 26 209 27 210
rect 25 209 26 210
rect 24 209 25 210
rect 23 209 24 210
rect 22 209 23 210
rect 21 209 22 210
rect 20 209 21 210
rect 19 209 20 210
rect 18 209 19 210
rect 17 209 18 210
rect 16 209 17 210
rect 15 209 16 210
rect 14 209 15 210
rect 13 209 14 210
rect 12 209 13 210
rect 11 209 12 210
rect 10 209 11 210
rect 9 209 10 210
rect 8 209 9 210
rect 7 209 8 210
rect 430 210 431 211
rect 429 210 430 211
rect 428 210 429 211
rect 427 210 428 211
rect 426 210 427 211
rect 425 210 426 211
rect 424 210 425 211
rect 423 210 424 211
rect 422 210 423 211
rect 421 210 422 211
rect 420 210 421 211
rect 419 210 420 211
rect 418 210 419 211
rect 417 210 418 211
rect 416 210 417 211
rect 415 210 416 211
rect 414 210 415 211
rect 413 210 414 211
rect 412 210 413 211
rect 411 210 412 211
rect 410 210 411 211
rect 409 210 410 211
rect 408 210 409 211
rect 407 210 408 211
rect 406 210 407 211
rect 405 210 406 211
rect 404 210 405 211
rect 403 210 404 211
rect 402 210 403 211
rect 401 210 402 211
rect 355 210 356 211
rect 354 210 355 211
rect 353 210 354 211
rect 352 210 353 211
rect 351 210 352 211
rect 350 210 351 211
rect 349 210 350 211
rect 348 210 349 211
rect 347 210 348 211
rect 346 210 347 211
rect 345 210 346 211
rect 344 210 345 211
rect 343 210 344 211
rect 342 210 343 211
rect 341 210 342 211
rect 340 210 341 211
rect 339 210 340 211
rect 338 210 339 211
rect 337 210 338 211
rect 336 210 337 211
rect 335 210 336 211
rect 334 210 335 211
rect 333 210 334 211
rect 332 210 333 211
rect 331 210 332 211
rect 330 210 331 211
rect 329 210 330 211
rect 328 210 329 211
rect 327 210 328 211
rect 326 210 327 211
rect 325 210 326 211
rect 324 210 325 211
rect 323 210 324 211
rect 322 210 323 211
rect 321 210 322 211
rect 320 210 321 211
rect 319 210 320 211
rect 318 210 319 211
rect 317 210 318 211
rect 316 210 317 211
rect 315 210 316 211
rect 314 210 315 211
rect 313 210 314 211
rect 312 210 313 211
rect 311 210 312 211
rect 310 210 311 211
rect 309 210 310 211
rect 308 210 309 211
rect 307 210 308 211
rect 306 210 307 211
rect 305 210 306 211
rect 304 210 305 211
rect 303 210 304 211
rect 302 210 303 211
rect 301 210 302 211
rect 300 210 301 211
rect 299 210 300 211
rect 298 210 299 211
rect 297 210 298 211
rect 296 210 297 211
rect 295 210 296 211
rect 294 210 295 211
rect 293 210 294 211
rect 292 210 293 211
rect 291 210 292 211
rect 290 210 291 211
rect 289 210 290 211
rect 288 210 289 211
rect 287 210 288 211
rect 286 210 287 211
rect 285 210 286 211
rect 284 210 285 211
rect 283 210 284 211
rect 282 210 283 211
rect 281 210 282 211
rect 280 210 281 211
rect 279 210 280 211
rect 278 210 279 211
rect 277 210 278 211
rect 276 210 277 211
rect 275 210 276 211
rect 274 210 275 211
rect 273 210 274 211
rect 272 210 273 211
rect 271 210 272 211
rect 270 210 271 211
rect 269 210 270 211
rect 268 210 269 211
rect 267 210 268 211
rect 266 210 267 211
rect 265 210 266 211
rect 264 210 265 211
rect 263 210 264 211
rect 262 210 263 211
rect 261 210 262 211
rect 260 210 261 211
rect 259 210 260 211
rect 258 210 259 211
rect 257 210 258 211
rect 256 210 257 211
rect 255 210 256 211
rect 254 210 255 211
rect 253 210 254 211
rect 252 210 253 211
rect 251 210 252 211
rect 250 210 251 211
rect 249 210 250 211
rect 248 210 249 211
rect 247 210 248 211
rect 246 210 247 211
rect 245 210 246 211
rect 244 210 245 211
rect 243 210 244 211
rect 242 210 243 211
rect 241 210 242 211
rect 240 210 241 211
rect 239 210 240 211
rect 238 210 239 211
rect 237 210 238 211
rect 236 210 237 211
rect 235 210 236 211
rect 234 210 235 211
rect 233 210 234 211
rect 232 210 233 211
rect 231 210 232 211
rect 230 210 231 211
rect 229 210 230 211
rect 228 210 229 211
rect 227 210 228 211
rect 226 210 227 211
rect 225 210 226 211
rect 224 210 225 211
rect 223 210 224 211
rect 222 210 223 211
rect 221 210 222 211
rect 220 210 221 211
rect 219 210 220 211
rect 218 210 219 211
rect 217 210 218 211
rect 216 210 217 211
rect 215 210 216 211
rect 214 210 215 211
rect 213 210 214 211
rect 212 210 213 211
rect 211 210 212 211
rect 210 210 211 211
rect 209 210 210 211
rect 208 210 209 211
rect 207 210 208 211
rect 206 210 207 211
rect 205 210 206 211
rect 204 210 205 211
rect 203 210 204 211
rect 202 210 203 211
rect 201 210 202 211
rect 200 210 201 211
rect 199 210 200 211
rect 198 210 199 211
rect 197 210 198 211
rect 196 210 197 211
rect 195 210 196 211
rect 194 210 195 211
rect 193 210 194 211
rect 154 210 155 211
rect 153 210 154 211
rect 152 210 153 211
rect 151 210 152 211
rect 150 210 151 211
rect 149 210 150 211
rect 148 210 149 211
rect 147 210 148 211
rect 146 210 147 211
rect 145 210 146 211
rect 144 210 145 211
rect 143 210 144 211
rect 142 210 143 211
rect 141 210 142 211
rect 140 210 141 211
rect 139 210 140 211
rect 138 210 139 211
rect 137 210 138 211
rect 136 210 137 211
rect 135 210 136 211
rect 134 210 135 211
rect 133 210 134 211
rect 132 210 133 211
rect 131 210 132 211
rect 130 210 131 211
rect 129 210 130 211
rect 128 210 129 211
rect 127 210 128 211
rect 126 210 127 211
rect 125 210 126 211
rect 124 210 125 211
rect 123 210 124 211
rect 122 210 123 211
rect 121 210 122 211
rect 120 210 121 211
rect 119 210 120 211
rect 118 210 119 211
rect 117 210 118 211
rect 116 210 117 211
rect 115 210 116 211
rect 114 210 115 211
rect 113 210 114 211
rect 112 210 113 211
rect 111 210 112 211
rect 110 210 111 211
rect 109 210 110 211
rect 108 210 109 211
rect 107 210 108 211
rect 106 210 107 211
rect 105 210 106 211
rect 104 210 105 211
rect 103 210 104 211
rect 102 210 103 211
rect 101 210 102 211
rect 100 210 101 211
rect 99 210 100 211
rect 98 210 99 211
rect 97 210 98 211
rect 96 210 97 211
rect 95 210 96 211
rect 94 210 95 211
rect 93 210 94 211
rect 92 210 93 211
rect 91 210 92 211
rect 90 210 91 211
rect 89 210 90 211
rect 88 210 89 211
rect 87 210 88 211
rect 86 210 87 211
rect 85 210 86 211
rect 84 210 85 211
rect 61 210 62 211
rect 60 210 61 211
rect 59 210 60 211
rect 58 210 59 211
rect 57 210 58 211
rect 56 210 57 211
rect 55 210 56 211
rect 54 210 55 211
rect 53 210 54 211
rect 52 210 53 211
rect 51 210 52 211
rect 50 210 51 211
rect 49 210 50 211
rect 48 210 49 211
rect 47 210 48 211
rect 46 210 47 211
rect 45 210 46 211
rect 44 210 45 211
rect 43 210 44 211
rect 42 210 43 211
rect 41 210 42 211
rect 40 210 41 211
rect 39 210 40 211
rect 38 210 39 211
rect 37 210 38 211
rect 36 210 37 211
rect 35 210 36 211
rect 34 210 35 211
rect 33 210 34 211
rect 32 210 33 211
rect 31 210 32 211
rect 30 210 31 211
rect 29 210 30 211
rect 28 210 29 211
rect 27 210 28 211
rect 26 210 27 211
rect 25 210 26 211
rect 24 210 25 211
rect 23 210 24 211
rect 22 210 23 211
rect 21 210 22 211
rect 20 210 21 211
rect 19 210 20 211
rect 18 210 19 211
rect 17 210 18 211
rect 16 210 17 211
rect 15 210 16 211
rect 14 210 15 211
rect 13 210 14 211
rect 12 210 13 211
rect 11 210 12 211
rect 10 210 11 211
rect 9 210 10 211
rect 8 210 9 211
rect 7 210 8 211
rect 431 211 432 212
rect 430 211 431 212
rect 429 211 430 212
rect 428 211 429 212
rect 427 211 428 212
rect 426 211 427 212
rect 425 211 426 212
rect 424 211 425 212
rect 423 211 424 212
rect 422 211 423 212
rect 421 211 422 212
rect 420 211 421 212
rect 419 211 420 212
rect 418 211 419 212
rect 417 211 418 212
rect 416 211 417 212
rect 415 211 416 212
rect 414 211 415 212
rect 413 211 414 212
rect 412 211 413 212
rect 411 211 412 212
rect 410 211 411 212
rect 409 211 410 212
rect 408 211 409 212
rect 407 211 408 212
rect 406 211 407 212
rect 405 211 406 212
rect 404 211 405 212
rect 403 211 404 212
rect 402 211 403 212
rect 401 211 402 212
rect 400 211 401 212
rect 356 211 357 212
rect 355 211 356 212
rect 354 211 355 212
rect 353 211 354 212
rect 352 211 353 212
rect 351 211 352 212
rect 350 211 351 212
rect 349 211 350 212
rect 348 211 349 212
rect 347 211 348 212
rect 346 211 347 212
rect 345 211 346 212
rect 344 211 345 212
rect 343 211 344 212
rect 342 211 343 212
rect 341 211 342 212
rect 340 211 341 212
rect 339 211 340 212
rect 338 211 339 212
rect 337 211 338 212
rect 336 211 337 212
rect 335 211 336 212
rect 334 211 335 212
rect 333 211 334 212
rect 332 211 333 212
rect 331 211 332 212
rect 330 211 331 212
rect 329 211 330 212
rect 328 211 329 212
rect 327 211 328 212
rect 326 211 327 212
rect 325 211 326 212
rect 324 211 325 212
rect 323 211 324 212
rect 322 211 323 212
rect 321 211 322 212
rect 320 211 321 212
rect 319 211 320 212
rect 318 211 319 212
rect 317 211 318 212
rect 316 211 317 212
rect 315 211 316 212
rect 314 211 315 212
rect 313 211 314 212
rect 312 211 313 212
rect 311 211 312 212
rect 310 211 311 212
rect 309 211 310 212
rect 308 211 309 212
rect 307 211 308 212
rect 306 211 307 212
rect 305 211 306 212
rect 304 211 305 212
rect 303 211 304 212
rect 302 211 303 212
rect 301 211 302 212
rect 300 211 301 212
rect 299 211 300 212
rect 298 211 299 212
rect 297 211 298 212
rect 296 211 297 212
rect 295 211 296 212
rect 294 211 295 212
rect 293 211 294 212
rect 292 211 293 212
rect 291 211 292 212
rect 290 211 291 212
rect 289 211 290 212
rect 288 211 289 212
rect 287 211 288 212
rect 286 211 287 212
rect 285 211 286 212
rect 284 211 285 212
rect 283 211 284 212
rect 282 211 283 212
rect 281 211 282 212
rect 280 211 281 212
rect 279 211 280 212
rect 278 211 279 212
rect 277 211 278 212
rect 276 211 277 212
rect 275 211 276 212
rect 274 211 275 212
rect 273 211 274 212
rect 272 211 273 212
rect 271 211 272 212
rect 270 211 271 212
rect 269 211 270 212
rect 268 211 269 212
rect 267 211 268 212
rect 266 211 267 212
rect 265 211 266 212
rect 264 211 265 212
rect 263 211 264 212
rect 262 211 263 212
rect 261 211 262 212
rect 260 211 261 212
rect 259 211 260 212
rect 258 211 259 212
rect 257 211 258 212
rect 256 211 257 212
rect 255 211 256 212
rect 254 211 255 212
rect 253 211 254 212
rect 252 211 253 212
rect 251 211 252 212
rect 250 211 251 212
rect 249 211 250 212
rect 248 211 249 212
rect 247 211 248 212
rect 246 211 247 212
rect 245 211 246 212
rect 244 211 245 212
rect 243 211 244 212
rect 242 211 243 212
rect 241 211 242 212
rect 240 211 241 212
rect 239 211 240 212
rect 238 211 239 212
rect 237 211 238 212
rect 236 211 237 212
rect 235 211 236 212
rect 234 211 235 212
rect 233 211 234 212
rect 232 211 233 212
rect 231 211 232 212
rect 230 211 231 212
rect 229 211 230 212
rect 228 211 229 212
rect 227 211 228 212
rect 226 211 227 212
rect 225 211 226 212
rect 224 211 225 212
rect 223 211 224 212
rect 222 211 223 212
rect 221 211 222 212
rect 220 211 221 212
rect 219 211 220 212
rect 218 211 219 212
rect 217 211 218 212
rect 216 211 217 212
rect 215 211 216 212
rect 214 211 215 212
rect 213 211 214 212
rect 212 211 213 212
rect 211 211 212 212
rect 210 211 211 212
rect 209 211 210 212
rect 208 211 209 212
rect 207 211 208 212
rect 206 211 207 212
rect 205 211 206 212
rect 204 211 205 212
rect 203 211 204 212
rect 202 211 203 212
rect 201 211 202 212
rect 200 211 201 212
rect 199 211 200 212
rect 198 211 199 212
rect 197 211 198 212
rect 196 211 197 212
rect 195 211 196 212
rect 194 211 195 212
rect 193 211 194 212
rect 192 211 193 212
rect 191 211 192 212
rect 151 211 152 212
rect 150 211 151 212
rect 149 211 150 212
rect 148 211 149 212
rect 147 211 148 212
rect 146 211 147 212
rect 145 211 146 212
rect 144 211 145 212
rect 143 211 144 212
rect 142 211 143 212
rect 141 211 142 212
rect 140 211 141 212
rect 139 211 140 212
rect 138 211 139 212
rect 137 211 138 212
rect 136 211 137 212
rect 135 211 136 212
rect 134 211 135 212
rect 133 211 134 212
rect 132 211 133 212
rect 131 211 132 212
rect 130 211 131 212
rect 129 211 130 212
rect 128 211 129 212
rect 127 211 128 212
rect 126 211 127 212
rect 125 211 126 212
rect 124 211 125 212
rect 123 211 124 212
rect 122 211 123 212
rect 121 211 122 212
rect 120 211 121 212
rect 119 211 120 212
rect 118 211 119 212
rect 117 211 118 212
rect 116 211 117 212
rect 115 211 116 212
rect 114 211 115 212
rect 113 211 114 212
rect 112 211 113 212
rect 111 211 112 212
rect 110 211 111 212
rect 109 211 110 212
rect 108 211 109 212
rect 107 211 108 212
rect 106 211 107 212
rect 105 211 106 212
rect 104 211 105 212
rect 103 211 104 212
rect 102 211 103 212
rect 101 211 102 212
rect 100 211 101 212
rect 99 211 100 212
rect 98 211 99 212
rect 97 211 98 212
rect 96 211 97 212
rect 95 211 96 212
rect 94 211 95 212
rect 93 211 94 212
rect 92 211 93 212
rect 91 211 92 212
rect 90 211 91 212
rect 89 211 90 212
rect 88 211 89 212
rect 87 211 88 212
rect 86 211 87 212
rect 62 211 63 212
rect 61 211 62 212
rect 60 211 61 212
rect 59 211 60 212
rect 58 211 59 212
rect 57 211 58 212
rect 56 211 57 212
rect 55 211 56 212
rect 54 211 55 212
rect 53 211 54 212
rect 52 211 53 212
rect 51 211 52 212
rect 50 211 51 212
rect 49 211 50 212
rect 48 211 49 212
rect 47 211 48 212
rect 46 211 47 212
rect 45 211 46 212
rect 44 211 45 212
rect 43 211 44 212
rect 42 211 43 212
rect 41 211 42 212
rect 40 211 41 212
rect 39 211 40 212
rect 38 211 39 212
rect 37 211 38 212
rect 36 211 37 212
rect 35 211 36 212
rect 34 211 35 212
rect 33 211 34 212
rect 32 211 33 212
rect 31 211 32 212
rect 30 211 31 212
rect 29 211 30 212
rect 28 211 29 212
rect 27 211 28 212
rect 26 211 27 212
rect 25 211 26 212
rect 24 211 25 212
rect 23 211 24 212
rect 22 211 23 212
rect 21 211 22 212
rect 20 211 21 212
rect 19 211 20 212
rect 18 211 19 212
rect 17 211 18 212
rect 16 211 17 212
rect 15 211 16 212
rect 14 211 15 212
rect 13 211 14 212
rect 12 211 13 212
rect 11 211 12 212
rect 10 211 11 212
rect 9 211 10 212
rect 8 211 9 212
rect 7 211 8 212
rect 6 211 7 212
rect 432 212 433 213
rect 431 212 432 213
rect 430 212 431 213
rect 429 212 430 213
rect 428 212 429 213
rect 427 212 428 213
rect 426 212 427 213
rect 425 212 426 213
rect 424 212 425 213
rect 423 212 424 213
rect 422 212 423 213
rect 421 212 422 213
rect 420 212 421 213
rect 419 212 420 213
rect 418 212 419 213
rect 417 212 418 213
rect 416 212 417 213
rect 415 212 416 213
rect 414 212 415 213
rect 413 212 414 213
rect 412 212 413 213
rect 411 212 412 213
rect 410 212 411 213
rect 409 212 410 213
rect 408 212 409 213
rect 407 212 408 213
rect 406 212 407 213
rect 405 212 406 213
rect 404 212 405 213
rect 403 212 404 213
rect 402 212 403 213
rect 401 212 402 213
rect 400 212 401 213
rect 399 212 400 213
rect 356 212 357 213
rect 355 212 356 213
rect 354 212 355 213
rect 353 212 354 213
rect 352 212 353 213
rect 351 212 352 213
rect 350 212 351 213
rect 349 212 350 213
rect 348 212 349 213
rect 347 212 348 213
rect 346 212 347 213
rect 345 212 346 213
rect 344 212 345 213
rect 343 212 344 213
rect 342 212 343 213
rect 341 212 342 213
rect 340 212 341 213
rect 339 212 340 213
rect 338 212 339 213
rect 337 212 338 213
rect 336 212 337 213
rect 335 212 336 213
rect 334 212 335 213
rect 333 212 334 213
rect 332 212 333 213
rect 331 212 332 213
rect 330 212 331 213
rect 329 212 330 213
rect 328 212 329 213
rect 327 212 328 213
rect 326 212 327 213
rect 325 212 326 213
rect 324 212 325 213
rect 323 212 324 213
rect 322 212 323 213
rect 321 212 322 213
rect 320 212 321 213
rect 319 212 320 213
rect 318 212 319 213
rect 317 212 318 213
rect 316 212 317 213
rect 315 212 316 213
rect 314 212 315 213
rect 313 212 314 213
rect 312 212 313 213
rect 311 212 312 213
rect 310 212 311 213
rect 309 212 310 213
rect 308 212 309 213
rect 307 212 308 213
rect 306 212 307 213
rect 305 212 306 213
rect 304 212 305 213
rect 303 212 304 213
rect 302 212 303 213
rect 301 212 302 213
rect 300 212 301 213
rect 299 212 300 213
rect 298 212 299 213
rect 297 212 298 213
rect 296 212 297 213
rect 295 212 296 213
rect 294 212 295 213
rect 293 212 294 213
rect 292 212 293 213
rect 291 212 292 213
rect 290 212 291 213
rect 289 212 290 213
rect 288 212 289 213
rect 287 212 288 213
rect 286 212 287 213
rect 285 212 286 213
rect 284 212 285 213
rect 283 212 284 213
rect 282 212 283 213
rect 281 212 282 213
rect 280 212 281 213
rect 279 212 280 213
rect 278 212 279 213
rect 277 212 278 213
rect 276 212 277 213
rect 275 212 276 213
rect 274 212 275 213
rect 273 212 274 213
rect 272 212 273 213
rect 271 212 272 213
rect 270 212 271 213
rect 269 212 270 213
rect 268 212 269 213
rect 267 212 268 213
rect 266 212 267 213
rect 265 212 266 213
rect 264 212 265 213
rect 263 212 264 213
rect 262 212 263 213
rect 261 212 262 213
rect 260 212 261 213
rect 259 212 260 213
rect 258 212 259 213
rect 257 212 258 213
rect 256 212 257 213
rect 255 212 256 213
rect 254 212 255 213
rect 253 212 254 213
rect 252 212 253 213
rect 251 212 252 213
rect 250 212 251 213
rect 249 212 250 213
rect 248 212 249 213
rect 247 212 248 213
rect 246 212 247 213
rect 245 212 246 213
rect 244 212 245 213
rect 243 212 244 213
rect 242 212 243 213
rect 241 212 242 213
rect 240 212 241 213
rect 239 212 240 213
rect 238 212 239 213
rect 237 212 238 213
rect 236 212 237 213
rect 235 212 236 213
rect 234 212 235 213
rect 233 212 234 213
rect 232 212 233 213
rect 231 212 232 213
rect 230 212 231 213
rect 229 212 230 213
rect 228 212 229 213
rect 227 212 228 213
rect 226 212 227 213
rect 225 212 226 213
rect 224 212 225 213
rect 223 212 224 213
rect 222 212 223 213
rect 221 212 222 213
rect 220 212 221 213
rect 219 212 220 213
rect 218 212 219 213
rect 217 212 218 213
rect 216 212 217 213
rect 215 212 216 213
rect 214 212 215 213
rect 213 212 214 213
rect 212 212 213 213
rect 211 212 212 213
rect 210 212 211 213
rect 209 212 210 213
rect 208 212 209 213
rect 207 212 208 213
rect 206 212 207 213
rect 205 212 206 213
rect 204 212 205 213
rect 203 212 204 213
rect 202 212 203 213
rect 201 212 202 213
rect 200 212 201 213
rect 199 212 200 213
rect 198 212 199 213
rect 197 212 198 213
rect 196 212 197 213
rect 195 212 196 213
rect 194 212 195 213
rect 193 212 194 213
rect 192 212 193 213
rect 191 212 192 213
rect 190 212 191 213
rect 149 212 150 213
rect 148 212 149 213
rect 147 212 148 213
rect 146 212 147 213
rect 145 212 146 213
rect 144 212 145 213
rect 143 212 144 213
rect 142 212 143 213
rect 141 212 142 213
rect 140 212 141 213
rect 139 212 140 213
rect 138 212 139 213
rect 137 212 138 213
rect 136 212 137 213
rect 135 212 136 213
rect 134 212 135 213
rect 133 212 134 213
rect 132 212 133 213
rect 131 212 132 213
rect 130 212 131 213
rect 129 212 130 213
rect 128 212 129 213
rect 127 212 128 213
rect 126 212 127 213
rect 125 212 126 213
rect 124 212 125 213
rect 123 212 124 213
rect 122 212 123 213
rect 121 212 122 213
rect 120 212 121 213
rect 119 212 120 213
rect 118 212 119 213
rect 117 212 118 213
rect 116 212 117 213
rect 115 212 116 213
rect 114 212 115 213
rect 113 212 114 213
rect 112 212 113 213
rect 111 212 112 213
rect 110 212 111 213
rect 109 212 110 213
rect 108 212 109 213
rect 107 212 108 213
rect 106 212 107 213
rect 105 212 106 213
rect 104 212 105 213
rect 103 212 104 213
rect 102 212 103 213
rect 101 212 102 213
rect 100 212 101 213
rect 99 212 100 213
rect 98 212 99 213
rect 97 212 98 213
rect 96 212 97 213
rect 95 212 96 213
rect 94 212 95 213
rect 93 212 94 213
rect 92 212 93 213
rect 91 212 92 213
rect 90 212 91 213
rect 89 212 90 213
rect 88 212 89 213
rect 63 212 64 213
rect 62 212 63 213
rect 61 212 62 213
rect 60 212 61 213
rect 59 212 60 213
rect 58 212 59 213
rect 57 212 58 213
rect 56 212 57 213
rect 55 212 56 213
rect 54 212 55 213
rect 53 212 54 213
rect 52 212 53 213
rect 51 212 52 213
rect 50 212 51 213
rect 49 212 50 213
rect 48 212 49 213
rect 47 212 48 213
rect 46 212 47 213
rect 45 212 46 213
rect 44 212 45 213
rect 43 212 44 213
rect 42 212 43 213
rect 41 212 42 213
rect 40 212 41 213
rect 39 212 40 213
rect 38 212 39 213
rect 37 212 38 213
rect 36 212 37 213
rect 35 212 36 213
rect 34 212 35 213
rect 33 212 34 213
rect 32 212 33 213
rect 31 212 32 213
rect 30 212 31 213
rect 29 212 30 213
rect 28 212 29 213
rect 27 212 28 213
rect 26 212 27 213
rect 25 212 26 213
rect 24 212 25 213
rect 23 212 24 213
rect 22 212 23 213
rect 21 212 22 213
rect 20 212 21 213
rect 19 212 20 213
rect 18 212 19 213
rect 17 212 18 213
rect 16 212 17 213
rect 15 212 16 213
rect 14 212 15 213
rect 13 212 14 213
rect 12 212 13 213
rect 11 212 12 213
rect 10 212 11 213
rect 9 212 10 213
rect 8 212 9 213
rect 7 212 8 213
rect 6 212 7 213
rect 433 213 434 214
rect 432 213 433 214
rect 431 213 432 214
rect 430 213 431 214
rect 429 213 430 214
rect 428 213 429 214
rect 427 213 428 214
rect 426 213 427 214
rect 425 213 426 214
rect 424 213 425 214
rect 423 213 424 214
rect 422 213 423 214
rect 421 213 422 214
rect 420 213 421 214
rect 419 213 420 214
rect 418 213 419 214
rect 417 213 418 214
rect 416 213 417 214
rect 415 213 416 214
rect 414 213 415 214
rect 413 213 414 214
rect 412 213 413 214
rect 411 213 412 214
rect 410 213 411 214
rect 409 213 410 214
rect 408 213 409 214
rect 407 213 408 214
rect 406 213 407 214
rect 405 213 406 214
rect 404 213 405 214
rect 403 213 404 214
rect 402 213 403 214
rect 401 213 402 214
rect 400 213 401 214
rect 399 213 400 214
rect 398 213 399 214
rect 357 213 358 214
rect 356 213 357 214
rect 355 213 356 214
rect 354 213 355 214
rect 353 213 354 214
rect 352 213 353 214
rect 351 213 352 214
rect 350 213 351 214
rect 349 213 350 214
rect 348 213 349 214
rect 347 213 348 214
rect 346 213 347 214
rect 345 213 346 214
rect 344 213 345 214
rect 343 213 344 214
rect 342 213 343 214
rect 341 213 342 214
rect 340 213 341 214
rect 339 213 340 214
rect 338 213 339 214
rect 337 213 338 214
rect 336 213 337 214
rect 335 213 336 214
rect 334 213 335 214
rect 333 213 334 214
rect 332 213 333 214
rect 331 213 332 214
rect 330 213 331 214
rect 329 213 330 214
rect 309 213 310 214
rect 308 213 309 214
rect 307 213 308 214
rect 306 213 307 214
rect 305 213 306 214
rect 304 213 305 214
rect 303 213 304 214
rect 302 213 303 214
rect 301 213 302 214
rect 300 213 301 214
rect 299 213 300 214
rect 298 213 299 214
rect 297 213 298 214
rect 296 213 297 214
rect 295 213 296 214
rect 294 213 295 214
rect 293 213 294 214
rect 292 213 293 214
rect 291 213 292 214
rect 290 213 291 214
rect 289 213 290 214
rect 288 213 289 214
rect 287 213 288 214
rect 286 213 287 214
rect 285 213 286 214
rect 284 213 285 214
rect 283 213 284 214
rect 282 213 283 214
rect 281 213 282 214
rect 280 213 281 214
rect 279 213 280 214
rect 278 213 279 214
rect 277 213 278 214
rect 276 213 277 214
rect 275 213 276 214
rect 274 213 275 214
rect 273 213 274 214
rect 272 213 273 214
rect 271 213 272 214
rect 270 213 271 214
rect 269 213 270 214
rect 268 213 269 214
rect 267 213 268 214
rect 266 213 267 214
rect 265 213 266 214
rect 264 213 265 214
rect 263 213 264 214
rect 262 213 263 214
rect 261 213 262 214
rect 260 213 261 214
rect 259 213 260 214
rect 258 213 259 214
rect 257 213 258 214
rect 256 213 257 214
rect 255 213 256 214
rect 254 213 255 214
rect 253 213 254 214
rect 252 213 253 214
rect 251 213 252 214
rect 250 213 251 214
rect 249 213 250 214
rect 248 213 249 214
rect 247 213 248 214
rect 246 213 247 214
rect 245 213 246 214
rect 244 213 245 214
rect 243 213 244 214
rect 242 213 243 214
rect 241 213 242 214
rect 240 213 241 214
rect 239 213 240 214
rect 238 213 239 214
rect 237 213 238 214
rect 236 213 237 214
rect 235 213 236 214
rect 234 213 235 214
rect 233 213 234 214
rect 232 213 233 214
rect 231 213 232 214
rect 230 213 231 214
rect 229 213 230 214
rect 228 213 229 214
rect 227 213 228 214
rect 226 213 227 214
rect 225 213 226 214
rect 224 213 225 214
rect 223 213 224 214
rect 222 213 223 214
rect 221 213 222 214
rect 220 213 221 214
rect 219 213 220 214
rect 218 213 219 214
rect 217 213 218 214
rect 216 213 217 214
rect 215 213 216 214
rect 214 213 215 214
rect 213 213 214 214
rect 212 213 213 214
rect 211 213 212 214
rect 210 213 211 214
rect 209 213 210 214
rect 208 213 209 214
rect 207 213 208 214
rect 206 213 207 214
rect 205 213 206 214
rect 204 213 205 214
rect 203 213 204 214
rect 202 213 203 214
rect 201 213 202 214
rect 200 213 201 214
rect 199 213 200 214
rect 198 213 199 214
rect 197 213 198 214
rect 196 213 197 214
rect 195 213 196 214
rect 194 213 195 214
rect 193 213 194 214
rect 192 213 193 214
rect 191 213 192 214
rect 190 213 191 214
rect 189 213 190 214
rect 188 213 189 214
rect 147 213 148 214
rect 146 213 147 214
rect 145 213 146 214
rect 144 213 145 214
rect 143 213 144 214
rect 142 213 143 214
rect 141 213 142 214
rect 140 213 141 214
rect 139 213 140 214
rect 138 213 139 214
rect 137 213 138 214
rect 136 213 137 214
rect 135 213 136 214
rect 134 213 135 214
rect 133 213 134 214
rect 132 213 133 214
rect 131 213 132 214
rect 130 213 131 214
rect 129 213 130 214
rect 128 213 129 214
rect 127 213 128 214
rect 126 213 127 214
rect 125 213 126 214
rect 124 213 125 214
rect 123 213 124 214
rect 122 213 123 214
rect 121 213 122 214
rect 120 213 121 214
rect 119 213 120 214
rect 118 213 119 214
rect 117 213 118 214
rect 116 213 117 214
rect 115 213 116 214
rect 114 213 115 214
rect 113 213 114 214
rect 112 213 113 214
rect 111 213 112 214
rect 110 213 111 214
rect 109 213 110 214
rect 108 213 109 214
rect 107 213 108 214
rect 106 213 107 214
rect 105 213 106 214
rect 104 213 105 214
rect 103 213 104 214
rect 102 213 103 214
rect 101 213 102 214
rect 100 213 101 214
rect 99 213 100 214
rect 98 213 99 214
rect 97 213 98 214
rect 96 213 97 214
rect 95 213 96 214
rect 94 213 95 214
rect 93 213 94 214
rect 92 213 93 214
rect 91 213 92 214
rect 64 213 65 214
rect 63 213 64 214
rect 62 213 63 214
rect 61 213 62 214
rect 60 213 61 214
rect 59 213 60 214
rect 58 213 59 214
rect 57 213 58 214
rect 56 213 57 214
rect 55 213 56 214
rect 54 213 55 214
rect 53 213 54 214
rect 52 213 53 214
rect 51 213 52 214
rect 50 213 51 214
rect 49 213 50 214
rect 48 213 49 214
rect 47 213 48 214
rect 46 213 47 214
rect 45 213 46 214
rect 44 213 45 214
rect 43 213 44 214
rect 42 213 43 214
rect 41 213 42 214
rect 40 213 41 214
rect 39 213 40 214
rect 38 213 39 214
rect 37 213 38 214
rect 36 213 37 214
rect 35 213 36 214
rect 34 213 35 214
rect 33 213 34 214
rect 32 213 33 214
rect 31 213 32 214
rect 30 213 31 214
rect 29 213 30 214
rect 28 213 29 214
rect 27 213 28 214
rect 26 213 27 214
rect 25 213 26 214
rect 24 213 25 214
rect 23 213 24 214
rect 22 213 23 214
rect 21 213 22 214
rect 20 213 21 214
rect 19 213 20 214
rect 18 213 19 214
rect 17 213 18 214
rect 16 213 17 214
rect 15 213 16 214
rect 14 213 15 214
rect 13 213 14 214
rect 12 213 13 214
rect 11 213 12 214
rect 10 213 11 214
rect 9 213 10 214
rect 8 213 9 214
rect 7 213 8 214
rect 6 213 7 214
rect 478 214 479 215
rect 458 214 459 215
rect 434 214 435 215
rect 433 214 434 215
rect 432 214 433 215
rect 431 214 432 215
rect 430 214 431 215
rect 429 214 430 215
rect 428 214 429 215
rect 427 214 428 215
rect 426 214 427 215
rect 425 214 426 215
rect 424 214 425 215
rect 423 214 424 215
rect 422 214 423 215
rect 421 214 422 215
rect 420 214 421 215
rect 419 214 420 215
rect 418 214 419 215
rect 417 214 418 215
rect 416 214 417 215
rect 415 214 416 215
rect 414 214 415 215
rect 413 214 414 215
rect 412 214 413 215
rect 411 214 412 215
rect 410 214 411 215
rect 409 214 410 215
rect 408 214 409 215
rect 407 214 408 215
rect 406 214 407 215
rect 405 214 406 215
rect 404 214 405 215
rect 403 214 404 215
rect 402 214 403 215
rect 401 214 402 215
rect 400 214 401 215
rect 399 214 400 215
rect 398 214 399 215
rect 397 214 398 215
rect 357 214 358 215
rect 356 214 357 215
rect 355 214 356 215
rect 354 214 355 215
rect 353 214 354 215
rect 352 214 353 215
rect 351 214 352 215
rect 350 214 351 215
rect 349 214 350 215
rect 348 214 349 215
rect 347 214 348 215
rect 346 214 347 215
rect 345 214 346 215
rect 344 214 345 215
rect 343 214 344 215
rect 342 214 343 215
rect 341 214 342 215
rect 340 214 341 215
rect 339 214 340 215
rect 338 214 339 215
rect 337 214 338 215
rect 336 214 337 215
rect 335 214 336 215
rect 303 214 304 215
rect 302 214 303 215
rect 301 214 302 215
rect 300 214 301 215
rect 299 214 300 215
rect 298 214 299 215
rect 297 214 298 215
rect 296 214 297 215
rect 295 214 296 215
rect 294 214 295 215
rect 293 214 294 215
rect 292 214 293 215
rect 291 214 292 215
rect 290 214 291 215
rect 289 214 290 215
rect 288 214 289 215
rect 287 214 288 215
rect 286 214 287 215
rect 285 214 286 215
rect 284 214 285 215
rect 283 214 284 215
rect 282 214 283 215
rect 281 214 282 215
rect 280 214 281 215
rect 279 214 280 215
rect 278 214 279 215
rect 277 214 278 215
rect 276 214 277 215
rect 275 214 276 215
rect 274 214 275 215
rect 273 214 274 215
rect 272 214 273 215
rect 271 214 272 215
rect 270 214 271 215
rect 269 214 270 215
rect 268 214 269 215
rect 267 214 268 215
rect 266 214 267 215
rect 265 214 266 215
rect 264 214 265 215
rect 263 214 264 215
rect 262 214 263 215
rect 261 214 262 215
rect 260 214 261 215
rect 259 214 260 215
rect 258 214 259 215
rect 257 214 258 215
rect 256 214 257 215
rect 255 214 256 215
rect 254 214 255 215
rect 253 214 254 215
rect 252 214 253 215
rect 251 214 252 215
rect 250 214 251 215
rect 249 214 250 215
rect 248 214 249 215
rect 247 214 248 215
rect 246 214 247 215
rect 245 214 246 215
rect 244 214 245 215
rect 243 214 244 215
rect 242 214 243 215
rect 241 214 242 215
rect 240 214 241 215
rect 239 214 240 215
rect 238 214 239 215
rect 237 214 238 215
rect 236 214 237 215
rect 235 214 236 215
rect 234 214 235 215
rect 233 214 234 215
rect 232 214 233 215
rect 231 214 232 215
rect 230 214 231 215
rect 229 214 230 215
rect 228 214 229 215
rect 227 214 228 215
rect 226 214 227 215
rect 225 214 226 215
rect 224 214 225 215
rect 223 214 224 215
rect 222 214 223 215
rect 221 214 222 215
rect 220 214 221 215
rect 219 214 220 215
rect 218 214 219 215
rect 217 214 218 215
rect 216 214 217 215
rect 215 214 216 215
rect 214 214 215 215
rect 213 214 214 215
rect 212 214 213 215
rect 211 214 212 215
rect 210 214 211 215
rect 209 214 210 215
rect 208 214 209 215
rect 207 214 208 215
rect 206 214 207 215
rect 205 214 206 215
rect 204 214 205 215
rect 203 214 204 215
rect 202 214 203 215
rect 201 214 202 215
rect 200 214 201 215
rect 199 214 200 215
rect 198 214 199 215
rect 197 214 198 215
rect 196 214 197 215
rect 195 214 196 215
rect 194 214 195 215
rect 193 214 194 215
rect 192 214 193 215
rect 191 214 192 215
rect 190 214 191 215
rect 189 214 190 215
rect 188 214 189 215
rect 187 214 188 215
rect 186 214 187 215
rect 146 214 147 215
rect 145 214 146 215
rect 144 214 145 215
rect 143 214 144 215
rect 142 214 143 215
rect 141 214 142 215
rect 140 214 141 215
rect 139 214 140 215
rect 138 214 139 215
rect 137 214 138 215
rect 136 214 137 215
rect 135 214 136 215
rect 134 214 135 215
rect 133 214 134 215
rect 132 214 133 215
rect 131 214 132 215
rect 130 214 131 215
rect 129 214 130 215
rect 128 214 129 215
rect 127 214 128 215
rect 126 214 127 215
rect 125 214 126 215
rect 124 214 125 215
rect 123 214 124 215
rect 122 214 123 215
rect 121 214 122 215
rect 120 214 121 215
rect 119 214 120 215
rect 118 214 119 215
rect 117 214 118 215
rect 116 214 117 215
rect 115 214 116 215
rect 114 214 115 215
rect 113 214 114 215
rect 112 214 113 215
rect 111 214 112 215
rect 110 214 111 215
rect 109 214 110 215
rect 108 214 109 215
rect 107 214 108 215
rect 106 214 107 215
rect 105 214 106 215
rect 104 214 105 215
rect 103 214 104 215
rect 102 214 103 215
rect 101 214 102 215
rect 100 214 101 215
rect 99 214 100 215
rect 98 214 99 215
rect 97 214 98 215
rect 96 214 97 215
rect 95 214 96 215
rect 94 214 95 215
rect 93 214 94 215
rect 65 214 66 215
rect 64 214 65 215
rect 63 214 64 215
rect 62 214 63 215
rect 61 214 62 215
rect 60 214 61 215
rect 59 214 60 215
rect 58 214 59 215
rect 57 214 58 215
rect 56 214 57 215
rect 55 214 56 215
rect 54 214 55 215
rect 53 214 54 215
rect 52 214 53 215
rect 51 214 52 215
rect 50 214 51 215
rect 49 214 50 215
rect 48 214 49 215
rect 47 214 48 215
rect 46 214 47 215
rect 45 214 46 215
rect 44 214 45 215
rect 43 214 44 215
rect 42 214 43 215
rect 41 214 42 215
rect 40 214 41 215
rect 39 214 40 215
rect 38 214 39 215
rect 37 214 38 215
rect 36 214 37 215
rect 35 214 36 215
rect 34 214 35 215
rect 33 214 34 215
rect 32 214 33 215
rect 31 214 32 215
rect 30 214 31 215
rect 29 214 30 215
rect 28 214 29 215
rect 27 214 28 215
rect 26 214 27 215
rect 25 214 26 215
rect 24 214 25 215
rect 23 214 24 215
rect 22 214 23 215
rect 21 214 22 215
rect 20 214 21 215
rect 19 214 20 215
rect 18 214 19 215
rect 17 214 18 215
rect 16 214 17 215
rect 15 214 16 215
rect 14 214 15 215
rect 13 214 14 215
rect 12 214 13 215
rect 11 214 12 215
rect 10 214 11 215
rect 9 214 10 215
rect 8 214 9 215
rect 7 214 8 215
rect 6 214 7 215
rect 478 215 479 216
rect 458 215 459 216
rect 434 215 435 216
rect 433 215 434 216
rect 432 215 433 216
rect 431 215 432 216
rect 430 215 431 216
rect 429 215 430 216
rect 428 215 429 216
rect 427 215 428 216
rect 426 215 427 216
rect 425 215 426 216
rect 424 215 425 216
rect 423 215 424 216
rect 422 215 423 216
rect 421 215 422 216
rect 420 215 421 216
rect 419 215 420 216
rect 418 215 419 216
rect 417 215 418 216
rect 416 215 417 216
rect 415 215 416 216
rect 414 215 415 216
rect 413 215 414 216
rect 412 215 413 216
rect 411 215 412 216
rect 410 215 411 216
rect 409 215 410 216
rect 408 215 409 216
rect 407 215 408 216
rect 406 215 407 216
rect 405 215 406 216
rect 404 215 405 216
rect 403 215 404 216
rect 402 215 403 216
rect 401 215 402 216
rect 400 215 401 216
rect 399 215 400 216
rect 398 215 399 216
rect 397 215 398 216
rect 358 215 359 216
rect 357 215 358 216
rect 356 215 357 216
rect 355 215 356 216
rect 354 215 355 216
rect 353 215 354 216
rect 352 215 353 216
rect 351 215 352 216
rect 350 215 351 216
rect 349 215 350 216
rect 348 215 349 216
rect 347 215 348 216
rect 346 215 347 216
rect 345 215 346 216
rect 344 215 345 216
rect 343 215 344 216
rect 342 215 343 216
rect 341 215 342 216
rect 340 215 341 216
rect 299 215 300 216
rect 298 215 299 216
rect 297 215 298 216
rect 296 215 297 216
rect 295 215 296 216
rect 294 215 295 216
rect 293 215 294 216
rect 292 215 293 216
rect 291 215 292 216
rect 290 215 291 216
rect 289 215 290 216
rect 288 215 289 216
rect 287 215 288 216
rect 286 215 287 216
rect 285 215 286 216
rect 284 215 285 216
rect 283 215 284 216
rect 282 215 283 216
rect 281 215 282 216
rect 280 215 281 216
rect 279 215 280 216
rect 278 215 279 216
rect 277 215 278 216
rect 276 215 277 216
rect 275 215 276 216
rect 274 215 275 216
rect 273 215 274 216
rect 272 215 273 216
rect 271 215 272 216
rect 270 215 271 216
rect 269 215 270 216
rect 268 215 269 216
rect 267 215 268 216
rect 266 215 267 216
rect 265 215 266 216
rect 264 215 265 216
rect 263 215 264 216
rect 262 215 263 216
rect 261 215 262 216
rect 260 215 261 216
rect 259 215 260 216
rect 258 215 259 216
rect 257 215 258 216
rect 256 215 257 216
rect 255 215 256 216
rect 254 215 255 216
rect 253 215 254 216
rect 252 215 253 216
rect 251 215 252 216
rect 250 215 251 216
rect 249 215 250 216
rect 248 215 249 216
rect 247 215 248 216
rect 246 215 247 216
rect 245 215 246 216
rect 244 215 245 216
rect 243 215 244 216
rect 242 215 243 216
rect 241 215 242 216
rect 240 215 241 216
rect 239 215 240 216
rect 238 215 239 216
rect 237 215 238 216
rect 236 215 237 216
rect 235 215 236 216
rect 234 215 235 216
rect 233 215 234 216
rect 232 215 233 216
rect 231 215 232 216
rect 230 215 231 216
rect 229 215 230 216
rect 228 215 229 216
rect 227 215 228 216
rect 226 215 227 216
rect 225 215 226 216
rect 224 215 225 216
rect 223 215 224 216
rect 222 215 223 216
rect 221 215 222 216
rect 220 215 221 216
rect 219 215 220 216
rect 218 215 219 216
rect 217 215 218 216
rect 216 215 217 216
rect 215 215 216 216
rect 214 215 215 216
rect 213 215 214 216
rect 212 215 213 216
rect 211 215 212 216
rect 210 215 211 216
rect 209 215 210 216
rect 208 215 209 216
rect 207 215 208 216
rect 206 215 207 216
rect 205 215 206 216
rect 204 215 205 216
rect 203 215 204 216
rect 202 215 203 216
rect 201 215 202 216
rect 200 215 201 216
rect 199 215 200 216
rect 198 215 199 216
rect 197 215 198 216
rect 196 215 197 216
rect 195 215 196 216
rect 194 215 195 216
rect 193 215 194 216
rect 192 215 193 216
rect 191 215 192 216
rect 190 215 191 216
rect 189 215 190 216
rect 188 215 189 216
rect 187 215 188 216
rect 186 215 187 216
rect 185 215 186 216
rect 184 215 185 216
rect 145 215 146 216
rect 144 215 145 216
rect 143 215 144 216
rect 142 215 143 216
rect 141 215 142 216
rect 140 215 141 216
rect 139 215 140 216
rect 138 215 139 216
rect 137 215 138 216
rect 136 215 137 216
rect 135 215 136 216
rect 134 215 135 216
rect 133 215 134 216
rect 132 215 133 216
rect 131 215 132 216
rect 130 215 131 216
rect 129 215 130 216
rect 128 215 129 216
rect 127 215 128 216
rect 126 215 127 216
rect 125 215 126 216
rect 124 215 125 216
rect 123 215 124 216
rect 122 215 123 216
rect 121 215 122 216
rect 120 215 121 216
rect 119 215 120 216
rect 118 215 119 216
rect 117 215 118 216
rect 116 215 117 216
rect 115 215 116 216
rect 114 215 115 216
rect 113 215 114 216
rect 112 215 113 216
rect 111 215 112 216
rect 110 215 111 216
rect 109 215 110 216
rect 108 215 109 216
rect 107 215 108 216
rect 106 215 107 216
rect 105 215 106 216
rect 104 215 105 216
rect 103 215 104 216
rect 102 215 103 216
rect 101 215 102 216
rect 100 215 101 216
rect 99 215 100 216
rect 98 215 99 216
rect 97 215 98 216
rect 96 215 97 216
rect 95 215 96 216
rect 66 215 67 216
rect 65 215 66 216
rect 64 215 65 216
rect 63 215 64 216
rect 62 215 63 216
rect 61 215 62 216
rect 60 215 61 216
rect 59 215 60 216
rect 58 215 59 216
rect 57 215 58 216
rect 56 215 57 216
rect 55 215 56 216
rect 54 215 55 216
rect 53 215 54 216
rect 52 215 53 216
rect 51 215 52 216
rect 50 215 51 216
rect 49 215 50 216
rect 48 215 49 216
rect 47 215 48 216
rect 46 215 47 216
rect 45 215 46 216
rect 44 215 45 216
rect 43 215 44 216
rect 42 215 43 216
rect 41 215 42 216
rect 40 215 41 216
rect 39 215 40 216
rect 38 215 39 216
rect 37 215 38 216
rect 36 215 37 216
rect 35 215 36 216
rect 34 215 35 216
rect 33 215 34 216
rect 32 215 33 216
rect 31 215 32 216
rect 30 215 31 216
rect 29 215 30 216
rect 28 215 29 216
rect 27 215 28 216
rect 26 215 27 216
rect 25 215 26 216
rect 24 215 25 216
rect 23 215 24 216
rect 22 215 23 216
rect 21 215 22 216
rect 20 215 21 216
rect 19 215 20 216
rect 18 215 19 216
rect 17 215 18 216
rect 16 215 17 216
rect 15 215 16 216
rect 14 215 15 216
rect 13 215 14 216
rect 12 215 13 216
rect 11 215 12 216
rect 10 215 11 216
rect 9 215 10 216
rect 8 215 9 216
rect 7 215 8 216
rect 6 215 7 216
rect 5 215 6 216
rect 478 216 479 217
rect 477 216 478 217
rect 476 216 477 217
rect 460 216 461 217
rect 459 216 460 217
rect 458 216 459 217
rect 435 216 436 217
rect 434 216 435 217
rect 433 216 434 217
rect 432 216 433 217
rect 431 216 432 217
rect 430 216 431 217
rect 429 216 430 217
rect 428 216 429 217
rect 427 216 428 217
rect 426 216 427 217
rect 425 216 426 217
rect 424 216 425 217
rect 423 216 424 217
rect 422 216 423 217
rect 421 216 422 217
rect 408 216 409 217
rect 407 216 408 217
rect 406 216 407 217
rect 405 216 406 217
rect 404 216 405 217
rect 403 216 404 217
rect 402 216 403 217
rect 401 216 402 217
rect 400 216 401 217
rect 399 216 400 217
rect 398 216 399 217
rect 397 216 398 217
rect 396 216 397 217
rect 358 216 359 217
rect 357 216 358 217
rect 356 216 357 217
rect 355 216 356 217
rect 354 216 355 217
rect 353 216 354 217
rect 352 216 353 217
rect 351 216 352 217
rect 350 216 351 217
rect 349 216 350 217
rect 348 216 349 217
rect 347 216 348 217
rect 346 216 347 217
rect 345 216 346 217
rect 344 216 345 217
rect 296 216 297 217
rect 295 216 296 217
rect 294 216 295 217
rect 293 216 294 217
rect 292 216 293 217
rect 291 216 292 217
rect 290 216 291 217
rect 289 216 290 217
rect 288 216 289 217
rect 287 216 288 217
rect 286 216 287 217
rect 285 216 286 217
rect 284 216 285 217
rect 283 216 284 217
rect 282 216 283 217
rect 281 216 282 217
rect 280 216 281 217
rect 279 216 280 217
rect 278 216 279 217
rect 277 216 278 217
rect 276 216 277 217
rect 275 216 276 217
rect 274 216 275 217
rect 273 216 274 217
rect 272 216 273 217
rect 271 216 272 217
rect 270 216 271 217
rect 269 216 270 217
rect 268 216 269 217
rect 267 216 268 217
rect 266 216 267 217
rect 265 216 266 217
rect 264 216 265 217
rect 263 216 264 217
rect 262 216 263 217
rect 261 216 262 217
rect 260 216 261 217
rect 259 216 260 217
rect 258 216 259 217
rect 257 216 258 217
rect 256 216 257 217
rect 255 216 256 217
rect 254 216 255 217
rect 253 216 254 217
rect 252 216 253 217
rect 251 216 252 217
rect 250 216 251 217
rect 249 216 250 217
rect 248 216 249 217
rect 247 216 248 217
rect 246 216 247 217
rect 245 216 246 217
rect 244 216 245 217
rect 243 216 244 217
rect 242 216 243 217
rect 241 216 242 217
rect 240 216 241 217
rect 239 216 240 217
rect 238 216 239 217
rect 237 216 238 217
rect 236 216 237 217
rect 235 216 236 217
rect 234 216 235 217
rect 233 216 234 217
rect 232 216 233 217
rect 231 216 232 217
rect 230 216 231 217
rect 229 216 230 217
rect 228 216 229 217
rect 227 216 228 217
rect 226 216 227 217
rect 225 216 226 217
rect 224 216 225 217
rect 223 216 224 217
rect 222 216 223 217
rect 221 216 222 217
rect 220 216 221 217
rect 219 216 220 217
rect 218 216 219 217
rect 217 216 218 217
rect 216 216 217 217
rect 215 216 216 217
rect 214 216 215 217
rect 213 216 214 217
rect 212 216 213 217
rect 211 216 212 217
rect 210 216 211 217
rect 209 216 210 217
rect 208 216 209 217
rect 207 216 208 217
rect 206 216 207 217
rect 205 216 206 217
rect 204 216 205 217
rect 203 216 204 217
rect 202 216 203 217
rect 201 216 202 217
rect 200 216 201 217
rect 199 216 200 217
rect 198 216 199 217
rect 197 216 198 217
rect 196 216 197 217
rect 195 216 196 217
rect 194 216 195 217
rect 193 216 194 217
rect 192 216 193 217
rect 191 216 192 217
rect 190 216 191 217
rect 189 216 190 217
rect 188 216 189 217
rect 187 216 188 217
rect 186 216 187 217
rect 185 216 186 217
rect 184 216 185 217
rect 183 216 184 217
rect 182 216 183 217
rect 181 216 182 217
rect 144 216 145 217
rect 143 216 144 217
rect 142 216 143 217
rect 141 216 142 217
rect 140 216 141 217
rect 139 216 140 217
rect 138 216 139 217
rect 137 216 138 217
rect 136 216 137 217
rect 135 216 136 217
rect 134 216 135 217
rect 133 216 134 217
rect 132 216 133 217
rect 131 216 132 217
rect 130 216 131 217
rect 129 216 130 217
rect 128 216 129 217
rect 127 216 128 217
rect 126 216 127 217
rect 125 216 126 217
rect 124 216 125 217
rect 123 216 124 217
rect 122 216 123 217
rect 121 216 122 217
rect 120 216 121 217
rect 119 216 120 217
rect 118 216 119 217
rect 117 216 118 217
rect 116 216 117 217
rect 115 216 116 217
rect 114 216 115 217
rect 113 216 114 217
rect 112 216 113 217
rect 111 216 112 217
rect 110 216 111 217
rect 109 216 110 217
rect 108 216 109 217
rect 107 216 108 217
rect 106 216 107 217
rect 105 216 106 217
rect 104 216 105 217
rect 103 216 104 217
rect 102 216 103 217
rect 101 216 102 217
rect 100 216 101 217
rect 99 216 100 217
rect 98 216 99 217
rect 97 216 98 217
rect 67 216 68 217
rect 66 216 67 217
rect 65 216 66 217
rect 64 216 65 217
rect 63 216 64 217
rect 62 216 63 217
rect 61 216 62 217
rect 60 216 61 217
rect 59 216 60 217
rect 58 216 59 217
rect 57 216 58 217
rect 56 216 57 217
rect 55 216 56 217
rect 54 216 55 217
rect 53 216 54 217
rect 52 216 53 217
rect 51 216 52 217
rect 50 216 51 217
rect 49 216 50 217
rect 48 216 49 217
rect 47 216 48 217
rect 46 216 47 217
rect 45 216 46 217
rect 44 216 45 217
rect 43 216 44 217
rect 42 216 43 217
rect 41 216 42 217
rect 40 216 41 217
rect 39 216 40 217
rect 38 216 39 217
rect 37 216 38 217
rect 36 216 37 217
rect 35 216 36 217
rect 34 216 35 217
rect 33 216 34 217
rect 32 216 33 217
rect 31 216 32 217
rect 30 216 31 217
rect 29 216 30 217
rect 28 216 29 217
rect 27 216 28 217
rect 26 216 27 217
rect 25 216 26 217
rect 24 216 25 217
rect 23 216 24 217
rect 22 216 23 217
rect 21 216 22 217
rect 20 216 21 217
rect 19 216 20 217
rect 18 216 19 217
rect 17 216 18 217
rect 16 216 17 217
rect 15 216 16 217
rect 14 216 15 217
rect 13 216 14 217
rect 12 216 13 217
rect 11 216 12 217
rect 10 216 11 217
rect 9 216 10 217
rect 8 216 9 217
rect 7 216 8 217
rect 6 216 7 217
rect 5 216 6 217
rect 478 217 479 218
rect 477 217 478 218
rect 476 217 477 218
rect 475 217 476 218
rect 474 217 475 218
rect 473 217 474 218
rect 472 217 473 218
rect 471 217 472 218
rect 470 217 471 218
rect 469 217 470 218
rect 468 217 469 218
rect 467 217 468 218
rect 466 217 467 218
rect 465 217 466 218
rect 464 217 465 218
rect 463 217 464 218
rect 462 217 463 218
rect 461 217 462 218
rect 460 217 461 218
rect 459 217 460 218
rect 458 217 459 218
rect 435 217 436 218
rect 434 217 435 218
rect 433 217 434 218
rect 432 217 433 218
rect 431 217 432 218
rect 430 217 431 218
rect 429 217 430 218
rect 428 217 429 218
rect 427 217 428 218
rect 426 217 427 218
rect 425 217 426 218
rect 404 217 405 218
rect 403 217 404 218
rect 402 217 403 218
rect 401 217 402 218
rect 400 217 401 218
rect 399 217 400 218
rect 398 217 399 218
rect 397 217 398 218
rect 396 217 397 218
rect 395 217 396 218
rect 359 217 360 218
rect 358 217 359 218
rect 357 217 358 218
rect 356 217 357 218
rect 355 217 356 218
rect 354 217 355 218
rect 353 217 354 218
rect 352 217 353 218
rect 351 217 352 218
rect 350 217 351 218
rect 349 217 350 218
rect 348 217 349 218
rect 347 217 348 218
rect 293 217 294 218
rect 292 217 293 218
rect 291 217 292 218
rect 290 217 291 218
rect 289 217 290 218
rect 288 217 289 218
rect 287 217 288 218
rect 286 217 287 218
rect 285 217 286 218
rect 284 217 285 218
rect 283 217 284 218
rect 282 217 283 218
rect 281 217 282 218
rect 280 217 281 218
rect 279 217 280 218
rect 278 217 279 218
rect 277 217 278 218
rect 276 217 277 218
rect 275 217 276 218
rect 274 217 275 218
rect 273 217 274 218
rect 272 217 273 218
rect 271 217 272 218
rect 270 217 271 218
rect 269 217 270 218
rect 268 217 269 218
rect 267 217 268 218
rect 266 217 267 218
rect 265 217 266 218
rect 264 217 265 218
rect 263 217 264 218
rect 262 217 263 218
rect 261 217 262 218
rect 260 217 261 218
rect 259 217 260 218
rect 258 217 259 218
rect 257 217 258 218
rect 256 217 257 218
rect 255 217 256 218
rect 254 217 255 218
rect 253 217 254 218
rect 252 217 253 218
rect 251 217 252 218
rect 250 217 251 218
rect 249 217 250 218
rect 248 217 249 218
rect 247 217 248 218
rect 246 217 247 218
rect 245 217 246 218
rect 244 217 245 218
rect 243 217 244 218
rect 242 217 243 218
rect 241 217 242 218
rect 240 217 241 218
rect 239 217 240 218
rect 238 217 239 218
rect 237 217 238 218
rect 236 217 237 218
rect 235 217 236 218
rect 234 217 235 218
rect 233 217 234 218
rect 232 217 233 218
rect 231 217 232 218
rect 230 217 231 218
rect 229 217 230 218
rect 228 217 229 218
rect 227 217 228 218
rect 226 217 227 218
rect 225 217 226 218
rect 224 217 225 218
rect 223 217 224 218
rect 222 217 223 218
rect 221 217 222 218
rect 220 217 221 218
rect 219 217 220 218
rect 218 217 219 218
rect 217 217 218 218
rect 216 217 217 218
rect 215 217 216 218
rect 214 217 215 218
rect 213 217 214 218
rect 212 217 213 218
rect 211 217 212 218
rect 210 217 211 218
rect 209 217 210 218
rect 208 217 209 218
rect 207 217 208 218
rect 206 217 207 218
rect 205 217 206 218
rect 204 217 205 218
rect 203 217 204 218
rect 202 217 203 218
rect 201 217 202 218
rect 200 217 201 218
rect 199 217 200 218
rect 198 217 199 218
rect 197 217 198 218
rect 196 217 197 218
rect 195 217 196 218
rect 194 217 195 218
rect 193 217 194 218
rect 192 217 193 218
rect 191 217 192 218
rect 190 217 191 218
rect 189 217 190 218
rect 188 217 189 218
rect 187 217 188 218
rect 186 217 187 218
rect 185 217 186 218
rect 184 217 185 218
rect 183 217 184 218
rect 182 217 183 218
rect 181 217 182 218
rect 180 217 181 218
rect 179 217 180 218
rect 143 217 144 218
rect 142 217 143 218
rect 141 217 142 218
rect 140 217 141 218
rect 139 217 140 218
rect 138 217 139 218
rect 137 217 138 218
rect 136 217 137 218
rect 135 217 136 218
rect 134 217 135 218
rect 133 217 134 218
rect 132 217 133 218
rect 131 217 132 218
rect 130 217 131 218
rect 129 217 130 218
rect 128 217 129 218
rect 127 217 128 218
rect 126 217 127 218
rect 125 217 126 218
rect 124 217 125 218
rect 123 217 124 218
rect 122 217 123 218
rect 121 217 122 218
rect 120 217 121 218
rect 119 217 120 218
rect 118 217 119 218
rect 117 217 118 218
rect 116 217 117 218
rect 115 217 116 218
rect 114 217 115 218
rect 113 217 114 218
rect 112 217 113 218
rect 111 217 112 218
rect 110 217 111 218
rect 109 217 110 218
rect 108 217 109 218
rect 107 217 108 218
rect 106 217 107 218
rect 105 217 106 218
rect 104 217 105 218
rect 103 217 104 218
rect 102 217 103 218
rect 101 217 102 218
rect 100 217 101 218
rect 99 217 100 218
rect 68 217 69 218
rect 67 217 68 218
rect 66 217 67 218
rect 65 217 66 218
rect 64 217 65 218
rect 63 217 64 218
rect 62 217 63 218
rect 61 217 62 218
rect 60 217 61 218
rect 59 217 60 218
rect 58 217 59 218
rect 57 217 58 218
rect 56 217 57 218
rect 55 217 56 218
rect 54 217 55 218
rect 53 217 54 218
rect 52 217 53 218
rect 51 217 52 218
rect 50 217 51 218
rect 49 217 50 218
rect 48 217 49 218
rect 47 217 48 218
rect 46 217 47 218
rect 45 217 46 218
rect 44 217 45 218
rect 43 217 44 218
rect 42 217 43 218
rect 41 217 42 218
rect 40 217 41 218
rect 39 217 40 218
rect 38 217 39 218
rect 37 217 38 218
rect 36 217 37 218
rect 35 217 36 218
rect 34 217 35 218
rect 33 217 34 218
rect 32 217 33 218
rect 31 217 32 218
rect 30 217 31 218
rect 29 217 30 218
rect 28 217 29 218
rect 27 217 28 218
rect 26 217 27 218
rect 25 217 26 218
rect 24 217 25 218
rect 23 217 24 218
rect 22 217 23 218
rect 21 217 22 218
rect 20 217 21 218
rect 19 217 20 218
rect 18 217 19 218
rect 17 217 18 218
rect 16 217 17 218
rect 15 217 16 218
rect 14 217 15 218
rect 13 217 14 218
rect 12 217 13 218
rect 11 217 12 218
rect 10 217 11 218
rect 9 217 10 218
rect 8 217 9 218
rect 7 217 8 218
rect 6 217 7 218
rect 5 217 6 218
rect 478 218 479 219
rect 477 218 478 219
rect 476 218 477 219
rect 475 218 476 219
rect 474 218 475 219
rect 473 218 474 219
rect 472 218 473 219
rect 471 218 472 219
rect 470 218 471 219
rect 469 218 470 219
rect 468 218 469 219
rect 467 218 468 219
rect 466 218 467 219
rect 465 218 466 219
rect 464 218 465 219
rect 463 218 464 219
rect 462 218 463 219
rect 461 218 462 219
rect 460 218 461 219
rect 459 218 460 219
rect 458 218 459 219
rect 436 218 437 219
rect 435 218 436 219
rect 434 218 435 219
rect 433 218 434 219
rect 432 218 433 219
rect 431 218 432 219
rect 430 218 431 219
rect 429 218 430 219
rect 428 218 429 219
rect 427 218 428 219
rect 402 218 403 219
rect 401 218 402 219
rect 400 218 401 219
rect 399 218 400 219
rect 398 218 399 219
rect 397 218 398 219
rect 396 218 397 219
rect 395 218 396 219
rect 359 218 360 219
rect 358 218 359 219
rect 357 218 358 219
rect 356 218 357 219
rect 355 218 356 219
rect 354 218 355 219
rect 353 218 354 219
rect 352 218 353 219
rect 351 218 352 219
rect 350 218 351 219
rect 291 218 292 219
rect 290 218 291 219
rect 289 218 290 219
rect 288 218 289 219
rect 287 218 288 219
rect 286 218 287 219
rect 285 218 286 219
rect 284 218 285 219
rect 283 218 284 219
rect 282 218 283 219
rect 281 218 282 219
rect 280 218 281 219
rect 279 218 280 219
rect 278 218 279 219
rect 277 218 278 219
rect 276 218 277 219
rect 275 218 276 219
rect 274 218 275 219
rect 273 218 274 219
rect 272 218 273 219
rect 271 218 272 219
rect 270 218 271 219
rect 269 218 270 219
rect 268 218 269 219
rect 267 218 268 219
rect 266 218 267 219
rect 265 218 266 219
rect 264 218 265 219
rect 263 218 264 219
rect 262 218 263 219
rect 261 218 262 219
rect 260 218 261 219
rect 259 218 260 219
rect 258 218 259 219
rect 257 218 258 219
rect 256 218 257 219
rect 255 218 256 219
rect 254 218 255 219
rect 253 218 254 219
rect 252 218 253 219
rect 251 218 252 219
rect 250 218 251 219
rect 249 218 250 219
rect 248 218 249 219
rect 247 218 248 219
rect 246 218 247 219
rect 245 218 246 219
rect 244 218 245 219
rect 243 218 244 219
rect 242 218 243 219
rect 241 218 242 219
rect 240 218 241 219
rect 239 218 240 219
rect 238 218 239 219
rect 237 218 238 219
rect 236 218 237 219
rect 235 218 236 219
rect 234 218 235 219
rect 233 218 234 219
rect 232 218 233 219
rect 231 218 232 219
rect 230 218 231 219
rect 229 218 230 219
rect 228 218 229 219
rect 227 218 228 219
rect 226 218 227 219
rect 225 218 226 219
rect 224 218 225 219
rect 223 218 224 219
rect 222 218 223 219
rect 221 218 222 219
rect 220 218 221 219
rect 219 218 220 219
rect 218 218 219 219
rect 217 218 218 219
rect 216 218 217 219
rect 215 218 216 219
rect 214 218 215 219
rect 213 218 214 219
rect 212 218 213 219
rect 211 218 212 219
rect 210 218 211 219
rect 209 218 210 219
rect 208 218 209 219
rect 207 218 208 219
rect 206 218 207 219
rect 205 218 206 219
rect 204 218 205 219
rect 203 218 204 219
rect 202 218 203 219
rect 201 218 202 219
rect 200 218 201 219
rect 199 218 200 219
rect 198 218 199 219
rect 197 218 198 219
rect 196 218 197 219
rect 195 218 196 219
rect 194 218 195 219
rect 193 218 194 219
rect 192 218 193 219
rect 191 218 192 219
rect 190 218 191 219
rect 189 218 190 219
rect 188 218 189 219
rect 187 218 188 219
rect 186 218 187 219
rect 185 218 186 219
rect 184 218 185 219
rect 183 218 184 219
rect 182 218 183 219
rect 181 218 182 219
rect 180 218 181 219
rect 179 218 180 219
rect 178 218 179 219
rect 177 218 178 219
rect 143 218 144 219
rect 142 218 143 219
rect 141 218 142 219
rect 140 218 141 219
rect 139 218 140 219
rect 138 218 139 219
rect 137 218 138 219
rect 136 218 137 219
rect 135 218 136 219
rect 134 218 135 219
rect 133 218 134 219
rect 132 218 133 219
rect 131 218 132 219
rect 130 218 131 219
rect 129 218 130 219
rect 128 218 129 219
rect 127 218 128 219
rect 126 218 127 219
rect 125 218 126 219
rect 124 218 125 219
rect 123 218 124 219
rect 122 218 123 219
rect 121 218 122 219
rect 120 218 121 219
rect 119 218 120 219
rect 118 218 119 219
rect 117 218 118 219
rect 116 218 117 219
rect 115 218 116 219
rect 114 218 115 219
rect 113 218 114 219
rect 112 218 113 219
rect 111 218 112 219
rect 110 218 111 219
rect 109 218 110 219
rect 108 218 109 219
rect 107 218 108 219
rect 106 218 107 219
rect 105 218 106 219
rect 104 218 105 219
rect 103 218 104 219
rect 102 218 103 219
rect 101 218 102 219
rect 69 218 70 219
rect 68 218 69 219
rect 67 218 68 219
rect 66 218 67 219
rect 65 218 66 219
rect 64 218 65 219
rect 63 218 64 219
rect 62 218 63 219
rect 61 218 62 219
rect 60 218 61 219
rect 59 218 60 219
rect 58 218 59 219
rect 57 218 58 219
rect 56 218 57 219
rect 55 218 56 219
rect 54 218 55 219
rect 53 218 54 219
rect 52 218 53 219
rect 51 218 52 219
rect 50 218 51 219
rect 49 218 50 219
rect 48 218 49 219
rect 47 218 48 219
rect 46 218 47 219
rect 45 218 46 219
rect 44 218 45 219
rect 43 218 44 219
rect 42 218 43 219
rect 41 218 42 219
rect 40 218 41 219
rect 39 218 40 219
rect 38 218 39 219
rect 37 218 38 219
rect 36 218 37 219
rect 35 218 36 219
rect 34 218 35 219
rect 33 218 34 219
rect 32 218 33 219
rect 31 218 32 219
rect 30 218 31 219
rect 29 218 30 219
rect 28 218 29 219
rect 27 218 28 219
rect 26 218 27 219
rect 25 218 26 219
rect 24 218 25 219
rect 23 218 24 219
rect 22 218 23 219
rect 21 218 22 219
rect 20 218 21 219
rect 19 218 20 219
rect 18 218 19 219
rect 17 218 18 219
rect 16 218 17 219
rect 15 218 16 219
rect 14 218 15 219
rect 13 218 14 219
rect 12 218 13 219
rect 11 218 12 219
rect 10 218 11 219
rect 9 218 10 219
rect 8 218 9 219
rect 7 218 8 219
rect 6 218 7 219
rect 5 218 6 219
rect 478 219 479 220
rect 477 219 478 220
rect 476 219 477 220
rect 475 219 476 220
rect 474 219 475 220
rect 473 219 474 220
rect 472 219 473 220
rect 471 219 472 220
rect 470 219 471 220
rect 469 219 470 220
rect 468 219 469 220
rect 467 219 468 220
rect 466 219 467 220
rect 465 219 466 220
rect 464 219 465 220
rect 463 219 464 220
rect 462 219 463 220
rect 461 219 462 220
rect 460 219 461 220
rect 459 219 460 220
rect 458 219 459 220
rect 436 219 437 220
rect 435 219 436 220
rect 434 219 435 220
rect 433 219 434 220
rect 432 219 433 220
rect 431 219 432 220
rect 430 219 431 220
rect 429 219 430 220
rect 401 219 402 220
rect 400 219 401 220
rect 399 219 400 220
rect 398 219 399 220
rect 397 219 398 220
rect 396 219 397 220
rect 395 219 396 220
rect 394 219 395 220
rect 359 219 360 220
rect 358 219 359 220
rect 357 219 358 220
rect 356 219 357 220
rect 355 219 356 220
rect 354 219 355 220
rect 353 219 354 220
rect 288 219 289 220
rect 287 219 288 220
rect 286 219 287 220
rect 285 219 286 220
rect 284 219 285 220
rect 283 219 284 220
rect 282 219 283 220
rect 281 219 282 220
rect 280 219 281 220
rect 279 219 280 220
rect 278 219 279 220
rect 277 219 278 220
rect 276 219 277 220
rect 275 219 276 220
rect 274 219 275 220
rect 273 219 274 220
rect 272 219 273 220
rect 271 219 272 220
rect 270 219 271 220
rect 269 219 270 220
rect 268 219 269 220
rect 267 219 268 220
rect 266 219 267 220
rect 265 219 266 220
rect 264 219 265 220
rect 263 219 264 220
rect 262 219 263 220
rect 261 219 262 220
rect 260 219 261 220
rect 259 219 260 220
rect 258 219 259 220
rect 257 219 258 220
rect 256 219 257 220
rect 255 219 256 220
rect 254 219 255 220
rect 253 219 254 220
rect 252 219 253 220
rect 251 219 252 220
rect 250 219 251 220
rect 249 219 250 220
rect 248 219 249 220
rect 247 219 248 220
rect 246 219 247 220
rect 245 219 246 220
rect 244 219 245 220
rect 243 219 244 220
rect 242 219 243 220
rect 241 219 242 220
rect 240 219 241 220
rect 239 219 240 220
rect 238 219 239 220
rect 237 219 238 220
rect 236 219 237 220
rect 235 219 236 220
rect 234 219 235 220
rect 233 219 234 220
rect 232 219 233 220
rect 231 219 232 220
rect 230 219 231 220
rect 229 219 230 220
rect 228 219 229 220
rect 227 219 228 220
rect 226 219 227 220
rect 225 219 226 220
rect 224 219 225 220
rect 223 219 224 220
rect 222 219 223 220
rect 221 219 222 220
rect 220 219 221 220
rect 219 219 220 220
rect 218 219 219 220
rect 217 219 218 220
rect 216 219 217 220
rect 215 219 216 220
rect 214 219 215 220
rect 213 219 214 220
rect 212 219 213 220
rect 211 219 212 220
rect 210 219 211 220
rect 209 219 210 220
rect 208 219 209 220
rect 207 219 208 220
rect 206 219 207 220
rect 205 219 206 220
rect 204 219 205 220
rect 203 219 204 220
rect 202 219 203 220
rect 201 219 202 220
rect 200 219 201 220
rect 199 219 200 220
rect 198 219 199 220
rect 197 219 198 220
rect 196 219 197 220
rect 195 219 196 220
rect 194 219 195 220
rect 193 219 194 220
rect 192 219 193 220
rect 191 219 192 220
rect 190 219 191 220
rect 189 219 190 220
rect 188 219 189 220
rect 187 219 188 220
rect 186 219 187 220
rect 185 219 186 220
rect 184 219 185 220
rect 183 219 184 220
rect 182 219 183 220
rect 181 219 182 220
rect 180 219 181 220
rect 179 219 180 220
rect 178 219 179 220
rect 177 219 178 220
rect 176 219 177 220
rect 175 219 176 220
rect 142 219 143 220
rect 141 219 142 220
rect 140 219 141 220
rect 139 219 140 220
rect 138 219 139 220
rect 137 219 138 220
rect 136 219 137 220
rect 135 219 136 220
rect 134 219 135 220
rect 133 219 134 220
rect 132 219 133 220
rect 131 219 132 220
rect 130 219 131 220
rect 129 219 130 220
rect 128 219 129 220
rect 127 219 128 220
rect 126 219 127 220
rect 125 219 126 220
rect 124 219 125 220
rect 123 219 124 220
rect 122 219 123 220
rect 121 219 122 220
rect 120 219 121 220
rect 119 219 120 220
rect 118 219 119 220
rect 117 219 118 220
rect 116 219 117 220
rect 115 219 116 220
rect 114 219 115 220
rect 113 219 114 220
rect 112 219 113 220
rect 111 219 112 220
rect 110 219 111 220
rect 109 219 110 220
rect 108 219 109 220
rect 107 219 108 220
rect 106 219 107 220
rect 105 219 106 220
rect 104 219 105 220
rect 103 219 104 220
rect 102 219 103 220
rect 70 219 71 220
rect 69 219 70 220
rect 68 219 69 220
rect 67 219 68 220
rect 66 219 67 220
rect 65 219 66 220
rect 64 219 65 220
rect 63 219 64 220
rect 62 219 63 220
rect 61 219 62 220
rect 60 219 61 220
rect 59 219 60 220
rect 58 219 59 220
rect 57 219 58 220
rect 56 219 57 220
rect 55 219 56 220
rect 54 219 55 220
rect 53 219 54 220
rect 52 219 53 220
rect 51 219 52 220
rect 50 219 51 220
rect 49 219 50 220
rect 48 219 49 220
rect 47 219 48 220
rect 46 219 47 220
rect 45 219 46 220
rect 44 219 45 220
rect 43 219 44 220
rect 42 219 43 220
rect 41 219 42 220
rect 40 219 41 220
rect 39 219 40 220
rect 38 219 39 220
rect 37 219 38 220
rect 36 219 37 220
rect 35 219 36 220
rect 34 219 35 220
rect 33 219 34 220
rect 32 219 33 220
rect 31 219 32 220
rect 30 219 31 220
rect 29 219 30 220
rect 28 219 29 220
rect 27 219 28 220
rect 26 219 27 220
rect 25 219 26 220
rect 24 219 25 220
rect 23 219 24 220
rect 22 219 23 220
rect 21 219 22 220
rect 20 219 21 220
rect 19 219 20 220
rect 18 219 19 220
rect 17 219 18 220
rect 16 219 17 220
rect 15 219 16 220
rect 14 219 15 220
rect 13 219 14 220
rect 12 219 13 220
rect 11 219 12 220
rect 10 219 11 220
rect 9 219 10 220
rect 8 219 9 220
rect 7 219 8 220
rect 6 219 7 220
rect 5 219 6 220
rect 478 220 479 221
rect 477 220 478 221
rect 476 220 477 221
rect 475 220 476 221
rect 474 220 475 221
rect 473 220 474 221
rect 472 220 473 221
rect 471 220 472 221
rect 470 220 471 221
rect 469 220 470 221
rect 468 220 469 221
rect 467 220 468 221
rect 466 220 467 221
rect 465 220 466 221
rect 464 220 465 221
rect 463 220 464 221
rect 462 220 463 221
rect 461 220 462 221
rect 460 220 461 221
rect 459 220 460 221
rect 458 220 459 221
rect 437 220 438 221
rect 436 220 437 221
rect 435 220 436 221
rect 434 220 435 221
rect 433 220 434 221
rect 432 220 433 221
rect 431 220 432 221
rect 430 220 431 221
rect 399 220 400 221
rect 398 220 399 221
rect 397 220 398 221
rect 396 220 397 221
rect 395 220 396 221
rect 394 220 395 221
rect 360 220 361 221
rect 359 220 360 221
rect 358 220 359 221
rect 357 220 358 221
rect 356 220 357 221
rect 287 220 288 221
rect 286 220 287 221
rect 285 220 286 221
rect 284 220 285 221
rect 283 220 284 221
rect 282 220 283 221
rect 281 220 282 221
rect 280 220 281 221
rect 279 220 280 221
rect 278 220 279 221
rect 277 220 278 221
rect 276 220 277 221
rect 275 220 276 221
rect 274 220 275 221
rect 273 220 274 221
rect 272 220 273 221
rect 271 220 272 221
rect 270 220 271 221
rect 269 220 270 221
rect 268 220 269 221
rect 267 220 268 221
rect 266 220 267 221
rect 265 220 266 221
rect 264 220 265 221
rect 263 220 264 221
rect 262 220 263 221
rect 261 220 262 221
rect 260 220 261 221
rect 259 220 260 221
rect 258 220 259 221
rect 257 220 258 221
rect 256 220 257 221
rect 255 220 256 221
rect 254 220 255 221
rect 253 220 254 221
rect 252 220 253 221
rect 251 220 252 221
rect 250 220 251 221
rect 249 220 250 221
rect 248 220 249 221
rect 247 220 248 221
rect 246 220 247 221
rect 245 220 246 221
rect 244 220 245 221
rect 243 220 244 221
rect 242 220 243 221
rect 241 220 242 221
rect 240 220 241 221
rect 239 220 240 221
rect 238 220 239 221
rect 237 220 238 221
rect 236 220 237 221
rect 235 220 236 221
rect 234 220 235 221
rect 233 220 234 221
rect 232 220 233 221
rect 231 220 232 221
rect 230 220 231 221
rect 229 220 230 221
rect 228 220 229 221
rect 227 220 228 221
rect 226 220 227 221
rect 225 220 226 221
rect 224 220 225 221
rect 223 220 224 221
rect 222 220 223 221
rect 221 220 222 221
rect 220 220 221 221
rect 219 220 220 221
rect 218 220 219 221
rect 217 220 218 221
rect 216 220 217 221
rect 215 220 216 221
rect 214 220 215 221
rect 213 220 214 221
rect 212 220 213 221
rect 211 220 212 221
rect 210 220 211 221
rect 209 220 210 221
rect 208 220 209 221
rect 207 220 208 221
rect 206 220 207 221
rect 205 220 206 221
rect 204 220 205 221
rect 203 220 204 221
rect 202 220 203 221
rect 201 220 202 221
rect 200 220 201 221
rect 199 220 200 221
rect 198 220 199 221
rect 197 220 198 221
rect 196 220 197 221
rect 195 220 196 221
rect 194 220 195 221
rect 193 220 194 221
rect 192 220 193 221
rect 191 220 192 221
rect 190 220 191 221
rect 189 220 190 221
rect 188 220 189 221
rect 187 220 188 221
rect 186 220 187 221
rect 185 220 186 221
rect 184 220 185 221
rect 183 220 184 221
rect 182 220 183 221
rect 181 220 182 221
rect 180 220 181 221
rect 179 220 180 221
rect 178 220 179 221
rect 177 220 178 221
rect 176 220 177 221
rect 175 220 176 221
rect 174 220 175 221
rect 173 220 174 221
rect 142 220 143 221
rect 141 220 142 221
rect 140 220 141 221
rect 139 220 140 221
rect 138 220 139 221
rect 137 220 138 221
rect 136 220 137 221
rect 135 220 136 221
rect 134 220 135 221
rect 133 220 134 221
rect 132 220 133 221
rect 131 220 132 221
rect 130 220 131 221
rect 129 220 130 221
rect 128 220 129 221
rect 127 220 128 221
rect 126 220 127 221
rect 125 220 126 221
rect 124 220 125 221
rect 123 220 124 221
rect 122 220 123 221
rect 121 220 122 221
rect 120 220 121 221
rect 119 220 120 221
rect 118 220 119 221
rect 117 220 118 221
rect 116 220 117 221
rect 115 220 116 221
rect 114 220 115 221
rect 113 220 114 221
rect 112 220 113 221
rect 111 220 112 221
rect 110 220 111 221
rect 109 220 110 221
rect 108 220 109 221
rect 107 220 108 221
rect 106 220 107 221
rect 105 220 106 221
rect 104 220 105 221
rect 71 220 72 221
rect 70 220 71 221
rect 69 220 70 221
rect 68 220 69 221
rect 67 220 68 221
rect 66 220 67 221
rect 65 220 66 221
rect 64 220 65 221
rect 63 220 64 221
rect 62 220 63 221
rect 61 220 62 221
rect 60 220 61 221
rect 59 220 60 221
rect 58 220 59 221
rect 57 220 58 221
rect 56 220 57 221
rect 55 220 56 221
rect 54 220 55 221
rect 53 220 54 221
rect 52 220 53 221
rect 51 220 52 221
rect 50 220 51 221
rect 49 220 50 221
rect 48 220 49 221
rect 47 220 48 221
rect 46 220 47 221
rect 45 220 46 221
rect 44 220 45 221
rect 43 220 44 221
rect 42 220 43 221
rect 41 220 42 221
rect 40 220 41 221
rect 39 220 40 221
rect 38 220 39 221
rect 37 220 38 221
rect 36 220 37 221
rect 35 220 36 221
rect 34 220 35 221
rect 33 220 34 221
rect 32 220 33 221
rect 31 220 32 221
rect 30 220 31 221
rect 29 220 30 221
rect 28 220 29 221
rect 27 220 28 221
rect 26 220 27 221
rect 25 220 26 221
rect 24 220 25 221
rect 23 220 24 221
rect 22 220 23 221
rect 21 220 22 221
rect 20 220 21 221
rect 19 220 20 221
rect 18 220 19 221
rect 17 220 18 221
rect 16 220 17 221
rect 15 220 16 221
rect 14 220 15 221
rect 13 220 14 221
rect 12 220 13 221
rect 11 220 12 221
rect 10 220 11 221
rect 9 220 10 221
rect 8 220 9 221
rect 7 220 8 221
rect 6 220 7 221
rect 5 220 6 221
rect 4 220 5 221
rect 478 221 479 222
rect 477 221 478 222
rect 469 221 470 222
rect 468 221 469 222
rect 459 221 460 222
rect 458 221 459 222
rect 437 221 438 222
rect 436 221 437 222
rect 435 221 436 222
rect 434 221 435 222
rect 433 221 434 222
rect 432 221 433 222
rect 398 221 399 222
rect 397 221 398 222
rect 396 221 397 222
rect 395 221 396 222
rect 394 221 395 222
rect 360 221 361 222
rect 359 221 360 222
rect 358 221 359 222
rect 285 221 286 222
rect 284 221 285 222
rect 283 221 284 222
rect 282 221 283 222
rect 281 221 282 222
rect 280 221 281 222
rect 279 221 280 222
rect 278 221 279 222
rect 277 221 278 222
rect 276 221 277 222
rect 275 221 276 222
rect 274 221 275 222
rect 273 221 274 222
rect 272 221 273 222
rect 271 221 272 222
rect 270 221 271 222
rect 269 221 270 222
rect 268 221 269 222
rect 267 221 268 222
rect 266 221 267 222
rect 265 221 266 222
rect 264 221 265 222
rect 263 221 264 222
rect 262 221 263 222
rect 261 221 262 222
rect 260 221 261 222
rect 259 221 260 222
rect 258 221 259 222
rect 257 221 258 222
rect 256 221 257 222
rect 255 221 256 222
rect 254 221 255 222
rect 253 221 254 222
rect 252 221 253 222
rect 251 221 252 222
rect 250 221 251 222
rect 249 221 250 222
rect 248 221 249 222
rect 247 221 248 222
rect 246 221 247 222
rect 245 221 246 222
rect 244 221 245 222
rect 243 221 244 222
rect 242 221 243 222
rect 241 221 242 222
rect 240 221 241 222
rect 239 221 240 222
rect 238 221 239 222
rect 237 221 238 222
rect 236 221 237 222
rect 235 221 236 222
rect 234 221 235 222
rect 233 221 234 222
rect 232 221 233 222
rect 231 221 232 222
rect 230 221 231 222
rect 229 221 230 222
rect 228 221 229 222
rect 227 221 228 222
rect 226 221 227 222
rect 225 221 226 222
rect 224 221 225 222
rect 223 221 224 222
rect 222 221 223 222
rect 221 221 222 222
rect 220 221 221 222
rect 219 221 220 222
rect 218 221 219 222
rect 217 221 218 222
rect 216 221 217 222
rect 215 221 216 222
rect 214 221 215 222
rect 213 221 214 222
rect 212 221 213 222
rect 211 221 212 222
rect 210 221 211 222
rect 209 221 210 222
rect 208 221 209 222
rect 207 221 208 222
rect 206 221 207 222
rect 205 221 206 222
rect 204 221 205 222
rect 203 221 204 222
rect 202 221 203 222
rect 201 221 202 222
rect 200 221 201 222
rect 199 221 200 222
rect 198 221 199 222
rect 197 221 198 222
rect 196 221 197 222
rect 195 221 196 222
rect 194 221 195 222
rect 193 221 194 222
rect 192 221 193 222
rect 191 221 192 222
rect 190 221 191 222
rect 189 221 190 222
rect 188 221 189 222
rect 187 221 188 222
rect 186 221 187 222
rect 185 221 186 222
rect 184 221 185 222
rect 183 221 184 222
rect 182 221 183 222
rect 181 221 182 222
rect 180 221 181 222
rect 179 221 180 222
rect 178 221 179 222
rect 177 221 178 222
rect 176 221 177 222
rect 175 221 176 222
rect 174 221 175 222
rect 173 221 174 222
rect 172 221 173 222
rect 171 221 172 222
rect 142 221 143 222
rect 141 221 142 222
rect 140 221 141 222
rect 139 221 140 222
rect 138 221 139 222
rect 137 221 138 222
rect 136 221 137 222
rect 135 221 136 222
rect 134 221 135 222
rect 133 221 134 222
rect 132 221 133 222
rect 131 221 132 222
rect 130 221 131 222
rect 129 221 130 222
rect 128 221 129 222
rect 127 221 128 222
rect 126 221 127 222
rect 125 221 126 222
rect 124 221 125 222
rect 123 221 124 222
rect 122 221 123 222
rect 121 221 122 222
rect 120 221 121 222
rect 119 221 120 222
rect 118 221 119 222
rect 117 221 118 222
rect 116 221 117 222
rect 115 221 116 222
rect 114 221 115 222
rect 113 221 114 222
rect 112 221 113 222
rect 111 221 112 222
rect 110 221 111 222
rect 109 221 110 222
rect 108 221 109 222
rect 107 221 108 222
rect 106 221 107 222
rect 105 221 106 222
rect 73 221 74 222
rect 72 221 73 222
rect 71 221 72 222
rect 70 221 71 222
rect 69 221 70 222
rect 68 221 69 222
rect 67 221 68 222
rect 66 221 67 222
rect 65 221 66 222
rect 64 221 65 222
rect 63 221 64 222
rect 62 221 63 222
rect 61 221 62 222
rect 60 221 61 222
rect 59 221 60 222
rect 58 221 59 222
rect 57 221 58 222
rect 56 221 57 222
rect 55 221 56 222
rect 54 221 55 222
rect 53 221 54 222
rect 52 221 53 222
rect 51 221 52 222
rect 50 221 51 222
rect 49 221 50 222
rect 48 221 49 222
rect 47 221 48 222
rect 46 221 47 222
rect 45 221 46 222
rect 44 221 45 222
rect 43 221 44 222
rect 42 221 43 222
rect 41 221 42 222
rect 40 221 41 222
rect 39 221 40 222
rect 38 221 39 222
rect 37 221 38 222
rect 36 221 37 222
rect 35 221 36 222
rect 34 221 35 222
rect 33 221 34 222
rect 32 221 33 222
rect 31 221 32 222
rect 30 221 31 222
rect 29 221 30 222
rect 28 221 29 222
rect 27 221 28 222
rect 26 221 27 222
rect 25 221 26 222
rect 24 221 25 222
rect 23 221 24 222
rect 22 221 23 222
rect 21 221 22 222
rect 20 221 21 222
rect 19 221 20 222
rect 18 221 19 222
rect 17 221 18 222
rect 16 221 17 222
rect 15 221 16 222
rect 14 221 15 222
rect 13 221 14 222
rect 12 221 13 222
rect 11 221 12 222
rect 10 221 11 222
rect 9 221 10 222
rect 8 221 9 222
rect 7 221 8 222
rect 6 221 7 222
rect 5 221 6 222
rect 4 221 5 222
rect 478 222 479 223
rect 469 222 470 223
rect 458 222 459 223
rect 437 222 438 223
rect 436 222 437 223
rect 435 222 436 223
rect 434 222 435 223
rect 433 222 434 223
rect 397 222 398 223
rect 396 222 397 223
rect 395 222 396 223
rect 394 222 395 223
rect 393 222 394 223
rect 360 222 361 223
rect 283 222 284 223
rect 282 222 283 223
rect 281 222 282 223
rect 280 222 281 223
rect 279 222 280 223
rect 278 222 279 223
rect 277 222 278 223
rect 276 222 277 223
rect 275 222 276 223
rect 274 222 275 223
rect 273 222 274 223
rect 272 222 273 223
rect 271 222 272 223
rect 270 222 271 223
rect 269 222 270 223
rect 268 222 269 223
rect 267 222 268 223
rect 266 222 267 223
rect 265 222 266 223
rect 264 222 265 223
rect 263 222 264 223
rect 262 222 263 223
rect 261 222 262 223
rect 260 222 261 223
rect 259 222 260 223
rect 258 222 259 223
rect 257 222 258 223
rect 256 222 257 223
rect 255 222 256 223
rect 254 222 255 223
rect 253 222 254 223
rect 252 222 253 223
rect 251 222 252 223
rect 250 222 251 223
rect 249 222 250 223
rect 248 222 249 223
rect 247 222 248 223
rect 246 222 247 223
rect 245 222 246 223
rect 244 222 245 223
rect 243 222 244 223
rect 242 222 243 223
rect 241 222 242 223
rect 240 222 241 223
rect 239 222 240 223
rect 238 222 239 223
rect 237 222 238 223
rect 236 222 237 223
rect 235 222 236 223
rect 234 222 235 223
rect 233 222 234 223
rect 232 222 233 223
rect 231 222 232 223
rect 230 222 231 223
rect 229 222 230 223
rect 228 222 229 223
rect 227 222 228 223
rect 226 222 227 223
rect 225 222 226 223
rect 224 222 225 223
rect 223 222 224 223
rect 222 222 223 223
rect 221 222 222 223
rect 220 222 221 223
rect 219 222 220 223
rect 218 222 219 223
rect 217 222 218 223
rect 216 222 217 223
rect 215 222 216 223
rect 214 222 215 223
rect 213 222 214 223
rect 212 222 213 223
rect 211 222 212 223
rect 210 222 211 223
rect 209 222 210 223
rect 208 222 209 223
rect 207 222 208 223
rect 206 222 207 223
rect 205 222 206 223
rect 204 222 205 223
rect 203 222 204 223
rect 202 222 203 223
rect 201 222 202 223
rect 200 222 201 223
rect 199 222 200 223
rect 198 222 199 223
rect 197 222 198 223
rect 196 222 197 223
rect 195 222 196 223
rect 194 222 195 223
rect 193 222 194 223
rect 192 222 193 223
rect 191 222 192 223
rect 190 222 191 223
rect 189 222 190 223
rect 188 222 189 223
rect 187 222 188 223
rect 186 222 187 223
rect 185 222 186 223
rect 184 222 185 223
rect 183 222 184 223
rect 182 222 183 223
rect 181 222 182 223
rect 180 222 181 223
rect 179 222 180 223
rect 178 222 179 223
rect 177 222 178 223
rect 176 222 177 223
rect 175 222 176 223
rect 174 222 175 223
rect 173 222 174 223
rect 172 222 173 223
rect 171 222 172 223
rect 170 222 171 223
rect 169 222 170 223
rect 142 222 143 223
rect 141 222 142 223
rect 140 222 141 223
rect 139 222 140 223
rect 138 222 139 223
rect 137 222 138 223
rect 136 222 137 223
rect 135 222 136 223
rect 134 222 135 223
rect 133 222 134 223
rect 132 222 133 223
rect 131 222 132 223
rect 130 222 131 223
rect 129 222 130 223
rect 128 222 129 223
rect 127 222 128 223
rect 126 222 127 223
rect 125 222 126 223
rect 124 222 125 223
rect 123 222 124 223
rect 122 222 123 223
rect 121 222 122 223
rect 120 222 121 223
rect 119 222 120 223
rect 118 222 119 223
rect 117 222 118 223
rect 116 222 117 223
rect 115 222 116 223
rect 114 222 115 223
rect 113 222 114 223
rect 112 222 113 223
rect 111 222 112 223
rect 110 222 111 223
rect 109 222 110 223
rect 108 222 109 223
rect 107 222 108 223
rect 74 222 75 223
rect 73 222 74 223
rect 72 222 73 223
rect 71 222 72 223
rect 70 222 71 223
rect 69 222 70 223
rect 68 222 69 223
rect 67 222 68 223
rect 66 222 67 223
rect 65 222 66 223
rect 64 222 65 223
rect 63 222 64 223
rect 62 222 63 223
rect 61 222 62 223
rect 60 222 61 223
rect 59 222 60 223
rect 58 222 59 223
rect 57 222 58 223
rect 56 222 57 223
rect 55 222 56 223
rect 54 222 55 223
rect 53 222 54 223
rect 52 222 53 223
rect 51 222 52 223
rect 50 222 51 223
rect 49 222 50 223
rect 48 222 49 223
rect 47 222 48 223
rect 46 222 47 223
rect 45 222 46 223
rect 44 222 45 223
rect 43 222 44 223
rect 42 222 43 223
rect 41 222 42 223
rect 40 222 41 223
rect 39 222 40 223
rect 38 222 39 223
rect 37 222 38 223
rect 36 222 37 223
rect 35 222 36 223
rect 34 222 35 223
rect 33 222 34 223
rect 32 222 33 223
rect 31 222 32 223
rect 30 222 31 223
rect 29 222 30 223
rect 28 222 29 223
rect 27 222 28 223
rect 26 222 27 223
rect 25 222 26 223
rect 24 222 25 223
rect 23 222 24 223
rect 22 222 23 223
rect 21 222 22 223
rect 20 222 21 223
rect 19 222 20 223
rect 18 222 19 223
rect 17 222 18 223
rect 16 222 17 223
rect 15 222 16 223
rect 14 222 15 223
rect 13 222 14 223
rect 12 222 13 223
rect 11 222 12 223
rect 10 222 11 223
rect 9 222 10 223
rect 8 222 9 223
rect 7 222 8 223
rect 6 222 7 223
rect 5 222 6 223
rect 4 222 5 223
rect 478 223 479 224
rect 470 223 471 224
rect 469 223 470 224
rect 468 223 469 224
rect 458 223 459 224
rect 437 223 438 224
rect 436 223 437 224
rect 435 223 436 224
rect 434 223 435 224
rect 433 223 434 224
rect 397 223 398 224
rect 396 223 397 224
rect 395 223 396 224
rect 394 223 395 224
rect 393 223 394 224
rect 282 223 283 224
rect 281 223 282 224
rect 280 223 281 224
rect 279 223 280 224
rect 278 223 279 224
rect 277 223 278 224
rect 276 223 277 224
rect 275 223 276 224
rect 274 223 275 224
rect 273 223 274 224
rect 272 223 273 224
rect 271 223 272 224
rect 270 223 271 224
rect 269 223 270 224
rect 268 223 269 224
rect 267 223 268 224
rect 266 223 267 224
rect 265 223 266 224
rect 264 223 265 224
rect 263 223 264 224
rect 262 223 263 224
rect 261 223 262 224
rect 260 223 261 224
rect 259 223 260 224
rect 258 223 259 224
rect 257 223 258 224
rect 256 223 257 224
rect 255 223 256 224
rect 254 223 255 224
rect 253 223 254 224
rect 252 223 253 224
rect 251 223 252 224
rect 250 223 251 224
rect 249 223 250 224
rect 248 223 249 224
rect 247 223 248 224
rect 246 223 247 224
rect 245 223 246 224
rect 244 223 245 224
rect 243 223 244 224
rect 242 223 243 224
rect 241 223 242 224
rect 240 223 241 224
rect 239 223 240 224
rect 238 223 239 224
rect 237 223 238 224
rect 236 223 237 224
rect 235 223 236 224
rect 234 223 235 224
rect 233 223 234 224
rect 232 223 233 224
rect 231 223 232 224
rect 230 223 231 224
rect 229 223 230 224
rect 228 223 229 224
rect 227 223 228 224
rect 226 223 227 224
rect 225 223 226 224
rect 224 223 225 224
rect 223 223 224 224
rect 222 223 223 224
rect 221 223 222 224
rect 220 223 221 224
rect 219 223 220 224
rect 218 223 219 224
rect 217 223 218 224
rect 216 223 217 224
rect 215 223 216 224
rect 214 223 215 224
rect 213 223 214 224
rect 212 223 213 224
rect 211 223 212 224
rect 210 223 211 224
rect 209 223 210 224
rect 208 223 209 224
rect 207 223 208 224
rect 206 223 207 224
rect 205 223 206 224
rect 204 223 205 224
rect 203 223 204 224
rect 202 223 203 224
rect 201 223 202 224
rect 200 223 201 224
rect 199 223 200 224
rect 198 223 199 224
rect 197 223 198 224
rect 196 223 197 224
rect 195 223 196 224
rect 194 223 195 224
rect 193 223 194 224
rect 192 223 193 224
rect 191 223 192 224
rect 190 223 191 224
rect 189 223 190 224
rect 188 223 189 224
rect 187 223 188 224
rect 186 223 187 224
rect 185 223 186 224
rect 184 223 185 224
rect 183 223 184 224
rect 182 223 183 224
rect 181 223 182 224
rect 180 223 181 224
rect 179 223 180 224
rect 178 223 179 224
rect 177 223 178 224
rect 176 223 177 224
rect 175 223 176 224
rect 174 223 175 224
rect 173 223 174 224
rect 172 223 173 224
rect 171 223 172 224
rect 170 223 171 224
rect 169 223 170 224
rect 168 223 169 224
rect 167 223 168 224
rect 142 223 143 224
rect 141 223 142 224
rect 140 223 141 224
rect 139 223 140 224
rect 138 223 139 224
rect 137 223 138 224
rect 136 223 137 224
rect 135 223 136 224
rect 134 223 135 224
rect 133 223 134 224
rect 132 223 133 224
rect 131 223 132 224
rect 130 223 131 224
rect 129 223 130 224
rect 128 223 129 224
rect 127 223 128 224
rect 126 223 127 224
rect 125 223 126 224
rect 124 223 125 224
rect 123 223 124 224
rect 122 223 123 224
rect 121 223 122 224
rect 120 223 121 224
rect 119 223 120 224
rect 118 223 119 224
rect 117 223 118 224
rect 116 223 117 224
rect 115 223 116 224
rect 114 223 115 224
rect 113 223 114 224
rect 112 223 113 224
rect 111 223 112 224
rect 110 223 111 224
rect 109 223 110 224
rect 108 223 109 224
rect 75 223 76 224
rect 74 223 75 224
rect 73 223 74 224
rect 72 223 73 224
rect 71 223 72 224
rect 70 223 71 224
rect 69 223 70 224
rect 68 223 69 224
rect 67 223 68 224
rect 66 223 67 224
rect 65 223 66 224
rect 64 223 65 224
rect 63 223 64 224
rect 62 223 63 224
rect 61 223 62 224
rect 60 223 61 224
rect 59 223 60 224
rect 58 223 59 224
rect 57 223 58 224
rect 56 223 57 224
rect 55 223 56 224
rect 54 223 55 224
rect 53 223 54 224
rect 52 223 53 224
rect 51 223 52 224
rect 50 223 51 224
rect 49 223 50 224
rect 48 223 49 224
rect 47 223 48 224
rect 46 223 47 224
rect 45 223 46 224
rect 44 223 45 224
rect 43 223 44 224
rect 42 223 43 224
rect 41 223 42 224
rect 40 223 41 224
rect 39 223 40 224
rect 38 223 39 224
rect 37 223 38 224
rect 36 223 37 224
rect 35 223 36 224
rect 34 223 35 224
rect 33 223 34 224
rect 32 223 33 224
rect 31 223 32 224
rect 30 223 31 224
rect 29 223 30 224
rect 28 223 29 224
rect 27 223 28 224
rect 26 223 27 224
rect 25 223 26 224
rect 24 223 25 224
rect 23 223 24 224
rect 22 223 23 224
rect 21 223 22 224
rect 20 223 21 224
rect 19 223 20 224
rect 18 223 19 224
rect 17 223 18 224
rect 16 223 17 224
rect 15 223 16 224
rect 14 223 15 224
rect 13 223 14 224
rect 12 223 13 224
rect 11 223 12 224
rect 10 223 11 224
rect 9 223 10 224
rect 8 223 9 224
rect 7 223 8 224
rect 6 223 7 224
rect 5 223 6 224
rect 4 223 5 224
rect 472 224 473 225
rect 471 224 472 225
rect 470 224 471 225
rect 469 224 470 225
rect 468 224 469 225
rect 459 224 460 225
rect 458 224 459 225
rect 438 224 439 225
rect 437 224 438 225
rect 436 224 437 225
rect 435 224 436 225
rect 434 224 435 225
rect 396 224 397 225
rect 395 224 396 225
rect 394 224 395 225
rect 393 224 394 225
rect 280 224 281 225
rect 279 224 280 225
rect 278 224 279 225
rect 277 224 278 225
rect 276 224 277 225
rect 275 224 276 225
rect 274 224 275 225
rect 273 224 274 225
rect 272 224 273 225
rect 271 224 272 225
rect 270 224 271 225
rect 269 224 270 225
rect 268 224 269 225
rect 267 224 268 225
rect 266 224 267 225
rect 265 224 266 225
rect 264 224 265 225
rect 263 224 264 225
rect 262 224 263 225
rect 261 224 262 225
rect 260 224 261 225
rect 259 224 260 225
rect 258 224 259 225
rect 257 224 258 225
rect 256 224 257 225
rect 255 224 256 225
rect 254 224 255 225
rect 253 224 254 225
rect 252 224 253 225
rect 251 224 252 225
rect 250 224 251 225
rect 249 224 250 225
rect 248 224 249 225
rect 247 224 248 225
rect 246 224 247 225
rect 245 224 246 225
rect 244 224 245 225
rect 243 224 244 225
rect 242 224 243 225
rect 241 224 242 225
rect 240 224 241 225
rect 239 224 240 225
rect 238 224 239 225
rect 237 224 238 225
rect 236 224 237 225
rect 235 224 236 225
rect 234 224 235 225
rect 233 224 234 225
rect 232 224 233 225
rect 231 224 232 225
rect 230 224 231 225
rect 229 224 230 225
rect 228 224 229 225
rect 227 224 228 225
rect 226 224 227 225
rect 225 224 226 225
rect 224 224 225 225
rect 223 224 224 225
rect 222 224 223 225
rect 221 224 222 225
rect 220 224 221 225
rect 219 224 220 225
rect 218 224 219 225
rect 217 224 218 225
rect 216 224 217 225
rect 215 224 216 225
rect 214 224 215 225
rect 213 224 214 225
rect 212 224 213 225
rect 211 224 212 225
rect 210 224 211 225
rect 209 224 210 225
rect 208 224 209 225
rect 207 224 208 225
rect 206 224 207 225
rect 205 224 206 225
rect 204 224 205 225
rect 203 224 204 225
rect 202 224 203 225
rect 201 224 202 225
rect 200 224 201 225
rect 199 224 200 225
rect 198 224 199 225
rect 197 224 198 225
rect 196 224 197 225
rect 195 224 196 225
rect 194 224 195 225
rect 193 224 194 225
rect 192 224 193 225
rect 191 224 192 225
rect 190 224 191 225
rect 189 224 190 225
rect 188 224 189 225
rect 187 224 188 225
rect 186 224 187 225
rect 185 224 186 225
rect 184 224 185 225
rect 183 224 184 225
rect 182 224 183 225
rect 181 224 182 225
rect 180 224 181 225
rect 179 224 180 225
rect 178 224 179 225
rect 177 224 178 225
rect 176 224 177 225
rect 175 224 176 225
rect 174 224 175 225
rect 173 224 174 225
rect 172 224 173 225
rect 171 224 172 225
rect 170 224 171 225
rect 169 224 170 225
rect 168 224 169 225
rect 167 224 168 225
rect 166 224 167 225
rect 165 224 166 225
rect 142 224 143 225
rect 141 224 142 225
rect 140 224 141 225
rect 139 224 140 225
rect 138 224 139 225
rect 137 224 138 225
rect 136 224 137 225
rect 135 224 136 225
rect 134 224 135 225
rect 133 224 134 225
rect 132 224 133 225
rect 131 224 132 225
rect 130 224 131 225
rect 129 224 130 225
rect 128 224 129 225
rect 127 224 128 225
rect 126 224 127 225
rect 125 224 126 225
rect 124 224 125 225
rect 123 224 124 225
rect 122 224 123 225
rect 121 224 122 225
rect 120 224 121 225
rect 119 224 120 225
rect 118 224 119 225
rect 117 224 118 225
rect 116 224 117 225
rect 115 224 116 225
rect 114 224 115 225
rect 113 224 114 225
rect 112 224 113 225
rect 111 224 112 225
rect 110 224 111 225
rect 109 224 110 225
rect 77 224 78 225
rect 76 224 77 225
rect 75 224 76 225
rect 74 224 75 225
rect 73 224 74 225
rect 72 224 73 225
rect 71 224 72 225
rect 70 224 71 225
rect 69 224 70 225
rect 68 224 69 225
rect 67 224 68 225
rect 66 224 67 225
rect 65 224 66 225
rect 64 224 65 225
rect 63 224 64 225
rect 62 224 63 225
rect 61 224 62 225
rect 60 224 61 225
rect 59 224 60 225
rect 58 224 59 225
rect 57 224 58 225
rect 56 224 57 225
rect 55 224 56 225
rect 54 224 55 225
rect 53 224 54 225
rect 52 224 53 225
rect 51 224 52 225
rect 50 224 51 225
rect 49 224 50 225
rect 48 224 49 225
rect 47 224 48 225
rect 46 224 47 225
rect 45 224 46 225
rect 44 224 45 225
rect 43 224 44 225
rect 42 224 43 225
rect 41 224 42 225
rect 40 224 41 225
rect 39 224 40 225
rect 38 224 39 225
rect 37 224 38 225
rect 36 224 37 225
rect 35 224 36 225
rect 34 224 35 225
rect 33 224 34 225
rect 32 224 33 225
rect 31 224 32 225
rect 30 224 31 225
rect 29 224 30 225
rect 28 224 29 225
rect 27 224 28 225
rect 26 224 27 225
rect 25 224 26 225
rect 24 224 25 225
rect 23 224 24 225
rect 22 224 23 225
rect 21 224 22 225
rect 20 224 21 225
rect 19 224 20 225
rect 18 224 19 225
rect 17 224 18 225
rect 16 224 17 225
rect 15 224 16 225
rect 14 224 15 225
rect 13 224 14 225
rect 12 224 13 225
rect 11 224 12 225
rect 10 224 11 225
rect 9 224 10 225
rect 8 224 9 225
rect 7 224 8 225
rect 6 224 7 225
rect 5 224 6 225
rect 4 224 5 225
rect 3 224 4 225
rect 474 225 475 226
rect 473 225 474 226
rect 472 225 473 226
rect 471 225 472 226
rect 470 225 471 226
rect 469 225 470 226
rect 468 225 469 226
rect 467 225 468 226
rect 459 225 460 226
rect 458 225 459 226
rect 438 225 439 226
rect 437 225 438 226
rect 436 225 437 226
rect 435 225 436 226
rect 395 225 396 226
rect 394 225 395 226
rect 393 225 394 226
rect 279 225 280 226
rect 278 225 279 226
rect 277 225 278 226
rect 276 225 277 226
rect 275 225 276 226
rect 274 225 275 226
rect 273 225 274 226
rect 272 225 273 226
rect 271 225 272 226
rect 270 225 271 226
rect 269 225 270 226
rect 268 225 269 226
rect 267 225 268 226
rect 266 225 267 226
rect 265 225 266 226
rect 264 225 265 226
rect 263 225 264 226
rect 262 225 263 226
rect 261 225 262 226
rect 260 225 261 226
rect 259 225 260 226
rect 258 225 259 226
rect 257 225 258 226
rect 256 225 257 226
rect 255 225 256 226
rect 254 225 255 226
rect 253 225 254 226
rect 252 225 253 226
rect 251 225 252 226
rect 250 225 251 226
rect 249 225 250 226
rect 248 225 249 226
rect 247 225 248 226
rect 246 225 247 226
rect 245 225 246 226
rect 244 225 245 226
rect 243 225 244 226
rect 242 225 243 226
rect 241 225 242 226
rect 240 225 241 226
rect 239 225 240 226
rect 238 225 239 226
rect 237 225 238 226
rect 236 225 237 226
rect 235 225 236 226
rect 234 225 235 226
rect 233 225 234 226
rect 232 225 233 226
rect 231 225 232 226
rect 230 225 231 226
rect 229 225 230 226
rect 228 225 229 226
rect 227 225 228 226
rect 226 225 227 226
rect 225 225 226 226
rect 224 225 225 226
rect 223 225 224 226
rect 222 225 223 226
rect 221 225 222 226
rect 220 225 221 226
rect 219 225 220 226
rect 218 225 219 226
rect 217 225 218 226
rect 216 225 217 226
rect 215 225 216 226
rect 214 225 215 226
rect 213 225 214 226
rect 212 225 213 226
rect 211 225 212 226
rect 210 225 211 226
rect 209 225 210 226
rect 208 225 209 226
rect 207 225 208 226
rect 206 225 207 226
rect 205 225 206 226
rect 204 225 205 226
rect 203 225 204 226
rect 202 225 203 226
rect 201 225 202 226
rect 200 225 201 226
rect 199 225 200 226
rect 198 225 199 226
rect 197 225 198 226
rect 196 225 197 226
rect 195 225 196 226
rect 194 225 195 226
rect 193 225 194 226
rect 192 225 193 226
rect 191 225 192 226
rect 190 225 191 226
rect 189 225 190 226
rect 188 225 189 226
rect 187 225 188 226
rect 186 225 187 226
rect 185 225 186 226
rect 184 225 185 226
rect 183 225 184 226
rect 182 225 183 226
rect 181 225 182 226
rect 180 225 181 226
rect 179 225 180 226
rect 178 225 179 226
rect 177 225 178 226
rect 176 225 177 226
rect 175 225 176 226
rect 174 225 175 226
rect 173 225 174 226
rect 172 225 173 226
rect 171 225 172 226
rect 170 225 171 226
rect 169 225 170 226
rect 168 225 169 226
rect 167 225 168 226
rect 166 225 167 226
rect 165 225 166 226
rect 164 225 165 226
rect 163 225 164 226
rect 162 225 163 226
rect 142 225 143 226
rect 141 225 142 226
rect 140 225 141 226
rect 139 225 140 226
rect 138 225 139 226
rect 137 225 138 226
rect 136 225 137 226
rect 135 225 136 226
rect 134 225 135 226
rect 133 225 134 226
rect 132 225 133 226
rect 131 225 132 226
rect 130 225 131 226
rect 129 225 130 226
rect 128 225 129 226
rect 127 225 128 226
rect 126 225 127 226
rect 125 225 126 226
rect 124 225 125 226
rect 123 225 124 226
rect 122 225 123 226
rect 121 225 122 226
rect 120 225 121 226
rect 119 225 120 226
rect 118 225 119 226
rect 117 225 118 226
rect 116 225 117 226
rect 115 225 116 226
rect 114 225 115 226
rect 113 225 114 226
rect 112 225 113 226
rect 111 225 112 226
rect 110 225 111 226
rect 78 225 79 226
rect 77 225 78 226
rect 76 225 77 226
rect 75 225 76 226
rect 74 225 75 226
rect 73 225 74 226
rect 72 225 73 226
rect 71 225 72 226
rect 70 225 71 226
rect 69 225 70 226
rect 68 225 69 226
rect 67 225 68 226
rect 66 225 67 226
rect 65 225 66 226
rect 64 225 65 226
rect 63 225 64 226
rect 62 225 63 226
rect 61 225 62 226
rect 60 225 61 226
rect 59 225 60 226
rect 58 225 59 226
rect 57 225 58 226
rect 56 225 57 226
rect 55 225 56 226
rect 54 225 55 226
rect 53 225 54 226
rect 52 225 53 226
rect 51 225 52 226
rect 50 225 51 226
rect 49 225 50 226
rect 48 225 49 226
rect 47 225 48 226
rect 46 225 47 226
rect 45 225 46 226
rect 44 225 45 226
rect 43 225 44 226
rect 42 225 43 226
rect 41 225 42 226
rect 40 225 41 226
rect 39 225 40 226
rect 38 225 39 226
rect 37 225 38 226
rect 36 225 37 226
rect 35 225 36 226
rect 34 225 35 226
rect 33 225 34 226
rect 32 225 33 226
rect 31 225 32 226
rect 30 225 31 226
rect 29 225 30 226
rect 28 225 29 226
rect 27 225 28 226
rect 26 225 27 226
rect 25 225 26 226
rect 24 225 25 226
rect 23 225 24 226
rect 22 225 23 226
rect 21 225 22 226
rect 20 225 21 226
rect 19 225 20 226
rect 18 225 19 226
rect 17 225 18 226
rect 16 225 17 226
rect 15 225 16 226
rect 14 225 15 226
rect 13 225 14 226
rect 12 225 13 226
rect 11 225 12 226
rect 10 225 11 226
rect 9 225 10 226
rect 8 225 9 226
rect 7 225 8 226
rect 6 225 7 226
rect 5 225 6 226
rect 4 225 5 226
rect 3 225 4 226
rect 476 226 477 227
rect 475 226 476 227
rect 474 226 475 227
rect 473 226 474 227
rect 472 226 473 227
rect 471 226 472 227
rect 470 226 471 227
rect 469 226 470 227
rect 468 226 469 227
rect 467 226 468 227
rect 466 226 467 227
rect 465 226 466 227
rect 462 226 463 227
rect 461 226 462 227
rect 460 226 461 227
rect 459 226 460 227
rect 458 226 459 227
rect 438 226 439 227
rect 437 226 438 227
rect 436 226 437 227
rect 435 226 436 227
rect 395 226 396 227
rect 394 226 395 227
rect 393 226 394 227
rect 392 226 393 227
rect 278 226 279 227
rect 277 226 278 227
rect 276 226 277 227
rect 275 226 276 227
rect 274 226 275 227
rect 273 226 274 227
rect 272 226 273 227
rect 271 226 272 227
rect 270 226 271 227
rect 269 226 270 227
rect 268 226 269 227
rect 267 226 268 227
rect 266 226 267 227
rect 265 226 266 227
rect 264 226 265 227
rect 263 226 264 227
rect 262 226 263 227
rect 261 226 262 227
rect 260 226 261 227
rect 259 226 260 227
rect 258 226 259 227
rect 257 226 258 227
rect 256 226 257 227
rect 255 226 256 227
rect 254 226 255 227
rect 253 226 254 227
rect 252 226 253 227
rect 251 226 252 227
rect 250 226 251 227
rect 249 226 250 227
rect 248 226 249 227
rect 247 226 248 227
rect 246 226 247 227
rect 245 226 246 227
rect 244 226 245 227
rect 243 226 244 227
rect 242 226 243 227
rect 241 226 242 227
rect 240 226 241 227
rect 239 226 240 227
rect 238 226 239 227
rect 237 226 238 227
rect 236 226 237 227
rect 235 226 236 227
rect 234 226 235 227
rect 233 226 234 227
rect 232 226 233 227
rect 231 226 232 227
rect 230 226 231 227
rect 229 226 230 227
rect 228 226 229 227
rect 227 226 228 227
rect 226 226 227 227
rect 225 226 226 227
rect 224 226 225 227
rect 223 226 224 227
rect 222 226 223 227
rect 221 226 222 227
rect 220 226 221 227
rect 219 226 220 227
rect 218 226 219 227
rect 217 226 218 227
rect 216 226 217 227
rect 215 226 216 227
rect 214 226 215 227
rect 213 226 214 227
rect 212 226 213 227
rect 211 226 212 227
rect 210 226 211 227
rect 209 226 210 227
rect 208 226 209 227
rect 207 226 208 227
rect 206 226 207 227
rect 205 226 206 227
rect 204 226 205 227
rect 203 226 204 227
rect 202 226 203 227
rect 201 226 202 227
rect 200 226 201 227
rect 199 226 200 227
rect 198 226 199 227
rect 197 226 198 227
rect 196 226 197 227
rect 195 226 196 227
rect 194 226 195 227
rect 193 226 194 227
rect 192 226 193 227
rect 191 226 192 227
rect 190 226 191 227
rect 189 226 190 227
rect 188 226 189 227
rect 187 226 188 227
rect 186 226 187 227
rect 185 226 186 227
rect 184 226 185 227
rect 183 226 184 227
rect 182 226 183 227
rect 181 226 182 227
rect 180 226 181 227
rect 179 226 180 227
rect 178 226 179 227
rect 177 226 178 227
rect 176 226 177 227
rect 175 226 176 227
rect 174 226 175 227
rect 173 226 174 227
rect 172 226 173 227
rect 171 226 172 227
rect 170 226 171 227
rect 169 226 170 227
rect 168 226 169 227
rect 167 226 168 227
rect 166 226 167 227
rect 165 226 166 227
rect 164 226 165 227
rect 163 226 164 227
rect 162 226 163 227
rect 161 226 162 227
rect 160 226 161 227
rect 142 226 143 227
rect 141 226 142 227
rect 140 226 141 227
rect 139 226 140 227
rect 138 226 139 227
rect 137 226 138 227
rect 136 226 137 227
rect 135 226 136 227
rect 134 226 135 227
rect 133 226 134 227
rect 132 226 133 227
rect 131 226 132 227
rect 130 226 131 227
rect 129 226 130 227
rect 128 226 129 227
rect 127 226 128 227
rect 126 226 127 227
rect 125 226 126 227
rect 124 226 125 227
rect 123 226 124 227
rect 122 226 123 227
rect 121 226 122 227
rect 120 226 121 227
rect 119 226 120 227
rect 118 226 119 227
rect 117 226 118 227
rect 116 226 117 227
rect 115 226 116 227
rect 114 226 115 227
rect 113 226 114 227
rect 112 226 113 227
rect 111 226 112 227
rect 110 226 111 227
rect 80 226 81 227
rect 79 226 80 227
rect 78 226 79 227
rect 77 226 78 227
rect 76 226 77 227
rect 75 226 76 227
rect 74 226 75 227
rect 73 226 74 227
rect 72 226 73 227
rect 71 226 72 227
rect 70 226 71 227
rect 69 226 70 227
rect 68 226 69 227
rect 67 226 68 227
rect 66 226 67 227
rect 65 226 66 227
rect 64 226 65 227
rect 63 226 64 227
rect 62 226 63 227
rect 61 226 62 227
rect 60 226 61 227
rect 59 226 60 227
rect 58 226 59 227
rect 57 226 58 227
rect 56 226 57 227
rect 55 226 56 227
rect 54 226 55 227
rect 53 226 54 227
rect 52 226 53 227
rect 51 226 52 227
rect 50 226 51 227
rect 49 226 50 227
rect 48 226 49 227
rect 47 226 48 227
rect 46 226 47 227
rect 45 226 46 227
rect 44 226 45 227
rect 43 226 44 227
rect 42 226 43 227
rect 41 226 42 227
rect 40 226 41 227
rect 39 226 40 227
rect 38 226 39 227
rect 37 226 38 227
rect 36 226 37 227
rect 35 226 36 227
rect 34 226 35 227
rect 33 226 34 227
rect 32 226 33 227
rect 31 226 32 227
rect 30 226 31 227
rect 29 226 30 227
rect 28 226 29 227
rect 27 226 28 227
rect 26 226 27 227
rect 25 226 26 227
rect 24 226 25 227
rect 23 226 24 227
rect 22 226 23 227
rect 21 226 22 227
rect 20 226 21 227
rect 19 226 20 227
rect 18 226 19 227
rect 17 226 18 227
rect 16 226 17 227
rect 15 226 16 227
rect 14 226 15 227
rect 13 226 14 227
rect 12 226 13 227
rect 11 226 12 227
rect 10 226 11 227
rect 9 226 10 227
rect 8 226 9 227
rect 7 226 8 227
rect 6 226 7 227
rect 5 226 6 227
rect 4 226 5 227
rect 3 226 4 227
rect 477 227 478 228
rect 476 227 477 228
rect 475 227 476 228
rect 474 227 475 228
rect 473 227 474 228
rect 472 227 473 228
rect 471 227 472 228
rect 470 227 471 228
rect 469 227 470 228
rect 468 227 469 228
rect 467 227 468 228
rect 466 227 467 228
rect 465 227 466 228
rect 464 227 465 228
rect 463 227 464 228
rect 462 227 463 228
rect 461 227 462 228
rect 460 227 461 228
rect 459 227 460 228
rect 458 227 459 228
rect 438 227 439 228
rect 437 227 438 228
rect 436 227 437 228
rect 435 227 436 228
rect 395 227 396 228
rect 394 227 395 228
rect 393 227 394 228
rect 392 227 393 228
rect 276 227 277 228
rect 275 227 276 228
rect 274 227 275 228
rect 273 227 274 228
rect 272 227 273 228
rect 271 227 272 228
rect 270 227 271 228
rect 269 227 270 228
rect 268 227 269 228
rect 267 227 268 228
rect 266 227 267 228
rect 265 227 266 228
rect 264 227 265 228
rect 263 227 264 228
rect 262 227 263 228
rect 261 227 262 228
rect 260 227 261 228
rect 259 227 260 228
rect 258 227 259 228
rect 257 227 258 228
rect 256 227 257 228
rect 255 227 256 228
rect 254 227 255 228
rect 253 227 254 228
rect 252 227 253 228
rect 251 227 252 228
rect 250 227 251 228
rect 249 227 250 228
rect 248 227 249 228
rect 247 227 248 228
rect 246 227 247 228
rect 245 227 246 228
rect 244 227 245 228
rect 243 227 244 228
rect 242 227 243 228
rect 241 227 242 228
rect 240 227 241 228
rect 239 227 240 228
rect 238 227 239 228
rect 237 227 238 228
rect 236 227 237 228
rect 235 227 236 228
rect 234 227 235 228
rect 233 227 234 228
rect 232 227 233 228
rect 231 227 232 228
rect 230 227 231 228
rect 229 227 230 228
rect 228 227 229 228
rect 227 227 228 228
rect 226 227 227 228
rect 225 227 226 228
rect 224 227 225 228
rect 223 227 224 228
rect 222 227 223 228
rect 221 227 222 228
rect 220 227 221 228
rect 219 227 220 228
rect 218 227 219 228
rect 217 227 218 228
rect 216 227 217 228
rect 215 227 216 228
rect 214 227 215 228
rect 213 227 214 228
rect 212 227 213 228
rect 211 227 212 228
rect 210 227 211 228
rect 209 227 210 228
rect 208 227 209 228
rect 207 227 208 228
rect 206 227 207 228
rect 205 227 206 228
rect 204 227 205 228
rect 203 227 204 228
rect 202 227 203 228
rect 201 227 202 228
rect 200 227 201 228
rect 199 227 200 228
rect 198 227 199 228
rect 197 227 198 228
rect 196 227 197 228
rect 195 227 196 228
rect 194 227 195 228
rect 193 227 194 228
rect 192 227 193 228
rect 191 227 192 228
rect 190 227 191 228
rect 189 227 190 228
rect 188 227 189 228
rect 187 227 188 228
rect 186 227 187 228
rect 185 227 186 228
rect 184 227 185 228
rect 183 227 184 228
rect 182 227 183 228
rect 181 227 182 228
rect 180 227 181 228
rect 179 227 180 228
rect 178 227 179 228
rect 177 227 178 228
rect 176 227 177 228
rect 175 227 176 228
rect 174 227 175 228
rect 173 227 174 228
rect 172 227 173 228
rect 171 227 172 228
rect 170 227 171 228
rect 169 227 170 228
rect 168 227 169 228
rect 167 227 168 228
rect 166 227 167 228
rect 165 227 166 228
rect 164 227 165 228
rect 163 227 164 228
rect 162 227 163 228
rect 161 227 162 228
rect 160 227 161 228
rect 142 227 143 228
rect 141 227 142 228
rect 140 227 141 228
rect 139 227 140 228
rect 138 227 139 228
rect 137 227 138 228
rect 136 227 137 228
rect 135 227 136 228
rect 134 227 135 228
rect 133 227 134 228
rect 132 227 133 228
rect 131 227 132 228
rect 130 227 131 228
rect 129 227 130 228
rect 128 227 129 228
rect 127 227 128 228
rect 126 227 127 228
rect 125 227 126 228
rect 124 227 125 228
rect 123 227 124 228
rect 122 227 123 228
rect 121 227 122 228
rect 120 227 121 228
rect 119 227 120 228
rect 118 227 119 228
rect 117 227 118 228
rect 116 227 117 228
rect 115 227 116 228
rect 114 227 115 228
rect 113 227 114 228
rect 112 227 113 228
rect 111 227 112 228
rect 81 227 82 228
rect 80 227 81 228
rect 79 227 80 228
rect 78 227 79 228
rect 77 227 78 228
rect 76 227 77 228
rect 75 227 76 228
rect 74 227 75 228
rect 73 227 74 228
rect 72 227 73 228
rect 71 227 72 228
rect 70 227 71 228
rect 69 227 70 228
rect 68 227 69 228
rect 67 227 68 228
rect 66 227 67 228
rect 65 227 66 228
rect 64 227 65 228
rect 63 227 64 228
rect 62 227 63 228
rect 61 227 62 228
rect 60 227 61 228
rect 59 227 60 228
rect 58 227 59 228
rect 57 227 58 228
rect 56 227 57 228
rect 55 227 56 228
rect 54 227 55 228
rect 53 227 54 228
rect 52 227 53 228
rect 51 227 52 228
rect 50 227 51 228
rect 49 227 50 228
rect 48 227 49 228
rect 47 227 48 228
rect 46 227 47 228
rect 45 227 46 228
rect 44 227 45 228
rect 43 227 44 228
rect 42 227 43 228
rect 41 227 42 228
rect 40 227 41 228
rect 39 227 40 228
rect 38 227 39 228
rect 37 227 38 228
rect 36 227 37 228
rect 35 227 36 228
rect 34 227 35 228
rect 33 227 34 228
rect 32 227 33 228
rect 31 227 32 228
rect 30 227 31 228
rect 29 227 30 228
rect 28 227 29 228
rect 27 227 28 228
rect 26 227 27 228
rect 25 227 26 228
rect 24 227 25 228
rect 23 227 24 228
rect 22 227 23 228
rect 21 227 22 228
rect 20 227 21 228
rect 19 227 20 228
rect 18 227 19 228
rect 17 227 18 228
rect 16 227 17 228
rect 15 227 16 228
rect 14 227 15 228
rect 13 227 14 228
rect 12 227 13 228
rect 11 227 12 228
rect 10 227 11 228
rect 9 227 10 228
rect 8 227 9 228
rect 7 227 8 228
rect 6 227 7 228
rect 5 227 6 228
rect 4 227 5 228
rect 3 227 4 228
rect 478 228 479 229
rect 477 228 478 229
rect 476 228 477 229
rect 475 228 476 229
rect 474 228 475 229
rect 473 228 474 229
rect 472 228 473 229
rect 471 228 472 229
rect 467 228 468 229
rect 466 228 467 229
rect 465 228 466 229
rect 464 228 465 229
rect 463 228 464 229
rect 462 228 463 229
rect 461 228 462 229
rect 460 228 461 229
rect 459 228 460 229
rect 458 228 459 229
rect 438 228 439 229
rect 437 228 438 229
rect 436 228 437 229
rect 394 228 395 229
rect 393 228 394 229
rect 392 228 393 229
rect 275 228 276 229
rect 274 228 275 229
rect 273 228 274 229
rect 272 228 273 229
rect 271 228 272 229
rect 270 228 271 229
rect 269 228 270 229
rect 268 228 269 229
rect 267 228 268 229
rect 266 228 267 229
rect 265 228 266 229
rect 264 228 265 229
rect 263 228 264 229
rect 262 228 263 229
rect 261 228 262 229
rect 260 228 261 229
rect 259 228 260 229
rect 258 228 259 229
rect 257 228 258 229
rect 256 228 257 229
rect 255 228 256 229
rect 254 228 255 229
rect 253 228 254 229
rect 252 228 253 229
rect 251 228 252 229
rect 250 228 251 229
rect 249 228 250 229
rect 248 228 249 229
rect 247 228 248 229
rect 246 228 247 229
rect 245 228 246 229
rect 244 228 245 229
rect 243 228 244 229
rect 242 228 243 229
rect 241 228 242 229
rect 240 228 241 229
rect 239 228 240 229
rect 238 228 239 229
rect 237 228 238 229
rect 236 228 237 229
rect 235 228 236 229
rect 234 228 235 229
rect 233 228 234 229
rect 232 228 233 229
rect 231 228 232 229
rect 230 228 231 229
rect 229 228 230 229
rect 228 228 229 229
rect 227 228 228 229
rect 226 228 227 229
rect 225 228 226 229
rect 224 228 225 229
rect 223 228 224 229
rect 222 228 223 229
rect 221 228 222 229
rect 220 228 221 229
rect 219 228 220 229
rect 218 228 219 229
rect 217 228 218 229
rect 216 228 217 229
rect 215 228 216 229
rect 214 228 215 229
rect 213 228 214 229
rect 212 228 213 229
rect 211 228 212 229
rect 210 228 211 229
rect 209 228 210 229
rect 208 228 209 229
rect 207 228 208 229
rect 206 228 207 229
rect 205 228 206 229
rect 204 228 205 229
rect 203 228 204 229
rect 202 228 203 229
rect 201 228 202 229
rect 200 228 201 229
rect 199 228 200 229
rect 198 228 199 229
rect 197 228 198 229
rect 196 228 197 229
rect 195 228 196 229
rect 194 228 195 229
rect 193 228 194 229
rect 192 228 193 229
rect 191 228 192 229
rect 190 228 191 229
rect 189 228 190 229
rect 188 228 189 229
rect 187 228 188 229
rect 186 228 187 229
rect 185 228 186 229
rect 184 228 185 229
rect 183 228 184 229
rect 182 228 183 229
rect 181 228 182 229
rect 180 228 181 229
rect 179 228 180 229
rect 178 228 179 229
rect 177 228 178 229
rect 176 228 177 229
rect 175 228 176 229
rect 174 228 175 229
rect 173 228 174 229
rect 172 228 173 229
rect 171 228 172 229
rect 170 228 171 229
rect 169 228 170 229
rect 168 228 169 229
rect 167 228 168 229
rect 166 228 167 229
rect 165 228 166 229
rect 164 228 165 229
rect 163 228 164 229
rect 162 228 163 229
rect 161 228 162 229
rect 143 228 144 229
rect 142 228 143 229
rect 141 228 142 229
rect 140 228 141 229
rect 139 228 140 229
rect 138 228 139 229
rect 137 228 138 229
rect 136 228 137 229
rect 135 228 136 229
rect 134 228 135 229
rect 133 228 134 229
rect 132 228 133 229
rect 131 228 132 229
rect 130 228 131 229
rect 129 228 130 229
rect 128 228 129 229
rect 127 228 128 229
rect 126 228 127 229
rect 125 228 126 229
rect 124 228 125 229
rect 123 228 124 229
rect 122 228 123 229
rect 121 228 122 229
rect 120 228 121 229
rect 119 228 120 229
rect 118 228 119 229
rect 117 228 118 229
rect 116 228 117 229
rect 115 228 116 229
rect 114 228 115 229
rect 113 228 114 229
rect 112 228 113 229
rect 83 228 84 229
rect 82 228 83 229
rect 81 228 82 229
rect 80 228 81 229
rect 79 228 80 229
rect 78 228 79 229
rect 77 228 78 229
rect 76 228 77 229
rect 75 228 76 229
rect 74 228 75 229
rect 73 228 74 229
rect 72 228 73 229
rect 71 228 72 229
rect 70 228 71 229
rect 69 228 70 229
rect 68 228 69 229
rect 67 228 68 229
rect 66 228 67 229
rect 65 228 66 229
rect 64 228 65 229
rect 63 228 64 229
rect 62 228 63 229
rect 61 228 62 229
rect 60 228 61 229
rect 59 228 60 229
rect 58 228 59 229
rect 57 228 58 229
rect 56 228 57 229
rect 55 228 56 229
rect 54 228 55 229
rect 53 228 54 229
rect 52 228 53 229
rect 51 228 52 229
rect 50 228 51 229
rect 49 228 50 229
rect 48 228 49 229
rect 47 228 48 229
rect 46 228 47 229
rect 45 228 46 229
rect 44 228 45 229
rect 43 228 44 229
rect 42 228 43 229
rect 41 228 42 229
rect 40 228 41 229
rect 39 228 40 229
rect 38 228 39 229
rect 37 228 38 229
rect 36 228 37 229
rect 35 228 36 229
rect 34 228 35 229
rect 33 228 34 229
rect 32 228 33 229
rect 31 228 32 229
rect 30 228 31 229
rect 29 228 30 229
rect 28 228 29 229
rect 27 228 28 229
rect 26 228 27 229
rect 25 228 26 229
rect 24 228 25 229
rect 23 228 24 229
rect 22 228 23 229
rect 21 228 22 229
rect 20 228 21 229
rect 19 228 20 229
rect 18 228 19 229
rect 17 228 18 229
rect 16 228 17 229
rect 15 228 16 229
rect 14 228 15 229
rect 13 228 14 229
rect 12 228 13 229
rect 11 228 12 229
rect 10 228 11 229
rect 9 228 10 229
rect 8 228 9 229
rect 7 228 8 229
rect 6 228 7 229
rect 5 228 6 229
rect 4 228 5 229
rect 3 228 4 229
rect 478 229 479 230
rect 477 229 478 230
rect 476 229 477 230
rect 475 229 476 230
rect 474 229 475 230
rect 473 229 474 230
rect 472 229 473 230
rect 467 229 468 230
rect 466 229 467 230
rect 465 229 466 230
rect 464 229 465 230
rect 463 229 464 230
rect 462 229 463 230
rect 461 229 462 230
rect 460 229 461 230
rect 459 229 460 230
rect 438 229 439 230
rect 437 229 438 230
rect 436 229 437 230
rect 394 229 395 230
rect 393 229 394 230
rect 392 229 393 230
rect 274 229 275 230
rect 273 229 274 230
rect 272 229 273 230
rect 271 229 272 230
rect 270 229 271 230
rect 269 229 270 230
rect 268 229 269 230
rect 267 229 268 230
rect 266 229 267 230
rect 265 229 266 230
rect 264 229 265 230
rect 263 229 264 230
rect 262 229 263 230
rect 261 229 262 230
rect 260 229 261 230
rect 259 229 260 230
rect 258 229 259 230
rect 257 229 258 230
rect 256 229 257 230
rect 255 229 256 230
rect 254 229 255 230
rect 253 229 254 230
rect 252 229 253 230
rect 251 229 252 230
rect 250 229 251 230
rect 249 229 250 230
rect 248 229 249 230
rect 247 229 248 230
rect 246 229 247 230
rect 245 229 246 230
rect 244 229 245 230
rect 243 229 244 230
rect 242 229 243 230
rect 241 229 242 230
rect 240 229 241 230
rect 239 229 240 230
rect 238 229 239 230
rect 237 229 238 230
rect 236 229 237 230
rect 235 229 236 230
rect 234 229 235 230
rect 233 229 234 230
rect 232 229 233 230
rect 231 229 232 230
rect 230 229 231 230
rect 229 229 230 230
rect 228 229 229 230
rect 227 229 228 230
rect 226 229 227 230
rect 225 229 226 230
rect 224 229 225 230
rect 223 229 224 230
rect 222 229 223 230
rect 221 229 222 230
rect 220 229 221 230
rect 219 229 220 230
rect 218 229 219 230
rect 217 229 218 230
rect 216 229 217 230
rect 215 229 216 230
rect 214 229 215 230
rect 213 229 214 230
rect 212 229 213 230
rect 211 229 212 230
rect 210 229 211 230
rect 209 229 210 230
rect 208 229 209 230
rect 207 229 208 230
rect 206 229 207 230
rect 205 229 206 230
rect 204 229 205 230
rect 203 229 204 230
rect 202 229 203 230
rect 201 229 202 230
rect 200 229 201 230
rect 199 229 200 230
rect 198 229 199 230
rect 197 229 198 230
rect 196 229 197 230
rect 195 229 196 230
rect 194 229 195 230
rect 193 229 194 230
rect 192 229 193 230
rect 191 229 192 230
rect 190 229 191 230
rect 189 229 190 230
rect 188 229 189 230
rect 187 229 188 230
rect 186 229 187 230
rect 185 229 186 230
rect 184 229 185 230
rect 183 229 184 230
rect 182 229 183 230
rect 181 229 182 230
rect 180 229 181 230
rect 179 229 180 230
rect 178 229 179 230
rect 177 229 178 230
rect 176 229 177 230
rect 175 229 176 230
rect 174 229 175 230
rect 173 229 174 230
rect 172 229 173 230
rect 171 229 172 230
rect 170 229 171 230
rect 169 229 170 230
rect 168 229 169 230
rect 167 229 168 230
rect 166 229 167 230
rect 165 229 166 230
rect 164 229 165 230
rect 163 229 164 230
rect 162 229 163 230
rect 143 229 144 230
rect 142 229 143 230
rect 141 229 142 230
rect 140 229 141 230
rect 139 229 140 230
rect 138 229 139 230
rect 137 229 138 230
rect 136 229 137 230
rect 135 229 136 230
rect 134 229 135 230
rect 133 229 134 230
rect 132 229 133 230
rect 131 229 132 230
rect 130 229 131 230
rect 129 229 130 230
rect 128 229 129 230
rect 127 229 128 230
rect 126 229 127 230
rect 125 229 126 230
rect 124 229 125 230
rect 123 229 124 230
rect 122 229 123 230
rect 121 229 122 230
rect 120 229 121 230
rect 119 229 120 230
rect 118 229 119 230
rect 117 229 118 230
rect 116 229 117 230
rect 115 229 116 230
rect 114 229 115 230
rect 113 229 114 230
rect 112 229 113 230
rect 85 229 86 230
rect 84 229 85 230
rect 83 229 84 230
rect 82 229 83 230
rect 81 229 82 230
rect 80 229 81 230
rect 79 229 80 230
rect 78 229 79 230
rect 77 229 78 230
rect 76 229 77 230
rect 75 229 76 230
rect 74 229 75 230
rect 73 229 74 230
rect 72 229 73 230
rect 71 229 72 230
rect 70 229 71 230
rect 69 229 70 230
rect 68 229 69 230
rect 67 229 68 230
rect 66 229 67 230
rect 65 229 66 230
rect 64 229 65 230
rect 63 229 64 230
rect 62 229 63 230
rect 61 229 62 230
rect 60 229 61 230
rect 59 229 60 230
rect 58 229 59 230
rect 57 229 58 230
rect 56 229 57 230
rect 55 229 56 230
rect 54 229 55 230
rect 53 229 54 230
rect 52 229 53 230
rect 51 229 52 230
rect 50 229 51 230
rect 49 229 50 230
rect 48 229 49 230
rect 47 229 48 230
rect 46 229 47 230
rect 45 229 46 230
rect 44 229 45 230
rect 43 229 44 230
rect 42 229 43 230
rect 41 229 42 230
rect 40 229 41 230
rect 39 229 40 230
rect 38 229 39 230
rect 37 229 38 230
rect 36 229 37 230
rect 35 229 36 230
rect 34 229 35 230
rect 33 229 34 230
rect 32 229 33 230
rect 31 229 32 230
rect 30 229 31 230
rect 29 229 30 230
rect 28 229 29 230
rect 27 229 28 230
rect 26 229 27 230
rect 25 229 26 230
rect 24 229 25 230
rect 23 229 24 230
rect 22 229 23 230
rect 21 229 22 230
rect 20 229 21 230
rect 19 229 20 230
rect 18 229 19 230
rect 17 229 18 230
rect 16 229 17 230
rect 15 229 16 230
rect 14 229 15 230
rect 13 229 14 230
rect 12 229 13 230
rect 11 229 12 230
rect 10 229 11 230
rect 9 229 10 230
rect 8 229 9 230
rect 7 229 8 230
rect 6 229 7 230
rect 5 229 6 230
rect 4 229 5 230
rect 3 229 4 230
rect 478 230 479 231
rect 477 230 478 231
rect 476 230 477 231
rect 475 230 476 231
rect 474 230 475 231
rect 466 230 467 231
rect 465 230 466 231
rect 464 230 465 231
rect 463 230 464 231
rect 462 230 463 231
rect 461 230 462 231
rect 460 230 461 231
rect 438 230 439 231
rect 437 230 438 231
rect 436 230 437 231
rect 418 230 419 231
rect 417 230 418 231
rect 416 230 417 231
rect 394 230 395 231
rect 393 230 394 231
rect 392 230 393 231
rect 273 230 274 231
rect 272 230 273 231
rect 271 230 272 231
rect 270 230 271 231
rect 269 230 270 231
rect 268 230 269 231
rect 267 230 268 231
rect 266 230 267 231
rect 265 230 266 231
rect 264 230 265 231
rect 263 230 264 231
rect 262 230 263 231
rect 261 230 262 231
rect 260 230 261 231
rect 259 230 260 231
rect 258 230 259 231
rect 257 230 258 231
rect 256 230 257 231
rect 255 230 256 231
rect 254 230 255 231
rect 253 230 254 231
rect 252 230 253 231
rect 251 230 252 231
rect 250 230 251 231
rect 249 230 250 231
rect 248 230 249 231
rect 247 230 248 231
rect 246 230 247 231
rect 245 230 246 231
rect 244 230 245 231
rect 243 230 244 231
rect 242 230 243 231
rect 241 230 242 231
rect 240 230 241 231
rect 239 230 240 231
rect 238 230 239 231
rect 237 230 238 231
rect 236 230 237 231
rect 235 230 236 231
rect 234 230 235 231
rect 233 230 234 231
rect 232 230 233 231
rect 231 230 232 231
rect 230 230 231 231
rect 229 230 230 231
rect 228 230 229 231
rect 227 230 228 231
rect 226 230 227 231
rect 225 230 226 231
rect 224 230 225 231
rect 223 230 224 231
rect 222 230 223 231
rect 221 230 222 231
rect 220 230 221 231
rect 219 230 220 231
rect 218 230 219 231
rect 217 230 218 231
rect 216 230 217 231
rect 215 230 216 231
rect 214 230 215 231
rect 213 230 214 231
rect 212 230 213 231
rect 211 230 212 231
rect 210 230 211 231
rect 209 230 210 231
rect 208 230 209 231
rect 207 230 208 231
rect 206 230 207 231
rect 205 230 206 231
rect 204 230 205 231
rect 203 230 204 231
rect 202 230 203 231
rect 201 230 202 231
rect 200 230 201 231
rect 199 230 200 231
rect 198 230 199 231
rect 197 230 198 231
rect 196 230 197 231
rect 195 230 196 231
rect 194 230 195 231
rect 193 230 194 231
rect 192 230 193 231
rect 191 230 192 231
rect 190 230 191 231
rect 189 230 190 231
rect 188 230 189 231
rect 187 230 188 231
rect 186 230 187 231
rect 185 230 186 231
rect 184 230 185 231
rect 183 230 184 231
rect 182 230 183 231
rect 181 230 182 231
rect 180 230 181 231
rect 179 230 180 231
rect 178 230 179 231
rect 177 230 178 231
rect 176 230 177 231
rect 175 230 176 231
rect 174 230 175 231
rect 173 230 174 231
rect 172 230 173 231
rect 171 230 172 231
rect 170 230 171 231
rect 169 230 170 231
rect 168 230 169 231
rect 167 230 168 231
rect 166 230 167 231
rect 165 230 166 231
rect 164 230 165 231
rect 163 230 164 231
rect 143 230 144 231
rect 142 230 143 231
rect 141 230 142 231
rect 140 230 141 231
rect 139 230 140 231
rect 138 230 139 231
rect 137 230 138 231
rect 136 230 137 231
rect 135 230 136 231
rect 134 230 135 231
rect 133 230 134 231
rect 132 230 133 231
rect 131 230 132 231
rect 130 230 131 231
rect 129 230 130 231
rect 128 230 129 231
rect 127 230 128 231
rect 126 230 127 231
rect 125 230 126 231
rect 124 230 125 231
rect 123 230 124 231
rect 122 230 123 231
rect 121 230 122 231
rect 120 230 121 231
rect 119 230 120 231
rect 118 230 119 231
rect 117 230 118 231
rect 116 230 117 231
rect 115 230 116 231
rect 114 230 115 231
rect 113 230 114 231
rect 87 230 88 231
rect 86 230 87 231
rect 85 230 86 231
rect 84 230 85 231
rect 83 230 84 231
rect 82 230 83 231
rect 81 230 82 231
rect 80 230 81 231
rect 79 230 80 231
rect 78 230 79 231
rect 77 230 78 231
rect 76 230 77 231
rect 75 230 76 231
rect 74 230 75 231
rect 73 230 74 231
rect 72 230 73 231
rect 71 230 72 231
rect 70 230 71 231
rect 69 230 70 231
rect 68 230 69 231
rect 67 230 68 231
rect 66 230 67 231
rect 65 230 66 231
rect 64 230 65 231
rect 63 230 64 231
rect 62 230 63 231
rect 61 230 62 231
rect 60 230 61 231
rect 59 230 60 231
rect 58 230 59 231
rect 57 230 58 231
rect 56 230 57 231
rect 55 230 56 231
rect 54 230 55 231
rect 53 230 54 231
rect 52 230 53 231
rect 51 230 52 231
rect 50 230 51 231
rect 49 230 50 231
rect 48 230 49 231
rect 47 230 48 231
rect 46 230 47 231
rect 45 230 46 231
rect 44 230 45 231
rect 43 230 44 231
rect 42 230 43 231
rect 41 230 42 231
rect 40 230 41 231
rect 39 230 40 231
rect 38 230 39 231
rect 37 230 38 231
rect 36 230 37 231
rect 35 230 36 231
rect 34 230 35 231
rect 33 230 34 231
rect 32 230 33 231
rect 31 230 32 231
rect 30 230 31 231
rect 29 230 30 231
rect 28 230 29 231
rect 27 230 28 231
rect 26 230 27 231
rect 25 230 26 231
rect 24 230 25 231
rect 21 230 22 231
rect 20 230 21 231
rect 19 230 20 231
rect 18 230 19 231
rect 17 230 18 231
rect 16 230 17 231
rect 15 230 16 231
rect 14 230 15 231
rect 13 230 14 231
rect 12 230 13 231
rect 11 230 12 231
rect 10 230 11 231
rect 9 230 10 231
rect 8 230 9 231
rect 7 230 8 231
rect 6 230 7 231
rect 5 230 6 231
rect 4 230 5 231
rect 3 230 4 231
rect 2 230 3 231
rect 479 231 480 232
rect 478 231 479 232
rect 477 231 478 232
rect 476 231 477 232
rect 438 231 439 232
rect 437 231 438 232
rect 436 231 437 232
rect 418 231 419 232
rect 417 231 418 232
rect 416 231 417 232
rect 394 231 395 232
rect 393 231 394 232
rect 392 231 393 232
rect 272 231 273 232
rect 271 231 272 232
rect 270 231 271 232
rect 269 231 270 232
rect 268 231 269 232
rect 267 231 268 232
rect 266 231 267 232
rect 265 231 266 232
rect 264 231 265 232
rect 263 231 264 232
rect 262 231 263 232
rect 261 231 262 232
rect 260 231 261 232
rect 259 231 260 232
rect 258 231 259 232
rect 257 231 258 232
rect 256 231 257 232
rect 255 231 256 232
rect 254 231 255 232
rect 253 231 254 232
rect 252 231 253 232
rect 251 231 252 232
rect 250 231 251 232
rect 249 231 250 232
rect 248 231 249 232
rect 247 231 248 232
rect 246 231 247 232
rect 245 231 246 232
rect 244 231 245 232
rect 243 231 244 232
rect 242 231 243 232
rect 241 231 242 232
rect 240 231 241 232
rect 239 231 240 232
rect 238 231 239 232
rect 237 231 238 232
rect 236 231 237 232
rect 235 231 236 232
rect 234 231 235 232
rect 233 231 234 232
rect 232 231 233 232
rect 231 231 232 232
rect 230 231 231 232
rect 229 231 230 232
rect 228 231 229 232
rect 227 231 228 232
rect 226 231 227 232
rect 225 231 226 232
rect 224 231 225 232
rect 223 231 224 232
rect 222 231 223 232
rect 221 231 222 232
rect 220 231 221 232
rect 219 231 220 232
rect 218 231 219 232
rect 217 231 218 232
rect 216 231 217 232
rect 215 231 216 232
rect 214 231 215 232
rect 213 231 214 232
rect 212 231 213 232
rect 211 231 212 232
rect 210 231 211 232
rect 209 231 210 232
rect 208 231 209 232
rect 207 231 208 232
rect 206 231 207 232
rect 205 231 206 232
rect 204 231 205 232
rect 203 231 204 232
rect 202 231 203 232
rect 201 231 202 232
rect 200 231 201 232
rect 199 231 200 232
rect 198 231 199 232
rect 197 231 198 232
rect 196 231 197 232
rect 195 231 196 232
rect 194 231 195 232
rect 193 231 194 232
rect 192 231 193 232
rect 191 231 192 232
rect 190 231 191 232
rect 189 231 190 232
rect 188 231 189 232
rect 187 231 188 232
rect 186 231 187 232
rect 185 231 186 232
rect 184 231 185 232
rect 183 231 184 232
rect 182 231 183 232
rect 181 231 182 232
rect 180 231 181 232
rect 179 231 180 232
rect 178 231 179 232
rect 177 231 178 232
rect 176 231 177 232
rect 175 231 176 232
rect 174 231 175 232
rect 173 231 174 232
rect 172 231 173 232
rect 171 231 172 232
rect 170 231 171 232
rect 169 231 170 232
rect 168 231 169 232
rect 167 231 168 232
rect 166 231 167 232
rect 165 231 166 232
rect 143 231 144 232
rect 142 231 143 232
rect 141 231 142 232
rect 140 231 141 232
rect 139 231 140 232
rect 138 231 139 232
rect 137 231 138 232
rect 136 231 137 232
rect 135 231 136 232
rect 134 231 135 232
rect 133 231 134 232
rect 132 231 133 232
rect 131 231 132 232
rect 130 231 131 232
rect 129 231 130 232
rect 128 231 129 232
rect 127 231 128 232
rect 126 231 127 232
rect 125 231 126 232
rect 124 231 125 232
rect 123 231 124 232
rect 122 231 123 232
rect 121 231 122 232
rect 120 231 121 232
rect 119 231 120 232
rect 118 231 119 232
rect 117 231 118 232
rect 116 231 117 232
rect 115 231 116 232
rect 114 231 115 232
rect 90 231 91 232
rect 89 231 90 232
rect 88 231 89 232
rect 87 231 88 232
rect 86 231 87 232
rect 85 231 86 232
rect 84 231 85 232
rect 83 231 84 232
rect 82 231 83 232
rect 81 231 82 232
rect 80 231 81 232
rect 79 231 80 232
rect 78 231 79 232
rect 77 231 78 232
rect 76 231 77 232
rect 75 231 76 232
rect 74 231 75 232
rect 73 231 74 232
rect 72 231 73 232
rect 71 231 72 232
rect 70 231 71 232
rect 69 231 70 232
rect 68 231 69 232
rect 67 231 68 232
rect 66 231 67 232
rect 65 231 66 232
rect 64 231 65 232
rect 63 231 64 232
rect 62 231 63 232
rect 61 231 62 232
rect 60 231 61 232
rect 59 231 60 232
rect 58 231 59 232
rect 57 231 58 232
rect 56 231 57 232
rect 55 231 56 232
rect 54 231 55 232
rect 53 231 54 232
rect 52 231 53 232
rect 51 231 52 232
rect 50 231 51 232
rect 49 231 50 232
rect 48 231 49 232
rect 47 231 48 232
rect 46 231 47 232
rect 45 231 46 232
rect 44 231 45 232
rect 43 231 44 232
rect 42 231 43 232
rect 41 231 42 232
rect 40 231 41 232
rect 39 231 40 232
rect 38 231 39 232
rect 37 231 38 232
rect 36 231 37 232
rect 35 231 36 232
rect 34 231 35 232
rect 33 231 34 232
rect 32 231 33 232
rect 31 231 32 232
rect 30 231 31 232
rect 29 231 30 232
rect 28 231 29 232
rect 27 231 28 232
rect 26 231 27 232
rect 25 231 26 232
rect 24 231 25 232
rect 20 231 21 232
rect 19 231 20 232
rect 18 231 19 232
rect 17 231 18 232
rect 16 231 17 232
rect 15 231 16 232
rect 14 231 15 232
rect 13 231 14 232
rect 12 231 13 232
rect 11 231 12 232
rect 10 231 11 232
rect 9 231 10 232
rect 8 231 9 232
rect 7 231 8 232
rect 6 231 7 232
rect 5 231 6 232
rect 4 231 5 232
rect 3 231 4 232
rect 2 231 3 232
rect 479 232 480 233
rect 478 232 479 233
rect 477 232 478 233
rect 438 232 439 233
rect 437 232 438 233
rect 436 232 437 233
rect 418 232 419 233
rect 417 232 418 233
rect 416 232 417 233
rect 394 232 395 233
rect 393 232 394 233
rect 392 232 393 233
rect 271 232 272 233
rect 270 232 271 233
rect 269 232 270 233
rect 268 232 269 233
rect 267 232 268 233
rect 266 232 267 233
rect 265 232 266 233
rect 264 232 265 233
rect 263 232 264 233
rect 262 232 263 233
rect 261 232 262 233
rect 260 232 261 233
rect 259 232 260 233
rect 258 232 259 233
rect 257 232 258 233
rect 256 232 257 233
rect 255 232 256 233
rect 254 232 255 233
rect 253 232 254 233
rect 252 232 253 233
rect 251 232 252 233
rect 250 232 251 233
rect 249 232 250 233
rect 248 232 249 233
rect 247 232 248 233
rect 246 232 247 233
rect 245 232 246 233
rect 244 232 245 233
rect 243 232 244 233
rect 242 232 243 233
rect 241 232 242 233
rect 240 232 241 233
rect 239 232 240 233
rect 238 232 239 233
rect 237 232 238 233
rect 236 232 237 233
rect 235 232 236 233
rect 234 232 235 233
rect 233 232 234 233
rect 232 232 233 233
rect 231 232 232 233
rect 230 232 231 233
rect 229 232 230 233
rect 228 232 229 233
rect 227 232 228 233
rect 226 232 227 233
rect 225 232 226 233
rect 224 232 225 233
rect 223 232 224 233
rect 222 232 223 233
rect 221 232 222 233
rect 220 232 221 233
rect 219 232 220 233
rect 218 232 219 233
rect 217 232 218 233
rect 216 232 217 233
rect 215 232 216 233
rect 214 232 215 233
rect 213 232 214 233
rect 212 232 213 233
rect 211 232 212 233
rect 210 232 211 233
rect 209 232 210 233
rect 208 232 209 233
rect 207 232 208 233
rect 206 232 207 233
rect 205 232 206 233
rect 204 232 205 233
rect 203 232 204 233
rect 202 232 203 233
rect 201 232 202 233
rect 200 232 201 233
rect 199 232 200 233
rect 198 232 199 233
rect 197 232 198 233
rect 196 232 197 233
rect 195 232 196 233
rect 194 232 195 233
rect 193 232 194 233
rect 192 232 193 233
rect 191 232 192 233
rect 190 232 191 233
rect 189 232 190 233
rect 188 232 189 233
rect 187 232 188 233
rect 186 232 187 233
rect 185 232 186 233
rect 184 232 185 233
rect 183 232 184 233
rect 182 232 183 233
rect 181 232 182 233
rect 180 232 181 233
rect 179 232 180 233
rect 178 232 179 233
rect 177 232 178 233
rect 176 232 177 233
rect 175 232 176 233
rect 174 232 175 233
rect 173 232 174 233
rect 172 232 173 233
rect 171 232 172 233
rect 170 232 171 233
rect 169 232 170 233
rect 168 232 169 233
rect 167 232 168 233
rect 166 232 167 233
rect 144 232 145 233
rect 143 232 144 233
rect 142 232 143 233
rect 141 232 142 233
rect 140 232 141 233
rect 139 232 140 233
rect 138 232 139 233
rect 137 232 138 233
rect 136 232 137 233
rect 135 232 136 233
rect 134 232 135 233
rect 133 232 134 233
rect 132 232 133 233
rect 131 232 132 233
rect 130 232 131 233
rect 129 232 130 233
rect 128 232 129 233
rect 127 232 128 233
rect 126 232 127 233
rect 125 232 126 233
rect 124 232 125 233
rect 123 232 124 233
rect 122 232 123 233
rect 121 232 122 233
rect 120 232 121 233
rect 119 232 120 233
rect 118 232 119 233
rect 117 232 118 233
rect 116 232 117 233
rect 115 232 116 233
rect 114 232 115 233
rect 92 232 93 233
rect 91 232 92 233
rect 90 232 91 233
rect 89 232 90 233
rect 88 232 89 233
rect 87 232 88 233
rect 86 232 87 233
rect 85 232 86 233
rect 84 232 85 233
rect 83 232 84 233
rect 82 232 83 233
rect 81 232 82 233
rect 80 232 81 233
rect 79 232 80 233
rect 78 232 79 233
rect 77 232 78 233
rect 76 232 77 233
rect 75 232 76 233
rect 74 232 75 233
rect 73 232 74 233
rect 72 232 73 233
rect 71 232 72 233
rect 70 232 71 233
rect 69 232 70 233
rect 68 232 69 233
rect 67 232 68 233
rect 66 232 67 233
rect 65 232 66 233
rect 64 232 65 233
rect 63 232 64 233
rect 62 232 63 233
rect 61 232 62 233
rect 60 232 61 233
rect 59 232 60 233
rect 58 232 59 233
rect 57 232 58 233
rect 56 232 57 233
rect 55 232 56 233
rect 54 232 55 233
rect 53 232 54 233
rect 52 232 53 233
rect 51 232 52 233
rect 50 232 51 233
rect 49 232 50 233
rect 48 232 49 233
rect 47 232 48 233
rect 46 232 47 233
rect 45 232 46 233
rect 44 232 45 233
rect 43 232 44 233
rect 42 232 43 233
rect 41 232 42 233
rect 40 232 41 233
rect 39 232 40 233
rect 38 232 39 233
rect 37 232 38 233
rect 36 232 37 233
rect 35 232 36 233
rect 34 232 35 233
rect 33 232 34 233
rect 32 232 33 233
rect 31 232 32 233
rect 30 232 31 233
rect 29 232 30 233
rect 28 232 29 233
rect 27 232 28 233
rect 26 232 27 233
rect 25 232 26 233
rect 20 232 21 233
rect 19 232 20 233
rect 18 232 19 233
rect 17 232 18 233
rect 16 232 17 233
rect 15 232 16 233
rect 14 232 15 233
rect 13 232 14 233
rect 12 232 13 233
rect 11 232 12 233
rect 10 232 11 233
rect 9 232 10 233
rect 8 232 9 233
rect 7 232 8 233
rect 6 232 7 233
rect 5 232 6 233
rect 4 232 5 233
rect 3 232 4 233
rect 2 232 3 233
rect 479 233 480 234
rect 478 233 479 234
rect 438 233 439 234
rect 437 233 438 234
rect 436 233 437 234
rect 419 233 420 234
rect 418 233 419 234
rect 417 233 418 234
rect 416 233 417 234
rect 394 233 395 234
rect 393 233 394 234
rect 392 233 393 234
rect 270 233 271 234
rect 269 233 270 234
rect 268 233 269 234
rect 267 233 268 234
rect 266 233 267 234
rect 265 233 266 234
rect 264 233 265 234
rect 263 233 264 234
rect 262 233 263 234
rect 261 233 262 234
rect 260 233 261 234
rect 259 233 260 234
rect 258 233 259 234
rect 257 233 258 234
rect 256 233 257 234
rect 255 233 256 234
rect 254 233 255 234
rect 253 233 254 234
rect 252 233 253 234
rect 251 233 252 234
rect 250 233 251 234
rect 249 233 250 234
rect 248 233 249 234
rect 247 233 248 234
rect 246 233 247 234
rect 245 233 246 234
rect 244 233 245 234
rect 243 233 244 234
rect 242 233 243 234
rect 241 233 242 234
rect 240 233 241 234
rect 239 233 240 234
rect 238 233 239 234
rect 237 233 238 234
rect 236 233 237 234
rect 235 233 236 234
rect 234 233 235 234
rect 233 233 234 234
rect 232 233 233 234
rect 231 233 232 234
rect 230 233 231 234
rect 229 233 230 234
rect 228 233 229 234
rect 227 233 228 234
rect 226 233 227 234
rect 225 233 226 234
rect 224 233 225 234
rect 223 233 224 234
rect 222 233 223 234
rect 221 233 222 234
rect 220 233 221 234
rect 219 233 220 234
rect 218 233 219 234
rect 217 233 218 234
rect 216 233 217 234
rect 215 233 216 234
rect 214 233 215 234
rect 213 233 214 234
rect 212 233 213 234
rect 211 233 212 234
rect 210 233 211 234
rect 209 233 210 234
rect 208 233 209 234
rect 207 233 208 234
rect 206 233 207 234
rect 205 233 206 234
rect 204 233 205 234
rect 203 233 204 234
rect 202 233 203 234
rect 201 233 202 234
rect 200 233 201 234
rect 199 233 200 234
rect 198 233 199 234
rect 197 233 198 234
rect 196 233 197 234
rect 195 233 196 234
rect 194 233 195 234
rect 193 233 194 234
rect 192 233 193 234
rect 191 233 192 234
rect 190 233 191 234
rect 189 233 190 234
rect 188 233 189 234
rect 187 233 188 234
rect 186 233 187 234
rect 185 233 186 234
rect 184 233 185 234
rect 183 233 184 234
rect 182 233 183 234
rect 181 233 182 234
rect 180 233 181 234
rect 179 233 180 234
rect 178 233 179 234
rect 177 233 178 234
rect 176 233 177 234
rect 175 233 176 234
rect 174 233 175 234
rect 173 233 174 234
rect 172 233 173 234
rect 171 233 172 234
rect 170 233 171 234
rect 169 233 170 234
rect 168 233 169 234
rect 144 233 145 234
rect 143 233 144 234
rect 142 233 143 234
rect 141 233 142 234
rect 140 233 141 234
rect 139 233 140 234
rect 138 233 139 234
rect 137 233 138 234
rect 136 233 137 234
rect 135 233 136 234
rect 134 233 135 234
rect 133 233 134 234
rect 132 233 133 234
rect 131 233 132 234
rect 130 233 131 234
rect 129 233 130 234
rect 128 233 129 234
rect 127 233 128 234
rect 126 233 127 234
rect 125 233 126 234
rect 124 233 125 234
rect 123 233 124 234
rect 122 233 123 234
rect 121 233 122 234
rect 120 233 121 234
rect 119 233 120 234
rect 118 233 119 234
rect 117 233 118 234
rect 116 233 117 234
rect 115 233 116 234
rect 94 233 95 234
rect 93 233 94 234
rect 92 233 93 234
rect 91 233 92 234
rect 90 233 91 234
rect 89 233 90 234
rect 88 233 89 234
rect 87 233 88 234
rect 86 233 87 234
rect 85 233 86 234
rect 84 233 85 234
rect 83 233 84 234
rect 82 233 83 234
rect 81 233 82 234
rect 80 233 81 234
rect 79 233 80 234
rect 78 233 79 234
rect 77 233 78 234
rect 76 233 77 234
rect 75 233 76 234
rect 74 233 75 234
rect 73 233 74 234
rect 72 233 73 234
rect 71 233 72 234
rect 70 233 71 234
rect 69 233 70 234
rect 68 233 69 234
rect 67 233 68 234
rect 66 233 67 234
rect 65 233 66 234
rect 64 233 65 234
rect 63 233 64 234
rect 62 233 63 234
rect 61 233 62 234
rect 60 233 61 234
rect 59 233 60 234
rect 58 233 59 234
rect 57 233 58 234
rect 56 233 57 234
rect 55 233 56 234
rect 54 233 55 234
rect 53 233 54 234
rect 52 233 53 234
rect 51 233 52 234
rect 50 233 51 234
rect 49 233 50 234
rect 48 233 49 234
rect 47 233 48 234
rect 46 233 47 234
rect 45 233 46 234
rect 44 233 45 234
rect 43 233 44 234
rect 42 233 43 234
rect 41 233 42 234
rect 40 233 41 234
rect 39 233 40 234
rect 38 233 39 234
rect 37 233 38 234
rect 36 233 37 234
rect 35 233 36 234
rect 34 233 35 234
rect 33 233 34 234
rect 32 233 33 234
rect 31 233 32 234
rect 30 233 31 234
rect 29 233 30 234
rect 28 233 29 234
rect 27 233 28 234
rect 26 233 27 234
rect 25 233 26 234
rect 20 233 21 234
rect 19 233 20 234
rect 18 233 19 234
rect 17 233 18 234
rect 16 233 17 234
rect 15 233 16 234
rect 14 233 15 234
rect 13 233 14 234
rect 12 233 13 234
rect 11 233 12 234
rect 10 233 11 234
rect 9 233 10 234
rect 8 233 9 234
rect 7 233 8 234
rect 6 233 7 234
rect 5 233 6 234
rect 4 233 5 234
rect 3 233 4 234
rect 2 233 3 234
rect 438 234 439 235
rect 437 234 438 235
rect 436 234 437 235
rect 419 234 420 235
rect 418 234 419 235
rect 417 234 418 235
rect 416 234 417 235
rect 394 234 395 235
rect 393 234 394 235
rect 392 234 393 235
rect 269 234 270 235
rect 268 234 269 235
rect 267 234 268 235
rect 266 234 267 235
rect 265 234 266 235
rect 264 234 265 235
rect 263 234 264 235
rect 262 234 263 235
rect 261 234 262 235
rect 260 234 261 235
rect 259 234 260 235
rect 258 234 259 235
rect 257 234 258 235
rect 256 234 257 235
rect 255 234 256 235
rect 254 234 255 235
rect 253 234 254 235
rect 252 234 253 235
rect 251 234 252 235
rect 250 234 251 235
rect 249 234 250 235
rect 248 234 249 235
rect 247 234 248 235
rect 246 234 247 235
rect 245 234 246 235
rect 244 234 245 235
rect 243 234 244 235
rect 242 234 243 235
rect 241 234 242 235
rect 240 234 241 235
rect 239 234 240 235
rect 238 234 239 235
rect 237 234 238 235
rect 236 234 237 235
rect 235 234 236 235
rect 234 234 235 235
rect 233 234 234 235
rect 232 234 233 235
rect 231 234 232 235
rect 230 234 231 235
rect 229 234 230 235
rect 228 234 229 235
rect 227 234 228 235
rect 226 234 227 235
rect 225 234 226 235
rect 224 234 225 235
rect 223 234 224 235
rect 222 234 223 235
rect 221 234 222 235
rect 220 234 221 235
rect 219 234 220 235
rect 218 234 219 235
rect 217 234 218 235
rect 216 234 217 235
rect 215 234 216 235
rect 214 234 215 235
rect 213 234 214 235
rect 212 234 213 235
rect 211 234 212 235
rect 210 234 211 235
rect 209 234 210 235
rect 208 234 209 235
rect 207 234 208 235
rect 206 234 207 235
rect 205 234 206 235
rect 204 234 205 235
rect 203 234 204 235
rect 202 234 203 235
rect 201 234 202 235
rect 200 234 201 235
rect 199 234 200 235
rect 198 234 199 235
rect 197 234 198 235
rect 196 234 197 235
rect 195 234 196 235
rect 194 234 195 235
rect 193 234 194 235
rect 192 234 193 235
rect 191 234 192 235
rect 190 234 191 235
rect 189 234 190 235
rect 188 234 189 235
rect 187 234 188 235
rect 186 234 187 235
rect 185 234 186 235
rect 184 234 185 235
rect 183 234 184 235
rect 182 234 183 235
rect 181 234 182 235
rect 180 234 181 235
rect 179 234 180 235
rect 178 234 179 235
rect 177 234 178 235
rect 176 234 177 235
rect 175 234 176 235
rect 174 234 175 235
rect 173 234 174 235
rect 172 234 173 235
rect 171 234 172 235
rect 170 234 171 235
rect 169 234 170 235
rect 145 234 146 235
rect 144 234 145 235
rect 143 234 144 235
rect 142 234 143 235
rect 141 234 142 235
rect 140 234 141 235
rect 139 234 140 235
rect 138 234 139 235
rect 137 234 138 235
rect 136 234 137 235
rect 135 234 136 235
rect 134 234 135 235
rect 133 234 134 235
rect 132 234 133 235
rect 131 234 132 235
rect 130 234 131 235
rect 129 234 130 235
rect 128 234 129 235
rect 127 234 128 235
rect 126 234 127 235
rect 125 234 126 235
rect 124 234 125 235
rect 123 234 124 235
rect 122 234 123 235
rect 121 234 122 235
rect 120 234 121 235
rect 119 234 120 235
rect 118 234 119 235
rect 117 234 118 235
rect 116 234 117 235
rect 115 234 116 235
rect 95 234 96 235
rect 94 234 95 235
rect 93 234 94 235
rect 92 234 93 235
rect 91 234 92 235
rect 90 234 91 235
rect 89 234 90 235
rect 88 234 89 235
rect 87 234 88 235
rect 86 234 87 235
rect 85 234 86 235
rect 84 234 85 235
rect 83 234 84 235
rect 82 234 83 235
rect 81 234 82 235
rect 80 234 81 235
rect 79 234 80 235
rect 78 234 79 235
rect 77 234 78 235
rect 76 234 77 235
rect 75 234 76 235
rect 74 234 75 235
rect 73 234 74 235
rect 72 234 73 235
rect 71 234 72 235
rect 70 234 71 235
rect 69 234 70 235
rect 68 234 69 235
rect 67 234 68 235
rect 66 234 67 235
rect 65 234 66 235
rect 64 234 65 235
rect 63 234 64 235
rect 62 234 63 235
rect 61 234 62 235
rect 60 234 61 235
rect 59 234 60 235
rect 58 234 59 235
rect 57 234 58 235
rect 56 234 57 235
rect 55 234 56 235
rect 54 234 55 235
rect 53 234 54 235
rect 52 234 53 235
rect 51 234 52 235
rect 50 234 51 235
rect 49 234 50 235
rect 48 234 49 235
rect 47 234 48 235
rect 46 234 47 235
rect 45 234 46 235
rect 44 234 45 235
rect 43 234 44 235
rect 42 234 43 235
rect 41 234 42 235
rect 40 234 41 235
rect 39 234 40 235
rect 38 234 39 235
rect 37 234 38 235
rect 36 234 37 235
rect 35 234 36 235
rect 34 234 35 235
rect 33 234 34 235
rect 32 234 33 235
rect 31 234 32 235
rect 30 234 31 235
rect 29 234 30 235
rect 28 234 29 235
rect 27 234 28 235
rect 26 234 27 235
rect 25 234 26 235
rect 19 234 20 235
rect 18 234 19 235
rect 17 234 18 235
rect 16 234 17 235
rect 15 234 16 235
rect 14 234 15 235
rect 13 234 14 235
rect 12 234 13 235
rect 11 234 12 235
rect 10 234 11 235
rect 9 234 10 235
rect 8 234 9 235
rect 7 234 8 235
rect 6 234 7 235
rect 5 234 6 235
rect 4 234 5 235
rect 3 234 4 235
rect 2 234 3 235
rect 438 235 439 236
rect 437 235 438 236
rect 436 235 437 236
rect 419 235 420 236
rect 418 235 419 236
rect 417 235 418 236
rect 416 235 417 236
rect 395 235 396 236
rect 394 235 395 236
rect 393 235 394 236
rect 392 235 393 236
rect 269 235 270 236
rect 268 235 269 236
rect 267 235 268 236
rect 266 235 267 236
rect 265 235 266 236
rect 264 235 265 236
rect 263 235 264 236
rect 262 235 263 236
rect 261 235 262 236
rect 260 235 261 236
rect 259 235 260 236
rect 258 235 259 236
rect 257 235 258 236
rect 256 235 257 236
rect 255 235 256 236
rect 254 235 255 236
rect 253 235 254 236
rect 252 235 253 236
rect 251 235 252 236
rect 250 235 251 236
rect 249 235 250 236
rect 248 235 249 236
rect 247 235 248 236
rect 246 235 247 236
rect 245 235 246 236
rect 244 235 245 236
rect 243 235 244 236
rect 242 235 243 236
rect 241 235 242 236
rect 240 235 241 236
rect 239 235 240 236
rect 238 235 239 236
rect 237 235 238 236
rect 236 235 237 236
rect 235 235 236 236
rect 234 235 235 236
rect 233 235 234 236
rect 232 235 233 236
rect 231 235 232 236
rect 230 235 231 236
rect 229 235 230 236
rect 228 235 229 236
rect 227 235 228 236
rect 226 235 227 236
rect 225 235 226 236
rect 224 235 225 236
rect 223 235 224 236
rect 222 235 223 236
rect 221 235 222 236
rect 220 235 221 236
rect 219 235 220 236
rect 218 235 219 236
rect 217 235 218 236
rect 216 235 217 236
rect 215 235 216 236
rect 214 235 215 236
rect 213 235 214 236
rect 212 235 213 236
rect 211 235 212 236
rect 210 235 211 236
rect 209 235 210 236
rect 208 235 209 236
rect 207 235 208 236
rect 206 235 207 236
rect 205 235 206 236
rect 204 235 205 236
rect 203 235 204 236
rect 202 235 203 236
rect 201 235 202 236
rect 200 235 201 236
rect 199 235 200 236
rect 198 235 199 236
rect 197 235 198 236
rect 196 235 197 236
rect 195 235 196 236
rect 194 235 195 236
rect 193 235 194 236
rect 192 235 193 236
rect 191 235 192 236
rect 190 235 191 236
rect 189 235 190 236
rect 188 235 189 236
rect 187 235 188 236
rect 186 235 187 236
rect 185 235 186 236
rect 184 235 185 236
rect 183 235 184 236
rect 182 235 183 236
rect 181 235 182 236
rect 180 235 181 236
rect 179 235 180 236
rect 178 235 179 236
rect 177 235 178 236
rect 176 235 177 236
rect 175 235 176 236
rect 174 235 175 236
rect 173 235 174 236
rect 172 235 173 236
rect 171 235 172 236
rect 145 235 146 236
rect 144 235 145 236
rect 143 235 144 236
rect 142 235 143 236
rect 141 235 142 236
rect 140 235 141 236
rect 139 235 140 236
rect 138 235 139 236
rect 137 235 138 236
rect 136 235 137 236
rect 135 235 136 236
rect 134 235 135 236
rect 133 235 134 236
rect 132 235 133 236
rect 131 235 132 236
rect 130 235 131 236
rect 129 235 130 236
rect 128 235 129 236
rect 127 235 128 236
rect 126 235 127 236
rect 125 235 126 236
rect 124 235 125 236
rect 123 235 124 236
rect 122 235 123 236
rect 121 235 122 236
rect 120 235 121 236
rect 119 235 120 236
rect 118 235 119 236
rect 117 235 118 236
rect 116 235 117 236
rect 115 235 116 236
rect 97 235 98 236
rect 96 235 97 236
rect 95 235 96 236
rect 94 235 95 236
rect 93 235 94 236
rect 92 235 93 236
rect 91 235 92 236
rect 90 235 91 236
rect 89 235 90 236
rect 88 235 89 236
rect 87 235 88 236
rect 86 235 87 236
rect 85 235 86 236
rect 84 235 85 236
rect 83 235 84 236
rect 82 235 83 236
rect 81 235 82 236
rect 80 235 81 236
rect 79 235 80 236
rect 78 235 79 236
rect 77 235 78 236
rect 76 235 77 236
rect 75 235 76 236
rect 74 235 75 236
rect 73 235 74 236
rect 72 235 73 236
rect 71 235 72 236
rect 70 235 71 236
rect 69 235 70 236
rect 68 235 69 236
rect 67 235 68 236
rect 66 235 67 236
rect 65 235 66 236
rect 64 235 65 236
rect 63 235 64 236
rect 62 235 63 236
rect 61 235 62 236
rect 60 235 61 236
rect 59 235 60 236
rect 58 235 59 236
rect 57 235 58 236
rect 56 235 57 236
rect 55 235 56 236
rect 54 235 55 236
rect 53 235 54 236
rect 52 235 53 236
rect 51 235 52 236
rect 50 235 51 236
rect 49 235 50 236
rect 48 235 49 236
rect 47 235 48 236
rect 46 235 47 236
rect 45 235 46 236
rect 44 235 45 236
rect 43 235 44 236
rect 42 235 43 236
rect 41 235 42 236
rect 40 235 41 236
rect 39 235 40 236
rect 38 235 39 236
rect 37 235 38 236
rect 36 235 37 236
rect 35 235 36 236
rect 34 235 35 236
rect 33 235 34 236
rect 32 235 33 236
rect 31 235 32 236
rect 30 235 31 236
rect 29 235 30 236
rect 28 235 29 236
rect 27 235 28 236
rect 26 235 27 236
rect 25 235 26 236
rect 19 235 20 236
rect 18 235 19 236
rect 17 235 18 236
rect 16 235 17 236
rect 15 235 16 236
rect 14 235 15 236
rect 13 235 14 236
rect 12 235 13 236
rect 11 235 12 236
rect 10 235 11 236
rect 9 235 10 236
rect 8 235 9 236
rect 7 235 8 236
rect 6 235 7 236
rect 5 235 6 236
rect 4 235 5 236
rect 3 235 4 236
rect 2 235 3 236
rect 438 236 439 237
rect 437 236 438 237
rect 436 236 437 237
rect 435 236 436 237
rect 420 236 421 237
rect 419 236 420 237
rect 418 236 419 237
rect 417 236 418 237
rect 416 236 417 237
rect 395 236 396 237
rect 394 236 395 237
rect 393 236 394 237
rect 392 236 393 237
rect 268 236 269 237
rect 267 236 268 237
rect 266 236 267 237
rect 265 236 266 237
rect 264 236 265 237
rect 263 236 264 237
rect 262 236 263 237
rect 261 236 262 237
rect 260 236 261 237
rect 259 236 260 237
rect 258 236 259 237
rect 257 236 258 237
rect 256 236 257 237
rect 255 236 256 237
rect 254 236 255 237
rect 253 236 254 237
rect 252 236 253 237
rect 251 236 252 237
rect 250 236 251 237
rect 249 236 250 237
rect 248 236 249 237
rect 247 236 248 237
rect 246 236 247 237
rect 245 236 246 237
rect 244 236 245 237
rect 243 236 244 237
rect 242 236 243 237
rect 241 236 242 237
rect 240 236 241 237
rect 239 236 240 237
rect 238 236 239 237
rect 237 236 238 237
rect 236 236 237 237
rect 235 236 236 237
rect 234 236 235 237
rect 233 236 234 237
rect 232 236 233 237
rect 231 236 232 237
rect 230 236 231 237
rect 229 236 230 237
rect 228 236 229 237
rect 227 236 228 237
rect 226 236 227 237
rect 225 236 226 237
rect 224 236 225 237
rect 223 236 224 237
rect 222 236 223 237
rect 221 236 222 237
rect 220 236 221 237
rect 219 236 220 237
rect 218 236 219 237
rect 217 236 218 237
rect 216 236 217 237
rect 215 236 216 237
rect 214 236 215 237
rect 213 236 214 237
rect 212 236 213 237
rect 211 236 212 237
rect 210 236 211 237
rect 209 236 210 237
rect 208 236 209 237
rect 207 236 208 237
rect 206 236 207 237
rect 205 236 206 237
rect 204 236 205 237
rect 203 236 204 237
rect 202 236 203 237
rect 201 236 202 237
rect 200 236 201 237
rect 199 236 200 237
rect 198 236 199 237
rect 197 236 198 237
rect 196 236 197 237
rect 195 236 196 237
rect 194 236 195 237
rect 193 236 194 237
rect 192 236 193 237
rect 191 236 192 237
rect 190 236 191 237
rect 189 236 190 237
rect 188 236 189 237
rect 187 236 188 237
rect 186 236 187 237
rect 185 236 186 237
rect 184 236 185 237
rect 183 236 184 237
rect 182 236 183 237
rect 181 236 182 237
rect 180 236 181 237
rect 179 236 180 237
rect 178 236 179 237
rect 177 236 178 237
rect 176 236 177 237
rect 175 236 176 237
rect 174 236 175 237
rect 173 236 174 237
rect 146 236 147 237
rect 145 236 146 237
rect 144 236 145 237
rect 143 236 144 237
rect 142 236 143 237
rect 141 236 142 237
rect 140 236 141 237
rect 139 236 140 237
rect 138 236 139 237
rect 137 236 138 237
rect 136 236 137 237
rect 135 236 136 237
rect 134 236 135 237
rect 133 236 134 237
rect 132 236 133 237
rect 131 236 132 237
rect 130 236 131 237
rect 129 236 130 237
rect 128 236 129 237
rect 127 236 128 237
rect 126 236 127 237
rect 125 236 126 237
rect 124 236 125 237
rect 123 236 124 237
rect 122 236 123 237
rect 121 236 122 237
rect 120 236 121 237
rect 119 236 120 237
rect 118 236 119 237
rect 117 236 118 237
rect 116 236 117 237
rect 98 236 99 237
rect 97 236 98 237
rect 96 236 97 237
rect 95 236 96 237
rect 94 236 95 237
rect 93 236 94 237
rect 92 236 93 237
rect 91 236 92 237
rect 90 236 91 237
rect 89 236 90 237
rect 88 236 89 237
rect 87 236 88 237
rect 86 236 87 237
rect 85 236 86 237
rect 84 236 85 237
rect 83 236 84 237
rect 82 236 83 237
rect 81 236 82 237
rect 80 236 81 237
rect 79 236 80 237
rect 78 236 79 237
rect 77 236 78 237
rect 76 236 77 237
rect 75 236 76 237
rect 74 236 75 237
rect 73 236 74 237
rect 72 236 73 237
rect 71 236 72 237
rect 70 236 71 237
rect 69 236 70 237
rect 68 236 69 237
rect 67 236 68 237
rect 66 236 67 237
rect 65 236 66 237
rect 64 236 65 237
rect 63 236 64 237
rect 62 236 63 237
rect 61 236 62 237
rect 60 236 61 237
rect 59 236 60 237
rect 58 236 59 237
rect 57 236 58 237
rect 56 236 57 237
rect 55 236 56 237
rect 54 236 55 237
rect 53 236 54 237
rect 52 236 53 237
rect 51 236 52 237
rect 50 236 51 237
rect 49 236 50 237
rect 48 236 49 237
rect 47 236 48 237
rect 46 236 47 237
rect 45 236 46 237
rect 44 236 45 237
rect 43 236 44 237
rect 42 236 43 237
rect 41 236 42 237
rect 40 236 41 237
rect 39 236 40 237
rect 38 236 39 237
rect 37 236 38 237
rect 36 236 37 237
rect 35 236 36 237
rect 34 236 35 237
rect 33 236 34 237
rect 32 236 33 237
rect 31 236 32 237
rect 30 236 31 237
rect 29 236 30 237
rect 28 236 29 237
rect 27 236 28 237
rect 26 236 27 237
rect 25 236 26 237
rect 19 236 20 237
rect 18 236 19 237
rect 17 236 18 237
rect 16 236 17 237
rect 15 236 16 237
rect 14 236 15 237
rect 13 236 14 237
rect 12 236 13 237
rect 11 236 12 237
rect 10 236 11 237
rect 9 236 10 237
rect 8 236 9 237
rect 7 236 8 237
rect 6 236 7 237
rect 5 236 6 237
rect 4 236 5 237
rect 3 236 4 237
rect 2 236 3 237
rect 438 237 439 238
rect 437 237 438 238
rect 436 237 437 238
rect 435 237 436 238
rect 434 237 435 238
rect 433 237 434 238
rect 432 237 433 238
rect 422 237 423 238
rect 421 237 422 238
rect 420 237 421 238
rect 419 237 420 238
rect 418 237 419 238
rect 417 237 418 238
rect 416 237 417 238
rect 395 237 396 238
rect 394 237 395 238
rect 393 237 394 238
rect 392 237 393 238
rect 306 237 307 238
rect 305 237 306 238
rect 304 237 305 238
rect 303 237 304 238
rect 302 237 303 238
rect 301 237 302 238
rect 300 237 301 238
rect 299 237 300 238
rect 298 237 299 238
rect 297 237 298 238
rect 296 237 297 238
rect 295 237 296 238
rect 294 237 295 238
rect 293 237 294 238
rect 292 237 293 238
rect 291 237 292 238
rect 290 237 291 238
rect 267 237 268 238
rect 266 237 267 238
rect 265 237 266 238
rect 264 237 265 238
rect 263 237 264 238
rect 262 237 263 238
rect 261 237 262 238
rect 260 237 261 238
rect 259 237 260 238
rect 258 237 259 238
rect 257 237 258 238
rect 256 237 257 238
rect 255 237 256 238
rect 254 237 255 238
rect 253 237 254 238
rect 252 237 253 238
rect 251 237 252 238
rect 250 237 251 238
rect 249 237 250 238
rect 248 237 249 238
rect 247 237 248 238
rect 246 237 247 238
rect 245 237 246 238
rect 244 237 245 238
rect 243 237 244 238
rect 242 237 243 238
rect 241 237 242 238
rect 240 237 241 238
rect 239 237 240 238
rect 238 237 239 238
rect 237 237 238 238
rect 236 237 237 238
rect 235 237 236 238
rect 234 237 235 238
rect 233 237 234 238
rect 232 237 233 238
rect 231 237 232 238
rect 230 237 231 238
rect 229 237 230 238
rect 228 237 229 238
rect 227 237 228 238
rect 226 237 227 238
rect 225 237 226 238
rect 224 237 225 238
rect 223 237 224 238
rect 222 237 223 238
rect 221 237 222 238
rect 220 237 221 238
rect 219 237 220 238
rect 218 237 219 238
rect 217 237 218 238
rect 216 237 217 238
rect 215 237 216 238
rect 214 237 215 238
rect 213 237 214 238
rect 212 237 213 238
rect 211 237 212 238
rect 210 237 211 238
rect 209 237 210 238
rect 208 237 209 238
rect 207 237 208 238
rect 206 237 207 238
rect 205 237 206 238
rect 204 237 205 238
rect 203 237 204 238
rect 202 237 203 238
rect 201 237 202 238
rect 200 237 201 238
rect 199 237 200 238
rect 198 237 199 238
rect 197 237 198 238
rect 196 237 197 238
rect 195 237 196 238
rect 194 237 195 238
rect 193 237 194 238
rect 192 237 193 238
rect 191 237 192 238
rect 190 237 191 238
rect 189 237 190 238
rect 188 237 189 238
rect 187 237 188 238
rect 186 237 187 238
rect 185 237 186 238
rect 184 237 185 238
rect 183 237 184 238
rect 182 237 183 238
rect 181 237 182 238
rect 180 237 181 238
rect 179 237 180 238
rect 178 237 179 238
rect 177 237 178 238
rect 176 237 177 238
rect 175 237 176 238
rect 174 237 175 238
rect 146 237 147 238
rect 145 237 146 238
rect 144 237 145 238
rect 143 237 144 238
rect 142 237 143 238
rect 141 237 142 238
rect 140 237 141 238
rect 139 237 140 238
rect 138 237 139 238
rect 137 237 138 238
rect 136 237 137 238
rect 135 237 136 238
rect 134 237 135 238
rect 133 237 134 238
rect 132 237 133 238
rect 131 237 132 238
rect 130 237 131 238
rect 129 237 130 238
rect 128 237 129 238
rect 127 237 128 238
rect 126 237 127 238
rect 125 237 126 238
rect 124 237 125 238
rect 123 237 124 238
rect 122 237 123 238
rect 121 237 122 238
rect 120 237 121 238
rect 119 237 120 238
rect 118 237 119 238
rect 117 237 118 238
rect 116 237 117 238
rect 99 237 100 238
rect 98 237 99 238
rect 97 237 98 238
rect 96 237 97 238
rect 95 237 96 238
rect 94 237 95 238
rect 93 237 94 238
rect 92 237 93 238
rect 91 237 92 238
rect 90 237 91 238
rect 89 237 90 238
rect 88 237 89 238
rect 87 237 88 238
rect 86 237 87 238
rect 85 237 86 238
rect 84 237 85 238
rect 83 237 84 238
rect 82 237 83 238
rect 81 237 82 238
rect 80 237 81 238
rect 79 237 80 238
rect 78 237 79 238
rect 77 237 78 238
rect 76 237 77 238
rect 75 237 76 238
rect 74 237 75 238
rect 73 237 74 238
rect 72 237 73 238
rect 71 237 72 238
rect 70 237 71 238
rect 69 237 70 238
rect 68 237 69 238
rect 67 237 68 238
rect 66 237 67 238
rect 65 237 66 238
rect 64 237 65 238
rect 63 237 64 238
rect 62 237 63 238
rect 61 237 62 238
rect 60 237 61 238
rect 59 237 60 238
rect 58 237 59 238
rect 57 237 58 238
rect 56 237 57 238
rect 55 237 56 238
rect 54 237 55 238
rect 53 237 54 238
rect 52 237 53 238
rect 51 237 52 238
rect 50 237 51 238
rect 49 237 50 238
rect 48 237 49 238
rect 47 237 48 238
rect 46 237 47 238
rect 45 237 46 238
rect 44 237 45 238
rect 43 237 44 238
rect 42 237 43 238
rect 41 237 42 238
rect 40 237 41 238
rect 39 237 40 238
rect 38 237 39 238
rect 37 237 38 238
rect 36 237 37 238
rect 35 237 36 238
rect 34 237 35 238
rect 33 237 34 238
rect 32 237 33 238
rect 31 237 32 238
rect 30 237 31 238
rect 29 237 30 238
rect 28 237 29 238
rect 27 237 28 238
rect 26 237 27 238
rect 19 237 20 238
rect 18 237 19 238
rect 17 237 18 238
rect 16 237 17 238
rect 15 237 16 238
rect 14 237 15 238
rect 13 237 14 238
rect 12 237 13 238
rect 11 237 12 238
rect 10 237 11 238
rect 9 237 10 238
rect 8 237 9 238
rect 7 237 8 238
rect 6 237 7 238
rect 5 237 6 238
rect 4 237 5 238
rect 3 237 4 238
rect 2 237 3 238
rect 438 238 439 239
rect 437 238 438 239
rect 436 238 437 239
rect 435 238 436 239
rect 434 238 435 239
rect 433 238 434 239
rect 432 238 433 239
rect 431 238 432 239
rect 430 238 431 239
rect 429 238 430 239
rect 428 238 429 239
rect 427 238 428 239
rect 426 238 427 239
rect 425 238 426 239
rect 424 238 425 239
rect 423 238 424 239
rect 422 238 423 239
rect 421 238 422 239
rect 420 238 421 239
rect 419 238 420 239
rect 418 238 419 239
rect 417 238 418 239
rect 416 238 417 239
rect 396 238 397 239
rect 395 238 396 239
rect 394 238 395 239
rect 393 238 394 239
rect 392 238 393 239
rect 314 238 315 239
rect 313 238 314 239
rect 312 238 313 239
rect 311 238 312 239
rect 310 238 311 239
rect 309 238 310 239
rect 308 238 309 239
rect 307 238 308 239
rect 306 238 307 239
rect 305 238 306 239
rect 304 238 305 239
rect 303 238 304 239
rect 302 238 303 239
rect 301 238 302 239
rect 300 238 301 239
rect 299 238 300 239
rect 298 238 299 239
rect 297 238 298 239
rect 296 238 297 239
rect 295 238 296 239
rect 294 238 295 239
rect 293 238 294 239
rect 292 238 293 239
rect 291 238 292 239
rect 290 238 291 239
rect 289 238 290 239
rect 288 238 289 239
rect 287 238 288 239
rect 286 238 287 239
rect 285 238 286 239
rect 284 238 285 239
rect 283 238 284 239
rect 266 238 267 239
rect 265 238 266 239
rect 264 238 265 239
rect 263 238 264 239
rect 262 238 263 239
rect 261 238 262 239
rect 260 238 261 239
rect 259 238 260 239
rect 258 238 259 239
rect 257 238 258 239
rect 256 238 257 239
rect 255 238 256 239
rect 254 238 255 239
rect 253 238 254 239
rect 252 238 253 239
rect 251 238 252 239
rect 250 238 251 239
rect 249 238 250 239
rect 248 238 249 239
rect 247 238 248 239
rect 246 238 247 239
rect 245 238 246 239
rect 244 238 245 239
rect 243 238 244 239
rect 242 238 243 239
rect 241 238 242 239
rect 240 238 241 239
rect 239 238 240 239
rect 238 238 239 239
rect 237 238 238 239
rect 236 238 237 239
rect 235 238 236 239
rect 234 238 235 239
rect 233 238 234 239
rect 232 238 233 239
rect 231 238 232 239
rect 230 238 231 239
rect 229 238 230 239
rect 228 238 229 239
rect 227 238 228 239
rect 226 238 227 239
rect 225 238 226 239
rect 224 238 225 239
rect 223 238 224 239
rect 222 238 223 239
rect 221 238 222 239
rect 220 238 221 239
rect 219 238 220 239
rect 218 238 219 239
rect 217 238 218 239
rect 216 238 217 239
rect 215 238 216 239
rect 214 238 215 239
rect 213 238 214 239
rect 212 238 213 239
rect 211 238 212 239
rect 210 238 211 239
rect 209 238 210 239
rect 208 238 209 239
rect 207 238 208 239
rect 206 238 207 239
rect 205 238 206 239
rect 204 238 205 239
rect 203 238 204 239
rect 202 238 203 239
rect 201 238 202 239
rect 200 238 201 239
rect 199 238 200 239
rect 198 238 199 239
rect 197 238 198 239
rect 196 238 197 239
rect 195 238 196 239
rect 194 238 195 239
rect 193 238 194 239
rect 192 238 193 239
rect 191 238 192 239
rect 190 238 191 239
rect 189 238 190 239
rect 188 238 189 239
rect 187 238 188 239
rect 186 238 187 239
rect 185 238 186 239
rect 184 238 185 239
rect 183 238 184 239
rect 182 238 183 239
rect 181 238 182 239
rect 180 238 181 239
rect 179 238 180 239
rect 178 238 179 239
rect 177 238 178 239
rect 147 238 148 239
rect 146 238 147 239
rect 145 238 146 239
rect 144 238 145 239
rect 143 238 144 239
rect 142 238 143 239
rect 141 238 142 239
rect 140 238 141 239
rect 139 238 140 239
rect 138 238 139 239
rect 137 238 138 239
rect 136 238 137 239
rect 135 238 136 239
rect 134 238 135 239
rect 133 238 134 239
rect 132 238 133 239
rect 131 238 132 239
rect 130 238 131 239
rect 129 238 130 239
rect 128 238 129 239
rect 127 238 128 239
rect 126 238 127 239
rect 125 238 126 239
rect 124 238 125 239
rect 123 238 124 239
rect 122 238 123 239
rect 121 238 122 239
rect 120 238 121 239
rect 119 238 120 239
rect 118 238 119 239
rect 117 238 118 239
rect 116 238 117 239
rect 100 238 101 239
rect 99 238 100 239
rect 98 238 99 239
rect 97 238 98 239
rect 96 238 97 239
rect 95 238 96 239
rect 94 238 95 239
rect 93 238 94 239
rect 92 238 93 239
rect 91 238 92 239
rect 90 238 91 239
rect 89 238 90 239
rect 88 238 89 239
rect 87 238 88 239
rect 86 238 87 239
rect 85 238 86 239
rect 84 238 85 239
rect 83 238 84 239
rect 82 238 83 239
rect 81 238 82 239
rect 80 238 81 239
rect 79 238 80 239
rect 78 238 79 239
rect 77 238 78 239
rect 76 238 77 239
rect 75 238 76 239
rect 74 238 75 239
rect 73 238 74 239
rect 72 238 73 239
rect 71 238 72 239
rect 70 238 71 239
rect 69 238 70 239
rect 68 238 69 239
rect 67 238 68 239
rect 66 238 67 239
rect 65 238 66 239
rect 64 238 65 239
rect 63 238 64 239
rect 62 238 63 239
rect 61 238 62 239
rect 60 238 61 239
rect 59 238 60 239
rect 58 238 59 239
rect 57 238 58 239
rect 56 238 57 239
rect 55 238 56 239
rect 54 238 55 239
rect 53 238 54 239
rect 52 238 53 239
rect 51 238 52 239
rect 50 238 51 239
rect 49 238 50 239
rect 48 238 49 239
rect 47 238 48 239
rect 46 238 47 239
rect 45 238 46 239
rect 44 238 45 239
rect 43 238 44 239
rect 42 238 43 239
rect 41 238 42 239
rect 40 238 41 239
rect 39 238 40 239
rect 38 238 39 239
rect 37 238 38 239
rect 36 238 37 239
rect 35 238 36 239
rect 34 238 35 239
rect 33 238 34 239
rect 32 238 33 239
rect 31 238 32 239
rect 30 238 31 239
rect 29 238 30 239
rect 28 238 29 239
rect 27 238 28 239
rect 26 238 27 239
rect 19 238 20 239
rect 18 238 19 239
rect 17 238 18 239
rect 16 238 17 239
rect 15 238 16 239
rect 14 238 15 239
rect 13 238 14 239
rect 12 238 13 239
rect 11 238 12 239
rect 10 238 11 239
rect 9 238 10 239
rect 8 238 9 239
rect 7 238 8 239
rect 6 238 7 239
rect 5 238 6 239
rect 4 238 5 239
rect 3 238 4 239
rect 2 238 3 239
rect 1 238 2 239
rect 437 239 438 240
rect 436 239 437 240
rect 435 239 436 240
rect 434 239 435 240
rect 433 239 434 240
rect 432 239 433 240
rect 431 239 432 240
rect 430 239 431 240
rect 429 239 430 240
rect 428 239 429 240
rect 427 239 428 240
rect 426 239 427 240
rect 425 239 426 240
rect 424 239 425 240
rect 423 239 424 240
rect 422 239 423 240
rect 421 239 422 240
rect 420 239 421 240
rect 419 239 420 240
rect 418 239 419 240
rect 417 239 418 240
rect 416 239 417 240
rect 397 239 398 240
rect 396 239 397 240
rect 395 239 396 240
rect 394 239 395 240
rect 393 239 394 240
rect 318 239 319 240
rect 317 239 318 240
rect 316 239 317 240
rect 315 239 316 240
rect 314 239 315 240
rect 313 239 314 240
rect 312 239 313 240
rect 311 239 312 240
rect 310 239 311 240
rect 309 239 310 240
rect 308 239 309 240
rect 307 239 308 240
rect 306 239 307 240
rect 305 239 306 240
rect 304 239 305 240
rect 303 239 304 240
rect 302 239 303 240
rect 301 239 302 240
rect 300 239 301 240
rect 299 239 300 240
rect 298 239 299 240
rect 297 239 298 240
rect 296 239 297 240
rect 295 239 296 240
rect 294 239 295 240
rect 293 239 294 240
rect 292 239 293 240
rect 291 239 292 240
rect 290 239 291 240
rect 289 239 290 240
rect 288 239 289 240
rect 287 239 288 240
rect 286 239 287 240
rect 285 239 286 240
rect 284 239 285 240
rect 283 239 284 240
rect 282 239 283 240
rect 281 239 282 240
rect 280 239 281 240
rect 279 239 280 240
rect 278 239 279 240
rect 265 239 266 240
rect 264 239 265 240
rect 263 239 264 240
rect 262 239 263 240
rect 261 239 262 240
rect 260 239 261 240
rect 259 239 260 240
rect 258 239 259 240
rect 257 239 258 240
rect 256 239 257 240
rect 255 239 256 240
rect 254 239 255 240
rect 253 239 254 240
rect 252 239 253 240
rect 251 239 252 240
rect 250 239 251 240
rect 249 239 250 240
rect 248 239 249 240
rect 247 239 248 240
rect 246 239 247 240
rect 245 239 246 240
rect 244 239 245 240
rect 243 239 244 240
rect 242 239 243 240
rect 241 239 242 240
rect 240 239 241 240
rect 239 239 240 240
rect 238 239 239 240
rect 237 239 238 240
rect 236 239 237 240
rect 235 239 236 240
rect 234 239 235 240
rect 233 239 234 240
rect 232 239 233 240
rect 231 239 232 240
rect 230 239 231 240
rect 229 239 230 240
rect 228 239 229 240
rect 227 239 228 240
rect 226 239 227 240
rect 225 239 226 240
rect 224 239 225 240
rect 223 239 224 240
rect 222 239 223 240
rect 221 239 222 240
rect 220 239 221 240
rect 219 239 220 240
rect 218 239 219 240
rect 217 239 218 240
rect 216 239 217 240
rect 215 239 216 240
rect 214 239 215 240
rect 213 239 214 240
rect 212 239 213 240
rect 211 239 212 240
rect 210 239 211 240
rect 209 239 210 240
rect 208 239 209 240
rect 207 239 208 240
rect 206 239 207 240
rect 205 239 206 240
rect 204 239 205 240
rect 203 239 204 240
rect 202 239 203 240
rect 201 239 202 240
rect 200 239 201 240
rect 199 239 200 240
rect 198 239 199 240
rect 197 239 198 240
rect 196 239 197 240
rect 195 239 196 240
rect 194 239 195 240
rect 193 239 194 240
rect 192 239 193 240
rect 191 239 192 240
rect 190 239 191 240
rect 189 239 190 240
rect 188 239 189 240
rect 187 239 188 240
rect 186 239 187 240
rect 185 239 186 240
rect 184 239 185 240
rect 183 239 184 240
rect 182 239 183 240
rect 181 239 182 240
rect 180 239 181 240
rect 179 239 180 240
rect 148 239 149 240
rect 147 239 148 240
rect 146 239 147 240
rect 145 239 146 240
rect 144 239 145 240
rect 143 239 144 240
rect 142 239 143 240
rect 141 239 142 240
rect 140 239 141 240
rect 139 239 140 240
rect 138 239 139 240
rect 137 239 138 240
rect 136 239 137 240
rect 135 239 136 240
rect 134 239 135 240
rect 133 239 134 240
rect 132 239 133 240
rect 131 239 132 240
rect 130 239 131 240
rect 129 239 130 240
rect 128 239 129 240
rect 127 239 128 240
rect 126 239 127 240
rect 125 239 126 240
rect 124 239 125 240
rect 123 239 124 240
rect 122 239 123 240
rect 121 239 122 240
rect 120 239 121 240
rect 119 239 120 240
rect 118 239 119 240
rect 117 239 118 240
rect 101 239 102 240
rect 100 239 101 240
rect 99 239 100 240
rect 98 239 99 240
rect 97 239 98 240
rect 96 239 97 240
rect 95 239 96 240
rect 94 239 95 240
rect 93 239 94 240
rect 92 239 93 240
rect 91 239 92 240
rect 90 239 91 240
rect 89 239 90 240
rect 88 239 89 240
rect 87 239 88 240
rect 86 239 87 240
rect 85 239 86 240
rect 84 239 85 240
rect 83 239 84 240
rect 82 239 83 240
rect 81 239 82 240
rect 80 239 81 240
rect 79 239 80 240
rect 78 239 79 240
rect 77 239 78 240
rect 76 239 77 240
rect 75 239 76 240
rect 74 239 75 240
rect 73 239 74 240
rect 72 239 73 240
rect 71 239 72 240
rect 70 239 71 240
rect 69 239 70 240
rect 68 239 69 240
rect 67 239 68 240
rect 66 239 67 240
rect 65 239 66 240
rect 64 239 65 240
rect 63 239 64 240
rect 62 239 63 240
rect 61 239 62 240
rect 60 239 61 240
rect 59 239 60 240
rect 58 239 59 240
rect 57 239 58 240
rect 56 239 57 240
rect 55 239 56 240
rect 54 239 55 240
rect 53 239 54 240
rect 52 239 53 240
rect 51 239 52 240
rect 50 239 51 240
rect 49 239 50 240
rect 48 239 49 240
rect 47 239 48 240
rect 46 239 47 240
rect 45 239 46 240
rect 44 239 45 240
rect 43 239 44 240
rect 42 239 43 240
rect 41 239 42 240
rect 40 239 41 240
rect 39 239 40 240
rect 38 239 39 240
rect 37 239 38 240
rect 36 239 37 240
rect 35 239 36 240
rect 34 239 35 240
rect 33 239 34 240
rect 32 239 33 240
rect 31 239 32 240
rect 30 239 31 240
rect 29 239 30 240
rect 28 239 29 240
rect 27 239 28 240
rect 26 239 27 240
rect 19 239 20 240
rect 18 239 19 240
rect 17 239 18 240
rect 16 239 17 240
rect 15 239 16 240
rect 14 239 15 240
rect 13 239 14 240
rect 12 239 13 240
rect 11 239 12 240
rect 10 239 11 240
rect 9 239 10 240
rect 8 239 9 240
rect 7 239 8 240
rect 6 239 7 240
rect 5 239 6 240
rect 4 239 5 240
rect 3 239 4 240
rect 2 239 3 240
rect 1 239 2 240
rect 437 240 438 241
rect 436 240 437 241
rect 435 240 436 241
rect 434 240 435 241
rect 433 240 434 241
rect 432 240 433 241
rect 431 240 432 241
rect 430 240 431 241
rect 429 240 430 241
rect 428 240 429 241
rect 427 240 428 241
rect 426 240 427 241
rect 425 240 426 241
rect 424 240 425 241
rect 423 240 424 241
rect 422 240 423 241
rect 421 240 422 241
rect 420 240 421 241
rect 419 240 420 241
rect 418 240 419 241
rect 417 240 418 241
rect 416 240 417 241
rect 398 240 399 241
rect 397 240 398 241
rect 396 240 397 241
rect 395 240 396 241
rect 394 240 395 241
rect 393 240 394 241
rect 322 240 323 241
rect 321 240 322 241
rect 320 240 321 241
rect 319 240 320 241
rect 318 240 319 241
rect 317 240 318 241
rect 316 240 317 241
rect 315 240 316 241
rect 314 240 315 241
rect 313 240 314 241
rect 312 240 313 241
rect 311 240 312 241
rect 310 240 311 241
rect 309 240 310 241
rect 308 240 309 241
rect 307 240 308 241
rect 306 240 307 241
rect 305 240 306 241
rect 304 240 305 241
rect 303 240 304 241
rect 302 240 303 241
rect 301 240 302 241
rect 300 240 301 241
rect 299 240 300 241
rect 298 240 299 241
rect 297 240 298 241
rect 296 240 297 241
rect 295 240 296 241
rect 294 240 295 241
rect 293 240 294 241
rect 292 240 293 241
rect 291 240 292 241
rect 290 240 291 241
rect 289 240 290 241
rect 288 240 289 241
rect 287 240 288 241
rect 286 240 287 241
rect 285 240 286 241
rect 284 240 285 241
rect 283 240 284 241
rect 282 240 283 241
rect 281 240 282 241
rect 280 240 281 241
rect 279 240 280 241
rect 278 240 279 241
rect 277 240 278 241
rect 276 240 277 241
rect 275 240 276 241
rect 274 240 275 241
rect 265 240 266 241
rect 264 240 265 241
rect 263 240 264 241
rect 262 240 263 241
rect 261 240 262 241
rect 260 240 261 241
rect 259 240 260 241
rect 258 240 259 241
rect 257 240 258 241
rect 256 240 257 241
rect 255 240 256 241
rect 254 240 255 241
rect 253 240 254 241
rect 252 240 253 241
rect 251 240 252 241
rect 250 240 251 241
rect 249 240 250 241
rect 248 240 249 241
rect 247 240 248 241
rect 246 240 247 241
rect 245 240 246 241
rect 244 240 245 241
rect 243 240 244 241
rect 242 240 243 241
rect 241 240 242 241
rect 240 240 241 241
rect 239 240 240 241
rect 238 240 239 241
rect 237 240 238 241
rect 236 240 237 241
rect 235 240 236 241
rect 234 240 235 241
rect 233 240 234 241
rect 232 240 233 241
rect 231 240 232 241
rect 230 240 231 241
rect 226 240 227 241
rect 225 240 226 241
rect 224 240 225 241
rect 223 240 224 241
rect 222 240 223 241
rect 221 240 222 241
rect 220 240 221 241
rect 219 240 220 241
rect 218 240 219 241
rect 217 240 218 241
rect 216 240 217 241
rect 215 240 216 241
rect 214 240 215 241
rect 213 240 214 241
rect 212 240 213 241
rect 211 240 212 241
rect 210 240 211 241
rect 209 240 210 241
rect 208 240 209 241
rect 207 240 208 241
rect 206 240 207 241
rect 205 240 206 241
rect 204 240 205 241
rect 203 240 204 241
rect 202 240 203 241
rect 201 240 202 241
rect 200 240 201 241
rect 199 240 200 241
rect 198 240 199 241
rect 197 240 198 241
rect 196 240 197 241
rect 195 240 196 241
rect 194 240 195 241
rect 193 240 194 241
rect 192 240 193 241
rect 191 240 192 241
rect 190 240 191 241
rect 189 240 190 241
rect 188 240 189 241
rect 187 240 188 241
rect 186 240 187 241
rect 185 240 186 241
rect 184 240 185 241
rect 183 240 184 241
rect 182 240 183 241
rect 148 240 149 241
rect 147 240 148 241
rect 146 240 147 241
rect 145 240 146 241
rect 144 240 145 241
rect 143 240 144 241
rect 142 240 143 241
rect 141 240 142 241
rect 140 240 141 241
rect 139 240 140 241
rect 138 240 139 241
rect 137 240 138 241
rect 136 240 137 241
rect 135 240 136 241
rect 134 240 135 241
rect 133 240 134 241
rect 132 240 133 241
rect 131 240 132 241
rect 130 240 131 241
rect 129 240 130 241
rect 128 240 129 241
rect 127 240 128 241
rect 126 240 127 241
rect 125 240 126 241
rect 124 240 125 241
rect 123 240 124 241
rect 122 240 123 241
rect 121 240 122 241
rect 120 240 121 241
rect 119 240 120 241
rect 118 240 119 241
rect 117 240 118 241
rect 102 240 103 241
rect 101 240 102 241
rect 100 240 101 241
rect 99 240 100 241
rect 98 240 99 241
rect 97 240 98 241
rect 96 240 97 241
rect 95 240 96 241
rect 94 240 95 241
rect 93 240 94 241
rect 92 240 93 241
rect 91 240 92 241
rect 90 240 91 241
rect 89 240 90 241
rect 88 240 89 241
rect 87 240 88 241
rect 86 240 87 241
rect 85 240 86 241
rect 84 240 85 241
rect 83 240 84 241
rect 82 240 83 241
rect 81 240 82 241
rect 80 240 81 241
rect 79 240 80 241
rect 78 240 79 241
rect 77 240 78 241
rect 76 240 77 241
rect 75 240 76 241
rect 74 240 75 241
rect 73 240 74 241
rect 72 240 73 241
rect 71 240 72 241
rect 70 240 71 241
rect 69 240 70 241
rect 68 240 69 241
rect 67 240 68 241
rect 66 240 67 241
rect 65 240 66 241
rect 64 240 65 241
rect 63 240 64 241
rect 62 240 63 241
rect 61 240 62 241
rect 60 240 61 241
rect 59 240 60 241
rect 58 240 59 241
rect 57 240 58 241
rect 56 240 57 241
rect 55 240 56 241
rect 54 240 55 241
rect 53 240 54 241
rect 52 240 53 241
rect 51 240 52 241
rect 50 240 51 241
rect 49 240 50 241
rect 48 240 49 241
rect 47 240 48 241
rect 46 240 47 241
rect 45 240 46 241
rect 44 240 45 241
rect 43 240 44 241
rect 42 240 43 241
rect 41 240 42 241
rect 40 240 41 241
rect 39 240 40 241
rect 38 240 39 241
rect 37 240 38 241
rect 36 240 37 241
rect 35 240 36 241
rect 34 240 35 241
rect 33 240 34 241
rect 32 240 33 241
rect 31 240 32 241
rect 30 240 31 241
rect 29 240 30 241
rect 28 240 29 241
rect 27 240 28 241
rect 19 240 20 241
rect 18 240 19 241
rect 17 240 18 241
rect 16 240 17 241
rect 15 240 16 241
rect 14 240 15 241
rect 13 240 14 241
rect 12 240 13 241
rect 11 240 12 241
rect 10 240 11 241
rect 9 240 10 241
rect 8 240 9 241
rect 7 240 8 241
rect 6 240 7 241
rect 5 240 6 241
rect 4 240 5 241
rect 3 240 4 241
rect 2 240 3 241
rect 1 240 2 241
rect 437 241 438 242
rect 436 241 437 242
rect 435 241 436 242
rect 434 241 435 242
rect 433 241 434 242
rect 432 241 433 242
rect 431 241 432 242
rect 430 241 431 242
rect 429 241 430 242
rect 428 241 429 242
rect 427 241 428 242
rect 426 241 427 242
rect 425 241 426 242
rect 424 241 425 242
rect 423 241 424 242
rect 422 241 423 242
rect 421 241 422 242
rect 420 241 421 242
rect 419 241 420 242
rect 418 241 419 242
rect 417 241 418 242
rect 416 241 417 242
rect 399 241 400 242
rect 398 241 399 242
rect 397 241 398 242
rect 396 241 397 242
rect 395 241 396 242
rect 394 241 395 242
rect 393 241 394 242
rect 325 241 326 242
rect 324 241 325 242
rect 323 241 324 242
rect 322 241 323 242
rect 321 241 322 242
rect 320 241 321 242
rect 319 241 320 242
rect 318 241 319 242
rect 317 241 318 242
rect 316 241 317 242
rect 315 241 316 242
rect 314 241 315 242
rect 313 241 314 242
rect 312 241 313 242
rect 311 241 312 242
rect 310 241 311 242
rect 309 241 310 242
rect 308 241 309 242
rect 307 241 308 242
rect 306 241 307 242
rect 305 241 306 242
rect 304 241 305 242
rect 303 241 304 242
rect 302 241 303 242
rect 301 241 302 242
rect 300 241 301 242
rect 299 241 300 242
rect 298 241 299 242
rect 297 241 298 242
rect 296 241 297 242
rect 295 241 296 242
rect 294 241 295 242
rect 293 241 294 242
rect 292 241 293 242
rect 291 241 292 242
rect 290 241 291 242
rect 289 241 290 242
rect 288 241 289 242
rect 287 241 288 242
rect 286 241 287 242
rect 285 241 286 242
rect 284 241 285 242
rect 283 241 284 242
rect 282 241 283 242
rect 281 241 282 242
rect 280 241 281 242
rect 279 241 280 242
rect 278 241 279 242
rect 277 241 278 242
rect 276 241 277 242
rect 275 241 276 242
rect 274 241 275 242
rect 273 241 274 242
rect 272 241 273 242
rect 271 241 272 242
rect 264 241 265 242
rect 263 241 264 242
rect 262 241 263 242
rect 261 241 262 242
rect 260 241 261 242
rect 259 241 260 242
rect 258 241 259 242
rect 257 241 258 242
rect 256 241 257 242
rect 255 241 256 242
rect 254 241 255 242
rect 253 241 254 242
rect 252 241 253 242
rect 251 241 252 242
rect 250 241 251 242
rect 249 241 250 242
rect 248 241 249 242
rect 247 241 248 242
rect 246 241 247 242
rect 245 241 246 242
rect 244 241 245 242
rect 243 241 244 242
rect 242 241 243 242
rect 241 241 242 242
rect 240 241 241 242
rect 239 241 240 242
rect 238 241 239 242
rect 237 241 238 242
rect 236 241 237 242
rect 235 241 236 242
rect 234 241 235 242
rect 233 241 234 242
rect 232 241 233 242
rect 231 241 232 242
rect 230 241 231 242
rect 222 241 223 242
rect 221 241 222 242
rect 220 241 221 242
rect 219 241 220 242
rect 218 241 219 242
rect 217 241 218 242
rect 216 241 217 242
rect 215 241 216 242
rect 214 241 215 242
rect 213 241 214 242
rect 212 241 213 242
rect 211 241 212 242
rect 210 241 211 242
rect 209 241 210 242
rect 208 241 209 242
rect 207 241 208 242
rect 206 241 207 242
rect 205 241 206 242
rect 204 241 205 242
rect 203 241 204 242
rect 202 241 203 242
rect 201 241 202 242
rect 200 241 201 242
rect 199 241 200 242
rect 198 241 199 242
rect 197 241 198 242
rect 196 241 197 242
rect 195 241 196 242
rect 194 241 195 242
rect 193 241 194 242
rect 192 241 193 242
rect 191 241 192 242
rect 190 241 191 242
rect 189 241 190 242
rect 188 241 189 242
rect 187 241 188 242
rect 186 241 187 242
rect 185 241 186 242
rect 149 241 150 242
rect 148 241 149 242
rect 147 241 148 242
rect 146 241 147 242
rect 145 241 146 242
rect 144 241 145 242
rect 143 241 144 242
rect 142 241 143 242
rect 141 241 142 242
rect 140 241 141 242
rect 139 241 140 242
rect 138 241 139 242
rect 137 241 138 242
rect 136 241 137 242
rect 135 241 136 242
rect 134 241 135 242
rect 133 241 134 242
rect 132 241 133 242
rect 131 241 132 242
rect 130 241 131 242
rect 129 241 130 242
rect 128 241 129 242
rect 127 241 128 242
rect 126 241 127 242
rect 125 241 126 242
rect 124 241 125 242
rect 123 241 124 242
rect 122 241 123 242
rect 121 241 122 242
rect 120 241 121 242
rect 119 241 120 242
rect 118 241 119 242
rect 117 241 118 242
rect 102 241 103 242
rect 101 241 102 242
rect 100 241 101 242
rect 99 241 100 242
rect 98 241 99 242
rect 97 241 98 242
rect 96 241 97 242
rect 95 241 96 242
rect 94 241 95 242
rect 93 241 94 242
rect 92 241 93 242
rect 91 241 92 242
rect 90 241 91 242
rect 89 241 90 242
rect 88 241 89 242
rect 87 241 88 242
rect 86 241 87 242
rect 85 241 86 242
rect 84 241 85 242
rect 83 241 84 242
rect 82 241 83 242
rect 81 241 82 242
rect 80 241 81 242
rect 79 241 80 242
rect 78 241 79 242
rect 77 241 78 242
rect 76 241 77 242
rect 75 241 76 242
rect 74 241 75 242
rect 73 241 74 242
rect 72 241 73 242
rect 71 241 72 242
rect 70 241 71 242
rect 69 241 70 242
rect 68 241 69 242
rect 67 241 68 242
rect 66 241 67 242
rect 65 241 66 242
rect 64 241 65 242
rect 63 241 64 242
rect 62 241 63 242
rect 61 241 62 242
rect 60 241 61 242
rect 59 241 60 242
rect 58 241 59 242
rect 57 241 58 242
rect 56 241 57 242
rect 55 241 56 242
rect 54 241 55 242
rect 53 241 54 242
rect 52 241 53 242
rect 51 241 52 242
rect 50 241 51 242
rect 49 241 50 242
rect 48 241 49 242
rect 47 241 48 242
rect 46 241 47 242
rect 45 241 46 242
rect 44 241 45 242
rect 43 241 44 242
rect 42 241 43 242
rect 41 241 42 242
rect 40 241 41 242
rect 39 241 40 242
rect 38 241 39 242
rect 37 241 38 242
rect 36 241 37 242
rect 35 241 36 242
rect 34 241 35 242
rect 33 241 34 242
rect 32 241 33 242
rect 31 241 32 242
rect 30 241 31 242
rect 29 241 30 242
rect 28 241 29 242
rect 27 241 28 242
rect 19 241 20 242
rect 18 241 19 242
rect 17 241 18 242
rect 16 241 17 242
rect 15 241 16 242
rect 14 241 15 242
rect 13 241 14 242
rect 12 241 13 242
rect 11 241 12 242
rect 10 241 11 242
rect 9 241 10 242
rect 8 241 9 242
rect 7 241 8 242
rect 6 241 7 242
rect 5 241 6 242
rect 4 241 5 242
rect 3 241 4 242
rect 2 241 3 242
rect 1 241 2 242
rect 477 242 478 243
rect 476 242 477 243
rect 475 242 476 243
rect 474 242 475 243
rect 473 242 474 243
rect 464 242 465 243
rect 463 242 464 243
rect 462 242 463 243
rect 437 242 438 243
rect 436 242 437 243
rect 435 242 436 243
rect 434 242 435 243
rect 433 242 434 243
rect 432 242 433 243
rect 431 242 432 243
rect 430 242 431 243
rect 429 242 430 243
rect 428 242 429 243
rect 427 242 428 243
rect 426 242 427 243
rect 425 242 426 243
rect 424 242 425 243
rect 423 242 424 243
rect 422 242 423 243
rect 421 242 422 243
rect 420 242 421 243
rect 419 242 420 243
rect 418 242 419 243
rect 417 242 418 243
rect 416 242 417 243
rect 400 242 401 243
rect 399 242 400 243
rect 398 242 399 243
rect 397 242 398 243
rect 396 242 397 243
rect 395 242 396 243
rect 394 242 395 243
rect 393 242 394 243
rect 325 242 326 243
rect 324 242 325 243
rect 323 242 324 243
rect 322 242 323 243
rect 321 242 322 243
rect 320 242 321 243
rect 319 242 320 243
rect 318 242 319 243
rect 317 242 318 243
rect 316 242 317 243
rect 315 242 316 243
rect 314 242 315 243
rect 313 242 314 243
rect 312 242 313 243
rect 311 242 312 243
rect 310 242 311 243
rect 309 242 310 243
rect 308 242 309 243
rect 307 242 308 243
rect 306 242 307 243
rect 305 242 306 243
rect 304 242 305 243
rect 303 242 304 243
rect 302 242 303 243
rect 301 242 302 243
rect 300 242 301 243
rect 299 242 300 243
rect 298 242 299 243
rect 297 242 298 243
rect 296 242 297 243
rect 295 242 296 243
rect 294 242 295 243
rect 293 242 294 243
rect 292 242 293 243
rect 291 242 292 243
rect 290 242 291 243
rect 289 242 290 243
rect 288 242 289 243
rect 287 242 288 243
rect 286 242 287 243
rect 285 242 286 243
rect 284 242 285 243
rect 283 242 284 243
rect 282 242 283 243
rect 281 242 282 243
rect 280 242 281 243
rect 279 242 280 243
rect 278 242 279 243
rect 277 242 278 243
rect 276 242 277 243
rect 275 242 276 243
rect 274 242 275 243
rect 273 242 274 243
rect 272 242 273 243
rect 271 242 272 243
rect 270 242 271 243
rect 269 242 270 243
rect 263 242 264 243
rect 262 242 263 243
rect 261 242 262 243
rect 260 242 261 243
rect 259 242 260 243
rect 258 242 259 243
rect 257 242 258 243
rect 256 242 257 243
rect 255 242 256 243
rect 254 242 255 243
rect 253 242 254 243
rect 252 242 253 243
rect 251 242 252 243
rect 250 242 251 243
rect 249 242 250 243
rect 248 242 249 243
rect 247 242 248 243
rect 246 242 247 243
rect 245 242 246 243
rect 244 242 245 243
rect 243 242 244 243
rect 242 242 243 243
rect 241 242 242 243
rect 240 242 241 243
rect 239 242 240 243
rect 238 242 239 243
rect 237 242 238 243
rect 236 242 237 243
rect 235 242 236 243
rect 234 242 235 243
rect 233 242 234 243
rect 232 242 233 243
rect 231 242 232 243
rect 230 242 231 243
rect 218 242 219 243
rect 217 242 218 243
rect 216 242 217 243
rect 215 242 216 243
rect 214 242 215 243
rect 213 242 214 243
rect 212 242 213 243
rect 211 242 212 243
rect 210 242 211 243
rect 209 242 210 243
rect 208 242 209 243
rect 207 242 208 243
rect 206 242 207 243
rect 205 242 206 243
rect 204 242 205 243
rect 203 242 204 243
rect 202 242 203 243
rect 201 242 202 243
rect 200 242 201 243
rect 199 242 200 243
rect 198 242 199 243
rect 197 242 198 243
rect 196 242 197 243
rect 195 242 196 243
rect 194 242 195 243
rect 193 242 194 243
rect 192 242 193 243
rect 191 242 192 243
rect 190 242 191 243
rect 189 242 190 243
rect 150 242 151 243
rect 149 242 150 243
rect 148 242 149 243
rect 147 242 148 243
rect 146 242 147 243
rect 145 242 146 243
rect 144 242 145 243
rect 143 242 144 243
rect 142 242 143 243
rect 141 242 142 243
rect 140 242 141 243
rect 139 242 140 243
rect 138 242 139 243
rect 137 242 138 243
rect 136 242 137 243
rect 135 242 136 243
rect 134 242 135 243
rect 133 242 134 243
rect 132 242 133 243
rect 131 242 132 243
rect 130 242 131 243
rect 129 242 130 243
rect 128 242 129 243
rect 127 242 128 243
rect 126 242 127 243
rect 125 242 126 243
rect 124 242 125 243
rect 123 242 124 243
rect 122 242 123 243
rect 121 242 122 243
rect 120 242 121 243
rect 119 242 120 243
rect 118 242 119 243
rect 117 242 118 243
rect 103 242 104 243
rect 102 242 103 243
rect 101 242 102 243
rect 100 242 101 243
rect 99 242 100 243
rect 98 242 99 243
rect 97 242 98 243
rect 96 242 97 243
rect 95 242 96 243
rect 94 242 95 243
rect 93 242 94 243
rect 92 242 93 243
rect 91 242 92 243
rect 90 242 91 243
rect 89 242 90 243
rect 88 242 89 243
rect 87 242 88 243
rect 86 242 87 243
rect 85 242 86 243
rect 84 242 85 243
rect 83 242 84 243
rect 82 242 83 243
rect 81 242 82 243
rect 80 242 81 243
rect 79 242 80 243
rect 78 242 79 243
rect 77 242 78 243
rect 76 242 77 243
rect 75 242 76 243
rect 74 242 75 243
rect 73 242 74 243
rect 72 242 73 243
rect 71 242 72 243
rect 70 242 71 243
rect 69 242 70 243
rect 68 242 69 243
rect 67 242 68 243
rect 66 242 67 243
rect 65 242 66 243
rect 64 242 65 243
rect 63 242 64 243
rect 62 242 63 243
rect 61 242 62 243
rect 60 242 61 243
rect 59 242 60 243
rect 58 242 59 243
rect 57 242 58 243
rect 56 242 57 243
rect 55 242 56 243
rect 54 242 55 243
rect 53 242 54 243
rect 52 242 53 243
rect 51 242 52 243
rect 50 242 51 243
rect 49 242 50 243
rect 48 242 49 243
rect 47 242 48 243
rect 46 242 47 243
rect 45 242 46 243
rect 44 242 45 243
rect 43 242 44 243
rect 42 242 43 243
rect 41 242 42 243
rect 40 242 41 243
rect 39 242 40 243
rect 38 242 39 243
rect 37 242 38 243
rect 36 242 37 243
rect 35 242 36 243
rect 34 242 35 243
rect 33 242 34 243
rect 32 242 33 243
rect 31 242 32 243
rect 30 242 31 243
rect 29 242 30 243
rect 28 242 29 243
rect 27 242 28 243
rect 19 242 20 243
rect 18 242 19 243
rect 17 242 18 243
rect 16 242 17 243
rect 15 242 16 243
rect 14 242 15 243
rect 13 242 14 243
rect 12 242 13 243
rect 11 242 12 243
rect 10 242 11 243
rect 9 242 10 243
rect 8 242 9 243
rect 7 242 8 243
rect 6 242 7 243
rect 5 242 6 243
rect 4 242 5 243
rect 3 242 4 243
rect 2 242 3 243
rect 1 242 2 243
rect 478 243 479 244
rect 477 243 478 244
rect 476 243 477 244
rect 475 243 476 244
rect 474 243 475 244
rect 466 243 467 244
rect 465 243 466 244
rect 464 243 465 244
rect 463 243 464 244
rect 462 243 463 244
rect 461 243 462 244
rect 460 243 461 244
rect 437 243 438 244
rect 436 243 437 244
rect 435 243 436 244
rect 434 243 435 244
rect 433 243 434 244
rect 432 243 433 244
rect 431 243 432 244
rect 430 243 431 244
rect 429 243 430 244
rect 428 243 429 244
rect 427 243 428 244
rect 426 243 427 244
rect 425 243 426 244
rect 424 243 425 244
rect 423 243 424 244
rect 422 243 423 244
rect 421 243 422 244
rect 420 243 421 244
rect 419 243 420 244
rect 418 243 419 244
rect 417 243 418 244
rect 416 243 417 244
rect 402 243 403 244
rect 401 243 402 244
rect 400 243 401 244
rect 399 243 400 244
rect 398 243 399 244
rect 397 243 398 244
rect 396 243 397 244
rect 395 243 396 244
rect 394 243 395 244
rect 393 243 394 244
rect 323 243 324 244
rect 322 243 323 244
rect 321 243 322 244
rect 320 243 321 244
rect 319 243 320 244
rect 318 243 319 244
rect 317 243 318 244
rect 316 243 317 244
rect 315 243 316 244
rect 314 243 315 244
rect 313 243 314 244
rect 312 243 313 244
rect 311 243 312 244
rect 310 243 311 244
rect 309 243 310 244
rect 308 243 309 244
rect 307 243 308 244
rect 306 243 307 244
rect 305 243 306 244
rect 304 243 305 244
rect 303 243 304 244
rect 302 243 303 244
rect 301 243 302 244
rect 300 243 301 244
rect 299 243 300 244
rect 298 243 299 244
rect 297 243 298 244
rect 296 243 297 244
rect 295 243 296 244
rect 294 243 295 244
rect 293 243 294 244
rect 292 243 293 244
rect 291 243 292 244
rect 290 243 291 244
rect 289 243 290 244
rect 288 243 289 244
rect 287 243 288 244
rect 286 243 287 244
rect 285 243 286 244
rect 284 243 285 244
rect 283 243 284 244
rect 282 243 283 244
rect 281 243 282 244
rect 280 243 281 244
rect 279 243 280 244
rect 278 243 279 244
rect 277 243 278 244
rect 276 243 277 244
rect 275 243 276 244
rect 274 243 275 244
rect 273 243 274 244
rect 272 243 273 244
rect 271 243 272 244
rect 270 243 271 244
rect 269 243 270 244
rect 268 243 269 244
rect 267 243 268 244
rect 263 243 264 244
rect 262 243 263 244
rect 261 243 262 244
rect 260 243 261 244
rect 259 243 260 244
rect 258 243 259 244
rect 257 243 258 244
rect 256 243 257 244
rect 255 243 256 244
rect 254 243 255 244
rect 253 243 254 244
rect 252 243 253 244
rect 251 243 252 244
rect 250 243 251 244
rect 249 243 250 244
rect 248 243 249 244
rect 247 243 248 244
rect 246 243 247 244
rect 245 243 246 244
rect 244 243 245 244
rect 243 243 244 244
rect 242 243 243 244
rect 241 243 242 244
rect 240 243 241 244
rect 239 243 240 244
rect 238 243 239 244
rect 237 243 238 244
rect 236 243 237 244
rect 235 243 236 244
rect 234 243 235 244
rect 233 243 234 244
rect 232 243 233 244
rect 231 243 232 244
rect 230 243 231 244
rect 212 243 213 244
rect 211 243 212 244
rect 210 243 211 244
rect 209 243 210 244
rect 208 243 209 244
rect 207 243 208 244
rect 206 243 207 244
rect 205 243 206 244
rect 204 243 205 244
rect 203 243 204 244
rect 202 243 203 244
rect 201 243 202 244
rect 200 243 201 244
rect 199 243 200 244
rect 198 243 199 244
rect 197 243 198 244
rect 196 243 197 244
rect 195 243 196 244
rect 194 243 195 244
rect 151 243 152 244
rect 150 243 151 244
rect 149 243 150 244
rect 148 243 149 244
rect 147 243 148 244
rect 146 243 147 244
rect 145 243 146 244
rect 144 243 145 244
rect 143 243 144 244
rect 142 243 143 244
rect 141 243 142 244
rect 140 243 141 244
rect 139 243 140 244
rect 138 243 139 244
rect 137 243 138 244
rect 136 243 137 244
rect 135 243 136 244
rect 134 243 135 244
rect 133 243 134 244
rect 132 243 133 244
rect 131 243 132 244
rect 130 243 131 244
rect 129 243 130 244
rect 128 243 129 244
rect 127 243 128 244
rect 126 243 127 244
rect 125 243 126 244
rect 124 243 125 244
rect 123 243 124 244
rect 122 243 123 244
rect 121 243 122 244
rect 120 243 121 244
rect 119 243 120 244
rect 118 243 119 244
rect 103 243 104 244
rect 102 243 103 244
rect 101 243 102 244
rect 100 243 101 244
rect 99 243 100 244
rect 98 243 99 244
rect 97 243 98 244
rect 96 243 97 244
rect 95 243 96 244
rect 94 243 95 244
rect 93 243 94 244
rect 92 243 93 244
rect 91 243 92 244
rect 90 243 91 244
rect 89 243 90 244
rect 88 243 89 244
rect 87 243 88 244
rect 86 243 87 244
rect 85 243 86 244
rect 84 243 85 244
rect 83 243 84 244
rect 82 243 83 244
rect 81 243 82 244
rect 80 243 81 244
rect 79 243 80 244
rect 78 243 79 244
rect 77 243 78 244
rect 76 243 77 244
rect 75 243 76 244
rect 74 243 75 244
rect 73 243 74 244
rect 72 243 73 244
rect 71 243 72 244
rect 70 243 71 244
rect 69 243 70 244
rect 68 243 69 244
rect 67 243 68 244
rect 66 243 67 244
rect 65 243 66 244
rect 64 243 65 244
rect 63 243 64 244
rect 62 243 63 244
rect 61 243 62 244
rect 60 243 61 244
rect 59 243 60 244
rect 58 243 59 244
rect 57 243 58 244
rect 56 243 57 244
rect 55 243 56 244
rect 54 243 55 244
rect 53 243 54 244
rect 52 243 53 244
rect 51 243 52 244
rect 50 243 51 244
rect 49 243 50 244
rect 48 243 49 244
rect 47 243 48 244
rect 46 243 47 244
rect 45 243 46 244
rect 44 243 45 244
rect 43 243 44 244
rect 42 243 43 244
rect 41 243 42 244
rect 40 243 41 244
rect 39 243 40 244
rect 38 243 39 244
rect 37 243 38 244
rect 36 243 37 244
rect 35 243 36 244
rect 34 243 35 244
rect 33 243 34 244
rect 32 243 33 244
rect 31 243 32 244
rect 30 243 31 244
rect 29 243 30 244
rect 28 243 29 244
rect 27 243 28 244
rect 19 243 20 244
rect 18 243 19 244
rect 17 243 18 244
rect 16 243 17 244
rect 15 243 16 244
rect 14 243 15 244
rect 13 243 14 244
rect 12 243 13 244
rect 11 243 12 244
rect 10 243 11 244
rect 9 243 10 244
rect 8 243 9 244
rect 7 243 8 244
rect 6 243 7 244
rect 5 243 6 244
rect 4 243 5 244
rect 3 243 4 244
rect 2 243 3 244
rect 1 243 2 244
rect 478 244 479 245
rect 477 244 478 245
rect 476 244 477 245
rect 475 244 476 245
rect 467 244 468 245
rect 466 244 467 245
rect 465 244 466 245
rect 464 244 465 245
rect 463 244 464 245
rect 462 244 463 245
rect 461 244 462 245
rect 460 244 461 245
rect 459 244 460 245
rect 436 244 437 245
rect 435 244 436 245
rect 434 244 435 245
rect 433 244 434 245
rect 432 244 433 245
rect 431 244 432 245
rect 430 244 431 245
rect 429 244 430 245
rect 428 244 429 245
rect 427 244 428 245
rect 426 244 427 245
rect 425 244 426 245
rect 424 244 425 245
rect 423 244 424 245
rect 422 244 423 245
rect 421 244 422 245
rect 420 244 421 245
rect 419 244 420 245
rect 418 244 419 245
rect 417 244 418 245
rect 416 244 417 245
rect 405 244 406 245
rect 404 244 405 245
rect 403 244 404 245
rect 402 244 403 245
rect 401 244 402 245
rect 400 244 401 245
rect 399 244 400 245
rect 398 244 399 245
rect 397 244 398 245
rect 396 244 397 245
rect 395 244 396 245
rect 394 244 395 245
rect 321 244 322 245
rect 320 244 321 245
rect 319 244 320 245
rect 318 244 319 245
rect 317 244 318 245
rect 316 244 317 245
rect 315 244 316 245
rect 314 244 315 245
rect 313 244 314 245
rect 312 244 313 245
rect 311 244 312 245
rect 310 244 311 245
rect 309 244 310 245
rect 308 244 309 245
rect 307 244 308 245
rect 306 244 307 245
rect 305 244 306 245
rect 304 244 305 245
rect 303 244 304 245
rect 302 244 303 245
rect 301 244 302 245
rect 300 244 301 245
rect 299 244 300 245
rect 298 244 299 245
rect 297 244 298 245
rect 296 244 297 245
rect 295 244 296 245
rect 294 244 295 245
rect 293 244 294 245
rect 292 244 293 245
rect 291 244 292 245
rect 290 244 291 245
rect 289 244 290 245
rect 288 244 289 245
rect 287 244 288 245
rect 286 244 287 245
rect 285 244 286 245
rect 284 244 285 245
rect 283 244 284 245
rect 282 244 283 245
rect 281 244 282 245
rect 280 244 281 245
rect 279 244 280 245
rect 278 244 279 245
rect 277 244 278 245
rect 276 244 277 245
rect 275 244 276 245
rect 274 244 275 245
rect 273 244 274 245
rect 272 244 273 245
rect 271 244 272 245
rect 270 244 271 245
rect 269 244 270 245
rect 268 244 269 245
rect 267 244 268 245
rect 266 244 267 245
rect 265 244 266 245
rect 262 244 263 245
rect 261 244 262 245
rect 260 244 261 245
rect 259 244 260 245
rect 258 244 259 245
rect 257 244 258 245
rect 256 244 257 245
rect 255 244 256 245
rect 254 244 255 245
rect 253 244 254 245
rect 252 244 253 245
rect 251 244 252 245
rect 250 244 251 245
rect 249 244 250 245
rect 248 244 249 245
rect 247 244 248 245
rect 246 244 247 245
rect 245 244 246 245
rect 244 244 245 245
rect 243 244 244 245
rect 242 244 243 245
rect 241 244 242 245
rect 240 244 241 245
rect 239 244 240 245
rect 238 244 239 245
rect 237 244 238 245
rect 236 244 237 245
rect 235 244 236 245
rect 234 244 235 245
rect 233 244 234 245
rect 232 244 233 245
rect 231 244 232 245
rect 230 244 231 245
rect 152 244 153 245
rect 151 244 152 245
rect 150 244 151 245
rect 149 244 150 245
rect 148 244 149 245
rect 147 244 148 245
rect 146 244 147 245
rect 145 244 146 245
rect 144 244 145 245
rect 143 244 144 245
rect 142 244 143 245
rect 141 244 142 245
rect 140 244 141 245
rect 139 244 140 245
rect 138 244 139 245
rect 137 244 138 245
rect 136 244 137 245
rect 135 244 136 245
rect 134 244 135 245
rect 133 244 134 245
rect 132 244 133 245
rect 131 244 132 245
rect 130 244 131 245
rect 129 244 130 245
rect 128 244 129 245
rect 127 244 128 245
rect 126 244 127 245
rect 125 244 126 245
rect 124 244 125 245
rect 123 244 124 245
rect 122 244 123 245
rect 121 244 122 245
rect 120 244 121 245
rect 119 244 120 245
rect 118 244 119 245
rect 104 244 105 245
rect 103 244 104 245
rect 102 244 103 245
rect 101 244 102 245
rect 100 244 101 245
rect 99 244 100 245
rect 98 244 99 245
rect 97 244 98 245
rect 96 244 97 245
rect 95 244 96 245
rect 94 244 95 245
rect 93 244 94 245
rect 92 244 93 245
rect 91 244 92 245
rect 90 244 91 245
rect 89 244 90 245
rect 88 244 89 245
rect 87 244 88 245
rect 86 244 87 245
rect 85 244 86 245
rect 84 244 85 245
rect 83 244 84 245
rect 82 244 83 245
rect 81 244 82 245
rect 80 244 81 245
rect 79 244 80 245
rect 78 244 79 245
rect 77 244 78 245
rect 76 244 77 245
rect 75 244 76 245
rect 74 244 75 245
rect 73 244 74 245
rect 72 244 73 245
rect 71 244 72 245
rect 70 244 71 245
rect 69 244 70 245
rect 68 244 69 245
rect 67 244 68 245
rect 66 244 67 245
rect 65 244 66 245
rect 64 244 65 245
rect 63 244 64 245
rect 62 244 63 245
rect 61 244 62 245
rect 60 244 61 245
rect 59 244 60 245
rect 58 244 59 245
rect 57 244 58 245
rect 56 244 57 245
rect 55 244 56 245
rect 54 244 55 245
rect 53 244 54 245
rect 52 244 53 245
rect 51 244 52 245
rect 50 244 51 245
rect 49 244 50 245
rect 48 244 49 245
rect 47 244 48 245
rect 46 244 47 245
rect 45 244 46 245
rect 44 244 45 245
rect 43 244 44 245
rect 42 244 43 245
rect 41 244 42 245
rect 40 244 41 245
rect 39 244 40 245
rect 38 244 39 245
rect 37 244 38 245
rect 36 244 37 245
rect 35 244 36 245
rect 34 244 35 245
rect 33 244 34 245
rect 32 244 33 245
rect 31 244 32 245
rect 30 244 31 245
rect 29 244 30 245
rect 28 244 29 245
rect 19 244 20 245
rect 18 244 19 245
rect 17 244 18 245
rect 16 244 17 245
rect 15 244 16 245
rect 14 244 15 245
rect 13 244 14 245
rect 12 244 13 245
rect 11 244 12 245
rect 10 244 11 245
rect 9 244 10 245
rect 8 244 9 245
rect 7 244 8 245
rect 6 244 7 245
rect 5 244 6 245
rect 4 244 5 245
rect 3 244 4 245
rect 2 244 3 245
rect 1 244 2 245
rect 479 245 480 246
rect 478 245 479 246
rect 477 245 478 246
rect 468 245 469 246
rect 467 245 468 246
rect 466 245 467 246
rect 465 245 466 246
rect 464 245 465 246
rect 463 245 464 246
rect 462 245 463 246
rect 461 245 462 246
rect 460 245 461 246
rect 459 245 460 246
rect 458 245 459 246
rect 436 245 437 246
rect 435 245 436 246
rect 434 245 435 246
rect 433 245 434 246
rect 432 245 433 246
rect 431 245 432 246
rect 430 245 431 246
rect 429 245 430 246
rect 428 245 429 246
rect 427 245 428 246
rect 426 245 427 246
rect 425 245 426 246
rect 424 245 425 246
rect 423 245 424 246
rect 422 245 423 246
rect 421 245 422 246
rect 420 245 421 246
rect 419 245 420 246
rect 418 245 419 246
rect 417 245 418 246
rect 416 245 417 246
rect 405 245 406 246
rect 404 245 405 246
rect 403 245 404 246
rect 402 245 403 246
rect 401 245 402 246
rect 400 245 401 246
rect 399 245 400 246
rect 398 245 399 246
rect 397 245 398 246
rect 396 245 397 246
rect 395 245 396 246
rect 394 245 395 246
rect 319 245 320 246
rect 318 245 319 246
rect 317 245 318 246
rect 316 245 317 246
rect 315 245 316 246
rect 314 245 315 246
rect 313 245 314 246
rect 312 245 313 246
rect 311 245 312 246
rect 310 245 311 246
rect 309 245 310 246
rect 308 245 309 246
rect 307 245 308 246
rect 306 245 307 246
rect 305 245 306 246
rect 304 245 305 246
rect 303 245 304 246
rect 302 245 303 246
rect 301 245 302 246
rect 300 245 301 246
rect 299 245 300 246
rect 298 245 299 246
rect 297 245 298 246
rect 296 245 297 246
rect 295 245 296 246
rect 294 245 295 246
rect 293 245 294 246
rect 292 245 293 246
rect 291 245 292 246
rect 290 245 291 246
rect 289 245 290 246
rect 288 245 289 246
rect 287 245 288 246
rect 286 245 287 246
rect 285 245 286 246
rect 284 245 285 246
rect 283 245 284 246
rect 282 245 283 246
rect 281 245 282 246
rect 280 245 281 246
rect 279 245 280 246
rect 278 245 279 246
rect 277 245 278 246
rect 276 245 277 246
rect 275 245 276 246
rect 274 245 275 246
rect 273 245 274 246
rect 272 245 273 246
rect 271 245 272 246
rect 270 245 271 246
rect 269 245 270 246
rect 268 245 269 246
rect 267 245 268 246
rect 266 245 267 246
rect 265 245 266 246
rect 264 245 265 246
rect 263 245 264 246
rect 261 245 262 246
rect 260 245 261 246
rect 259 245 260 246
rect 258 245 259 246
rect 257 245 258 246
rect 256 245 257 246
rect 255 245 256 246
rect 254 245 255 246
rect 253 245 254 246
rect 252 245 253 246
rect 251 245 252 246
rect 250 245 251 246
rect 249 245 250 246
rect 248 245 249 246
rect 247 245 248 246
rect 246 245 247 246
rect 245 245 246 246
rect 244 245 245 246
rect 243 245 244 246
rect 242 245 243 246
rect 241 245 242 246
rect 240 245 241 246
rect 239 245 240 246
rect 238 245 239 246
rect 237 245 238 246
rect 236 245 237 246
rect 235 245 236 246
rect 234 245 235 246
rect 233 245 234 246
rect 232 245 233 246
rect 231 245 232 246
rect 230 245 231 246
rect 153 245 154 246
rect 152 245 153 246
rect 151 245 152 246
rect 150 245 151 246
rect 149 245 150 246
rect 148 245 149 246
rect 147 245 148 246
rect 146 245 147 246
rect 145 245 146 246
rect 144 245 145 246
rect 143 245 144 246
rect 142 245 143 246
rect 141 245 142 246
rect 140 245 141 246
rect 139 245 140 246
rect 138 245 139 246
rect 137 245 138 246
rect 136 245 137 246
rect 135 245 136 246
rect 134 245 135 246
rect 133 245 134 246
rect 132 245 133 246
rect 131 245 132 246
rect 130 245 131 246
rect 129 245 130 246
rect 128 245 129 246
rect 127 245 128 246
rect 126 245 127 246
rect 125 245 126 246
rect 124 245 125 246
rect 123 245 124 246
rect 122 245 123 246
rect 121 245 122 246
rect 120 245 121 246
rect 119 245 120 246
rect 118 245 119 246
rect 104 245 105 246
rect 103 245 104 246
rect 102 245 103 246
rect 101 245 102 246
rect 100 245 101 246
rect 99 245 100 246
rect 98 245 99 246
rect 97 245 98 246
rect 96 245 97 246
rect 95 245 96 246
rect 94 245 95 246
rect 93 245 94 246
rect 92 245 93 246
rect 91 245 92 246
rect 90 245 91 246
rect 89 245 90 246
rect 88 245 89 246
rect 87 245 88 246
rect 86 245 87 246
rect 85 245 86 246
rect 84 245 85 246
rect 83 245 84 246
rect 82 245 83 246
rect 81 245 82 246
rect 80 245 81 246
rect 79 245 80 246
rect 78 245 79 246
rect 77 245 78 246
rect 76 245 77 246
rect 75 245 76 246
rect 74 245 75 246
rect 73 245 74 246
rect 72 245 73 246
rect 71 245 72 246
rect 70 245 71 246
rect 69 245 70 246
rect 68 245 69 246
rect 67 245 68 246
rect 66 245 67 246
rect 65 245 66 246
rect 64 245 65 246
rect 63 245 64 246
rect 62 245 63 246
rect 61 245 62 246
rect 60 245 61 246
rect 59 245 60 246
rect 58 245 59 246
rect 57 245 58 246
rect 56 245 57 246
rect 55 245 56 246
rect 54 245 55 246
rect 53 245 54 246
rect 52 245 53 246
rect 51 245 52 246
rect 50 245 51 246
rect 49 245 50 246
rect 48 245 49 246
rect 47 245 48 246
rect 46 245 47 246
rect 45 245 46 246
rect 44 245 45 246
rect 43 245 44 246
rect 42 245 43 246
rect 41 245 42 246
rect 40 245 41 246
rect 39 245 40 246
rect 38 245 39 246
rect 37 245 38 246
rect 36 245 37 246
rect 35 245 36 246
rect 34 245 35 246
rect 33 245 34 246
rect 32 245 33 246
rect 31 245 32 246
rect 30 245 31 246
rect 29 245 30 246
rect 28 245 29 246
rect 19 245 20 246
rect 18 245 19 246
rect 17 245 18 246
rect 16 245 17 246
rect 15 245 16 246
rect 14 245 15 246
rect 13 245 14 246
rect 12 245 13 246
rect 11 245 12 246
rect 10 245 11 246
rect 9 245 10 246
rect 8 245 9 246
rect 7 245 8 246
rect 6 245 7 246
rect 5 245 6 246
rect 4 245 5 246
rect 3 245 4 246
rect 2 245 3 246
rect 1 245 2 246
rect 479 246 480 247
rect 478 246 479 247
rect 469 246 470 247
rect 468 246 469 247
rect 467 246 468 247
rect 466 246 467 247
rect 465 246 466 247
rect 464 246 465 247
rect 463 246 464 247
rect 460 246 461 247
rect 459 246 460 247
rect 458 246 459 247
rect 436 246 437 247
rect 435 246 436 247
rect 434 246 435 247
rect 433 246 434 247
rect 432 246 433 247
rect 431 246 432 247
rect 430 246 431 247
rect 429 246 430 247
rect 428 246 429 247
rect 427 246 428 247
rect 426 246 427 247
rect 425 246 426 247
rect 424 246 425 247
rect 423 246 424 247
rect 422 246 423 247
rect 421 246 422 247
rect 420 246 421 247
rect 419 246 420 247
rect 418 246 419 247
rect 417 246 418 247
rect 416 246 417 247
rect 405 246 406 247
rect 404 246 405 247
rect 403 246 404 247
rect 402 246 403 247
rect 401 246 402 247
rect 400 246 401 247
rect 399 246 400 247
rect 398 246 399 247
rect 397 246 398 247
rect 317 246 318 247
rect 316 246 317 247
rect 315 246 316 247
rect 314 246 315 247
rect 313 246 314 247
rect 312 246 313 247
rect 311 246 312 247
rect 310 246 311 247
rect 309 246 310 247
rect 308 246 309 247
rect 307 246 308 247
rect 306 246 307 247
rect 305 246 306 247
rect 304 246 305 247
rect 303 246 304 247
rect 302 246 303 247
rect 301 246 302 247
rect 300 246 301 247
rect 299 246 300 247
rect 298 246 299 247
rect 297 246 298 247
rect 296 246 297 247
rect 295 246 296 247
rect 294 246 295 247
rect 293 246 294 247
rect 292 246 293 247
rect 291 246 292 247
rect 290 246 291 247
rect 289 246 290 247
rect 288 246 289 247
rect 287 246 288 247
rect 286 246 287 247
rect 285 246 286 247
rect 284 246 285 247
rect 283 246 284 247
rect 282 246 283 247
rect 281 246 282 247
rect 280 246 281 247
rect 279 246 280 247
rect 278 246 279 247
rect 277 246 278 247
rect 276 246 277 247
rect 275 246 276 247
rect 274 246 275 247
rect 273 246 274 247
rect 272 246 273 247
rect 271 246 272 247
rect 270 246 271 247
rect 269 246 270 247
rect 268 246 269 247
rect 267 246 268 247
rect 266 246 267 247
rect 265 246 266 247
rect 264 246 265 247
rect 263 246 264 247
rect 262 246 263 247
rect 261 246 262 247
rect 260 246 261 247
rect 259 246 260 247
rect 258 246 259 247
rect 257 246 258 247
rect 256 246 257 247
rect 255 246 256 247
rect 254 246 255 247
rect 253 246 254 247
rect 252 246 253 247
rect 251 246 252 247
rect 250 246 251 247
rect 249 246 250 247
rect 248 246 249 247
rect 247 246 248 247
rect 246 246 247 247
rect 245 246 246 247
rect 244 246 245 247
rect 243 246 244 247
rect 242 246 243 247
rect 241 246 242 247
rect 240 246 241 247
rect 239 246 240 247
rect 238 246 239 247
rect 237 246 238 247
rect 236 246 237 247
rect 235 246 236 247
rect 234 246 235 247
rect 233 246 234 247
rect 232 246 233 247
rect 231 246 232 247
rect 230 246 231 247
rect 154 246 155 247
rect 153 246 154 247
rect 152 246 153 247
rect 151 246 152 247
rect 150 246 151 247
rect 149 246 150 247
rect 148 246 149 247
rect 147 246 148 247
rect 146 246 147 247
rect 145 246 146 247
rect 144 246 145 247
rect 143 246 144 247
rect 142 246 143 247
rect 141 246 142 247
rect 140 246 141 247
rect 139 246 140 247
rect 138 246 139 247
rect 137 246 138 247
rect 136 246 137 247
rect 135 246 136 247
rect 134 246 135 247
rect 133 246 134 247
rect 132 246 133 247
rect 131 246 132 247
rect 130 246 131 247
rect 129 246 130 247
rect 128 246 129 247
rect 127 246 128 247
rect 126 246 127 247
rect 125 246 126 247
rect 124 246 125 247
rect 123 246 124 247
rect 122 246 123 247
rect 121 246 122 247
rect 120 246 121 247
rect 119 246 120 247
rect 118 246 119 247
rect 105 246 106 247
rect 104 246 105 247
rect 103 246 104 247
rect 102 246 103 247
rect 101 246 102 247
rect 100 246 101 247
rect 99 246 100 247
rect 98 246 99 247
rect 97 246 98 247
rect 96 246 97 247
rect 95 246 96 247
rect 94 246 95 247
rect 93 246 94 247
rect 92 246 93 247
rect 91 246 92 247
rect 90 246 91 247
rect 89 246 90 247
rect 88 246 89 247
rect 87 246 88 247
rect 86 246 87 247
rect 85 246 86 247
rect 84 246 85 247
rect 83 246 84 247
rect 82 246 83 247
rect 81 246 82 247
rect 80 246 81 247
rect 79 246 80 247
rect 78 246 79 247
rect 77 246 78 247
rect 76 246 77 247
rect 75 246 76 247
rect 74 246 75 247
rect 73 246 74 247
rect 72 246 73 247
rect 71 246 72 247
rect 70 246 71 247
rect 69 246 70 247
rect 68 246 69 247
rect 67 246 68 247
rect 66 246 67 247
rect 65 246 66 247
rect 64 246 65 247
rect 63 246 64 247
rect 62 246 63 247
rect 61 246 62 247
rect 60 246 61 247
rect 59 246 60 247
rect 58 246 59 247
rect 57 246 58 247
rect 56 246 57 247
rect 55 246 56 247
rect 54 246 55 247
rect 53 246 54 247
rect 52 246 53 247
rect 51 246 52 247
rect 50 246 51 247
rect 49 246 50 247
rect 48 246 49 247
rect 47 246 48 247
rect 46 246 47 247
rect 45 246 46 247
rect 44 246 45 247
rect 43 246 44 247
rect 42 246 43 247
rect 41 246 42 247
rect 40 246 41 247
rect 39 246 40 247
rect 38 246 39 247
rect 37 246 38 247
rect 36 246 37 247
rect 35 246 36 247
rect 34 246 35 247
rect 33 246 34 247
rect 32 246 33 247
rect 31 246 32 247
rect 30 246 31 247
rect 29 246 30 247
rect 28 246 29 247
rect 19 246 20 247
rect 18 246 19 247
rect 17 246 18 247
rect 16 246 17 247
rect 15 246 16 247
rect 14 246 15 247
rect 13 246 14 247
rect 12 246 13 247
rect 11 246 12 247
rect 10 246 11 247
rect 9 246 10 247
rect 8 246 9 247
rect 7 246 8 247
rect 6 246 7 247
rect 5 246 6 247
rect 4 246 5 247
rect 3 246 4 247
rect 2 246 3 247
rect 1 246 2 247
rect 479 247 480 248
rect 478 247 479 248
rect 469 247 470 248
rect 468 247 469 248
rect 467 247 468 248
rect 466 247 467 248
rect 465 247 466 248
rect 464 247 465 248
rect 458 247 459 248
rect 457 247 458 248
rect 420 247 421 248
rect 419 247 420 248
rect 418 247 419 248
rect 417 247 418 248
rect 416 247 417 248
rect 316 247 317 248
rect 315 247 316 248
rect 314 247 315 248
rect 313 247 314 248
rect 312 247 313 248
rect 311 247 312 248
rect 310 247 311 248
rect 309 247 310 248
rect 308 247 309 248
rect 307 247 308 248
rect 306 247 307 248
rect 305 247 306 248
rect 304 247 305 248
rect 303 247 304 248
rect 302 247 303 248
rect 301 247 302 248
rect 300 247 301 248
rect 299 247 300 248
rect 298 247 299 248
rect 297 247 298 248
rect 296 247 297 248
rect 295 247 296 248
rect 294 247 295 248
rect 293 247 294 248
rect 292 247 293 248
rect 291 247 292 248
rect 290 247 291 248
rect 289 247 290 248
rect 288 247 289 248
rect 287 247 288 248
rect 286 247 287 248
rect 285 247 286 248
rect 284 247 285 248
rect 283 247 284 248
rect 282 247 283 248
rect 281 247 282 248
rect 280 247 281 248
rect 279 247 280 248
rect 278 247 279 248
rect 277 247 278 248
rect 276 247 277 248
rect 275 247 276 248
rect 274 247 275 248
rect 273 247 274 248
rect 272 247 273 248
rect 271 247 272 248
rect 270 247 271 248
rect 269 247 270 248
rect 268 247 269 248
rect 267 247 268 248
rect 266 247 267 248
rect 265 247 266 248
rect 264 247 265 248
rect 263 247 264 248
rect 262 247 263 248
rect 261 247 262 248
rect 260 247 261 248
rect 259 247 260 248
rect 258 247 259 248
rect 257 247 258 248
rect 256 247 257 248
rect 255 247 256 248
rect 254 247 255 248
rect 253 247 254 248
rect 252 247 253 248
rect 251 247 252 248
rect 250 247 251 248
rect 249 247 250 248
rect 248 247 249 248
rect 247 247 248 248
rect 246 247 247 248
rect 245 247 246 248
rect 244 247 245 248
rect 243 247 244 248
rect 242 247 243 248
rect 241 247 242 248
rect 240 247 241 248
rect 239 247 240 248
rect 238 247 239 248
rect 237 247 238 248
rect 236 247 237 248
rect 235 247 236 248
rect 234 247 235 248
rect 233 247 234 248
rect 232 247 233 248
rect 231 247 232 248
rect 230 247 231 248
rect 229 247 230 248
rect 155 247 156 248
rect 154 247 155 248
rect 153 247 154 248
rect 152 247 153 248
rect 151 247 152 248
rect 150 247 151 248
rect 149 247 150 248
rect 148 247 149 248
rect 147 247 148 248
rect 146 247 147 248
rect 145 247 146 248
rect 144 247 145 248
rect 143 247 144 248
rect 142 247 143 248
rect 141 247 142 248
rect 140 247 141 248
rect 139 247 140 248
rect 138 247 139 248
rect 137 247 138 248
rect 136 247 137 248
rect 135 247 136 248
rect 134 247 135 248
rect 133 247 134 248
rect 132 247 133 248
rect 131 247 132 248
rect 130 247 131 248
rect 129 247 130 248
rect 128 247 129 248
rect 127 247 128 248
rect 126 247 127 248
rect 125 247 126 248
rect 124 247 125 248
rect 123 247 124 248
rect 122 247 123 248
rect 121 247 122 248
rect 120 247 121 248
rect 119 247 120 248
rect 118 247 119 248
rect 105 247 106 248
rect 104 247 105 248
rect 103 247 104 248
rect 102 247 103 248
rect 101 247 102 248
rect 100 247 101 248
rect 99 247 100 248
rect 98 247 99 248
rect 97 247 98 248
rect 96 247 97 248
rect 95 247 96 248
rect 94 247 95 248
rect 93 247 94 248
rect 92 247 93 248
rect 91 247 92 248
rect 90 247 91 248
rect 89 247 90 248
rect 88 247 89 248
rect 87 247 88 248
rect 86 247 87 248
rect 85 247 86 248
rect 84 247 85 248
rect 83 247 84 248
rect 82 247 83 248
rect 81 247 82 248
rect 80 247 81 248
rect 79 247 80 248
rect 78 247 79 248
rect 77 247 78 248
rect 76 247 77 248
rect 75 247 76 248
rect 74 247 75 248
rect 73 247 74 248
rect 72 247 73 248
rect 71 247 72 248
rect 70 247 71 248
rect 69 247 70 248
rect 68 247 69 248
rect 67 247 68 248
rect 66 247 67 248
rect 65 247 66 248
rect 64 247 65 248
rect 63 247 64 248
rect 62 247 63 248
rect 61 247 62 248
rect 60 247 61 248
rect 59 247 60 248
rect 58 247 59 248
rect 57 247 58 248
rect 56 247 57 248
rect 55 247 56 248
rect 54 247 55 248
rect 53 247 54 248
rect 52 247 53 248
rect 51 247 52 248
rect 50 247 51 248
rect 49 247 50 248
rect 48 247 49 248
rect 47 247 48 248
rect 46 247 47 248
rect 45 247 46 248
rect 44 247 45 248
rect 43 247 44 248
rect 42 247 43 248
rect 41 247 42 248
rect 40 247 41 248
rect 39 247 40 248
rect 38 247 39 248
rect 37 247 38 248
rect 36 247 37 248
rect 35 247 36 248
rect 34 247 35 248
rect 33 247 34 248
rect 32 247 33 248
rect 31 247 32 248
rect 30 247 31 248
rect 29 247 30 248
rect 19 247 20 248
rect 18 247 19 248
rect 17 247 18 248
rect 16 247 17 248
rect 15 247 16 248
rect 14 247 15 248
rect 13 247 14 248
rect 12 247 13 248
rect 11 247 12 248
rect 10 247 11 248
rect 9 247 10 248
rect 8 247 9 248
rect 7 247 8 248
rect 6 247 7 248
rect 5 247 6 248
rect 4 247 5 248
rect 3 247 4 248
rect 2 247 3 248
rect 1 247 2 248
rect 479 248 480 249
rect 478 248 479 249
rect 470 248 471 249
rect 469 248 470 249
rect 468 248 469 249
rect 467 248 468 249
rect 466 248 467 249
rect 465 248 466 249
rect 458 248 459 249
rect 457 248 458 249
rect 419 248 420 249
rect 418 248 419 249
rect 417 248 418 249
rect 416 248 417 249
rect 314 248 315 249
rect 313 248 314 249
rect 312 248 313 249
rect 311 248 312 249
rect 310 248 311 249
rect 309 248 310 249
rect 308 248 309 249
rect 307 248 308 249
rect 306 248 307 249
rect 305 248 306 249
rect 304 248 305 249
rect 303 248 304 249
rect 302 248 303 249
rect 301 248 302 249
rect 300 248 301 249
rect 299 248 300 249
rect 298 248 299 249
rect 297 248 298 249
rect 296 248 297 249
rect 295 248 296 249
rect 294 248 295 249
rect 293 248 294 249
rect 292 248 293 249
rect 291 248 292 249
rect 290 248 291 249
rect 289 248 290 249
rect 288 248 289 249
rect 287 248 288 249
rect 286 248 287 249
rect 285 248 286 249
rect 284 248 285 249
rect 283 248 284 249
rect 282 248 283 249
rect 281 248 282 249
rect 280 248 281 249
rect 279 248 280 249
rect 278 248 279 249
rect 277 248 278 249
rect 276 248 277 249
rect 275 248 276 249
rect 274 248 275 249
rect 273 248 274 249
rect 272 248 273 249
rect 271 248 272 249
rect 270 248 271 249
rect 269 248 270 249
rect 268 248 269 249
rect 267 248 268 249
rect 266 248 267 249
rect 265 248 266 249
rect 264 248 265 249
rect 263 248 264 249
rect 262 248 263 249
rect 261 248 262 249
rect 260 248 261 249
rect 259 248 260 249
rect 258 248 259 249
rect 257 248 258 249
rect 256 248 257 249
rect 255 248 256 249
rect 254 248 255 249
rect 253 248 254 249
rect 252 248 253 249
rect 251 248 252 249
rect 250 248 251 249
rect 249 248 250 249
rect 248 248 249 249
rect 247 248 248 249
rect 246 248 247 249
rect 245 248 246 249
rect 244 248 245 249
rect 243 248 244 249
rect 242 248 243 249
rect 241 248 242 249
rect 240 248 241 249
rect 239 248 240 249
rect 238 248 239 249
rect 237 248 238 249
rect 236 248 237 249
rect 235 248 236 249
rect 234 248 235 249
rect 233 248 234 249
rect 232 248 233 249
rect 231 248 232 249
rect 230 248 231 249
rect 229 248 230 249
rect 156 248 157 249
rect 155 248 156 249
rect 154 248 155 249
rect 153 248 154 249
rect 152 248 153 249
rect 151 248 152 249
rect 150 248 151 249
rect 149 248 150 249
rect 148 248 149 249
rect 147 248 148 249
rect 146 248 147 249
rect 145 248 146 249
rect 144 248 145 249
rect 143 248 144 249
rect 142 248 143 249
rect 141 248 142 249
rect 140 248 141 249
rect 139 248 140 249
rect 138 248 139 249
rect 137 248 138 249
rect 136 248 137 249
rect 135 248 136 249
rect 134 248 135 249
rect 133 248 134 249
rect 132 248 133 249
rect 131 248 132 249
rect 130 248 131 249
rect 129 248 130 249
rect 128 248 129 249
rect 127 248 128 249
rect 126 248 127 249
rect 125 248 126 249
rect 124 248 125 249
rect 123 248 124 249
rect 122 248 123 249
rect 121 248 122 249
rect 120 248 121 249
rect 119 248 120 249
rect 106 248 107 249
rect 105 248 106 249
rect 104 248 105 249
rect 103 248 104 249
rect 102 248 103 249
rect 101 248 102 249
rect 100 248 101 249
rect 99 248 100 249
rect 98 248 99 249
rect 97 248 98 249
rect 96 248 97 249
rect 95 248 96 249
rect 94 248 95 249
rect 93 248 94 249
rect 92 248 93 249
rect 91 248 92 249
rect 90 248 91 249
rect 89 248 90 249
rect 88 248 89 249
rect 87 248 88 249
rect 86 248 87 249
rect 85 248 86 249
rect 84 248 85 249
rect 83 248 84 249
rect 82 248 83 249
rect 81 248 82 249
rect 80 248 81 249
rect 79 248 80 249
rect 78 248 79 249
rect 77 248 78 249
rect 76 248 77 249
rect 75 248 76 249
rect 74 248 75 249
rect 73 248 74 249
rect 72 248 73 249
rect 71 248 72 249
rect 70 248 71 249
rect 69 248 70 249
rect 68 248 69 249
rect 67 248 68 249
rect 66 248 67 249
rect 65 248 66 249
rect 64 248 65 249
rect 63 248 64 249
rect 62 248 63 249
rect 61 248 62 249
rect 60 248 61 249
rect 59 248 60 249
rect 58 248 59 249
rect 57 248 58 249
rect 56 248 57 249
rect 55 248 56 249
rect 54 248 55 249
rect 53 248 54 249
rect 52 248 53 249
rect 51 248 52 249
rect 50 248 51 249
rect 49 248 50 249
rect 48 248 49 249
rect 47 248 48 249
rect 46 248 47 249
rect 45 248 46 249
rect 44 248 45 249
rect 43 248 44 249
rect 42 248 43 249
rect 41 248 42 249
rect 40 248 41 249
rect 39 248 40 249
rect 38 248 39 249
rect 37 248 38 249
rect 36 248 37 249
rect 35 248 36 249
rect 34 248 35 249
rect 33 248 34 249
rect 32 248 33 249
rect 31 248 32 249
rect 30 248 31 249
rect 29 248 30 249
rect 19 248 20 249
rect 18 248 19 249
rect 17 248 18 249
rect 16 248 17 249
rect 15 248 16 249
rect 14 248 15 249
rect 13 248 14 249
rect 12 248 13 249
rect 11 248 12 249
rect 10 248 11 249
rect 9 248 10 249
rect 8 248 9 249
rect 7 248 8 249
rect 6 248 7 249
rect 5 248 6 249
rect 4 248 5 249
rect 3 248 4 249
rect 2 248 3 249
rect 1 248 2 249
rect 479 249 480 250
rect 478 249 479 250
rect 470 249 471 250
rect 469 249 470 250
rect 468 249 469 250
rect 467 249 468 250
rect 466 249 467 250
rect 458 249 459 250
rect 457 249 458 250
rect 418 249 419 250
rect 417 249 418 250
rect 416 249 417 250
rect 313 249 314 250
rect 312 249 313 250
rect 311 249 312 250
rect 310 249 311 250
rect 309 249 310 250
rect 308 249 309 250
rect 307 249 308 250
rect 306 249 307 250
rect 305 249 306 250
rect 304 249 305 250
rect 303 249 304 250
rect 302 249 303 250
rect 301 249 302 250
rect 300 249 301 250
rect 299 249 300 250
rect 298 249 299 250
rect 297 249 298 250
rect 296 249 297 250
rect 295 249 296 250
rect 294 249 295 250
rect 293 249 294 250
rect 292 249 293 250
rect 291 249 292 250
rect 290 249 291 250
rect 289 249 290 250
rect 288 249 289 250
rect 287 249 288 250
rect 286 249 287 250
rect 285 249 286 250
rect 284 249 285 250
rect 283 249 284 250
rect 282 249 283 250
rect 281 249 282 250
rect 280 249 281 250
rect 279 249 280 250
rect 278 249 279 250
rect 277 249 278 250
rect 276 249 277 250
rect 275 249 276 250
rect 274 249 275 250
rect 273 249 274 250
rect 272 249 273 250
rect 271 249 272 250
rect 270 249 271 250
rect 269 249 270 250
rect 268 249 269 250
rect 267 249 268 250
rect 266 249 267 250
rect 265 249 266 250
rect 264 249 265 250
rect 263 249 264 250
rect 262 249 263 250
rect 261 249 262 250
rect 260 249 261 250
rect 259 249 260 250
rect 258 249 259 250
rect 257 249 258 250
rect 256 249 257 250
rect 255 249 256 250
rect 254 249 255 250
rect 253 249 254 250
rect 252 249 253 250
rect 251 249 252 250
rect 250 249 251 250
rect 249 249 250 250
rect 248 249 249 250
rect 247 249 248 250
rect 246 249 247 250
rect 245 249 246 250
rect 244 249 245 250
rect 243 249 244 250
rect 242 249 243 250
rect 241 249 242 250
rect 240 249 241 250
rect 239 249 240 250
rect 238 249 239 250
rect 237 249 238 250
rect 236 249 237 250
rect 235 249 236 250
rect 234 249 235 250
rect 233 249 234 250
rect 232 249 233 250
rect 231 249 232 250
rect 230 249 231 250
rect 229 249 230 250
rect 157 249 158 250
rect 156 249 157 250
rect 155 249 156 250
rect 154 249 155 250
rect 153 249 154 250
rect 152 249 153 250
rect 151 249 152 250
rect 150 249 151 250
rect 149 249 150 250
rect 148 249 149 250
rect 147 249 148 250
rect 146 249 147 250
rect 145 249 146 250
rect 144 249 145 250
rect 143 249 144 250
rect 142 249 143 250
rect 141 249 142 250
rect 140 249 141 250
rect 139 249 140 250
rect 138 249 139 250
rect 137 249 138 250
rect 136 249 137 250
rect 135 249 136 250
rect 134 249 135 250
rect 133 249 134 250
rect 132 249 133 250
rect 131 249 132 250
rect 130 249 131 250
rect 129 249 130 250
rect 128 249 129 250
rect 127 249 128 250
rect 126 249 127 250
rect 125 249 126 250
rect 124 249 125 250
rect 123 249 124 250
rect 122 249 123 250
rect 121 249 122 250
rect 120 249 121 250
rect 119 249 120 250
rect 106 249 107 250
rect 105 249 106 250
rect 104 249 105 250
rect 103 249 104 250
rect 102 249 103 250
rect 101 249 102 250
rect 100 249 101 250
rect 99 249 100 250
rect 98 249 99 250
rect 97 249 98 250
rect 96 249 97 250
rect 95 249 96 250
rect 94 249 95 250
rect 93 249 94 250
rect 92 249 93 250
rect 91 249 92 250
rect 90 249 91 250
rect 89 249 90 250
rect 88 249 89 250
rect 87 249 88 250
rect 86 249 87 250
rect 85 249 86 250
rect 84 249 85 250
rect 83 249 84 250
rect 82 249 83 250
rect 81 249 82 250
rect 80 249 81 250
rect 79 249 80 250
rect 78 249 79 250
rect 77 249 78 250
rect 76 249 77 250
rect 75 249 76 250
rect 74 249 75 250
rect 73 249 74 250
rect 72 249 73 250
rect 71 249 72 250
rect 70 249 71 250
rect 69 249 70 250
rect 68 249 69 250
rect 67 249 68 250
rect 66 249 67 250
rect 65 249 66 250
rect 64 249 65 250
rect 63 249 64 250
rect 62 249 63 250
rect 61 249 62 250
rect 60 249 61 250
rect 59 249 60 250
rect 58 249 59 250
rect 57 249 58 250
rect 56 249 57 250
rect 55 249 56 250
rect 54 249 55 250
rect 53 249 54 250
rect 52 249 53 250
rect 51 249 52 250
rect 50 249 51 250
rect 49 249 50 250
rect 48 249 49 250
rect 47 249 48 250
rect 46 249 47 250
rect 45 249 46 250
rect 44 249 45 250
rect 43 249 44 250
rect 42 249 43 250
rect 41 249 42 250
rect 40 249 41 250
rect 39 249 40 250
rect 38 249 39 250
rect 37 249 38 250
rect 36 249 37 250
rect 35 249 36 250
rect 34 249 35 250
rect 33 249 34 250
rect 32 249 33 250
rect 31 249 32 250
rect 30 249 31 250
rect 29 249 30 250
rect 19 249 20 250
rect 18 249 19 250
rect 17 249 18 250
rect 16 249 17 250
rect 15 249 16 250
rect 14 249 15 250
rect 13 249 14 250
rect 12 249 13 250
rect 11 249 12 250
rect 10 249 11 250
rect 9 249 10 250
rect 8 249 9 250
rect 7 249 8 250
rect 6 249 7 250
rect 5 249 6 250
rect 4 249 5 250
rect 3 249 4 250
rect 2 249 3 250
rect 1 249 2 250
rect 479 250 480 251
rect 478 250 479 251
rect 471 250 472 251
rect 470 250 471 251
rect 469 250 470 251
rect 468 250 469 251
rect 467 250 468 251
rect 466 250 467 251
rect 458 250 459 251
rect 457 250 458 251
rect 418 250 419 251
rect 417 250 418 251
rect 311 250 312 251
rect 310 250 311 251
rect 309 250 310 251
rect 308 250 309 251
rect 307 250 308 251
rect 306 250 307 251
rect 305 250 306 251
rect 304 250 305 251
rect 303 250 304 251
rect 302 250 303 251
rect 301 250 302 251
rect 300 250 301 251
rect 299 250 300 251
rect 298 250 299 251
rect 297 250 298 251
rect 296 250 297 251
rect 295 250 296 251
rect 294 250 295 251
rect 293 250 294 251
rect 292 250 293 251
rect 291 250 292 251
rect 290 250 291 251
rect 289 250 290 251
rect 288 250 289 251
rect 287 250 288 251
rect 286 250 287 251
rect 285 250 286 251
rect 284 250 285 251
rect 283 250 284 251
rect 282 250 283 251
rect 281 250 282 251
rect 280 250 281 251
rect 279 250 280 251
rect 278 250 279 251
rect 277 250 278 251
rect 276 250 277 251
rect 275 250 276 251
rect 274 250 275 251
rect 273 250 274 251
rect 272 250 273 251
rect 271 250 272 251
rect 270 250 271 251
rect 269 250 270 251
rect 268 250 269 251
rect 267 250 268 251
rect 266 250 267 251
rect 265 250 266 251
rect 264 250 265 251
rect 263 250 264 251
rect 262 250 263 251
rect 261 250 262 251
rect 260 250 261 251
rect 259 250 260 251
rect 258 250 259 251
rect 257 250 258 251
rect 256 250 257 251
rect 255 250 256 251
rect 254 250 255 251
rect 253 250 254 251
rect 252 250 253 251
rect 251 250 252 251
rect 250 250 251 251
rect 249 250 250 251
rect 248 250 249 251
rect 247 250 248 251
rect 246 250 247 251
rect 245 250 246 251
rect 244 250 245 251
rect 243 250 244 251
rect 242 250 243 251
rect 241 250 242 251
rect 240 250 241 251
rect 239 250 240 251
rect 238 250 239 251
rect 237 250 238 251
rect 236 250 237 251
rect 235 250 236 251
rect 234 250 235 251
rect 233 250 234 251
rect 232 250 233 251
rect 231 250 232 251
rect 230 250 231 251
rect 229 250 230 251
rect 158 250 159 251
rect 157 250 158 251
rect 156 250 157 251
rect 155 250 156 251
rect 154 250 155 251
rect 153 250 154 251
rect 152 250 153 251
rect 151 250 152 251
rect 150 250 151 251
rect 149 250 150 251
rect 148 250 149 251
rect 147 250 148 251
rect 146 250 147 251
rect 145 250 146 251
rect 144 250 145 251
rect 143 250 144 251
rect 142 250 143 251
rect 141 250 142 251
rect 140 250 141 251
rect 139 250 140 251
rect 138 250 139 251
rect 137 250 138 251
rect 136 250 137 251
rect 135 250 136 251
rect 134 250 135 251
rect 133 250 134 251
rect 132 250 133 251
rect 131 250 132 251
rect 130 250 131 251
rect 129 250 130 251
rect 128 250 129 251
rect 127 250 128 251
rect 126 250 127 251
rect 125 250 126 251
rect 124 250 125 251
rect 123 250 124 251
rect 122 250 123 251
rect 121 250 122 251
rect 120 250 121 251
rect 119 250 120 251
rect 106 250 107 251
rect 105 250 106 251
rect 104 250 105 251
rect 103 250 104 251
rect 102 250 103 251
rect 101 250 102 251
rect 100 250 101 251
rect 99 250 100 251
rect 98 250 99 251
rect 97 250 98 251
rect 96 250 97 251
rect 95 250 96 251
rect 94 250 95 251
rect 93 250 94 251
rect 92 250 93 251
rect 91 250 92 251
rect 90 250 91 251
rect 89 250 90 251
rect 88 250 89 251
rect 87 250 88 251
rect 86 250 87 251
rect 85 250 86 251
rect 84 250 85 251
rect 83 250 84 251
rect 82 250 83 251
rect 81 250 82 251
rect 80 250 81 251
rect 79 250 80 251
rect 78 250 79 251
rect 77 250 78 251
rect 76 250 77 251
rect 75 250 76 251
rect 74 250 75 251
rect 73 250 74 251
rect 72 250 73 251
rect 71 250 72 251
rect 70 250 71 251
rect 69 250 70 251
rect 68 250 69 251
rect 67 250 68 251
rect 66 250 67 251
rect 65 250 66 251
rect 64 250 65 251
rect 63 250 64 251
rect 62 250 63 251
rect 61 250 62 251
rect 60 250 61 251
rect 59 250 60 251
rect 58 250 59 251
rect 57 250 58 251
rect 56 250 57 251
rect 55 250 56 251
rect 54 250 55 251
rect 53 250 54 251
rect 52 250 53 251
rect 51 250 52 251
rect 50 250 51 251
rect 49 250 50 251
rect 48 250 49 251
rect 47 250 48 251
rect 46 250 47 251
rect 45 250 46 251
rect 44 250 45 251
rect 43 250 44 251
rect 42 250 43 251
rect 41 250 42 251
rect 40 250 41 251
rect 39 250 40 251
rect 38 250 39 251
rect 37 250 38 251
rect 36 250 37 251
rect 35 250 36 251
rect 34 250 35 251
rect 33 250 34 251
rect 32 250 33 251
rect 31 250 32 251
rect 30 250 31 251
rect 19 250 20 251
rect 18 250 19 251
rect 17 250 18 251
rect 16 250 17 251
rect 15 250 16 251
rect 14 250 15 251
rect 13 250 14 251
rect 12 250 13 251
rect 11 250 12 251
rect 10 250 11 251
rect 9 250 10 251
rect 8 250 9 251
rect 7 250 8 251
rect 6 250 7 251
rect 5 250 6 251
rect 4 250 5 251
rect 3 250 4 251
rect 2 250 3 251
rect 1 250 2 251
rect 478 251 479 252
rect 477 251 478 252
rect 472 251 473 252
rect 471 251 472 252
rect 470 251 471 252
rect 469 251 470 252
rect 468 251 469 252
rect 467 251 468 252
rect 458 251 459 252
rect 457 251 458 252
rect 310 251 311 252
rect 309 251 310 252
rect 308 251 309 252
rect 307 251 308 252
rect 306 251 307 252
rect 305 251 306 252
rect 304 251 305 252
rect 303 251 304 252
rect 302 251 303 252
rect 301 251 302 252
rect 300 251 301 252
rect 299 251 300 252
rect 298 251 299 252
rect 297 251 298 252
rect 296 251 297 252
rect 295 251 296 252
rect 294 251 295 252
rect 293 251 294 252
rect 292 251 293 252
rect 291 251 292 252
rect 290 251 291 252
rect 289 251 290 252
rect 288 251 289 252
rect 287 251 288 252
rect 286 251 287 252
rect 285 251 286 252
rect 284 251 285 252
rect 283 251 284 252
rect 282 251 283 252
rect 281 251 282 252
rect 280 251 281 252
rect 279 251 280 252
rect 278 251 279 252
rect 277 251 278 252
rect 276 251 277 252
rect 275 251 276 252
rect 274 251 275 252
rect 273 251 274 252
rect 272 251 273 252
rect 271 251 272 252
rect 270 251 271 252
rect 269 251 270 252
rect 268 251 269 252
rect 267 251 268 252
rect 266 251 267 252
rect 265 251 266 252
rect 264 251 265 252
rect 263 251 264 252
rect 262 251 263 252
rect 261 251 262 252
rect 260 251 261 252
rect 259 251 260 252
rect 258 251 259 252
rect 257 251 258 252
rect 256 251 257 252
rect 255 251 256 252
rect 254 251 255 252
rect 253 251 254 252
rect 252 251 253 252
rect 251 251 252 252
rect 250 251 251 252
rect 249 251 250 252
rect 248 251 249 252
rect 247 251 248 252
rect 246 251 247 252
rect 245 251 246 252
rect 244 251 245 252
rect 243 251 244 252
rect 242 251 243 252
rect 241 251 242 252
rect 240 251 241 252
rect 239 251 240 252
rect 238 251 239 252
rect 237 251 238 252
rect 236 251 237 252
rect 235 251 236 252
rect 234 251 235 252
rect 233 251 234 252
rect 232 251 233 252
rect 231 251 232 252
rect 230 251 231 252
rect 229 251 230 252
rect 228 251 229 252
rect 160 251 161 252
rect 159 251 160 252
rect 158 251 159 252
rect 157 251 158 252
rect 156 251 157 252
rect 155 251 156 252
rect 154 251 155 252
rect 153 251 154 252
rect 152 251 153 252
rect 151 251 152 252
rect 150 251 151 252
rect 149 251 150 252
rect 148 251 149 252
rect 147 251 148 252
rect 146 251 147 252
rect 145 251 146 252
rect 144 251 145 252
rect 143 251 144 252
rect 142 251 143 252
rect 141 251 142 252
rect 140 251 141 252
rect 139 251 140 252
rect 138 251 139 252
rect 137 251 138 252
rect 136 251 137 252
rect 135 251 136 252
rect 134 251 135 252
rect 133 251 134 252
rect 132 251 133 252
rect 131 251 132 252
rect 130 251 131 252
rect 129 251 130 252
rect 128 251 129 252
rect 127 251 128 252
rect 126 251 127 252
rect 125 251 126 252
rect 124 251 125 252
rect 123 251 124 252
rect 122 251 123 252
rect 121 251 122 252
rect 120 251 121 252
rect 119 251 120 252
rect 106 251 107 252
rect 105 251 106 252
rect 104 251 105 252
rect 103 251 104 252
rect 102 251 103 252
rect 101 251 102 252
rect 100 251 101 252
rect 99 251 100 252
rect 98 251 99 252
rect 97 251 98 252
rect 96 251 97 252
rect 95 251 96 252
rect 94 251 95 252
rect 93 251 94 252
rect 92 251 93 252
rect 91 251 92 252
rect 90 251 91 252
rect 89 251 90 252
rect 88 251 89 252
rect 87 251 88 252
rect 86 251 87 252
rect 85 251 86 252
rect 84 251 85 252
rect 83 251 84 252
rect 82 251 83 252
rect 81 251 82 252
rect 80 251 81 252
rect 79 251 80 252
rect 78 251 79 252
rect 77 251 78 252
rect 76 251 77 252
rect 75 251 76 252
rect 74 251 75 252
rect 73 251 74 252
rect 72 251 73 252
rect 71 251 72 252
rect 70 251 71 252
rect 69 251 70 252
rect 68 251 69 252
rect 67 251 68 252
rect 66 251 67 252
rect 65 251 66 252
rect 64 251 65 252
rect 63 251 64 252
rect 62 251 63 252
rect 61 251 62 252
rect 60 251 61 252
rect 59 251 60 252
rect 58 251 59 252
rect 57 251 58 252
rect 56 251 57 252
rect 55 251 56 252
rect 54 251 55 252
rect 53 251 54 252
rect 52 251 53 252
rect 51 251 52 252
rect 50 251 51 252
rect 49 251 50 252
rect 48 251 49 252
rect 47 251 48 252
rect 46 251 47 252
rect 45 251 46 252
rect 44 251 45 252
rect 43 251 44 252
rect 42 251 43 252
rect 41 251 42 252
rect 40 251 41 252
rect 39 251 40 252
rect 38 251 39 252
rect 37 251 38 252
rect 36 251 37 252
rect 35 251 36 252
rect 34 251 35 252
rect 33 251 34 252
rect 32 251 33 252
rect 31 251 32 252
rect 30 251 31 252
rect 19 251 20 252
rect 18 251 19 252
rect 17 251 18 252
rect 16 251 17 252
rect 15 251 16 252
rect 14 251 15 252
rect 13 251 14 252
rect 12 251 13 252
rect 11 251 12 252
rect 10 251 11 252
rect 9 251 10 252
rect 8 251 9 252
rect 7 251 8 252
rect 6 251 7 252
rect 5 251 6 252
rect 4 251 5 252
rect 3 251 4 252
rect 2 251 3 252
rect 1 251 2 252
rect 478 252 479 253
rect 477 252 478 253
rect 476 252 477 253
rect 475 252 476 253
rect 474 252 475 253
rect 473 252 474 253
rect 472 252 473 253
rect 471 252 472 253
rect 470 252 471 253
rect 469 252 470 253
rect 468 252 469 253
rect 467 252 468 253
rect 459 252 460 253
rect 458 252 459 253
rect 457 252 458 253
rect 309 252 310 253
rect 308 252 309 253
rect 307 252 308 253
rect 306 252 307 253
rect 305 252 306 253
rect 304 252 305 253
rect 303 252 304 253
rect 302 252 303 253
rect 301 252 302 253
rect 300 252 301 253
rect 299 252 300 253
rect 298 252 299 253
rect 297 252 298 253
rect 296 252 297 253
rect 295 252 296 253
rect 294 252 295 253
rect 293 252 294 253
rect 292 252 293 253
rect 291 252 292 253
rect 290 252 291 253
rect 289 252 290 253
rect 288 252 289 253
rect 287 252 288 253
rect 286 252 287 253
rect 285 252 286 253
rect 284 252 285 253
rect 283 252 284 253
rect 282 252 283 253
rect 281 252 282 253
rect 280 252 281 253
rect 279 252 280 253
rect 278 252 279 253
rect 277 252 278 253
rect 276 252 277 253
rect 275 252 276 253
rect 274 252 275 253
rect 273 252 274 253
rect 272 252 273 253
rect 271 252 272 253
rect 270 252 271 253
rect 269 252 270 253
rect 268 252 269 253
rect 267 252 268 253
rect 266 252 267 253
rect 265 252 266 253
rect 264 252 265 253
rect 263 252 264 253
rect 262 252 263 253
rect 261 252 262 253
rect 260 252 261 253
rect 259 252 260 253
rect 258 252 259 253
rect 257 252 258 253
rect 256 252 257 253
rect 255 252 256 253
rect 254 252 255 253
rect 253 252 254 253
rect 252 252 253 253
rect 251 252 252 253
rect 250 252 251 253
rect 249 252 250 253
rect 248 252 249 253
rect 247 252 248 253
rect 246 252 247 253
rect 245 252 246 253
rect 244 252 245 253
rect 243 252 244 253
rect 242 252 243 253
rect 241 252 242 253
rect 240 252 241 253
rect 239 252 240 253
rect 238 252 239 253
rect 237 252 238 253
rect 236 252 237 253
rect 235 252 236 253
rect 234 252 235 253
rect 233 252 234 253
rect 232 252 233 253
rect 231 252 232 253
rect 230 252 231 253
rect 229 252 230 253
rect 228 252 229 253
rect 162 252 163 253
rect 161 252 162 253
rect 160 252 161 253
rect 159 252 160 253
rect 158 252 159 253
rect 157 252 158 253
rect 156 252 157 253
rect 155 252 156 253
rect 154 252 155 253
rect 153 252 154 253
rect 152 252 153 253
rect 151 252 152 253
rect 150 252 151 253
rect 149 252 150 253
rect 148 252 149 253
rect 147 252 148 253
rect 146 252 147 253
rect 145 252 146 253
rect 144 252 145 253
rect 143 252 144 253
rect 142 252 143 253
rect 141 252 142 253
rect 140 252 141 253
rect 139 252 140 253
rect 138 252 139 253
rect 137 252 138 253
rect 136 252 137 253
rect 135 252 136 253
rect 134 252 135 253
rect 133 252 134 253
rect 132 252 133 253
rect 131 252 132 253
rect 130 252 131 253
rect 129 252 130 253
rect 128 252 129 253
rect 127 252 128 253
rect 126 252 127 253
rect 125 252 126 253
rect 124 252 125 253
rect 123 252 124 253
rect 122 252 123 253
rect 121 252 122 253
rect 120 252 121 253
rect 119 252 120 253
rect 107 252 108 253
rect 106 252 107 253
rect 105 252 106 253
rect 104 252 105 253
rect 103 252 104 253
rect 102 252 103 253
rect 101 252 102 253
rect 100 252 101 253
rect 99 252 100 253
rect 98 252 99 253
rect 97 252 98 253
rect 96 252 97 253
rect 95 252 96 253
rect 94 252 95 253
rect 93 252 94 253
rect 92 252 93 253
rect 91 252 92 253
rect 90 252 91 253
rect 89 252 90 253
rect 88 252 89 253
rect 87 252 88 253
rect 86 252 87 253
rect 85 252 86 253
rect 84 252 85 253
rect 83 252 84 253
rect 82 252 83 253
rect 81 252 82 253
rect 80 252 81 253
rect 79 252 80 253
rect 78 252 79 253
rect 77 252 78 253
rect 76 252 77 253
rect 75 252 76 253
rect 74 252 75 253
rect 73 252 74 253
rect 72 252 73 253
rect 71 252 72 253
rect 70 252 71 253
rect 69 252 70 253
rect 68 252 69 253
rect 67 252 68 253
rect 66 252 67 253
rect 65 252 66 253
rect 64 252 65 253
rect 63 252 64 253
rect 62 252 63 253
rect 61 252 62 253
rect 60 252 61 253
rect 59 252 60 253
rect 58 252 59 253
rect 57 252 58 253
rect 56 252 57 253
rect 52 252 53 253
rect 51 252 52 253
rect 50 252 51 253
rect 49 252 50 253
rect 48 252 49 253
rect 47 252 48 253
rect 46 252 47 253
rect 45 252 46 253
rect 44 252 45 253
rect 43 252 44 253
rect 42 252 43 253
rect 41 252 42 253
rect 40 252 41 253
rect 39 252 40 253
rect 38 252 39 253
rect 37 252 38 253
rect 36 252 37 253
rect 35 252 36 253
rect 34 252 35 253
rect 33 252 34 253
rect 32 252 33 253
rect 31 252 32 253
rect 30 252 31 253
rect 20 252 21 253
rect 19 252 20 253
rect 18 252 19 253
rect 17 252 18 253
rect 16 252 17 253
rect 15 252 16 253
rect 14 252 15 253
rect 13 252 14 253
rect 12 252 13 253
rect 11 252 12 253
rect 10 252 11 253
rect 9 252 10 253
rect 8 252 9 253
rect 7 252 8 253
rect 6 252 7 253
rect 5 252 6 253
rect 4 252 5 253
rect 3 252 4 253
rect 2 252 3 253
rect 1 252 2 253
rect 477 253 478 254
rect 476 253 477 254
rect 475 253 476 254
rect 474 253 475 254
rect 473 253 474 254
rect 472 253 473 254
rect 471 253 472 254
rect 470 253 471 254
rect 469 253 470 254
rect 468 253 469 254
rect 461 253 462 254
rect 460 253 461 254
rect 459 253 460 254
rect 458 253 459 254
rect 307 253 308 254
rect 306 253 307 254
rect 305 253 306 254
rect 304 253 305 254
rect 303 253 304 254
rect 302 253 303 254
rect 301 253 302 254
rect 300 253 301 254
rect 299 253 300 254
rect 298 253 299 254
rect 297 253 298 254
rect 296 253 297 254
rect 295 253 296 254
rect 294 253 295 254
rect 293 253 294 254
rect 292 253 293 254
rect 291 253 292 254
rect 290 253 291 254
rect 289 253 290 254
rect 288 253 289 254
rect 287 253 288 254
rect 286 253 287 254
rect 285 253 286 254
rect 284 253 285 254
rect 283 253 284 254
rect 282 253 283 254
rect 281 253 282 254
rect 280 253 281 254
rect 279 253 280 254
rect 278 253 279 254
rect 277 253 278 254
rect 276 253 277 254
rect 275 253 276 254
rect 274 253 275 254
rect 273 253 274 254
rect 272 253 273 254
rect 271 253 272 254
rect 270 253 271 254
rect 269 253 270 254
rect 268 253 269 254
rect 267 253 268 254
rect 266 253 267 254
rect 265 253 266 254
rect 264 253 265 254
rect 263 253 264 254
rect 262 253 263 254
rect 261 253 262 254
rect 260 253 261 254
rect 259 253 260 254
rect 258 253 259 254
rect 257 253 258 254
rect 256 253 257 254
rect 255 253 256 254
rect 254 253 255 254
rect 253 253 254 254
rect 252 253 253 254
rect 251 253 252 254
rect 250 253 251 254
rect 249 253 250 254
rect 248 253 249 254
rect 247 253 248 254
rect 246 253 247 254
rect 245 253 246 254
rect 244 253 245 254
rect 243 253 244 254
rect 242 253 243 254
rect 241 253 242 254
rect 240 253 241 254
rect 239 253 240 254
rect 238 253 239 254
rect 237 253 238 254
rect 236 253 237 254
rect 235 253 236 254
rect 234 253 235 254
rect 233 253 234 254
rect 232 253 233 254
rect 231 253 232 254
rect 230 253 231 254
rect 229 253 230 254
rect 228 253 229 254
rect 164 253 165 254
rect 163 253 164 254
rect 162 253 163 254
rect 161 253 162 254
rect 160 253 161 254
rect 159 253 160 254
rect 158 253 159 254
rect 157 253 158 254
rect 156 253 157 254
rect 155 253 156 254
rect 154 253 155 254
rect 153 253 154 254
rect 152 253 153 254
rect 151 253 152 254
rect 150 253 151 254
rect 149 253 150 254
rect 148 253 149 254
rect 147 253 148 254
rect 146 253 147 254
rect 145 253 146 254
rect 144 253 145 254
rect 143 253 144 254
rect 142 253 143 254
rect 141 253 142 254
rect 140 253 141 254
rect 139 253 140 254
rect 138 253 139 254
rect 137 253 138 254
rect 136 253 137 254
rect 135 253 136 254
rect 134 253 135 254
rect 133 253 134 254
rect 132 253 133 254
rect 131 253 132 254
rect 130 253 131 254
rect 129 253 130 254
rect 128 253 129 254
rect 127 253 128 254
rect 126 253 127 254
rect 125 253 126 254
rect 124 253 125 254
rect 123 253 124 254
rect 122 253 123 254
rect 121 253 122 254
rect 120 253 121 254
rect 107 253 108 254
rect 106 253 107 254
rect 105 253 106 254
rect 104 253 105 254
rect 103 253 104 254
rect 102 253 103 254
rect 101 253 102 254
rect 100 253 101 254
rect 99 253 100 254
rect 98 253 99 254
rect 97 253 98 254
rect 96 253 97 254
rect 95 253 96 254
rect 94 253 95 254
rect 93 253 94 254
rect 92 253 93 254
rect 91 253 92 254
rect 90 253 91 254
rect 89 253 90 254
rect 88 253 89 254
rect 87 253 88 254
rect 86 253 87 254
rect 85 253 86 254
rect 84 253 85 254
rect 83 253 84 254
rect 82 253 83 254
rect 81 253 82 254
rect 80 253 81 254
rect 79 253 80 254
rect 78 253 79 254
rect 77 253 78 254
rect 76 253 77 254
rect 75 253 76 254
rect 74 253 75 254
rect 73 253 74 254
rect 72 253 73 254
rect 71 253 72 254
rect 70 253 71 254
rect 69 253 70 254
rect 68 253 69 254
rect 67 253 68 254
rect 66 253 67 254
rect 65 253 66 254
rect 64 253 65 254
rect 63 253 64 254
rect 62 253 63 254
rect 61 253 62 254
rect 52 253 53 254
rect 51 253 52 254
rect 50 253 51 254
rect 49 253 50 254
rect 48 253 49 254
rect 47 253 48 254
rect 46 253 47 254
rect 45 253 46 254
rect 44 253 45 254
rect 43 253 44 254
rect 42 253 43 254
rect 41 253 42 254
rect 40 253 41 254
rect 39 253 40 254
rect 38 253 39 254
rect 37 253 38 254
rect 36 253 37 254
rect 35 253 36 254
rect 34 253 35 254
rect 33 253 34 254
rect 32 253 33 254
rect 31 253 32 254
rect 20 253 21 254
rect 19 253 20 254
rect 18 253 19 254
rect 17 253 18 254
rect 16 253 17 254
rect 15 253 16 254
rect 14 253 15 254
rect 13 253 14 254
rect 12 253 13 254
rect 11 253 12 254
rect 10 253 11 254
rect 9 253 10 254
rect 8 253 9 254
rect 7 253 8 254
rect 6 253 7 254
rect 5 253 6 254
rect 4 253 5 254
rect 3 253 4 254
rect 2 253 3 254
rect 1 253 2 254
rect 476 254 477 255
rect 475 254 476 255
rect 474 254 475 255
rect 473 254 474 255
rect 472 254 473 255
rect 471 254 472 255
rect 470 254 471 255
rect 469 254 470 255
rect 462 254 463 255
rect 461 254 462 255
rect 460 254 461 255
rect 459 254 460 255
rect 458 254 459 255
rect 306 254 307 255
rect 305 254 306 255
rect 304 254 305 255
rect 303 254 304 255
rect 302 254 303 255
rect 301 254 302 255
rect 300 254 301 255
rect 299 254 300 255
rect 298 254 299 255
rect 297 254 298 255
rect 296 254 297 255
rect 295 254 296 255
rect 294 254 295 255
rect 293 254 294 255
rect 292 254 293 255
rect 291 254 292 255
rect 290 254 291 255
rect 289 254 290 255
rect 288 254 289 255
rect 287 254 288 255
rect 286 254 287 255
rect 285 254 286 255
rect 284 254 285 255
rect 283 254 284 255
rect 282 254 283 255
rect 281 254 282 255
rect 280 254 281 255
rect 279 254 280 255
rect 278 254 279 255
rect 277 254 278 255
rect 276 254 277 255
rect 275 254 276 255
rect 274 254 275 255
rect 273 254 274 255
rect 272 254 273 255
rect 271 254 272 255
rect 270 254 271 255
rect 269 254 270 255
rect 268 254 269 255
rect 267 254 268 255
rect 266 254 267 255
rect 265 254 266 255
rect 264 254 265 255
rect 263 254 264 255
rect 262 254 263 255
rect 261 254 262 255
rect 260 254 261 255
rect 259 254 260 255
rect 258 254 259 255
rect 257 254 258 255
rect 256 254 257 255
rect 255 254 256 255
rect 254 254 255 255
rect 253 254 254 255
rect 252 254 253 255
rect 251 254 252 255
rect 250 254 251 255
rect 249 254 250 255
rect 248 254 249 255
rect 247 254 248 255
rect 246 254 247 255
rect 245 254 246 255
rect 244 254 245 255
rect 243 254 244 255
rect 242 254 243 255
rect 241 254 242 255
rect 240 254 241 255
rect 239 254 240 255
rect 238 254 239 255
rect 237 254 238 255
rect 236 254 237 255
rect 235 254 236 255
rect 234 254 235 255
rect 233 254 234 255
rect 232 254 233 255
rect 231 254 232 255
rect 230 254 231 255
rect 229 254 230 255
rect 228 254 229 255
rect 166 254 167 255
rect 165 254 166 255
rect 164 254 165 255
rect 163 254 164 255
rect 162 254 163 255
rect 161 254 162 255
rect 160 254 161 255
rect 159 254 160 255
rect 158 254 159 255
rect 157 254 158 255
rect 156 254 157 255
rect 155 254 156 255
rect 154 254 155 255
rect 153 254 154 255
rect 152 254 153 255
rect 151 254 152 255
rect 150 254 151 255
rect 149 254 150 255
rect 148 254 149 255
rect 147 254 148 255
rect 146 254 147 255
rect 145 254 146 255
rect 144 254 145 255
rect 143 254 144 255
rect 142 254 143 255
rect 141 254 142 255
rect 140 254 141 255
rect 139 254 140 255
rect 138 254 139 255
rect 137 254 138 255
rect 136 254 137 255
rect 135 254 136 255
rect 134 254 135 255
rect 133 254 134 255
rect 132 254 133 255
rect 131 254 132 255
rect 130 254 131 255
rect 129 254 130 255
rect 128 254 129 255
rect 127 254 128 255
rect 126 254 127 255
rect 125 254 126 255
rect 124 254 125 255
rect 123 254 124 255
rect 122 254 123 255
rect 121 254 122 255
rect 120 254 121 255
rect 107 254 108 255
rect 106 254 107 255
rect 105 254 106 255
rect 104 254 105 255
rect 103 254 104 255
rect 102 254 103 255
rect 101 254 102 255
rect 100 254 101 255
rect 99 254 100 255
rect 98 254 99 255
rect 97 254 98 255
rect 96 254 97 255
rect 95 254 96 255
rect 94 254 95 255
rect 93 254 94 255
rect 92 254 93 255
rect 91 254 92 255
rect 90 254 91 255
rect 89 254 90 255
rect 88 254 89 255
rect 87 254 88 255
rect 86 254 87 255
rect 85 254 86 255
rect 84 254 85 255
rect 83 254 84 255
rect 82 254 83 255
rect 81 254 82 255
rect 80 254 81 255
rect 79 254 80 255
rect 78 254 79 255
rect 77 254 78 255
rect 76 254 77 255
rect 75 254 76 255
rect 74 254 75 255
rect 73 254 74 255
rect 72 254 73 255
rect 71 254 72 255
rect 70 254 71 255
rect 69 254 70 255
rect 68 254 69 255
rect 67 254 68 255
rect 66 254 67 255
rect 65 254 66 255
rect 64 254 65 255
rect 63 254 64 255
rect 52 254 53 255
rect 51 254 52 255
rect 50 254 51 255
rect 49 254 50 255
rect 48 254 49 255
rect 47 254 48 255
rect 46 254 47 255
rect 45 254 46 255
rect 44 254 45 255
rect 43 254 44 255
rect 42 254 43 255
rect 41 254 42 255
rect 40 254 41 255
rect 39 254 40 255
rect 38 254 39 255
rect 37 254 38 255
rect 36 254 37 255
rect 35 254 36 255
rect 34 254 35 255
rect 33 254 34 255
rect 32 254 33 255
rect 31 254 32 255
rect 20 254 21 255
rect 19 254 20 255
rect 18 254 19 255
rect 17 254 18 255
rect 16 254 17 255
rect 15 254 16 255
rect 14 254 15 255
rect 13 254 14 255
rect 12 254 13 255
rect 11 254 12 255
rect 10 254 11 255
rect 9 254 10 255
rect 8 254 9 255
rect 7 254 8 255
rect 6 254 7 255
rect 5 254 6 255
rect 4 254 5 255
rect 3 254 4 255
rect 2 254 3 255
rect 1 254 2 255
rect 475 255 476 256
rect 474 255 475 256
rect 473 255 474 256
rect 472 255 473 256
rect 471 255 472 256
rect 470 255 471 256
rect 305 255 306 256
rect 304 255 305 256
rect 303 255 304 256
rect 302 255 303 256
rect 301 255 302 256
rect 300 255 301 256
rect 299 255 300 256
rect 298 255 299 256
rect 297 255 298 256
rect 296 255 297 256
rect 295 255 296 256
rect 294 255 295 256
rect 293 255 294 256
rect 292 255 293 256
rect 291 255 292 256
rect 290 255 291 256
rect 289 255 290 256
rect 288 255 289 256
rect 287 255 288 256
rect 286 255 287 256
rect 285 255 286 256
rect 284 255 285 256
rect 283 255 284 256
rect 282 255 283 256
rect 281 255 282 256
rect 280 255 281 256
rect 279 255 280 256
rect 278 255 279 256
rect 277 255 278 256
rect 276 255 277 256
rect 275 255 276 256
rect 274 255 275 256
rect 273 255 274 256
rect 272 255 273 256
rect 271 255 272 256
rect 270 255 271 256
rect 269 255 270 256
rect 268 255 269 256
rect 267 255 268 256
rect 266 255 267 256
rect 265 255 266 256
rect 264 255 265 256
rect 263 255 264 256
rect 262 255 263 256
rect 261 255 262 256
rect 260 255 261 256
rect 259 255 260 256
rect 258 255 259 256
rect 257 255 258 256
rect 256 255 257 256
rect 255 255 256 256
rect 254 255 255 256
rect 253 255 254 256
rect 252 255 253 256
rect 251 255 252 256
rect 250 255 251 256
rect 249 255 250 256
rect 248 255 249 256
rect 247 255 248 256
rect 246 255 247 256
rect 245 255 246 256
rect 244 255 245 256
rect 243 255 244 256
rect 242 255 243 256
rect 241 255 242 256
rect 240 255 241 256
rect 239 255 240 256
rect 238 255 239 256
rect 237 255 238 256
rect 236 255 237 256
rect 235 255 236 256
rect 234 255 235 256
rect 233 255 234 256
rect 232 255 233 256
rect 231 255 232 256
rect 230 255 231 256
rect 229 255 230 256
rect 228 255 229 256
rect 227 255 228 256
rect 168 255 169 256
rect 167 255 168 256
rect 166 255 167 256
rect 165 255 166 256
rect 164 255 165 256
rect 163 255 164 256
rect 162 255 163 256
rect 161 255 162 256
rect 160 255 161 256
rect 159 255 160 256
rect 158 255 159 256
rect 157 255 158 256
rect 156 255 157 256
rect 155 255 156 256
rect 154 255 155 256
rect 153 255 154 256
rect 152 255 153 256
rect 151 255 152 256
rect 150 255 151 256
rect 149 255 150 256
rect 148 255 149 256
rect 147 255 148 256
rect 146 255 147 256
rect 145 255 146 256
rect 144 255 145 256
rect 143 255 144 256
rect 142 255 143 256
rect 141 255 142 256
rect 140 255 141 256
rect 139 255 140 256
rect 138 255 139 256
rect 137 255 138 256
rect 136 255 137 256
rect 135 255 136 256
rect 134 255 135 256
rect 133 255 134 256
rect 132 255 133 256
rect 131 255 132 256
rect 130 255 131 256
rect 129 255 130 256
rect 128 255 129 256
rect 127 255 128 256
rect 126 255 127 256
rect 125 255 126 256
rect 124 255 125 256
rect 123 255 124 256
rect 122 255 123 256
rect 121 255 122 256
rect 120 255 121 256
rect 107 255 108 256
rect 106 255 107 256
rect 105 255 106 256
rect 104 255 105 256
rect 103 255 104 256
rect 102 255 103 256
rect 101 255 102 256
rect 100 255 101 256
rect 99 255 100 256
rect 98 255 99 256
rect 97 255 98 256
rect 96 255 97 256
rect 95 255 96 256
rect 94 255 95 256
rect 93 255 94 256
rect 92 255 93 256
rect 91 255 92 256
rect 90 255 91 256
rect 89 255 90 256
rect 88 255 89 256
rect 87 255 88 256
rect 86 255 87 256
rect 85 255 86 256
rect 84 255 85 256
rect 83 255 84 256
rect 82 255 83 256
rect 81 255 82 256
rect 80 255 81 256
rect 79 255 80 256
rect 78 255 79 256
rect 77 255 78 256
rect 76 255 77 256
rect 75 255 76 256
rect 74 255 75 256
rect 73 255 74 256
rect 72 255 73 256
rect 71 255 72 256
rect 70 255 71 256
rect 69 255 70 256
rect 68 255 69 256
rect 67 255 68 256
rect 66 255 67 256
rect 65 255 66 256
rect 53 255 54 256
rect 52 255 53 256
rect 51 255 52 256
rect 50 255 51 256
rect 49 255 50 256
rect 48 255 49 256
rect 47 255 48 256
rect 46 255 47 256
rect 45 255 46 256
rect 44 255 45 256
rect 43 255 44 256
rect 42 255 43 256
rect 41 255 42 256
rect 40 255 41 256
rect 39 255 40 256
rect 38 255 39 256
rect 37 255 38 256
rect 36 255 37 256
rect 35 255 36 256
rect 34 255 35 256
rect 33 255 34 256
rect 32 255 33 256
rect 31 255 32 256
rect 20 255 21 256
rect 19 255 20 256
rect 18 255 19 256
rect 17 255 18 256
rect 16 255 17 256
rect 15 255 16 256
rect 14 255 15 256
rect 13 255 14 256
rect 12 255 13 256
rect 11 255 12 256
rect 10 255 11 256
rect 9 255 10 256
rect 8 255 9 256
rect 7 255 8 256
rect 6 255 7 256
rect 5 255 6 256
rect 4 255 5 256
rect 3 255 4 256
rect 2 255 3 256
rect 1 255 2 256
rect 304 256 305 257
rect 303 256 304 257
rect 302 256 303 257
rect 301 256 302 257
rect 300 256 301 257
rect 299 256 300 257
rect 298 256 299 257
rect 297 256 298 257
rect 296 256 297 257
rect 295 256 296 257
rect 294 256 295 257
rect 293 256 294 257
rect 292 256 293 257
rect 291 256 292 257
rect 290 256 291 257
rect 289 256 290 257
rect 288 256 289 257
rect 287 256 288 257
rect 286 256 287 257
rect 285 256 286 257
rect 284 256 285 257
rect 283 256 284 257
rect 282 256 283 257
rect 281 256 282 257
rect 280 256 281 257
rect 279 256 280 257
rect 278 256 279 257
rect 277 256 278 257
rect 276 256 277 257
rect 275 256 276 257
rect 274 256 275 257
rect 273 256 274 257
rect 272 256 273 257
rect 271 256 272 257
rect 270 256 271 257
rect 269 256 270 257
rect 268 256 269 257
rect 267 256 268 257
rect 266 256 267 257
rect 265 256 266 257
rect 264 256 265 257
rect 263 256 264 257
rect 262 256 263 257
rect 261 256 262 257
rect 260 256 261 257
rect 259 256 260 257
rect 258 256 259 257
rect 257 256 258 257
rect 256 256 257 257
rect 255 256 256 257
rect 254 256 255 257
rect 253 256 254 257
rect 252 256 253 257
rect 251 256 252 257
rect 250 256 251 257
rect 249 256 250 257
rect 248 256 249 257
rect 247 256 248 257
rect 246 256 247 257
rect 245 256 246 257
rect 244 256 245 257
rect 243 256 244 257
rect 242 256 243 257
rect 241 256 242 257
rect 240 256 241 257
rect 239 256 240 257
rect 238 256 239 257
rect 237 256 238 257
rect 236 256 237 257
rect 235 256 236 257
rect 234 256 235 257
rect 233 256 234 257
rect 232 256 233 257
rect 231 256 232 257
rect 230 256 231 257
rect 229 256 230 257
rect 228 256 229 257
rect 227 256 228 257
rect 171 256 172 257
rect 170 256 171 257
rect 169 256 170 257
rect 168 256 169 257
rect 167 256 168 257
rect 166 256 167 257
rect 165 256 166 257
rect 164 256 165 257
rect 163 256 164 257
rect 162 256 163 257
rect 161 256 162 257
rect 160 256 161 257
rect 159 256 160 257
rect 158 256 159 257
rect 157 256 158 257
rect 156 256 157 257
rect 155 256 156 257
rect 154 256 155 257
rect 153 256 154 257
rect 152 256 153 257
rect 151 256 152 257
rect 150 256 151 257
rect 149 256 150 257
rect 148 256 149 257
rect 147 256 148 257
rect 146 256 147 257
rect 145 256 146 257
rect 144 256 145 257
rect 143 256 144 257
rect 142 256 143 257
rect 141 256 142 257
rect 140 256 141 257
rect 139 256 140 257
rect 138 256 139 257
rect 137 256 138 257
rect 136 256 137 257
rect 135 256 136 257
rect 134 256 135 257
rect 133 256 134 257
rect 132 256 133 257
rect 131 256 132 257
rect 130 256 131 257
rect 129 256 130 257
rect 128 256 129 257
rect 127 256 128 257
rect 126 256 127 257
rect 125 256 126 257
rect 124 256 125 257
rect 123 256 124 257
rect 122 256 123 257
rect 121 256 122 257
rect 120 256 121 257
rect 107 256 108 257
rect 106 256 107 257
rect 105 256 106 257
rect 104 256 105 257
rect 103 256 104 257
rect 102 256 103 257
rect 101 256 102 257
rect 100 256 101 257
rect 99 256 100 257
rect 98 256 99 257
rect 97 256 98 257
rect 96 256 97 257
rect 95 256 96 257
rect 94 256 95 257
rect 93 256 94 257
rect 92 256 93 257
rect 91 256 92 257
rect 90 256 91 257
rect 89 256 90 257
rect 88 256 89 257
rect 87 256 88 257
rect 86 256 87 257
rect 85 256 86 257
rect 84 256 85 257
rect 83 256 84 257
rect 82 256 83 257
rect 81 256 82 257
rect 80 256 81 257
rect 79 256 80 257
rect 78 256 79 257
rect 77 256 78 257
rect 76 256 77 257
rect 75 256 76 257
rect 74 256 75 257
rect 73 256 74 257
rect 72 256 73 257
rect 71 256 72 257
rect 70 256 71 257
rect 69 256 70 257
rect 68 256 69 257
rect 67 256 68 257
rect 66 256 67 257
rect 53 256 54 257
rect 52 256 53 257
rect 51 256 52 257
rect 50 256 51 257
rect 49 256 50 257
rect 48 256 49 257
rect 47 256 48 257
rect 46 256 47 257
rect 45 256 46 257
rect 44 256 45 257
rect 43 256 44 257
rect 42 256 43 257
rect 41 256 42 257
rect 40 256 41 257
rect 39 256 40 257
rect 38 256 39 257
rect 37 256 38 257
rect 36 256 37 257
rect 35 256 36 257
rect 34 256 35 257
rect 33 256 34 257
rect 32 256 33 257
rect 20 256 21 257
rect 19 256 20 257
rect 18 256 19 257
rect 17 256 18 257
rect 16 256 17 257
rect 15 256 16 257
rect 14 256 15 257
rect 13 256 14 257
rect 12 256 13 257
rect 11 256 12 257
rect 10 256 11 257
rect 9 256 10 257
rect 8 256 9 257
rect 7 256 8 257
rect 6 256 7 257
rect 5 256 6 257
rect 4 256 5 257
rect 3 256 4 257
rect 2 256 3 257
rect 1 256 2 257
rect 303 257 304 258
rect 302 257 303 258
rect 301 257 302 258
rect 300 257 301 258
rect 299 257 300 258
rect 298 257 299 258
rect 297 257 298 258
rect 296 257 297 258
rect 295 257 296 258
rect 294 257 295 258
rect 293 257 294 258
rect 292 257 293 258
rect 291 257 292 258
rect 290 257 291 258
rect 289 257 290 258
rect 288 257 289 258
rect 287 257 288 258
rect 286 257 287 258
rect 285 257 286 258
rect 284 257 285 258
rect 283 257 284 258
rect 282 257 283 258
rect 281 257 282 258
rect 280 257 281 258
rect 279 257 280 258
rect 278 257 279 258
rect 277 257 278 258
rect 276 257 277 258
rect 275 257 276 258
rect 274 257 275 258
rect 273 257 274 258
rect 272 257 273 258
rect 271 257 272 258
rect 270 257 271 258
rect 269 257 270 258
rect 268 257 269 258
rect 267 257 268 258
rect 266 257 267 258
rect 265 257 266 258
rect 264 257 265 258
rect 263 257 264 258
rect 262 257 263 258
rect 261 257 262 258
rect 260 257 261 258
rect 259 257 260 258
rect 258 257 259 258
rect 257 257 258 258
rect 256 257 257 258
rect 255 257 256 258
rect 254 257 255 258
rect 253 257 254 258
rect 252 257 253 258
rect 251 257 252 258
rect 250 257 251 258
rect 249 257 250 258
rect 248 257 249 258
rect 247 257 248 258
rect 246 257 247 258
rect 245 257 246 258
rect 244 257 245 258
rect 243 257 244 258
rect 242 257 243 258
rect 241 257 242 258
rect 240 257 241 258
rect 239 257 240 258
rect 238 257 239 258
rect 237 257 238 258
rect 236 257 237 258
rect 235 257 236 258
rect 234 257 235 258
rect 233 257 234 258
rect 232 257 233 258
rect 231 257 232 258
rect 230 257 231 258
rect 229 257 230 258
rect 228 257 229 258
rect 227 257 228 258
rect 175 257 176 258
rect 174 257 175 258
rect 173 257 174 258
rect 172 257 173 258
rect 171 257 172 258
rect 170 257 171 258
rect 169 257 170 258
rect 168 257 169 258
rect 167 257 168 258
rect 166 257 167 258
rect 165 257 166 258
rect 164 257 165 258
rect 163 257 164 258
rect 162 257 163 258
rect 161 257 162 258
rect 160 257 161 258
rect 159 257 160 258
rect 158 257 159 258
rect 157 257 158 258
rect 156 257 157 258
rect 155 257 156 258
rect 154 257 155 258
rect 153 257 154 258
rect 152 257 153 258
rect 151 257 152 258
rect 150 257 151 258
rect 149 257 150 258
rect 148 257 149 258
rect 147 257 148 258
rect 146 257 147 258
rect 145 257 146 258
rect 144 257 145 258
rect 143 257 144 258
rect 142 257 143 258
rect 141 257 142 258
rect 140 257 141 258
rect 139 257 140 258
rect 138 257 139 258
rect 137 257 138 258
rect 136 257 137 258
rect 135 257 136 258
rect 134 257 135 258
rect 133 257 134 258
rect 132 257 133 258
rect 131 257 132 258
rect 130 257 131 258
rect 129 257 130 258
rect 128 257 129 258
rect 127 257 128 258
rect 126 257 127 258
rect 125 257 126 258
rect 124 257 125 258
rect 123 257 124 258
rect 122 257 123 258
rect 121 257 122 258
rect 120 257 121 258
rect 108 257 109 258
rect 107 257 108 258
rect 106 257 107 258
rect 105 257 106 258
rect 104 257 105 258
rect 103 257 104 258
rect 102 257 103 258
rect 101 257 102 258
rect 100 257 101 258
rect 99 257 100 258
rect 98 257 99 258
rect 97 257 98 258
rect 96 257 97 258
rect 95 257 96 258
rect 94 257 95 258
rect 93 257 94 258
rect 92 257 93 258
rect 91 257 92 258
rect 90 257 91 258
rect 89 257 90 258
rect 88 257 89 258
rect 87 257 88 258
rect 86 257 87 258
rect 85 257 86 258
rect 84 257 85 258
rect 83 257 84 258
rect 82 257 83 258
rect 81 257 82 258
rect 80 257 81 258
rect 79 257 80 258
rect 78 257 79 258
rect 77 257 78 258
rect 76 257 77 258
rect 75 257 76 258
rect 74 257 75 258
rect 73 257 74 258
rect 72 257 73 258
rect 71 257 72 258
rect 70 257 71 258
rect 69 257 70 258
rect 68 257 69 258
rect 67 257 68 258
rect 53 257 54 258
rect 52 257 53 258
rect 51 257 52 258
rect 50 257 51 258
rect 49 257 50 258
rect 48 257 49 258
rect 47 257 48 258
rect 46 257 47 258
rect 45 257 46 258
rect 44 257 45 258
rect 43 257 44 258
rect 42 257 43 258
rect 41 257 42 258
rect 40 257 41 258
rect 39 257 40 258
rect 38 257 39 258
rect 37 257 38 258
rect 36 257 37 258
rect 35 257 36 258
rect 34 257 35 258
rect 33 257 34 258
rect 32 257 33 258
rect 21 257 22 258
rect 20 257 21 258
rect 19 257 20 258
rect 18 257 19 258
rect 17 257 18 258
rect 16 257 17 258
rect 15 257 16 258
rect 14 257 15 258
rect 13 257 14 258
rect 12 257 13 258
rect 11 257 12 258
rect 10 257 11 258
rect 9 257 10 258
rect 8 257 9 258
rect 7 257 8 258
rect 6 257 7 258
rect 5 257 6 258
rect 4 257 5 258
rect 3 257 4 258
rect 2 257 3 258
rect 1 257 2 258
rect 302 258 303 259
rect 301 258 302 259
rect 300 258 301 259
rect 299 258 300 259
rect 298 258 299 259
rect 297 258 298 259
rect 296 258 297 259
rect 295 258 296 259
rect 294 258 295 259
rect 293 258 294 259
rect 292 258 293 259
rect 291 258 292 259
rect 290 258 291 259
rect 289 258 290 259
rect 288 258 289 259
rect 287 258 288 259
rect 286 258 287 259
rect 285 258 286 259
rect 284 258 285 259
rect 283 258 284 259
rect 282 258 283 259
rect 281 258 282 259
rect 280 258 281 259
rect 279 258 280 259
rect 278 258 279 259
rect 277 258 278 259
rect 276 258 277 259
rect 275 258 276 259
rect 274 258 275 259
rect 273 258 274 259
rect 272 258 273 259
rect 271 258 272 259
rect 270 258 271 259
rect 269 258 270 259
rect 268 258 269 259
rect 267 258 268 259
rect 266 258 267 259
rect 265 258 266 259
rect 264 258 265 259
rect 263 258 264 259
rect 262 258 263 259
rect 261 258 262 259
rect 260 258 261 259
rect 259 258 260 259
rect 258 258 259 259
rect 257 258 258 259
rect 256 258 257 259
rect 255 258 256 259
rect 254 258 255 259
rect 253 258 254 259
rect 252 258 253 259
rect 251 258 252 259
rect 250 258 251 259
rect 249 258 250 259
rect 248 258 249 259
rect 247 258 248 259
rect 246 258 247 259
rect 245 258 246 259
rect 244 258 245 259
rect 243 258 244 259
rect 242 258 243 259
rect 241 258 242 259
rect 240 258 241 259
rect 239 258 240 259
rect 238 258 239 259
rect 237 258 238 259
rect 236 258 237 259
rect 235 258 236 259
rect 234 258 235 259
rect 233 258 234 259
rect 232 258 233 259
rect 231 258 232 259
rect 230 258 231 259
rect 229 258 230 259
rect 228 258 229 259
rect 227 258 228 259
rect 226 258 227 259
rect 179 258 180 259
rect 178 258 179 259
rect 177 258 178 259
rect 176 258 177 259
rect 175 258 176 259
rect 174 258 175 259
rect 173 258 174 259
rect 172 258 173 259
rect 171 258 172 259
rect 170 258 171 259
rect 169 258 170 259
rect 168 258 169 259
rect 167 258 168 259
rect 166 258 167 259
rect 165 258 166 259
rect 164 258 165 259
rect 163 258 164 259
rect 162 258 163 259
rect 161 258 162 259
rect 160 258 161 259
rect 159 258 160 259
rect 158 258 159 259
rect 157 258 158 259
rect 156 258 157 259
rect 155 258 156 259
rect 154 258 155 259
rect 153 258 154 259
rect 152 258 153 259
rect 151 258 152 259
rect 150 258 151 259
rect 149 258 150 259
rect 148 258 149 259
rect 147 258 148 259
rect 146 258 147 259
rect 145 258 146 259
rect 144 258 145 259
rect 143 258 144 259
rect 142 258 143 259
rect 141 258 142 259
rect 140 258 141 259
rect 139 258 140 259
rect 138 258 139 259
rect 137 258 138 259
rect 136 258 137 259
rect 135 258 136 259
rect 134 258 135 259
rect 133 258 134 259
rect 132 258 133 259
rect 131 258 132 259
rect 130 258 131 259
rect 129 258 130 259
rect 128 258 129 259
rect 127 258 128 259
rect 126 258 127 259
rect 125 258 126 259
rect 124 258 125 259
rect 123 258 124 259
rect 122 258 123 259
rect 121 258 122 259
rect 120 258 121 259
rect 108 258 109 259
rect 107 258 108 259
rect 106 258 107 259
rect 105 258 106 259
rect 104 258 105 259
rect 103 258 104 259
rect 102 258 103 259
rect 101 258 102 259
rect 100 258 101 259
rect 99 258 100 259
rect 98 258 99 259
rect 97 258 98 259
rect 96 258 97 259
rect 95 258 96 259
rect 94 258 95 259
rect 93 258 94 259
rect 92 258 93 259
rect 91 258 92 259
rect 90 258 91 259
rect 89 258 90 259
rect 88 258 89 259
rect 87 258 88 259
rect 86 258 87 259
rect 85 258 86 259
rect 84 258 85 259
rect 83 258 84 259
rect 82 258 83 259
rect 81 258 82 259
rect 80 258 81 259
rect 79 258 80 259
rect 78 258 79 259
rect 77 258 78 259
rect 76 258 77 259
rect 75 258 76 259
rect 74 258 75 259
rect 73 258 74 259
rect 72 258 73 259
rect 71 258 72 259
rect 70 258 71 259
rect 69 258 70 259
rect 68 258 69 259
rect 53 258 54 259
rect 52 258 53 259
rect 51 258 52 259
rect 50 258 51 259
rect 49 258 50 259
rect 48 258 49 259
rect 47 258 48 259
rect 46 258 47 259
rect 45 258 46 259
rect 44 258 45 259
rect 43 258 44 259
rect 42 258 43 259
rect 41 258 42 259
rect 40 258 41 259
rect 39 258 40 259
rect 38 258 39 259
rect 37 258 38 259
rect 36 258 37 259
rect 35 258 36 259
rect 34 258 35 259
rect 33 258 34 259
rect 32 258 33 259
rect 21 258 22 259
rect 20 258 21 259
rect 19 258 20 259
rect 18 258 19 259
rect 17 258 18 259
rect 16 258 17 259
rect 15 258 16 259
rect 14 258 15 259
rect 13 258 14 259
rect 12 258 13 259
rect 11 258 12 259
rect 10 258 11 259
rect 9 258 10 259
rect 8 258 9 259
rect 7 258 8 259
rect 6 258 7 259
rect 5 258 6 259
rect 4 258 5 259
rect 3 258 4 259
rect 2 258 3 259
rect 1 258 2 259
rect 301 259 302 260
rect 300 259 301 260
rect 299 259 300 260
rect 298 259 299 260
rect 297 259 298 260
rect 296 259 297 260
rect 295 259 296 260
rect 294 259 295 260
rect 293 259 294 260
rect 292 259 293 260
rect 291 259 292 260
rect 290 259 291 260
rect 289 259 290 260
rect 288 259 289 260
rect 287 259 288 260
rect 286 259 287 260
rect 285 259 286 260
rect 284 259 285 260
rect 283 259 284 260
rect 282 259 283 260
rect 281 259 282 260
rect 280 259 281 260
rect 279 259 280 260
rect 278 259 279 260
rect 277 259 278 260
rect 276 259 277 260
rect 275 259 276 260
rect 274 259 275 260
rect 273 259 274 260
rect 272 259 273 260
rect 271 259 272 260
rect 270 259 271 260
rect 269 259 270 260
rect 268 259 269 260
rect 267 259 268 260
rect 266 259 267 260
rect 265 259 266 260
rect 264 259 265 260
rect 263 259 264 260
rect 262 259 263 260
rect 261 259 262 260
rect 260 259 261 260
rect 259 259 260 260
rect 258 259 259 260
rect 257 259 258 260
rect 256 259 257 260
rect 255 259 256 260
rect 254 259 255 260
rect 253 259 254 260
rect 252 259 253 260
rect 251 259 252 260
rect 250 259 251 260
rect 249 259 250 260
rect 248 259 249 260
rect 247 259 248 260
rect 246 259 247 260
rect 245 259 246 260
rect 244 259 245 260
rect 243 259 244 260
rect 242 259 243 260
rect 241 259 242 260
rect 240 259 241 260
rect 239 259 240 260
rect 238 259 239 260
rect 237 259 238 260
rect 236 259 237 260
rect 235 259 236 260
rect 234 259 235 260
rect 233 259 234 260
rect 232 259 233 260
rect 231 259 232 260
rect 230 259 231 260
rect 229 259 230 260
rect 228 259 229 260
rect 227 259 228 260
rect 226 259 227 260
rect 183 259 184 260
rect 182 259 183 260
rect 181 259 182 260
rect 180 259 181 260
rect 179 259 180 260
rect 178 259 179 260
rect 177 259 178 260
rect 176 259 177 260
rect 175 259 176 260
rect 174 259 175 260
rect 173 259 174 260
rect 172 259 173 260
rect 171 259 172 260
rect 170 259 171 260
rect 169 259 170 260
rect 168 259 169 260
rect 167 259 168 260
rect 166 259 167 260
rect 165 259 166 260
rect 164 259 165 260
rect 163 259 164 260
rect 162 259 163 260
rect 161 259 162 260
rect 160 259 161 260
rect 159 259 160 260
rect 158 259 159 260
rect 157 259 158 260
rect 156 259 157 260
rect 155 259 156 260
rect 154 259 155 260
rect 153 259 154 260
rect 152 259 153 260
rect 151 259 152 260
rect 150 259 151 260
rect 149 259 150 260
rect 148 259 149 260
rect 147 259 148 260
rect 146 259 147 260
rect 145 259 146 260
rect 144 259 145 260
rect 143 259 144 260
rect 142 259 143 260
rect 141 259 142 260
rect 140 259 141 260
rect 139 259 140 260
rect 138 259 139 260
rect 137 259 138 260
rect 136 259 137 260
rect 135 259 136 260
rect 134 259 135 260
rect 133 259 134 260
rect 132 259 133 260
rect 131 259 132 260
rect 130 259 131 260
rect 129 259 130 260
rect 128 259 129 260
rect 127 259 128 260
rect 126 259 127 260
rect 125 259 126 260
rect 124 259 125 260
rect 123 259 124 260
rect 122 259 123 260
rect 121 259 122 260
rect 108 259 109 260
rect 107 259 108 260
rect 106 259 107 260
rect 105 259 106 260
rect 104 259 105 260
rect 103 259 104 260
rect 102 259 103 260
rect 101 259 102 260
rect 100 259 101 260
rect 99 259 100 260
rect 98 259 99 260
rect 97 259 98 260
rect 96 259 97 260
rect 95 259 96 260
rect 94 259 95 260
rect 93 259 94 260
rect 92 259 93 260
rect 91 259 92 260
rect 90 259 91 260
rect 89 259 90 260
rect 88 259 89 260
rect 87 259 88 260
rect 86 259 87 260
rect 85 259 86 260
rect 84 259 85 260
rect 83 259 84 260
rect 82 259 83 260
rect 81 259 82 260
rect 80 259 81 260
rect 79 259 80 260
rect 78 259 79 260
rect 77 259 78 260
rect 76 259 77 260
rect 75 259 76 260
rect 74 259 75 260
rect 73 259 74 260
rect 72 259 73 260
rect 71 259 72 260
rect 70 259 71 260
rect 69 259 70 260
rect 54 259 55 260
rect 53 259 54 260
rect 52 259 53 260
rect 51 259 52 260
rect 50 259 51 260
rect 49 259 50 260
rect 48 259 49 260
rect 47 259 48 260
rect 46 259 47 260
rect 45 259 46 260
rect 44 259 45 260
rect 43 259 44 260
rect 42 259 43 260
rect 41 259 42 260
rect 40 259 41 260
rect 39 259 40 260
rect 38 259 39 260
rect 37 259 38 260
rect 36 259 37 260
rect 35 259 36 260
rect 34 259 35 260
rect 33 259 34 260
rect 21 259 22 260
rect 20 259 21 260
rect 19 259 20 260
rect 18 259 19 260
rect 17 259 18 260
rect 16 259 17 260
rect 15 259 16 260
rect 14 259 15 260
rect 13 259 14 260
rect 12 259 13 260
rect 11 259 12 260
rect 10 259 11 260
rect 9 259 10 260
rect 8 259 9 260
rect 7 259 8 260
rect 6 259 7 260
rect 5 259 6 260
rect 4 259 5 260
rect 3 259 4 260
rect 2 259 3 260
rect 1 259 2 260
rect 300 260 301 261
rect 299 260 300 261
rect 298 260 299 261
rect 297 260 298 261
rect 296 260 297 261
rect 295 260 296 261
rect 294 260 295 261
rect 293 260 294 261
rect 292 260 293 261
rect 291 260 292 261
rect 290 260 291 261
rect 289 260 290 261
rect 288 260 289 261
rect 287 260 288 261
rect 286 260 287 261
rect 285 260 286 261
rect 284 260 285 261
rect 283 260 284 261
rect 282 260 283 261
rect 281 260 282 261
rect 280 260 281 261
rect 279 260 280 261
rect 278 260 279 261
rect 277 260 278 261
rect 276 260 277 261
rect 275 260 276 261
rect 274 260 275 261
rect 273 260 274 261
rect 272 260 273 261
rect 271 260 272 261
rect 270 260 271 261
rect 269 260 270 261
rect 268 260 269 261
rect 267 260 268 261
rect 266 260 267 261
rect 265 260 266 261
rect 264 260 265 261
rect 263 260 264 261
rect 262 260 263 261
rect 261 260 262 261
rect 260 260 261 261
rect 259 260 260 261
rect 258 260 259 261
rect 257 260 258 261
rect 256 260 257 261
rect 255 260 256 261
rect 254 260 255 261
rect 253 260 254 261
rect 252 260 253 261
rect 251 260 252 261
rect 250 260 251 261
rect 249 260 250 261
rect 248 260 249 261
rect 247 260 248 261
rect 246 260 247 261
rect 245 260 246 261
rect 244 260 245 261
rect 243 260 244 261
rect 242 260 243 261
rect 241 260 242 261
rect 240 260 241 261
rect 239 260 240 261
rect 238 260 239 261
rect 237 260 238 261
rect 236 260 237 261
rect 235 260 236 261
rect 234 260 235 261
rect 233 260 234 261
rect 232 260 233 261
rect 231 260 232 261
rect 230 260 231 261
rect 229 260 230 261
rect 228 260 229 261
rect 227 260 228 261
rect 226 260 227 261
rect 205 260 206 261
rect 204 260 205 261
rect 203 260 204 261
rect 202 260 203 261
rect 201 260 202 261
rect 200 260 201 261
rect 190 260 191 261
rect 189 260 190 261
rect 188 260 189 261
rect 187 260 188 261
rect 186 260 187 261
rect 185 260 186 261
rect 184 260 185 261
rect 183 260 184 261
rect 182 260 183 261
rect 181 260 182 261
rect 180 260 181 261
rect 179 260 180 261
rect 178 260 179 261
rect 177 260 178 261
rect 176 260 177 261
rect 175 260 176 261
rect 174 260 175 261
rect 173 260 174 261
rect 172 260 173 261
rect 171 260 172 261
rect 170 260 171 261
rect 169 260 170 261
rect 168 260 169 261
rect 167 260 168 261
rect 166 260 167 261
rect 165 260 166 261
rect 164 260 165 261
rect 163 260 164 261
rect 162 260 163 261
rect 161 260 162 261
rect 160 260 161 261
rect 159 260 160 261
rect 158 260 159 261
rect 157 260 158 261
rect 156 260 157 261
rect 155 260 156 261
rect 154 260 155 261
rect 153 260 154 261
rect 152 260 153 261
rect 151 260 152 261
rect 150 260 151 261
rect 149 260 150 261
rect 148 260 149 261
rect 147 260 148 261
rect 146 260 147 261
rect 145 260 146 261
rect 144 260 145 261
rect 143 260 144 261
rect 142 260 143 261
rect 141 260 142 261
rect 140 260 141 261
rect 139 260 140 261
rect 138 260 139 261
rect 137 260 138 261
rect 136 260 137 261
rect 135 260 136 261
rect 134 260 135 261
rect 133 260 134 261
rect 132 260 133 261
rect 131 260 132 261
rect 130 260 131 261
rect 129 260 130 261
rect 128 260 129 261
rect 127 260 128 261
rect 126 260 127 261
rect 125 260 126 261
rect 124 260 125 261
rect 123 260 124 261
rect 122 260 123 261
rect 121 260 122 261
rect 108 260 109 261
rect 107 260 108 261
rect 106 260 107 261
rect 105 260 106 261
rect 104 260 105 261
rect 103 260 104 261
rect 102 260 103 261
rect 101 260 102 261
rect 100 260 101 261
rect 99 260 100 261
rect 98 260 99 261
rect 97 260 98 261
rect 96 260 97 261
rect 95 260 96 261
rect 94 260 95 261
rect 93 260 94 261
rect 92 260 93 261
rect 91 260 92 261
rect 90 260 91 261
rect 89 260 90 261
rect 88 260 89 261
rect 87 260 88 261
rect 86 260 87 261
rect 85 260 86 261
rect 84 260 85 261
rect 83 260 84 261
rect 82 260 83 261
rect 81 260 82 261
rect 80 260 81 261
rect 79 260 80 261
rect 78 260 79 261
rect 77 260 78 261
rect 76 260 77 261
rect 75 260 76 261
rect 74 260 75 261
rect 73 260 74 261
rect 72 260 73 261
rect 71 260 72 261
rect 70 260 71 261
rect 54 260 55 261
rect 53 260 54 261
rect 52 260 53 261
rect 51 260 52 261
rect 50 260 51 261
rect 49 260 50 261
rect 48 260 49 261
rect 47 260 48 261
rect 46 260 47 261
rect 45 260 46 261
rect 44 260 45 261
rect 43 260 44 261
rect 42 260 43 261
rect 41 260 42 261
rect 40 260 41 261
rect 39 260 40 261
rect 38 260 39 261
rect 37 260 38 261
rect 36 260 37 261
rect 35 260 36 261
rect 34 260 35 261
rect 33 260 34 261
rect 22 260 23 261
rect 21 260 22 261
rect 20 260 21 261
rect 19 260 20 261
rect 18 260 19 261
rect 17 260 18 261
rect 16 260 17 261
rect 15 260 16 261
rect 14 260 15 261
rect 13 260 14 261
rect 12 260 13 261
rect 11 260 12 261
rect 10 260 11 261
rect 9 260 10 261
rect 8 260 9 261
rect 7 260 8 261
rect 6 260 7 261
rect 5 260 6 261
rect 4 260 5 261
rect 3 260 4 261
rect 2 260 3 261
rect 1 260 2 261
rect 300 261 301 262
rect 299 261 300 262
rect 298 261 299 262
rect 297 261 298 262
rect 296 261 297 262
rect 295 261 296 262
rect 294 261 295 262
rect 293 261 294 262
rect 292 261 293 262
rect 291 261 292 262
rect 290 261 291 262
rect 289 261 290 262
rect 288 261 289 262
rect 287 261 288 262
rect 286 261 287 262
rect 285 261 286 262
rect 284 261 285 262
rect 283 261 284 262
rect 282 261 283 262
rect 281 261 282 262
rect 280 261 281 262
rect 279 261 280 262
rect 278 261 279 262
rect 277 261 278 262
rect 276 261 277 262
rect 275 261 276 262
rect 274 261 275 262
rect 273 261 274 262
rect 272 261 273 262
rect 271 261 272 262
rect 270 261 271 262
rect 269 261 270 262
rect 268 261 269 262
rect 267 261 268 262
rect 266 261 267 262
rect 265 261 266 262
rect 264 261 265 262
rect 263 261 264 262
rect 262 261 263 262
rect 261 261 262 262
rect 260 261 261 262
rect 259 261 260 262
rect 258 261 259 262
rect 257 261 258 262
rect 256 261 257 262
rect 255 261 256 262
rect 254 261 255 262
rect 253 261 254 262
rect 252 261 253 262
rect 251 261 252 262
rect 250 261 251 262
rect 249 261 250 262
rect 248 261 249 262
rect 247 261 248 262
rect 246 261 247 262
rect 245 261 246 262
rect 244 261 245 262
rect 243 261 244 262
rect 242 261 243 262
rect 241 261 242 262
rect 240 261 241 262
rect 239 261 240 262
rect 238 261 239 262
rect 237 261 238 262
rect 236 261 237 262
rect 235 261 236 262
rect 234 261 235 262
rect 233 261 234 262
rect 232 261 233 262
rect 231 261 232 262
rect 230 261 231 262
rect 229 261 230 262
rect 228 261 229 262
rect 227 261 228 262
rect 226 261 227 262
rect 225 261 226 262
rect 204 261 205 262
rect 203 261 204 262
rect 202 261 203 262
rect 201 261 202 262
rect 200 261 201 262
rect 199 261 200 262
rect 198 261 199 262
rect 197 261 198 262
rect 196 261 197 262
rect 195 261 196 262
rect 194 261 195 262
rect 193 261 194 262
rect 192 261 193 262
rect 191 261 192 262
rect 190 261 191 262
rect 189 261 190 262
rect 188 261 189 262
rect 187 261 188 262
rect 186 261 187 262
rect 185 261 186 262
rect 184 261 185 262
rect 183 261 184 262
rect 182 261 183 262
rect 181 261 182 262
rect 180 261 181 262
rect 179 261 180 262
rect 178 261 179 262
rect 177 261 178 262
rect 176 261 177 262
rect 175 261 176 262
rect 174 261 175 262
rect 173 261 174 262
rect 172 261 173 262
rect 171 261 172 262
rect 170 261 171 262
rect 169 261 170 262
rect 168 261 169 262
rect 167 261 168 262
rect 166 261 167 262
rect 165 261 166 262
rect 164 261 165 262
rect 163 261 164 262
rect 162 261 163 262
rect 161 261 162 262
rect 160 261 161 262
rect 159 261 160 262
rect 158 261 159 262
rect 157 261 158 262
rect 156 261 157 262
rect 155 261 156 262
rect 154 261 155 262
rect 153 261 154 262
rect 152 261 153 262
rect 151 261 152 262
rect 150 261 151 262
rect 149 261 150 262
rect 148 261 149 262
rect 147 261 148 262
rect 146 261 147 262
rect 145 261 146 262
rect 144 261 145 262
rect 143 261 144 262
rect 142 261 143 262
rect 141 261 142 262
rect 140 261 141 262
rect 139 261 140 262
rect 138 261 139 262
rect 137 261 138 262
rect 136 261 137 262
rect 135 261 136 262
rect 134 261 135 262
rect 133 261 134 262
rect 132 261 133 262
rect 131 261 132 262
rect 130 261 131 262
rect 129 261 130 262
rect 128 261 129 262
rect 127 261 128 262
rect 126 261 127 262
rect 125 261 126 262
rect 124 261 125 262
rect 123 261 124 262
rect 122 261 123 262
rect 121 261 122 262
rect 108 261 109 262
rect 107 261 108 262
rect 106 261 107 262
rect 105 261 106 262
rect 104 261 105 262
rect 103 261 104 262
rect 102 261 103 262
rect 101 261 102 262
rect 100 261 101 262
rect 99 261 100 262
rect 98 261 99 262
rect 97 261 98 262
rect 96 261 97 262
rect 95 261 96 262
rect 94 261 95 262
rect 93 261 94 262
rect 92 261 93 262
rect 91 261 92 262
rect 90 261 91 262
rect 89 261 90 262
rect 88 261 89 262
rect 87 261 88 262
rect 86 261 87 262
rect 85 261 86 262
rect 84 261 85 262
rect 83 261 84 262
rect 82 261 83 262
rect 81 261 82 262
rect 80 261 81 262
rect 79 261 80 262
rect 78 261 79 262
rect 77 261 78 262
rect 76 261 77 262
rect 75 261 76 262
rect 74 261 75 262
rect 73 261 74 262
rect 72 261 73 262
rect 71 261 72 262
rect 70 261 71 262
rect 55 261 56 262
rect 54 261 55 262
rect 53 261 54 262
rect 52 261 53 262
rect 51 261 52 262
rect 50 261 51 262
rect 49 261 50 262
rect 48 261 49 262
rect 47 261 48 262
rect 46 261 47 262
rect 45 261 46 262
rect 44 261 45 262
rect 43 261 44 262
rect 42 261 43 262
rect 41 261 42 262
rect 40 261 41 262
rect 39 261 40 262
rect 38 261 39 262
rect 37 261 38 262
rect 36 261 37 262
rect 35 261 36 262
rect 34 261 35 262
rect 33 261 34 262
rect 22 261 23 262
rect 21 261 22 262
rect 20 261 21 262
rect 19 261 20 262
rect 18 261 19 262
rect 17 261 18 262
rect 16 261 17 262
rect 15 261 16 262
rect 14 261 15 262
rect 13 261 14 262
rect 12 261 13 262
rect 11 261 12 262
rect 10 261 11 262
rect 9 261 10 262
rect 8 261 9 262
rect 7 261 8 262
rect 6 261 7 262
rect 5 261 6 262
rect 4 261 5 262
rect 3 261 4 262
rect 2 261 3 262
rect 1 261 2 262
rect 299 262 300 263
rect 298 262 299 263
rect 297 262 298 263
rect 296 262 297 263
rect 295 262 296 263
rect 294 262 295 263
rect 293 262 294 263
rect 292 262 293 263
rect 291 262 292 263
rect 290 262 291 263
rect 289 262 290 263
rect 288 262 289 263
rect 287 262 288 263
rect 286 262 287 263
rect 285 262 286 263
rect 284 262 285 263
rect 283 262 284 263
rect 282 262 283 263
rect 281 262 282 263
rect 280 262 281 263
rect 279 262 280 263
rect 278 262 279 263
rect 277 262 278 263
rect 276 262 277 263
rect 275 262 276 263
rect 274 262 275 263
rect 273 262 274 263
rect 272 262 273 263
rect 271 262 272 263
rect 270 262 271 263
rect 269 262 270 263
rect 268 262 269 263
rect 267 262 268 263
rect 266 262 267 263
rect 265 262 266 263
rect 264 262 265 263
rect 263 262 264 263
rect 262 262 263 263
rect 261 262 262 263
rect 260 262 261 263
rect 259 262 260 263
rect 258 262 259 263
rect 257 262 258 263
rect 256 262 257 263
rect 255 262 256 263
rect 254 262 255 263
rect 253 262 254 263
rect 252 262 253 263
rect 251 262 252 263
rect 250 262 251 263
rect 249 262 250 263
rect 248 262 249 263
rect 247 262 248 263
rect 246 262 247 263
rect 245 262 246 263
rect 244 262 245 263
rect 243 262 244 263
rect 242 262 243 263
rect 241 262 242 263
rect 240 262 241 263
rect 239 262 240 263
rect 238 262 239 263
rect 237 262 238 263
rect 236 262 237 263
rect 235 262 236 263
rect 234 262 235 263
rect 233 262 234 263
rect 232 262 233 263
rect 231 262 232 263
rect 230 262 231 263
rect 229 262 230 263
rect 228 262 229 263
rect 227 262 228 263
rect 226 262 227 263
rect 225 262 226 263
rect 204 262 205 263
rect 203 262 204 263
rect 202 262 203 263
rect 201 262 202 263
rect 200 262 201 263
rect 199 262 200 263
rect 198 262 199 263
rect 197 262 198 263
rect 196 262 197 263
rect 195 262 196 263
rect 194 262 195 263
rect 193 262 194 263
rect 192 262 193 263
rect 191 262 192 263
rect 190 262 191 263
rect 189 262 190 263
rect 188 262 189 263
rect 187 262 188 263
rect 186 262 187 263
rect 185 262 186 263
rect 184 262 185 263
rect 183 262 184 263
rect 182 262 183 263
rect 181 262 182 263
rect 180 262 181 263
rect 179 262 180 263
rect 178 262 179 263
rect 177 262 178 263
rect 176 262 177 263
rect 175 262 176 263
rect 174 262 175 263
rect 173 262 174 263
rect 172 262 173 263
rect 171 262 172 263
rect 170 262 171 263
rect 169 262 170 263
rect 168 262 169 263
rect 167 262 168 263
rect 166 262 167 263
rect 165 262 166 263
rect 164 262 165 263
rect 163 262 164 263
rect 162 262 163 263
rect 161 262 162 263
rect 160 262 161 263
rect 159 262 160 263
rect 158 262 159 263
rect 157 262 158 263
rect 156 262 157 263
rect 155 262 156 263
rect 154 262 155 263
rect 153 262 154 263
rect 152 262 153 263
rect 151 262 152 263
rect 150 262 151 263
rect 149 262 150 263
rect 148 262 149 263
rect 147 262 148 263
rect 146 262 147 263
rect 145 262 146 263
rect 144 262 145 263
rect 143 262 144 263
rect 142 262 143 263
rect 141 262 142 263
rect 140 262 141 263
rect 139 262 140 263
rect 138 262 139 263
rect 137 262 138 263
rect 136 262 137 263
rect 135 262 136 263
rect 134 262 135 263
rect 133 262 134 263
rect 132 262 133 263
rect 131 262 132 263
rect 130 262 131 263
rect 129 262 130 263
rect 128 262 129 263
rect 127 262 128 263
rect 126 262 127 263
rect 125 262 126 263
rect 124 262 125 263
rect 123 262 124 263
rect 122 262 123 263
rect 121 262 122 263
rect 108 262 109 263
rect 107 262 108 263
rect 106 262 107 263
rect 105 262 106 263
rect 104 262 105 263
rect 103 262 104 263
rect 102 262 103 263
rect 101 262 102 263
rect 100 262 101 263
rect 99 262 100 263
rect 98 262 99 263
rect 97 262 98 263
rect 96 262 97 263
rect 95 262 96 263
rect 94 262 95 263
rect 93 262 94 263
rect 92 262 93 263
rect 91 262 92 263
rect 90 262 91 263
rect 89 262 90 263
rect 88 262 89 263
rect 87 262 88 263
rect 86 262 87 263
rect 85 262 86 263
rect 84 262 85 263
rect 83 262 84 263
rect 82 262 83 263
rect 81 262 82 263
rect 80 262 81 263
rect 79 262 80 263
rect 78 262 79 263
rect 77 262 78 263
rect 76 262 77 263
rect 75 262 76 263
rect 74 262 75 263
rect 73 262 74 263
rect 72 262 73 263
rect 71 262 72 263
rect 55 262 56 263
rect 54 262 55 263
rect 53 262 54 263
rect 52 262 53 263
rect 51 262 52 263
rect 50 262 51 263
rect 49 262 50 263
rect 48 262 49 263
rect 47 262 48 263
rect 46 262 47 263
rect 45 262 46 263
rect 44 262 45 263
rect 43 262 44 263
rect 42 262 43 263
rect 41 262 42 263
rect 40 262 41 263
rect 39 262 40 263
rect 38 262 39 263
rect 37 262 38 263
rect 36 262 37 263
rect 35 262 36 263
rect 34 262 35 263
rect 33 262 34 263
rect 22 262 23 263
rect 21 262 22 263
rect 20 262 21 263
rect 19 262 20 263
rect 18 262 19 263
rect 17 262 18 263
rect 16 262 17 263
rect 15 262 16 263
rect 14 262 15 263
rect 13 262 14 263
rect 12 262 13 263
rect 11 262 12 263
rect 10 262 11 263
rect 9 262 10 263
rect 8 262 9 263
rect 7 262 8 263
rect 6 262 7 263
rect 5 262 6 263
rect 4 262 5 263
rect 3 262 4 263
rect 2 262 3 263
rect 1 262 2 263
rect 298 263 299 264
rect 297 263 298 264
rect 296 263 297 264
rect 295 263 296 264
rect 294 263 295 264
rect 293 263 294 264
rect 292 263 293 264
rect 291 263 292 264
rect 290 263 291 264
rect 289 263 290 264
rect 288 263 289 264
rect 287 263 288 264
rect 286 263 287 264
rect 285 263 286 264
rect 284 263 285 264
rect 283 263 284 264
rect 282 263 283 264
rect 281 263 282 264
rect 280 263 281 264
rect 279 263 280 264
rect 278 263 279 264
rect 277 263 278 264
rect 276 263 277 264
rect 275 263 276 264
rect 274 263 275 264
rect 273 263 274 264
rect 272 263 273 264
rect 271 263 272 264
rect 270 263 271 264
rect 269 263 270 264
rect 268 263 269 264
rect 267 263 268 264
rect 266 263 267 264
rect 265 263 266 264
rect 264 263 265 264
rect 263 263 264 264
rect 262 263 263 264
rect 261 263 262 264
rect 260 263 261 264
rect 259 263 260 264
rect 258 263 259 264
rect 257 263 258 264
rect 256 263 257 264
rect 255 263 256 264
rect 254 263 255 264
rect 253 263 254 264
rect 252 263 253 264
rect 251 263 252 264
rect 250 263 251 264
rect 249 263 250 264
rect 248 263 249 264
rect 247 263 248 264
rect 246 263 247 264
rect 245 263 246 264
rect 244 263 245 264
rect 243 263 244 264
rect 242 263 243 264
rect 241 263 242 264
rect 240 263 241 264
rect 239 263 240 264
rect 238 263 239 264
rect 237 263 238 264
rect 236 263 237 264
rect 235 263 236 264
rect 234 263 235 264
rect 233 263 234 264
rect 232 263 233 264
rect 231 263 232 264
rect 230 263 231 264
rect 229 263 230 264
rect 228 263 229 264
rect 227 263 228 264
rect 226 263 227 264
rect 225 263 226 264
rect 204 263 205 264
rect 203 263 204 264
rect 202 263 203 264
rect 201 263 202 264
rect 200 263 201 264
rect 199 263 200 264
rect 198 263 199 264
rect 197 263 198 264
rect 196 263 197 264
rect 195 263 196 264
rect 194 263 195 264
rect 193 263 194 264
rect 192 263 193 264
rect 191 263 192 264
rect 190 263 191 264
rect 189 263 190 264
rect 188 263 189 264
rect 187 263 188 264
rect 186 263 187 264
rect 185 263 186 264
rect 184 263 185 264
rect 183 263 184 264
rect 182 263 183 264
rect 181 263 182 264
rect 180 263 181 264
rect 179 263 180 264
rect 178 263 179 264
rect 177 263 178 264
rect 176 263 177 264
rect 175 263 176 264
rect 174 263 175 264
rect 173 263 174 264
rect 172 263 173 264
rect 171 263 172 264
rect 170 263 171 264
rect 169 263 170 264
rect 168 263 169 264
rect 167 263 168 264
rect 166 263 167 264
rect 165 263 166 264
rect 164 263 165 264
rect 163 263 164 264
rect 162 263 163 264
rect 161 263 162 264
rect 160 263 161 264
rect 159 263 160 264
rect 158 263 159 264
rect 157 263 158 264
rect 156 263 157 264
rect 155 263 156 264
rect 154 263 155 264
rect 153 263 154 264
rect 152 263 153 264
rect 151 263 152 264
rect 150 263 151 264
rect 149 263 150 264
rect 148 263 149 264
rect 147 263 148 264
rect 146 263 147 264
rect 145 263 146 264
rect 144 263 145 264
rect 143 263 144 264
rect 142 263 143 264
rect 141 263 142 264
rect 140 263 141 264
rect 139 263 140 264
rect 138 263 139 264
rect 137 263 138 264
rect 136 263 137 264
rect 135 263 136 264
rect 134 263 135 264
rect 133 263 134 264
rect 132 263 133 264
rect 131 263 132 264
rect 130 263 131 264
rect 129 263 130 264
rect 128 263 129 264
rect 127 263 128 264
rect 126 263 127 264
rect 125 263 126 264
rect 124 263 125 264
rect 123 263 124 264
rect 122 263 123 264
rect 109 263 110 264
rect 108 263 109 264
rect 107 263 108 264
rect 106 263 107 264
rect 105 263 106 264
rect 104 263 105 264
rect 103 263 104 264
rect 102 263 103 264
rect 101 263 102 264
rect 100 263 101 264
rect 99 263 100 264
rect 98 263 99 264
rect 97 263 98 264
rect 96 263 97 264
rect 95 263 96 264
rect 94 263 95 264
rect 93 263 94 264
rect 92 263 93 264
rect 91 263 92 264
rect 90 263 91 264
rect 89 263 90 264
rect 88 263 89 264
rect 87 263 88 264
rect 86 263 87 264
rect 85 263 86 264
rect 84 263 85 264
rect 83 263 84 264
rect 82 263 83 264
rect 81 263 82 264
rect 80 263 81 264
rect 79 263 80 264
rect 78 263 79 264
rect 77 263 78 264
rect 76 263 77 264
rect 75 263 76 264
rect 74 263 75 264
rect 73 263 74 264
rect 72 263 73 264
rect 55 263 56 264
rect 54 263 55 264
rect 53 263 54 264
rect 52 263 53 264
rect 51 263 52 264
rect 50 263 51 264
rect 49 263 50 264
rect 48 263 49 264
rect 47 263 48 264
rect 46 263 47 264
rect 45 263 46 264
rect 44 263 45 264
rect 43 263 44 264
rect 42 263 43 264
rect 41 263 42 264
rect 40 263 41 264
rect 39 263 40 264
rect 38 263 39 264
rect 37 263 38 264
rect 36 263 37 264
rect 35 263 36 264
rect 34 263 35 264
rect 22 263 23 264
rect 21 263 22 264
rect 20 263 21 264
rect 19 263 20 264
rect 18 263 19 264
rect 17 263 18 264
rect 16 263 17 264
rect 15 263 16 264
rect 14 263 15 264
rect 13 263 14 264
rect 12 263 13 264
rect 11 263 12 264
rect 10 263 11 264
rect 9 263 10 264
rect 8 263 9 264
rect 7 263 8 264
rect 6 263 7 264
rect 5 263 6 264
rect 4 263 5 264
rect 3 263 4 264
rect 2 263 3 264
rect 1 263 2 264
rect 478 264 479 265
rect 458 264 459 265
rect 297 264 298 265
rect 296 264 297 265
rect 295 264 296 265
rect 294 264 295 265
rect 293 264 294 265
rect 292 264 293 265
rect 291 264 292 265
rect 290 264 291 265
rect 289 264 290 265
rect 288 264 289 265
rect 287 264 288 265
rect 286 264 287 265
rect 285 264 286 265
rect 284 264 285 265
rect 283 264 284 265
rect 282 264 283 265
rect 281 264 282 265
rect 280 264 281 265
rect 279 264 280 265
rect 278 264 279 265
rect 277 264 278 265
rect 276 264 277 265
rect 275 264 276 265
rect 274 264 275 265
rect 273 264 274 265
rect 272 264 273 265
rect 271 264 272 265
rect 270 264 271 265
rect 269 264 270 265
rect 268 264 269 265
rect 267 264 268 265
rect 266 264 267 265
rect 265 264 266 265
rect 264 264 265 265
rect 263 264 264 265
rect 262 264 263 265
rect 261 264 262 265
rect 260 264 261 265
rect 259 264 260 265
rect 258 264 259 265
rect 257 264 258 265
rect 256 264 257 265
rect 255 264 256 265
rect 254 264 255 265
rect 253 264 254 265
rect 252 264 253 265
rect 251 264 252 265
rect 250 264 251 265
rect 249 264 250 265
rect 248 264 249 265
rect 247 264 248 265
rect 246 264 247 265
rect 245 264 246 265
rect 244 264 245 265
rect 243 264 244 265
rect 242 264 243 265
rect 241 264 242 265
rect 240 264 241 265
rect 239 264 240 265
rect 238 264 239 265
rect 237 264 238 265
rect 236 264 237 265
rect 235 264 236 265
rect 234 264 235 265
rect 233 264 234 265
rect 232 264 233 265
rect 231 264 232 265
rect 230 264 231 265
rect 229 264 230 265
rect 228 264 229 265
rect 227 264 228 265
rect 226 264 227 265
rect 225 264 226 265
rect 224 264 225 265
rect 203 264 204 265
rect 202 264 203 265
rect 201 264 202 265
rect 200 264 201 265
rect 199 264 200 265
rect 198 264 199 265
rect 197 264 198 265
rect 196 264 197 265
rect 195 264 196 265
rect 194 264 195 265
rect 193 264 194 265
rect 192 264 193 265
rect 191 264 192 265
rect 190 264 191 265
rect 189 264 190 265
rect 188 264 189 265
rect 187 264 188 265
rect 186 264 187 265
rect 185 264 186 265
rect 184 264 185 265
rect 183 264 184 265
rect 182 264 183 265
rect 181 264 182 265
rect 180 264 181 265
rect 179 264 180 265
rect 178 264 179 265
rect 177 264 178 265
rect 176 264 177 265
rect 175 264 176 265
rect 174 264 175 265
rect 173 264 174 265
rect 172 264 173 265
rect 171 264 172 265
rect 170 264 171 265
rect 169 264 170 265
rect 168 264 169 265
rect 167 264 168 265
rect 166 264 167 265
rect 165 264 166 265
rect 164 264 165 265
rect 163 264 164 265
rect 162 264 163 265
rect 161 264 162 265
rect 160 264 161 265
rect 159 264 160 265
rect 158 264 159 265
rect 157 264 158 265
rect 156 264 157 265
rect 155 264 156 265
rect 154 264 155 265
rect 153 264 154 265
rect 152 264 153 265
rect 151 264 152 265
rect 150 264 151 265
rect 149 264 150 265
rect 148 264 149 265
rect 147 264 148 265
rect 146 264 147 265
rect 145 264 146 265
rect 144 264 145 265
rect 143 264 144 265
rect 142 264 143 265
rect 141 264 142 265
rect 140 264 141 265
rect 139 264 140 265
rect 138 264 139 265
rect 137 264 138 265
rect 136 264 137 265
rect 135 264 136 265
rect 134 264 135 265
rect 133 264 134 265
rect 132 264 133 265
rect 131 264 132 265
rect 130 264 131 265
rect 129 264 130 265
rect 128 264 129 265
rect 127 264 128 265
rect 126 264 127 265
rect 125 264 126 265
rect 124 264 125 265
rect 123 264 124 265
rect 122 264 123 265
rect 109 264 110 265
rect 108 264 109 265
rect 107 264 108 265
rect 106 264 107 265
rect 105 264 106 265
rect 104 264 105 265
rect 103 264 104 265
rect 102 264 103 265
rect 101 264 102 265
rect 100 264 101 265
rect 99 264 100 265
rect 98 264 99 265
rect 97 264 98 265
rect 96 264 97 265
rect 95 264 96 265
rect 94 264 95 265
rect 93 264 94 265
rect 92 264 93 265
rect 91 264 92 265
rect 90 264 91 265
rect 89 264 90 265
rect 88 264 89 265
rect 87 264 88 265
rect 86 264 87 265
rect 85 264 86 265
rect 84 264 85 265
rect 83 264 84 265
rect 82 264 83 265
rect 81 264 82 265
rect 80 264 81 265
rect 79 264 80 265
rect 78 264 79 265
rect 77 264 78 265
rect 76 264 77 265
rect 75 264 76 265
rect 74 264 75 265
rect 73 264 74 265
rect 72 264 73 265
rect 56 264 57 265
rect 55 264 56 265
rect 54 264 55 265
rect 53 264 54 265
rect 52 264 53 265
rect 51 264 52 265
rect 50 264 51 265
rect 49 264 50 265
rect 48 264 49 265
rect 47 264 48 265
rect 46 264 47 265
rect 45 264 46 265
rect 44 264 45 265
rect 43 264 44 265
rect 42 264 43 265
rect 41 264 42 265
rect 40 264 41 265
rect 39 264 40 265
rect 38 264 39 265
rect 37 264 38 265
rect 36 264 37 265
rect 35 264 36 265
rect 34 264 35 265
rect 23 264 24 265
rect 22 264 23 265
rect 21 264 22 265
rect 20 264 21 265
rect 19 264 20 265
rect 18 264 19 265
rect 17 264 18 265
rect 16 264 17 265
rect 15 264 16 265
rect 14 264 15 265
rect 13 264 14 265
rect 12 264 13 265
rect 11 264 12 265
rect 10 264 11 265
rect 9 264 10 265
rect 8 264 9 265
rect 7 264 8 265
rect 6 264 7 265
rect 5 264 6 265
rect 4 264 5 265
rect 3 264 4 265
rect 2 264 3 265
rect 1 264 2 265
rect 478 265 479 266
rect 458 265 459 266
rect 297 265 298 266
rect 296 265 297 266
rect 295 265 296 266
rect 294 265 295 266
rect 293 265 294 266
rect 292 265 293 266
rect 291 265 292 266
rect 290 265 291 266
rect 289 265 290 266
rect 288 265 289 266
rect 287 265 288 266
rect 286 265 287 266
rect 285 265 286 266
rect 284 265 285 266
rect 283 265 284 266
rect 282 265 283 266
rect 281 265 282 266
rect 280 265 281 266
rect 279 265 280 266
rect 278 265 279 266
rect 277 265 278 266
rect 276 265 277 266
rect 275 265 276 266
rect 274 265 275 266
rect 273 265 274 266
rect 272 265 273 266
rect 271 265 272 266
rect 270 265 271 266
rect 269 265 270 266
rect 268 265 269 266
rect 267 265 268 266
rect 266 265 267 266
rect 265 265 266 266
rect 264 265 265 266
rect 263 265 264 266
rect 262 265 263 266
rect 261 265 262 266
rect 260 265 261 266
rect 259 265 260 266
rect 258 265 259 266
rect 257 265 258 266
rect 256 265 257 266
rect 255 265 256 266
rect 254 265 255 266
rect 253 265 254 266
rect 252 265 253 266
rect 251 265 252 266
rect 250 265 251 266
rect 249 265 250 266
rect 248 265 249 266
rect 247 265 248 266
rect 246 265 247 266
rect 245 265 246 266
rect 244 265 245 266
rect 243 265 244 266
rect 242 265 243 266
rect 241 265 242 266
rect 240 265 241 266
rect 239 265 240 266
rect 238 265 239 266
rect 237 265 238 266
rect 236 265 237 266
rect 235 265 236 266
rect 234 265 235 266
rect 233 265 234 266
rect 232 265 233 266
rect 231 265 232 266
rect 230 265 231 266
rect 229 265 230 266
rect 228 265 229 266
rect 227 265 228 266
rect 226 265 227 266
rect 225 265 226 266
rect 224 265 225 266
rect 203 265 204 266
rect 202 265 203 266
rect 201 265 202 266
rect 200 265 201 266
rect 199 265 200 266
rect 198 265 199 266
rect 197 265 198 266
rect 196 265 197 266
rect 195 265 196 266
rect 194 265 195 266
rect 193 265 194 266
rect 192 265 193 266
rect 191 265 192 266
rect 190 265 191 266
rect 189 265 190 266
rect 188 265 189 266
rect 187 265 188 266
rect 186 265 187 266
rect 185 265 186 266
rect 184 265 185 266
rect 183 265 184 266
rect 182 265 183 266
rect 181 265 182 266
rect 180 265 181 266
rect 179 265 180 266
rect 178 265 179 266
rect 177 265 178 266
rect 176 265 177 266
rect 175 265 176 266
rect 174 265 175 266
rect 173 265 174 266
rect 172 265 173 266
rect 171 265 172 266
rect 170 265 171 266
rect 169 265 170 266
rect 168 265 169 266
rect 167 265 168 266
rect 166 265 167 266
rect 165 265 166 266
rect 164 265 165 266
rect 163 265 164 266
rect 162 265 163 266
rect 161 265 162 266
rect 160 265 161 266
rect 159 265 160 266
rect 158 265 159 266
rect 157 265 158 266
rect 156 265 157 266
rect 155 265 156 266
rect 154 265 155 266
rect 153 265 154 266
rect 152 265 153 266
rect 151 265 152 266
rect 150 265 151 266
rect 149 265 150 266
rect 148 265 149 266
rect 147 265 148 266
rect 146 265 147 266
rect 145 265 146 266
rect 144 265 145 266
rect 143 265 144 266
rect 142 265 143 266
rect 141 265 142 266
rect 140 265 141 266
rect 139 265 140 266
rect 138 265 139 266
rect 137 265 138 266
rect 136 265 137 266
rect 135 265 136 266
rect 134 265 135 266
rect 133 265 134 266
rect 132 265 133 266
rect 131 265 132 266
rect 130 265 131 266
rect 129 265 130 266
rect 128 265 129 266
rect 127 265 128 266
rect 126 265 127 266
rect 125 265 126 266
rect 124 265 125 266
rect 123 265 124 266
rect 122 265 123 266
rect 109 265 110 266
rect 108 265 109 266
rect 107 265 108 266
rect 106 265 107 266
rect 105 265 106 266
rect 104 265 105 266
rect 103 265 104 266
rect 102 265 103 266
rect 101 265 102 266
rect 100 265 101 266
rect 99 265 100 266
rect 98 265 99 266
rect 97 265 98 266
rect 96 265 97 266
rect 95 265 96 266
rect 94 265 95 266
rect 93 265 94 266
rect 92 265 93 266
rect 91 265 92 266
rect 90 265 91 266
rect 89 265 90 266
rect 88 265 89 266
rect 87 265 88 266
rect 86 265 87 266
rect 85 265 86 266
rect 84 265 85 266
rect 83 265 84 266
rect 82 265 83 266
rect 81 265 82 266
rect 80 265 81 266
rect 79 265 80 266
rect 78 265 79 266
rect 77 265 78 266
rect 76 265 77 266
rect 75 265 76 266
rect 74 265 75 266
rect 73 265 74 266
rect 56 265 57 266
rect 55 265 56 266
rect 54 265 55 266
rect 53 265 54 266
rect 52 265 53 266
rect 51 265 52 266
rect 50 265 51 266
rect 49 265 50 266
rect 48 265 49 266
rect 47 265 48 266
rect 46 265 47 266
rect 45 265 46 266
rect 44 265 45 266
rect 43 265 44 266
rect 42 265 43 266
rect 41 265 42 266
rect 40 265 41 266
rect 39 265 40 266
rect 38 265 39 266
rect 37 265 38 266
rect 36 265 37 266
rect 35 265 36 266
rect 34 265 35 266
rect 23 265 24 266
rect 22 265 23 266
rect 21 265 22 266
rect 20 265 21 266
rect 19 265 20 266
rect 18 265 19 266
rect 17 265 18 266
rect 16 265 17 266
rect 15 265 16 266
rect 14 265 15 266
rect 13 265 14 266
rect 12 265 13 266
rect 11 265 12 266
rect 10 265 11 266
rect 9 265 10 266
rect 8 265 9 266
rect 7 265 8 266
rect 6 265 7 266
rect 5 265 6 266
rect 4 265 5 266
rect 3 265 4 266
rect 2 265 3 266
rect 1 265 2 266
rect 478 266 479 267
rect 477 266 478 267
rect 459 266 460 267
rect 458 266 459 267
rect 296 266 297 267
rect 295 266 296 267
rect 294 266 295 267
rect 293 266 294 267
rect 292 266 293 267
rect 291 266 292 267
rect 290 266 291 267
rect 289 266 290 267
rect 288 266 289 267
rect 287 266 288 267
rect 286 266 287 267
rect 285 266 286 267
rect 284 266 285 267
rect 283 266 284 267
rect 282 266 283 267
rect 281 266 282 267
rect 280 266 281 267
rect 279 266 280 267
rect 278 266 279 267
rect 277 266 278 267
rect 276 266 277 267
rect 275 266 276 267
rect 274 266 275 267
rect 273 266 274 267
rect 272 266 273 267
rect 271 266 272 267
rect 270 266 271 267
rect 269 266 270 267
rect 268 266 269 267
rect 267 266 268 267
rect 266 266 267 267
rect 265 266 266 267
rect 264 266 265 267
rect 263 266 264 267
rect 262 266 263 267
rect 261 266 262 267
rect 260 266 261 267
rect 259 266 260 267
rect 258 266 259 267
rect 257 266 258 267
rect 256 266 257 267
rect 255 266 256 267
rect 254 266 255 267
rect 253 266 254 267
rect 252 266 253 267
rect 251 266 252 267
rect 250 266 251 267
rect 249 266 250 267
rect 248 266 249 267
rect 247 266 248 267
rect 246 266 247 267
rect 245 266 246 267
rect 244 266 245 267
rect 243 266 244 267
rect 242 266 243 267
rect 241 266 242 267
rect 240 266 241 267
rect 239 266 240 267
rect 238 266 239 267
rect 237 266 238 267
rect 236 266 237 267
rect 235 266 236 267
rect 234 266 235 267
rect 233 266 234 267
rect 232 266 233 267
rect 231 266 232 267
rect 230 266 231 267
rect 229 266 230 267
rect 228 266 229 267
rect 227 266 228 267
rect 226 266 227 267
rect 225 266 226 267
rect 224 266 225 267
rect 223 266 224 267
rect 202 266 203 267
rect 201 266 202 267
rect 200 266 201 267
rect 199 266 200 267
rect 198 266 199 267
rect 197 266 198 267
rect 196 266 197 267
rect 195 266 196 267
rect 194 266 195 267
rect 193 266 194 267
rect 192 266 193 267
rect 191 266 192 267
rect 190 266 191 267
rect 189 266 190 267
rect 188 266 189 267
rect 187 266 188 267
rect 186 266 187 267
rect 185 266 186 267
rect 184 266 185 267
rect 183 266 184 267
rect 182 266 183 267
rect 181 266 182 267
rect 180 266 181 267
rect 179 266 180 267
rect 178 266 179 267
rect 177 266 178 267
rect 176 266 177 267
rect 175 266 176 267
rect 174 266 175 267
rect 173 266 174 267
rect 172 266 173 267
rect 171 266 172 267
rect 170 266 171 267
rect 169 266 170 267
rect 168 266 169 267
rect 167 266 168 267
rect 166 266 167 267
rect 165 266 166 267
rect 164 266 165 267
rect 163 266 164 267
rect 162 266 163 267
rect 161 266 162 267
rect 160 266 161 267
rect 159 266 160 267
rect 158 266 159 267
rect 157 266 158 267
rect 156 266 157 267
rect 155 266 156 267
rect 154 266 155 267
rect 153 266 154 267
rect 152 266 153 267
rect 151 266 152 267
rect 150 266 151 267
rect 149 266 150 267
rect 148 266 149 267
rect 147 266 148 267
rect 146 266 147 267
rect 145 266 146 267
rect 144 266 145 267
rect 143 266 144 267
rect 142 266 143 267
rect 141 266 142 267
rect 140 266 141 267
rect 139 266 140 267
rect 138 266 139 267
rect 137 266 138 267
rect 136 266 137 267
rect 135 266 136 267
rect 134 266 135 267
rect 133 266 134 267
rect 132 266 133 267
rect 131 266 132 267
rect 130 266 131 267
rect 129 266 130 267
rect 128 266 129 267
rect 127 266 128 267
rect 126 266 127 267
rect 125 266 126 267
rect 124 266 125 267
rect 123 266 124 267
rect 122 266 123 267
rect 109 266 110 267
rect 108 266 109 267
rect 107 266 108 267
rect 106 266 107 267
rect 105 266 106 267
rect 104 266 105 267
rect 103 266 104 267
rect 102 266 103 267
rect 101 266 102 267
rect 100 266 101 267
rect 99 266 100 267
rect 98 266 99 267
rect 97 266 98 267
rect 96 266 97 267
rect 95 266 96 267
rect 94 266 95 267
rect 93 266 94 267
rect 92 266 93 267
rect 91 266 92 267
rect 90 266 91 267
rect 89 266 90 267
rect 88 266 89 267
rect 87 266 88 267
rect 86 266 87 267
rect 85 266 86 267
rect 84 266 85 267
rect 83 266 84 267
rect 82 266 83 267
rect 81 266 82 267
rect 80 266 81 267
rect 79 266 80 267
rect 78 266 79 267
rect 77 266 78 267
rect 76 266 77 267
rect 75 266 76 267
rect 74 266 75 267
rect 73 266 74 267
rect 57 266 58 267
rect 56 266 57 267
rect 55 266 56 267
rect 54 266 55 267
rect 53 266 54 267
rect 52 266 53 267
rect 51 266 52 267
rect 50 266 51 267
rect 49 266 50 267
rect 48 266 49 267
rect 47 266 48 267
rect 46 266 47 267
rect 45 266 46 267
rect 44 266 45 267
rect 43 266 44 267
rect 42 266 43 267
rect 41 266 42 267
rect 40 266 41 267
rect 39 266 40 267
rect 38 266 39 267
rect 37 266 38 267
rect 36 266 37 267
rect 35 266 36 267
rect 34 266 35 267
rect 23 266 24 267
rect 22 266 23 267
rect 21 266 22 267
rect 20 266 21 267
rect 19 266 20 267
rect 18 266 19 267
rect 17 266 18 267
rect 16 266 17 267
rect 15 266 16 267
rect 14 266 15 267
rect 13 266 14 267
rect 12 266 13 267
rect 11 266 12 267
rect 10 266 11 267
rect 9 266 10 267
rect 8 266 9 267
rect 7 266 8 267
rect 6 266 7 267
rect 5 266 6 267
rect 4 266 5 267
rect 3 266 4 267
rect 2 266 3 267
rect 1 266 2 267
rect 478 267 479 268
rect 477 267 478 268
rect 476 267 477 268
rect 475 267 476 268
rect 474 267 475 268
rect 473 267 474 268
rect 472 267 473 268
rect 471 267 472 268
rect 470 267 471 268
rect 469 267 470 268
rect 468 267 469 268
rect 467 267 468 268
rect 466 267 467 268
rect 465 267 466 268
rect 464 267 465 268
rect 463 267 464 268
rect 462 267 463 268
rect 461 267 462 268
rect 460 267 461 268
rect 459 267 460 268
rect 458 267 459 268
rect 295 267 296 268
rect 294 267 295 268
rect 293 267 294 268
rect 292 267 293 268
rect 291 267 292 268
rect 290 267 291 268
rect 289 267 290 268
rect 288 267 289 268
rect 287 267 288 268
rect 286 267 287 268
rect 285 267 286 268
rect 284 267 285 268
rect 283 267 284 268
rect 282 267 283 268
rect 281 267 282 268
rect 280 267 281 268
rect 279 267 280 268
rect 278 267 279 268
rect 277 267 278 268
rect 276 267 277 268
rect 275 267 276 268
rect 274 267 275 268
rect 273 267 274 268
rect 272 267 273 268
rect 271 267 272 268
rect 270 267 271 268
rect 269 267 270 268
rect 268 267 269 268
rect 267 267 268 268
rect 266 267 267 268
rect 265 267 266 268
rect 264 267 265 268
rect 263 267 264 268
rect 262 267 263 268
rect 261 267 262 268
rect 260 267 261 268
rect 259 267 260 268
rect 258 267 259 268
rect 257 267 258 268
rect 256 267 257 268
rect 255 267 256 268
rect 254 267 255 268
rect 253 267 254 268
rect 252 267 253 268
rect 251 267 252 268
rect 250 267 251 268
rect 249 267 250 268
rect 248 267 249 268
rect 247 267 248 268
rect 246 267 247 268
rect 245 267 246 268
rect 244 267 245 268
rect 243 267 244 268
rect 242 267 243 268
rect 241 267 242 268
rect 240 267 241 268
rect 239 267 240 268
rect 238 267 239 268
rect 237 267 238 268
rect 236 267 237 268
rect 235 267 236 268
rect 234 267 235 268
rect 233 267 234 268
rect 232 267 233 268
rect 231 267 232 268
rect 230 267 231 268
rect 229 267 230 268
rect 228 267 229 268
rect 227 267 228 268
rect 226 267 227 268
rect 225 267 226 268
rect 224 267 225 268
rect 223 267 224 268
rect 202 267 203 268
rect 201 267 202 268
rect 200 267 201 268
rect 199 267 200 268
rect 198 267 199 268
rect 197 267 198 268
rect 196 267 197 268
rect 195 267 196 268
rect 194 267 195 268
rect 193 267 194 268
rect 192 267 193 268
rect 191 267 192 268
rect 190 267 191 268
rect 189 267 190 268
rect 188 267 189 268
rect 187 267 188 268
rect 186 267 187 268
rect 185 267 186 268
rect 184 267 185 268
rect 183 267 184 268
rect 182 267 183 268
rect 181 267 182 268
rect 180 267 181 268
rect 179 267 180 268
rect 178 267 179 268
rect 177 267 178 268
rect 176 267 177 268
rect 175 267 176 268
rect 174 267 175 268
rect 173 267 174 268
rect 172 267 173 268
rect 171 267 172 268
rect 170 267 171 268
rect 169 267 170 268
rect 168 267 169 268
rect 167 267 168 268
rect 166 267 167 268
rect 165 267 166 268
rect 164 267 165 268
rect 163 267 164 268
rect 162 267 163 268
rect 161 267 162 268
rect 160 267 161 268
rect 159 267 160 268
rect 158 267 159 268
rect 157 267 158 268
rect 156 267 157 268
rect 155 267 156 268
rect 154 267 155 268
rect 153 267 154 268
rect 152 267 153 268
rect 151 267 152 268
rect 150 267 151 268
rect 149 267 150 268
rect 148 267 149 268
rect 147 267 148 268
rect 146 267 147 268
rect 145 267 146 268
rect 144 267 145 268
rect 143 267 144 268
rect 142 267 143 268
rect 141 267 142 268
rect 140 267 141 268
rect 139 267 140 268
rect 138 267 139 268
rect 137 267 138 268
rect 136 267 137 268
rect 135 267 136 268
rect 134 267 135 268
rect 133 267 134 268
rect 132 267 133 268
rect 131 267 132 268
rect 130 267 131 268
rect 129 267 130 268
rect 128 267 129 268
rect 127 267 128 268
rect 126 267 127 268
rect 125 267 126 268
rect 124 267 125 268
rect 123 267 124 268
rect 109 267 110 268
rect 108 267 109 268
rect 107 267 108 268
rect 106 267 107 268
rect 105 267 106 268
rect 104 267 105 268
rect 103 267 104 268
rect 102 267 103 268
rect 101 267 102 268
rect 100 267 101 268
rect 99 267 100 268
rect 98 267 99 268
rect 97 267 98 268
rect 96 267 97 268
rect 95 267 96 268
rect 94 267 95 268
rect 93 267 94 268
rect 92 267 93 268
rect 91 267 92 268
rect 90 267 91 268
rect 89 267 90 268
rect 88 267 89 268
rect 87 267 88 268
rect 86 267 87 268
rect 85 267 86 268
rect 84 267 85 268
rect 83 267 84 268
rect 82 267 83 268
rect 81 267 82 268
rect 80 267 81 268
rect 79 267 80 268
rect 78 267 79 268
rect 77 267 78 268
rect 76 267 77 268
rect 75 267 76 268
rect 74 267 75 268
rect 57 267 58 268
rect 56 267 57 268
rect 55 267 56 268
rect 54 267 55 268
rect 53 267 54 268
rect 52 267 53 268
rect 51 267 52 268
rect 50 267 51 268
rect 49 267 50 268
rect 48 267 49 268
rect 47 267 48 268
rect 46 267 47 268
rect 45 267 46 268
rect 44 267 45 268
rect 43 267 44 268
rect 42 267 43 268
rect 41 267 42 268
rect 40 267 41 268
rect 39 267 40 268
rect 38 267 39 268
rect 37 267 38 268
rect 36 267 37 268
rect 35 267 36 268
rect 23 267 24 268
rect 22 267 23 268
rect 21 267 22 268
rect 20 267 21 268
rect 19 267 20 268
rect 18 267 19 268
rect 17 267 18 268
rect 16 267 17 268
rect 15 267 16 268
rect 14 267 15 268
rect 13 267 14 268
rect 12 267 13 268
rect 11 267 12 268
rect 10 267 11 268
rect 9 267 10 268
rect 8 267 9 268
rect 7 267 8 268
rect 6 267 7 268
rect 5 267 6 268
rect 4 267 5 268
rect 3 267 4 268
rect 2 267 3 268
rect 1 267 2 268
rect 478 268 479 269
rect 477 268 478 269
rect 476 268 477 269
rect 475 268 476 269
rect 474 268 475 269
rect 473 268 474 269
rect 472 268 473 269
rect 471 268 472 269
rect 470 268 471 269
rect 469 268 470 269
rect 468 268 469 269
rect 467 268 468 269
rect 466 268 467 269
rect 465 268 466 269
rect 464 268 465 269
rect 463 268 464 269
rect 462 268 463 269
rect 461 268 462 269
rect 460 268 461 269
rect 459 268 460 269
rect 458 268 459 269
rect 295 268 296 269
rect 294 268 295 269
rect 293 268 294 269
rect 292 268 293 269
rect 291 268 292 269
rect 290 268 291 269
rect 289 268 290 269
rect 288 268 289 269
rect 287 268 288 269
rect 286 268 287 269
rect 285 268 286 269
rect 284 268 285 269
rect 283 268 284 269
rect 282 268 283 269
rect 281 268 282 269
rect 280 268 281 269
rect 279 268 280 269
rect 278 268 279 269
rect 277 268 278 269
rect 276 268 277 269
rect 275 268 276 269
rect 274 268 275 269
rect 273 268 274 269
rect 272 268 273 269
rect 271 268 272 269
rect 270 268 271 269
rect 269 268 270 269
rect 268 268 269 269
rect 267 268 268 269
rect 266 268 267 269
rect 265 268 266 269
rect 264 268 265 269
rect 263 268 264 269
rect 262 268 263 269
rect 261 268 262 269
rect 260 268 261 269
rect 259 268 260 269
rect 258 268 259 269
rect 257 268 258 269
rect 256 268 257 269
rect 255 268 256 269
rect 254 268 255 269
rect 253 268 254 269
rect 252 268 253 269
rect 251 268 252 269
rect 250 268 251 269
rect 249 268 250 269
rect 248 268 249 269
rect 247 268 248 269
rect 246 268 247 269
rect 245 268 246 269
rect 244 268 245 269
rect 243 268 244 269
rect 242 268 243 269
rect 241 268 242 269
rect 240 268 241 269
rect 239 268 240 269
rect 238 268 239 269
rect 237 268 238 269
rect 236 268 237 269
rect 235 268 236 269
rect 234 268 235 269
rect 233 268 234 269
rect 232 268 233 269
rect 231 268 232 269
rect 230 268 231 269
rect 229 268 230 269
rect 228 268 229 269
rect 227 268 228 269
rect 226 268 227 269
rect 225 268 226 269
rect 224 268 225 269
rect 223 268 224 269
rect 202 268 203 269
rect 201 268 202 269
rect 200 268 201 269
rect 199 268 200 269
rect 198 268 199 269
rect 197 268 198 269
rect 196 268 197 269
rect 195 268 196 269
rect 194 268 195 269
rect 193 268 194 269
rect 192 268 193 269
rect 191 268 192 269
rect 190 268 191 269
rect 189 268 190 269
rect 188 268 189 269
rect 187 268 188 269
rect 186 268 187 269
rect 185 268 186 269
rect 184 268 185 269
rect 183 268 184 269
rect 182 268 183 269
rect 181 268 182 269
rect 180 268 181 269
rect 179 268 180 269
rect 178 268 179 269
rect 177 268 178 269
rect 176 268 177 269
rect 175 268 176 269
rect 174 268 175 269
rect 173 268 174 269
rect 172 268 173 269
rect 171 268 172 269
rect 170 268 171 269
rect 169 268 170 269
rect 168 268 169 269
rect 167 268 168 269
rect 166 268 167 269
rect 165 268 166 269
rect 164 268 165 269
rect 163 268 164 269
rect 162 268 163 269
rect 161 268 162 269
rect 160 268 161 269
rect 159 268 160 269
rect 158 268 159 269
rect 157 268 158 269
rect 156 268 157 269
rect 155 268 156 269
rect 154 268 155 269
rect 153 268 154 269
rect 152 268 153 269
rect 151 268 152 269
rect 150 268 151 269
rect 149 268 150 269
rect 148 268 149 269
rect 147 268 148 269
rect 146 268 147 269
rect 145 268 146 269
rect 144 268 145 269
rect 143 268 144 269
rect 142 268 143 269
rect 141 268 142 269
rect 140 268 141 269
rect 139 268 140 269
rect 138 268 139 269
rect 137 268 138 269
rect 136 268 137 269
rect 135 268 136 269
rect 134 268 135 269
rect 133 268 134 269
rect 132 268 133 269
rect 131 268 132 269
rect 130 268 131 269
rect 129 268 130 269
rect 128 268 129 269
rect 127 268 128 269
rect 126 268 127 269
rect 125 268 126 269
rect 124 268 125 269
rect 123 268 124 269
rect 109 268 110 269
rect 108 268 109 269
rect 107 268 108 269
rect 106 268 107 269
rect 105 268 106 269
rect 104 268 105 269
rect 103 268 104 269
rect 102 268 103 269
rect 101 268 102 269
rect 100 268 101 269
rect 99 268 100 269
rect 98 268 99 269
rect 97 268 98 269
rect 96 268 97 269
rect 95 268 96 269
rect 94 268 95 269
rect 93 268 94 269
rect 92 268 93 269
rect 91 268 92 269
rect 90 268 91 269
rect 89 268 90 269
rect 88 268 89 269
rect 87 268 88 269
rect 86 268 87 269
rect 85 268 86 269
rect 84 268 85 269
rect 83 268 84 269
rect 82 268 83 269
rect 81 268 82 269
rect 80 268 81 269
rect 79 268 80 269
rect 78 268 79 269
rect 77 268 78 269
rect 76 268 77 269
rect 75 268 76 269
rect 74 268 75 269
rect 57 268 58 269
rect 56 268 57 269
rect 55 268 56 269
rect 54 268 55 269
rect 53 268 54 269
rect 52 268 53 269
rect 51 268 52 269
rect 50 268 51 269
rect 49 268 50 269
rect 48 268 49 269
rect 47 268 48 269
rect 46 268 47 269
rect 45 268 46 269
rect 44 268 45 269
rect 43 268 44 269
rect 42 268 43 269
rect 41 268 42 269
rect 40 268 41 269
rect 39 268 40 269
rect 38 268 39 269
rect 37 268 38 269
rect 36 268 37 269
rect 35 268 36 269
rect 23 268 24 269
rect 22 268 23 269
rect 21 268 22 269
rect 20 268 21 269
rect 19 268 20 269
rect 18 268 19 269
rect 17 268 18 269
rect 16 268 17 269
rect 15 268 16 269
rect 14 268 15 269
rect 13 268 14 269
rect 12 268 13 269
rect 11 268 12 269
rect 10 268 11 269
rect 9 268 10 269
rect 8 268 9 269
rect 7 268 8 269
rect 6 268 7 269
rect 5 268 6 269
rect 4 268 5 269
rect 3 268 4 269
rect 2 268 3 269
rect 1 268 2 269
rect 478 269 479 270
rect 477 269 478 270
rect 476 269 477 270
rect 475 269 476 270
rect 474 269 475 270
rect 473 269 474 270
rect 472 269 473 270
rect 471 269 472 270
rect 470 269 471 270
rect 469 269 470 270
rect 468 269 469 270
rect 467 269 468 270
rect 466 269 467 270
rect 465 269 466 270
rect 464 269 465 270
rect 463 269 464 270
rect 462 269 463 270
rect 461 269 462 270
rect 460 269 461 270
rect 459 269 460 270
rect 458 269 459 270
rect 294 269 295 270
rect 293 269 294 270
rect 292 269 293 270
rect 291 269 292 270
rect 290 269 291 270
rect 289 269 290 270
rect 288 269 289 270
rect 287 269 288 270
rect 286 269 287 270
rect 285 269 286 270
rect 284 269 285 270
rect 283 269 284 270
rect 282 269 283 270
rect 281 269 282 270
rect 280 269 281 270
rect 279 269 280 270
rect 278 269 279 270
rect 277 269 278 270
rect 276 269 277 270
rect 275 269 276 270
rect 274 269 275 270
rect 273 269 274 270
rect 272 269 273 270
rect 271 269 272 270
rect 270 269 271 270
rect 269 269 270 270
rect 268 269 269 270
rect 267 269 268 270
rect 266 269 267 270
rect 265 269 266 270
rect 264 269 265 270
rect 263 269 264 270
rect 262 269 263 270
rect 261 269 262 270
rect 260 269 261 270
rect 259 269 260 270
rect 258 269 259 270
rect 257 269 258 270
rect 256 269 257 270
rect 255 269 256 270
rect 254 269 255 270
rect 253 269 254 270
rect 252 269 253 270
rect 251 269 252 270
rect 250 269 251 270
rect 249 269 250 270
rect 248 269 249 270
rect 247 269 248 270
rect 246 269 247 270
rect 245 269 246 270
rect 244 269 245 270
rect 243 269 244 270
rect 242 269 243 270
rect 241 269 242 270
rect 240 269 241 270
rect 239 269 240 270
rect 238 269 239 270
rect 237 269 238 270
rect 236 269 237 270
rect 235 269 236 270
rect 234 269 235 270
rect 233 269 234 270
rect 232 269 233 270
rect 231 269 232 270
rect 230 269 231 270
rect 229 269 230 270
rect 228 269 229 270
rect 227 269 228 270
rect 226 269 227 270
rect 225 269 226 270
rect 224 269 225 270
rect 223 269 224 270
rect 222 269 223 270
rect 201 269 202 270
rect 200 269 201 270
rect 199 269 200 270
rect 198 269 199 270
rect 197 269 198 270
rect 196 269 197 270
rect 195 269 196 270
rect 194 269 195 270
rect 193 269 194 270
rect 192 269 193 270
rect 191 269 192 270
rect 190 269 191 270
rect 189 269 190 270
rect 188 269 189 270
rect 187 269 188 270
rect 186 269 187 270
rect 185 269 186 270
rect 184 269 185 270
rect 183 269 184 270
rect 182 269 183 270
rect 181 269 182 270
rect 180 269 181 270
rect 179 269 180 270
rect 178 269 179 270
rect 177 269 178 270
rect 176 269 177 270
rect 175 269 176 270
rect 174 269 175 270
rect 173 269 174 270
rect 172 269 173 270
rect 171 269 172 270
rect 170 269 171 270
rect 169 269 170 270
rect 168 269 169 270
rect 167 269 168 270
rect 166 269 167 270
rect 165 269 166 270
rect 164 269 165 270
rect 163 269 164 270
rect 162 269 163 270
rect 161 269 162 270
rect 160 269 161 270
rect 159 269 160 270
rect 158 269 159 270
rect 157 269 158 270
rect 156 269 157 270
rect 155 269 156 270
rect 154 269 155 270
rect 153 269 154 270
rect 152 269 153 270
rect 151 269 152 270
rect 150 269 151 270
rect 149 269 150 270
rect 148 269 149 270
rect 147 269 148 270
rect 146 269 147 270
rect 145 269 146 270
rect 144 269 145 270
rect 143 269 144 270
rect 142 269 143 270
rect 141 269 142 270
rect 140 269 141 270
rect 139 269 140 270
rect 138 269 139 270
rect 137 269 138 270
rect 136 269 137 270
rect 135 269 136 270
rect 134 269 135 270
rect 133 269 134 270
rect 132 269 133 270
rect 131 269 132 270
rect 130 269 131 270
rect 129 269 130 270
rect 128 269 129 270
rect 127 269 128 270
rect 126 269 127 270
rect 125 269 126 270
rect 124 269 125 270
rect 110 269 111 270
rect 109 269 110 270
rect 108 269 109 270
rect 107 269 108 270
rect 106 269 107 270
rect 105 269 106 270
rect 104 269 105 270
rect 103 269 104 270
rect 102 269 103 270
rect 101 269 102 270
rect 100 269 101 270
rect 99 269 100 270
rect 98 269 99 270
rect 97 269 98 270
rect 96 269 97 270
rect 95 269 96 270
rect 94 269 95 270
rect 93 269 94 270
rect 92 269 93 270
rect 91 269 92 270
rect 90 269 91 270
rect 89 269 90 270
rect 88 269 89 270
rect 87 269 88 270
rect 86 269 87 270
rect 85 269 86 270
rect 84 269 85 270
rect 83 269 84 270
rect 82 269 83 270
rect 81 269 82 270
rect 80 269 81 270
rect 79 269 80 270
rect 78 269 79 270
rect 77 269 78 270
rect 76 269 77 270
rect 75 269 76 270
rect 58 269 59 270
rect 57 269 58 270
rect 56 269 57 270
rect 55 269 56 270
rect 54 269 55 270
rect 53 269 54 270
rect 52 269 53 270
rect 51 269 52 270
rect 50 269 51 270
rect 49 269 50 270
rect 48 269 49 270
rect 47 269 48 270
rect 46 269 47 270
rect 45 269 46 270
rect 44 269 45 270
rect 43 269 44 270
rect 42 269 43 270
rect 41 269 42 270
rect 40 269 41 270
rect 39 269 40 270
rect 38 269 39 270
rect 37 269 38 270
rect 36 269 37 270
rect 35 269 36 270
rect 24 269 25 270
rect 23 269 24 270
rect 22 269 23 270
rect 21 269 22 270
rect 20 269 21 270
rect 19 269 20 270
rect 18 269 19 270
rect 17 269 18 270
rect 16 269 17 270
rect 15 269 16 270
rect 14 269 15 270
rect 13 269 14 270
rect 12 269 13 270
rect 11 269 12 270
rect 10 269 11 270
rect 9 269 10 270
rect 8 269 9 270
rect 7 269 8 270
rect 6 269 7 270
rect 5 269 6 270
rect 4 269 5 270
rect 3 269 4 270
rect 2 269 3 270
rect 1 269 2 270
rect 478 270 479 271
rect 477 270 478 271
rect 476 270 477 271
rect 475 270 476 271
rect 474 270 475 271
rect 473 270 474 271
rect 472 270 473 271
rect 471 270 472 271
rect 470 270 471 271
rect 469 270 470 271
rect 468 270 469 271
rect 467 270 468 271
rect 466 270 467 271
rect 465 270 466 271
rect 464 270 465 271
rect 463 270 464 271
rect 462 270 463 271
rect 461 270 462 271
rect 460 270 461 271
rect 459 270 460 271
rect 458 270 459 271
rect 293 270 294 271
rect 292 270 293 271
rect 291 270 292 271
rect 290 270 291 271
rect 289 270 290 271
rect 288 270 289 271
rect 287 270 288 271
rect 286 270 287 271
rect 285 270 286 271
rect 284 270 285 271
rect 283 270 284 271
rect 282 270 283 271
rect 281 270 282 271
rect 280 270 281 271
rect 279 270 280 271
rect 278 270 279 271
rect 277 270 278 271
rect 276 270 277 271
rect 275 270 276 271
rect 274 270 275 271
rect 273 270 274 271
rect 272 270 273 271
rect 271 270 272 271
rect 270 270 271 271
rect 269 270 270 271
rect 268 270 269 271
rect 267 270 268 271
rect 266 270 267 271
rect 265 270 266 271
rect 264 270 265 271
rect 263 270 264 271
rect 262 270 263 271
rect 261 270 262 271
rect 260 270 261 271
rect 259 270 260 271
rect 258 270 259 271
rect 257 270 258 271
rect 256 270 257 271
rect 255 270 256 271
rect 254 270 255 271
rect 253 270 254 271
rect 252 270 253 271
rect 251 270 252 271
rect 250 270 251 271
rect 249 270 250 271
rect 248 270 249 271
rect 247 270 248 271
rect 246 270 247 271
rect 245 270 246 271
rect 244 270 245 271
rect 243 270 244 271
rect 242 270 243 271
rect 241 270 242 271
rect 240 270 241 271
rect 239 270 240 271
rect 238 270 239 271
rect 237 270 238 271
rect 236 270 237 271
rect 235 270 236 271
rect 234 270 235 271
rect 233 270 234 271
rect 232 270 233 271
rect 231 270 232 271
rect 230 270 231 271
rect 229 270 230 271
rect 228 270 229 271
rect 227 270 228 271
rect 226 270 227 271
rect 225 270 226 271
rect 224 270 225 271
rect 223 270 224 271
rect 222 270 223 271
rect 201 270 202 271
rect 200 270 201 271
rect 199 270 200 271
rect 198 270 199 271
rect 197 270 198 271
rect 196 270 197 271
rect 195 270 196 271
rect 194 270 195 271
rect 193 270 194 271
rect 192 270 193 271
rect 191 270 192 271
rect 190 270 191 271
rect 189 270 190 271
rect 188 270 189 271
rect 187 270 188 271
rect 186 270 187 271
rect 185 270 186 271
rect 184 270 185 271
rect 183 270 184 271
rect 182 270 183 271
rect 181 270 182 271
rect 180 270 181 271
rect 179 270 180 271
rect 178 270 179 271
rect 177 270 178 271
rect 176 270 177 271
rect 175 270 176 271
rect 174 270 175 271
rect 173 270 174 271
rect 172 270 173 271
rect 171 270 172 271
rect 170 270 171 271
rect 169 270 170 271
rect 168 270 169 271
rect 167 270 168 271
rect 166 270 167 271
rect 165 270 166 271
rect 164 270 165 271
rect 163 270 164 271
rect 162 270 163 271
rect 161 270 162 271
rect 160 270 161 271
rect 159 270 160 271
rect 158 270 159 271
rect 157 270 158 271
rect 156 270 157 271
rect 155 270 156 271
rect 154 270 155 271
rect 153 270 154 271
rect 152 270 153 271
rect 151 270 152 271
rect 150 270 151 271
rect 149 270 150 271
rect 148 270 149 271
rect 147 270 148 271
rect 146 270 147 271
rect 145 270 146 271
rect 144 270 145 271
rect 143 270 144 271
rect 142 270 143 271
rect 141 270 142 271
rect 140 270 141 271
rect 139 270 140 271
rect 138 270 139 271
rect 137 270 138 271
rect 136 270 137 271
rect 135 270 136 271
rect 134 270 135 271
rect 133 270 134 271
rect 132 270 133 271
rect 131 270 132 271
rect 130 270 131 271
rect 129 270 130 271
rect 128 270 129 271
rect 127 270 128 271
rect 126 270 127 271
rect 125 270 126 271
rect 124 270 125 271
rect 110 270 111 271
rect 109 270 110 271
rect 108 270 109 271
rect 107 270 108 271
rect 106 270 107 271
rect 105 270 106 271
rect 104 270 105 271
rect 103 270 104 271
rect 102 270 103 271
rect 101 270 102 271
rect 100 270 101 271
rect 99 270 100 271
rect 98 270 99 271
rect 97 270 98 271
rect 96 270 97 271
rect 95 270 96 271
rect 94 270 95 271
rect 93 270 94 271
rect 92 270 93 271
rect 91 270 92 271
rect 90 270 91 271
rect 89 270 90 271
rect 88 270 89 271
rect 87 270 88 271
rect 86 270 87 271
rect 85 270 86 271
rect 84 270 85 271
rect 83 270 84 271
rect 82 270 83 271
rect 81 270 82 271
rect 80 270 81 271
rect 79 270 80 271
rect 78 270 79 271
rect 77 270 78 271
rect 76 270 77 271
rect 75 270 76 271
rect 58 270 59 271
rect 57 270 58 271
rect 56 270 57 271
rect 55 270 56 271
rect 54 270 55 271
rect 53 270 54 271
rect 52 270 53 271
rect 51 270 52 271
rect 50 270 51 271
rect 49 270 50 271
rect 48 270 49 271
rect 47 270 48 271
rect 46 270 47 271
rect 45 270 46 271
rect 44 270 45 271
rect 43 270 44 271
rect 42 270 43 271
rect 41 270 42 271
rect 40 270 41 271
rect 39 270 40 271
rect 38 270 39 271
rect 37 270 38 271
rect 36 270 37 271
rect 35 270 36 271
rect 24 270 25 271
rect 23 270 24 271
rect 22 270 23 271
rect 21 270 22 271
rect 20 270 21 271
rect 19 270 20 271
rect 18 270 19 271
rect 17 270 18 271
rect 16 270 17 271
rect 15 270 16 271
rect 14 270 15 271
rect 13 270 14 271
rect 12 270 13 271
rect 11 270 12 271
rect 10 270 11 271
rect 9 270 10 271
rect 8 270 9 271
rect 7 270 8 271
rect 6 270 7 271
rect 5 270 6 271
rect 4 270 5 271
rect 3 270 4 271
rect 2 270 3 271
rect 1 270 2 271
rect 478 271 479 272
rect 477 271 478 272
rect 476 271 477 272
rect 475 271 476 272
rect 474 271 475 272
rect 473 271 474 272
rect 472 271 473 272
rect 471 271 472 272
rect 470 271 471 272
rect 469 271 470 272
rect 468 271 469 272
rect 467 271 468 272
rect 466 271 467 272
rect 465 271 466 272
rect 464 271 465 272
rect 463 271 464 272
rect 462 271 463 272
rect 461 271 462 272
rect 460 271 461 272
rect 459 271 460 272
rect 458 271 459 272
rect 292 271 293 272
rect 291 271 292 272
rect 290 271 291 272
rect 289 271 290 272
rect 288 271 289 272
rect 287 271 288 272
rect 286 271 287 272
rect 285 271 286 272
rect 284 271 285 272
rect 283 271 284 272
rect 282 271 283 272
rect 281 271 282 272
rect 280 271 281 272
rect 279 271 280 272
rect 278 271 279 272
rect 277 271 278 272
rect 276 271 277 272
rect 275 271 276 272
rect 274 271 275 272
rect 273 271 274 272
rect 272 271 273 272
rect 271 271 272 272
rect 270 271 271 272
rect 269 271 270 272
rect 268 271 269 272
rect 267 271 268 272
rect 266 271 267 272
rect 265 271 266 272
rect 264 271 265 272
rect 263 271 264 272
rect 262 271 263 272
rect 261 271 262 272
rect 260 271 261 272
rect 259 271 260 272
rect 258 271 259 272
rect 257 271 258 272
rect 256 271 257 272
rect 255 271 256 272
rect 254 271 255 272
rect 253 271 254 272
rect 252 271 253 272
rect 251 271 252 272
rect 250 271 251 272
rect 249 271 250 272
rect 248 271 249 272
rect 247 271 248 272
rect 246 271 247 272
rect 245 271 246 272
rect 244 271 245 272
rect 243 271 244 272
rect 242 271 243 272
rect 241 271 242 272
rect 240 271 241 272
rect 239 271 240 272
rect 238 271 239 272
rect 237 271 238 272
rect 236 271 237 272
rect 235 271 236 272
rect 234 271 235 272
rect 233 271 234 272
rect 232 271 233 272
rect 231 271 232 272
rect 230 271 231 272
rect 229 271 230 272
rect 228 271 229 272
rect 227 271 228 272
rect 226 271 227 272
rect 225 271 226 272
rect 224 271 225 272
rect 223 271 224 272
rect 222 271 223 272
rect 221 271 222 272
rect 200 271 201 272
rect 199 271 200 272
rect 198 271 199 272
rect 197 271 198 272
rect 196 271 197 272
rect 195 271 196 272
rect 194 271 195 272
rect 193 271 194 272
rect 192 271 193 272
rect 191 271 192 272
rect 190 271 191 272
rect 189 271 190 272
rect 188 271 189 272
rect 187 271 188 272
rect 186 271 187 272
rect 185 271 186 272
rect 184 271 185 272
rect 183 271 184 272
rect 182 271 183 272
rect 181 271 182 272
rect 180 271 181 272
rect 179 271 180 272
rect 178 271 179 272
rect 177 271 178 272
rect 176 271 177 272
rect 175 271 176 272
rect 174 271 175 272
rect 173 271 174 272
rect 172 271 173 272
rect 171 271 172 272
rect 170 271 171 272
rect 169 271 170 272
rect 168 271 169 272
rect 167 271 168 272
rect 166 271 167 272
rect 165 271 166 272
rect 164 271 165 272
rect 163 271 164 272
rect 162 271 163 272
rect 161 271 162 272
rect 160 271 161 272
rect 159 271 160 272
rect 158 271 159 272
rect 157 271 158 272
rect 156 271 157 272
rect 155 271 156 272
rect 154 271 155 272
rect 153 271 154 272
rect 152 271 153 272
rect 151 271 152 272
rect 150 271 151 272
rect 149 271 150 272
rect 148 271 149 272
rect 147 271 148 272
rect 146 271 147 272
rect 145 271 146 272
rect 144 271 145 272
rect 143 271 144 272
rect 142 271 143 272
rect 141 271 142 272
rect 140 271 141 272
rect 139 271 140 272
rect 138 271 139 272
rect 137 271 138 272
rect 136 271 137 272
rect 135 271 136 272
rect 134 271 135 272
rect 133 271 134 272
rect 132 271 133 272
rect 131 271 132 272
rect 130 271 131 272
rect 129 271 130 272
rect 128 271 129 272
rect 127 271 128 272
rect 126 271 127 272
rect 125 271 126 272
rect 124 271 125 272
rect 110 271 111 272
rect 109 271 110 272
rect 108 271 109 272
rect 107 271 108 272
rect 106 271 107 272
rect 105 271 106 272
rect 104 271 105 272
rect 103 271 104 272
rect 102 271 103 272
rect 101 271 102 272
rect 100 271 101 272
rect 99 271 100 272
rect 98 271 99 272
rect 97 271 98 272
rect 96 271 97 272
rect 95 271 96 272
rect 94 271 95 272
rect 93 271 94 272
rect 92 271 93 272
rect 91 271 92 272
rect 90 271 91 272
rect 89 271 90 272
rect 88 271 89 272
rect 87 271 88 272
rect 86 271 87 272
rect 85 271 86 272
rect 84 271 85 272
rect 83 271 84 272
rect 82 271 83 272
rect 81 271 82 272
rect 80 271 81 272
rect 79 271 80 272
rect 78 271 79 272
rect 77 271 78 272
rect 76 271 77 272
rect 59 271 60 272
rect 58 271 59 272
rect 57 271 58 272
rect 56 271 57 272
rect 55 271 56 272
rect 54 271 55 272
rect 53 271 54 272
rect 52 271 53 272
rect 51 271 52 272
rect 50 271 51 272
rect 49 271 50 272
rect 48 271 49 272
rect 47 271 48 272
rect 46 271 47 272
rect 45 271 46 272
rect 44 271 45 272
rect 43 271 44 272
rect 42 271 43 272
rect 41 271 42 272
rect 40 271 41 272
rect 39 271 40 272
rect 38 271 39 272
rect 37 271 38 272
rect 36 271 37 272
rect 35 271 36 272
rect 24 271 25 272
rect 23 271 24 272
rect 22 271 23 272
rect 21 271 22 272
rect 20 271 21 272
rect 19 271 20 272
rect 18 271 19 272
rect 17 271 18 272
rect 16 271 17 272
rect 15 271 16 272
rect 14 271 15 272
rect 13 271 14 272
rect 12 271 13 272
rect 11 271 12 272
rect 10 271 11 272
rect 9 271 10 272
rect 8 271 9 272
rect 7 271 8 272
rect 6 271 7 272
rect 5 271 6 272
rect 4 271 5 272
rect 3 271 4 272
rect 2 271 3 272
rect 1 271 2 272
rect 478 272 479 273
rect 458 272 459 273
rect 437 272 438 273
rect 436 272 437 273
rect 395 272 396 273
rect 394 272 395 273
rect 393 272 394 273
rect 292 272 293 273
rect 291 272 292 273
rect 290 272 291 273
rect 289 272 290 273
rect 288 272 289 273
rect 287 272 288 273
rect 286 272 287 273
rect 285 272 286 273
rect 284 272 285 273
rect 283 272 284 273
rect 282 272 283 273
rect 281 272 282 273
rect 280 272 281 273
rect 279 272 280 273
rect 278 272 279 273
rect 277 272 278 273
rect 276 272 277 273
rect 275 272 276 273
rect 274 272 275 273
rect 273 272 274 273
rect 272 272 273 273
rect 271 272 272 273
rect 270 272 271 273
rect 269 272 270 273
rect 268 272 269 273
rect 267 272 268 273
rect 266 272 267 273
rect 265 272 266 273
rect 264 272 265 273
rect 263 272 264 273
rect 262 272 263 273
rect 261 272 262 273
rect 260 272 261 273
rect 259 272 260 273
rect 258 272 259 273
rect 257 272 258 273
rect 256 272 257 273
rect 255 272 256 273
rect 254 272 255 273
rect 253 272 254 273
rect 252 272 253 273
rect 251 272 252 273
rect 250 272 251 273
rect 249 272 250 273
rect 248 272 249 273
rect 247 272 248 273
rect 246 272 247 273
rect 245 272 246 273
rect 244 272 245 273
rect 243 272 244 273
rect 242 272 243 273
rect 241 272 242 273
rect 240 272 241 273
rect 239 272 240 273
rect 238 272 239 273
rect 237 272 238 273
rect 236 272 237 273
rect 235 272 236 273
rect 234 272 235 273
rect 233 272 234 273
rect 232 272 233 273
rect 231 272 232 273
rect 230 272 231 273
rect 229 272 230 273
rect 228 272 229 273
rect 227 272 228 273
rect 226 272 227 273
rect 225 272 226 273
rect 224 272 225 273
rect 223 272 224 273
rect 222 272 223 273
rect 221 272 222 273
rect 200 272 201 273
rect 199 272 200 273
rect 198 272 199 273
rect 197 272 198 273
rect 196 272 197 273
rect 195 272 196 273
rect 194 272 195 273
rect 193 272 194 273
rect 192 272 193 273
rect 191 272 192 273
rect 190 272 191 273
rect 189 272 190 273
rect 188 272 189 273
rect 187 272 188 273
rect 186 272 187 273
rect 185 272 186 273
rect 184 272 185 273
rect 183 272 184 273
rect 182 272 183 273
rect 181 272 182 273
rect 180 272 181 273
rect 179 272 180 273
rect 178 272 179 273
rect 177 272 178 273
rect 176 272 177 273
rect 175 272 176 273
rect 174 272 175 273
rect 173 272 174 273
rect 172 272 173 273
rect 171 272 172 273
rect 170 272 171 273
rect 169 272 170 273
rect 168 272 169 273
rect 167 272 168 273
rect 166 272 167 273
rect 165 272 166 273
rect 164 272 165 273
rect 163 272 164 273
rect 162 272 163 273
rect 161 272 162 273
rect 160 272 161 273
rect 159 272 160 273
rect 158 272 159 273
rect 157 272 158 273
rect 156 272 157 273
rect 155 272 156 273
rect 154 272 155 273
rect 153 272 154 273
rect 152 272 153 273
rect 151 272 152 273
rect 150 272 151 273
rect 149 272 150 273
rect 148 272 149 273
rect 147 272 148 273
rect 146 272 147 273
rect 145 272 146 273
rect 144 272 145 273
rect 143 272 144 273
rect 142 272 143 273
rect 141 272 142 273
rect 140 272 141 273
rect 139 272 140 273
rect 138 272 139 273
rect 137 272 138 273
rect 136 272 137 273
rect 135 272 136 273
rect 134 272 135 273
rect 133 272 134 273
rect 132 272 133 273
rect 131 272 132 273
rect 130 272 131 273
rect 129 272 130 273
rect 128 272 129 273
rect 127 272 128 273
rect 126 272 127 273
rect 125 272 126 273
rect 110 272 111 273
rect 109 272 110 273
rect 108 272 109 273
rect 107 272 108 273
rect 106 272 107 273
rect 105 272 106 273
rect 104 272 105 273
rect 103 272 104 273
rect 102 272 103 273
rect 101 272 102 273
rect 100 272 101 273
rect 99 272 100 273
rect 98 272 99 273
rect 97 272 98 273
rect 96 272 97 273
rect 95 272 96 273
rect 94 272 95 273
rect 93 272 94 273
rect 92 272 93 273
rect 91 272 92 273
rect 90 272 91 273
rect 89 272 90 273
rect 88 272 89 273
rect 87 272 88 273
rect 86 272 87 273
rect 85 272 86 273
rect 84 272 85 273
rect 83 272 84 273
rect 82 272 83 273
rect 81 272 82 273
rect 80 272 81 273
rect 79 272 80 273
rect 78 272 79 273
rect 77 272 78 273
rect 76 272 77 273
rect 59 272 60 273
rect 58 272 59 273
rect 57 272 58 273
rect 56 272 57 273
rect 55 272 56 273
rect 54 272 55 273
rect 53 272 54 273
rect 52 272 53 273
rect 51 272 52 273
rect 50 272 51 273
rect 49 272 50 273
rect 48 272 49 273
rect 47 272 48 273
rect 46 272 47 273
rect 45 272 46 273
rect 44 272 45 273
rect 43 272 44 273
rect 42 272 43 273
rect 41 272 42 273
rect 40 272 41 273
rect 39 272 40 273
rect 38 272 39 273
rect 37 272 38 273
rect 36 272 37 273
rect 35 272 36 273
rect 24 272 25 273
rect 23 272 24 273
rect 22 272 23 273
rect 21 272 22 273
rect 20 272 21 273
rect 19 272 20 273
rect 18 272 19 273
rect 17 272 18 273
rect 16 272 17 273
rect 15 272 16 273
rect 14 272 15 273
rect 13 272 14 273
rect 12 272 13 273
rect 11 272 12 273
rect 10 272 11 273
rect 9 272 10 273
rect 8 272 9 273
rect 7 272 8 273
rect 6 272 7 273
rect 5 272 6 273
rect 4 272 5 273
rect 3 272 4 273
rect 2 272 3 273
rect 1 272 2 273
rect 478 273 479 274
rect 458 273 459 274
rect 437 273 438 274
rect 436 273 437 274
rect 435 273 436 274
rect 395 273 396 274
rect 394 273 395 274
rect 393 273 394 274
rect 291 273 292 274
rect 290 273 291 274
rect 289 273 290 274
rect 288 273 289 274
rect 287 273 288 274
rect 286 273 287 274
rect 285 273 286 274
rect 284 273 285 274
rect 283 273 284 274
rect 282 273 283 274
rect 281 273 282 274
rect 280 273 281 274
rect 279 273 280 274
rect 278 273 279 274
rect 277 273 278 274
rect 276 273 277 274
rect 275 273 276 274
rect 274 273 275 274
rect 273 273 274 274
rect 272 273 273 274
rect 271 273 272 274
rect 270 273 271 274
rect 269 273 270 274
rect 268 273 269 274
rect 267 273 268 274
rect 266 273 267 274
rect 265 273 266 274
rect 264 273 265 274
rect 263 273 264 274
rect 262 273 263 274
rect 261 273 262 274
rect 260 273 261 274
rect 259 273 260 274
rect 258 273 259 274
rect 257 273 258 274
rect 256 273 257 274
rect 255 273 256 274
rect 254 273 255 274
rect 253 273 254 274
rect 252 273 253 274
rect 251 273 252 274
rect 250 273 251 274
rect 249 273 250 274
rect 248 273 249 274
rect 247 273 248 274
rect 246 273 247 274
rect 245 273 246 274
rect 244 273 245 274
rect 243 273 244 274
rect 242 273 243 274
rect 241 273 242 274
rect 240 273 241 274
rect 239 273 240 274
rect 238 273 239 274
rect 237 273 238 274
rect 236 273 237 274
rect 235 273 236 274
rect 234 273 235 274
rect 233 273 234 274
rect 232 273 233 274
rect 231 273 232 274
rect 230 273 231 274
rect 229 273 230 274
rect 228 273 229 274
rect 227 273 228 274
rect 226 273 227 274
rect 225 273 226 274
rect 224 273 225 274
rect 223 273 224 274
rect 222 273 223 274
rect 221 273 222 274
rect 220 273 221 274
rect 199 273 200 274
rect 198 273 199 274
rect 197 273 198 274
rect 196 273 197 274
rect 195 273 196 274
rect 194 273 195 274
rect 193 273 194 274
rect 192 273 193 274
rect 191 273 192 274
rect 190 273 191 274
rect 189 273 190 274
rect 188 273 189 274
rect 187 273 188 274
rect 186 273 187 274
rect 185 273 186 274
rect 184 273 185 274
rect 183 273 184 274
rect 182 273 183 274
rect 181 273 182 274
rect 180 273 181 274
rect 179 273 180 274
rect 178 273 179 274
rect 177 273 178 274
rect 176 273 177 274
rect 175 273 176 274
rect 174 273 175 274
rect 173 273 174 274
rect 172 273 173 274
rect 171 273 172 274
rect 170 273 171 274
rect 169 273 170 274
rect 168 273 169 274
rect 167 273 168 274
rect 166 273 167 274
rect 165 273 166 274
rect 164 273 165 274
rect 163 273 164 274
rect 162 273 163 274
rect 161 273 162 274
rect 160 273 161 274
rect 159 273 160 274
rect 158 273 159 274
rect 157 273 158 274
rect 156 273 157 274
rect 155 273 156 274
rect 154 273 155 274
rect 153 273 154 274
rect 152 273 153 274
rect 151 273 152 274
rect 150 273 151 274
rect 149 273 150 274
rect 148 273 149 274
rect 147 273 148 274
rect 146 273 147 274
rect 145 273 146 274
rect 144 273 145 274
rect 143 273 144 274
rect 142 273 143 274
rect 141 273 142 274
rect 140 273 141 274
rect 139 273 140 274
rect 138 273 139 274
rect 137 273 138 274
rect 136 273 137 274
rect 135 273 136 274
rect 134 273 135 274
rect 133 273 134 274
rect 132 273 133 274
rect 131 273 132 274
rect 130 273 131 274
rect 129 273 130 274
rect 128 273 129 274
rect 127 273 128 274
rect 126 273 127 274
rect 125 273 126 274
rect 110 273 111 274
rect 109 273 110 274
rect 108 273 109 274
rect 107 273 108 274
rect 106 273 107 274
rect 105 273 106 274
rect 104 273 105 274
rect 103 273 104 274
rect 102 273 103 274
rect 101 273 102 274
rect 100 273 101 274
rect 99 273 100 274
rect 98 273 99 274
rect 97 273 98 274
rect 96 273 97 274
rect 95 273 96 274
rect 94 273 95 274
rect 93 273 94 274
rect 92 273 93 274
rect 91 273 92 274
rect 90 273 91 274
rect 89 273 90 274
rect 88 273 89 274
rect 87 273 88 274
rect 86 273 87 274
rect 85 273 86 274
rect 84 273 85 274
rect 83 273 84 274
rect 82 273 83 274
rect 81 273 82 274
rect 80 273 81 274
rect 79 273 80 274
rect 78 273 79 274
rect 77 273 78 274
rect 60 273 61 274
rect 59 273 60 274
rect 58 273 59 274
rect 57 273 58 274
rect 56 273 57 274
rect 55 273 56 274
rect 54 273 55 274
rect 53 273 54 274
rect 52 273 53 274
rect 51 273 52 274
rect 50 273 51 274
rect 49 273 50 274
rect 48 273 49 274
rect 47 273 48 274
rect 46 273 47 274
rect 45 273 46 274
rect 44 273 45 274
rect 43 273 44 274
rect 42 273 43 274
rect 41 273 42 274
rect 40 273 41 274
rect 39 273 40 274
rect 38 273 39 274
rect 37 273 38 274
rect 36 273 37 274
rect 25 273 26 274
rect 24 273 25 274
rect 23 273 24 274
rect 22 273 23 274
rect 21 273 22 274
rect 20 273 21 274
rect 19 273 20 274
rect 18 273 19 274
rect 17 273 18 274
rect 16 273 17 274
rect 15 273 16 274
rect 14 273 15 274
rect 13 273 14 274
rect 12 273 13 274
rect 11 273 12 274
rect 10 273 11 274
rect 9 273 10 274
rect 8 273 9 274
rect 7 273 8 274
rect 6 273 7 274
rect 5 273 6 274
rect 4 273 5 274
rect 3 273 4 274
rect 2 273 3 274
rect 1 273 2 274
rect 437 274 438 275
rect 436 274 437 275
rect 435 274 436 275
rect 395 274 396 275
rect 394 274 395 275
rect 393 274 394 275
rect 290 274 291 275
rect 289 274 290 275
rect 288 274 289 275
rect 287 274 288 275
rect 286 274 287 275
rect 285 274 286 275
rect 284 274 285 275
rect 283 274 284 275
rect 282 274 283 275
rect 281 274 282 275
rect 280 274 281 275
rect 279 274 280 275
rect 278 274 279 275
rect 277 274 278 275
rect 276 274 277 275
rect 275 274 276 275
rect 274 274 275 275
rect 273 274 274 275
rect 272 274 273 275
rect 271 274 272 275
rect 270 274 271 275
rect 269 274 270 275
rect 268 274 269 275
rect 267 274 268 275
rect 266 274 267 275
rect 265 274 266 275
rect 264 274 265 275
rect 263 274 264 275
rect 262 274 263 275
rect 261 274 262 275
rect 260 274 261 275
rect 259 274 260 275
rect 258 274 259 275
rect 257 274 258 275
rect 256 274 257 275
rect 255 274 256 275
rect 254 274 255 275
rect 253 274 254 275
rect 252 274 253 275
rect 251 274 252 275
rect 250 274 251 275
rect 249 274 250 275
rect 248 274 249 275
rect 247 274 248 275
rect 246 274 247 275
rect 245 274 246 275
rect 244 274 245 275
rect 243 274 244 275
rect 242 274 243 275
rect 241 274 242 275
rect 240 274 241 275
rect 239 274 240 275
rect 238 274 239 275
rect 237 274 238 275
rect 236 274 237 275
rect 235 274 236 275
rect 234 274 235 275
rect 233 274 234 275
rect 232 274 233 275
rect 231 274 232 275
rect 230 274 231 275
rect 229 274 230 275
rect 228 274 229 275
rect 227 274 228 275
rect 226 274 227 275
rect 225 274 226 275
rect 224 274 225 275
rect 223 274 224 275
rect 222 274 223 275
rect 221 274 222 275
rect 220 274 221 275
rect 199 274 200 275
rect 198 274 199 275
rect 197 274 198 275
rect 196 274 197 275
rect 195 274 196 275
rect 194 274 195 275
rect 193 274 194 275
rect 192 274 193 275
rect 191 274 192 275
rect 190 274 191 275
rect 189 274 190 275
rect 188 274 189 275
rect 187 274 188 275
rect 186 274 187 275
rect 185 274 186 275
rect 184 274 185 275
rect 183 274 184 275
rect 182 274 183 275
rect 181 274 182 275
rect 180 274 181 275
rect 179 274 180 275
rect 178 274 179 275
rect 177 274 178 275
rect 176 274 177 275
rect 175 274 176 275
rect 174 274 175 275
rect 173 274 174 275
rect 172 274 173 275
rect 171 274 172 275
rect 170 274 171 275
rect 169 274 170 275
rect 168 274 169 275
rect 167 274 168 275
rect 166 274 167 275
rect 165 274 166 275
rect 164 274 165 275
rect 163 274 164 275
rect 162 274 163 275
rect 161 274 162 275
rect 160 274 161 275
rect 159 274 160 275
rect 158 274 159 275
rect 157 274 158 275
rect 156 274 157 275
rect 155 274 156 275
rect 154 274 155 275
rect 153 274 154 275
rect 152 274 153 275
rect 151 274 152 275
rect 150 274 151 275
rect 149 274 150 275
rect 148 274 149 275
rect 147 274 148 275
rect 146 274 147 275
rect 145 274 146 275
rect 144 274 145 275
rect 143 274 144 275
rect 142 274 143 275
rect 141 274 142 275
rect 140 274 141 275
rect 139 274 140 275
rect 138 274 139 275
rect 137 274 138 275
rect 136 274 137 275
rect 135 274 136 275
rect 134 274 135 275
rect 133 274 134 275
rect 132 274 133 275
rect 131 274 132 275
rect 130 274 131 275
rect 129 274 130 275
rect 128 274 129 275
rect 127 274 128 275
rect 126 274 127 275
rect 125 274 126 275
rect 111 274 112 275
rect 110 274 111 275
rect 109 274 110 275
rect 108 274 109 275
rect 107 274 108 275
rect 106 274 107 275
rect 105 274 106 275
rect 104 274 105 275
rect 103 274 104 275
rect 102 274 103 275
rect 101 274 102 275
rect 100 274 101 275
rect 99 274 100 275
rect 98 274 99 275
rect 97 274 98 275
rect 96 274 97 275
rect 95 274 96 275
rect 94 274 95 275
rect 93 274 94 275
rect 92 274 93 275
rect 91 274 92 275
rect 90 274 91 275
rect 89 274 90 275
rect 88 274 89 275
rect 87 274 88 275
rect 86 274 87 275
rect 85 274 86 275
rect 84 274 85 275
rect 83 274 84 275
rect 82 274 83 275
rect 81 274 82 275
rect 80 274 81 275
rect 79 274 80 275
rect 78 274 79 275
rect 77 274 78 275
rect 60 274 61 275
rect 59 274 60 275
rect 58 274 59 275
rect 57 274 58 275
rect 56 274 57 275
rect 55 274 56 275
rect 54 274 55 275
rect 53 274 54 275
rect 52 274 53 275
rect 51 274 52 275
rect 50 274 51 275
rect 49 274 50 275
rect 48 274 49 275
rect 47 274 48 275
rect 46 274 47 275
rect 45 274 46 275
rect 44 274 45 275
rect 43 274 44 275
rect 42 274 43 275
rect 41 274 42 275
rect 40 274 41 275
rect 39 274 40 275
rect 38 274 39 275
rect 37 274 38 275
rect 36 274 37 275
rect 25 274 26 275
rect 24 274 25 275
rect 23 274 24 275
rect 22 274 23 275
rect 21 274 22 275
rect 20 274 21 275
rect 19 274 20 275
rect 18 274 19 275
rect 17 274 18 275
rect 16 274 17 275
rect 15 274 16 275
rect 14 274 15 275
rect 13 274 14 275
rect 12 274 13 275
rect 11 274 12 275
rect 10 274 11 275
rect 9 274 10 275
rect 8 274 9 275
rect 7 274 8 275
rect 6 274 7 275
rect 5 274 6 275
rect 4 274 5 275
rect 3 274 4 275
rect 2 274 3 275
rect 1 274 2 275
rect 437 275 438 276
rect 436 275 437 276
rect 435 275 436 276
rect 395 275 396 276
rect 394 275 395 276
rect 393 275 394 276
rect 289 275 290 276
rect 288 275 289 276
rect 287 275 288 276
rect 286 275 287 276
rect 285 275 286 276
rect 284 275 285 276
rect 283 275 284 276
rect 282 275 283 276
rect 281 275 282 276
rect 280 275 281 276
rect 279 275 280 276
rect 278 275 279 276
rect 277 275 278 276
rect 276 275 277 276
rect 275 275 276 276
rect 274 275 275 276
rect 273 275 274 276
rect 272 275 273 276
rect 271 275 272 276
rect 270 275 271 276
rect 269 275 270 276
rect 268 275 269 276
rect 267 275 268 276
rect 266 275 267 276
rect 265 275 266 276
rect 264 275 265 276
rect 263 275 264 276
rect 262 275 263 276
rect 261 275 262 276
rect 260 275 261 276
rect 259 275 260 276
rect 258 275 259 276
rect 257 275 258 276
rect 256 275 257 276
rect 255 275 256 276
rect 254 275 255 276
rect 253 275 254 276
rect 252 275 253 276
rect 251 275 252 276
rect 250 275 251 276
rect 249 275 250 276
rect 248 275 249 276
rect 247 275 248 276
rect 246 275 247 276
rect 245 275 246 276
rect 244 275 245 276
rect 243 275 244 276
rect 242 275 243 276
rect 241 275 242 276
rect 240 275 241 276
rect 239 275 240 276
rect 238 275 239 276
rect 237 275 238 276
rect 236 275 237 276
rect 235 275 236 276
rect 234 275 235 276
rect 233 275 234 276
rect 232 275 233 276
rect 231 275 232 276
rect 230 275 231 276
rect 229 275 230 276
rect 228 275 229 276
rect 227 275 228 276
rect 226 275 227 276
rect 225 275 226 276
rect 224 275 225 276
rect 223 275 224 276
rect 222 275 223 276
rect 221 275 222 276
rect 220 275 221 276
rect 198 275 199 276
rect 197 275 198 276
rect 196 275 197 276
rect 195 275 196 276
rect 194 275 195 276
rect 193 275 194 276
rect 192 275 193 276
rect 191 275 192 276
rect 190 275 191 276
rect 189 275 190 276
rect 188 275 189 276
rect 187 275 188 276
rect 186 275 187 276
rect 185 275 186 276
rect 184 275 185 276
rect 183 275 184 276
rect 182 275 183 276
rect 181 275 182 276
rect 180 275 181 276
rect 179 275 180 276
rect 178 275 179 276
rect 177 275 178 276
rect 176 275 177 276
rect 175 275 176 276
rect 174 275 175 276
rect 173 275 174 276
rect 172 275 173 276
rect 171 275 172 276
rect 170 275 171 276
rect 169 275 170 276
rect 168 275 169 276
rect 167 275 168 276
rect 166 275 167 276
rect 165 275 166 276
rect 164 275 165 276
rect 163 275 164 276
rect 162 275 163 276
rect 161 275 162 276
rect 160 275 161 276
rect 159 275 160 276
rect 158 275 159 276
rect 157 275 158 276
rect 156 275 157 276
rect 155 275 156 276
rect 154 275 155 276
rect 153 275 154 276
rect 152 275 153 276
rect 151 275 152 276
rect 150 275 151 276
rect 149 275 150 276
rect 148 275 149 276
rect 147 275 148 276
rect 146 275 147 276
rect 145 275 146 276
rect 144 275 145 276
rect 143 275 144 276
rect 142 275 143 276
rect 141 275 142 276
rect 140 275 141 276
rect 139 275 140 276
rect 138 275 139 276
rect 137 275 138 276
rect 136 275 137 276
rect 135 275 136 276
rect 134 275 135 276
rect 133 275 134 276
rect 132 275 133 276
rect 131 275 132 276
rect 130 275 131 276
rect 129 275 130 276
rect 128 275 129 276
rect 127 275 128 276
rect 126 275 127 276
rect 111 275 112 276
rect 110 275 111 276
rect 109 275 110 276
rect 108 275 109 276
rect 107 275 108 276
rect 106 275 107 276
rect 105 275 106 276
rect 104 275 105 276
rect 103 275 104 276
rect 102 275 103 276
rect 101 275 102 276
rect 100 275 101 276
rect 99 275 100 276
rect 98 275 99 276
rect 97 275 98 276
rect 96 275 97 276
rect 95 275 96 276
rect 94 275 95 276
rect 93 275 94 276
rect 92 275 93 276
rect 91 275 92 276
rect 90 275 91 276
rect 89 275 90 276
rect 88 275 89 276
rect 87 275 88 276
rect 86 275 87 276
rect 85 275 86 276
rect 84 275 85 276
rect 83 275 84 276
rect 82 275 83 276
rect 81 275 82 276
rect 80 275 81 276
rect 79 275 80 276
rect 78 275 79 276
rect 77 275 78 276
rect 60 275 61 276
rect 59 275 60 276
rect 58 275 59 276
rect 57 275 58 276
rect 56 275 57 276
rect 55 275 56 276
rect 54 275 55 276
rect 53 275 54 276
rect 52 275 53 276
rect 51 275 52 276
rect 50 275 51 276
rect 49 275 50 276
rect 48 275 49 276
rect 47 275 48 276
rect 46 275 47 276
rect 45 275 46 276
rect 44 275 45 276
rect 43 275 44 276
rect 42 275 43 276
rect 41 275 42 276
rect 40 275 41 276
rect 39 275 40 276
rect 38 275 39 276
rect 37 275 38 276
rect 36 275 37 276
rect 25 275 26 276
rect 24 275 25 276
rect 23 275 24 276
rect 22 275 23 276
rect 21 275 22 276
rect 20 275 21 276
rect 19 275 20 276
rect 18 275 19 276
rect 17 275 18 276
rect 16 275 17 276
rect 15 275 16 276
rect 14 275 15 276
rect 13 275 14 276
rect 12 275 13 276
rect 11 275 12 276
rect 10 275 11 276
rect 9 275 10 276
rect 8 275 9 276
rect 7 275 8 276
rect 6 275 7 276
rect 5 275 6 276
rect 4 275 5 276
rect 3 275 4 276
rect 2 275 3 276
rect 1 275 2 276
rect 437 276 438 277
rect 436 276 437 277
rect 435 276 436 277
rect 396 276 397 277
rect 395 276 396 277
rect 394 276 395 277
rect 393 276 394 277
rect 288 276 289 277
rect 287 276 288 277
rect 286 276 287 277
rect 285 276 286 277
rect 284 276 285 277
rect 283 276 284 277
rect 282 276 283 277
rect 281 276 282 277
rect 280 276 281 277
rect 279 276 280 277
rect 278 276 279 277
rect 277 276 278 277
rect 276 276 277 277
rect 275 276 276 277
rect 274 276 275 277
rect 273 276 274 277
rect 272 276 273 277
rect 271 276 272 277
rect 270 276 271 277
rect 269 276 270 277
rect 268 276 269 277
rect 267 276 268 277
rect 266 276 267 277
rect 265 276 266 277
rect 264 276 265 277
rect 263 276 264 277
rect 262 276 263 277
rect 261 276 262 277
rect 260 276 261 277
rect 259 276 260 277
rect 258 276 259 277
rect 257 276 258 277
rect 256 276 257 277
rect 255 276 256 277
rect 254 276 255 277
rect 253 276 254 277
rect 252 276 253 277
rect 251 276 252 277
rect 250 276 251 277
rect 249 276 250 277
rect 248 276 249 277
rect 247 276 248 277
rect 246 276 247 277
rect 245 276 246 277
rect 244 276 245 277
rect 243 276 244 277
rect 242 276 243 277
rect 241 276 242 277
rect 240 276 241 277
rect 239 276 240 277
rect 238 276 239 277
rect 237 276 238 277
rect 236 276 237 277
rect 235 276 236 277
rect 234 276 235 277
rect 233 276 234 277
rect 232 276 233 277
rect 231 276 232 277
rect 230 276 231 277
rect 229 276 230 277
rect 228 276 229 277
rect 227 276 228 277
rect 226 276 227 277
rect 225 276 226 277
rect 224 276 225 277
rect 223 276 224 277
rect 222 276 223 277
rect 221 276 222 277
rect 220 276 221 277
rect 219 276 220 277
rect 197 276 198 277
rect 196 276 197 277
rect 195 276 196 277
rect 194 276 195 277
rect 193 276 194 277
rect 192 276 193 277
rect 191 276 192 277
rect 190 276 191 277
rect 189 276 190 277
rect 188 276 189 277
rect 187 276 188 277
rect 186 276 187 277
rect 185 276 186 277
rect 184 276 185 277
rect 183 276 184 277
rect 182 276 183 277
rect 181 276 182 277
rect 180 276 181 277
rect 179 276 180 277
rect 178 276 179 277
rect 177 276 178 277
rect 176 276 177 277
rect 175 276 176 277
rect 174 276 175 277
rect 173 276 174 277
rect 172 276 173 277
rect 171 276 172 277
rect 170 276 171 277
rect 169 276 170 277
rect 168 276 169 277
rect 167 276 168 277
rect 166 276 167 277
rect 165 276 166 277
rect 164 276 165 277
rect 163 276 164 277
rect 162 276 163 277
rect 161 276 162 277
rect 160 276 161 277
rect 159 276 160 277
rect 158 276 159 277
rect 157 276 158 277
rect 156 276 157 277
rect 155 276 156 277
rect 154 276 155 277
rect 153 276 154 277
rect 152 276 153 277
rect 151 276 152 277
rect 150 276 151 277
rect 149 276 150 277
rect 148 276 149 277
rect 147 276 148 277
rect 146 276 147 277
rect 145 276 146 277
rect 144 276 145 277
rect 143 276 144 277
rect 142 276 143 277
rect 141 276 142 277
rect 140 276 141 277
rect 139 276 140 277
rect 138 276 139 277
rect 137 276 138 277
rect 136 276 137 277
rect 135 276 136 277
rect 134 276 135 277
rect 133 276 134 277
rect 132 276 133 277
rect 131 276 132 277
rect 130 276 131 277
rect 129 276 130 277
rect 128 276 129 277
rect 127 276 128 277
rect 126 276 127 277
rect 111 276 112 277
rect 110 276 111 277
rect 109 276 110 277
rect 108 276 109 277
rect 107 276 108 277
rect 106 276 107 277
rect 105 276 106 277
rect 104 276 105 277
rect 103 276 104 277
rect 102 276 103 277
rect 101 276 102 277
rect 100 276 101 277
rect 99 276 100 277
rect 98 276 99 277
rect 97 276 98 277
rect 96 276 97 277
rect 95 276 96 277
rect 94 276 95 277
rect 93 276 94 277
rect 92 276 93 277
rect 91 276 92 277
rect 90 276 91 277
rect 89 276 90 277
rect 88 276 89 277
rect 87 276 88 277
rect 86 276 87 277
rect 85 276 86 277
rect 84 276 85 277
rect 83 276 84 277
rect 82 276 83 277
rect 81 276 82 277
rect 80 276 81 277
rect 79 276 80 277
rect 78 276 79 277
rect 61 276 62 277
rect 60 276 61 277
rect 59 276 60 277
rect 58 276 59 277
rect 57 276 58 277
rect 56 276 57 277
rect 55 276 56 277
rect 54 276 55 277
rect 53 276 54 277
rect 52 276 53 277
rect 51 276 52 277
rect 50 276 51 277
rect 49 276 50 277
rect 48 276 49 277
rect 47 276 48 277
rect 46 276 47 277
rect 45 276 46 277
rect 44 276 45 277
rect 43 276 44 277
rect 42 276 43 277
rect 41 276 42 277
rect 40 276 41 277
rect 39 276 40 277
rect 38 276 39 277
rect 37 276 38 277
rect 36 276 37 277
rect 25 276 26 277
rect 24 276 25 277
rect 23 276 24 277
rect 22 276 23 277
rect 21 276 22 277
rect 20 276 21 277
rect 19 276 20 277
rect 18 276 19 277
rect 17 276 18 277
rect 16 276 17 277
rect 15 276 16 277
rect 14 276 15 277
rect 13 276 14 277
rect 12 276 13 277
rect 11 276 12 277
rect 10 276 11 277
rect 9 276 10 277
rect 8 276 9 277
rect 7 276 8 277
rect 6 276 7 277
rect 5 276 6 277
rect 4 276 5 277
rect 3 276 4 277
rect 2 276 3 277
rect 1 276 2 277
rect 437 277 438 278
rect 436 277 437 278
rect 435 277 436 278
rect 434 277 435 278
rect 433 277 434 278
rect 397 277 398 278
rect 396 277 397 278
rect 395 277 396 278
rect 394 277 395 278
rect 393 277 394 278
rect 288 277 289 278
rect 287 277 288 278
rect 286 277 287 278
rect 285 277 286 278
rect 284 277 285 278
rect 283 277 284 278
rect 282 277 283 278
rect 281 277 282 278
rect 280 277 281 278
rect 279 277 280 278
rect 278 277 279 278
rect 277 277 278 278
rect 276 277 277 278
rect 275 277 276 278
rect 274 277 275 278
rect 273 277 274 278
rect 272 277 273 278
rect 271 277 272 278
rect 270 277 271 278
rect 269 277 270 278
rect 268 277 269 278
rect 267 277 268 278
rect 266 277 267 278
rect 265 277 266 278
rect 264 277 265 278
rect 263 277 264 278
rect 262 277 263 278
rect 261 277 262 278
rect 260 277 261 278
rect 259 277 260 278
rect 258 277 259 278
rect 257 277 258 278
rect 256 277 257 278
rect 255 277 256 278
rect 254 277 255 278
rect 253 277 254 278
rect 252 277 253 278
rect 251 277 252 278
rect 250 277 251 278
rect 249 277 250 278
rect 248 277 249 278
rect 247 277 248 278
rect 246 277 247 278
rect 245 277 246 278
rect 244 277 245 278
rect 243 277 244 278
rect 242 277 243 278
rect 241 277 242 278
rect 240 277 241 278
rect 239 277 240 278
rect 238 277 239 278
rect 237 277 238 278
rect 236 277 237 278
rect 235 277 236 278
rect 234 277 235 278
rect 233 277 234 278
rect 232 277 233 278
rect 231 277 232 278
rect 230 277 231 278
rect 229 277 230 278
rect 228 277 229 278
rect 227 277 228 278
rect 226 277 227 278
rect 225 277 226 278
rect 224 277 225 278
rect 223 277 224 278
rect 222 277 223 278
rect 221 277 222 278
rect 220 277 221 278
rect 219 277 220 278
rect 197 277 198 278
rect 196 277 197 278
rect 195 277 196 278
rect 194 277 195 278
rect 193 277 194 278
rect 192 277 193 278
rect 191 277 192 278
rect 190 277 191 278
rect 189 277 190 278
rect 188 277 189 278
rect 187 277 188 278
rect 186 277 187 278
rect 185 277 186 278
rect 184 277 185 278
rect 183 277 184 278
rect 182 277 183 278
rect 181 277 182 278
rect 180 277 181 278
rect 179 277 180 278
rect 178 277 179 278
rect 177 277 178 278
rect 176 277 177 278
rect 175 277 176 278
rect 174 277 175 278
rect 173 277 174 278
rect 172 277 173 278
rect 171 277 172 278
rect 170 277 171 278
rect 169 277 170 278
rect 168 277 169 278
rect 167 277 168 278
rect 166 277 167 278
rect 165 277 166 278
rect 164 277 165 278
rect 163 277 164 278
rect 162 277 163 278
rect 161 277 162 278
rect 160 277 161 278
rect 159 277 160 278
rect 158 277 159 278
rect 157 277 158 278
rect 156 277 157 278
rect 155 277 156 278
rect 154 277 155 278
rect 153 277 154 278
rect 152 277 153 278
rect 151 277 152 278
rect 150 277 151 278
rect 149 277 150 278
rect 148 277 149 278
rect 147 277 148 278
rect 146 277 147 278
rect 145 277 146 278
rect 144 277 145 278
rect 143 277 144 278
rect 142 277 143 278
rect 141 277 142 278
rect 140 277 141 278
rect 139 277 140 278
rect 138 277 139 278
rect 137 277 138 278
rect 136 277 137 278
rect 135 277 136 278
rect 134 277 135 278
rect 133 277 134 278
rect 132 277 133 278
rect 131 277 132 278
rect 130 277 131 278
rect 129 277 130 278
rect 128 277 129 278
rect 127 277 128 278
rect 112 277 113 278
rect 111 277 112 278
rect 110 277 111 278
rect 109 277 110 278
rect 108 277 109 278
rect 107 277 108 278
rect 106 277 107 278
rect 105 277 106 278
rect 104 277 105 278
rect 103 277 104 278
rect 102 277 103 278
rect 101 277 102 278
rect 100 277 101 278
rect 99 277 100 278
rect 98 277 99 278
rect 97 277 98 278
rect 96 277 97 278
rect 95 277 96 278
rect 94 277 95 278
rect 93 277 94 278
rect 92 277 93 278
rect 91 277 92 278
rect 90 277 91 278
rect 89 277 90 278
rect 88 277 89 278
rect 87 277 88 278
rect 86 277 87 278
rect 85 277 86 278
rect 84 277 85 278
rect 83 277 84 278
rect 82 277 83 278
rect 81 277 82 278
rect 80 277 81 278
rect 79 277 80 278
rect 78 277 79 278
rect 61 277 62 278
rect 60 277 61 278
rect 59 277 60 278
rect 58 277 59 278
rect 57 277 58 278
rect 56 277 57 278
rect 55 277 56 278
rect 54 277 55 278
rect 53 277 54 278
rect 52 277 53 278
rect 51 277 52 278
rect 50 277 51 278
rect 49 277 50 278
rect 48 277 49 278
rect 47 277 48 278
rect 46 277 47 278
rect 45 277 46 278
rect 44 277 45 278
rect 43 277 44 278
rect 42 277 43 278
rect 41 277 42 278
rect 40 277 41 278
rect 39 277 40 278
rect 38 277 39 278
rect 37 277 38 278
rect 36 277 37 278
rect 25 277 26 278
rect 24 277 25 278
rect 23 277 24 278
rect 22 277 23 278
rect 21 277 22 278
rect 20 277 21 278
rect 19 277 20 278
rect 18 277 19 278
rect 17 277 18 278
rect 16 277 17 278
rect 15 277 16 278
rect 14 277 15 278
rect 13 277 14 278
rect 12 277 13 278
rect 11 277 12 278
rect 10 277 11 278
rect 9 277 10 278
rect 8 277 9 278
rect 7 277 8 278
rect 6 277 7 278
rect 5 277 6 278
rect 4 277 5 278
rect 3 277 4 278
rect 2 277 3 278
rect 1 277 2 278
rect 437 278 438 279
rect 436 278 437 279
rect 435 278 436 279
rect 434 278 435 279
rect 433 278 434 279
rect 432 278 433 279
rect 431 278 432 279
rect 430 278 431 279
rect 429 278 430 279
rect 428 278 429 279
rect 427 278 428 279
rect 426 278 427 279
rect 425 278 426 279
rect 424 278 425 279
rect 423 278 424 279
rect 422 278 423 279
rect 421 278 422 279
rect 420 278 421 279
rect 419 278 420 279
rect 418 278 419 279
rect 417 278 418 279
rect 416 278 417 279
rect 415 278 416 279
rect 414 278 415 279
rect 413 278 414 279
rect 412 278 413 279
rect 411 278 412 279
rect 410 278 411 279
rect 409 278 410 279
rect 408 278 409 279
rect 407 278 408 279
rect 406 278 407 279
rect 405 278 406 279
rect 404 278 405 279
rect 403 278 404 279
rect 402 278 403 279
rect 401 278 402 279
rect 400 278 401 279
rect 399 278 400 279
rect 398 278 399 279
rect 397 278 398 279
rect 396 278 397 279
rect 395 278 396 279
rect 394 278 395 279
rect 393 278 394 279
rect 287 278 288 279
rect 286 278 287 279
rect 285 278 286 279
rect 284 278 285 279
rect 283 278 284 279
rect 282 278 283 279
rect 281 278 282 279
rect 280 278 281 279
rect 279 278 280 279
rect 278 278 279 279
rect 277 278 278 279
rect 276 278 277 279
rect 275 278 276 279
rect 274 278 275 279
rect 273 278 274 279
rect 272 278 273 279
rect 271 278 272 279
rect 270 278 271 279
rect 269 278 270 279
rect 268 278 269 279
rect 267 278 268 279
rect 266 278 267 279
rect 265 278 266 279
rect 264 278 265 279
rect 263 278 264 279
rect 262 278 263 279
rect 261 278 262 279
rect 260 278 261 279
rect 259 278 260 279
rect 258 278 259 279
rect 257 278 258 279
rect 256 278 257 279
rect 255 278 256 279
rect 254 278 255 279
rect 253 278 254 279
rect 252 278 253 279
rect 251 278 252 279
rect 250 278 251 279
rect 249 278 250 279
rect 248 278 249 279
rect 247 278 248 279
rect 246 278 247 279
rect 245 278 246 279
rect 244 278 245 279
rect 243 278 244 279
rect 242 278 243 279
rect 241 278 242 279
rect 240 278 241 279
rect 239 278 240 279
rect 238 278 239 279
rect 237 278 238 279
rect 236 278 237 279
rect 235 278 236 279
rect 234 278 235 279
rect 233 278 234 279
rect 232 278 233 279
rect 231 278 232 279
rect 230 278 231 279
rect 229 278 230 279
rect 228 278 229 279
rect 227 278 228 279
rect 226 278 227 279
rect 225 278 226 279
rect 224 278 225 279
rect 223 278 224 279
rect 222 278 223 279
rect 221 278 222 279
rect 220 278 221 279
rect 219 278 220 279
rect 218 278 219 279
rect 196 278 197 279
rect 195 278 196 279
rect 194 278 195 279
rect 193 278 194 279
rect 192 278 193 279
rect 191 278 192 279
rect 190 278 191 279
rect 189 278 190 279
rect 188 278 189 279
rect 187 278 188 279
rect 186 278 187 279
rect 185 278 186 279
rect 184 278 185 279
rect 183 278 184 279
rect 182 278 183 279
rect 181 278 182 279
rect 180 278 181 279
rect 179 278 180 279
rect 178 278 179 279
rect 177 278 178 279
rect 176 278 177 279
rect 175 278 176 279
rect 174 278 175 279
rect 173 278 174 279
rect 172 278 173 279
rect 171 278 172 279
rect 170 278 171 279
rect 169 278 170 279
rect 168 278 169 279
rect 167 278 168 279
rect 166 278 167 279
rect 165 278 166 279
rect 164 278 165 279
rect 163 278 164 279
rect 162 278 163 279
rect 161 278 162 279
rect 160 278 161 279
rect 159 278 160 279
rect 158 278 159 279
rect 157 278 158 279
rect 156 278 157 279
rect 155 278 156 279
rect 154 278 155 279
rect 153 278 154 279
rect 152 278 153 279
rect 151 278 152 279
rect 150 278 151 279
rect 149 278 150 279
rect 148 278 149 279
rect 147 278 148 279
rect 146 278 147 279
rect 145 278 146 279
rect 144 278 145 279
rect 143 278 144 279
rect 142 278 143 279
rect 141 278 142 279
rect 140 278 141 279
rect 139 278 140 279
rect 138 278 139 279
rect 137 278 138 279
rect 136 278 137 279
rect 135 278 136 279
rect 134 278 135 279
rect 133 278 134 279
rect 132 278 133 279
rect 131 278 132 279
rect 130 278 131 279
rect 129 278 130 279
rect 128 278 129 279
rect 127 278 128 279
rect 112 278 113 279
rect 111 278 112 279
rect 110 278 111 279
rect 109 278 110 279
rect 108 278 109 279
rect 107 278 108 279
rect 106 278 107 279
rect 105 278 106 279
rect 104 278 105 279
rect 103 278 104 279
rect 102 278 103 279
rect 101 278 102 279
rect 100 278 101 279
rect 99 278 100 279
rect 98 278 99 279
rect 97 278 98 279
rect 96 278 97 279
rect 95 278 96 279
rect 94 278 95 279
rect 93 278 94 279
rect 92 278 93 279
rect 91 278 92 279
rect 90 278 91 279
rect 89 278 90 279
rect 88 278 89 279
rect 87 278 88 279
rect 86 278 87 279
rect 85 278 86 279
rect 84 278 85 279
rect 83 278 84 279
rect 82 278 83 279
rect 81 278 82 279
rect 80 278 81 279
rect 79 278 80 279
rect 78 278 79 279
rect 62 278 63 279
rect 61 278 62 279
rect 60 278 61 279
rect 59 278 60 279
rect 58 278 59 279
rect 57 278 58 279
rect 56 278 57 279
rect 55 278 56 279
rect 54 278 55 279
rect 53 278 54 279
rect 52 278 53 279
rect 51 278 52 279
rect 50 278 51 279
rect 49 278 50 279
rect 48 278 49 279
rect 47 278 48 279
rect 46 278 47 279
rect 45 278 46 279
rect 44 278 45 279
rect 43 278 44 279
rect 42 278 43 279
rect 41 278 42 279
rect 40 278 41 279
rect 39 278 40 279
rect 38 278 39 279
rect 37 278 38 279
rect 36 278 37 279
rect 26 278 27 279
rect 25 278 26 279
rect 24 278 25 279
rect 23 278 24 279
rect 22 278 23 279
rect 21 278 22 279
rect 20 278 21 279
rect 19 278 20 279
rect 18 278 19 279
rect 17 278 18 279
rect 16 278 17 279
rect 15 278 16 279
rect 14 278 15 279
rect 13 278 14 279
rect 12 278 13 279
rect 11 278 12 279
rect 10 278 11 279
rect 9 278 10 279
rect 8 278 9 279
rect 7 278 8 279
rect 6 278 7 279
rect 5 278 6 279
rect 4 278 5 279
rect 3 278 4 279
rect 2 278 3 279
rect 1 278 2 279
rect 437 279 438 280
rect 436 279 437 280
rect 435 279 436 280
rect 434 279 435 280
rect 433 279 434 280
rect 432 279 433 280
rect 431 279 432 280
rect 430 279 431 280
rect 429 279 430 280
rect 428 279 429 280
rect 427 279 428 280
rect 426 279 427 280
rect 425 279 426 280
rect 424 279 425 280
rect 423 279 424 280
rect 422 279 423 280
rect 421 279 422 280
rect 420 279 421 280
rect 419 279 420 280
rect 418 279 419 280
rect 417 279 418 280
rect 416 279 417 280
rect 415 279 416 280
rect 414 279 415 280
rect 413 279 414 280
rect 412 279 413 280
rect 411 279 412 280
rect 410 279 411 280
rect 409 279 410 280
rect 408 279 409 280
rect 407 279 408 280
rect 406 279 407 280
rect 405 279 406 280
rect 404 279 405 280
rect 403 279 404 280
rect 402 279 403 280
rect 401 279 402 280
rect 400 279 401 280
rect 399 279 400 280
rect 398 279 399 280
rect 397 279 398 280
rect 396 279 397 280
rect 395 279 396 280
rect 394 279 395 280
rect 393 279 394 280
rect 286 279 287 280
rect 285 279 286 280
rect 284 279 285 280
rect 283 279 284 280
rect 282 279 283 280
rect 281 279 282 280
rect 280 279 281 280
rect 279 279 280 280
rect 278 279 279 280
rect 277 279 278 280
rect 276 279 277 280
rect 275 279 276 280
rect 274 279 275 280
rect 273 279 274 280
rect 272 279 273 280
rect 271 279 272 280
rect 270 279 271 280
rect 269 279 270 280
rect 268 279 269 280
rect 267 279 268 280
rect 266 279 267 280
rect 265 279 266 280
rect 264 279 265 280
rect 263 279 264 280
rect 262 279 263 280
rect 261 279 262 280
rect 260 279 261 280
rect 259 279 260 280
rect 258 279 259 280
rect 257 279 258 280
rect 256 279 257 280
rect 255 279 256 280
rect 254 279 255 280
rect 253 279 254 280
rect 252 279 253 280
rect 251 279 252 280
rect 250 279 251 280
rect 249 279 250 280
rect 248 279 249 280
rect 247 279 248 280
rect 246 279 247 280
rect 245 279 246 280
rect 244 279 245 280
rect 243 279 244 280
rect 242 279 243 280
rect 241 279 242 280
rect 240 279 241 280
rect 239 279 240 280
rect 238 279 239 280
rect 237 279 238 280
rect 236 279 237 280
rect 235 279 236 280
rect 234 279 235 280
rect 233 279 234 280
rect 232 279 233 280
rect 231 279 232 280
rect 230 279 231 280
rect 229 279 230 280
rect 228 279 229 280
rect 227 279 228 280
rect 226 279 227 280
rect 225 279 226 280
rect 224 279 225 280
rect 223 279 224 280
rect 222 279 223 280
rect 221 279 222 280
rect 220 279 221 280
rect 219 279 220 280
rect 218 279 219 280
rect 196 279 197 280
rect 195 279 196 280
rect 194 279 195 280
rect 193 279 194 280
rect 192 279 193 280
rect 191 279 192 280
rect 190 279 191 280
rect 189 279 190 280
rect 188 279 189 280
rect 187 279 188 280
rect 186 279 187 280
rect 185 279 186 280
rect 184 279 185 280
rect 183 279 184 280
rect 182 279 183 280
rect 181 279 182 280
rect 180 279 181 280
rect 179 279 180 280
rect 178 279 179 280
rect 177 279 178 280
rect 176 279 177 280
rect 175 279 176 280
rect 174 279 175 280
rect 173 279 174 280
rect 172 279 173 280
rect 171 279 172 280
rect 170 279 171 280
rect 169 279 170 280
rect 168 279 169 280
rect 167 279 168 280
rect 166 279 167 280
rect 165 279 166 280
rect 164 279 165 280
rect 163 279 164 280
rect 162 279 163 280
rect 161 279 162 280
rect 160 279 161 280
rect 159 279 160 280
rect 158 279 159 280
rect 157 279 158 280
rect 156 279 157 280
rect 155 279 156 280
rect 154 279 155 280
rect 153 279 154 280
rect 152 279 153 280
rect 151 279 152 280
rect 150 279 151 280
rect 149 279 150 280
rect 148 279 149 280
rect 147 279 148 280
rect 146 279 147 280
rect 145 279 146 280
rect 144 279 145 280
rect 143 279 144 280
rect 142 279 143 280
rect 141 279 142 280
rect 140 279 141 280
rect 139 279 140 280
rect 138 279 139 280
rect 137 279 138 280
rect 136 279 137 280
rect 135 279 136 280
rect 134 279 135 280
rect 133 279 134 280
rect 132 279 133 280
rect 131 279 132 280
rect 130 279 131 280
rect 129 279 130 280
rect 128 279 129 280
rect 112 279 113 280
rect 111 279 112 280
rect 110 279 111 280
rect 109 279 110 280
rect 108 279 109 280
rect 107 279 108 280
rect 106 279 107 280
rect 105 279 106 280
rect 104 279 105 280
rect 103 279 104 280
rect 102 279 103 280
rect 101 279 102 280
rect 100 279 101 280
rect 99 279 100 280
rect 98 279 99 280
rect 97 279 98 280
rect 96 279 97 280
rect 95 279 96 280
rect 94 279 95 280
rect 93 279 94 280
rect 92 279 93 280
rect 91 279 92 280
rect 90 279 91 280
rect 89 279 90 280
rect 88 279 89 280
rect 87 279 88 280
rect 86 279 87 280
rect 85 279 86 280
rect 84 279 85 280
rect 83 279 84 280
rect 82 279 83 280
rect 81 279 82 280
rect 80 279 81 280
rect 79 279 80 280
rect 78 279 79 280
rect 62 279 63 280
rect 61 279 62 280
rect 60 279 61 280
rect 59 279 60 280
rect 58 279 59 280
rect 57 279 58 280
rect 56 279 57 280
rect 55 279 56 280
rect 54 279 55 280
rect 53 279 54 280
rect 52 279 53 280
rect 51 279 52 280
rect 50 279 51 280
rect 49 279 50 280
rect 48 279 49 280
rect 47 279 48 280
rect 46 279 47 280
rect 45 279 46 280
rect 44 279 45 280
rect 43 279 44 280
rect 42 279 43 280
rect 41 279 42 280
rect 40 279 41 280
rect 39 279 40 280
rect 38 279 39 280
rect 37 279 38 280
rect 36 279 37 280
rect 26 279 27 280
rect 25 279 26 280
rect 24 279 25 280
rect 23 279 24 280
rect 22 279 23 280
rect 21 279 22 280
rect 20 279 21 280
rect 19 279 20 280
rect 18 279 19 280
rect 17 279 18 280
rect 16 279 17 280
rect 15 279 16 280
rect 14 279 15 280
rect 13 279 14 280
rect 12 279 13 280
rect 11 279 12 280
rect 10 279 11 280
rect 9 279 10 280
rect 8 279 9 280
rect 7 279 8 280
rect 6 279 7 280
rect 5 279 6 280
rect 4 279 5 280
rect 3 279 4 280
rect 2 279 3 280
rect 1 279 2 280
rect 437 280 438 281
rect 436 280 437 281
rect 435 280 436 281
rect 434 280 435 281
rect 433 280 434 281
rect 432 280 433 281
rect 431 280 432 281
rect 430 280 431 281
rect 429 280 430 281
rect 428 280 429 281
rect 427 280 428 281
rect 426 280 427 281
rect 425 280 426 281
rect 424 280 425 281
rect 423 280 424 281
rect 422 280 423 281
rect 421 280 422 281
rect 420 280 421 281
rect 419 280 420 281
rect 418 280 419 281
rect 417 280 418 281
rect 416 280 417 281
rect 415 280 416 281
rect 414 280 415 281
rect 413 280 414 281
rect 412 280 413 281
rect 411 280 412 281
rect 410 280 411 281
rect 409 280 410 281
rect 408 280 409 281
rect 407 280 408 281
rect 406 280 407 281
rect 405 280 406 281
rect 404 280 405 281
rect 403 280 404 281
rect 402 280 403 281
rect 401 280 402 281
rect 400 280 401 281
rect 399 280 400 281
rect 398 280 399 281
rect 397 280 398 281
rect 396 280 397 281
rect 395 280 396 281
rect 394 280 395 281
rect 393 280 394 281
rect 285 280 286 281
rect 284 280 285 281
rect 283 280 284 281
rect 282 280 283 281
rect 281 280 282 281
rect 280 280 281 281
rect 279 280 280 281
rect 278 280 279 281
rect 277 280 278 281
rect 276 280 277 281
rect 275 280 276 281
rect 274 280 275 281
rect 273 280 274 281
rect 272 280 273 281
rect 271 280 272 281
rect 270 280 271 281
rect 269 280 270 281
rect 268 280 269 281
rect 267 280 268 281
rect 266 280 267 281
rect 265 280 266 281
rect 264 280 265 281
rect 263 280 264 281
rect 262 280 263 281
rect 261 280 262 281
rect 260 280 261 281
rect 259 280 260 281
rect 258 280 259 281
rect 257 280 258 281
rect 256 280 257 281
rect 255 280 256 281
rect 254 280 255 281
rect 253 280 254 281
rect 252 280 253 281
rect 251 280 252 281
rect 250 280 251 281
rect 249 280 250 281
rect 248 280 249 281
rect 247 280 248 281
rect 246 280 247 281
rect 245 280 246 281
rect 244 280 245 281
rect 243 280 244 281
rect 242 280 243 281
rect 241 280 242 281
rect 240 280 241 281
rect 239 280 240 281
rect 238 280 239 281
rect 237 280 238 281
rect 236 280 237 281
rect 235 280 236 281
rect 234 280 235 281
rect 233 280 234 281
rect 232 280 233 281
rect 231 280 232 281
rect 230 280 231 281
rect 229 280 230 281
rect 228 280 229 281
rect 227 280 228 281
rect 226 280 227 281
rect 225 280 226 281
rect 224 280 225 281
rect 223 280 224 281
rect 222 280 223 281
rect 221 280 222 281
rect 220 280 221 281
rect 219 280 220 281
rect 218 280 219 281
rect 217 280 218 281
rect 195 280 196 281
rect 194 280 195 281
rect 193 280 194 281
rect 192 280 193 281
rect 191 280 192 281
rect 190 280 191 281
rect 189 280 190 281
rect 188 280 189 281
rect 187 280 188 281
rect 186 280 187 281
rect 185 280 186 281
rect 184 280 185 281
rect 183 280 184 281
rect 182 280 183 281
rect 181 280 182 281
rect 180 280 181 281
rect 179 280 180 281
rect 178 280 179 281
rect 177 280 178 281
rect 176 280 177 281
rect 175 280 176 281
rect 174 280 175 281
rect 173 280 174 281
rect 172 280 173 281
rect 171 280 172 281
rect 170 280 171 281
rect 169 280 170 281
rect 168 280 169 281
rect 167 280 168 281
rect 166 280 167 281
rect 165 280 166 281
rect 164 280 165 281
rect 163 280 164 281
rect 162 280 163 281
rect 161 280 162 281
rect 160 280 161 281
rect 159 280 160 281
rect 158 280 159 281
rect 157 280 158 281
rect 156 280 157 281
rect 155 280 156 281
rect 154 280 155 281
rect 153 280 154 281
rect 152 280 153 281
rect 151 280 152 281
rect 150 280 151 281
rect 149 280 150 281
rect 148 280 149 281
rect 147 280 148 281
rect 146 280 147 281
rect 145 280 146 281
rect 144 280 145 281
rect 143 280 144 281
rect 142 280 143 281
rect 141 280 142 281
rect 140 280 141 281
rect 139 280 140 281
rect 138 280 139 281
rect 137 280 138 281
rect 136 280 137 281
rect 135 280 136 281
rect 134 280 135 281
rect 133 280 134 281
rect 132 280 133 281
rect 131 280 132 281
rect 130 280 131 281
rect 129 280 130 281
rect 128 280 129 281
rect 113 280 114 281
rect 112 280 113 281
rect 111 280 112 281
rect 110 280 111 281
rect 109 280 110 281
rect 108 280 109 281
rect 107 280 108 281
rect 106 280 107 281
rect 105 280 106 281
rect 104 280 105 281
rect 103 280 104 281
rect 102 280 103 281
rect 101 280 102 281
rect 100 280 101 281
rect 99 280 100 281
rect 98 280 99 281
rect 97 280 98 281
rect 96 280 97 281
rect 95 280 96 281
rect 94 280 95 281
rect 93 280 94 281
rect 92 280 93 281
rect 91 280 92 281
rect 90 280 91 281
rect 89 280 90 281
rect 88 280 89 281
rect 87 280 88 281
rect 86 280 87 281
rect 85 280 86 281
rect 84 280 85 281
rect 83 280 84 281
rect 82 280 83 281
rect 81 280 82 281
rect 80 280 81 281
rect 79 280 80 281
rect 62 280 63 281
rect 61 280 62 281
rect 60 280 61 281
rect 59 280 60 281
rect 58 280 59 281
rect 57 280 58 281
rect 56 280 57 281
rect 55 280 56 281
rect 54 280 55 281
rect 53 280 54 281
rect 52 280 53 281
rect 51 280 52 281
rect 50 280 51 281
rect 49 280 50 281
rect 48 280 49 281
rect 47 280 48 281
rect 46 280 47 281
rect 45 280 46 281
rect 44 280 45 281
rect 43 280 44 281
rect 42 280 43 281
rect 41 280 42 281
rect 40 280 41 281
rect 39 280 40 281
rect 38 280 39 281
rect 37 280 38 281
rect 36 280 37 281
rect 26 280 27 281
rect 25 280 26 281
rect 24 280 25 281
rect 23 280 24 281
rect 22 280 23 281
rect 21 280 22 281
rect 20 280 21 281
rect 19 280 20 281
rect 18 280 19 281
rect 17 280 18 281
rect 16 280 17 281
rect 15 280 16 281
rect 14 280 15 281
rect 13 280 14 281
rect 12 280 13 281
rect 11 280 12 281
rect 10 280 11 281
rect 9 280 10 281
rect 8 280 9 281
rect 7 280 8 281
rect 6 280 7 281
rect 5 280 6 281
rect 4 280 5 281
rect 3 280 4 281
rect 2 280 3 281
rect 1 280 2 281
rect 437 281 438 282
rect 436 281 437 282
rect 435 281 436 282
rect 434 281 435 282
rect 433 281 434 282
rect 432 281 433 282
rect 431 281 432 282
rect 430 281 431 282
rect 429 281 430 282
rect 428 281 429 282
rect 427 281 428 282
rect 426 281 427 282
rect 425 281 426 282
rect 424 281 425 282
rect 423 281 424 282
rect 422 281 423 282
rect 421 281 422 282
rect 420 281 421 282
rect 419 281 420 282
rect 418 281 419 282
rect 417 281 418 282
rect 416 281 417 282
rect 415 281 416 282
rect 414 281 415 282
rect 413 281 414 282
rect 412 281 413 282
rect 411 281 412 282
rect 410 281 411 282
rect 409 281 410 282
rect 408 281 409 282
rect 407 281 408 282
rect 406 281 407 282
rect 405 281 406 282
rect 404 281 405 282
rect 403 281 404 282
rect 402 281 403 282
rect 401 281 402 282
rect 400 281 401 282
rect 399 281 400 282
rect 398 281 399 282
rect 397 281 398 282
rect 396 281 397 282
rect 395 281 396 282
rect 394 281 395 282
rect 393 281 394 282
rect 284 281 285 282
rect 283 281 284 282
rect 282 281 283 282
rect 281 281 282 282
rect 280 281 281 282
rect 279 281 280 282
rect 278 281 279 282
rect 277 281 278 282
rect 276 281 277 282
rect 275 281 276 282
rect 274 281 275 282
rect 273 281 274 282
rect 272 281 273 282
rect 271 281 272 282
rect 270 281 271 282
rect 269 281 270 282
rect 268 281 269 282
rect 267 281 268 282
rect 266 281 267 282
rect 265 281 266 282
rect 264 281 265 282
rect 263 281 264 282
rect 262 281 263 282
rect 261 281 262 282
rect 260 281 261 282
rect 259 281 260 282
rect 258 281 259 282
rect 257 281 258 282
rect 256 281 257 282
rect 255 281 256 282
rect 254 281 255 282
rect 253 281 254 282
rect 252 281 253 282
rect 251 281 252 282
rect 250 281 251 282
rect 249 281 250 282
rect 248 281 249 282
rect 247 281 248 282
rect 246 281 247 282
rect 245 281 246 282
rect 244 281 245 282
rect 243 281 244 282
rect 242 281 243 282
rect 241 281 242 282
rect 240 281 241 282
rect 239 281 240 282
rect 238 281 239 282
rect 237 281 238 282
rect 236 281 237 282
rect 235 281 236 282
rect 234 281 235 282
rect 233 281 234 282
rect 232 281 233 282
rect 231 281 232 282
rect 230 281 231 282
rect 229 281 230 282
rect 228 281 229 282
rect 227 281 228 282
rect 226 281 227 282
rect 225 281 226 282
rect 224 281 225 282
rect 223 281 224 282
rect 222 281 223 282
rect 221 281 222 282
rect 220 281 221 282
rect 219 281 220 282
rect 218 281 219 282
rect 217 281 218 282
rect 194 281 195 282
rect 193 281 194 282
rect 192 281 193 282
rect 191 281 192 282
rect 190 281 191 282
rect 189 281 190 282
rect 188 281 189 282
rect 187 281 188 282
rect 186 281 187 282
rect 185 281 186 282
rect 184 281 185 282
rect 183 281 184 282
rect 182 281 183 282
rect 181 281 182 282
rect 180 281 181 282
rect 179 281 180 282
rect 178 281 179 282
rect 177 281 178 282
rect 176 281 177 282
rect 175 281 176 282
rect 174 281 175 282
rect 173 281 174 282
rect 172 281 173 282
rect 171 281 172 282
rect 170 281 171 282
rect 169 281 170 282
rect 168 281 169 282
rect 167 281 168 282
rect 166 281 167 282
rect 165 281 166 282
rect 164 281 165 282
rect 163 281 164 282
rect 162 281 163 282
rect 161 281 162 282
rect 160 281 161 282
rect 159 281 160 282
rect 158 281 159 282
rect 157 281 158 282
rect 156 281 157 282
rect 155 281 156 282
rect 154 281 155 282
rect 153 281 154 282
rect 152 281 153 282
rect 151 281 152 282
rect 150 281 151 282
rect 149 281 150 282
rect 148 281 149 282
rect 147 281 148 282
rect 146 281 147 282
rect 145 281 146 282
rect 144 281 145 282
rect 143 281 144 282
rect 142 281 143 282
rect 141 281 142 282
rect 140 281 141 282
rect 139 281 140 282
rect 138 281 139 282
rect 137 281 138 282
rect 136 281 137 282
rect 135 281 136 282
rect 134 281 135 282
rect 133 281 134 282
rect 132 281 133 282
rect 131 281 132 282
rect 130 281 131 282
rect 129 281 130 282
rect 113 281 114 282
rect 112 281 113 282
rect 111 281 112 282
rect 110 281 111 282
rect 109 281 110 282
rect 108 281 109 282
rect 107 281 108 282
rect 106 281 107 282
rect 105 281 106 282
rect 104 281 105 282
rect 103 281 104 282
rect 102 281 103 282
rect 101 281 102 282
rect 100 281 101 282
rect 99 281 100 282
rect 98 281 99 282
rect 97 281 98 282
rect 96 281 97 282
rect 95 281 96 282
rect 94 281 95 282
rect 93 281 94 282
rect 92 281 93 282
rect 91 281 92 282
rect 90 281 91 282
rect 89 281 90 282
rect 88 281 89 282
rect 87 281 88 282
rect 86 281 87 282
rect 85 281 86 282
rect 84 281 85 282
rect 83 281 84 282
rect 82 281 83 282
rect 81 281 82 282
rect 80 281 81 282
rect 79 281 80 282
rect 63 281 64 282
rect 62 281 63 282
rect 61 281 62 282
rect 60 281 61 282
rect 59 281 60 282
rect 58 281 59 282
rect 57 281 58 282
rect 56 281 57 282
rect 55 281 56 282
rect 54 281 55 282
rect 53 281 54 282
rect 52 281 53 282
rect 51 281 52 282
rect 50 281 51 282
rect 49 281 50 282
rect 48 281 49 282
rect 47 281 48 282
rect 46 281 47 282
rect 45 281 46 282
rect 44 281 45 282
rect 43 281 44 282
rect 42 281 43 282
rect 41 281 42 282
rect 40 281 41 282
rect 39 281 40 282
rect 38 281 39 282
rect 37 281 38 282
rect 36 281 37 282
rect 26 281 27 282
rect 25 281 26 282
rect 24 281 25 282
rect 23 281 24 282
rect 22 281 23 282
rect 21 281 22 282
rect 20 281 21 282
rect 19 281 20 282
rect 18 281 19 282
rect 17 281 18 282
rect 16 281 17 282
rect 15 281 16 282
rect 14 281 15 282
rect 13 281 14 282
rect 12 281 13 282
rect 11 281 12 282
rect 10 281 11 282
rect 9 281 10 282
rect 8 281 9 282
rect 7 281 8 282
rect 6 281 7 282
rect 5 281 6 282
rect 4 281 5 282
rect 3 281 4 282
rect 2 281 3 282
rect 1 281 2 282
rect 462 282 463 283
rect 437 282 438 283
rect 436 282 437 283
rect 435 282 436 283
rect 434 282 435 283
rect 433 282 434 283
rect 432 282 433 283
rect 431 282 432 283
rect 430 282 431 283
rect 429 282 430 283
rect 428 282 429 283
rect 427 282 428 283
rect 426 282 427 283
rect 425 282 426 283
rect 424 282 425 283
rect 423 282 424 283
rect 422 282 423 283
rect 421 282 422 283
rect 420 282 421 283
rect 419 282 420 283
rect 418 282 419 283
rect 417 282 418 283
rect 416 282 417 283
rect 415 282 416 283
rect 414 282 415 283
rect 413 282 414 283
rect 412 282 413 283
rect 411 282 412 283
rect 410 282 411 283
rect 409 282 410 283
rect 408 282 409 283
rect 407 282 408 283
rect 406 282 407 283
rect 405 282 406 283
rect 404 282 405 283
rect 403 282 404 283
rect 402 282 403 283
rect 401 282 402 283
rect 400 282 401 283
rect 399 282 400 283
rect 398 282 399 283
rect 397 282 398 283
rect 396 282 397 283
rect 395 282 396 283
rect 394 282 395 283
rect 393 282 394 283
rect 283 282 284 283
rect 282 282 283 283
rect 281 282 282 283
rect 280 282 281 283
rect 279 282 280 283
rect 278 282 279 283
rect 277 282 278 283
rect 276 282 277 283
rect 275 282 276 283
rect 274 282 275 283
rect 273 282 274 283
rect 272 282 273 283
rect 271 282 272 283
rect 270 282 271 283
rect 269 282 270 283
rect 268 282 269 283
rect 267 282 268 283
rect 266 282 267 283
rect 265 282 266 283
rect 264 282 265 283
rect 263 282 264 283
rect 262 282 263 283
rect 261 282 262 283
rect 260 282 261 283
rect 259 282 260 283
rect 258 282 259 283
rect 257 282 258 283
rect 256 282 257 283
rect 255 282 256 283
rect 254 282 255 283
rect 253 282 254 283
rect 252 282 253 283
rect 251 282 252 283
rect 250 282 251 283
rect 249 282 250 283
rect 248 282 249 283
rect 247 282 248 283
rect 246 282 247 283
rect 245 282 246 283
rect 244 282 245 283
rect 243 282 244 283
rect 242 282 243 283
rect 241 282 242 283
rect 240 282 241 283
rect 239 282 240 283
rect 238 282 239 283
rect 237 282 238 283
rect 236 282 237 283
rect 235 282 236 283
rect 234 282 235 283
rect 233 282 234 283
rect 232 282 233 283
rect 231 282 232 283
rect 230 282 231 283
rect 229 282 230 283
rect 228 282 229 283
rect 227 282 228 283
rect 226 282 227 283
rect 225 282 226 283
rect 224 282 225 283
rect 223 282 224 283
rect 222 282 223 283
rect 221 282 222 283
rect 220 282 221 283
rect 219 282 220 283
rect 218 282 219 283
rect 217 282 218 283
rect 216 282 217 283
rect 194 282 195 283
rect 193 282 194 283
rect 192 282 193 283
rect 191 282 192 283
rect 190 282 191 283
rect 189 282 190 283
rect 188 282 189 283
rect 187 282 188 283
rect 186 282 187 283
rect 185 282 186 283
rect 184 282 185 283
rect 183 282 184 283
rect 182 282 183 283
rect 181 282 182 283
rect 180 282 181 283
rect 179 282 180 283
rect 178 282 179 283
rect 177 282 178 283
rect 176 282 177 283
rect 175 282 176 283
rect 174 282 175 283
rect 173 282 174 283
rect 172 282 173 283
rect 171 282 172 283
rect 170 282 171 283
rect 169 282 170 283
rect 168 282 169 283
rect 167 282 168 283
rect 166 282 167 283
rect 165 282 166 283
rect 164 282 165 283
rect 163 282 164 283
rect 162 282 163 283
rect 161 282 162 283
rect 160 282 161 283
rect 159 282 160 283
rect 158 282 159 283
rect 157 282 158 283
rect 156 282 157 283
rect 155 282 156 283
rect 154 282 155 283
rect 153 282 154 283
rect 152 282 153 283
rect 151 282 152 283
rect 150 282 151 283
rect 149 282 150 283
rect 148 282 149 283
rect 147 282 148 283
rect 146 282 147 283
rect 145 282 146 283
rect 144 282 145 283
rect 143 282 144 283
rect 142 282 143 283
rect 141 282 142 283
rect 140 282 141 283
rect 139 282 140 283
rect 138 282 139 283
rect 137 282 138 283
rect 136 282 137 283
rect 135 282 136 283
rect 134 282 135 283
rect 133 282 134 283
rect 132 282 133 283
rect 131 282 132 283
rect 130 282 131 283
rect 129 282 130 283
rect 113 282 114 283
rect 112 282 113 283
rect 111 282 112 283
rect 110 282 111 283
rect 109 282 110 283
rect 108 282 109 283
rect 107 282 108 283
rect 106 282 107 283
rect 105 282 106 283
rect 104 282 105 283
rect 103 282 104 283
rect 102 282 103 283
rect 101 282 102 283
rect 100 282 101 283
rect 99 282 100 283
rect 98 282 99 283
rect 97 282 98 283
rect 96 282 97 283
rect 95 282 96 283
rect 94 282 95 283
rect 93 282 94 283
rect 92 282 93 283
rect 91 282 92 283
rect 90 282 91 283
rect 89 282 90 283
rect 88 282 89 283
rect 87 282 88 283
rect 86 282 87 283
rect 85 282 86 283
rect 84 282 85 283
rect 83 282 84 283
rect 82 282 83 283
rect 81 282 82 283
rect 80 282 81 283
rect 79 282 80 283
rect 63 282 64 283
rect 62 282 63 283
rect 61 282 62 283
rect 60 282 61 283
rect 59 282 60 283
rect 58 282 59 283
rect 57 282 58 283
rect 56 282 57 283
rect 55 282 56 283
rect 54 282 55 283
rect 53 282 54 283
rect 52 282 53 283
rect 51 282 52 283
rect 50 282 51 283
rect 49 282 50 283
rect 48 282 49 283
rect 47 282 48 283
rect 46 282 47 283
rect 45 282 46 283
rect 44 282 45 283
rect 43 282 44 283
rect 42 282 43 283
rect 41 282 42 283
rect 40 282 41 283
rect 39 282 40 283
rect 38 282 39 283
rect 37 282 38 283
rect 36 282 37 283
rect 26 282 27 283
rect 25 282 26 283
rect 24 282 25 283
rect 23 282 24 283
rect 22 282 23 283
rect 21 282 22 283
rect 20 282 21 283
rect 19 282 20 283
rect 18 282 19 283
rect 17 282 18 283
rect 16 282 17 283
rect 15 282 16 283
rect 14 282 15 283
rect 13 282 14 283
rect 12 282 13 283
rect 11 282 12 283
rect 10 282 11 283
rect 9 282 10 283
rect 8 282 9 283
rect 7 282 8 283
rect 6 282 7 283
rect 5 282 6 283
rect 4 282 5 283
rect 3 282 4 283
rect 2 282 3 283
rect 1 282 2 283
rect 463 283 464 284
rect 462 283 463 284
rect 461 283 462 284
rect 460 283 461 284
rect 459 283 460 284
rect 458 283 459 284
rect 457 283 458 284
rect 437 283 438 284
rect 436 283 437 284
rect 435 283 436 284
rect 434 283 435 284
rect 433 283 434 284
rect 432 283 433 284
rect 431 283 432 284
rect 430 283 431 284
rect 429 283 430 284
rect 428 283 429 284
rect 427 283 428 284
rect 426 283 427 284
rect 425 283 426 284
rect 424 283 425 284
rect 423 283 424 284
rect 422 283 423 284
rect 421 283 422 284
rect 420 283 421 284
rect 419 283 420 284
rect 418 283 419 284
rect 417 283 418 284
rect 416 283 417 284
rect 415 283 416 284
rect 414 283 415 284
rect 413 283 414 284
rect 412 283 413 284
rect 411 283 412 284
rect 410 283 411 284
rect 409 283 410 284
rect 408 283 409 284
rect 407 283 408 284
rect 406 283 407 284
rect 405 283 406 284
rect 404 283 405 284
rect 403 283 404 284
rect 402 283 403 284
rect 401 283 402 284
rect 400 283 401 284
rect 399 283 400 284
rect 398 283 399 284
rect 397 283 398 284
rect 396 283 397 284
rect 395 283 396 284
rect 394 283 395 284
rect 393 283 394 284
rect 282 283 283 284
rect 281 283 282 284
rect 280 283 281 284
rect 279 283 280 284
rect 278 283 279 284
rect 277 283 278 284
rect 276 283 277 284
rect 275 283 276 284
rect 274 283 275 284
rect 273 283 274 284
rect 272 283 273 284
rect 271 283 272 284
rect 270 283 271 284
rect 269 283 270 284
rect 268 283 269 284
rect 267 283 268 284
rect 266 283 267 284
rect 265 283 266 284
rect 264 283 265 284
rect 263 283 264 284
rect 262 283 263 284
rect 261 283 262 284
rect 260 283 261 284
rect 259 283 260 284
rect 258 283 259 284
rect 257 283 258 284
rect 256 283 257 284
rect 255 283 256 284
rect 254 283 255 284
rect 253 283 254 284
rect 252 283 253 284
rect 251 283 252 284
rect 250 283 251 284
rect 249 283 250 284
rect 248 283 249 284
rect 247 283 248 284
rect 246 283 247 284
rect 245 283 246 284
rect 244 283 245 284
rect 243 283 244 284
rect 242 283 243 284
rect 241 283 242 284
rect 240 283 241 284
rect 239 283 240 284
rect 238 283 239 284
rect 237 283 238 284
rect 236 283 237 284
rect 235 283 236 284
rect 234 283 235 284
rect 233 283 234 284
rect 232 283 233 284
rect 231 283 232 284
rect 230 283 231 284
rect 229 283 230 284
rect 228 283 229 284
rect 227 283 228 284
rect 226 283 227 284
rect 225 283 226 284
rect 224 283 225 284
rect 223 283 224 284
rect 222 283 223 284
rect 221 283 222 284
rect 220 283 221 284
rect 219 283 220 284
rect 218 283 219 284
rect 217 283 218 284
rect 216 283 217 284
rect 215 283 216 284
rect 193 283 194 284
rect 192 283 193 284
rect 191 283 192 284
rect 190 283 191 284
rect 189 283 190 284
rect 188 283 189 284
rect 187 283 188 284
rect 186 283 187 284
rect 185 283 186 284
rect 184 283 185 284
rect 183 283 184 284
rect 182 283 183 284
rect 181 283 182 284
rect 180 283 181 284
rect 179 283 180 284
rect 178 283 179 284
rect 177 283 178 284
rect 176 283 177 284
rect 175 283 176 284
rect 174 283 175 284
rect 173 283 174 284
rect 172 283 173 284
rect 171 283 172 284
rect 170 283 171 284
rect 169 283 170 284
rect 168 283 169 284
rect 167 283 168 284
rect 166 283 167 284
rect 165 283 166 284
rect 164 283 165 284
rect 163 283 164 284
rect 162 283 163 284
rect 161 283 162 284
rect 160 283 161 284
rect 159 283 160 284
rect 158 283 159 284
rect 157 283 158 284
rect 156 283 157 284
rect 155 283 156 284
rect 154 283 155 284
rect 153 283 154 284
rect 152 283 153 284
rect 151 283 152 284
rect 150 283 151 284
rect 149 283 150 284
rect 148 283 149 284
rect 147 283 148 284
rect 146 283 147 284
rect 145 283 146 284
rect 144 283 145 284
rect 143 283 144 284
rect 142 283 143 284
rect 141 283 142 284
rect 140 283 141 284
rect 139 283 140 284
rect 138 283 139 284
rect 137 283 138 284
rect 136 283 137 284
rect 135 283 136 284
rect 134 283 135 284
rect 133 283 134 284
rect 132 283 133 284
rect 131 283 132 284
rect 130 283 131 284
rect 114 283 115 284
rect 113 283 114 284
rect 112 283 113 284
rect 111 283 112 284
rect 110 283 111 284
rect 109 283 110 284
rect 108 283 109 284
rect 107 283 108 284
rect 106 283 107 284
rect 105 283 106 284
rect 104 283 105 284
rect 103 283 104 284
rect 102 283 103 284
rect 101 283 102 284
rect 100 283 101 284
rect 99 283 100 284
rect 98 283 99 284
rect 97 283 98 284
rect 96 283 97 284
rect 95 283 96 284
rect 94 283 95 284
rect 93 283 94 284
rect 92 283 93 284
rect 91 283 92 284
rect 90 283 91 284
rect 89 283 90 284
rect 88 283 89 284
rect 87 283 88 284
rect 86 283 87 284
rect 85 283 86 284
rect 84 283 85 284
rect 83 283 84 284
rect 82 283 83 284
rect 81 283 82 284
rect 80 283 81 284
rect 64 283 65 284
rect 63 283 64 284
rect 62 283 63 284
rect 61 283 62 284
rect 60 283 61 284
rect 59 283 60 284
rect 58 283 59 284
rect 57 283 58 284
rect 56 283 57 284
rect 55 283 56 284
rect 54 283 55 284
rect 53 283 54 284
rect 52 283 53 284
rect 51 283 52 284
rect 50 283 51 284
rect 49 283 50 284
rect 48 283 49 284
rect 47 283 48 284
rect 46 283 47 284
rect 45 283 46 284
rect 44 283 45 284
rect 43 283 44 284
rect 42 283 43 284
rect 41 283 42 284
rect 40 283 41 284
rect 39 283 40 284
rect 38 283 39 284
rect 37 283 38 284
rect 36 283 37 284
rect 26 283 27 284
rect 25 283 26 284
rect 24 283 25 284
rect 23 283 24 284
rect 22 283 23 284
rect 21 283 22 284
rect 20 283 21 284
rect 19 283 20 284
rect 18 283 19 284
rect 17 283 18 284
rect 16 283 17 284
rect 15 283 16 284
rect 14 283 15 284
rect 13 283 14 284
rect 12 283 13 284
rect 11 283 12 284
rect 10 283 11 284
rect 9 283 10 284
rect 8 283 9 284
rect 7 283 8 284
rect 6 283 7 284
rect 5 283 6 284
rect 4 283 5 284
rect 3 283 4 284
rect 2 283 3 284
rect 1 283 2 284
rect 460 284 461 285
rect 459 284 460 285
rect 458 284 459 285
rect 457 284 458 285
rect 437 284 438 285
rect 436 284 437 285
rect 435 284 436 285
rect 434 284 435 285
rect 433 284 434 285
rect 432 284 433 285
rect 431 284 432 285
rect 430 284 431 285
rect 429 284 430 285
rect 428 284 429 285
rect 427 284 428 285
rect 426 284 427 285
rect 425 284 426 285
rect 424 284 425 285
rect 423 284 424 285
rect 422 284 423 285
rect 421 284 422 285
rect 420 284 421 285
rect 419 284 420 285
rect 418 284 419 285
rect 417 284 418 285
rect 416 284 417 285
rect 415 284 416 285
rect 414 284 415 285
rect 413 284 414 285
rect 412 284 413 285
rect 411 284 412 285
rect 410 284 411 285
rect 409 284 410 285
rect 408 284 409 285
rect 407 284 408 285
rect 406 284 407 285
rect 405 284 406 285
rect 404 284 405 285
rect 403 284 404 285
rect 402 284 403 285
rect 401 284 402 285
rect 400 284 401 285
rect 399 284 400 285
rect 398 284 399 285
rect 397 284 398 285
rect 396 284 397 285
rect 395 284 396 285
rect 394 284 395 285
rect 393 284 394 285
rect 282 284 283 285
rect 281 284 282 285
rect 280 284 281 285
rect 279 284 280 285
rect 278 284 279 285
rect 277 284 278 285
rect 276 284 277 285
rect 275 284 276 285
rect 274 284 275 285
rect 273 284 274 285
rect 272 284 273 285
rect 271 284 272 285
rect 270 284 271 285
rect 269 284 270 285
rect 268 284 269 285
rect 267 284 268 285
rect 266 284 267 285
rect 265 284 266 285
rect 264 284 265 285
rect 263 284 264 285
rect 262 284 263 285
rect 261 284 262 285
rect 260 284 261 285
rect 259 284 260 285
rect 258 284 259 285
rect 257 284 258 285
rect 256 284 257 285
rect 255 284 256 285
rect 254 284 255 285
rect 253 284 254 285
rect 252 284 253 285
rect 251 284 252 285
rect 250 284 251 285
rect 249 284 250 285
rect 248 284 249 285
rect 247 284 248 285
rect 246 284 247 285
rect 245 284 246 285
rect 244 284 245 285
rect 243 284 244 285
rect 242 284 243 285
rect 241 284 242 285
rect 240 284 241 285
rect 239 284 240 285
rect 238 284 239 285
rect 237 284 238 285
rect 236 284 237 285
rect 235 284 236 285
rect 234 284 235 285
rect 233 284 234 285
rect 232 284 233 285
rect 231 284 232 285
rect 230 284 231 285
rect 229 284 230 285
rect 228 284 229 285
rect 227 284 228 285
rect 226 284 227 285
rect 225 284 226 285
rect 224 284 225 285
rect 223 284 224 285
rect 222 284 223 285
rect 221 284 222 285
rect 220 284 221 285
rect 219 284 220 285
rect 218 284 219 285
rect 217 284 218 285
rect 216 284 217 285
rect 215 284 216 285
rect 192 284 193 285
rect 191 284 192 285
rect 190 284 191 285
rect 189 284 190 285
rect 188 284 189 285
rect 187 284 188 285
rect 186 284 187 285
rect 185 284 186 285
rect 184 284 185 285
rect 183 284 184 285
rect 182 284 183 285
rect 181 284 182 285
rect 180 284 181 285
rect 179 284 180 285
rect 178 284 179 285
rect 177 284 178 285
rect 176 284 177 285
rect 175 284 176 285
rect 174 284 175 285
rect 173 284 174 285
rect 172 284 173 285
rect 171 284 172 285
rect 170 284 171 285
rect 169 284 170 285
rect 168 284 169 285
rect 167 284 168 285
rect 166 284 167 285
rect 165 284 166 285
rect 164 284 165 285
rect 163 284 164 285
rect 162 284 163 285
rect 161 284 162 285
rect 160 284 161 285
rect 159 284 160 285
rect 158 284 159 285
rect 157 284 158 285
rect 156 284 157 285
rect 155 284 156 285
rect 154 284 155 285
rect 153 284 154 285
rect 152 284 153 285
rect 151 284 152 285
rect 150 284 151 285
rect 149 284 150 285
rect 148 284 149 285
rect 147 284 148 285
rect 146 284 147 285
rect 145 284 146 285
rect 144 284 145 285
rect 143 284 144 285
rect 142 284 143 285
rect 141 284 142 285
rect 140 284 141 285
rect 139 284 140 285
rect 138 284 139 285
rect 137 284 138 285
rect 136 284 137 285
rect 135 284 136 285
rect 134 284 135 285
rect 133 284 134 285
rect 132 284 133 285
rect 131 284 132 285
rect 130 284 131 285
rect 114 284 115 285
rect 113 284 114 285
rect 112 284 113 285
rect 111 284 112 285
rect 110 284 111 285
rect 109 284 110 285
rect 108 284 109 285
rect 107 284 108 285
rect 106 284 107 285
rect 105 284 106 285
rect 104 284 105 285
rect 103 284 104 285
rect 102 284 103 285
rect 101 284 102 285
rect 100 284 101 285
rect 99 284 100 285
rect 98 284 99 285
rect 97 284 98 285
rect 96 284 97 285
rect 95 284 96 285
rect 94 284 95 285
rect 93 284 94 285
rect 92 284 93 285
rect 91 284 92 285
rect 90 284 91 285
rect 89 284 90 285
rect 88 284 89 285
rect 87 284 88 285
rect 86 284 87 285
rect 85 284 86 285
rect 84 284 85 285
rect 83 284 84 285
rect 82 284 83 285
rect 81 284 82 285
rect 80 284 81 285
rect 64 284 65 285
rect 63 284 64 285
rect 62 284 63 285
rect 61 284 62 285
rect 60 284 61 285
rect 59 284 60 285
rect 58 284 59 285
rect 57 284 58 285
rect 56 284 57 285
rect 55 284 56 285
rect 54 284 55 285
rect 53 284 54 285
rect 52 284 53 285
rect 51 284 52 285
rect 50 284 51 285
rect 49 284 50 285
rect 48 284 49 285
rect 47 284 48 285
rect 46 284 47 285
rect 45 284 46 285
rect 44 284 45 285
rect 43 284 44 285
rect 42 284 43 285
rect 41 284 42 285
rect 40 284 41 285
rect 39 284 40 285
rect 38 284 39 285
rect 37 284 38 285
rect 36 284 37 285
rect 26 284 27 285
rect 25 284 26 285
rect 24 284 25 285
rect 23 284 24 285
rect 22 284 23 285
rect 21 284 22 285
rect 20 284 21 285
rect 19 284 20 285
rect 18 284 19 285
rect 17 284 18 285
rect 16 284 17 285
rect 15 284 16 285
rect 14 284 15 285
rect 13 284 14 285
rect 12 284 13 285
rect 11 284 12 285
rect 10 284 11 285
rect 9 284 10 285
rect 8 284 9 285
rect 7 284 8 285
rect 6 284 7 285
rect 5 284 6 285
rect 4 284 5 285
rect 3 284 4 285
rect 2 284 3 285
rect 1 284 2 285
rect 459 285 460 286
rect 458 285 459 286
rect 437 285 438 286
rect 436 285 437 286
rect 435 285 436 286
rect 434 285 435 286
rect 433 285 434 286
rect 432 285 433 286
rect 431 285 432 286
rect 430 285 431 286
rect 429 285 430 286
rect 428 285 429 286
rect 427 285 428 286
rect 426 285 427 286
rect 425 285 426 286
rect 424 285 425 286
rect 423 285 424 286
rect 422 285 423 286
rect 421 285 422 286
rect 420 285 421 286
rect 419 285 420 286
rect 418 285 419 286
rect 417 285 418 286
rect 416 285 417 286
rect 415 285 416 286
rect 414 285 415 286
rect 413 285 414 286
rect 412 285 413 286
rect 411 285 412 286
rect 410 285 411 286
rect 409 285 410 286
rect 408 285 409 286
rect 407 285 408 286
rect 406 285 407 286
rect 405 285 406 286
rect 404 285 405 286
rect 403 285 404 286
rect 402 285 403 286
rect 401 285 402 286
rect 400 285 401 286
rect 399 285 400 286
rect 398 285 399 286
rect 397 285 398 286
rect 396 285 397 286
rect 395 285 396 286
rect 394 285 395 286
rect 393 285 394 286
rect 281 285 282 286
rect 280 285 281 286
rect 279 285 280 286
rect 278 285 279 286
rect 277 285 278 286
rect 276 285 277 286
rect 275 285 276 286
rect 274 285 275 286
rect 273 285 274 286
rect 272 285 273 286
rect 271 285 272 286
rect 270 285 271 286
rect 269 285 270 286
rect 268 285 269 286
rect 267 285 268 286
rect 266 285 267 286
rect 265 285 266 286
rect 264 285 265 286
rect 263 285 264 286
rect 262 285 263 286
rect 261 285 262 286
rect 260 285 261 286
rect 259 285 260 286
rect 258 285 259 286
rect 257 285 258 286
rect 256 285 257 286
rect 255 285 256 286
rect 254 285 255 286
rect 253 285 254 286
rect 252 285 253 286
rect 251 285 252 286
rect 250 285 251 286
rect 249 285 250 286
rect 248 285 249 286
rect 247 285 248 286
rect 246 285 247 286
rect 245 285 246 286
rect 244 285 245 286
rect 243 285 244 286
rect 242 285 243 286
rect 241 285 242 286
rect 240 285 241 286
rect 239 285 240 286
rect 238 285 239 286
rect 237 285 238 286
rect 236 285 237 286
rect 235 285 236 286
rect 234 285 235 286
rect 233 285 234 286
rect 232 285 233 286
rect 231 285 232 286
rect 230 285 231 286
rect 229 285 230 286
rect 228 285 229 286
rect 227 285 228 286
rect 226 285 227 286
rect 225 285 226 286
rect 224 285 225 286
rect 223 285 224 286
rect 222 285 223 286
rect 221 285 222 286
rect 220 285 221 286
rect 219 285 220 286
rect 218 285 219 286
rect 217 285 218 286
rect 216 285 217 286
rect 215 285 216 286
rect 214 285 215 286
rect 192 285 193 286
rect 191 285 192 286
rect 190 285 191 286
rect 189 285 190 286
rect 188 285 189 286
rect 187 285 188 286
rect 186 285 187 286
rect 185 285 186 286
rect 184 285 185 286
rect 183 285 184 286
rect 182 285 183 286
rect 181 285 182 286
rect 180 285 181 286
rect 179 285 180 286
rect 178 285 179 286
rect 177 285 178 286
rect 176 285 177 286
rect 175 285 176 286
rect 174 285 175 286
rect 173 285 174 286
rect 172 285 173 286
rect 171 285 172 286
rect 170 285 171 286
rect 169 285 170 286
rect 168 285 169 286
rect 167 285 168 286
rect 166 285 167 286
rect 165 285 166 286
rect 164 285 165 286
rect 163 285 164 286
rect 162 285 163 286
rect 161 285 162 286
rect 160 285 161 286
rect 159 285 160 286
rect 158 285 159 286
rect 157 285 158 286
rect 156 285 157 286
rect 155 285 156 286
rect 154 285 155 286
rect 153 285 154 286
rect 152 285 153 286
rect 151 285 152 286
rect 150 285 151 286
rect 149 285 150 286
rect 148 285 149 286
rect 147 285 148 286
rect 146 285 147 286
rect 145 285 146 286
rect 144 285 145 286
rect 143 285 144 286
rect 142 285 143 286
rect 141 285 142 286
rect 140 285 141 286
rect 139 285 140 286
rect 138 285 139 286
rect 137 285 138 286
rect 136 285 137 286
rect 135 285 136 286
rect 134 285 135 286
rect 133 285 134 286
rect 132 285 133 286
rect 131 285 132 286
rect 114 285 115 286
rect 113 285 114 286
rect 112 285 113 286
rect 111 285 112 286
rect 110 285 111 286
rect 109 285 110 286
rect 108 285 109 286
rect 107 285 108 286
rect 106 285 107 286
rect 105 285 106 286
rect 104 285 105 286
rect 103 285 104 286
rect 102 285 103 286
rect 101 285 102 286
rect 100 285 101 286
rect 99 285 100 286
rect 98 285 99 286
rect 97 285 98 286
rect 96 285 97 286
rect 95 285 96 286
rect 94 285 95 286
rect 93 285 94 286
rect 92 285 93 286
rect 91 285 92 286
rect 90 285 91 286
rect 89 285 90 286
rect 88 285 89 286
rect 87 285 88 286
rect 86 285 87 286
rect 85 285 86 286
rect 84 285 85 286
rect 83 285 84 286
rect 82 285 83 286
rect 81 285 82 286
rect 80 285 81 286
rect 64 285 65 286
rect 63 285 64 286
rect 62 285 63 286
rect 61 285 62 286
rect 60 285 61 286
rect 59 285 60 286
rect 58 285 59 286
rect 57 285 58 286
rect 56 285 57 286
rect 55 285 56 286
rect 54 285 55 286
rect 53 285 54 286
rect 52 285 53 286
rect 51 285 52 286
rect 50 285 51 286
rect 49 285 50 286
rect 48 285 49 286
rect 47 285 48 286
rect 46 285 47 286
rect 45 285 46 286
rect 44 285 45 286
rect 43 285 44 286
rect 42 285 43 286
rect 41 285 42 286
rect 40 285 41 286
rect 39 285 40 286
rect 38 285 39 286
rect 37 285 38 286
rect 36 285 37 286
rect 27 285 28 286
rect 26 285 27 286
rect 25 285 26 286
rect 24 285 25 286
rect 23 285 24 286
rect 22 285 23 286
rect 21 285 22 286
rect 20 285 21 286
rect 19 285 20 286
rect 18 285 19 286
rect 17 285 18 286
rect 16 285 17 286
rect 15 285 16 286
rect 14 285 15 286
rect 13 285 14 286
rect 12 285 13 286
rect 11 285 12 286
rect 10 285 11 286
rect 9 285 10 286
rect 8 285 9 286
rect 7 285 8 286
rect 6 285 7 286
rect 5 285 6 286
rect 4 285 5 286
rect 3 285 4 286
rect 2 285 3 286
rect 1 285 2 286
rect 458 286 459 287
rect 437 286 438 287
rect 436 286 437 287
rect 435 286 436 287
rect 434 286 435 287
rect 433 286 434 287
rect 432 286 433 287
rect 431 286 432 287
rect 430 286 431 287
rect 429 286 430 287
rect 428 286 429 287
rect 427 286 428 287
rect 426 286 427 287
rect 425 286 426 287
rect 424 286 425 287
rect 423 286 424 287
rect 422 286 423 287
rect 421 286 422 287
rect 420 286 421 287
rect 419 286 420 287
rect 418 286 419 287
rect 417 286 418 287
rect 416 286 417 287
rect 415 286 416 287
rect 414 286 415 287
rect 413 286 414 287
rect 412 286 413 287
rect 411 286 412 287
rect 410 286 411 287
rect 409 286 410 287
rect 408 286 409 287
rect 407 286 408 287
rect 406 286 407 287
rect 405 286 406 287
rect 404 286 405 287
rect 403 286 404 287
rect 402 286 403 287
rect 401 286 402 287
rect 400 286 401 287
rect 399 286 400 287
rect 398 286 399 287
rect 397 286 398 287
rect 396 286 397 287
rect 395 286 396 287
rect 394 286 395 287
rect 393 286 394 287
rect 280 286 281 287
rect 279 286 280 287
rect 278 286 279 287
rect 277 286 278 287
rect 276 286 277 287
rect 275 286 276 287
rect 274 286 275 287
rect 273 286 274 287
rect 272 286 273 287
rect 271 286 272 287
rect 270 286 271 287
rect 269 286 270 287
rect 268 286 269 287
rect 267 286 268 287
rect 266 286 267 287
rect 265 286 266 287
rect 264 286 265 287
rect 263 286 264 287
rect 262 286 263 287
rect 261 286 262 287
rect 260 286 261 287
rect 259 286 260 287
rect 258 286 259 287
rect 257 286 258 287
rect 256 286 257 287
rect 255 286 256 287
rect 254 286 255 287
rect 253 286 254 287
rect 252 286 253 287
rect 251 286 252 287
rect 250 286 251 287
rect 249 286 250 287
rect 248 286 249 287
rect 247 286 248 287
rect 246 286 247 287
rect 245 286 246 287
rect 244 286 245 287
rect 243 286 244 287
rect 242 286 243 287
rect 241 286 242 287
rect 240 286 241 287
rect 239 286 240 287
rect 238 286 239 287
rect 237 286 238 287
rect 236 286 237 287
rect 235 286 236 287
rect 234 286 235 287
rect 233 286 234 287
rect 232 286 233 287
rect 231 286 232 287
rect 230 286 231 287
rect 229 286 230 287
rect 228 286 229 287
rect 227 286 228 287
rect 226 286 227 287
rect 225 286 226 287
rect 224 286 225 287
rect 223 286 224 287
rect 222 286 223 287
rect 221 286 222 287
rect 220 286 221 287
rect 219 286 220 287
rect 218 286 219 287
rect 217 286 218 287
rect 216 286 217 287
rect 215 286 216 287
rect 214 286 215 287
rect 191 286 192 287
rect 190 286 191 287
rect 189 286 190 287
rect 188 286 189 287
rect 187 286 188 287
rect 186 286 187 287
rect 185 286 186 287
rect 184 286 185 287
rect 183 286 184 287
rect 182 286 183 287
rect 181 286 182 287
rect 180 286 181 287
rect 179 286 180 287
rect 178 286 179 287
rect 177 286 178 287
rect 176 286 177 287
rect 175 286 176 287
rect 174 286 175 287
rect 173 286 174 287
rect 172 286 173 287
rect 171 286 172 287
rect 170 286 171 287
rect 169 286 170 287
rect 168 286 169 287
rect 167 286 168 287
rect 166 286 167 287
rect 165 286 166 287
rect 164 286 165 287
rect 163 286 164 287
rect 162 286 163 287
rect 161 286 162 287
rect 160 286 161 287
rect 159 286 160 287
rect 158 286 159 287
rect 157 286 158 287
rect 156 286 157 287
rect 155 286 156 287
rect 154 286 155 287
rect 153 286 154 287
rect 152 286 153 287
rect 151 286 152 287
rect 150 286 151 287
rect 149 286 150 287
rect 148 286 149 287
rect 147 286 148 287
rect 146 286 147 287
rect 145 286 146 287
rect 144 286 145 287
rect 143 286 144 287
rect 142 286 143 287
rect 141 286 142 287
rect 140 286 141 287
rect 139 286 140 287
rect 138 286 139 287
rect 137 286 138 287
rect 136 286 137 287
rect 135 286 136 287
rect 134 286 135 287
rect 133 286 134 287
rect 132 286 133 287
rect 131 286 132 287
rect 115 286 116 287
rect 114 286 115 287
rect 113 286 114 287
rect 112 286 113 287
rect 111 286 112 287
rect 110 286 111 287
rect 109 286 110 287
rect 108 286 109 287
rect 107 286 108 287
rect 106 286 107 287
rect 105 286 106 287
rect 104 286 105 287
rect 103 286 104 287
rect 102 286 103 287
rect 101 286 102 287
rect 100 286 101 287
rect 99 286 100 287
rect 98 286 99 287
rect 97 286 98 287
rect 96 286 97 287
rect 95 286 96 287
rect 94 286 95 287
rect 93 286 94 287
rect 92 286 93 287
rect 91 286 92 287
rect 90 286 91 287
rect 89 286 90 287
rect 88 286 89 287
rect 87 286 88 287
rect 86 286 87 287
rect 85 286 86 287
rect 84 286 85 287
rect 83 286 84 287
rect 82 286 83 287
rect 81 286 82 287
rect 80 286 81 287
rect 64 286 65 287
rect 63 286 64 287
rect 62 286 63 287
rect 61 286 62 287
rect 60 286 61 287
rect 59 286 60 287
rect 58 286 59 287
rect 57 286 58 287
rect 56 286 57 287
rect 55 286 56 287
rect 54 286 55 287
rect 53 286 54 287
rect 52 286 53 287
rect 51 286 52 287
rect 50 286 51 287
rect 49 286 50 287
rect 48 286 49 287
rect 47 286 48 287
rect 46 286 47 287
rect 45 286 46 287
rect 44 286 45 287
rect 43 286 44 287
rect 42 286 43 287
rect 41 286 42 287
rect 40 286 41 287
rect 39 286 40 287
rect 38 286 39 287
rect 37 286 38 287
rect 36 286 37 287
rect 27 286 28 287
rect 26 286 27 287
rect 25 286 26 287
rect 24 286 25 287
rect 23 286 24 287
rect 22 286 23 287
rect 21 286 22 287
rect 20 286 21 287
rect 19 286 20 287
rect 18 286 19 287
rect 17 286 18 287
rect 16 286 17 287
rect 15 286 16 287
rect 14 286 15 287
rect 13 286 14 287
rect 12 286 13 287
rect 11 286 12 287
rect 10 286 11 287
rect 9 286 10 287
rect 8 286 9 287
rect 7 286 8 287
rect 6 286 7 287
rect 5 286 6 287
rect 4 286 5 287
rect 3 286 4 287
rect 2 286 3 287
rect 1 286 2 287
rect 478 287 479 288
rect 458 287 459 288
rect 437 287 438 288
rect 436 287 437 288
rect 435 287 436 288
rect 434 287 435 288
rect 433 287 434 288
rect 432 287 433 288
rect 416 287 417 288
rect 415 287 416 288
rect 414 287 415 288
rect 413 287 414 288
rect 412 287 413 288
rect 399 287 400 288
rect 398 287 399 288
rect 397 287 398 288
rect 396 287 397 288
rect 395 287 396 288
rect 394 287 395 288
rect 393 287 394 288
rect 279 287 280 288
rect 278 287 279 288
rect 277 287 278 288
rect 276 287 277 288
rect 275 287 276 288
rect 274 287 275 288
rect 273 287 274 288
rect 272 287 273 288
rect 271 287 272 288
rect 270 287 271 288
rect 269 287 270 288
rect 268 287 269 288
rect 267 287 268 288
rect 266 287 267 288
rect 265 287 266 288
rect 264 287 265 288
rect 263 287 264 288
rect 262 287 263 288
rect 261 287 262 288
rect 260 287 261 288
rect 259 287 260 288
rect 258 287 259 288
rect 257 287 258 288
rect 256 287 257 288
rect 255 287 256 288
rect 254 287 255 288
rect 253 287 254 288
rect 252 287 253 288
rect 251 287 252 288
rect 250 287 251 288
rect 249 287 250 288
rect 248 287 249 288
rect 247 287 248 288
rect 246 287 247 288
rect 245 287 246 288
rect 244 287 245 288
rect 243 287 244 288
rect 242 287 243 288
rect 241 287 242 288
rect 240 287 241 288
rect 239 287 240 288
rect 238 287 239 288
rect 237 287 238 288
rect 236 287 237 288
rect 235 287 236 288
rect 234 287 235 288
rect 233 287 234 288
rect 232 287 233 288
rect 231 287 232 288
rect 230 287 231 288
rect 229 287 230 288
rect 228 287 229 288
rect 227 287 228 288
rect 226 287 227 288
rect 225 287 226 288
rect 224 287 225 288
rect 223 287 224 288
rect 222 287 223 288
rect 221 287 222 288
rect 220 287 221 288
rect 219 287 220 288
rect 218 287 219 288
rect 217 287 218 288
rect 216 287 217 288
rect 215 287 216 288
rect 214 287 215 288
rect 213 287 214 288
rect 190 287 191 288
rect 189 287 190 288
rect 188 287 189 288
rect 187 287 188 288
rect 186 287 187 288
rect 185 287 186 288
rect 184 287 185 288
rect 183 287 184 288
rect 182 287 183 288
rect 181 287 182 288
rect 180 287 181 288
rect 179 287 180 288
rect 178 287 179 288
rect 177 287 178 288
rect 176 287 177 288
rect 175 287 176 288
rect 174 287 175 288
rect 173 287 174 288
rect 172 287 173 288
rect 171 287 172 288
rect 170 287 171 288
rect 169 287 170 288
rect 168 287 169 288
rect 167 287 168 288
rect 166 287 167 288
rect 165 287 166 288
rect 164 287 165 288
rect 163 287 164 288
rect 162 287 163 288
rect 161 287 162 288
rect 160 287 161 288
rect 159 287 160 288
rect 158 287 159 288
rect 157 287 158 288
rect 156 287 157 288
rect 155 287 156 288
rect 154 287 155 288
rect 153 287 154 288
rect 152 287 153 288
rect 151 287 152 288
rect 150 287 151 288
rect 149 287 150 288
rect 148 287 149 288
rect 147 287 148 288
rect 146 287 147 288
rect 145 287 146 288
rect 144 287 145 288
rect 143 287 144 288
rect 142 287 143 288
rect 141 287 142 288
rect 140 287 141 288
rect 139 287 140 288
rect 138 287 139 288
rect 137 287 138 288
rect 136 287 137 288
rect 135 287 136 288
rect 134 287 135 288
rect 133 287 134 288
rect 132 287 133 288
rect 115 287 116 288
rect 114 287 115 288
rect 113 287 114 288
rect 112 287 113 288
rect 111 287 112 288
rect 110 287 111 288
rect 109 287 110 288
rect 108 287 109 288
rect 107 287 108 288
rect 106 287 107 288
rect 105 287 106 288
rect 104 287 105 288
rect 103 287 104 288
rect 102 287 103 288
rect 101 287 102 288
rect 100 287 101 288
rect 99 287 100 288
rect 98 287 99 288
rect 97 287 98 288
rect 96 287 97 288
rect 95 287 96 288
rect 94 287 95 288
rect 93 287 94 288
rect 92 287 93 288
rect 91 287 92 288
rect 90 287 91 288
rect 89 287 90 288
rect 88 287 89 288
rect 87 287 88 288
rect 86 287 87 288
rect 85 287 86 288
rect 84 287 85 288
rect 83 287 84 288
rect 82 287 83 288
rect 81 287 82 288
rect 65 287 66 288
rect 64 287 65 288
rect 63 287 64 288
rect 62 287 63 288
rect 61 287 62 288
rect 60 287 61 288
rect 59 287 60 288
rect 58 287 59 288
rect 57 287 58 288
rect 56 287 57 288
rect 55 287 56 288
rect 54 287 55 288
rect 53 287 54 288
rect 52 287 53 288
rect 51 287 52 288
rect 50 287 51 288
rect 49 287 50 288
rect 48 287 49 288
rect 47 287 48 288
rect 46 287 47 288
rect 45 287 46 288
rect 44 287 45 288
rect 43 287 44 288
rect 42 287 43 288
rect 41 287 42 288
rect 40 287 41 288
rect 39 287 40 288
rect 38 287 39 288
rect 37 287 38 288
rect 36 287 37 288
rect 27 287 28 288
rect 26 287 27 288
rect 25 287 26 288
rect 24 287 25 288
rect 23 287 24 288
rect 22 287 23 288
rect 21 287 22 288
rect 20 287 21 288
rect 19 287 20 288
rect 18 287 19 288
rect 17 287 18 288
rect 16 287 17 288
rect 15 287 16 288
rect 14 287 15 288
rect 13 287 14 288
rect 12 287 13 288
rect 11 287 12 288
rect 10 287 11 288
rect 9 287 10 288
rect 8 287 9 288
rect 7 287 8 288
rect 6 287 7 288
rect 5 287 6 288
rect 4 287 5 288
rect 3 287 4 288
rect 2 287 3 288
rect 1 287 2 288
rect 478 288 479 289
rect 458 288 459 289
rect 437 288 438 289
rect 436 288 437 289
rect 435 288 436 289
rect 434 288 435 289
rect 415 288 416 289
rect 414 288 415 289
rect 413 288 414 289
rect 412 288 413 289
rect 396 288 397 289
rect 395 288 396 289
rect 394 288 395 289
rect 393 288 394 289
rect 278 288 279 289
rect 277 288 278 289
rect 276 288 277 289
rect 275 288 276 289
rect 274 288 275 289
rect 273 288 274 289
rect 272 288 273 289
rect 271 288 272 289
rect 270 288 271 289
rect 269 288 270 289
rect 268 288 269 289
rect 267 288 268 289
rect 266 288 267 289
rect 265 288 266 289
rect 264 288 265 289
rect 263 288 264 289
rect 262 288 263 289
rect 261 288 262 289
rect 260 288 261 289
rect 259 288 260 289
rect 258 288 259 289
rect 257 288 258 289
rect 256 288 257 289
rect 255 288 256 289
rect 254 288 255 289
rect 253 288 254 289
rect 252 288 253 289
rect 251 288 252 289
rect 250 288 251 289
rect 249 288 250 289
rect 248 288 249 289
rect 247 288 248 289
rect 246 288 247 289
rect 245 288 246 289
rect 244 288 245 289
rect 243 288 244 289
rect 242 288 243 289
rect 241 288 242 289
rect 240 288 241 289
rect 239 288 240 289
rect 238 288 239 289
rect 237 288 238 289
rect 236 288 237 289
rect 235 288 236 289
rect 234 288 235 289
rect 233 288 234 289
rect 232 288 233 289
rect 231 288 232 289
rect 230 288 231 289
rect 229 288 230 289
rect 228 288 229 289
rect 227 288 228 289
rect 226 288 227 289
rect 225 288 226 289
rect 224 288 225 289
rect 223 288 224 289
rect 222 288 223 289
rect 221 288 222 289
rect 220 288 221 289
rect 219 288 220 289
rect 218 288 219 289
rect 217 288 218 289
rect 216 288 217 289
rect 215 288 216 289
rect 214 288 215 289
rect 213 288 214 289
rect 189 288 190 289
rect 188 288 189 289
rect 187 288 188 289
rect 186 288 187 289
rect 185 288 186 289
rect 184 288 185 289
rect 183 288 184 289
rect 182 288 183 289
rect 181 288 182 289
rect 180 288 181 289
rect 179 288 180 289
rect 178 288 179 289
rect 177 288 178 289
rect 176 288 177 289
rect 175 288 176 289
rect 174 288 175 289
rect 173 288 174 289
rect 172 288 173 289
rect 171 288 172 289
rect 170 288 171 289
rect 169 288 170 289
rect 168 288 169 289
rect 167 288 168 289
rect 166 288 167 289
rect 165 288 166 289
rect 164 288 165 289
rect 163 288 164 289
rect 162 288 163 289
rect 161 288 162 289
rect 160 288 161 289
rect 159 288 160 289
rect 158 288 159 289
rect 157 288 158 289
rect 156 288 157 289
rect 155 288 156 289
rect 154 288 155 289
rect 153 288 154 289
rect 152 288 153 289
rect 151 288 152 289
rect 150 288 151 289
rect 149 288 150 289
rect 148 288 149 289
rect 147 288 148 289
rect 146 288 147 289
rect 145 288 146 289
rect 144 288 145 289
rect 143 288 144 289
rect 142 288 143 289
rect 141 288 142 289
rect 140 288 141 289
rect 139 288 140 289
rect 138 288 139 289
rect 137 288 138 289
rect 136 288 137 289
rect 135 288 136 289
rect 134 288 135 289
rect 133 288 134 289
rect 116 288 117 289
rect 115 288 116 289
rect 114 288 115 289
rect 113 288 114 289
rect 112 288 113 289
rect 111 288 112 289
rect 110 288 111 289
rect 109 288 110 289
rect 108 288 109 289
rect 107 288 108 289
rect 106 288 107 289
rect 105 288 106 289
rect 104 288 105 289
rect 103 288 104 289
rect 102 288 103 289
rect 101 288 102 289
rect 100 288 101 289
rect 99 288 100 289
rect 98 288 99 289
rect 97 288 98 289
rect 96 288 97 289
rect 95 288 96 289
rect 94 288 95 289
rect 93 288 94 289
rect 92 288 93 289
rect 91 288 92 289
rect 90 288 91 289
rect 89 288 90 289
rect 88 288 89 289
rect 87 288 88 289
rect 86 288 87 289
rect 85 288 86 289
rect 84 288 85 289
rect 83 288 84 289
rect 82 288 83 289
rect 81 288 82 289
rect 65 288 66 289
rect 64 288 65 289
rect 63 288 64 289
rect 62 288 63 289
rect 61 288 62 289
rect 60 288 61 289
rect 59 288 60 289
rect 58 288 59 289
rect 57 288 58 289
rect 56 288 57 289
rect 55 288 56 289
rect 54 288 55 289
rect 53 288 54 289
rect 52 288 53 289
rect 51 288 52 289
rect 50 288 51 289
rect 49 288 50 289
rect 48 288 49 289
rect 47 288 48 289
rect 46 288 47 289
rect 45 288 46 289
rect 44 288 45 289
rect 43 288 44 289
rect 42 288 43 289
rect 41 288 42 289
rect 40 288 41 289
rect 39 288 40 289
rect 38 288 39 289
rect 37 288 38 289
rect 36 288 37 289
rect 27 288 28 289
rect 26 288 27 289
rect 25 288 26 289
rect 24 288 25 289
rect 23 288 24 289
rect 22 288 23 289
rect 21 288 22 289
rect 20 288 21 289
rect 19 288 20 289
rect 18 288 19 289
rect 17 288 18 289
rect 16 288 17 289
rect 15 288 16 289
rect 14 288 15 289
rect 13 288 14 289
rect 12 288 13 289
rect 11 288 12 289
rect 10 288 11 289
rect 9 288 10 289
rect 8 288 9 289
rect 7 288 8 289
rect 6 288 7 289
rect 5 288 6 289
rect 4 288 5 289
rect 3 288 4 289
rect 2 288 3 289
rect 1 288 2 289
rect 478 289 479 290
rect 477 289 478 290
rect 458 289 459 290
rect 437 289 438 290
rect 436 289 437 290
rect 435 289 436 290
rect 415 289 416 290
rect 414 289 415 290
rect 413 289 414 290
rect 412 289 413 290
rect 395 289 396 290
rect 394 289 395 290
rect 393 289 394 290
rect 277 289 278 290
rect 276 289 277 290
rect 275 289 276 290
rect 274 289 275 290
rect 273 289 274 290
rect 272 289 273 290
rect 271 289 272 290
rect 270 289 271 290
rect 269 289 270 290
rect 268 289 269 290
rect 267 289 268 290
rect 266 289 267 290
rect 265 289 266 290
rect 264 289 265 290
rect 263 289 264 290
rect 262 289 263 290
rect 261 289 262 290
rect 260 289 261 290
rect 259 289 260 290
rect 258 289 259 290
rect 257 289 258 290
rect 256 289 257 290
rect 255 289 256 290
rect 254 289 255 290
rect 253 289 254 290
rect 252 289 253 290
rect 251 289 252 290
rect 250 289 251 290
rect 249 289 250 290
rect 248 289 249 290
rect 247 289 248 290
rect 246 289 247 290
rect 245 289 246 290
rect 244 289 245 290
rect 243 289 244 290
rect 242 289 243 290
rect 241 289 242 290
rect 240 289 241 290
rect 239 289 240 290
rect 238 289 239 290
rect 237 289 238 290
rect 236 289 237 290
rect 235 289 236 290
rect 234 289 235 290
rect 233 289 234 290
rect 232 289 233 290
rect 231 289 232 290
rect 230 289 231 290
rect 229 289 230 290
rect 228 289 229 290
rect 227 289 228 290
rect 226 289 227 290
rect 225 289 226 290
rect 224 289 225 290
rect 223 289 224 290
rect 222 289 223 290
rect 221 289 222 290
rect 220 289 221 290
rect 219 289 220 290
rect 218 289 219 290
rect 217 289 218 290
rect 216 289 217 290
rect 215 289 216 290
rect 214 289 215 290
rect 213 289 214 290
rect 212 289 213 290
rect 189 289 190 290
rect 188 289 189 290
rect 187 289 188 290
rect 186 289 187 290
rect 185 289 186 290
rect 184 289 185 290
rect 183 289 184 290
rect 182 289 183 290
rect 181 289 182 290
rect 180 289 181 290
rect 179 289 180 290
rect 178 289 179 290
rect 177 289 178 290
rect 176 289 177 290
rect 175 289 176 290
rect 174 289 175 290
rect 173 289 174 290
rect 172 289 173 290
rect 171 289 172 290
rect 170 289 171 290
rect 169 289 170 290
rect 168 289 169 290
rect 167 289 168 290
rect 166 289 167 290
rect 165 289 166 290
rect 164 289 165 290
rect 163 289 164 290
rect 162 289 163 290
rect 161 289 162 290
rect 160 289 161 290
rect 159 289 160 290
rect 158 289 159 290
rect 157 289 158 290
rect 156 289 157 290
rect 155 289 156 290
rect 154 289 155 290
rect 153 289 154 290
rect 152 289 153 290
rect 151 289 152 290
rect 150 289 151 290
rect 149 289 150 290
rect 148 289 149 290
rect 147 289 148 290
rect 146 289 147 290
rect 145 289 146 290
rect 144 289 145 290
rect 143 289 144 290
rect 142 289 143 290
rect 141 289 142 290
rect 140 289 141 290
rect 139 289 140 290
rect 138 289 139 290
rect 137 289 138 290
rect 136 289 137 290
rect 135 289 136 290
rect 134 289 135 290
rect 133 289 134 290
rect 116 289 117 290
rect 115 289 116 290
rect 114 289 115 290
rect 113 289 114 290
rect 112 289 113 290
rect 111 289 112 290
rect 110 289 111 290
rect 109 289 110 290
rect 108 289 109 290
rect 107 289 108 290
rect 106 289 107 290
rect 105 289 106 290
rect 104 289 105 290
rect 103 289 104 290
rect 102 289 103 290
rect 101 289 102 290
rect 100 289 101 290
rect 99 289 100 290
rect 98 289 99 290
rect 97 289 98 290
rect 96 289 97 290
rect 95 289 96 290
rect 94 289 95 290
rect 93 289 94 290
rect 92 289 93 290
rect 91 289 92 290
rect 90 289 91 290
rect 89 289 90 290
rect 88 289 89 290
rect 87 289 88 290
rect 86 289 87 290
rect 85 289 86 290
rect 84 289 85 290
rect 83 289 84 290
rect 82 289 83 290
rect 81 289 82 290
rect 65 289 66 290
rect 64 289 65 290
rect 63 289 64 290
rect 62 289 63 290
rect 61 289 62 290
rect 60 289 61 290
rect 59 289 60 290
rect 58 289 59 290
rect 57 289 58 290
rect 56 289 57 290
rect 55 289 56 290
rect 54 289 55 290
rect 53 289 54 290
rect 52 289 53 290
rect 51 289 52 290
rect 50 289 51 290
rect 49 289 50 290
rect 48 289 49 290
rect 47 289 48 290
rect 46 289 47 290
rect 45 289 46 290
rect 44 289 45 290
rect 43 289 44 290
rect 42 289 43 290
rect 41 289 42 290
rect 40 289 41 290
rect 39 289 40 290
rect 38 289 39 290
rect 37 289 38 290
rect 36 289 37 290
rect 27 289 28 290
rect 26 289 27 290
rect 25 289 26 290
rect 24 289 25 290
rect 23 289 24 290
rect 22 289 23 290
rect 21 289 22 290
rect 20 289 21 290
rect 19 289 20 290
rect 18 289 19 290
rect 17 289 18 290
rect 16 289 17 290
rect 15 289 16 290
rect 14 289 15 290
rect 13 289 14 290
rect 12 289 13 290
rect 11 289 12 290
rect 10 289 11 290
rect 9 289 10 290
rect 8 289 9 290
rect 7 289 8 290
rect 6 289 7 290
rect 5 289 6 290
rect 4 289 5 290
rect 3 289 4 290
rect 2 289 3 290
rect 1 289 2 290
rect 478 290 479 291
rect 477 290 478 291
rect 476 290 477 291
rect 475 290 476 291
rect 474 290 475 291
rect 473 290 474 291
rect 472 290 473 291
rect 471 290 472 291
rect 470 290 471 291
rect 469 290 470 291
rect 468 290 469 291
rect 467 290 468 291
rect 466 290 467 291
rect 465 290 466 291
rect 464 290 465 291
rect 463 290 464 291
rect 462 290 463 291
rect 461 290 462 291
rect 460 290 461 291
rect 459 290 460 291
rect 458 290 459 291
rect 437 290 438 291
rect 436 290 437 291
rect 435 290 436 291
rect 415 290 416 291
rect 414 290 415 291
rect 413 290 414 291
rect 412 290 413 291
rect 395 290 396 291
rect 394 290 395 291
rect 393 290 394 291
rect 276 290 277 291
rect 275 290 276 291
rect 274 290 275 291
rect 273 290 274 291
rect 272 290 273 291
rect 271 290 272 291
rect 270 290 271 291
rect 269 290 270 291
rect 268 290 269 291
rect 267 290 268 291
rect 266 290 267 291
rect 265 290 266 291
rect 264 290 265 291
rect 263 290 264 291
rect 262 290 263 291
rect 261 290 262 291
rect 260 290 261 291
rect 259 290 260 291
rect 258 290 259 291
rect 257 290 258 291
rect 256 290 257 291
rect 255 290 256 291
rect 254 290 255 291
rect 253 290 254 291
rect 252 290 253 291
rect 251 290 252 291
rect 250 290 251 291
rect 249 290 250 291
rect 248 290 249 291
rect 247 290 248 291
rect 246 290 247 291
rect 245 290 246 291
rect 244 290 245 291
rect 243 290 244 291
rect 242 290 243 291
rect 241 290 242 291
rect 240 290 241 291
rect 239 290 240 291
rect 238 290 239 291
rect 237 290 238 291
rect 236 290 237 291
rect 235 290 236 291
rect 234 290 235 291
rect 233 290 234 291
rect 232 290 233 291
rect 231 290 232 291
rect 230 290 231 291
rect 229 290 230 291
rect 228 290 229 291
rect 227 290 228 291
rect 226 290 227 291
rect 225 290 226 291
rect 224 290 225 291
rect 223 290 224 291
rect 222 290 223 291
rect 221 290 222 291
rect 220 290 221 291
rect 219 290 220 291
rect 218 290 219 291
rect 217 290 218 291
rect 216 290 217 291
rect 215 290 216 291
rect 214 290 215 291
rect 213 290 214 291
rect 212 290 213 291
rect 211 290 212 291
rect 188 290 189 291
rect 187 290 188 291
rect 186 290 187 291
rect 185 290 186 291
rect 184 290 185 291
rect 183 290 184 291
rect 182 290 183 291
rect 181 290 182 291
rect 180 290 181 291
rect 179 290 180 291
rect 178 290 179 291
rect 177 290 178 291
rect 176 290 177 291
rect 175 290 176 291
rect 174 290 175 291
rect 173 290 174 291
rect 172 290 173 291
rect 171 290 172 291
rect 170 290 171 291
rect 169 290 170 291
rect 168 290 169 291
rect 167 290 168 291
rect 166 290 167 291
rect 165 290 166 291
rect 164 290 165 291
rect 163 290 164 291
rect 162 290 163 291
rect 161 290 162 291
rect 160 290 161 291
rect 159 290 160 291
rect 158 290 159 291
rect 157 290 158 291
rect 156 290 157 291
rect 155 290 156 291
rect 154 290 155 291
rect 153 290 154 291
rect 152 290 153 291
rect 151 290 152 291
rect 150 290 151 291
rect 149 290 150 291
rect 148 290 149 291
rect 147 290 148 291
rect 146 290 147 291
rect 145 290 146 291
rect 144 290 145 291
rect 143 290 144 291
rect 142 290 143 291
rect 141 290 142 291
rect 140 290 141 291
rect 139 290 140 291
rect 138 290 139 291
rect 137 290 138 291
rect 136 290 137 291
rect 135 290 136 291
rect 134 290 135 291
rect 116 290 117 291
rect 115 290 116 291
rect 114 290 115 291
rect 113 290 114 291
rect 112 290 113 291
rect 111 290 112 291
rect 110 290 111 291
rect 109 290 110 291
rect 108 290 109 291
rect 107 290 108 291
rect 106 290 107 291
rect 105 290 106 291
rect 104 290 105 291
rect 103 290 104 291
rect 102 290 103 291
rect 101 290 102 291
rect 100 290 101 291
rect 99 290 100 291
rect 98 290 99 291
rect 97 290 98 291
rect 96 290 97 291
rect 95 290 96 291
rect 94 290 95 291
rect 93 290 94 291
rect 92 290 93 291
rect 91 290 92 291
rect 90 290 91 291
rect 89 290 90 291
rect 88 290 89 291
rect 87 290 88 291
rect 86 290 87 291
rect 85 290 86 291
rect 84 290 85 291
rect 83 290 84 291
rect 82 290 83 291
rect 81 290 82 291
rect 65 290 66 291
rect 64 290 65 291
rect 63 290 64 291
rect 62 290 63 291
rect 61 290 62 291
rect 60 290 61 291
rect 59 290 60 291
rect 58 290 59 291
rect 57 290 58 291
rect 56 290 57 291
rect 55 290 56 291
rect 54 290 55 291
rect 53 290 54 291
rect 52 290 53 291
rect 51 290 52 291
rect 50 290 51 291
rect 49 290 50 291
rect 48 290 49 291
rect 47 290 48 291
rect 46 290 47 291
rect 45 290 46 291
rect 44 290 45 291
rect 43 290 44 291
rect 42 290 43 291
rect 41 290 42 291
rect 40 290 41 291
rect 39 290 40 291
rect 38 290 39 291
rect 37 290 38 291
rect 27 290 28 291
rect 26 290 27 291
rect 25 290 26 291
rect 24 290 25 291
rect 23 290 24 291
rect 22 290 23 291
rect 21 290 22 291
rect 20 290 21 291
rect 19 290 20 291
rect 18 290 19 291
rect 17 290 18 291
rect 16 290 17 291
rect 15 290 16 291
rect 14 290 15 291
rect 13 290 14 291
rect 12 290 13 291
rect 11 290 12 291
rect 10 290 11 291
rect 9 290 10 291
rect 8 290 9 291
rect 7 290 8 291
rect 6 290 7 291
rect 5 290 6 291
rect 4 290 5 291
rect 3 290 4 291
rect 2 290 3 291
rect 1 290 2 291
rect 478 291 479 292
rect 477 291 478 292
rect 476 291 477 292
rect 475 291 476 292
rect 474 291 475 292
rect 473 291 474 292
rect 472 291 473 292
rect 471 291 472 292
rect 470 291 471 292
rect 469 291 470 292
rect 468 291 469 292
rect 467 291 468 292
rect 466 291 467 292
rect 465 291 466 292
rect 464 291 465 292
rect 463 291 464 292
rect 462 291 463 292
rect 461 291 462 292
rect 460 291 461 292
rect 459 291 460 292
rect 458 291 459 292
rect 437 291 438 292
rect 436 291 437 292
rect 435 291 436 292
rect 415 291 416 292
rect 414 291 415 292
rect 413 291 414 292
rect 412 291 413 292
rect 395 291 396 292
rect 394 291 395 292
rect 393 291 394 292
rect 275 291 276 292
rect 274 291 275 292
rect 273 291 274 292
rect 272 291 273 292
rect 271 291 272 292
rect 270 291 271 292
rect 269 291 270 292
rect 268 291 269 292
rect 267 291 268 292
rect 266 291 267 292
rect 265 291 266 292
rect 264 291 265 292
rect 263 291 264 292
rect 262 291 263 292
rect 261 291 262 292
rect 260 291 261 292
rect 259 291 260 292
rect 258 291 259 292
rect 257 291 258 292
rect 256 291 257 292
rect 255 291 256 292
rect 254 291 255 292
rect 253 291 254 292
rect 252 291 253 292
rect 251 291 252 292
rect 250 291 251 292
rect 249 291 250 292
rect 248 291 249 292
rect 247 291 248 292
rect 246 291 247 292
rect 245 291 246 292
rect 244 291 245 292
rect 243 291 244 292
rect 242 291 243 292
rect 241 291 242 292
rect 240 291 241 292
rect 239 291 240 292
rect 238 291 239 292
rect 237 291 238 292
rect 236 291 237 292
rect 235 291 236 292
rect 234 291 235 292
rect 233 291 234 292
rect 232 291 233 292
rect 231 291 232 292
rect 230 291 231 292
rect 229 291 230 292
rect 228 291 229 292
rect 227 291 228 292
rect 226 291 227 292
rect 225 291 226 292
rect 224 291 225 292
rect 223 291 224 292
rect 222 291 223 292
rect 221 291 222 292
rect 220 291 221 292
rect 219 291 220 292
rect 218 291 219 292
rect 217 291 218 292
rect 216 291 217 292
rect 215 291 216 292
rect 214 291 215 292
rect 213 291 214 292
rect 212 291 213 292
rect 211 291 212 292
rect 187 291 188 292
rect 186 291 187 292
rect 185 291 186 292
rect 184 291 185 292
rect 183 291 184 292
rect 182 291 183 292
rect 181 291 182 292
rect 180 291 181 292
rect 179 291 180 292
rect 178 291 179 292
rect 177 291 178 292
rect 176 291 177 292
rect 175 291 176 292
rect 174 291 175 292
rect 173 291 174 292
rect 172 291 173 292
rect 171 291 172 292
rect 170 291 171 292
rect 169 291 170 292
rect 168 291 169 292
rect 167 291 168 292
rect 166 291 167 292
rect 165 291 166 292
rect 164 291 165 292
rect 163 291 164 292
rect 162 291 163 292
rect 161 291 162 292
rect 160 291 161 292
rect 159 291 160 292
rect 158 291 159 292
rect 157 291 158 292
rect 156 291 157 292
rect 155 291 156 292
rect 154 291 155 292
rect 153 291 154 292
rect 152 291 153 292
rect 151 291 152 292
rect 150 291 151 292
rect 149 291 150 292
rect 148 291 149 292
rect 147 291 148 292
rect 146 291 147 292
rect 145 291 146 292
rect 144 291 145 292
rect 143 291 144 292
rect 142 291 143 292
rect 141 291 142 292
rect 140 291 141 292
rect 139 291 140 292
rect 138 291 139 292
rect 137 291 138 292
rect 136 291 137 292
rect 135 291 136 292
rect 117 291 118 292
rect 116 291 117 292
rect 115 291 116 292
rect 114 291 115 292
rect 113 291 114 292
rect 112 291 113 292
rect 111 291 112 292
rect 110 291 111 292
rect 109 291 110 292
rect 108 291 109 292
rect 107 291 108 292
rect 106 291 107 292
rect 105 291 106 292
rect 104 291 105 292
rect 103 291 104 292
rect 102 291 103 292
rect 101 291 102 292
rect 100 291 101 292
rect 99 291 100 292
rect 98 291 99 292
rect 97 291 98 292
rect 96 291 97 292
rect 95 291 96 292
rect 94 291 95 292
rect 93 291 94 292
rect 92 291 93 292
rect 91 291 92 292
rect 90 291 91 292
rect 89 291 90 292
rect 88 291 89 292
rect 87 291 88 292
rect 86 291 87 292
rect 85 291 86 292
rect 84 291 85 292
rect 83 291 84 292
rect 82 291 83 292
rect 66 291 67 292
rect 65 291 66 292
rect 64 291 65 292
rect 63 291 64 292
rect 62 291 63 292
rect 61 291 62 292
rect 60 291 61 292
rect 59 291 60 292
rect 58 291 59 292
rect 57 291 58 292
rect 56 291 57 292
rect 55 291 56 292
rect 54 291 55 292
rect 53 291 54 292
rect 52 291 53 292
rect 51 291 52 292
rect 50 291 51 292
rect 49 291 50 292
rect 48 291 49 292
rect 47 291 48 292
rect 46 291 47 292
rect 45 291 46 292
rect 44 291 45 292
rect 43 291 44 292
rect 42 291 43 292
rect 41 291 42 292
rect 40 291 41 292
rect 39 291 40 292
rect 38 291 39 292
rect 37 291 38 292
rect 27 291 28 292
rect 26 291 27 292
rect 25 291 26 292
rect 24 291 25 292
rect 23 291 24 292
rect 22 291 23 292
rect 21 291 22 292
rect 20 291 21 292
rect 19 291 20 292
rect 18 291 19 292
rect 17 291 18 292
rect 16 291 17 292
rect 15 291 16 292
rect 14 291 15 292
rect 13 291 14 292
rect 12 291 13 292
rect 11 291 12 292
rect 10 291 11 292
rect 9 291 10 292
rect 8 291 9 292
rect 7 291 8 292
rect 6 291 7 292
rect 5 291 6 292
rect 4 291 5 292
rect 3 291 4 292
rect 2 291 3 292
rect 1 291 2 292
rect 478 292 479 293
rect 477 292 478 293
rect 476 292 477 293
rect 475 292 476 293
rect 474 292 475 293
rect 473 292 474 293
rect 472 292 473 293
rect 471 292 472 293
rect 470 292 471 293
rect 469 292 470 293
rect 468 292 469 293
rect 467 292 468 293
rect 466 292 467 293
rect 465 292 466 293
rect 464 292 465 293
rect 463 292 464 293
rect 462 292 463 293
rect 461 292 462 293
rect 460 292 461 293
rect 459 292 460 293
rect 458 292 459 293
rect 437 292 438 293
rect 436 292 437 293
rect 415 292 416 293
rect 414 292 415 293
rect 413 292 414 293
rect 412 292 413 293
rect 395 292 396 293
rect 394 292 395 293
rect 393 292 394 293
rect 274 292 275 293
rect 273 292 274 293
rect 272 292 273 293
rect 271 292 272 293
rect 270 292 271 293
rect 269 292 270 293
rect 268 292 269 293
rect 267 292 268 293
rect 266 292 267 293
rect 265 292 266 293
rect 264 292 265 293
rect 263 292 264 293
rect 262 292 263 293
rect 261 292 262 293
rect 260 292 261 293
rect 259 292 260 293
rect 258 292 259 293
rect 257 292 258 293
rect 256 292 257 293
rect 255 292 256 293
rect 254 292 255 293
rect 253 292 254 293
rect 252 292 253 293
rect 251 292 252 293
rect 250 292 251 293
rect 249 292 250 293
rect 248 292 249 293
rect 247 292 248 293
rect 246 292 247 293
rect 245 292 246 293
rect 244 292 245 293
rect 243 292 244 293
rect 242 292 243 293
rect 241 292 242 293
rect 240 292 241 293
rect 239 292 240 293
rect 238 292 239 293
rect 237 292 238 293
rect 236 292 237 293
rect 235 292 236 293
rect 234 292 235 293
rect 233 292 234 293
rect 232 292 233 293
rect 231 292 232 293
rect 230 292 231 293
rect 229 292 230 293
rect 228 292 229 293
rect 227 292 228 293
rect 226 292 227 293
rect 225 292 226 293
rect 224 292 225 293
rect 223 292 224 293
rect 222 292 223 293
rect 221 292 222 293
rect 220 292 221 293
rect 219 292 220 293
rect 218 292 219 293
rect 217 292 218 293
rect 216 292 217 293
rect 215 292 216 293
rect 214 292 215 293
rect 213 292 214 293
rect 212 292 213 293
rect 211 292 212 293
rect 210 292 211 293
rect 186 292 187 293
rect 185 292 186 293
rect 184 292 185 293
rect 183 292 184 293
rect 182 292 183 293
rect 181 292 182 293
rect 180 292 181 293
rect 179 292 180 293
rect 178 292 179 293
rect 177 292 178 293
rect 176 292 177 293
rect 175 292 176 293
rect 174 292 175 293
rect 173 292 174 293
rect 172 292 173 293
rect 171 292 172 293
rect 170 292 171 293
rect 169 292 170 293
rect 168 292 169 293
rect 167 292 168 293
rect 166 292 167 293
rect 165 292 166 293
rect 164 292 165 293
rect 163 292 164 293
rect 162 292 163 293
rect 161 292 162 293
rect 160 292 161 293
rect 159 292 160 293
rect 158 292 159 293
rect 157 292 158 293
rect 156 292 157 293
rect 155 292 156 293
rect 154 292 155 293
rect 153 292 154 293
rect 152 292 153 293
rect 151 292 152 293
rect 150 292 151 293
rect 149 292 150 293
rect 148 292 149 293
rect 147 292 148 293
rect 146 292 147 293
rect 145 292 146 293
rect 144 292 145 293
rect 143 292 144 293
rect 142 292 143 293
rect 141 292 142 293
rect 140 292 141 293
rect 139 292 140 293
rect 138 292 139 293
rect 137 292 138 293
rect 136 292 137 293
rect 117 292 118 293
rect 116 292 117 293
rect 115 292 116 293
rect 114 292 115 293
rect 113 292 114 293
rect 112 292 113 293
rect 111 292 112 293
rect 110 292 111 293
rect 109 292 110 293
rect 108 292 109 293
rect 107 292 108 293
rect 106 292 107 293
rect 105 292 106 293
rect 104 292 105 293
rect 103 292 104 293
rect 102 292 103 293
rect 101 292 102 293
rect 100 292 101 293
rect 99 292 100 293
rect 98 292 99 293
rect 97 292 98 293
rect 96 292 97 293
rect 95 292 96 293
rect 94 292 95 293
rect 93 292 94 293
rect 92 292 93 293
rect 91 292 92 293
rect 90 292 91 293
rect 89 292 90 293
rect 88 292 89 293
rect 87 292 88 293
rect 86 292 87 293
rect 85 292 86 293
rect 84 292 85 293
rect 83 292 84 293
rect 82 292 83 293
rect 66 292 67 293
rect 65 292 66 293
rect 64 292 65 293
rect 63 292 64 293
rect 62 292 63 293
rect 61 292 62 293
rect 60 292 61 293
rect 59 292 60 293
rect 58 292 59 293
rect 57 292 58 293
rect 56 292 57 293
rect 55 292 56 293
rect 54 292 55 293
rect 53 292 54 293
rect 52 292 53 293
rect 51 292 52 293
rect 50 292 51 293
rect 49 292 50 293
rect 48 292 49 293
rect 47 292 48 293
rect 46 292 47 293
rect 45 292 46 293
rect 44 292 45 293
rect 43 292 44 293
rect 42 292 43 293
rect 41 292 42 293
rect 40 292 41 293
rect 39 292 40 293
rect 38 292 39 293
rect 37 292 38 293
rect 27 292 28 293
rect 26 292 27 293
rect 25 292 26 293
rect 24 292 25 293
rect 23 292 24 293
rect 22 292 23 293
rect 21 292 22 293
rect 20 292 21 293
rect 19 292 20 293
rect 18 292 19 293
rect 17 292 18 293
rect 16 292 17 293
rect 15 292 16 293
rect 14 292 15 293
rect 13 292 14 293
rect 12 292 13 293
rect 11 292 12 293
rect 10 292 11 293
rect 9 292 10 293
rect 8 292 9 293
rect 7 292 8 293
rect 6 292 7 293
rect 5 292 6 293
rect 4 292 5 293
rect 3 292 4 293
rect 2 292 3 293
rect 1 292 2 293
rect 478 293 479 294
rect 477 293 478 294
rect 476 293 477 294
rect 475 293 476 294
rect 474 293 475 294
rect 473 293 474 294
rect 472 293 473 294
rect 471 293 472 294
rect 470 293 471 294
rect 469 293 470 294
rect 468 293 469 294
rect 467 293 468 294
rect 466 293 467 294
rect 465 293 466 294
rect 464 293 465 294
rect 463 293 464 294
rect 462 293 463 294
rect 461 293 462 294
rect 460 293 461 294
rect 459 293 460 294
rect 458 293 459 294
rect 415 293 416 294
rect 414 293 415 294
rect 413 293 414 294
rect 412 293 413 294
rect 273 293 274 294
rect 272 293 273 294
rect 271 293 272 294
rect 270 293 271 294
rect 269 293 270 294
rect 268 293 269 294
rect 267 293 268 294
rect 266 293 267 294
rect 265 293 266 294
rect 264 293 265 294
rect 263 293 264 294
rect 262 293 263 294
rect 261 293 262 294
rect 260 293 261 294
rect 259 293 260 294
rect 258 293 259 294
rect 257 293 258 294
rect 256 293 257 294
rect 255 293 256 294
rect 254 293 255 294
rect 253 293 254 294
rect 252 293 253 294
rect 251 293 252 294
rect 250 293 251 294
rect 249 293 250 294
rect 248 293 249 294
rect 247 293 248 294
rect 246 293 247 294
rect 245 293 246 294
rect 244 293 245 294
rect 243 293 244 294
rect 242 293 243 294
rect 241 293 242 294
rect 240 293 241 294
rect 239 293 240 294
rect 238 293 239 294
rect 237 293 238 294
rect 236 293 237 294
rect 235 293 236 294
rect 234 293 235 294
rect 233 293 234 294
rect 232 293 233 294
rect 231 293 232 294
rect 230 293 231 294
rect 229 293 230 294
rect 228 293 229 294
rect 227 293 228 294
rect 226 293 227 294
rect 225 293 226 294
rect 224 293 225 294
rect 223 293 224 294
rect 222 293 223 294
rect 221 293 222 294
rect 220 293 221 294
rect 219 293 220 294
rect 218 293 219 294
rect 217 293 218 294
rect 216 293 217 294
rect 215 293 216 294
rect 214 293 215 294
rect 213 293 214 294
rect 212 293 213 294
rect 211 293 212 294
rect 210 293 211 294
rect 209 293 210 294
rect 185 293 186 294
rect 184 293 185 294
rect 183 293 184 294
rect 182 293 183 294
rect 181 293 182 294
rect 180 293 181 294
rect 179 293 180 294
rect 178 293 179 294
rect 177 293 178 294
rect 176 293 177 294
rect 175 293 176 294
rect 174 293 175 294
rect 173 293 174 294
rect 172 293 173 294
rect 171 293 172 294
rect 170 293 171 294
rect 169 293 170 294
rect 168 293 169 294
rect 167 293 168 294
rect 166 293 167 294
rect 165 293 166 294
rect 164 293 165 294
rect 163 293 164 294
rect 162 293 163 294
rect 161 293 162 294
rect 160 293 161 294
rect 159 293 160 294
rect 158 293 159 294
rect 157 293 158 294
rect 156 293 157 294
rect 155 293 156 294
rect 154 293 155 294
rect 153 293 154 294
rect 152 293 153 294
rect 151 293 152 294
rect 150 293 151 294
rect 149 293 150 294
rect 148 293 149 294
rect 147 293 148 294
rect 146 293 147 294
rect 145 293 146 294
rect 144 293 145 294
rect 143 293 144 294
rect 142 293 143 294
rect 141 293 142 294
rect 140 293 141 294
rect 139 293 140 294
rect 138 293 139 294
rect 137 293 138 294
rect 118 293 119 294
rect 117 293 118 294
rect 116 293 117 294
rect 115 293 116 294
rect 114 293 115 294
rect 113 293 114 294
rect 112 293 113 294
rect 111 293 112 294
rect 110 293 111 294
rect 109 293 110 294
rect 108 293 109 294
rect 107 293 108 294
rect 106 293 107 294
rect 105 293 106 294
rect 104 293 105 294
rect 103 293 104 294
rect 102 293 103 294
rect 101 293 102 294
rect 100 293 101 294
rect 99 293 100 294
rect 98 293 99 294
rect 97 293 98 294
rect 96 293 97 294
rect 95 293 96 294
rect 94 293 95 294
rect 93 293 94 294
rect 92 293 93 294
rect 91 293 92 294
rect 90 293 91 294
rect 89 293 90 294
rect 88 293 89 294
rect 87 293 88 294
rect 86 293 87 294
rect 85 293 86 294
rect 84 293 85 294
rect 83 293 84 294
rect 82 293 83 294
rect 66 293 67 294
rect 65 293 66 294
rect 64 293 65 294
rect 63 293 64 294
rect 62 293 63 294
rect 61 293 62 294
rect 60 293 61 294
rect 59 293 60 294
rect 58 293 59 294
rect 57 293 58 294
rect 56 293 57 294
rect 55 293 56 294
rect 54 293 55 294
rect 53 293 54 294
rect 52 293 53 294
rect 51 293 52 294
rect 50 293 51 294
rect 49 293 50 294
rect 48 293 49 294
rect 47 293 48 294
rect 46 293 47 294
rect 45 293 46 294
rect 44 293 45 294
rect 43 293 44 294
rect 42 293 43 294
rect 41 293 42 294
rect 40 293 41 294
rect 39 293 40 294
rect 38 293 39 294
rect 37 293 38 294
rect 27 293 28 294
rect 26 293 27 294
rect 25 293 26 294
rect 24 293 25 294
rect 23 293 24 294
rect 22 293 23 294
rect 21 293 22 294
rect 20 293 21 294
rect 19 293 20 294
rect 18 293 19 294
rect 17 293 18 294
rect 16 293 17 294
rect 15 293 16 294
rect 14 293 15 294
rect 13 293 14 294
rect 12 293 13 294
rect 11 293 12 294
rect 10 293 11 294
rect 9 293 10 294
rect 8 293 9 294
rect 7 293 8 294
rect 6 293 7 294
rect 5 293 6 294
rect 4 293 5 294
rect 3 293 4 294
rect 2 293 3 294
rect 1 293 2 294
rect 478 294 479 295
rect 477 294 478 295
rect 476 294 477 295
rect 475 294 476 295
rect 474 294 475 295
rect 473 294 474 295
rect 472 294 473 295
rect 471 294 472 295
rect 470 294 471 295
rect 469 294 470 295
rect 468 294 469 295
rect 467 294 468 295
rect 466 294 467 295
rect 465 294 466 295
rect 464 294 465 295
rect 463 294 464 295
rect 462 294 463 295
rect 461 294 462 295
rect 460 294 461 295
rect 459 294 460 295
rect 458 294 459 295
rect 415 294 416 295
rect 414 294 415 295
rect 413 294 414 295
rect 412 294 413 295
rect 271 294 272 295
rect 270 294 271 295
rect 269 294 270 295
rect 268 294 269 295
rect 267 294 268 295
rect 266 294 267 295
rect 265 294 266 295
rect 264 294 265 295
rect 263 294 264 295
rect 262 294 263 295
rect 261 294 262 295
rect 260 294 261 295
rect 259 294 260 295
rect 258 294 259 295
rect 257 294 258 295
rect 256 294 257 295
rect 255 294 256 295
rect 254 294 255 295
rect 253 294 254 295
rect 252 294 253 295
rect 251 294 252 295
rect 250 294 251 295
rect 249 294 250 295
rect 248 294 249 295
rect 247 294 248 295
rect 246 294 247 295
rect 245 294 246 295
rect 244 294 245 295
rect 243 294 244 295
rect 242 294 243 295
rect 241 294 242 295
rect 240 294 241 295
rect 239 294 240 295
rect 238 294 239 295
rect 237 294 238 295
rect 236 294 237 295
rect 235 294 236 295
rect 234 294 235 295
rect 233 294 234 295
rect 232 294 233 295
rect 231 294 232 295
rect 230 294 231 295
rect 229 294 230 295
rect 228 294 229 295
rect 227 294 228 295
rect 226 294 227 295
rect 225 294 226 295
rect 224 294 225 295
rect 223 294 224 295
rect 222 294 223 295
rect 221 294 222 295
rect 220 294 221 295
rect 219 294 220 295
rect 218 294 219 295
rect 217 294 218 295
rect 216 294 217 295
rect 215 294 216 295
rect 214 294 215 295
rect 213 294 214 295
rect 212 294 213 295
rect 211 294 212 295
rect 210 294 211 295
rect 209 294 210 295
rect 184 294 185 295
rect 183 294 184 295
rect 182 294 183 295
rect 181 294 182 295
rect 180 294 181 295
rect 179 294 180 295
rect 178 294 179 295
rect 177 294 178 295
rect 176 294 177 295
rect 175 294 176 295
rect 174 294 175 295
rect 173 294 174 295
rect 172 294 173 295
rect 171 294 172 295
rect 170 294 171 295
rect 169 294 170 295
rect 168 294 169 295
rect 167 294 168 295
rect 166 294 167 295
rect 165 294 166 295
rect 164 294 165 295
rect 163 294 164 295
rect 162 294 163 295
rect 161 294 162 295
rect 160 294 161 295
rect 159 294 160 295
rect 158 294 159 295
rect 157 294 158 295
rect 156 294 157 295
rect 155 294 156 295
rect 154 294 155 295
rect 153 294 154 295
rect 152 294 153 295
rect 151 294 152 295
rect 150 294 151 295
rect 149 294 150 295
rect 148 294 149 295
rect 147 294 148 295
rect 146 294 147 295
rect 145 294 146 295
rect 144 294 145 295
rect 143 294 144 295
rect 142 294 143 295
rect 141 294 142 295
rect 140 294 141 295
rect 139 294 140 295
rect 138 294 139 295
rect 118 294 119 295
rect 117 294 118 295
rect 116 294 117 295
rect 115 294 116 295
rect 114 294 115 295
rect 113 294 114 295
rect 112 294 113 295
rect 111 294 112 295
rect 110 294 111 295
rect 109 294 110 295
rect 108 294 109 295
rect 107 294 108 295
rect 106 294 107 295
rect 105 294 106 295
rect 104 294 105 295
rect 103 294 104 295
rect 102 294 103 295
rect 101 294 102 295
rect 100 294 101 295
rect 99 294 100 295
rect 98 294 99 295
rect 97 294 98 295
rect 96 294 97 295
rect 95 294 96 295
rect 94 294 95 295
rect 93 294 94 295
rect 92 294 93 295
rect 91 294 92 295
rect 90 294 91 295
rect 89 294 90 295
rect 88 294 89 295
rect 87 294 88 295
rect 86 294 87 295
rect 85 294 86 295
rect 84 294 85 295
rect 83 294 84 295
rect 82 294 83 295
rect 66 294 67 295
rect 65 294 66 295
rect 64 294 65 295
rect 63 294 64 295
rect 62 294 63 295
rect 61 294 62 295
rect 60 294 61 295
rect 59 294 60 295
rect 58 294 59 295
rect 57 294 58 295
rect 56 294 57 295
rect 55 294 56 295
rect 54 294 55 295
rect 53 294 54 295
rect 52 294 53 295
rect 51 294 52 295
rect 50 294 51 295
rect 49 294 50 295
rect 48 294 49 295
rect 47 294 48 295
rect 46 294 47 295
rect 45 294 46 295
rect 44 294 45 295
rect 43 294 44 295
rect 42 294 43 295
rect 41 294 42 295
rect 40 294 41 295
rect 39 294 40 295
rect 38 294 39 295
rect 37 294 38 295
rect 27 294 28 295
rect 26 294 27 295
rect 25 294 26 295
rect 24 294 25 295
rect 23 294 24 295
rect 22 294 23 295
rect 21 294 22 295
rect 20 294 21 295
rect 19 294 20 295
rect 18 294 19 295
rect 17 294 18 295
rect 16 294 17 295
rect 15 294 16 295
rect 14 294 15 295
rect 13 294 14 295
rect 12 294 13 295
rect 11 294 12 295
rect 10 294 11 295
rect 9 294 10 295
rect 8 294 9 295
rect 7 294 8 295
rect 6 294 7 295
rect 5 294 6 295
rect 4 294 5 295
rect 3 294 4 295
rect 2 294 3 295
rect 478 295 479 296
rect 458 295 459 296
rect 415 295 416 296
rect 414 295 415 296
rect 413 295 414 296
rect 412 295 413 296
rect 270 295 271 296
rect 269 295 270 296
rect 268 295 269 296
rect 267 295 268 296
rect 266 295 267 296
rect 265 295 266 296
rect 264 295 265 296
rect 263 295 264 296
rect 262 295 263 296
rect 261 295 262 296
rect 260 295 261 296
rect 259 295 260 296
rect 258 295 259 296
rect 257 295 258 296
rect 256 295 257 296
rect 255 295 256 296
rect 254 295 255 296
rect 253 295 254 296
rect 252 295 253 296
rect 251 295 252 296
rect 250 295 251 296
rect 249 295 250 296
rect 248 295 249 296
rect 247 295 248 296
rect 246 295 247 296
rect 245 295 246 296
rect 244 295 245 296
rect 243 295 244 296
rect 242 295 243 296
rect 241 295 242 296
rect 240 295 241 296
rect 239 295 240 296
rect 238 295 239 296
rect 237 295 238 296
rect 236 295 237 296
rect 235 295 236 296
rect 234 295 235 296
rect 233 295 234 296
rect 232 295 233 296
rect 231 295 232 296
rect 230 295 231 296
rect 229 295 230 296
rect 228 295 229 296
rect 227 295 228 296
rect 226 295 227 296
rect 225 295 226 296
rect 224 295 225 296
rect 223 295 224 296
rect 222 295 223 296
rect 221 295 222 296
rect 220 295 221 296
rect 219 295 220 296
rect 218 295 219 296
rect 217 295 218 296
rect 216 295 217 296
rect 215 295 216 296
rect 214 295 215 296
rect 213 295 214 296
rect 212 295 213 296
rect 211 295 212 296
rect 210 295 211 296
rect 209 295 210 296
rect 208 295 209 296
rect 183 295 184 296
rect 182 295 183 296
rect 181 295 182 296
rect 180 295 181 296
rect 179 295 180 296
rect 178 295 179 296
rect 177 295 178 296
rect 176 295 177 296
rect 175 295 176 296
rect 174 295 175 296
rect 173 295 174 296
rect 172 295 173 296
rect 171 295 172 296
rect 170 295 171 296
rect 169 295 170 296
rect 168 295 169 296
rect 167 295 168 296
rect 166 295 167 296
rect 165 295 166 296
rect 164 295 165 296
rect 163 295 164 296
rect 162 295 163 296
rect 161 295 162 296
rect 160 295 161 296
rect 159 295 160 296
rect 158 295 159 296
rect 157 295 158 296
rect 156 295 157 296
rect 155 295 156 296
rect 154 295 155 296
rect 153 295 154 296
rect 152 295 153 296
rect 151 295 152 296
rect 150 295 151 296
rect 149 295 150 296
rect 148 295 149 296
rect 147 295 148 296
rect 146 295 147 296
rect 145 295 146 296
rect 144 295 145 296
rect 143 295 144 296
rect 142 295 143 296
rect 141 295 142 296
rect 140 295 141 296
rect 139 295 140 296
rect 118 295 119 296
rect 117 295 118 296
rect 116 295 117 296
rect 115 295 116 296
rect 114 295 115 296
rect 113 295 114 296
rect 112 295 113 296
rect 111 295 112 296
rect 110 295 111 296
rect 109 295 110 296
rect 108 295 109 296
rect 107 295 108 296
rect 106 295 107 296
rect 105 295 106 296
rect 104 295 105 296
rect 103 295 104 296
rect 102 295 103 296
rect 101 295 102 296
rect 100 295 101 296
rect 99 295 100 296
rect 98 295 99 296
rect 97 295 98 296
rect 96 295 97 296
rect 95 295 96 296
rect 94 295 95 296
rect 93 295 94 296
rect 92 295 93 296
rect 91 295 92 296
rect 90 295 91 296
rect 89 295 90 296
rect 88 295 89 296
rect 87 295 88 296
rect 86 295 87 296
rect 85 295 86 296
rect 84 295 85 296
rect 83 295 84 296
rect 82 295 83 296
rect 66 295 67 296
rect 65 295 66 296
rect 64 295 65 296
rect 63 295 64 296
rect 62 295 63 296
rect 61 295 62 296
rect 60 295 61 296
rect 59 295 60 296
rect 58 295 59 296
rect 57 295 58 296
rect 56 295 57 296
rect 55 295 56 296
rect 54 295 55 296
rect 53 295 54 296
rect 52 295 53 296
rect 51 295 52 296
rect 50 295 51 296
rect 49 295 50 296
rect 48 295 49 296
rect 47 295 48 296
rect 46 295 47 296
rect 45 295 46 296
rect 44 295 45 296
rect 43 295 44 296
rect 42 295 43 296
rect 41 295 42 296
rect 40 295 41 296
rect 39 295 40 296
rect 38 295 39 296
rect 28 295 29 296
rect 27 295 28 296
rect 26 295 27 296
rect 25 295 26 296
rect 24 295 25 296
rect 23 295 24 296
rect 22 295 23 296
rect 21 295 22 296
rect 20 295 21 296
rect 19 295 20 296
rect 18 295 19 296
rect 17 295 18 296
rect 16 295 17 296
rect 15 295 16 296
rect 14 295 15 296
rect 13 295 14 296
rect 12 295 13 296
rect 11 295 12 296
rect 10 295 11 296
rect 9 295 10 296
rect 8 295 9 296
rect 7 295 8 296
rect 6 295 7 296
rect 5 295 6 296
rect 4 295 5 296
rect 3 295 4 296
rect 2 295 3 296
rect 478 296 479 297
rect 458 296 459 297
rect 415 296 416 297
rect 414 296 415 297
rect 413 296 414 297
rect 412 296 413 297
rect 269 296 270 297
rect 268 296 269 297
rect 267 296 268 297
rect 266 296 267 297
rect 265 296 266 297
rect 264 296 265 297
rect 263 296 264 297
rect 262 296 263 297
rect 261 296 262 297
rect 260 296 261 297
rect 259 296 260 297
rect 258 296 259 297
rect 257 296 258 297
rect 256 296 257 297
rect 255 296 256 297
rect 254 296 255 297
rect 253 296 254 297
rect 252 296 253 297
rect 251 296 252 297
rect 250 296 251 297
rect 249 296 250 297
rect 248 296 249 297
rect 247 296 248 297
rect 246 296 247 297
rect 245 296 246 297
rect 244 296 245 297
rect 243 296 244 297
rect 242 296 243 297
rect 241 296 242 297
rect 240 296 241 297
rect 239 296 240 297
rect 238 296 239 297
rect 237 296 238 297
rect 236 296 237 297
rect 235 296 236 297
rect 234 296 235 297
rect 233 296 234 297
rect 232 296 233 297
rect 231 296 232 297
rect 230 296 231 297
rect 229 296 230 297
rect 228 296 229 297
rect 227 296 228 297
rect 226 296 227 297
rect 225 296 226 297
rect 224 296 225 297
rect 223 296 224 297
rect 222 296 223 297
rect 221 296 222 297
rect 220 296 221 297
rect 219 296 220 297
rect 218 296 219 297
rect 217 296 218 297
rect 216 296 217 297
rect 215 296 216 297
rect 214 296 215 297
rect 213 296 214 297
rect 212 296 213 297
rect 211 296 212 297
rect 210 296 211 297
rect 209 296 210 297
rect 208 296 209 297
rect 207 296 208 297
rect 182 296 183 297
rect 181 296 182 297
rect 180 296 181 297
rect 179 296 180 297
rect 178 296 179 297
rect 177 296 178 297
rect 176 296 177 297
rect 175 296 176 297
rect 174 296 175 297
rect 173 296 174 297
rect 172 296 173 297
rect 171 296 172 297
rect 170 296 171 297
rect 169 296 170 297
rect 168 296 169 297
rect 167 296 168 297
rect 166 296 167 297
rect 165 296 166 297
rect 164 296 165 297
rect 163 296 164 297
rect 162 296 163 297
rect 161 296 162 297
rect 160 296 161 297
rect 159 296 160 297
rect 158 296 159 297
rect 157 296 158 297
rect 156 296 157 297
rect 155 296 156 297
rect 154 296 155 297
rect 153 296 154 297
rect 152 296 153 297
rect 151 296 152 297
rect 150 296 151 297
rect 149 296 150 297
rect 148 296 149 297
rect 147 296 148 297
rect 146 296 147 297
rect 145 296 146 297
rect 144 296 145 297
rect 143 296 144 297
rect 142 296 143 297
rect 141 296 142 297
rect 140 296 141 297
rect 119 296 120 297
rect 118 296 119 297
rect 117 296 118 297
rect 116 296 117 297
rect 115 296 116 297
rect 114 296 115 297
rect 113 296 114 297
rect 112 296 113 297
rect 111 296 112 297
rect 110 296 111 297
rect 109 296 110 297
rect 108 296 109 297
rect 107 296 108 297
rect 106 296 107 297
rect 105 296 106 297
rect 104 296 105 297
rect 103 296 104 297
rect 102 296 103 297
rect 101 296 102 297
rect 100 296 101 297
rect 99 296 100 297
rect 98 296 99 297
rect 97 296 98 297
rect 96 296 97 297
rect 95 296 96 297
rect 94 296 95 297
rect 93 296 94 297
rect 92 296 93 297
rect 91 296 92 297
rect 90 296 91 297
rect 89 296 90 297
rect 88 296 89 297
rect 87 296 88 297
rect 86 296 87 297
rect 85 296 86 297
rect 84 296 85 297
rect 83 296 84 297
rect 66 296 67 297
rect 65 296 66 297
rect 64 296 65 297
rect 63 296 64 297
rect 62 296 63 297
rect 61 296 62 297
rect 60 296 61 297
rect 59 296 60 297
rect 58 296 59 297
rect 57 296 58 297
rect 56 296 57 297
rect 55 296 56 297
rect 54 296 55 297
rect 53 296 54 297
rect 52 296 53 297
rect 51 296 52 297
rect 50 296 51 297
rect 49 296 50 297
rect 48 296 49 297
rect 47 296 48 297
rect 46 296 47 297
rect 45 296 46 297
rect 44 296 45 297
rect 43 296 44 297
rect 42 296 43 297
rect 41 296 42 297
rect 40 296 41 297
rect 39 296 40 297
rect 38 296 39 297
rect 28 296 29 297
rect 27 296 28 297
rect 26 296 27 297
rect 25 296 26 297
rect 24 296 25 297
rect 23 296 24 297
rect 22 296 23 297
rect 21 296 22 297
rect 20 296 21 297
rect 19 296 20 297
rect 18 296 19 297
rect 17 296 18 297
rect 16 296 17 297
rect 15 296 16 297
rect 14 296 15 297
rect 13 296 14 297
rect 12 296 13 297
rect 11 296 12 297
rect 10 296 11 297
rect 9 296 10 297
rect 8 296 9 297
rect 7 296 8 297
rect 6 296 7 297
rect 5 296 6 297
rect 4 296 5 297
rect 3 296 4 297
rect 2 296 3 297
rect 478 297 479 298
rect 458 297 459 298
rect 415 297 416 298
rect 414 297 415 298
rect 413 297 414 298
rect 412 297 413 298
rect 268 297 269 298
rect 267 297 268 298
rect 266 297 267 298
rect 265 297 266 298
rect 264 297 265 298
rect 263 297 264 298
rect 262 297 263 298
rect 261 297 262 298
rect 260 297 261 298
rect 259 297 260 298
rect 258 297 259 298
rect 257 297 258 298
rect 256 297 257 298
rect 255 297 256 298
rect 254 297 255 298
rect 253 297 254 298
rect 252 297 253 298
rect 251 297 252 298
rect 250 297 251 298
rect 249 297 250 298
rect 248 297 249 298
rect 247 297 248 298
rect 246 297 247 298
rect 245 297 246 298
rect 244 297 245 298
rect 243 297 244 298
rect 242 297 243 298
rect 241 297 242 298
rect 240 297 241 298
rect 239 297 240 298
rect 238 297 239 298
rect 237 297 238 298
rect 236 297 237 298
rect 235 297 236 298
rect 234 297 235 298
rect 233 297 234 298
rect 232 297 233 298
rect 231 297 232 298
rect 230 297 231 298
rect 229 297 230 298
rect 228 297 229 298
rect 227 297 228 298
rect 226 297 227 298
rect 225 297 226 298
rect 224 297 225 298
rect 223 297 224 298
rect 222 297 223 298
rect 221 297 222 298
rect 220 297 221 298
rect 219 297 220 298
rect 218 297 219 298
rect 217 297 218 298
rect 216 297 217 298
rect 215 297 216 298
rect 214 297 215 298
rect 213 297 214 298
rect 212 297 213 298
rect 211 297 212 298
rect 210 297 211 298
rect 209 297 210 298
rect 208 297 209 298
rect 207 297 208 298
rect 180 297 181 298
rect 179 297 180 298
rect 178 297 179 298
rect 177 297 178 298
rect 176 297 177 298
rect 175 297 176 298
rect 174 297 175 298
rect 173 297 174 298
rect 172 297 173 298
rect 171 297 172 298
rect 170 297 171 298
rect 169 297 170 298
rect 168 297 169 298
rect 167 297 168 298
rect 166 297 167 298
rect 165 297 166 298
rect 164 297 165 298
rect 163 297 164 298
rect 162 297 163 298
rect 161 297 162 298
rect 160 297 161 298
rect 159 297 160 298
rect 158 297 159 298
rect 157 297 158 298
rect 156 297 157 298
rect 155 297 156 298
rect 154 297 155 298
rect 153 297 154 298
rect 152 297 153 298
rect 151 297 152 298
rect 150 297 151 298
rect 149 297 150 298
rect 148 297 149 298
rect 147 297 148 298
rect 146 297 147 298
rect 145 297 146 298
rect 144 297 145 298
rect 143 297 144 298
rect 142 297 143 298
rect 141 297 142 298
rect 119 297 120 298
rect 118 297 119 298
rect 117 297 118 298
rect 116 297 117 298
rect 115 297 116 298
rect 114 297 115 298
rect 113 297 114 298
rect 112 297 113 298
rect 111 297 112 298
rect 110 297 111 298
rect 109 297 110 298
rect 108 297 109 298
rect 107 297 108 298
rect 106 297 107 298
rect 105 297 106 298
rect 104 297 105 298
rect 103 297 104 298
rect 102 297 103 298
rect 101 297 102 298
rect 100 297 101 298
rect 99 297 100 298
rect 98 297 99 298
rect 97 297 98 298
rect 96 297 97 298
rect 95 297 96 298
rect 94 297 95 298
rect 93 297 94 298
rect 92 297 93 298
rect 91 297 92 298
rect 90 297 91 298
rect 89 297 90 298
rect 88 297 89 298
rect 87 297 88 298
rect 86 297 87 298
rect 85 297 86 298
rect 84 297 85 298
rect 83 297 84 298
rect 67 297 68 298
rect 66 297 67 298
rect 65 297 66 298
rect 64 297 65 298
rect 63 297 64 298
rect 62 297 63 298
rect 61 297 62 298
rect 60 297 61 298
rect 59 297 60 298
rect 58 297 59 298
rect 57 297 58 298
rect 56 297 57 298
rect 55 297 56 298
rect 54 297 55 298
rect 53 297 54 298
rect 52 297 53 298
rect 51 297 52 298
rect 50 297 51 298
rect 49 297 50 298
rect 48 297 49 298
rect 47 297 48 298
rect 46 297 47 298
rect 45 297 46 298
rect 44 297 45 298
rect 43 297 44 298
rect 42 297 43 298
rect 41 297 42 298
rect 40 297 41 298
rect 39 297 40 298
rect 38 297 39 298
rect 28 297 29 298
rect 27 297 28 298
rect 26 297 27 298
rect 25 297 26 298
rect 24 297 25 298
rect 23 297 24 298
rect 22 297 23 298
rect 21 297 22 298
rect 20 297 21 298
rect 19 297 20 298
rect 18 297 19 298
rect 17 297 18 298
rect 16 297 17 298
rect 15 297 16 298
rect 14 297 15 298
rect 13 297 14 298
rect 12 297 13 298
rect 11 297 12 298
rect 10 297 11 298
rect 9 297 10 298
rect 8 297 9 298
rect 7 297 8 298
rect 6 297 7 298
rect 5 297 6 298
rect 4 297 5 298
rect 3 297 4 298
rect 459 298 460 299
rect 458 298 459 299
rect 415 298 416 299
rect 414 298 415 299
rect 413 298 414 299
rect 412 298 413 299
rect 267 298 268 299
rect 266 298 267 299
rect 265 298 266 299
rect 264 298 265 299
rect 263 298 264 299
rect 262 298 263 299
rect 261 298 262 299
rect 260 298 261 299
rect 259 298 260 299
rect 258 298 259 299
rect 257 298 258 299
rect 256 298 257 299
rect 255 298 256 299
rect 254 298 255 299
rect 253 298 254 299
rect 252 298 253 299
rect 251 298 252 299
rect 250 298 251 299
rect 249 298 250 299
rect 248 298 249 299
rect 247 298 248 299
rect 246 298 247 299
rect 245 298 246 299
rect 244 298 245 299
rect 243 298 244 299
rect 242 298 243 299
rect 241 298 242 299
rect 240 298 241 299
rect 239 298 240 299
rect 238 298 239 299
rect 237 298 238 299
rect 236 298 237 299
rect 235 298 236 299
rect 234 298 235 299
rect 233 298 234 299
rect 232 298 233 299
rect 231 298 232 299
rect 230 298 231 299
rect 229 298 230 299
rect 228 298 229 299
rect 227 298 228 299
rect 226 298 227 299
rect 225 298 226 299
rect 224 298 225 299
rect 223 298 224 299
rect 222 298 223 299
rect 221 298 222 299
rect 220 298 221 299
rect 219 298 220 299
rect 218 298 219 299
rect 217 298 218 299
rect 216 298 217 299
rect 215 298 216 299
rect 214 298 215 299
rect 213 298 214 299
rect 212 298 213 299
rect 211 298 212 299
rect 210 298 211 299
rect 209 298 210 299
rect 208 298 209 299
rect 207 298 208 299
rect 206 298 207 299
rect 179 298 180 299
rect 178 298 179 299
rect 177 298 178 299
rect 176 298 177 299
rect 175 298 176 299
rect 174 298 175 299
rect 173 298 174 299
rect 172 298 173 299
rect 171 298 172 299
rect 170 298 171 299
rect 169 298 170 299
rect 168 298 169 299
rect 167 298 168 299
rect 166 298 167 299
rect 165 298 166 299
rect 164 298 165 299
rect 163 298 164 299
rect 162 298 163 299
rect 161 298 162 299
rect 160 298 161 299
rect 159 298 160 299
rect 158 298 159 299
rect 157 298 158 299
rect 156 298 157 299
rect 155 298 156 299
rect 154 298 155 299
rect 153 298 154 299
rect 152 298 153 299
rect 151 298 152 299
rect 150 298 151 299
rect 149 298 150 299
rect 148 298 149 299
rect 147 298 148 299
rect 146 298 147 299
rect 145 298 146 299
rect 144 298 145 299
rect 143 298 144 299
rect 142 298 143 299
rect 119 298 120 299
rect 118 298 119 299
rect 117 298 118 299
rect 116 298 117 299
rect 115 298 116 299
rect 114 298 115 299
rect 113 298 114 299
rect 112 298 113 299
rect 111 298 112 299
rect 110 298 111 299
rect 109 298 110 299
rect 108 298 109 299
rect 107 298 108 299
rect 106 298 107 299
rect 105 298 106 299
rect 104 298 105 299
rect 103 298 104 299
rect 102 298 103 299
rect 101 298 102 299
rect 100 298 101 299
rect 99 298 100 299
rect 98 298 99 299
rect 97 298 98 299
rect 96 298 97 299
rect 95 298 96 299
rect 94 298 95 299
rect 93 298 94 299
rect 92 298 93 299
rect 91 298 92 299
rect 90 298 91 299
rect 89 298 90 299
rect 88 298 89 299
rect 87 298 88 299
rect 86 298 87 299
rect 85 298 86 299
rect 84 298 85 299
rect 83 298 84 299
rect 67 298 68 299
rect 66 298 67 299
rect 65 298 66 299
rect 64 298 65 299
rect 63 298 64 299
rect 62 298 63 299
rect 61 298 62 299
rect 60 298 61 299
rect 59 298 60 299
rect 58 298 59 299
rect 57 298 58 299
rect 56 298 57 299
rect 55 298 56 299
rect 54 298 55 299
rect 53 298 54 299
rect 52 298 53 299
rect 51 298 52 299
rect 50 298 51 299
rect 49 298 50 299
rect 48 298 49 299
rect 47 298 48 299
rect 46 298 47 299
rect 45 298 46 299
rect 44 298 45 299
rect 43 298 44 299
rect 42 298 43 299
rect 41 298 42 299
rect 40 298 41 299
rect 39 298 40 299
rect 38 298 39 299
rect 28 298 29 299
rect 27 298 28 299
rect 26 298 27 299
rect 25 298 26 299
rect 24 298 25 299
rect 23 298 24 299
rect 22 298 23 299
rect 21 298 22 299
rect 20 298 21 299
rect 19 298 20 299
rect 18 298 19 299
rect 17 298 18 299
rect 16 298 17 299
rect 15 298 16 299
rect 14 298 15 299
rect 13 298 14 299
rect 12 298 13 299
rect 11 298 12 299
rect 10 298 11 299
rect 9 298 10 299
rect 8 298 9 299
rect 7 298 8 299
rect 6 298 7 299
rect 5 298 6 299
rect 4 298 5 299
rect 3 298 4 299
rect 460 299 461 300
rect 459 299 460 300
rect 458 299 459 300
rect 415 299 416 300
rect 414 299 415 300
rect 413 299 414 300
rect 412 299 413 300
rect 266 299 267 300
rect 265 299 266 300
rect 264 299 265 300
rect 263 299 264 300
rect 262 299 263 300
rect 261 299 262 300
rect 260 299 261 300
rect 259 299 260 300
rect 258 299 259 300
rect 257 299 258 300
rect 256 299 257 300
rect 255 299 256 300
rect 254 299 255 300
rect 253 299 254 300
rect 252 299 253 300
rect 251 299 252 300
rect 250 299 251 300
rect 249 299 250 300
rect 248 299 249 300
rect 247 299 248 300
rect 246 299 247 300
rect 245 299 246 300
rect 244 299 245 300
rect 243 299 244 300
rect 242 299 243 300
rect 241 299 242 300
rect 240 299 241 300
rect 239 299 240 300
rect 238 299 239 300
rect 237 299 238 300
rect 236 299 237 300
rect 235 299 236 300
rect 234 299 235 300
rect 233 299 234 300
rect 232 299 233 300
rect 231 299 232 300
rect 230 299 231 300
rect 229 299 230 300
rect 228 299 229 300
rect 227 299 228 300
rect 226 299 227 300
rect 225 299 226 300
rect 224 299 225 300
rect 223 299 224 300
rect 222 299 223 300
rect 221 299 222 300
rect 220 299 221 300
rect 219 299 220 300
rect 218 299 219 300
rect 217 299 218 300
rect 216 299 217 300
rect 215 299 216 300
rect 214 299 215 300
rect 213 299 214 300
rect 212 299 213 300
rect 211 299 212 300
rect 210 299 211 300
rect 209 299 210 300
rect 208 299 209 300
rect 207 299 208 300
rect 206 299 207 300
rect 205 299 206 300
rect 178 299 179 300
rect 177 299 178 300
rect 176 299 177 300
rect 175 299 176 300
rect 174 299 175 300
rect 173 299 174 300
rect 172 299 173 300
rect 171 299 172 300
rect 170 299 171 300
rect 169 299 170 300
rect 168 299 169 300
rect 167 299 168 300
rect 166 299 167 300
rect 165 299 166 300
rect 164 299 165 300
rect 163 299 164 300
rect 162 299 163 300
rect 161 299 162 300
rect 160 299 161 300
rect 159 299 160 300
rect 158 299 159 300
rect 157 299 158 300
rect 156 299 157 300
rect 155 299 156 300
rect 154 299 155 300
rect 153 299 154 300
rect 152 299 153 300
rect 151 299 152 300
rect 150 299 151 300
rect 149 299 150 300
rect 148 299 149 300
rect 147 299 148 300
rect 146 299 147 300
rect 145 299 146 300
rect 144 299 145 300
rect 120 299 121 300
rect 119 299 120 300
rect 118 299 119 300
rect 117 299 118 300
rect 116 299 117 300
rect 115 299 116 300
rect 114 299 115 300
rect 113 299 114 300
rect 112 299 113 300
rect 111 299 112 300
rect 110 299 111 300
rect 109 299 110 300
rect 108 299 109 300
rect 107 299 108 300
rect 106 299 107 300
rect 105 299 106 300
rect 104 299 105 300
rect 103 299 104 300
rect 102 299 103 300
rect 101 299 102 300
rect 100 299 101 300
rect 99 299 100 300
rect 98 299 99 300
rect 97 299 98 300
rect 96 299 97 300
rect 95 299 96 300
rect 94 299 95 300
rect 93 299 94 300
rect 92 299 93 300
rect 91 299 92 300
rect 90 299 91 300
rect 89 299 90 300
rect 88 299 89 300
rect 87 299 88 300
rect 86 299 87 300
rect 85 299 86 300
rect 84 299 85 300
rect 83 299 84 300
rect 67 299 68 300
rect 66 299 67 300
rect 65 299 66 300
rect 64 299 65 300
rect 63 299 64 300
rect 62 299 63 300
rect 61 299 62 300
rect 60 299 61 300
rect 59 299 60 300
rect 58 299 59 300
rect 57 299 58 300
rect 56 299 57 300
rect 55 299 56 300
rect 54 299 55 300
rect 53 299 54 300
rect 52 299 53 300
rect 51 299 52 300
rect 50 299 51 300
rect 49 299 50 300
rect 48 299 49 300
rect 47 299 48 300
rect 46 299 47 300
rect 45 299 46 300
rect 44 299 45 300
rect 43 299 44 300
rect 42 299 43 300
rect 41 299 42 300
rect 40 299 41 300
rect 39 299 40 300
rect 28 299 29 300
rect 27 299 28 300
rect 26 299 27 300
rect 25 299 26 300
rect 24 299 25 300
rect 23 299 24 300
rect 22 299 23 300
rect 21 299 22 300
rect 20 299 21 300
rect 19 299 20 300
rect 18 299 19 300
rect 17 299 18 300
rect 16 299 17 300
rect 15 299 16 300
rect 14 299 15 300
rect 13 299 14 300
rect 12 299 13 300
rect 11 299 12 300
rect 10 299 11 300
rect 9 299 10 300
rect 8 299 9 300
rect 7 299 8 300
rect 6 299 7 300
rect 5 299 6 300
rect 4 299 5 300
rect 3 299 4 300
rect 462 300 463 301
rect 461 300 462 301
rect 460 300 461 301
rect 459 300 460 301
rect 458 300 459 301
rect 457 300 458 301
rect 437 300 438 301
rect 436 300 437 301
rect 415 300 416 301
rect 414 300 415 301
rect 413 300 414 301
rect 412 300 413 301
rect 394 300 395 301
rect 393 300 394 301
rect 264 300 265 301
rect 263 300 264 301
rect 262 300 263 301
rect 261 300 262 301
rect 260 300 261 301
rect 259 300 260 301
rect 258 300 259 301
rect 257 300 258 301
rect 256 300 257 301
rect 255 300 256 301
rect 254 300 255 301
rect 253 300 254 301
rect 252 300 253 301
rect 251 300 252 301
rect 250 300 251 301
rect 249 300 250 301
rect 248 300 249 301
rect 247 300 248 301
rect 246 300 247 301
rect 245 300 246 301
rect 244 300 245 301
rect 243 300 244 301
rect 242 300 243 301
rect 241 300 242 301
rect 240 300 241 301
rect 239 300 240 301
rect 238 300 239 301
rect 237 300 238 301
rect 236 300 237 301
rect 235 300 236 301
rect 234 300 235 301
rect 233 300 234 301
rect 232 300 233 301
rect 231 300 232 301
rect 230 300 231 301
rect 229 300 230 301
rect 228 300 229 301
rect 227 300 228 301
rect 226 300 227 301
rect 225 300 226 301
rect 224 300 225 301
rect 223 300 224 301
rect 222 300 223 301
rect 221 300 222 301
rect 220 300 221 301
rect 219 300 220 301
rect 218 300 219 301
rect 217 300 218 301
rect 216 300 217 301
rect 215 300 216 301
rect 214 300 215 301
rect 213 300 214 301
rect 212 300 213 301
rect 211 300 212 301
rect 210 300 211 301
rect 209 300 210 301
rect 208 300 209 301
rect 207 300 208 301
rect 206 300 207 301
rect 205 300 206 301
rect 176 300 177 301
rect 175 300 176 301
rect 174 300 175 301
rect 173 300 174 301
rect 172 300 173 301
rect 171 300 172 301
rect 170 300 171 301
rect 169 300 170 301
rect 168 300 169 301
rect 167 300 168 301
rect 166 300 167 301
rect 165 300 166 301
rect 164 300 165 301
rect 163 300 164 301
rect 162 300 163 301
rect 161 300 162 301
rect 160 300 161 301
rect 159 300 160 301
rect 158 300 159 301
rect 157 300 158 301
rect 156 300 157 301
rect 155 300 156 301
rect 154 300 155 301
rect 153 300 154 301
rect 152 300 153 301
rect 151 300 152 301
rect 150 300 151 301
rect 149 300 150 301
rect 148 300 149 301
rect 147 300 148 301
rect 146 300 147 301
rect 145 300 146 301
rect 120 300 121 301
rect 119 300 120 301
rect 118 300 119 301
rect 117 300 118 301
rect 116 300 117 301
rect 115 300 116 301
rect 114 300 115 301
rect 113 300 114 301
rect 112 300 113 301
rect 111 300 112 301
rect 110 300 111 301
rect 109 300 110 301
rect 108 300 109 301
rect 107 300 108 301
rect 106 300 107 301
rect 105 300 106 301
rect 104 300 105 301
rect 103 300 104 301
rect 102 300 103 301
rect 101 300 102 301
rect 100 300 101 301
rect 99 300 100 301
rect 98 300 99 301
rect 97 300 98 301
rect 96 300 97 301
rect 95 300 96 301
rect 94 300 95 301
rect 93 300 94 301
rect 92 300 93 301
rect 91 300 92 301
rect 90 300 91 301
rect 89 300 90 301
rect 88 300 89 301
rect 87 300 88 301
rect 86 300 87 301
rect 85 300 86 301
rect 84 300 85 301
rect 67 300 68 301
rect 66 300 67 301
rect 65 300 66 301
rect 64 300 65 301
rect 63 300 64 301
rect 62 300 63 301
rect 61 300 62 301
rect 60 300 61 301
rect 59 300 60 301
rect 58 300 59 301
rect 57 300 58 301
rect 56 300 57 301
rect 55 300 56 301
rect 54 300 55 301
rect 53 300 54 301
rect 52 300 53 301
rect 51 300 52 301
rect 50 300 51 301
rect 49 300 50 301
rect 48 300 49 301
rect 47 300 48 301
rect 46 300 47 301
rect 45 300 46 301
rect 44 300 45 301
rect 43 300 44 301
rect 42 300 43 301
rect 41 300 42 301
rect 40 300 41 301
rect 39 300 40 301
rect 28 300 29 301
rect 27 300 28 301
rect 26 300 27 301
rect 25 300 26 301
rect 24 300 25 301
rect 23 300 24 301
rect 22 300 23 301
rect 21 300 22 301
rect 20 300 21 301
rect 19 300 20 301
rect 18 300 19 301
rect 17 300 18 301
rect 16 300 17 301
rect 15 300 16 301
rect 14 300 15 301
rect 13 300 14 301
rect 12 300 13 301
rect 11 300 12 301
rect 10 300 11 301
rect 9 300 10 301
rect 8 300 9 301
rect 7 300 8 301
rect 6 300 7 301
rect 5 300 6 301
rect 4 300 5 301
rect 462 301 463 302
rect 461 301 462 302
rect 460 301 461 302
rect 459 301 460 302
rect 458 301 459 302
rect 457 301 458 302
rect 437 301 438 302
rect 436 301 437 302
rect 435 301 436 302
rect 415 301 416 302
rect 414 301 415 302
rect 413 301 414 302
rect 412 301 413 302
rect 395 301 396 302
rect 394 301 395 302
rect 393 301 394 302
rect 263 301 264 302
rect 262 301 263 302
rect 261 301 262 302
rect 260 301 261 302
rect 259 301 260 302
rect 258 301 259 302
rect 257 301 258 302
rect 256 301 257 302
rect 255 301 256 302
rect 254 301 255 302
rect 253 301 254 302
rect 252 301 253 302
rect 251 301 252 302
rect 250 301 251 302
rect 249 301 250 302
rect 248 301 249 302
rect 247 301 248 302
rect 246 301 247 302
rect 245 301 246 302
rect 244 301 245 302
rect 243 301 244 302
rect 242 301 243 302
rect 241 301 242 302
rect 240 301 241 302
rect 239 301 240 302
rect 238 301 239 302
rect 237 301 238 302
rect 236 301 237 302
rect 235 301 236 302
rect 234 301 235 302
rect 233 301 234 302
rect 232 301 233 302
rect 231 301 232 302
rect 230 301 231 302
rect 229 301 230 302
rect 228 301 229 302
rect 227 301 228 302
rect 226 301 227 302
rect 225 301 226 302
rect 224 301 225 302
rect 223 301 224 302
rect 222 301 223 302
rect 221 301 222 302
rect 220 301 221 302
rect 219 301 220 302
rect 218 301 219 302
rect 217 301 218 302
rect 216 301 217 302
rect 215 301 216 302
rect 214 301 215 302
rect 213 301 214 302
rect 212 301 213 302
rect 211 301 212 302
rect 210 301 211 302
rect 209 301 210 302
rect 208 301 209 302
rect 207 301 208 302
rect 206 301 207 302
rect 205 301 206 302
rect 204 301 205 302
rect 175 301 176 302
rect 174 301 175 302
rect 173 301 174 302
rect 172 301 173 302
rect 171 301 172 302
rect 170 301 171 302
rect 169 301 170 302
rect 168 301 169 302
rect 167 301 168 302
rect 166 301 167 302
rect 165 301 166 302
rect 164 301 165 302
rect 163 301 164 302
rect 162 301 163 302
rect 161 301 162 302
rect 160 301 161 302
rect 159 301 160 302
rect 158 301 159 302
rect 157 301 158 302
rect 156 301 157 302
rect 155 301 156 302
rect 154 301 155 302
rect 153 301 154 302
rect 152 301 153 302
rect 151 301 152 302
rect 150 301 151 302
rect 149 301 150 302
rect 148 301 149 302
rect 147 301 148 302
rect 121 301 122 302
rect 120 301 121 302
rect 119 301 120 302
rect 118 301 119 302
rect 117 301 118 302
rect 116 301 117 302
rect 115 301 116 302
rect 114 301 115 302
rect 113 301 114 302
rect 112 301 113 302
rect 111 301 112 302
rect 110 301 111 302
rect 109 301 110 302
rect 108 301 109 302
rect 107 301 108 302
rect 106 301 107 302
rect 105 301 106 302
rect 104 301 105 302
rect 103 301 104 302
rect 102 301 103 302
rect 101 301 102 302
rect 100 301 101 302
rect 99 301 100 302
rect 98 301 99 302
rect 97 301 98 302
rect 96 301 97 302
rect 95 301 96 302
rect 94 301 95 302
rect 93 301 94 302
rect 92 301 93 302
rect 91 301 92 302
rect 90 301 91 302
rect 89 301 90 302
rect 88 301 89 302
rect 87 301 88 302
rect 86 301 87 302
rect 85 301 86 302
rect 84 301 85 302
rect 68 301 69 302
rect 67 301 68 302
rect 66 301 67 302
rect 65 301 66 302
rect 64 301 65 302
rect 63 301 64 302
rect 62 301 63 302
rect 61 301 62 302
rect 60 301 61 302
rect 59 301 60 302
rect 58 301 59 302
rect 57 301 58 302
rect 56 301 57 302
rect 55 301 56 302
rect 54 301 55 302
rect 53 301 54 302
rect 52 301 53 302
rect 51 301 52 302
rect 50 301 51 302
rect 49 301 50 302
rect 48 301 49 302
rect 47 301 48 302
rect 46 301 47 302
rect 45 301 46 302
rect 44 301 45 302
rect 43 301 44 302
rect 42 301 43 302
rect 41 301 42 302
rect 40 301 41 302
rect 39 301 40 302
rect 29 301 30 302
rect 28 301 29 302
rect 27 301 28 302
rect 26 301 27 302
rect 25 301 26 302
rect 24 301 25 302
rect 23 301 24 302
rect 22 301 23 302
rect 21 301 22 302
rect 20 301 21 302
rect 19 301 20 302
rect 18 301 19 302
rect 17 301 18 302
rect 16 301 17 302
rect 15 301 16 302
rect 14 301 15 302
rect 13 301 14 302
rect 12 301 13 302
rect 11 301 12 302
rect 10 301 11 302
rect 9 301 10 302
rect 8 301 9 302
rect 7 301 8 302
rect 6 301 7 302
rect 5 301 6 302
rect 4 301 5 302
rect 437 302 438 303
rect 436 302 437 303
rect 435 302 436 303
rect 415 302 416 303
rect 414 302 415 303
rect 413 302 414 303
rect 412 302 413 303
rect 395 302 396 303
rect 394 302 395 303
rect 393 302 394 303
rect 262 302 263 303
rect 261 302 262 303
rect 260 302 261 303
rect 259 302 260 303
rect 258 302 259 303
rect 257 302 258 303
rect 256 302 257 303
rect 255 302 256 303
rect 254 302 255 303
rect 253 302 254 303
rect 252 302 253 303
rect 251 302 252 303
rect 250 302 251 303
rect 249 302 250 303
rect 248 302 249 303
rect 247 302 248 303
rect 246 302 247 303
rect 245 302 246 303
rect 244 302 245 303
rect 243 302 244 303
rect 242 302 243 303
rect 241 302 242 303
rect 240 302 241 303
rect 239 302 240 303
rect 238 302 239 303
rect 237 302 238 303
rect 236 302 237 303
rect 235 302 236 303
rect 234 302 235 303
rect 233 302 234 303
rect 232 302 233 303
rect 231 302 232 303
rect 230 302 231 303
rect 229 302 230 303
rect 228 302 229 303
rect 227 302 228 303
rect 226 302 227 303
rect 225 302 226 303
rect 224 302 225 303
rect 223 302 224 303
rect 222 302 223 303
rect 221 302 222 303
rect 220 302 221 303
rect 219 302 220 303
rect 218 302 219 303
rect 217 302 218 303
rect 216 302 217 303
rect 215 302 216 303
rect 214 302 215 303
rect 213 302 214 303
rect 212 302 213 303
rect 211 302 212 303
rect 210 302 211 303
rect 209 302 210 303
rect 208 302 209 303
rect 207 302 208 303
rect 206 302 207 303
rect 205 302 206 303
rect 204 302 205 303
rect 203 302 204 303
rect 173 302 174 303
rect 172 302 173 303
rect 171 302 172 303
rect 170 302 171 303
rect 169 302 170 303
rect 168 302 169 303
rect 167 302 168 303
rect 166 302 167 303
rect 165 302 166 303
rect 164 302 165 303
rect 163 302 164 303
rect 162 302 163 303
rect 161 302 162 303
rect 160 302 161 303
rect 159 302 160 303
rect 158 302 159 303
rect 157 302 158 303
rect 156 302 157 303
rect 155 302 156 303
rect 154 302 155 303
rect 153 302 154 303
rect 152 302 153 303
rect 151 302 152 303
rect 150 302 151 303
rect 149 302 150 303
rect 121 302 122 303
rect 120 302 121 303
rect 119 302 120 303
rect 118 302 119 303
rect 117 302 118 303
rect 116 302 117 303
rect 115 302 116 303
rect 114 302 115 303
rect 113 302 114 303
rect 112 302 113 303
rect 111 302 112 303
rect 110 302 111 303
rect 109 302 110 303
rect 108 302 109 303
rect 107 302 108 303
rect 106 302 107 303
rect 105 302 106 303
rect 104 302 105 303
rect 103 302 104 303
rect 102 302 103 303
rect 101 302 102 303
rect 100 302 101 303
rect 99 302 100 303
rect 98 302 99 303
rect 97 302 98 303
rect 96 302 97 303
rect 95 302 96 303
rect 94 302 95 303
rect 93 302 94 303
rect 92 302 93 303
rect 91 302 92 303
rect 90 302 91 303
rect 89 302 90 303
rect 88 302 89 303
rect 87 302 88 303
rect 86 302 87 303
rect 85 302 86 303
rect 84 302 85 303
rect 68 302 69 303
rect 67 302 68 303
rect 66 302 67 303
rect 65 302 66 303
rect 64 302 65 303
rect 63 302 64 303
rect 62 302 63 303
rect 61 302 62 303
rect 60 302 61 303
rect 59 302 60 303
rect 58 302 59 303
rect 57 302 58 303
rect 56 302 57 303
rect 55 302 56 303
rect 54 302 55 303
rect 53 302 54 303
rect 52 302 53 303
rect 51 302 52 303
rect 50 302 51 303
rect 49 302 50 303
rect 48 302 49 303
rect 47 302 48 303
rect 46 302 47 303
rect 45 302 46 303
rect 44 302 45 303
rect 43 302 44 303
rect 42 302 43 303
rect 41 302 42 303
rect 40 302 41 303
rect 29 302 30 303
rect 28 302 29 303
rect 27 302 28 303
rect 26 302 27 303
rect 25 302 26 303
rect 24 302 25 303
rect 23 302 24 303
rect 22 302 23 303
rect 21 302 22 303
rect 20 302 21 303
rect 19 302 20 303
rect 18 302 19 303
rect 17 302 18 303
rect 16 302 17 303
rect 15 302 16 303
rect 14 302 15 303
rect 13 302 14 303
rect 12 302 13 303
rect 11 302 12 303
rect 10 302 11 303
rect 9 302 10 303
rect 8 302 9 303
rect 7 302 8 303
rect 6 302 7 303
rect 5 302 6 303
rect 437 303 438 304
rect 436 303 437 304
rect 435 303 436 304
rect 415 303 416 304
rect 414 303 415 304
rect 413 303 414 304
rect 412 303 413 304
rect 395 303 396 304
rect 394 303 395 304
rect 393 303 394 304
rect 260 303 261 304
rect 259 303 260 304
rect 258 303 259 304
rect 257 303 258 304
rect 256 303 257 304
rect 255 303 256 304
rect 254 303 255 304
rect 253 303 254 304
rect 252 303 253 304
rect 251 303 252 304
rect 250 303 251 304
rect 249 303 250 304
rect 248 303 249 304
rect 247 303 248 304
rect 246 303 247 304
rect 245 303 246 304
rect 244 303 245 304
rect 243 303 244 304
rect 242 303 243 304
rect 241 303 242 304
rect 240 303 241 304
rect 239 303 240 304
rect 238 303 239 304
rect 237 303 238 304
rect 236 303 237 304
rect 235 303 236 304
rect 234 303 235 304
rect 233 303 234 304
rect 232 303 233 304
rect 231 303 232 304
rect 230 303 231 304
rect 229 303 230 304
rect 228 303 229 304
rect 227 303 228 304
rect 226 303 227 304
rect 225 303 226 304
rect 224 303 225 304
rect 223 303 224 304
rect 222 303 223 304
rect 221 303 222 304
rect 220 303 221 304
rect 219 303 220 304
rect 218 303 219 304
rect 217 303 218 304
rect 216 303 217 304
rect 215 303 216 304
rect 214 303 215 304
rect 213 303 214 304
rect 212 303 213 304
rect 211 303 212 304
rect 210 303 211 304
rect 209 303 210 304
rect 208 303 209 304
rect 207 303 208 304
rect 206 303 207 304
rect 205 303 206 304
rect 204 303 205 304
rect 203 303 204 304
rect 202 303 203 304
rect 171 303 172 304
rect 170 303 171 304
rect 169 303 170 304
rect 168 303 169 304
rect 167 303 168 304
rect 166 303 167 304
rect 165 303 166 304
rect 164 303 165 304
rect 163 303 164 304
rect 162 303 163 304
rect 161 303 162 304
rect 160 303 161 304
rect 159 303 160 304
rect 158 303 159 304
rect 157 303 158 304
rect 156 303 157 304
rect 155 303 156 304
rect 154 303 155 304
rect 153 303 154 304
rect 152 303 153 304
rect 151 303 152 304
rect 122 303 123 304
rect 121 303 122 304
rect 120 303 121 304
rect 119 303 120 304
rect 118 303 119 304
rect 117 303 118 304
rect 116 303 117 304
rect 115 303 116 304
rect 114 303 115 304
rect 113 303 114 304
rect 112 303 113 304
rect 111 303 112 304
rect 110 303 111 304
rect 109 303 110 304
rect 108 303 109 304
rect 107 303 108 304
rect 106 303 107 304
rect 105 303 106 304
rect 104 303 105 304
rect 103 303 104 304
rect 102 303 103 304
rect 101 303 102 304
rect 100 303 101 304
rect 99 303 100 304
rect 98 303 99 304
rect 97 303 98 304
rect 96 303 97 304
rect 95 303 96 304
rect 94 303 95 304
rect 93 303 94 304
rect 92 303 93 304
rect 91 303 92 304
rect 90 303 91 304
rect 89 303 90 304
rect 88 303 89 304
rect 87 303 88 304
rect 86 303 87 304
rect 85 303 86 304
rect 68 303 69 304
rect 67 303 68 304
rect 66 303 67 304
rect 65 303 66 304
rect 64 303 65 304
rect 63 303 64 304
rect 62 303 63 304
rect 61 303 62 304
rect 60 303 61 304
rect 59 303 60 304
rect 58 303 59 304
rect 57 303 58 304
rect 56 303 57 304
rect 55 303 56 304
rect 54 303 55 304
rect 53 303 54 304
rect 52 303 53 304
rect 51 303 52 304
rect 50 303 51 304
rect 49 303 50 304
rect 48 303 49 304
rect 47 303 48 304
rect 46 303 47 304
rect 45 303 46 304
rect 44 303 45 304
rect 43 303 44 304
rect 42 303 43 304
rect 41 303 42 304
rect 40 303 41 304
rect 29 303 30 304
rect 28 303 29 304
rect 27 303 28 304
rect 26 303 27 304
rect 25 303 26 304
rect 24 303 25 304
rect 23 303 24 304
rect 22 303 23 304
rect 21 303 22 304
rect 20 303 21 304
rect 19 303 20 304
rect 18 303 19 304
rect 17 303 18 304
rect 16 303 17 304
rect 15 303 16 304
rect 14 303 15 304
rect 13 303 14 304
rect 12 303 13 304
rect 11 303 12 304
rect 10 303 11 304
rect 9 303 10 304
rect 8 303 9 304
rect 7 303 8 304
rect 6 303 7 304
rect 5 303 6 304
rect 437 304 438 305
rect 436 304 437 305
rect 435 304 436 305
rect 415 304 416 305
rect 414 304 415 305
rect 413 304 414 305
rect 412 304 413 305
rect 395 304 396 305
rect 394 304 395 305
rect 393 304 394 305
rect 259 304 260 305
rect 258 304 259 305
rect 257 304 258 305
rect 256 304 257 305
rect 255 304 256 305
rect 254 304 255 305
rect 253 304 254 305
rect 252 304 253 305
rect 251 304 252 305
rect 250 304 251 305
rect 249 304 250 305
rect 248 304 249 305
rect 247 304 248 305
rect 246 304 247 305
rect 245 304 246 305
rect 244 304 245 305
rect 243 304 244 305
rect 242 304 243 305
rect 241 304 242 305
rect 240 304 241 305
rect 239 304 240 305
rect 238 304 239 305
rect 237 304 238 305
rect 236 304 237 305
rect 235 304 236 305
rect 234 304 235 305
rect 233 304 234 305
rect 232 304 233 305
rect 231 304 232 305
rect 230 304 231 305
rect 229 304 230 305
rect 228 304 229 305
rect 227 304 228 305
rect 226 304 227 305
rect 225 304 226 305
rect 224 304 225 305
rect 223 304 224 305
rect 222 304 223 305
rect 221 304 222 305
rect 220 304 221 305
rect 219 304 220 305
rect 218 304 219 305
rect 217 304 218 305
rect 216 304 217 305
rect 215 304 216 305
rect 214 304 215 305
rect 213 304 214 305
rect 212 304 213 305
rect 211 304 212 305
rect 210 304 211 305
rect 209 304 210 305
rect 208 304 209 305
rect 207 304 208 305
rect 206 304 207 305
rect 205 304 206 305
rect 204 304 205 305
rect 203 304 204 305
rect 202 304 203 305
rect 201 304 202 305
rect 168 304 169 305
rect 167 304 168 305
rect 166 304 167 305
rect 165 304 166 305
rect 164 304 165 305
rect 163 304 164 305
rect 162 304 163 305
rect 161 304 162 305
rect 160 304 161 305
rect 159 304 160 305
rect 158 304 159 305
rect 157 304 158 305
rect 156 304 157 305
rect 155 304 156 305
rect 154 304 155 305
rect 123 304 124 305
rect 122 304 123 305
rect 121 304 122 305
rect 120 304 121 305
rect 119 304 120 305
rect 118 304 119 305
rect 117 304 118 305
rect 116 304 117 305
rect 115 304 116 305
rect 114 304 115 305
rect 113 304 114 305
rect 112 304 113 305
rect 111 304 112 305
rect 110 304 111 305
rect 109 304 110 305
rect 108 304 109 305
rect 107 304 108 305
rect 106 304 107 305
rect 105 304 106 305
rect 104 304 105 305
rect 103 304 104 305
rect 102 304 103 305
rect 101 304 102 305
rect 100 304 101 305
rect 99 304 100 305
rect 98 304 99 305
rect 97 304 98 305
rect 96 304 97 305
rect 95 304 96 305
rect 94 304 95 305
rect 93 304 94 305
rect 92 304 93 305
rect 91 304 92 305
rect 90 304 91 305
rect 89 304 90 305
rect 88 304 89 305
rect 87 304 88 305
rect 86 304 87 305
rect 85 304 86 305
rect 69 304 70 305
rect 68 304 69 305
rect 67 304 68 305
rect 66 304 67 305
rect 65 304 66 305
rect 64 304 65 305
rect 63 304 64 305
rect 62 304 63 305
rect 61 304 62 305
rect 60 304 61 305
rect 59 304 60 305
rect 58 304 59 305
rect 57 304 58 305
rect 56 304 57 305
rect 55 304 56 305
rect 54 304 55 305
rect 53 304 54 305
rect 52 304 53 305
rect 51 304 52 305
rect 50 304 51 305
rect 49 304 50 305
rect 48 304 49 305
rect 47 304 48 305
rect 46 304 47 305
rect 45 304 46 305
rect 44 304 45 305
rect 43 304 44 305
rect 42 304 43 305
rect 41 304 42 305
rect 40 304 41 305
rect 29 304 30 305
rect 28 304 29 305
rect 27 304 28 305
rect 26 304 27 305
rect 25 304 26 305
rect 24 304 25 305
rect 23 304 24 305
rect 22 304 23 305
rect 21 304 22 305
rect 20 304 21 305
rect 19 304 20 305
rect 18 304 19 305
rect 17 304 18 305
rect 16 304 17 305
rect 15 304 16 305
rect 14 304 15 305
rect 13 304 14 305
rect 12 304 13 305
rect 11 304 12 305
rect 10 304 11 305
rect 9 304 10 305
rect 8 304 9 305
rect 7 304 8 305
rect 6 304 7 305
rect 437 305 438 306
rect 436 305 437 306
rect 435 305 436 306
rect 434 305 435 306
rect 415 305 416 306
rect 414 305 415 306
rect 413 305 414 306
rect 412 305 413 306
rect 397 305 398 306
rect 396 305 397 306
rect 395 305 396 306
rect 394 305 395 306
rect 393 305 394 306
rect 257 305 258 306
rect 256 305 257 306
rect 255 305 256 306
rect 254 305 255 306
rect 253 305 254 306
rect 252 305 253 306
rect 251 305 252 306
rect 250 305 251 306
rect 249 305 250 306
rect 248 305 249 306
rect 247 305 248 306
rect 246 305 247 306
rect 245 305 246 306
rect 244 305 245 306
rect 243 305 244 306
rect 242 305 243 306
rect 241 305 242 306
rect 240 305 241 306
rect 239 305 240 306
rect 238 305 239 306
rect 237 305 238 306
rect 236 305 237 306
rect 235 305 236 306
rect 234 305 235 306
rect 233 305 234 306
rect 232 305 233 306
rect 231 305 232 306
rect 230 305 231 306
rect 229 305 230 306
rect 228 305 229 306
rect 227 305 228 306
rect 226 305 227 306
rect 225 305 226 306
rect 224 305 225 306
rect 223 305 224 306
rect 222 305 223 306
rect 221 305 222 306
rect 220 305 221 306
rect 219 305 220 306
rect 218 305 219 306
rect 217 305 218 306
rect 216 305 217 306
rect 215 305 216 306
rect 214 305 215 306
rect 213 305 214 306
rect 212 305 213 306
rect 211 305 212 306
rect 210 305 211 306
rect 209 305 210 306
rect 208 305 209 306
rect 207 305 208 306
rect 206 305 207 306
rect 205 305 206 306
rect 204 305 205 306
rect 203 305 204 306
rect 202 305 203 306
rect 201 305 202 306
rect 162 305 163 306
rect 161 305 162 306
rect 160 305 161 306
rect 123 305 124 306
rect 122 305 123 306
rect 121 305 122 306
rect 120 305 121 306
rect 119 305 120 306
rect 118 305 119 306
rect 117 305 118 306
rect 116 305 117 306
rect 115 305 116 306
rect 114 305 115 306
rect 113 305 114 306
rect 112 305 113 306
rect 111 305 112 306
rect 110 305 111 306
rect 109 305 110 306
rect 108 305 109 306
rect 107 305 108 306
rect 106 305 107 306
rect 105 305 106 306
rect 104 305 105 306
rect 103 305 104 306
rect 102 305 103 306
rect 101 305 102 306
rect 100 305 101 306
rect 99 305 100 306
rect 98 305 99 306
rect 97 305 98 306
rect 96 305 97 306
rect 95 305 96 306
rect 94 305 95 306
rect 93 305 94 306
rect 92 305 93 306
rect 91 305 92 306
rect 90 305 91 306
rect 89 305 90 306
rect 88 305 89 306
rect 87 305 88 306
rect 86 305 87 306
rect 69 305 70 306
rect 68 305 69 306
rect 67 305 68 306
rect 66 305 67 306
rect 65 305 66 306
rect 64 305 65 306
rect 63 305 64 306
rect 62 305 63 306
rect 61 305 62 306
rect 60 305 61 306
rect 59 305 60 306
rect 58 305 59 306
rect 57 305 58 306
rect 56 305 57 306
rect 55 305 56 306
rect 54 305 55 306
rect 53 305 54 306
rect 52 305 53 306
rect 51 305 52 306
rect 50 305 51 306
rect 49 305 50 306
rect 48 305 49 306
rect 47 305 48 306
rect 46 305 47 306
rect 45 305 46 306
rect 44 305 45 306
rect 43 305 44 306
rect 42 305 43 306
rect 41 305 42 306
rect 30 305 31 306
rect 29 305 30 306
rect 28 305 29 306
rect 27 305 28 306
rect 26 305 27 306
rect 25 305 26 306
rect 24 305 25 306
rect 23 305 24 306
rect 22 305 23 306
rect 21 305 22 306
rect 20 305 21 306
rect 19 305 20 306
rect 18 305 19 306
rect 17 305 18 306
rect 16 305 17 306
rect 15 305 16 306
rect 14 305 15 306
rect 13 305 14 306
rect 12 305 13 306
rect 11 305 12 306
rect 10 305 11 306
rect 9 305 10 306
rect 8 305 9 306
rect 7 305 8 306
rect 6 305 7 306
rect 437 306 438 307
rect 436 306 437 307
rect 435 306 436 307
rect 434 306 435 307
rect 433 306 434 307
rect 432 306 433 307
rect 431 306 432 307
rect 430 306 431 307
rect 429 306 430 307
rect 428 306 429 307
rect 427 306 428 307
rect 426 306 427 307
rect 425 306 426 307
rect 424 306 425 307
rect 423 306 424 307
rect 422 306 423 307
rect 421 306 422 307
rect 420 306 421 307
rect 419 306 420 307
rect 418 306 419 307
rect 417 306 418 307
rect 416 306 417 307
rect 415 306 416 307
rect 414 306 415 307
rect 413 306 414 307
rect 412 306 413 307
rect 411 306 412 307
rect 410 306 411 307
rect 409 306 410 307
rect 408 306 409 307
rect 407 306 408 307
rect 406 306 407 307
rect 405 306 406 307
rect 404 306 405 307
rect 403 306 404 307
rect 402 306 403 307
rect 401 306 402 307
rect 400 306 401 307
rect 399 306 400 307
rect 398 306 399 307
rect 397 306 398 307
rect 396 306 397 307
rect 395 306 396 307
rect 394 306 395 307
rect 393 306 394 307
rect 256 306 257 307
rect 255 306 256 307
rect 254 306 255 307
rect 253 306 254 307
rect 252 306 253 307
rect 251 306 252 307
rect 250 306 251 307
rect 249 306 250 307
rect 248 306 249 307
rect 247 306 248 307
rect 246 306 247 307
rect 245 306 246 307
rect 244 306 245 307
rect 243 306 244 307
rect 242 306 243 307
rect 241 306 242 307
rect 240 306 241 307
rect 239 306 240 307
rect 238 306 239 307
rect 237 306 238 307
rect 236 306 237 307
rect 235 306 236 307
rect 234 306 235 307
rect 233 306 234 307
rect 232 306 233 307
rect 231 306 232 307
rect 230 306 231 307
rect 229 306 230 307
rect 228 306 229 307
rect 227 306 228 307
rect 226 306 227 307
rect 225 306 226 307
rect 224 306 225 307
rect 223 306 224 307
rect 222 306 223 307
rect 221 306 222 307
rect 220 306 221 307
rect 219 306 220 307
rect 218 306 219 307
rect 217 306 218 307
rect 216 306 217 307
rect 215 306 216 307
rect 214 306 215 307
rect 213 306 214 307
rect 212 306 213 307
rect 211 306 212 307
rect 210 306 211 307
rect 209 306 210 307
rect 208 306 209 307
rect 207 306 208 307
rect 206 306 207 307
rect 205 306 206 307
rect 204 306 205 307
rect 203 306 204 307
rect 202 306 203 307
rect 201 306 202 307
rect 200 306 201 307
rect 124 306 125 307
rect 123 306 124 307
rect 122 306 123 307
rect 121 306 122 307
rect 120 306 121 307
rect 119 306 120 307
rect 118 306 119 307
rect 117 306 118 307
rect 116 306 117 307
rect 115 306 116 307
rect 114 306 115 307
rect 113 306 114 307
rect 112 306 113 307
rect 111 306 112 307
rect 110 306 111 307
rect 109 306 110 307
rect 108 306 109 307
rect 107 306 108 307
rect 106 306 107 307
rect 105 306 106 307
rect 104 306 105 307
rect 103 306 104 307
rect 102 306 103 307
rect 101 306 102 307
rect 100 306 101 307
rect 99 306 100 307
rect 98 306 99 307
rect 97 306 98 307
rect 96 306 97 307
rect 95 306 96 307
rect 94 306 95 307
rect 93 306 94 307
rect 92 306 93 307
rect 91 306 92 307
rect 90 306 91 307
rect 89 306 90 307
rect 88 306 89 307
rect 87 306 88 307
rect 86 306 87 307
rect 70 306 71 307
rect 69 306 70 307
rect 68 306 69 307
rect 67 306 68 307
rect 66 306 67 307
rect 65 306 66 307
rect 64 306 65 307
rect 63 306 64 307
rect 62 306 63 307
rect 61 306 62 307
rect 60 306 61 307
rect 59 306 60 307
rect 58 306 59 307
rect 57 306 58 307
rect 56 306 57 307
rect 55 306 56 307
rect 54 306 55 307
rect 53 306 54 307
rect 52 306 53 307
rect 51 306 52 307
rect 50 306 51 307
rect 49 306 50 307
rect 48 306 49 307
rect 47 306 48 307
rect 46 306 47 307
rect 45 306 46 307
rect 44 306 45 307
rect 43 306 44 307
rect 42 306 43 307
rect 41 306 42 307
rect 30 306 31 307
rect 29 306 30 307
rect 28 306 29 307
rect 27 306 28 307
rect 26 306 27 307
rect 25 306 26 307
rect 24 306 25 307
rect 23 306 24 307
rect 22 306 23 307
rect 21 306 22 307
rect 20 306 21 307
rect 19 306 20 307
rect 18 306 19 307
rect 17 306 18 307
rect 16 306 17 307
rect 15 306 16 307
rect 14 306 15 307
rect 13 306 14 307
rect 12 306 13 307
rect 11 306 12 307
rect 10 306 11 307
rect 9 306 10 307
rect 8 306 9 307
rect 7 306 8 307
rect 437 307 438 308
rect 436 307 437 308
rect 435 307 436 308
rect 434 307 435 308
rect 433 307 434 308
rect 432 307 433 308
rect 431 307 432 308
rect 430 307 431 308
rect 429 307 430 308
rect 428 307 429 308
rect 427 307 428 308
rect 426 307 427 308
rect 425 307 426 308
rect 424 307 425 308
rect 423 307 424 308
rect 422 307 423 308
rect 421 307 422 308
rect 420 307 421 308
rect 419 307 420 308
rect 418 307 419 308
rect 417 307 418 308
rect 416 307 417 308
rect 415 307 416 308
rect 414 307 415 308
rect 413 307 414 308
rect 412 307 413 308
rect 411 307 412 308
rect 410 307 411 308
rect 409 307 410 308
rect 408 307 409 308
rect 407 307 408 308
rect 406 307 407 308
rect 405 307 406 308
rect 404 307 405 308
rect 403 307 404 308
rect 402 307 403 308
rect 401 307 402 308
rect 400 307 401 308
rect 399 307 400 308
rect 398 307 399 308
rect 397 307 398 308
rect 396 307 397 308
rect 395 307 396 308
rect 394 307 395 308
rect 393 307 394 308
rect 254 307 255 308
rect 253 307 254 308
rect 252 307 253 308
rect 251 307 252 308
rect 250 307 251 308
rect 249 307 250 308
rect 248 307 249 308
rect 247 307 248 308
rect 246 307 247 308
rect 245 307 246 308
rect 244 307 245 308
rect 243 307 244 308
rect 242 307 243 308
rect 241 307 242 308
rect 240 307 241 308
rect 239 307 240 308
rect 238 307 239 308
rect 237 307 238 308
rect 236 307 237 308
rect 235 307 236 308
rect 234 307 235 308
rect 233 307 234 308
rect 232 307 233 308
rect 231 307 232 308
rect 230 307 231 308
rect 229 307 230 308
rect 228 307 229 308
rect 227 307 228 308
rect 226 307 227 308
rect 225 307 226 308
rect 224 307 225 308
rect 223 307 224 308
rect 222 307 223 308
rect 221 307 222 308
rect 220 307 221 308
rect 219 307 220 308
rect 218 307 219 308
rect 217 307 218 308
rect 216 307 217 308
rect 215 307 216 308
rect 214 307 215 308
rect 213 307 214 308
rect 212 307 213 308
rect 211 307 212 308
rect 210 307 211 308
rect 209 307 210 308
rect 208 307 209 308
rect 207 307 208 308
rect 206 307 207 308
rect 205 307 206 308
rect 204 307 205 308
rect 203 307 204 308
rect 202 307 203 308
rect 201 307 202 308
rect 200 307 201 308
rect 199 307 200 308
rect 125 307 126 308
rect 124 307 125 308
rect 123 307 124 308
rect 122 307 123 308
rect 121 307 122 308
rect 120 307 121 308
rect 119 307 120 308
rect 118 307 119 308
rect 117 307 118 308
rect 116 307 117 308
rect 115 307 116 308
rect 114 307 115 308
rect 113 307 114 308
rect 112 307 113 308
rect 111 307 112 308
rect 110 307 111 308
rect 109 307 110 308
rect 108 307 109 308
rect 107 307 108 308
rect 106 307 107 308
rect 105 307 106 308
rect 104 307 105 308
rect 103 307 104 308
rect 102 307 103 308
rect 101 307 102 308
rect 100 307 101 308
rect 99 307 100 308
rect 98 307 99 308
rect 97 307 98 308
rect 96 307 97 308
rect 95 307 96 308
rect 94 307 95 308
rect 93 307 94 308
rect 92 307 93 308
rect 91 307 92 308
rect 90 307 91 308
rect 89 307 90 308
rect 88 307 89 308
rect 87 307 88 308
rect 70 307 71 308
rect 69 307 70 308
rect 68 307 69 308
rect 67 307 68 308
rect 66 307 67 308
rect 65 307 66 308
rect 64 307 65 308
rect 63 307 64 308
rect 62 307 63 308
rect 61 307 62 308
rect 60 307 61 308
rect 59 307 60 308
rect 58 307 59 308
rect 57 307 58 308
rect 56 307 57 308
rect 55 307 56 308
rect 54 307 55 308
rect 53 307 54 308
rect 52 307 53 308
rect 51 307 52 308
rect 50 307 51 308
rect 49 307 50 308
rect 48 307 49 308
rect 47 307 48 308
rect 46 307 47 308
rect 45 307 46 308
rect 44 307 45 308
rect 43 307 44 308
rect 42 307 43 308
rect 41 307 42 308
rect 30 307 31 308
rect 29 307 30 308
rect 28 307 29 308
rect 27 307 28 308
rect 26 307 27 308
rect 25 307 26 308
rect 24 307 25 308
rect 23 307 24 308
rect 22 307 23 308
rect 21 307 22 308
rect 20 307 21 308
rect 19 307 20 308
rect 18 307 19 308
rect 17 307 18 308
rect 16 307 17 308
rect 15 307 16 308
rect 14 307 15 308
rect 13 307 14 308
rect 12 307 13 308
rect 11 307 12 308
rect 10 307 11 308
rect 9 307 10 308
rect 8 307 9 308
rect 437 308 438 309
rect 436 308 437 309
rect 435 308 436 309
rect 434 308 435 309
rect 433 308 434 309
rect 432 308 433 309
rect 431 308 432 309
rect 430 308 431 309
rect 429 308 430 309
rect 428 308 429 309
rect 427 308 428 309
rect 426 308 427 309
rect 425 308 426 309
rect 424 308 425 309
rect 423 308 424 309
rect 422 308 423 309
rect 421 308 422 309
rect 420 308 421 309
rect 419 308 420 309
rect 418 308 419 309
rect 417 308 418 309
rect 416 308 417 309
rect 415 308 416 309
rect 414 308 415 309
rect 413 308 414 309
rect 412 308 413 309
rect 411 308 412 309
rect 410 308 411 309
rect 409 308 410 309
rect 408 308 409 309
rect 407 308 408 309
rect 406 308 407 309
rect 405 308 406 309
rect 404 308 405 309
rect 403 308 404 309
rect 402 308 403 309
rect 401 308 402 309
rect 400 308 401 309
rect 399 308 400 309
rect 398 308 399 309
rect 397 308 398 309
rect 396 308 397 309
rect 395 308 396 309
rect 394 308 395 309
rect 393 308 394 309
rect 252 308 253 309
rect 251 308 252 309
rect 250 308 251 309
rect 249 308 250 309
rect 248 308 249 309
rect 247 308 248 309
rect 246 308 247 309
rect 245 308 246 309
rect 244 308 245 309
rect 243 308 244 309
rect 242 308 243 309
rect 241 308 242 309
rect 240 308 241 309
rect 239 308 240 309
rect 238 308 239 309
rect 237 308 238 309
rect 236 308 237 309
rect 235 308 236 309
rect 234 308 235 309
rect 233 308 234 309
rect 232 308 233 309
rect 231 308 232 309
rect 230 308 231 309
rect 229 308 230 309
rect 228 308 229 309
rect 227 308 228 309
rect 226 308 227 309
rect 225 308 226 309
rect 224 308 225 309
rect 223 308 224 309
rect 222 308 223 309
rect 221 308 222 309
rect 220 308 221 309
rect 219 308 220 309
rect 218 308 219 309
rect 217 308 218 309
rect 216 308 217 309
rect 215 308 216 309
rect 214 308 215 309
rect 213 308 214 309
rect 212 308 213 309
rect 211 308 212 309
rect 210 308 211 309
rect 209 308 210 309
rect 208 308 209 309
rect 207 308 208 309
rect 206 308 207 309
rect 205 308 206 309
rect 204 308 205 309
rect 203 308 204 309
rect 202 308 203 309
rect 201 308 202 309
rect 200 308 201 309
rect 199 308 200 309
rect 198 308 199 309
rect 126 308 127 309
rect 125 308 126 309
rect 124 308 125 309
rect 123 308 124 309
rect 122 308 123 309
rect 121 308 122 309
rect 120 308 121 309
rect 119 308 120 309
rect 118 308 119 309
rect 117 308 118 309
rect 116 308 117 309
rect 115 308 116 309
rect 114 308 115 309
rect 113 308 114 309
rect 112 308 113 309
rect 111 308 112 309
rect 110 308 111 309
rect 109 308 110 309
rect 108 308 109 309
rect 107 308 108 309
rect 106 308 107 309
rect 105 308 106 309
rect 104 308 105 309
rect 103 308 104 309
rect 102 308 103 309
rect 101 308 102 309
rect 100 308 101 309
rect 99 308 100 309
rect 98 308 99 309
rect 97 308 98 309
rect 96 308 97 309
rect 95 308 96 309
rect 94 308 95 309
rect 93 308 94 309
rect 92 308 93 309
rect 91 308 92 309
rect 90 308 91 309
rect 89 308 90 309
rect 88 308 89 309
rect 87 308 88 309
rect 70 308 71 309
rect 69 308 70 309
rect 68 308 69 309
rect 67 308 68 309
rect 66 308 67 309
rect 65 308 66 309
rect 64 308 65 309
rect 63 308 64 309
rect 62 308 63 309
rect 61 308 62 309
rect 60 308 61 309
rect 59 308 60 309
rect 58 308 59 309
rect 57 308 58 309
rect 56 308 57 309
rect 55 308 56 309
rect 54 308 55 309
rect 53 308 54 309
rect 52 308 53 309
rect 51 308 52 309
rect 50 308 51 309
rect 49 308 50 309
rect 48 308 49 309
rect 47 308 48 309
rect 46 308 47 309
rect 45 308 46 309
rect 44 308 45 309
rect 43 308 44 309
rect 42 308 43 309
rect 30 308 31 309
rect 29 308 30 309
rect 28 308 29 309
rect 27 308 28 309
rect 26 308 27 309
rect 25 308 26 309
rect 24 308 25 309
rect 23 308 24 309
rect 22 308 23 309
rect 21 308 22 309
rect 20 308 21 309
rect 19 308 20 309
rect 18 308 19 309
rect 17 308 18 309
rect 16 308 17 309
rect 15 308 16 309
rect 14 308 15 309
rect 13 308 14 309
rect 12 308 13 309
rect 11 308 12 309
rect 10 308 11 309
rect 9 308 10 309
rect 8 308 9 309
rect 437 309 438 310
rect 436 309 437 310
rect 435 309 436 310
rect 434 309 435 310
rect 433 309 434 310
rect 432 309 433 310
rect 431 309 432 310
rect 430 309 431 310
rect 429 309 430 310
rect 428 309 429 310
rect 427 309 428 310
rect 426 309 427 310
rect 425 309 426 310
rect 424 309 425 310
rect 423 309 424 310
rect 422 309 423 310
rect 421 309 422 310
rect 420 309 421 310
rect 419 309 420 310
rect 418 309 419 310
rect 417 309 418 310
rect 416 309 417 310
rect 415 309 416 310
rect 414 309 415 310
rect 413 309 414 310
rect 412 309 413 310
rect 411 309 412 310
rect 410 309 411 310
rect 409 309 410 310
rect 408 309 409 310
rect 407 309 408 310
rect 406 309 407 310
rect 405 309 406 310
rect 404 309 405 310
rect 403 309 404 310
rect 402 309 403 310
rect 401 309 402 310
rect 400 309 401 310
rect 399 309 400 310
rect 398 309 399 310
rect 397 309 398 310
rect 396 309 397 310
rect 395 309 396 310
rect 394 309 395 310
rect 393 309 394 310
rect 251 309 252 310
rect 250 309 251 310
rect 249 309 250 310
rect 248 309 249 310
rect 247 309 248 310
rect 246 309 247 310
rect 245 309 246 310
rect 244 309 245 310
rect 243 309 244 310
rect 242 309 243 310
rect 241 309 242 310
rect 240 309 241 310
rect 239 309 240 310
rect 238 309 239 310
rect 237 309 238 310
rect 236 309 237 310
rect 235 309 236 310
rect 234 309 235 310
rect 233 309 234 310
rect 232 309 233 310
rect 231 309 232 310
rect 230 309 231 310
rect 229 309 230 310
rect 228 309 229 310
rect 227 309 228 310
rect 226 309 227 310
rect 225 309 226 310
rect 224 309 225 310
rect 223 309 224 310
rect 222 309 223 310
rect 221 309 222 310
rect 220 309 221 310
rect 219 309 220 310
rect 218 309 219 310
rect 217 309 218 310
rect 216 309 217 310
rect 215 309 216 310
rect 214 309 215 310
rect 213 309 214 310
rect 212 309 213 310
rect 211 309 212 310
rect 210 309 211 310
rect 209 309 210 310
rect 208 309 209 310
rect 207 309 208 310
rect 206 309 207 310
rect 205 309 206 310
rect 204 309 205 310
rect 203 309 204 310
rect 202 309 203 310
rect 201 309 202 310
rect 200 309 201 310
rect 199 309 200 310
rect 198 309 199 310
rect 197 309 198 310
rect 127 309 128 310
rect 126 309 127 310
rect 125 309 126 310
rect 124 309 125 310
rect 123 309 124 310
rect 122 309 123 310
rect 121 309 122 310
rect 120 309 121 310
rect 119 309 120 310
rect 118 309 119 310
rect 117 309 118 310
rect 116 309 117 310
rect 115 309 116 310
rect 114 309 115 310
rect 113 309 114 310
rect 112 309 113 310
rect 111 309 112 310
rect 110 309 111 310
rect 109 309 110 310
rect 108 309 109 310
rect 107 309 108 310
rect 106 309 107 310
rect 105 309 106 310
rect 104 309 105 310
rect 103 309 104 310
rect 102 309 103 310
rect 101 309 102 310
rect 100 309 101 310
rect 99 309 100 310
rect 98 309 99 310
rect 97 309 98 310
rect 96 309 97 310
rect 95 309 96 310
rect 94 309 95 310
rect 93 309 94 310
rect 92 309 93 310
rect 91 309 92 310
rect 90 309 91 310
rect 89 309 90 310
rect 88 309 89 310
rect 71 309 72 310
rect 70 309 71 310
rect 69 309 70 310
rect 68 309 69 310
rect 67 309 68 310
rect 66 309 67 310
rect 65 309 66 310
rect 64 309 65 310
rect 63 309 64 310
rect 62 309 63 310
rect 61 309 62 310
rect 60 309 61 310
rect 59 309 60 310
rect 58 309 59 310
rect 57 309 58 310
rect 56 309 57 310
rect 55 309 56 310
rect 54 309 55 310
rect 53 309 54 310
rect 52 309 53 310
rect 51 309 52 310
rect 50 309 51 310
rect 49 309 50 310
rect 48 309 49 310
rect 47 309 48 310
rect 46 309 47 310
rect 45 309 46 310
rect 44 309 45 310
rect 43 309 44 310
rect 42 309 43 310
rect 31 309 32 310
rect 30 309 31 310
rect 29 309 30 310
rect 28 309 29 310
rect 27 309 28 310
rect 26 309 27 310
rect 25 309 26 310
rect 24 309 25 310
rect 23 309 24 310
rect 22 309 23 310
rect 21 309 22 310
rect 20 309 21 310
rect 19 309 20 310
rect 18 309 19 310
rect 17 309 18 310
rect 16 309 17 310
rect 15 309 16 310
rect 14 309 15 310
rect 13 309 14 310
rect 12 309 13 310
rect 11 309 12 310
rect 10 309 11 310
rect 9 309 10 310
rect 458 310 459 311
rect 437 310 438 311
rect 436 310 437 311
rect 435 310 436 311
rect 434 310 435 311
rect 433 310 434 311
rect 432 310 433 311
rect 431 310 432 311
rect 430 310 431 311
rect 429 310 430 311
rect 428 310 429 311
rect 427 310 428 311
rect 426 310 427 311
rect 425 310 426 311
rect 424 310 425 311
rect 423 310 424 311
rect 422 310 423 311
rect 421 310 422 311
rect 420 310 421 311
rect 419 310 420 311
rect 418 310 419 311
rect 417 310 418 311
rect 416 310 417 311
rect 415 310 416 311
rect 414 310 415 311
rect 413 310 414 311
rect 412 310 413 311
rect 411 310 412 311
rect 410 310 411 311
rect 409 310 410 311
rect 408 310 409 311
rect 407 310 408 311
rect 406 310 407 311
rect 405 310 406 311
rect 404 310 405 311
rect 403 310 404 311
rect 402 310 403 311
rect 401 310 402 311
rect 400 310 401 311
rect 399 310 400 311
rect 398 310 399 311
rect 397 310 398 311
rect 396 310 397 311
rect 395 310 396 311
rect 394 310 395 311
rect 393 310 394 311
rect 249 310 250 311
rect 248 310 249 311
rect 247 310 248 311
rect 246 310 247 311
rect 245 310 246 311
rect 244 310 245 311
rect 243 310 244 311
rect 242 310 243 311
rect 241 310 242 311
rect 240 310 241 311
rect 239 310 240 311
rect 238 310 239 311
rect 237 310 238 311
rect 236 310 237 311
rect 235 310 236 311
rect 234 310 235 311
rect 233 310 234 311
rect 232 310 233 311
rect 231 310 232 311
rect 230 310 231 311
rect 229 310 230 311
rect 228 310 229 311
rect 227 310 228 311
rect 226 310 227 311
rect 225 310 226 311
rect 224 310 225 311
rect 223 310 224 311
rect 222 310 223 311
rect 221 310 222 311
rect 220 310 221 311
rect 219 310 220 311
rect 218 310 219 311
rect 217 310 218 311
rect 216 310 217 311
rect 215 310 216 311
rect 214 310 215 311
rect 213 310 214 311
rect 212 310 213 311
rect 211 310 212 311
rect 210 310 211 311
rect 209 310 210 311
rect 208 310 209 311
rect 207 310 208 311
rect 206 310 207 311
rect 205 310 206 311
rect 204 310 205 311
rect 203 310 204 311
rect 202 310 203 311
rect 201 310 202 311
rect 200 310 201 311
rect 199 310 200 311
rect 198 310 199 311
rect 197 310 198 311
rect 196 310 197 311
rect 128 310 129 311
rect 127 310 128 311
rect 126 310 127 311
rect 125 310 126 311
rect 124 310 125 311
rect 123 310 124 311
rect 122 310 123 311
rect 121 310 122 311
rect 120 310 121 311
rect 119 310 120 311
rect 118 310 119 311
rect 117 310 118 311
rect 116 310 117 311
rect 115 310 116 311
rect 114 310 115 311
rect 113 310 114 311
rect 112 310 113 311
rect 111 310 112 311
rect 110 310 111 311
rect 109 310 110 311
rect 108 310 109 311
rect 107 310 108 311
rect 106 310 107 311
rect 105 310 106 311
rect 104 310 105 311
rect 103 310 104 311
rect 102 310 103 311
rect 101 310 102 311
rect 100 310 101 311
rect 99 310 100 311
rect 98 310 99 311
rect 97 310 98 311
rect 96 310 97 311
rect 95 310 96 311
rect 94 310 95 311
rect 93 310 94 311
rect 92 310 93 311
rect 91 310 92 311
rect 90 310 91 311
rect 89 310 90 311
rect 71 310 72 311
rect 70 310 71 311
rect 69 310 70 311
rect 68 310 69 311
rect 67 310 68 311
rect 66 310 67 311
rect 65 310 66 311
rect 64 310 65 311
rect 63 310 64 311
rect 62 310 63 311
rect 61 310 62 311
rect 60 310 61 311
rect 59 310 60 311
rect 58 310 59 311
rect 57 310 58 311
rect 56 310 57 311
rect 55 310 56 311
rect 54 310 55 311
rect 53 310 54 311
rect 52 310 53 311
rect 51 310 52 311
rect 50 310 51 311
rect 49 310 50 311
rect 48 310 49 311
rect 47 310 48 311
rect 46 310 47 311
rect 45 310 46 311
rect 44 310 45 311
rect 43 310 44 311
rect 42 310 43 311
rect 31 310 32 311
rect 30 310 31 311
rect 29 310 30 311
rect 28 310 29 311
rect 27 310 28 311
rect 26 310 27 311
rect 25 310 26 311
rect 24 310 25 311
rect 23 310 24 311
rect 22 310 23 311
rect 21 310 22 311
rect 20 310 21 311
rect 19 310 20 311
rect 18 310 19 311
rect 17 310 18 311
rect 16 310 17 311
rect 15 310 16 311
rect 14 310 15 311
rect 13 310 14 311
rect 12 310 13 311
rect 11 310 12 311
rect 10 310 11 311
rect 458 311 459 312
rect 437 311 438 312
rect 436 311 437 312
rect 435 311 436 312
rect 434 311 435 312
rect 433 311 434 312
rect 432 311 433 312
rect 431 311 432 312
rect 430 311 431 312
rect 429 311 430 312
rect 428 311 429 312
rect 427 311 428 312
rect 426 311 427 312
rect 425 311 426 312
rect 424 311 425 312
rect 423 311 424 312
rect 422 311 423 312
rect 421 311 422 312
rect 420 311 421 312
rect 419 311 420 312
rect 418 311 419 312
rect 417 311 418 312
rect 416 311 417 312
rect 415 311 416 312
rect 414 311 415 312
rect 413 311 414 312
rect 412 311 413 312
rect 411 311 412 312
rect 410 311 411 312
rect 409 311 410 312
rect 408 311 409 312
rect 407 311 408 312
rect 406 311 407 312
rect 405 311 406 312
rect 404 311 405 312
rect 403 311 404 312
rect 402 311 403 312
rect 401 311 402 312
rect 400 311 401 312
rect 399 311 400 312
rect 398 311 399 312
rect 397 311 398 312
rect 396 311 397 312
rect 395 311 396 312
rect 394 311 395 312
rect 393 311 394 312
rect 247 311 248 312
rect 246 311 247 312
rect 245 311 246 312
rect 244 311 245 312
rect 243 311 244 312
rect 242 311 243 312
rect 241 311 242 312
rect 240 311 241 312
rect 239 311 240 312
rect 238 311 239 312
rect 237 311 238 312
rect 236 311 237 312
rect 235 311 236 312
rect 234 311 235 312
rect 233 311 234 312
rect 232 311 233 312
rect 231 311 232 312
rect 230 311 231 312
rect 229 311 230 312
rect 228 311 229 312
rect 227 311 228 312
rect 226 311 227 312
rect 225 311 226 312
rect 224 311 225 312
rect 223 311 224 312
rect 222 311 223 312
rect 221 311 222 312
rect 220 311 221 312
rect 219 311 220 312
rect 218 311 219 312
rect 217 311 218 312
rect 216 311 217 312
rect 215 311 216 312
rect 214 311 215 312
rect 213 311 214 312
rect 212 311 213 312
rect 211 311 212 312
rect 210 311 211 312
rect 209 311 210 312
rect 208 311 209 312
rect 207 311 208 312
rect 206 311 207 312
rect 205 311 206 312
rect 204 311 205 312
rect 203 311 204 312
rect 202 311 203 312
rect 201 311 202 312
rect 200 311 201 312
rect 199 311 200 312
rect 198 311 199 312
rect 197 311 198 312
rect 196 311 197 312
rect 195 311 196 312
rect 129 311 130 312
rect 128 311 129 312
rect 127 311 128 312
rect 126 311 127 312
rect 125 311 126 312
rect 124 311 125 312
rect 123 311 124 312
rect 122 311 123 312
rect 121 311 122 312
rect 120 311 121 312
rect 119 311 120 312
rect 118 311 119 312
rect 117 311 118 312
rect 116 311 117 312
rect 115 311 116 312
rect 114 311 115 312
rect 113 311 114 312
rect 112 311 113 312
rect 111 311 112 312
rect 110 311 111 312
rect 109 311 110 312
rect 108 311 109 312
rect 107 311 108 312
rect 106 311 107 312
rect 105 311 106 312
rect 104 311 105 312
rect 103 311 104 312
rect 102 311 103 312
rect 101 311 102 312
rect 100 311 101 312
rect 99 311 100 312
rect 98 311 99 312
rect 97 311 98 312
rect 96 311 97 312
rect 95 311 96 312
rect 94 311 95 312
rect 93 311 94 312
rect 92 311 93 312
rect 91 311 92 312
rect 90 311 91 312
rect 89 311 90 312
rect 72 311 73 312
rect 71 311 72 312
rect 70 311 71 312
rect 69 311 70 312
rect 68 311 69 312
rect 67 311 68 312
rect 66 311 67 312
rect 65 311 66 312
rect 64 311 65 312
rect 63 311 64 312
rect 62 311 63 312
rect 61 311 62 312
rect 60 311 61 312
rect 59 311 60 312
rect 58 311 59 312
rect 57 311 58 312
rect 56 311 57 312
rect 55 311 56 312
rect 54 311 55 312
rect 53 311 54 312
rect 52 311 53 312
rect 51 311 52 312
rect 50 311 51 312
rect 49 311 50 312
rect 48 311 49 312
rect 47 311 48 312
rect 46 311 47 312
rect 45 311 46 312
rect 44 311 45 312
rect 43 311 44 312
rect 31 311 32 312
rect 30 311 31 312
rect 29 311 30 312
rect 28 311 29 312
rect 27 311 28 312
rect 26 311 27 312
rect 25 311 26 312
rect 24 311 25 312
rect 23 311 24 312
rect 22 311 23 312
rect 21 311 22 312
rect 20 311 21 312
rect 19 311 20 312
rect 18 311 19 312
rect 17 311 18 312
rect 16 311 17 312
rect 15 311 16 312
rect 14 311 15 312
rect 13 311 14 312
rect 12 311 13 312
rect 11 311 12 312
rect 10 311 11 312
rect 459 312 460 313
rect 458 312 459 313
rect 437 312 438 313
rect 436 312 437 313
rect 435 312 436 313
rect 434 312 435 313
rect 433 312 434 313
rect 432 312 433 313
rect 431 312 432 313
rect 430 312 431 313
rect 429 312 430 313
rect 428 312 429 313
rect 427 312 428 313
rect 426 312 427 313
rect 425 312 426 313
rect 424 312 425 313
rect 423 312 424 313
rect 422 312 423 313
rect 421 312 422 313
rect 420 312 421 313
rect 419 312 420 313
rect 418 312 419 313
rect 417 312 418 313
rect 416 312 417 313
rect 415 312 416 313
rect 414 312 415 313
rect 413 312 414 313
rect 412 312 413 313
rect 411 312 412 313
rect 410 312 411 313
rect 409 312 410 313
rect 408 312 409 313
rect 407 312 408 313
rect 406 312 407 313
rect 405 312 406 313
rect 404 312 405 313
rect 403 312 404 313
rect 402 312 403 313
rect 401 312 402 313
rect 400 312 401 313
rect 399 312 400 313
rect 398 312 399 313
rect 397 312 398 313
rect 396 312 397 313
rect 395 312 396 313
rect 394 312 395 313
rect 393 312 394 313
rect 245 312 246 313
rect 244 312 245 313
rect 243 312 244 313
rect 242 312 243 313
rect 241 312 242 313
rect 240 312 241 313
rect 239 312 240 313
rect 238 312 239 313
rect 237 312 238 313
rect 236 312 237 313
rect 235 312 236 313
rect 234 312 235 313
rect 233 312 234 313
rect 232 312 233 313
rect 231 312 232 313
rect 230 312 231 313
rect 229 312 230 313
rect 228 312 229 313
rect 227 312 228 313
rect 226 312 227 313
rect 225 312 226 313
rect 224 312 225 313
rect 223 312 224 313
rect 222 312 223 313
rect 221 312 222 313
rect 220 312 221 313
rect 219 312 220 313
rect 218 312 219 313
rect 217 312 218 313
rect 216 312 217 313
rect 215 312 216 313
rect 214 312 215 313
rect 213 312 214 313
rect 212 312 213 313
rect 211 312 212 313
rect 210 312 211 313
rect 209 312 210 313
rect 208 312 209 313
rect 207 312 208 313
rect 206 312 207 313
rect 205 312 206 313
rect 204 312 205 313
rect 203 312 204 313
rect 202 312 203 313
rect 201 312 202 313
rect 200 312 201 313
rect 199 312 200 313
rect 198 312 199 313
rect 197 312 198 313
rect 196 312 197 313
rect 195 312 196 313
rect 194 312 195 313
rect 130 312 131 313
rect 129 312 130 313
rect 128 312 129 313
rect 127 312 128 313
rect 126 312 127 313
rect 125 312 126 313
rect 124 312 125 313
rect 123 312 124 313
rect 122 312 123 313
rect 121 312 122 313
rect 120 312 121 313
rect 119 312 120 313
rect 118 312 119 313
rect 117 312 118 313
rect 116 312 117 313
rect 115 312 116 313
rect 114 312 115 313
rect 113 312 114 313
rect 112 312 113 313
rect 111 312 112 313
rect 110 312 111 313
rect 109 312 110 313
rect 108 312 109 313
rect 107 312 108 313
rect 106 312 107 313
rect 105 312 106 313
rect 104 312 105 313
rect 103 312 104 313
rect 102 312 103 313
rect 101 312 102 313
rect 100 312 101 313
rect 99 312 100 313
rect 98 312 99 313
rect 97 312 98 313
rect 96 312 97 313
rect 95 312 96 313
rect 94 312 95 313
rect 93 312 94 313
rect 92 312 93 313
rect 91 312 92 313
rect 90 312 91 313
rect 72 312 73 313
rect 71 312 72 313
rect 70 312 71 313
rect 69 312 70 313
rect 68 312 69 313
rect 67 312 68 313
rect 66 312 67 313
rect 65 312 66 313
rect 64 312 65 313
rect 63 312 64 313
rect 62 312 63 313
rect 61 312 62 313
rect 60 312 61 313
rect 59 312 60 313
rect 58 312 59 313
rect 57 312 58 313
rect 56 312 57 313
rect 55 312 56 313
rect 54 312 55 313
rect 53 312 54 313
rect 52 312 53 313
rect 51 312 52 313
rect 50 312 51 313
rect 49 312 50 313
rect 48 312 49 313
rect 47 312 48 313
rect 46 312 47 313
rect 45 312 46 313
rect 44 312 45 313
rect 43 312 44 313
rect 31 312 32 313
rect 30 312 31 313
rect 29 312 30 313
rect 28 312 29 313
rect 27 312 28 313
rect 26 312 27 313
rect 25 312 26 313
rect 24 312 25 313
rect 23 312 24 313
rect 22 312 23 313
rect 21 312 22 313
rect 20 312 21 313
rect 19 312 20 313
rect 18 312 19 313
rect 17 312 18 313
rect 16 312 17 313
rect 15 312 16 313
rect 14 312 15 313
rect 13 312 14 313
rect 12 312 13 313
rect 11 312 12 313
rect 461 313 462 314
rect 460 313 461 314
rect 459 313 460 314
rect 458 313 459 314
rect 437 313 438 314
rect 436 313 437 314
rect 435 313 436 314
rect 434 313 435 314
rect 433 313 434 314
rect 432 313 433 314
rect 431 313 432 314
rect 430 313 431 314
rect 429 313 430 314
rect 428 313 429 314
rect 427 313 428 314
rect 426 313 427 314
rect 425 313 426 314
rect 424 313 425 314
rect 423 313 424 314
rect 422 313 423 314
rect 421 313 422 314
rect 420 313 421 314
rect 419 313 420 314
rect 418 313 419 314
rect 417 313 418 314
rect 416 313 417 314
rect 415 313 416 314
rect 414 313 415 314
rect 413 313 414 314
rect 412 313 413 314
rect 411 313 412 314
rect 410 313 411 314
rect 409 313 410 314
rect 408 313 409 314
rect 407 313 408 314
rect 406 313 407 314
rect 405 313 406 314
rect 404 313 405 314
rect 403 313 404 314
rect 402 313 403 314
rect 401 313 402 314
rect 400 313 401 314
rect 399 313 400 314
rect 398 313 399 314
rect 397 313 398 314
rect 396 313 397 314
rect 395 313 396 314
rect 394 313 395 314
rect 393 313 394 314
rect 243 313 244 314
rect 242 313 243 314
rect 241 313 242 314
rect 240 313 241 314
rect 239 313 240 314
rect 238 313 239 314
rect 237 313 238 314
rect 236 313 237 314
rect 235 313 236 314
rect 234 313 235 314
rect 233 313 234 314
rect 232 313 233 314
rect 231 313 232 314
rect 230 313 231 314
rect 229 313 230 314
rect 228 313 229 314
rect 227 313 228 314
rect 226 313 227 314
rect 225 313 226 314
rect 224 313 225 314
rect 223 313 224 314
rect 222 313 223 314
rect 221 313 222 314
rect 220 313 221 314
rect 219 313 220 314
rect 218 313 219 314
rect 217 313 218 314
rect 216 313 217 314
rect 215 313 216 314
rect 214 313 215 314
rect 213 313 214 314
rect 212 313 213 314
rect 211 313 212 314
rect 210 313 211 314
rect 209 313 210 314
rect 208 313 209 314
rect 207 313 208 314
rect 206 313 207 314
rect 205 313 206 314
rect 204 313 205 314
rect 203 313 204 314
rect 202 313 203 314
rect 201 313 202 314
rect 200 313 201 314
rect 199 313 200 314
rect 198 313 199 314
rect 197 313 198 314
rect 196 313 197 314
rect 195 313 196 314
rect 194 313 195 314
rect 193 313 194 314
rect 131 313 132 314
rect 130 313 131 314
rect 129 313 130 314
rect 128 313 129 314
rect 127 313 128 314
rect 126 313 127 314
rect 125 313 126 314
rect 124 313 125 314
rect 123 313 124 314
rect 122 313 123 314
rect 121 313 122 314
rect 120 313 121 314
rect 119 313 120 314
rect 118 313 119 314
rect 117 313 118 314
rect 116 313 117 314
rect 115 313 116 314
rect 114 313 115 314
rect 113 313 114 314
rect 112 313 113 314
rect 111 313 112 314
rect 110 313 111 314
rect 109 313 110 314
rect 108 313 109 314
rect 107 313 108 314
rect 106 313 107 314
rect 105 313 106 314
rect 104 313 105 314
rect 103 313 104 314
rect 102 313 103 314
rect 101 313 102 314
rect 100 313 101 314
rect 99 313 100 314
rect 98 313 99 314
rect 97 313 98 314
rect 96 313 97 314
rect 95 313 96 314
rect 94 313 95 314
rect 93 313 94 314
rect 92 313 93 314
rect 91 313 92 314
rect 90 313 91 314
rect 73 313 74 314
rect 72 313 73 314
rect 71 313 72 314
rect 70 313 71 314
rect 69 313 70 314
rect 68 313 69 314
rect 67 313 68 314
rect 66 313 67 314
rect 65 313 66 314
rect 64 313 65 314
rect 63 313 64 314
rect 62 313 63 314
rect 61 313 62 314
rect 60 313 61 314
rect 59 313 60 314
rect 58 313 59 314
rect 57 313 58 314
rect 56 313 57 314
rect 55 313 56 314
rect 54 313 55 314
rect 53 313 54 314
rect 52 313 53 314
rect 51 313 52 314
rect 50 313 51 314
rect 49 313 50 314
rect 48 313 49 314
rect 47 313 48 314
rect 46 313 47 314
rect 45 313 46 314
rect 44 313 45 314
rect 43 313 44 314
rect 32 313 33 314
rect 31 313 32 314
rect 30 313 31 314
rect 29 313 30 314
rect 28 313 29 314
rect 27 313 28 314
rect 26 313 27 314
rect 25 313 26 314
rect 24 313 25 314
rect 23 313 24 314
rect 22 313 23 314
rect 21 313 22 314
rect 20 313 21 314
rect 19 313 20 314
rect 18 313 19 314
rect 17 313 18 314
rect 16 313 17 314
rect 15 313 16 314
rect 14 313 15 314
rect 13 313 14 314
rect 12 313 13 314
rect 11 313 12 314
rect 463 314 464 315
rect 462 314 463 315
rect 461 314 462 315
rect 460 314 461 315
rect 459 314 460 315
rect 458 314 459 315
rect 437 314 438 315
rect 436 314 437 315
rect 435 314 436 315
rect 434 314 435 315
rect 433 314 434 315
rect 432 314 433 315
rect 431 314 432 315
rect 430 314 431 315
rect 429 314 430 315
rect 428 314 429 315
rect 427 314 428 315
rect 426 314 427 315
rect 425 314 426 315
rect 424 314 425 315
rect 423 314 424 315
rect 422 314 423 315
rect 421 314 422 315
rect 420 314 421 315
rect 419 314 420 315
rect 418 314 419 315
rect 417 314 418 315
rect 416 314 417 315
rect 415 314 416 315
rect 414 314 415 315
rect 413 314 414 315
rect 412 314 413 315
rect 411 314 412 315
rect 410 314 411 315
rect 409 314 410 315
rect 408 314 409 315
rect 407 314 408 315
rect 406 314 407 315
rect 405 314 406 315
rect 404 314 405 315
rect 403 314 404 315
rect 402 314 403 315
rect 401 314 402 315
rect 400 314 401 315
rect 399 314 400 315
rect 398 314 399 315
rect 397 314 398 315
rect 396 314 397 315
rect 395 314 396 315
rect 394 314 395 315
rect 393 314 394 315
rect 240 314 241 315
rect 239 314 240 315
rect 238 314 239 315
rect 237 314 238 315
rect 236 314 237 315
rect 235 314 236 315
rect 234 314 235 315
rect 233 314 234 315
rect 232 314 233 315
rect 231 314 232 315
rect 230 314 231 315
rect 229 314 230 315
rect 228 314 229 315
rect 227 314 228 315
rect 226 314 227 315
rect 225 314 226 315
rect 224 314 225 315
rect 223 314 224 315
rect 222 314 223 315
rect 221 314 222 315
rect 220 314 221 315
rect 219 314 220 315
rect 218 314 219 315
rect 217 314 218 315
rect 216 314 217 315
rect 215 314 216 315
rect 214 314 215 315
rect 213 314 214 315
rect 212 314 213 315
rect 211 314 212 315
rect 210 314 211 315
rect 209 314 210 315
rect 208 314 209 315
rect 207 314 208 315
rect 206 314 207 315
rect 205 314 206 315
rect 204 314 205 315
rect 203 314 204 315
rect 202 314 203 315
rect 201 314 202 315
rect 200 314 201 315
rect 199 314 200 315
rect 198 314 199 315
rect 197 314 198 315
rect 196 314 197 315
rect 195 314 196 315
rect 194 314 195 315
rect 193 314 194 315
rect 192 314 193 315
rect 132 314 133 315
rect 131 314 132 315
rect 130 314 131 315
rect 129 314 130 315
rect 128 314 129 315
rect 127 314 128 315
rect 126 314 127 315
rect 125 314 126 315
rect 124 314 125 315
rect 123 314 124 315
rect 122 314 123 315
rect 121 314 122 315
rect 120 314 121 315
rect 119 314 120 315
rect 118 314 119 315
rect 117 314 118 315
rect 116 314 117 315
rect 115 314 116 315
rect 114 314 115 315
rect 113 314 114 315
rect 112 314 113 315
rect 111 314 112 315
rect 110 314 111 315
rect 109 314 110 315
rect 108 314 109 315
rect 107 314 108 315
rect 106 314 107 315
rect 105 314 106 315
rect 104 314 105 315
rect 103 314 104 315
rect 102 314 103 315
rect 101 314 102 315
rect 100 314 101 315
rect 99 314 100 315
rect 98 314 99 315
rect 97 314 98 315
rect 96 314 97 315
rect 95 314 96 315
rect 94 314 95 315
rect 93 314 94 315
rect 92 314 93 315
rect 91 314 92 315
rect 73 314 74 315
rect 72 314 73 315
rect 71 314 72 315
rect 70 314 71 315
rect 69 314 70 315
rect 68 314 69 315
rect 67 314 68 315
rect 66 314 67 315
rect 65 314 66 315
rect 64 314 65 315
rect 63 314 64 315
rect 62 314 63 315
rect 61 314 62 315
rect 60 314 61 315
rect 59 314 60 315
rect 58 314 59 315
rect 57 314 58 315
rect 56 314 57 315
rect 55 314 56 315
rect 54 314 55 315
rect 53 314 54 315
rect 52 314 53 315
rect 51 314 52 315
rect 50 314 51 315
rect 49 314 50 315
rect 48 314 49 315
rect 47 314 48 315
rect 46 314 47 315
rect 45 314 46 315
rect 44 314 45 315
rect 32 314 33 315
rect 31 314 32 315
rect 30 314 31 315
rect 29 314 30 315
rect 28 314 29 315
rect 27 314 28 315
rect 26 314 27 315
rect 25 314 26 315
rect 24 314 25 315
rect 23 314 24 315
rect 22 314 23 315
rect 21 314 22 315
rect 20 314 21 315
rect 19 314 20 315
rect 18 314 19 315
rect 17 314 18 315
rect 16 314 17 315
rect 15 314 16 315
rect 14 314 15 315
rect 13 314 14 315
rect 12 314 13 315
rect 478 315 479 316
rect 464 315 465 316
rect 463 315 464 316
rect 462 315 463 316
rect 461 315 462 316
rect 460 315 461 316
rect 459 315 460 316
rect 458 315 459 316
rect 437 315 438 316
rect 436 315 437 316
rect 435 315 436 316
rect 434 315 435 316
rect 433 315 434 316
rect 432 315 433 316
rect 431 315 432 316
rect 430 315 431 316
rect 429 315 430 316
rect 428 315 429 316
rect 427 315 428 316
rect 426 315 427 316
rect 425 315 426 316
rect 424 315 425 316
rect 423 315 424 316
rect 422 315 423 316
rect 421 315 422 316
rect 420 315 421 316
rect 419 315 420 316
rect 418 315 419 316
rect 417 315 418 316
rect 416 315 417 316
rect 415 315 416 316
rect 414 315 415 316
rect 413 315 414 316
rect 412 315 413 316
rect 411 315 412 316
rect 410 315 411 316
rect 409 315 410 316
rect 408 315 409 316
rect 407 315 408 316
rect 406 315 407 316
rect 405 315 406 316
rect 404 315 405 316
rect 403 315 404 316
rect 402 315 403 316
rect 401 315 402 316
rect 400 315 401 316
rect 399 315 400 316
rect 398 315 399 316
rect 397 315 398 316
rect 396 315 397 316
rect 395 315 396 316
rect 394 315 395 316
rect 393 315 394 316
rect 238 315 239 316
rect 237 315 238 316
rect 236 315 237 316
rect 235 315 236 316
rect 234 315 235 316
rect 233 315 234 316
rect 232 315 233 316
rect 231 315 232 316
rect 230 315 231 316
rect 229 315 230 316
rect 228 315 229 316
rect 227 315 228 316
rect 226 315 227 316
rect 225 315 226 316
rect 224 315 225 316
rect 223 315 224 316
rect 222 315 223 316
rect 221 315 222 316
rect 220 315 221 316
rect 219 315 220 316
rect 218 315 219 316
rect 217 315 218 316
rect 216 315 217 316
rect 215 315 216 316
rect 214 315 215 316
rect 213 315 214 316
rect 212 315 213 316
rect 211 315 212 316
rect 210 315 211 316
rect 209 315 210 316
rect 208 315 209 316
rect 207 315 208 316
rect 206 315 207 316
rect 205 315 206 316
rect 204 315 205 316
rect 203 315 204 316
rect 202 315 203 316
rect 201 315 202 316
rect 200 315 201 316
rect 199 315 200 316
rect 198 315 199 316
rect 197 315 198 316
rect 196 315 197 316
rect 195 315 196 316
rect 194 315 195 316
rect 193 315 194 316
rect 192 315 193 316
rect 191 315 192 316
rect 134 315 135 316
rect 133 315 134 316
rect 132 315 133 316
rect 131 315 132 316
rect 130 315 131 316
rect 129 315 130 316
rect 128 315 129 316
rect 127 315 128 316
rect 126 315 127 316
rect 125 315 126 316
rect 124 315 125 316
rect 123 315 124 316
rect 122 315 123 316
rect 121 315 122 316
rect 120 315 121 316
rect 119 315 120 316
rect 118 315 119 316
rect 117 315 118 316
rect 116 315 117 316
rect 115 315 116 316
rect 114 315 115 316
rect 113 315 114 316
rect 112 315 113 316
rect 111 315 112 316
rect 110 315 111 316
rect 109 315 110 316
rect 108 315 109 316
rect 107 315 108 316
rect 106 315 107 316
rect 105 315 106 316
rect 104 315 105 316
rect 103 315 104 316
rect 102 315 103 316
rect 101 315 102 316
rect 100 315 101 316
rect 99 315 100 316
rect 98 315 99 316
rect 97 315 98 316
rect 96 315 97 316
rect 95 315 96 316
rect 94 315 95 316
rect 93 315 94 316
rect 92 315 93 316
rect 74 315 75 316
rect 73 315 74 316
rect 72 315 73 316
rect 71 315 72 316
rect 70 315 71 316
rect 69 315 70 316
rect 68 315 69 316
rect 67 315 68 316
rect 66 315 67 316
rect 65 315 66 316
rect 64 315 65 316
rect 63 315 64 316
rect 62 315 63 316
rect 61 315 62 316
rect 60 315 61 316
rect 59 315 60 316
rect 58 315 59 316
rect 57 315 58 316
rect 56 315 57 316
rect 55 315 56 316
rect 54 315 55 316
rect 53 315 54 316
rect 52 315 53 316
rect 51 315 52 316
rect 50 315 51 316
rect 49 315 50 316
rect 48 315 49 316
rect 47 315 48 316
rect 46 315 47 316
rect 45 315 46 316
rect 44 315 45 316
rect 32 315 33 316
rect 31 315 32 316
rect 30 315 31 316
rect 29 315 30 316
rect 28 315 29 316
rect 27 315 28 316
rect 26 315 27 316
rect 25 315 26 316
rect 24 315 25 316
rect 23 315 24 316
rect 22 315 23 316
rect 21 315 22 316
rect 20 315 21 316
rect 19 315 20 316
rect 18 315 19 316
rect 17 315 18 316
rect 16 315 17 316
rect 15 315 16 316
rect 14 315 15 316
rect 13 315 14 316
rect 478 316 479 317
rect 466 316 467 317
rect 465 316 466 317
rect 464 316 465 317
rect 463 316 464 317
rect 462 316 463 317
rect 461 316 462 317
rect 460 316 461 317
rect 459 316 460 317
rect 458 316 459 317
rect 437 316 438 317
rect 436 316 437 317
rect 435 316 436 317
rect 434 316 435 317
rect 396 316 397 317
rect 395 316 396 317
rect 394 316 395 317
rect 393 316 394 317
rect 235 316 236 317
rect 234 316 235 317
rect 233 316 234 317
rect 232 316 233 317
rect 231 316 232 317
rect 230 316 231 317
rect 229 316 230 317
rect 228 316 229 317
rect 227 316 228 317
rect 226 316 227 317
rect 225 316 226 317
rect 224 316 225 317
rect 223 316 224 317
rect 222 316 223 317
rect 221 316 222 317
rect 220 316 221 317
rect 219 316 220 317
rect 218 316 219 317
rect 217 316 218 317
rect 216 316 217 317
rect 215 316 216 317
rect 214 316 215 317
rect 213 316 214 317
rect 212 316 213 317
rect 211 316 212 317
rect 210 316 211 317
rect 209 316 210 317
rect 208 316 209 317
rect 207 316 208 317
rect 206 316 207 317
rect 205 316 206 317
rect 204 316 205 317
rect 203 316 204 317
rect 202 316 203 317
rect 201 316 202 317
rect 200 316 201 317
rect 199 316 200 317
rect 198 316 199 317
rect 197 316 198 317
rect 196 316 197 317
rect 195 316 196 317
rect 194 316 195 317
rect 193 316 194 317
rect 192 316 193 317
rect 191 316 192 317
rect 190 316 191 317
rect 135 316 136 317
rect 134 316 135 317
rect 133 316 134 317
rect 132 316 133 317
rect 131 316 132 317
rect 130 316 131 317
rect 129 316 130 317
rect 128 316 129 317
rect 127 316 128 317
rect 126 316 127 317
rect 125 316 126 317
rect 124 316 125 317
rect 123 316 124 317
rect 122 316 123 317
rect 121 316 122 317
rect 120 316 121 317
rect 119 316 120 317
rect 118 316 119 317
rect 117 316 118 317
rect 116 316 117 317
rect 115 316 116 317
rect 114 316 115 317
rect 113 316 114 317
rect 112 316 113 317
rect 111 316 112 317
rect 110 316 111 317
rect 109 316 110 317
rect 108 316 109 317
rect 107 316 108 317
rect 106 316 107 317
rect 105 316 106 317
rect 104 316 105 317
rect 103 316 104 317
rect 102 316 103 317
rect 101 316 102 317
rect 100 316 101 317
rect 99 316 100 317
rect 98 316 99 317
rect 97 316 98 317
rect 96 316 97 317
rect 95 316 96 317
rect 94 316 95 317
rect 93 316 94 317
rect 92 316 93 317
rect 74 316 75 317
rect 73 316 74 317
rect 72 316 73 317
rect 71 316 72 317
rect 70 316 71 317
rect 69 316 70 317
rect 68 316 69 317
rect 67 316 68 317
rect 66 316 67 317
rect 65 316 66 317
rect 64 316 65 317
rect 63 316 64 317
rect 62 316 63 317
rect 61 316 62 317
rect 60 316 61 317
rect 59 316 60 317
rect 58 316 59 317
rect 57 316 58 317
rect 56 316 57 317
rect 55 316 56 317
rect 54 316 55 317
rect 53 316 54 317
rect 52 316 53 317
rect 51 316 52 317
rect 50 316 51 317
rect 49 316 50 317
rect 48 316 49 317
rect 47 316 48 317
rect 46 316 47 317
rect 45 316 46 317
rect 44 316 45 317
rect 33 316 34 317
rect 32 316 33 317
rect 31 316 32 317
rect 30 316 31 317
rect 29 316 30 317
rect 28 316 29 317
rect 27 316 28 317
rect 26 316 27 317
rect 25 316 26 317
rect 24 316 25 317
rect 23 316 24 317
rect 22 316 23 317
rect 21 316 22 317
rect 20 316 21 317
rect 19 316 20 317
rect 18 316 19 317
rect 17 316 18 317
rect 16 316 17 317
rect 15 316 16 317
rect 14 316 15 317
rect 478 317 479 318
rect 477 317 478 318
rect 468 317 469 318
rect 467 317 468 318
rect 466 317 467 318
rect 465 317 466 318
rect 464 317 465 318
rect 463 317 464 318
rect 462 317 463 318
rect 461 317 462 318
rect 460 317 461 318
rect 459 317 460 318
rect 458 317 459 318
rect 437 317 438 318
rect 436 317 437 318
rect 435 317 436 318
rect 395 317 396 318
rect 394 317 395 318
rect 393 317 394 318
rect 232 317 233 318
rect 231 317 232 318
rect 230 317 231 318
rect 229 317 230 318
rect 228 317 229 318
rect 227 317 228 318
rect 226 317 227 318
rect 225 317 226 318
rect 224 317 225 318
rect 223 317 224 318
rect 222 317 223 318
rect 221 317 222 318
rect 220 317 221 318
rect 219 317 220 318
rect 218 317 219 318
rect 217 317 218 318
rect 216 317 217 318
rect 215 317 216 318
rect 214 317 215 318
rect 213 317 214 318
rect 212 317 213 318
rect 211 317 212 318
rect 210 317 211 318
rect 209 317 210 318
rect 208 317 209 318
rect 207 317 208 318
rect 206 317 207 318
rect 205 317 206 318
rect 204 317 205 318
rect 203 317 204 318
rect 202 317 203 318
rect 201 317 202 318
rect 200 317 201 318
rect 199 317 200 318
rect 198 317 199 318
rect 197 317 198 318
rect 196 317 197 318
rect 195 317 196 318
rect 194 317 195 318
rect 193 317 194 318
rect 192 317 193 318
rect 191 317 192 318
rect 190 317 191 318
rect 189 317 190 318
rect 136 317 137 318
rect 135 317 136 318
rect 134 317 135 318
rect 133 317 134 318
rect 132 317 133 318
rect 131 317 132 318
rect 130 317 131 318
rect 129 317 130 318
rect 128 317 129 318
rect 127 317 128 318
rect 126 317 127 318
rect 125 317 126 318
rect 124 317 125 318
rect 123 317 124 318
rect 122 317 123 318
rect 121 317 122 318
rect 120 317 121 318
rect 119 317 120 318
rect 118 317 119 318
rect 117 317 118 318
rect 116 317 117 318
rect 115 317 116 318
rect 114 317 115 318
rect 113 317 114 318
rect 112 317 113 318
rect 111 317 112 318
rect 110 317 111 318
rect 109 317 110 318
rect 108 317 109 318
rect 107 317 108 318
rect 106 317 107 318
rect 105 317 106 318
rect 104 317 105 318
rect 103 317 104 318
rect 102 317 103 318
rect 101 317 102 318
rect 100 317 101 318
rect 99 317 100 318
rect 98 317 99 318
rect 97 317 98 318
rect 96 317 97 318
rect 95 317 96 318
rect 94 317 95 318
rect 93 317 94 318
rect 75 317 76 318
rect 74 317 75 318
rect 73 317 74 318
rect 72 317 73 318
rect 71 317 72 318
rect 70 317 71 318
rect 69 317 70 318
rect 68 317 69 318
rect 67 317 68 318
rect 66 317 67 318
rect 65 317 66 318
rect 64 317 65 318
rect 63 317 64 318
rect 62 317 63 318
rect 61 317 62 318
rect 60 317 61 318
rect 59 317 60 318
rect 58 317 59 318
rect 57 317 58 318
rect 56 317 57 318
rect 55 317 56 318
rect 54 317 55 318
rect 53 317 54 318
rect 52 317 53 318
rect 51 317 52 318
rect 50 317 51 318
rect 49 317 50 318
rect 48 317 49 318
rect 47 317 48 318
rect 46 317 47 318
rect 45 317 46 318
rect 33 317 34 318
rect 32 317 33 318
rect 31 317 32 318
rect 30 317 31 318
rect 29 317 30 318
rect 28 317 29 318
rect 27 317 28 318
rect 26 317 27 318
rect 25 317 26 318
rect 24 317 25 318
rect 23 317 24 318
rect 22 317 23 318
rect 21 317 22 318
rect 20 317 21 318
rect 19 317 20 318
rect 18 317 19 318
rect 17 317 18 318
rect 16 317 17 318
rect 15 317 16 318
rect 14 317 15 318
rect 478 318 479 319
rect 477 318 478 319
rect 476 318 477 319
rect 475 318 476 319
rect 474 318 475 319
rect 473 318 474 319
rect 472 318 473 319
rect 471 318 472 319
rect 470 318 471 319
rect 469 318 470 319
rect 468 318 469 319
rect 467 318 468 319
rect 466 318 467 319
rect 465 318 466 319
rect 464 318 465 319
rect 463 318 464 319
rect 462 318 463 319
rect 458 318 459 319
rect 437 318 438 319
rect 436 318 437 319
rect 435 318 436 319
rect 395 318 396 319
rect 394 318 395 319
rect 393 318 394 319
rect 228 318 229 319
rect 227 318 228 319
rect 226 318 227 319
rect 225 318 226 319
rect 224 318 225 319
rect 223 318 224 319
rect 222 318 223 319
rect 221 318 222 319
rect 220 318 221 319
rect 219 318 220 319
rect 218 318 219 319
rect 217 318 218 319
rect 216 318 217 319
rect 215 318 216 319
rect 214 318 215 319
rect 213 318 214 319
rect 212 318 213 319
rect 211 318 212 319
rect 210 318 211 319
rect 209 318 210 319
rect 208 318 209 319
rect 207 318 208 319
rect 206 318 207 319
rect 205 318 206 319
rect 204 318 205 319
rect 203 318 204 319
rect 202 318 203 319
rect 201 318 202 319
rect 200 318 201 319
rect 199 318 200 319
rect 198 318 199 319
rect 197 318 198 319
rect 196 318 197 319
rect 195 318 196 319
rect 194 318 195 319
rect 193 318 194 319
rect 192 318 193 319
rect 191 318 192 319
rect 190 318 191 319
rect 189 318 190 319
rect 188 318 189 319
rect 138 318 139 319
rect 137 318 138 319
rect 136 318 137 319
rect 135 318 136 319
rect 134 318 135 319
rect 133 318 134 319
rect 132 318 133 319
rect 131 318 132 319
rect 130 318 131 319
rect 129 318 130 319
rect 128 318 129 319
rect 127 318 128 319
rect 126 318 127 319
rect 125 318 126 319
rect 124 318 125 319
rect 123 318 124 319
rect 122 318 123 319
rect 121 318 122 319
rect 120 318 121 319
rect 119 318 120 319
rect 118 318 119 319
rect 117 318 118 319
rect 116 318 117 319
rect 115 318 116 319
rect 114 318 115 319
rect 113 318 114 319
rect 112 318 113 319
rect 111 318 112 319
rect 110 318 111 319
rect 109 318 110 319
rect 108 318 109 319
rect 107 318 108 319
rect 106 318 107 319
rect 105 318 106 319
rect 104 318 105 319
rect 103 318 104 319
rect 102 318 103 319
rect 101 318 102 319
rect 100 318 101 319
rect 99 318 100 319
rect 98 318 99 319
rect 97 318 98 319
rect 96 318 97 319
rect 95 318 96 319
rect 94 318 95 319
rect 75 318 76 319
rect 74 318 75 319
rect 73 318 74 319
rect 72 318 73 319
rect 71 318 72 319
rect 70 318 71 319
rect 69 318 70 319
rect 68 318 69 319
rect 67 318 68 319
rect 66 318 67 319
rect 65 318 66 319
rect 64 318 65 319
rect 63 318 64 319
rect 62 318 63 319
rect 61 318 62 319
rect 60 318 61 319
rect 59 318 60 319
rect 58 318 59 319
rect 57 318 58 319
rect 56 318 57 319
rect 55 318 56 319
rect 54 318 55 319
rect 53 318 54 319
rect 52 318 53 319
rect 51 318 52 319
rect 50 318 51 319
rect 49 318 50 319
rect 48 318 49 319
rect 47 318 48 319
rect 46 318 47 319
rect 45 318 46 319
rect 33 318 34 319
rect 32 318 33 319
rect 31 318 32 319
rect 30 318 31 319
rect 29 318 30 319
rect 28 318 29 319
rect 27 318 28 319
rect 26 318 27 319
rect 25 318 26 319
rect 24 318 25 319
rect 23 318 24 319
rect 22 318 23 319
rect 21 318 22 319
rect 20 318 21 319
rect 19 318 20 319
rect 18 318 19 319
rect 17 318 18 319
rect 16 318 17 319
rect 15 318 16 319
rect 478 319 479 320
rect 477 319 478 320
rect 476 319 477 320
rect 475 319 476 320
rect 474 319 475 320
rect 473 319 474 320
rect 472 319 473 320
rect 471 319 472 320
rect 470 319 471 320
rect 469 319 470 320
rect 468 319 469 320
rect 467 319 468 320
rect 466 319 467 320
rect 465 319 466 320
rect 464 319 465 320
rect 458 319 459 320
rect 437 319 438 320
rect 436 319 437 320
rect 435 319 436 320
rect 395 319 396 320
rect 394 319 395 320
rect 393 319 394 320
rect 224 319 225 320
rect 223 319 224 320
rect 222 319 223 320
rect 221 319 222 320
rect 220 319 221 320
rect 219 319 220 320
rect 218 319 219 320
rect 217 319 218 320
rect 216 319 217 320
rect 215 319 216 320
rect 214 319 215 320
rect 213 319 214 320
rect 212 319 213 320
rect 211 319 212 320
rect 210 319 211 320
rect 209 319 210 320
rect 208 319 209 320
rect 207 319 208 320
rect 206 319 207 320
rect 205 319 206 320
rect 204 319 205 320
rect 203 319 204 320
rect 202 319 203 320
rect 201 319 202 320
rect 200 319 201 320
rect 199 319 200 320
rect 198 319 199 320
rect 197 319 198 320
rect 196 319 197 320
rect 195 319 196 320
rect 194 319 195 320
rect 193 319 194 320
rect 192 319 193 320
rect 191 319 192 320
rect 140 319 141 320
rect 139 319 140 320
rect 138 319 139 320
rect 137 319 138 320
rect 136 319 137 320
rect 135 319 136 320
rect 134 319 135 320
rect 133 319 134 320
rect 132 319 133 320
rect 131 319 132 320
rect 130 319 131 320
rect 129 319 130 320
rect 128 319 129 320
rect 127 319 128 320
rect 126 319 127 320
rect 125 319 126 320
rect 124 319 125 320
rect 123 319 124 320
rect 122 319 123 320
rect 121 319 122 320
rect 120 319 121 320
rect 119 319 120 320
rect 118 319 119 320
rect 117 319 118 320
rect 116 319 117 320
rect 115 319 116 320
rect 114 319 115 320
rect 113 319 114 320
rect 112 319 113 320
rect 111 319 112 320
rect 110 319 111 320
rect 109 319 110 320
rect 108 319 109 320
rect 107 319 108 320
rect 106 319 107 320
rect 105 319 106 320
rect 104 319 105 320
rect 103 319 104 320
rect 102 319 103 320
rect 101 319 102 320
rect 100 319 101 320
rect 99 319 100 320
rect 98 319 99 320
rect 97 319 98 320
rect 96 319 97 320
rect 95 319 96 320
rect 76 319 77 320
rect 75 319 76 320
rect 74 319 75 320
rect 73 319 74 320
rect 72 319 73 320
rect 71 319 72 320
rect 70 319 71 320
rect 69 319 70 320
rect 68 319 69 320
rect 67 319 68 320
rect 66 319 67 320
rect 65 319 66 320
rect 64 319 65 320
rect 63 319 64 320
rect 62 319 63 320
rect 61 319 62 320
rect 60 319 61 320
rect 59 319 60 320
rect 58 319 59 320
rect 57 319 58 320
rect 56 319 57 320
rect 55 319 56 320
rect 54 319 55 320
rect 53 319 54 320
rect 52 319 53 320
rect 51 319 52 320
rect 50 319 51 320
rect 49 319 50 320
rect 48 319 49 320
rect 47 319 48 320
rect 46 319 47 320
rect 45 319 46 320
rect 33 319 34 320
rect 32 319 33 320
rect 31 319 32 320
rect 30 319 31 320
rect 29 319 30 320
rect 28 319 29 320
rect 27 319 28 320
rect 26 319 27 320
rect 25 319 26 320
rect 24 319 25 320
rect 23 319 24 320
rect 22 319 23 320
rect 21 319 22 320
rect 20 319 21 320
rect 19 319 20 320
rect 18 319 19 320
rect 17 319 18 320
rect 16 319 17 320
rect 478 320 479 321
rect 477 320 478 321
rect 476 320 477 321
rect 475 320 476 321
rect 474 320 475 321
rect 473 320 474 321
rect 472 320 473 321
rect 471 320 472 321
rect 470 320 471 321
rect 469 320 470 321
rect 468 320 469 321
rect 467 320 468 321
rect 466 320 467 321
rect 437 320 438 321
rect 436 320 437 321
rect 435 320 436 321
rect 395 320 396 321
rect 394 320 395 321
rect 393 320 394 321
rect 217 320 218 321
rect 216 320 217 321
rect 215 320 216 321
rect 214 320 215 321
rect 213 320 214 321
rect 212 320 213 321
rect 211 320 212 321
rect 210 320 211 321
rect 209 320 210 321
rect 208 320 209 321
rect 207 320 208 321
rect 206 320 207 321
rect 205 320 206 321
rect 204 320 205 321
rect 203 320 204 321
rect 202 320 203 321
rect 201 320 202 321
rect 200 320 201 321
rect 199 320 200 321
rect 198 320 199 321
rect 141 320 142 321
rect 140 320 141 321
rect 139 320 140 321
rect 138 320 139 321
rect 137 320 138 321
rect 136 320 137 321
rect 135 320 136 321
rect 134 320 135 321
rect 133 320 134 321
rect 132 320 133 321
rect 131 320 132 321
rect 130 320 131 321
rect 129 320 130 321
rect 128 320 129 321
rect 127 320 128 321
rect 126 320 127 321
rect 125 320 126 321
rect 124 320 125 321
rect 123 320 124 321
rect 122 320 123 321
rect 121 320 122 321
rect 120 320 121 321
rect 119 320 120 321
rect 118 320 119 321
rect 117 320 118 321
rect 116 320 117 321
rect 115 320 116 321
rect 114 320 115 321
rect 113 320 114 321
rect 112 320 113 321
rect 111 320 112 321
rect 110 320 111 321
rect 109 320 110 321
rect 108 320 109 321
rect 107 320 108 321
rect 106 320 107 321
rect 105 320 106 321
rect 104 320 105 321
rect 103 320 104 321
rect 102 320 103 321
rect 101 320 102 321
rect 100 320 101 321
rect 99 320 100 321
rect 98 320 99 321
rect 97 320 98 321
rect 96 320 97 321
rect 95 320 96 321
rect 77 320 78 321
rect 76 320 77 321
rect 75 320 76 321
rect 74 320 75 321
rect 73 320 74 321
rect 72 320 73 321
rect 71 320 72 321
rect 70 320 71 321
rect 69 320 70 321
rect 68 320 69 321
rect 67 320 68 321
rect 66 320 67 321
rect 65 320 66 321
rect 64 320 65 321
rect 63 320 64 321
rect 62 320 63 321
rect 61 320 62 321
rect 60 320 61 321
rect 59 320 60 321
rect 58 320 59 321
rect 57 320 58 321
rect 56 320 57 321
rect 55 320 56 321
rect 54 320 55 321
rect 53 320 54 321
rect 52 320 53 321
rect 51 320 52 321
rect 50 320 51 321
rect 49 320 50 321
rect 48 320 49 321
rect 47 320 48 321
rect 46 320 47 321
rect 34 320 35 321
rect 33 320 34 321
rect 32 320 33 321
rect 31 320 32 321
rect 30 320 31 321
rect 29 320 30 321
rect 28 320 29 321
rect 27 320 28 321
rect 26 320 27 321
rect 25 320 26 321
rect 24 320 25 321
rect 23 320 24 321
rect 22 320 23 321
rect 21 320 22 321
rect 20 320 21 321
rect 19 320 20 321
rect 18 320 19 321
rect 17 320 18 321
rect 16 320 17 321
rect 478 321 479 322
rect 477 321 478 322
rect 476 321 477 322
rect 475 321 476 322
rect 474 321 475 322
rect 473 321 474 322
rect 472 321 473 322
rect 471 321 472 322
rect 470 321 471 322
rect 469 321 470 322
rect 468 321 469 322
rect 467 321 468 322
rect 143 321 144 322
rect 142 321 143 322
rect 141 321 142 322
rect 140 321 141 322
rect 139 321 140 322
rect 138 321 139 322
rect 137 321 138 322
rect 136 321 137 322
rect 135 321 136 322
rect 134 321 135 322
rect 133 321 134 322
rect 132 321 133 322
rect 131 321 132 322
rect 130 321 131 322
rect 129 321 130 322
rect 128 321 129 322
rect 127 321 128 322
rect 126 321 127 322
rect 125 321 126 322
rect 124 321 125 322
rect 123 321 124 322
rect 122 321 123 322
rect 121 321 122 322
rect 120 321 121 322
rect 119 321 120 322
rect 118 321 119 322
rect 117 321 118 322
rect 116 321 117 322
rect 115 321 116 322
rect 114 321 115 322
rect 113 321 114 322
rect 112 321 113 322
rect 111 321 112 322
rect 110 321 111 322
rect 109 321 110 322
rect 108 321 109 322
rect 107 321 108 322
rect 106 321 107 322
rect 105 321 106 322
rect 104 321 105 322
rect 103 321 104 322
rect 102 321 103 322
rect 101 321 102 322
rect 100 321 101 322
rect 99 321 100 322
rect 98 321 99 322
rect 97 321 98 322
rect 96 321 97 322
rect 77 321 78 322
rect 76 321 77 322
rect 75 321 76 322
rect 74 321 75 322
rect 73 321 74 322
rect 72 321 73 322
rect 71 321 72 322
rect 70 321 71 322
rect 69 321 70 322
rect 68 321 69 322
rect 67 321 68 322
rect 66 321 67 322
rect 65 321 66 322
rect 64 321 65 322
rect 63 321 64 322
rect 62 321 63 322
rect 61 321 62 322
rect 60 321 61 322
rect 59 321 60 322
rect 58 321 59 322
rect 57 321 58 322
rect 56 321 57 322
rect 55 321 56 322
rect 54 321 55 322
rect 53 321 54 322
rect 52 321 53 322
rect 51 321 52 322
rect 50 321 51 322
rect 49 321 50 322
rect 48 321 49 322
rect 47 321 48 322
rect 46 321 47 322
rect 34 321 35 322
rect 33 321 34 322
rect 32 321 33 322
rect 31 321 32 322
rect 30 321 31 322
rect 29 321 30 322
rect 28 321 29 322
rect 27 321 28 322
rect 26 321 27 322
rect 25 321 26 322
rect 24 321 25 322
rect 23 321 24 322
rect 22 321 23 322
rect 21 321 22 322
rect 20 321 21 322
rect 19 321 20 322
rect 18 321 19 322
rect 17 321 18 322
rect 478 322 479 323
rect 477 322 478 323
rect 476 322 477 323
rect 475 322 476 323
rect 474 322 475 323
rect 473 322 474 323
rect 472 322 473 323
rect 471 322 472 323
rect 470 322 471 323
rect 469 322 470 323
rect 468 322 469 323
rect 467 322 468 323
rect 466 322 467 323
rect 145 322 146 323
rect 144 322 145 323
rect 143 322 144 323
rect 142 322 143 323
rect 141 322 142 323
rect 140 322 141 323
rect 139 322 140 323
rect 138 322 139 323
rect 137 322 138 323
rect 136 322 137 323
rect 135 322 136 323
rect 134 322 135 323
rect 133 322 134 323
rect 132 322 133 323
rect 131 322 132 323
rect 130 322 131 323
rect 129 322 130 323
rect 128 322 129 323
rect 127 322 128 323
rect 126 322 127 323
rect 125 322 126 323
rect 124 322 125 323
rect 123 322 124 323
rect 122 322 123 323
rect 121 322 122 323
rect 120 322 121 323
rect 119 322 120 323
rect 118 322 119 323
rect 117 322 118 323
rect 116 322 117 323
rect 115 322 116 323
rect 114 322 115 323
rect 113 322 114 323
rect 112 322 113 323
rect 111 322 112 323
rect 110 322 111 323
rect 109 322 110 323
rect 108 322 109 323
rect 107 322 108 323
rect 106 322 107 323
rect 105 322 106 323
rect 104 322 105 323
rect 103 322 104 323
rect 102 322 103 323
rect 101 322 102 323
rect 100 322 101 323
rect 99 322 100 323
rect 98 322 99 323
rect 97 322 98 323
rect 78 322 79 323
rect 77 322 78 323
rect 76 322 77 323
rect 75 322 76 323
rect 74 322 75 323
rect 73 322 74 323
rect 72 322 73 323
rect 71 322 72 323
rect 70 322 71 323
rect 69 322 70 323
rect 68 322 69 323
rect 67 322 68 323
rect 66 322 67 323
rect 65 322 66 323
rect 64 322 65 323
rect 63 322 64 323
rect 62 322 63 323
rect 61 322 62 323
rect 60 322 61 323
rect 59 322 60 323
rect 58 322 59 323
rect 57 322 58 323
rect 56 322 57 323
rect 55 322 56 323
rect 54 322 55 323
rect 53 322 54 323
rect 52 322 53 323
rect 51 322 52 323
rect 50 322 51 323
rect 49 322 50 323
rect 48 322 49 323
rect 47 322 48 323
rect 46 322 47 323
rect 34 322 35 323
rect 33 322 34 323
rect 32 322 33 323
rect 31 322 32 323
rect 30 322 31 323
rect 29 322 30 323
rect 28 322 29 323
rect 27 322 28 323
rect 26 322 27 323
rect 25 322 26 323
rect 24 322 25 323
rect 23 322 24 323
rect 22 322 23 323
rect 21 322 22 323
rect 20 322 21 323
rect 19 322 20 323
rect 18 322 19 323
rect 478 323 479 324
rect 467 323 468 324
rect 466 323 467 324
rect 465 323 466 324
rect 464 323 465 324
rect 458 323 459 324
rect 147 323 148 324
rect 146 323 147 324
rect 145 323 146 324
rect 144 323 145 324
rect 143 323 144 324
rect 142 323 143 324
rect 141 323 142 324
rect 140 323 141 324
rect 139 323 140 324
rect 138 323 139 324
rect 137 323 138 324
rect 136 323 137 324
rect 135 323 136 324
rect 134 323 135 324
rect 133 323 134 324
rect 132 323 133 324
rect 131 323 132 324
rect 130 323 131 324
rect 129 323 130 324
rect 128 323 129 324
rect 127 323 128 324
rect 126 323 127 324
rect 125 323 126 324
rect 124 323 125 324
rect 123 323 124 324
rect 122 323 123 324
rect 121 323 122 324
rect 120 323 121 324
rect 119 323 120 324
rect 118 323 119 324
rect 117 323 118 324
rect 116 323 117 324
rect 115 323 116 324
rect 114 323 115 324
rect 113 323 114 324
rect 112 323 113 324
rect 111 323 112 324
rect 110 323 111 324
rect 109 323 110 324
rect 108 323 109 324
rect 107 323 108 324
rect 106 323 107 324
rect 105 323 106 324
rect 104 323 105 324
rect 103 323 104 324
rect 102 323 103 324
rect 101 323 102 324
rect 100 323 101 324
rect 99 323 100 324
rect 98 323 99 324
rect 78 323 79 324
rect 77 323 78 324
rect 76 323 77 324
rect 75 323 76 324
rect 74 323 75 324
rect 73 323 74 324
rect 72 323 73 324
rect 71 323 72 324
rect 70 323 71 324
rect 69 323 70 324
rect 68 323 69 324
rect 67 323 68 324
rect 66 323 67 324
rect 65 323 66 324
rect 64 323 65 324
rect 63 323 64 324
rect 62 323 63 324
rect 61 323 62 324
rect 60 323 61 324
rect 59 323 60 324
rect 58 323 59 324
rect 57 323 58 324
rect 56 323 57 324
rect 55 323 56 324
rect 54 323 55 324
rect 53 323 54 324
rect 52 323 53 324
rect 51 323 52 324
rect 50 323 51 324
rect 49 323 50 324
rect 48 323 49 324
rect 47 323 48 324
rect 35 323 36 324
rect 34 323 35 324
rect 33 323 34 324
rect 32 323 33 324
rect 31 323 32 324
rect 30 323 31 324
rect 29 323 30 324
rect 28 323 29 324
rect 27 323 28 324
rect 26 323 27 324
rect 25 323 26 324
rect 24 323 25 324
rect 23 323 24 324
rect 22 323 23 324
rect 21 323 22 324
rect 20 323 21 324
rect 19 323 20 324
rect 478 324 479 325
rect 465 324 466 325
rect 464 324 465 325
rect 463 324 464 325
rect 462 324 463 325
rect 458 324 459 325
rect 149 324 150 325
rect 148 324 149 325
rect 147 324 148 325
rect 146 324 147 325
rect 145 324 146 325
rect 144 324 145 325
rect 143 324 144 325
rect 142 324 143 325
rect 141 324 142 325
rect 140 324 141 325
rect 139 324 140 325
rect 138 324 139 325
rect 137 324 138 325
rect 136 324 137 325
rect 135 324 136 325
rect 134 324 135 325
rect 133 324 134 325
rect 132 324 133 325
rect 131 324 132 325
rect 130 324 131 325
rect 129 324 130 325
rect 128 324 129 325
rect 127 324 128 325
rect 126 324 127 325
rect 125 324 126 325
rect 124 324 125 325
rect 123 324 124 325
rect 122 324 123 325
rect 121 324 122 325
rect 120 324 121 325
rect 119 324 120 325
rect 118 324 119 325
rect 117 324 118 325
rect 116 324 117 325
rect 115 324 116 325
rect 114 324 115 325
rect 113 324 114 325
rect 112 324 113 325
rect 111 324 112 325
rect 110 324 111 325
rect 109 324 110 325
rect 108 324 109 325
rect 107 324 108 325
rect 106 324 107 325
rect 105 324 106 325
rect 104 324 105 325
rect 103 324 104 325
rect 102 324 103 325
rect 101 324 102 325
rect 100 324 101 325
rect 99 324 100 325
rect 98 324 99 325
rect 79 324 80 325
rect 78 324 79 325
rect 77 324 78 325
rect 76 324 77 325
rect 75 324 76 325
rect 74 324 75 325
rect 73 324 74 325
rect 72 324 73 325
rect 71 324 72 325
rect 70 324 71 325
rect 69 324 70 325
rect 68 324 69 325
rect 67 324 68 325
rect 66 324 67 325
rect 65 324 66 325
rect 64 324 65 325
rect 63 324 64 325
rect 62 324 63 325
rect 61 324 62 325
rect 60 324 61 325
rect 59 324 60 325
rect 58 324 59 325
rect 57 324 58 325
rect 56 324 57 325
rect 55 324 56 325
rect 54 324 55 325
rect 53 324 54 325
rect 52 324 53 325
rect 51 324 52 325
rect 50 324 51 325
rect 49 324 50 325
rect 48 324 49 325
rect 47 324 48 325
rect 35 324 36 325
rect 34 324 35 325
rect 33 324 34 325
rect 32 324 33 325
rect 31 324 32 325
rect 30 324 31 325
rect 29 324 30 325
rect 28 324 29 325
rect 27 324 28 325
rect 26 324 27 325
rect 25 324 26 325
rect 24 324 25 325
rect 23 324 24 325
rect 22 324 23 325
rect 21 324 22 325
rect 20 324 21 325
rect 478 325 479 326
rect 463 325 464 326
rect 462 325 463 326
rect 461 325 462 326
rect 460 325 461 326
rect 459 325 460 326
rect 458 325 459 326
rect 151 325 152 326
rect 150 325 151 326
rect 149 325 150 326
rect 148 325 149 326
rect 147 325 148 326
rect 146 325 147 326
rect 145 325 146 326
rect 144 325 145 326
rect 143 325 144 326
rect 142 325 143 326
rect 141 325 142 326
rect 140 325 141 326
rect 139 325 140 326
rect 138 325 139 326
rect 137 325 138 326
rect 136 325 137 326
rect 135 325 136 326
rect 134 325 135 326
rect 133 325 134 326
rect 132 325 133 326
rect 131 325 132 326
rect 130 325 131 326
rect 129 325 130 326
rect 128 325 129 326
rect 127 325 128 326
rect 126 325 127 326
rect 125 325 126 326
rect 124 325 125 326
rect 123 325 124 326
rect 122 325 123 326
rect 121 325 122 326
rect 120 325 121 326
rect 119 325 120 326
rect 118 325 119 326
rect 117 325 118 326
rect 116 325 117 326
rect 115 325 116 326
rect 114 325 115 326
rect 113 325 114 326
rect 112 325 113 326
rect 111 325 112 326
rect 110 325 111 326
rect 109 325 110 326
rect 108 325 109 326
rect 107 325 108 326
rect 106 325 107 326
rect 105 325 106 326
rect 104 325 105 326
rect 103 325 104 326
rect 102 325 103 326
rect 101 325 102 326
rect 100 325 101 326
rect 99 325 100 326
rect 80 325 81 326
rect 79 325 80 326
rect 78 325 79 326
rect 77 325 78 326
rect 76 325 77 326
rect 75 325 76 326
rect 74 325 75 326
rect 73 325 74 326
rect 72 325 73 326
rect 71 325 72 326
rect 70 325 71 326
rect 69 325 70 326
rect 68 325 69 326
rect 67 325 68 326
rect 66 325 67 326
rect 65 325 66 326
rect 64 325 65 326
rect 63 325 64 326
rect 62 325 63 326
rect 61 325 62 326
rect 60 325 61 326
rect 59 325 60 326
rect 58 325 59 326
rect 57 325 58 326
rect 56 325 57 326
rect 55 325 56 326
rect 54 325 55 326
rect 53 325 54 326
rect 52 325 53 326
rect 51 325 52 326
rect 50 325 51 326
rect 49 325 50 326
rect 48 325 49 326
rect 35 325 36 326
rect 34 325 35 326
rect 33 325 34 326
rect 32 325 33 326
rect 31 325 32 326
rect 30 325 31 326
rect 29 325 30 326
rect 28 325 29 326
rect 27 325 28 326
rect 26 325 27 326
rect 25 325 26 326
rect 24 325 25 326
rect 23 325 24 326
rect 22 325 23 326
rect 21 325 22 326
rect 20 325 21 326
rect 461 326 462 327
rect 460 326 461 327
rect 459 326 460 327
rect 458 326 459 327
rect 154 326 155 327
rect 153 326 154 327
rect 152 326 153 327
rect 151 326 152 327
rect 150 326 151 327
rect 149 326 150 327
rect 148 326 149 327
rect 147 326 148 327
rect 146 326 147 327
rect 145 326 146 327
rect 144 326 145 327
rect 143 326 144 327
rect 142 326 143 327
rect 141 326 142 327
rect 140 326 141 327
rect 139 326 140 327
rect 138 326 139 327
rect 137 326 138 327
rect 136 326 137 327
rect 135 326 136 327
rect 134 326 135 327
rect 133 326 134 327
rect 132 326 133 327
rect 131 326 132 327
rect 130 326 131 327
rect 129 326 130 327
rect 128 326 129 327
rect 127 326 128 327
rect 126 326 127 327
rect 125 326 126 327
rect 124 326 125 327
rect 123 326 124 327
rect 122 326 123 327
rect 121 326 122 327
rect 120 326 121 327
rect 119 326 120 327
rect 118 326 119 327
rect 117 326 118 327
rect 116 326 117 327
rect 115 326 116 327
rect 114 326 115 327
rect 113 326 114 327
rect 112 326 113 327
rect 111 326 112 327
rect 110 326 111 327
rect 109 326 110 327
rect 108 326 109 327
rect 107 326 108 327
rect 106 326 107 327
rect 105 326 106 327
rect 104 326 105 327
rect 103 326 104 327
rect 102 326 103 327
rect 101 326 102 327
rect 100 326 101 327
rect 80 326 81 327
rect 79 326 80 327
rect 78 326 79 327
rect 77 326 78 327
rect 76 326 77 327
rect 75 326 76 327
rect 74 326 75 327
rect 73 326 74 327
rect 72 326 73 327
rect 71 326 72 327
rect 70 326 71 327
rect 69 326 70 327
rect 68 326 69 327
rect 67 326 68 327
rect 66 326 67 327
rect 65 326 66 327
rect 64 326 65 327
rect 63 326 64 327
rect 62 326 63 327
rect 61 326 62 327
rect 60 326 61 327
rect 59 326 60 327
rect 58 326 59 327
rect 57 326 58 327
rect 56 326 57 327
rect 55 326 56 327
rect 54 326 55 327
rect 53 326 54 327
rect 52 326 53 327
rect 51 326 52 327
rect 50 326 51 327
rect 49 326 50 327
rect 48 326 49 327
rect 36 326 37 327
rect 35 326 36 327
rect 34 326 35 327
rect 33 326 34 327
rect 32 326 33 327
rect 31 326 32 327
rect 30 326 31 327
rect 29 326 30 327
rect 28 326 29 327
rect 27 326 28 327
rect 26 326 27 327
rect 25 326 26 327
rect 24 326 25 327
rect 23 326 24 327
rect 22 326 23 327
rect 21 326 22 327
rect 460 327 461 328
rect 459 327 460 328
rect 458 327 459 328
rect 156 327 157 328
rect 155 327 156 328
rect 154 327 155 328
rect 153 327 154 328
rect 152 327 153 328
rect 151 327 152 328
rect 150 327 151 328
rect 149 327 150 328
rect 148 327 149 328
rect 147 327 148 328
rect 146 327 147 328
rect 145 327 146 328
rect 144 327 145 328
rect 143 327 144 328
rect 142 327 143 328
rect 141 327 142 328
rect 140 327 141 328
rect 139 327 140 328
rect 138 327 139 328
rect 137 327 138 328
rect 136 327 137 328
rect 135 327 136 328
rect 134 327 135 328
rect 133 327 134 328
rect 132 327 133 328
rect 131 327 132 328
rect 130 327 131 328
rect 129 327 130 328
rect 128 327 129 328
rect 127 327 128 328
rect 126 327 127 328
rect 125 327 126 328
rect 124 327 125 328
rect 123 327 124 328
rect 122 327 123 328
rect 121 327 122 328
rect 120 327 121 328
rect 119 327 120 328
rect 118 327 119 328
rect 117 327 118 328
rect 116 327 117 328
rect 115 327 116 328
rect 114 327 115 328
rect 113 327 114 328
rect 112 327 113 328
rect 111 327 112 328
rect 110 327 111 328
rect 109 327 110 328
rect 108 327 109 328
rect 107 327 108 328
rect 106 327 107 328
rect 105 327 106 328
rect 104 327 105 328
rect 103 327 104 328
rect 102 327 103 328
rect 101 327 102 328
rect 81 327 82 328
rect 80 327 81 328
rect 79 327 80 328
rect 78 327 79 328
rect 77 327 78 328
rect 76 327 77 328
rect 75 327 76 328
rect 74 327 75 328
rect 73 327 74 328
rect 72 327 73 328
rect 71 327 72 328
rect 70 327 71 328
rect 69 327 70 328
rect 68 327 69 328
rect 67 327 68 328
rect 66 327 67 328
rect 65 327 66 328
rect 64 327 65 328
rect 63 327 64 328
rect 62 327 63 328
rect 61 327 62 328
rect 60 327 61 328
rect 59 327 60 328
rect 58 327 59 328
rect 57 327 58 328
rect 56 327 57 328
rect 55 327 56 328
rect 54 327 55 328
rect 53 327 54 328
rect 52 327 53 328
rect 51 327 52 328
rect 50 327 51 328
rect 49 327 50 328
rect 48 327 49 328
rect 36 327 37 328
rect 35 327 36 328
rect 34 327 35 328
rect 33 327 34 328
rect 32 327 33 328
rect 31 327 32 328
rect 30 327 31 328
rect 29 327 30 328
rect 28 327 29 328
rect 27 327 28 328
rect 26 327 27 328
rect 25 327 26 328
rect 24 327 25 328
rect 23 327 24 328
rect 22 327 23 328
rect 459 328 460 329
rect 458 328 459 329
rect 159 328 160 329
rect 158 328 159 329
rect 157 328 158 329
rect 156 328 157 329
rect 155 328 156 329
rect 154 328 155 329
rect 153 328 154 329
rect 152 328 153 329
rect 151 328 152 329
rect 150 328 151 329
rect 149 328 150 329
rect 148 328 149 329
rect 147 328 148 329
rect 146 328 147 329
rect 145 328 146 329
rect 144 328 145 329
rect 143 328 144 329
rect 142 328 143 329
rect 141 328 142 329
rect 140 328 141 329
rect 139 328 140 329
rect 138 328 139 329
rect 137 328 138 329
rect 136 328 137 329
rect 135 328 136 329
rect 134 328 135 329
rect 133 328 134 329
rect 132 328 133 329
rect 131 328 132 329
rect 130 328 131 329
rect 129 328 130 329
rect 128 328 129 329
rect 127 328 128 329
rect 126 328 127 329
rect 125 328 126 329
rect 124 328 125 329
rect 123 328 124 329
rect 122 328 123 329
rect 121 328 122 329
rect 120 328 121 329
rect 119 328 120 329
rect 118 328 119 329
rect 117 328 118 329
rect 116 328 117 329
rect 115 328 116 329
rect 114 328 115 329
rect 113 328 114 329
rect 112 328 113 329
rect 111 328 112 329
rect 110 328 111 329
rect 109 328 110 329
rect 108 328 109 329
rect 107 328 108 329
rect 106 328 107 329
rect 105 328 106 329
rect 104 328 105 329
rect 103 328 104 329
rect 102 328 103 329
rect 82 328 83 329
rect 81 328 82 329
rect 80 328 81 329
rect 79 328 80 329
rect 78 328 79 329
rect 77 328 78 329
rect 76 328 77 329
rect 75 328 76 329
rect 74 328 75 329
rect 73 328 74 329
rect 72 328 73 329
rect 71 328 72 329
rect 70 328 71 329
rect 69 328 70 329
rect 68 328 69 329
rect 67 328 68 329
rect 66 328 67 329
rect 65 328 66 329
rect 64 328 65 329
rect 63 328 64 329
rect 62 328 63 329
rect 61 328 62 329
rect 60 328 61 329
rect 59 328 60 329
rect 58 328 59 329
rect 57 328 58 329
rect 56 328 57 329
rect 55 328 56 329
rect 54 328 55 329
rect 53 328 54 329
rect 52 328 53 329
rect 51 328 52 329
rect 50 328 51 329
rect 49 328 50 329
rect 37 328 38 329
rect 36 328 37 329
rect 35 328 36 329
rect 34 328 35 329
rect 33 328 34 329
rect 32 328 33 329
rect 31 328 32 329
rect 30 328 31 329
rect 29 328 30 329
rect 28 328 29 329
rect 27 328 28 329
rect 26 328 27 329
rect 25 328 26 329
rect 24 328 25 329
rect 23 328 24 329
rect 458 329 459 330
rect 437 329 438 330
rect 436 329 437 330
rect 435 329 436 330
rect 162 329 163 330
rect 161 329 162 330
rect 160 329 161 330
rect 159 329 160 330
rect 158 329 159 330
rect 157 329 158 330
rect 156 329 157 330
rect 155 329 156 330
rect 154 329 155 330
rect 153 329 154 330
rect 152 329 153 330
rect 151 329 152 330
rect 150 329 151 330
rect 149 329 150 330
rect 148 329 149 330
rect 147 329 148 330
rect 146 329 147 330
rect 145 329 146 330
rect 144 329 145 330
rect 143 329 144 330
rect 142 329 143 330
rect 141 329 142 330
rect 140 329 141 330
rect 139 329 140 330
rect 138 329 139 330
rect 137 329 138 330
rect 136 329 137 330
rect 135 329 136 330
rect 134 329 135 330
rect 133 329 134 330
rect 132 329 133 330
rect 131 329 132 330
rect 130 329 131 330
rect 129 329 130 330
rect 128 329 129 330
rect 127 329 128 330
rect 126 329 127 330
rect 125 329 126 330
rect 124 329 125 330
rect 123 329 124 330
rect 122 329 123 330
rect 121 329 122 330
rect 120 329 121 330
rect 119 329 120 330
rect 118 329 119 330
rect 117 329 118 330
rect 116 329 117 330
rect 115 329 116 330
rect 114 329 115 330
rect 113 329 114 330
rect 112 329 113 330
rect 111 329 112 330
rect 110 329 111 330
rect 109 329 110 330
rect 108 329 109 330
rect 107 329 108 330
rect 106 329 107 330
rect 105 329 106 330
rect 104 329 105 330
rect 103 329 104 330
rect 102 329 103 330
rect 82 329 83 330
rect 81 329 82 330
rect 80 329 81 330
rect 79 329 80 330
rect 78 329 79 330
rect 77 329 78 330
rect 76 329 77 330
rect 75 329 76 330
rect 74 329 75 330
rect 73 329 74 330
rect 72 329 73 330
rect 71 329 72 330
rect 70 329 71 330
rect 69 329 70 330
rect 68 329 69 330
rect 67 329 68 330
rect 66 329 67 330
rect 65 329 66 330
rect 64 329 65 330
rect 63 329 64 330
rect 62 329 63 330
rect 61 329 62 330
rect 60 329 61 330
rect 59 329 60 330
rect 58 329 59 330
rect 57 329 58 330
rect 56 329 57 330
rect 55 329 56 330
rect 54 329 55 330
rect 53 329 54 330
rect 52 329 53 330
rect 51 329 52 330
rect 50 329 51 330
rect 49 329 50 330
rect 37 329 38 330
rect 36 329 37 330
rect 35 329 36 330
rect 34 329 35 330
rect 33 329 34 330
rect 32 329 33 330
rect 31 329 32 330
rect 30 329 31 330
rect 29 329 30 330
rect 28 329 29 330
rect 27 329 28 330
rect 26 329 27 330
rect 25 329 26 330
rect 24 329 25 330
rect 458 330 459 331
rect 437 330 438 331
rect 436 330 437 331
rect 435 330 436 331
rect 395 330 396 331
rect 394 330 395 331
rect 393 330 394 331
rect 165 330 166 331
rect 164 330 165 331
rect 163 330 164 331
rect 162 330 163 331
rect 161 330 162 331
rect 160 330 161 331
rect 159 330 160 331
rect 158 330 159 331
rect 157 330 158 331
rect 156 330 157 331
rect 155 330 156 331
rect 154 330 155 331
rect 153 330 154 331
rect 152 330 153 331
rect 151 330 152 331
rect 150 330 151 331
rect 149 330 150 331
rect 148 330 149 331
rect 147 330 148 331
rect 146 330 147 331
rect 145 330 146 331
rect 144 330 145 331
rect 143 330 144 331
rect 142 330 143 331
rect 141 330 142 331
rect 140 330 141 331
rect 139 330 140 331
rect 138 330 139 331
rect 137 330 138 331
rect 136 330 137 331
rect 135 330 136 331
rect 134 330 135 331
rect 133 330 134 331
rect 132 330 133 331
rect 131 330 132 331
rect 130 330 131 331
rect 129 330 130 331
rect 128 330 129 331
rect 127 330 128 331
rect 126 330 127 331
rect 125 330 126 331
rect 124 330 125 331
rect 123 330 124 331
rect 122 330 123 331
rect 121 330 122 331
rect 120 330 121 331
rect 119 330 120 331
rect 118 330 119 331
rect 117 330 118 331
rect 116 330 117 331
rect 115 330 116 331
rect 114 330 115 331
rect 113 330 114 331
rect 112 330 113 331
rect 111 330 112 331
rect 110 330 111 331
rect 109 330 110 331
rect 108 330 109 331
rect 107 330 108 331
rect 106 330 107 331
rect 105 330 106 331
rect 104 330 105 331
rect 103 330 104 331
rect 83 330 84 331
rect 82 330 83 331
rect 81 330 82 331
rect 80 330 81 331
rect 79 330 80 331
rect 78 330 79 331
rect 77 330 78 331
rect 76 330 77 331
rect 75 330 76 331
rect 74 330 75 331
rect 73 330 74 331
rect 72 330 73 331
rect 71 330 72 331
rect 70 330 71 331
rect 69 330 70 331
rect 68 330 69 331
rect 67 330 68 331
rect 66 330 67 331
rect 65 330 66 331
rect 64 330 65 331
rect 63 330 64 331
rect 62 330 63 331
rect 61 330 62 331
rect 60 330 61 331
rect 59 330 60 331
rect 58 330 59 331
rect 57 330 58 331
rect 56 330 57 331
rect 55 330 56 331
rect 54 330 55 331
rect 53 330 54 331
rect 52 330 53 331
rect 51 330 52 331
rect 50 330 51 331
rect 49 330 50 331
rect 37 330 38 331
rect 36 330 37 331
rect 35 330 36 331
rect 34 330 35 331
rect 33 330 34 331
rect 32 330 33 331
rect 31 330 32 331
rect 30 330 31 331
rect 29 330 30 331
rect 28 330 29 331
rect 27 330 28 331
rect 26 330 27 331
rect 25 330 26 331
rect 437 331 438 332
rect 436 331 437 332
rect 435 331 436 332
rect 395 331 396 332
rect 394 331 395 332
rect 393 331 394 332
rect 168 331 169 332
rect 167 331 168 332
rect 166 331 167 332
rect 165 331 166 332
rect 164 331 165 332
rect 163 331 164 332
rect 162 331 163 332
rect 161 331 162 332
rect 160 331 161 332
rect 159 331 160 332
rect 158 331 159 332
rect 157 331 158 332
rect 156 331 157 332
rect 155 331 156 332
rect 154 331 155 332
rect 153 331 154 332
rect 152 331 153 332
rect 151 331 152 332
rect 150 331 151 332
rect 149 331 150 332
rect 148 331 149 332
rect 147 331 148 332
rect 146 331 147 332
rect 145 331 146 332
rect 144 331 145 332
rect 143 331 144 332
rect 142 331 143 332
rect 141 331 142 332
rect 140 331 141 332
rect 139 331 140 332
rect 138 331 139 332
rect 137 331 138 332
rect 136 331 137 332
rect 135 331 136 332
rect 134 331 135 332
rect 133 331 134 332
rect 132 331 133 332
rect 131 331 132 332
rect 130 331 131 332
rect 129 331 130 332
rect 128 331 129 332
rect 127 331 128 332
rect 126 331 127 332
rect 125 331 126 332
rect 124 331 125 332
rect 123 331 124 332
rect 122 331 123 332
rect 121 331 122 332
rect 120 331 121 332
rect 119 331 120 332
rect 118 331 119 332
rect 117 331 118 332
rect 116 331 117 332
rect 115 331 116 332
rect 114 331 115 332
rect 113 331 114 332
rect 112 331 113 332
rect 111 331 112 332
rect 110 331 111 332
rect 109 331 110 332
rect 108 331 109 332
rect 107 331 108 332
rect 106 331 107 332
rect 105 331 106 332
rect 104 331 105 332
rect 84 331 85 332
rect 83 331 84 332
rect 82 331 83 332
rect 81 331 82 332
rect 80 331 81 332
rect 79 331 80 332
rect 78 331 79 332
rect 77 331 78 332
rect 76 331 77 332
rect 75 331 76 332
rect 74 331 75 332
rect 73 331 74 332
rect 72 331 73 332
rect 71 331 72 332
rect 70 331 71 332
rect 69 331 70 332
rect 68 331 69 332
rect 67 331 68 332
rect 66 331 67 332
rect 65 331 66 332
rect 64 331 65 332
rect 63 331 64 332
rect 62 331 63 332
rect 61 331 62 332
rect 60 331 61 332
rect 59 331 60 332
rect 58 331 59 332
rect 57 331 58 332
rect 56 331 57 332
rect 55 331 56 332
rect 54 331 55 332
rect 53 331 54 332
rect 52 331 53 332
rect 51 331 52 332
rect 50 331 51 332
rect 38 331 39 332
rect 37 331 38 332
rect 36 331 37 332
rect 35 331 36 332
rect 34 331 35 332
rect 33 331 34 332
rect 32 331 33 332
rect 31 331 32 332
rect 30 331 31 332
rect 29 331 30 332
rect 28 331 29 332
rect 27 331 28 332
rect 26 331 27 332
rect 437 332 438 333
rect 436 332 437 333
rect 435 332 436 333
rect 395 332 396 333
rect 394 332 395 333
rect 393 332 394 333
rect 172 332 173 333
rect 171 332 172 333
rect 170 332 171 333
rect 169 332 170 333
rect 168 332 169 333
rect 167 332 168 333
rect 166 332 167 333
rect 165 332 166 333
rect 164 332 165 333
rect 163 332 164 333
rect 162 332 163 333
rect 161 332 162 333
rect 160 332 161 333
rect 159 332 160 333
rect 158 332 159 333
rect 157 332 158 333
rect 156 332 157 333
rect 155 332 156 333
rect 154 332 155 333
rect 153 332 154 333
rect 152 332 153 333
rect 151 332 152 333
rect 150 332 151 333
rect 149 332 150 333
rect 148 332 149 333
rect 147 332 148 333
rect 146 332 147 333
rect 145 332 146 333
rect 144 332 145 333
rect 143 332 144 333
rect 142 332 143 333
rect 141 332 142 333
rect 140 332 141 333
rect 139 332 140 333
rect 138 332 139 333
rect 137 332 138 333
rect 136 332 137 333
rect 135 332 136 333
rect 134 332 135 333
rect 133 332 134 333
rect 132 332 133 333
rect 131 332 132 333
rect 130 332 131 333
rect 129 332 130 333
rect 128 332 129 333
rect 127 332 128 333
rect 126 332 127 333
rect 125 332 126 333
rect 124 332 125 333
rect 123 332 124 333
rect 122 332 123 333
rect 121 332 122 333
rect 120 332 121 333
rect 119 332 120 333
rect 118 332 119 333
rect 117 332 118 333
rect 116 332 117 333
rect 115 332 116 333
rect 114 332 115 333
rect 113 332 114 333
rect 112 332 113 333
rect 111 332 112 333
rect 110 332 111 333
rect 109 332 110 333
rect 108 332 109 333
rect 107 332 108 333
rect 106 332 107 333
rect 105 332 106 333
rect 85 332 86 333
rect 84 332 85 333
rect 83 332 84 333
rect 82 332 83 333
rect 81 332 82 333
rect 80 332 81 333
rect 79 332 80 333
rect 78 332 79 333
rect 77 332 78 333
rect 76 332 77 333
rect 75 332 76 333
rect 74 332 75 333
rect 73 332 74 333
rect 72 332 73 333
rect 71 332 72 333
rect 70 332 71 333
rect 69 332 70 333
rect 68 332 69 333
rect 67 332 68 333
rect 66 332 67 333
rect 65 332 66 333
rect 64 332 65 333
rect 63 332 64 333
rect 62 332 63 333
rect 61 332 62 333
rect 60 332 61 333
rect 59 332 60 333
rect 58 332 59 333
rect 57 332 58 333
rect 56 332 57 333
rect 55 332 56 333
rect 54 332 55 333
rect 53 332 54 333
rect 52 332 53 333
rect 51 332 52 333
rect 50 332 51 333
rect 38 332 39 333
rect 37 332 38 333
rect 36 332 37 333
rect 35 332 36 333
rect 34 332 35 333
rect 33 332 34 333
rect 32 332 33 333
rect 31 332 32 333
rect 30 332 31 333
rect 29 332 30 333
rect 28 332 29 333
rect 27 332 28 333
rect 437 333 438 334
rect 436 333 437 334
rect 435 333 436 334
rect 395 333 396 334
rect 394 333 395 334
rect 393 333 394 334
rect 176 333 177 334
rect 175 333 176 334
rect 174 333 175 334
rect 173 333 174 334
rect 172 333 173 334
rect 171 333 172 334
rect 170 333 171 334
rect 169 333 170 334
rect 168 333 169 334
rect 167 333 168 334
rect 166 333 167 334
rect 165 333 166 334
rect 164 333 165 334
rect 163 333 164 334
rect 162 333 163 334
rect 161 333 162 334
rect 160 333 161 334
rect 159 333 160 334
rect 158 333 159 334
rect 157 333 158 334
rect 156 333 157 334
rect 155 333 156 334
rect 154 333 155 334
rect 153 333 154 334
rect 152 333 153 334
rect 151 333 152 334
rect 150 333 151 334
rect 149 333 150 334
rect 148 333 149 334
rect 147 333 148 334
rect 146 333 147 334
rect 145 333 146 334
rect 144 333 145 334
rect 143 333 144 334
rect 142 333 143 334
rect 141 333 142 334
rect 140 333 141 334
rect 139 333 140 334
rect 138 333 139 334
rect 137 333 138 334
rect 136 333 137 334
rect 135 333 136 334
rect 134 333 135 334
rect 133 333 134 334
rect 132 333 133 334
rect 131 333 132 334
rect 130 333 131 334
rect 129 333 130 334
rect 128 333 129 334
rect 127 333 128 334
rect 126 333 127 334
rect 125 333 126 334
rect 124 333 125 334
rect 123 333 124 334
rect 122 333 123 334
rect 121 333 122 334
rect 120 333 121 334
rect 119 333 120 334
rect 118 333 119 334
rect 117 333 118 334
rect 116 333 117 334
rect 115 333 116 334
rect 114 333 115 334
rect 113 333 114 334
rect 112 333 113 334
rect 111 333 112 334
rect 110 333 111 334
rect 109 333 110 334
rect 108 333 109 334
rect 107 333 108 334
rect 106 333 107 334
rect 85 333 86 334
rect 84 333 85 334
rect 83 333 84 334
rect 82 333 83 334
rect 81 333 82 334
rect 80 333 81 334
rect 79 333 80 334
rect 78 333 79 334
rect 77 333 78 334
rect 76 333 77 334
rect 75 333 76 334
rect 74 333 75 334
rect 73 333 74 334
rect 72 333 73 334
rect 71 333 72 334
rect 70 333 71 334
rect 69 333 70 334
rect 68 333 69 334
rect 67 333 68 334
rect 66 333 67 334
rect 65 333 66 334
rect 64 333 65 334
rect 63 333 64 334
rect 62 333 63 334
rect 61 333 62 334
rect 60 333 61 334
rect 59 333 60 334
rect 58 333 59 334
rect 57 333 58 334
rect 56 333 57 334
rect 55 333 56 334
rect 54 333 55 334
rect 53 333 54 334
rect 52 333 53 334
rect 51 333 52 334
rect 38 333 39 334
rect 37 333 38 334
rect 36 333 37 334
rect 35 333 36 334
rect 34 333 35 334
rect 33 333 34 334
rect 32 333 33 334
rect 31 333 32 334
rect 30 333 31 334
rect 29 333 30 334
rect 28 333 29 334
rect 437 334 438 335
rect 436 334 437 335
rect 435 334 436 335
rect 434 334 435 335
rect 396 334 397 335
rect 395 334 396 335
rect 394 334 395 335
rect 393 334 394 335
rect 175 334 176 335
rect 174 334 175 335
rect 173 334 174 335
rect 172 334 173 335
rect 171 334 172 335
rect 170 334 171 335
rect 169 334 170 335
rect 168 334 169 335
rect 167 334 168 335
rect 166 334 167 335
rect 165 334 166 335
rect 164 334 165 335
rect 163 334 164 335
rect 162 334 163 335
rect 161 334 162 335
rect 160 334 161 335
rect 159 334 160 335
rect 158 334 159 335
rect 157 334 158 335
rect 156 334 157 335
rect 155 334 156 335
rect 154 334 155 335
rect 153 334 154 335
rect 152 334 153 335
rect 151 334 152 335
rect 150 334 151 335
rect 149 334 150 335
rect 148 334 149 335
rect 147 334 148 335
rect 146 334 147 335
rect 145 334 146 335
rect 144 334 145 335
rect 143 334 144 335
rect 142 334 143 335
rect 141 334 142 335
rect 140 334 141 335
rect 139 334 140 335
rect 138 334 139 335
rect 137 334 138 335
rect 136 334 137 335
rect 135 334 136 335
rect 134 334 135 335
rect 133 334 134 335
rect 132 334 133 335
rect 131 334 132 335
rect 130 334 131 335
rect 129 334 130 335
rect 128 334 129 335
rect 127 334 128 335
rect 126 334 127 335
rect 125 334 126 335
rect 124 334 125 335
rect 123 334 124 335
rect 122 334 123 335
rect 121 334 122 335
rect 120 334 121 335
rect 119 334 120 335
rect 118 334 119 335
rect 117 334 118 335
rect 116 334 117 335
rect 115 334 116 335
rect 114 334 115 335
rect 113 334 114 335
rect 112 334 113 335
rect 111 334 112 335
rect 110 334 111 335
rect 109 334 110 335
rect 108 334 109 335
rect 107 334 108 335
rect 86 334 87 335
rect 85 334 86 335
rect 84 334 85 335
rect 83 334 84 335
rect 82 334 83 335
rect 81 334 82 335
rect 80 334 81 335
rect 79 334 80 335
rect 78 334 79 335
rect 77 334 78 335
rect 76 334 77 335
rect 75 334 76 335
rect 74 334 75 335
rect 73 334 74 335
rect 72 334 73 335
rect 71 334 72 335
rect 70 334 71 335
rect 69 334 70 335
rect 68 334 69 335
rect 67 334 68 335
rect 66 334 67 335
rect 65 334 66 335
rect 64 334 65 335
rect 63 334 64 335
rect 62 334 63 335
rect 61 334 62 335
rect 60 334 61 335
rect 59 334 60 335
rect 58 334 59 335
rect 57 334 58 335
rect 56 334 57 335
rect 55 334 56 335
rect 54 334 55 335
rect 53 334 54 335
rect 52 334 53 335
rect 51 334 52 335
rect 39 334 40 335
rect 38 334 39 335
rect 37 334 38 335
rect 36 334 37 335
rect 35 334 36 335
rect 34 334 35 335
rect 33 334 34 335
rect 32 334 33 335
rect 31 334 32 335
rect 30 334 31 335
rect 29 334 30 335
rect 437 335 438 336
rect 436 335 437 336
rect 435 335 436 336
rect 434 335 435 336
rect 433 335 434 336
rect 432 335 433 336
rect 431 335 432 336
rect 430 335 431 336
rect 429 335 430 336
rect 428 335 429 336
rect 427 335 428 336
rect 426 335 427 336
rect 425 335 426 336
rect 424 335 425 336
rect 423 335 424 336
rect 422 335 423 336
rect 421 335 422 336
rect 420 335 421 336
rect 419 335 420 336
rect 418 335 419 336
rect 417 335 418 336
rect 416 335 417 336
rect 415 335 416 336
rect 414 335 415 336
rect 413 335 414 336
rect 412 335 413 336
rect 411 335 412 336
rect 410 335 411 336
rect 409 335 410 336
rect 408 335 409 336
rect 407 335 408 336
rect 406 335 407 336
rect 405 335 406 336
rect 404 335 405 336
rect 403 335 404 336
rect 402 335 403 336
rect 401 335 402 336
rect 400 335 401 336
rect 399 335 400 336
rect 398 335 399 336
rect 397 335 398 336
rect 396 335 397 336
rect 395 335 396 336
rect 394 335 395 336
rect 393 335 394 336
rect 174 335 175 336
rect 173 335 174 336
rect 172 335 173 336
rect 171 335 172 336
rect 170 335 171 336
rect 169 335 170 336
rect 168 335 169 336
rect 167 335 168 336
rect 166 335 167 336
rect 165 335 166 336
rect 164 335 165 336
rect 163 335 164 336
rect 162 335 163 336
rect 161 335 162 336
rect 160 335 161 336
rect 159 335 160 336
rect 158 335 159 336
rect 157 335 158 336
rect 156 335 157 336
rect 155 335 156 336
rect 154 335 155 336
rect 153 335 154 336
rect 152 335 153 336
rect 151 335 152 336
rect 150 335 151 336
rect 149 335 150 336
rect 148 335 149 336
rect 147 335 148 336
rect 146 335 147 336
rect 145 335 146 336
rect 144 335 145 336
rect 143 335 144 336
rect 142 335 143 336
rect 141 335 142 336
rect 140 335 141 336
rect 139 335 140 336
rect 138 335 139 336
rect 137 335 138 336
rect 136 335 137 336
rect 135 335 136 336
rect 134 335 135 336
rect 133 335 134 336
rect 132 335 133 336
rect 131 335 132 336
rect 130 335 131 336
rect 129 335 130 336
rect 128 335 129 336
rect 127 335 128 336
rect 126 335 127 336
rect 125 335 126 336
rect 124 335 125 336
rect 123 335 124 336
rect 122 335 123 336
rect 121 335 122 336
rect 120 335 121 336
rect 119 335 120 336
rect 118 335 119 336
rect 117 335 118 336
rect 116 335 117 336
rect 115 335 116 336
rect 114 335 115 336
rect 113 335 114 336
rect 112 335 113 336
rect 111 335 112 336
rect 110 335 111 336
rect 109 335 110 336
rect 108 335 109 336
rect 87 335 88 336
rect 86 335 87 336
rect 85 335 86 336
rect 84 335 85 336
rect 83 335 84 336
rect 82 335 83 336
rect 81 335 82 336
rect 80 335 81 336
rect 79 335 80 336
rect 78 335 79 336
rect 77 335 78 336
rect 76 335 77 336
rect 75 335 76 336
rect 74 335 75 336
rect 73 335 74 336
rect 72 335 73 336
rect 71 335 72 336
rect 70 335 71 336
rect 69 335 70 336
rect 68 335 69 336
rect 67 335 68 336
rect 66 335 67 336
rect 65 335 66 336
rect 64 335 65 336
rect 63 335 64 336
rect 62 335 63 336
rect 61 335 62 336
rect 60 335 61 336
rect 59 335 60 336
rect 58 335 59 336
rect 57 335 58 336
rect 56 335 57 336
rect 55 335 56 336
rect 54 335 55 336
rect 53 335 54 336
rect 52 335 53 336
rect 51 335 52 336
rect 39 335 40 336
rect 38 335 39 336
rect 37 335 38 336
rect 36 335 37 336
rect 35 335 36 336
rect 34 335 35 336
rect 33 335 34 336
rect 32 335 33 336
rect 31 335 32 336
rect 30 335 31 336
rect 437 336 438 337
rect 436 336 437 337
rect 435 336 436 337
rect 434 336 435 337
rect 433 336 434 337
rect 432 336 433 337
rect 431 336 432 337
rect 430 336 431 337
rect 429 336 430 337
rect 428 336 429 337
rect 427 336 428 337
rect 426 336 427 337
rect 425 336 426 337
rect 424 336 425 337
rect 423 336 424 337
rect 422 336 423 337
rect 421 336 422 337
rect 420 336 421 337
rect 419 336 420 337
rect 418 336 419 337
rect 417 336 418 337
rect 416 336 417 337
rect 415 336 416 337
rect 414 336 415 337
rect 413 336 414 337
rect 412 336 413 337
rect 411 336 412 337
rect 410 336 411 337
rect 409 336 410 337
rect 408 336 409 337
rect 407 336 408 337
rect 406 336 407 337
rect 405 336 406 337
rect 404 336 405 337
rect 403 336 404 337
rect 402 336 403 337
rect 401 336 402 337
rect 400 336 401 337
rect 399 336 400 337
rect 398 336 399 337
rect 397 336 398 337
rect 396 336 397 337
rect 395 336 396 337
rect 394 336 395 337
rect 393 336 394 337
rect 173 336 174 337
rect 172 336 173 337
rect 171 336 172 337
rect 170 336 171 337
rect 169 336 170 337
rect 168 336 169 337
rect 167 336 168 337
rect 166 336 167 337
rect 165 336 166 337
rect 164 336 165 337
rect 163 336 164 337
rect 162 336 163 337
rect 161 336 162 337
rect 160 336 161 337
rect 159 336 160 337
rect 158 336 159 337
rect 157 336 158 337
rect 156 336 157 337
rect 155 336 156 337
rect 154 336 155 337
rect 153 336 154 337
rect 152 336 153 337
rect 151 336 152 337
rect 150 336 151 337
rect 149 336 150 337
rect 148 336 149 337
rect 147 336 148 337
rect 146 336 147 337
rect 145 336 146 337
rect 144 336 145 337
rect 143 336 144 337
rect 142 336 143 337
rect 141 336 142 337
rect 140 336 141 337
rect 139 336 140 337
rect 138 336 139 337
rect 137 336 138 337
rect 136 336 137 337
rect 135 336 136 337
rect 134 336 135 337
rect 133 336 134 337
rect 132 336 133 337
rect 131 336 132 337
rect 130 336 131 337
rect 129 336 130 337
rect 128 336 129 337
rect 127 336 128 337
rect 126 336 127 337
rect 125 336 126 337
rect 124 336 125 337
rect 123 336 124 337
rect 122 336 123 337
rect 121 336 122 337
rect 120 336 121 337
rect 119 336 120 337
rect 118 336 119 337
rect 117 336 118 337
rect 116 336 117 337
rect 115 336 116 337
rect 114 336 115 337
rect 113 336 114 337
rect 112 336 113 337
rect 111 336 112 337
rect 110 336 111 337
rect 109 336 110 337
rect 88 336 89 337
rect 87 336 88 337
rect 86 336 87 337
rect 85 336 86 337
rect 84 336 85 337
rect 83 336 84 337
rect 82 336 83 337
rect 81 336 82 337
rect 80 336 81 337
rect 79 336 80 337
rect 78 336 79 337
rect 77 336 78 337
rect 76 336 77 337
rect 75 336 76 337
rect 74 336 75 337
rect 73 336 74 337
rect 72 336 73 337
rect 71 336 72 337
rect 70 336 71 337
rect 69 336 70 337
rect 68 336 69 337
rect 67 336 68 337
rect 66 336 67 337
rect 65 336 66 337
rect 64 336 65 337
rect 63 336 64 337
rect 62 336 63 337
rect 61 336 62 337
rect 60 336 61 337
rect 59 336 60 337
rect 58 336 59 337
rect 57 336 58 337
rect 56 336 57 337
rect 55 336 56 337
rect 54 336 55 337
rect 53 336 54 337
rect 52 336 53 337
rect 40 336 41 337
rect 39 336 40 337
rect 38 336 39 337
rect 37 336 38 337
rect 36 336 37 337
rect 35 336 36 337
rect 34 336 35 337
rect 33 336 34 337
rect 32 336 33 337
rect 31 336 32 337
rect 437 337 438 338
rect 436 337 437 338
rect 435 337 436 338
rect 434 337 435 338
rect 433 337 434 338
rect 432 337 433 338
rect 431 337 432 338
rect 430 337 431 338
rect 429 337 430 338
rect 428 337 429 338
rect 427 337 428 338
rect 426 337 427 338
rect 425 337 426 338
rect 424 337 425 338
rect 423 337 424 338
rect 422 337 423 338
rect 421 337 422 338
rect 420 337 421 338
rect 419 337 420 338
rect 418 337 419 338
rect 417 337 418 338
rect 416 337 417 338
rect 415 337 416 338
rect 414 337 415 338
rect 413 337 414 338
rect 412 337 413 338
rect 411 337 412 338
rect 410 337 411 338
rect 409 337 410 338
rect 408 337 409 338
rect 407 337 408 338
rect 406 337 407 338
rect 405 337 406 338
rect 404 337 405 338
rect 403 337 404 338
rect 402 337 403 338
rect 401 337 402 338
rect 400 337 401 338
rect 399 337 400 338
rect 398 337 399 338
rect 397 337 398 338
rect 396 337 397 338
rect 395 337 396 338
rect 394 337 395 338
rect 393 337 394 338
rect 172 337 173 338
rect 171 337 172 338
rect 170 337 171 338
rect 169 337 170 338
rect 168 337 169 338
rect 167 337 168 338
rect 166 337 167 338
rect 165 337 166 338
rect 164 337 165 338
rect 163 337 164 338
rect 162 337 163 338
rect 161 337 162 338
rect 160 337 161 338
rect 159 337 160 338
rect 158 337 159 338
rect 157 337 158 338
rect 156 337 157 338
rect 155 337 156 338
rect 154 337 155 338
rect 153 337 154 338
rect 152 337 153 338
rect 151 337 152 338
rect 150 337 151 338
rect 149 337 150 338
rect 148 337 149 338
rect 147 337 148 338
rect 146 337 147 338
rect 145 337 146 338
rect 144 337 145 338
rect 143 337 144 338
rect 142 337 143 338
rect 141 337 142 338
rect 140 337 141 338
rect 139 337 140 338
rect 138 337 139 338
rect 137 337 138 338
rect 136 337 137 338
rect 135 337 136 338
rect 134 337 135 338
rect 133 337 134 338
rect 132 337 133 338
rect 131 337 132 338
rect 130 337 131 338
rect 129 337 130 338
rect 128 337 129 338
rect 127 337 128 338
rect 126 337 127 338
rect 125 337 126 338
rect 124 337 125 338
rect 123 337 124 338
rect 122 337 123 338
rect 121 337 122 338
rect 120 337 121 338
rect 119 337 120 338
rect 118 337 119 338
rect 117 337 118 338
rect 116 337 117 338
rect 115 337 116 338
rect 114 337 115 338
rect 113 337 114 338
rect 112 337 113 338
rect 111 337 112 338
rect 110 337 111 338
rect 89 337 90 338
rect 88 337 89 338
rect 87 337 88 338
rect 86 337 87 338
rect 85 337 86 338
rect 84 337 85 338
rect 83 337 84 338
rect 82 337 83 338
rect 81 337 82 338
rect 80 337 81 338
rect 79 337 80 338
rect 78 337 79 338
rect 77 337 78 338
rect 76 337 77 338
rect 75 337 76 338
rect 74 337 75 338
rect 73 337 74 338
rect 72 337 73 338
rect 71 337 72 338
rect 70 337 71 338
rect 69 337 70 338
rect 68 337 69 338
rect 67 337 68 338
rect 66 337 67 338
rect 65 337 66 338
rect 64 337 65 338
rect 63 337 64 338
rect 62 337 63 338
rect 61 337 62 338
rect 60 337 61 338
rect 59 337 60 338
rect 58 337 59 338
rect 57 337 58 338
rect 56 337 57 338
rect 55 337 56 338
rect 54 337 55 338
rect 53 337 54 338
rect 52 337 53 338
rect 40 337 41 338
rect 39 337 40 338
rect 38 337 39 338
rect 37 337 38 338
rect 36 337 37 338
rect 35 337 36 338
rect 34 337 35 338
rect 33 337 34 338
rect 32 337 33 338
rect 437 338 438 339
rect 436 338 437 339
rect 435 338 436 339
rect 434 338 435 339
rect 433 338 434 339
rect 432 338 433 339
rect 431 338 432 339
rect 430 338 431 339
rect 429 338 430 339
rect 428 338 429 339
rect 427 338 428 339
rect 426 338 427 339
rect 425 338 426 339
rect 424 338 425 339
rect 423 338 424 339
rect 422 338 423 339
rect 421 338 422 339
rect 420 338 421 339
rect 419 338 420 339
rect 418 338 419 339
rect 417 338 418 339
rect 416 338 417 339
rect 415 338 416 339
rect 414 338 415 339
rect 413 338 414 339
rect 412 338 413 339
rect 411 338 412 339
rect 410 338 411 339
rect 409 338 410 339
rect 408 338 409 339
rect 407 338 408 339
rect 406 338 407 339
rect 405 338 406 339
rect 404 338 405 339
rect 403 338 404 339
rect 402 338 403 339
rect 401 338 402 339
rect 400 338 401 339
rect 399 338 400 339
rect 398 338 399 339
rect 397 338 398 339
rect 396 338 397 339
rect 395 338 396 339
rect 394 338 395 339
rect 393 338 394 339
rect 170 338 171 339
rect 169 338 170 339
rect 168 338 169 339
rect 167 338 168 339
rect 166 338 167 339
rect 165 338 166 339
rect 164 338 165 339
rect 163 338 164 339
rect 162 338 163 339
rect 161 338 162 339
rect 160 338 161 339
rect 159 338 160 339
rect 158 338 159 339
rect 157 338 158 339
rect 156 338 157 339
rect 155 338 156 339
rect 154 338 155 339
rect 153 338 154 339
rect 152 338 153 339
rect 151 338 152 339
rect 150 338 151 339
rect 149 338 150 339
rect 148 338 149 339
rect 147 338 148 339
rect 146 338 147 339
rect 145 338 146 339
rect 144 338 145 339
rect 143 338 144 339
rect 142 338 143 339
rect 141 338 142 339
rect 140 338 141 339
rect 139 338 140 339
rect 138 338 139 339
rect 137 338 138 339
rect 136 338 137 339
rect 135 338 136 339
rect 134 338 135 339
rect 133 338 134 339
rect 132 338 133 339
rect 131 338 132 339
rect 130 338 131 339
rect 129 338 130 339
rect 128 338 129 339
rect 127 338 128 339
rect 126 338 127 339
rect 125 338 126 339
rect 124 338 125 339
rect 123 338 124 339
rect 122 338 123 339
rect 121 338 122 339
rect 120 338 121 339
rect 119 338 120 339
rect 118 338 119 339
rect 117 338 118 339
rect 116 338 117 339
rect 115 338 116 339
rect 114 338 115 339
rect 113 338 114 339
rect 112 338 113 339
rect 111 338 112 339
rect 89 338 90 339
rect 88 338 89 339
rect 87 338 88 339
rect 86 338 87 339
rect 85 338 86 339
rect 84 338 85 339
rect 83 338 84 339
rect 82 338 83 339
rect 81 338 82 339
rect 80 338 81 339
rect 79 338 80 339
rect 78 338 79 339
rect 77 338 78 339
rect 76 338 77 339
rect 75 338 76 339
rect 74 338 75 339
rect 73 338 74 339
rect 72 338 73 339
rect 71 338 72 339
rect 70 338 71 339
rect 69 338 70 339
rect 68 338 69 339
rect 67 338 68 339
rect 66 338 67 339
rect 65 338 66 339
rect 64 338 65 339
rect 63 338 64 339
rect 62 338 63 339
rect 61 338 62 339
rect 60 338 61 339
rect 59 338 60 339
rect 58 338 59 339
rect 57 338 58 339
rect 56 338 57 339
rect 55 338 56 339
rect 54 338 55 339
rect 53 338 54 339
rect 41 338 42 339
rect 40 338 41 339
rect 39 338 40 339
rect 38 338 39 339
rect 37 338 38 339
rect 36 338 37 339
rect 35 338 36 339
rect 34 338 35 339
rect 33 338 34 339
rect 437 339 438 340
rect 436 339 437 340
rect 435 339 436 340
rect 434 339 435 340
rect 433 339 434 340
rect 432 339 433 340
rect 431 339 432 340
rect 430 339 431 340
rect 429 339 430 340
rect 428 339 429 340
rect 427 339 428 340
rect 426 339 427 340
rect 425 339 426 340
rect 424 339 425 340
rect 423 339 424 340
rect 422 339 423 340
rect 421 339 422 340
rect 420 339 421 340
rect 419 339 420 340
rect 418 339 419 340
rect 417 339 418 340
rect 416 339 417 340
rect 415 339 416 340
rect 414 339 415 340
rect 413 339 414 340
rect 412 339 413 340
rect 411 339 412 340
rect 410 339 411 340
rect 409 339 410 340
rect 408 339 409 340
rect 407 339 408 340
rect 406 339 407 340
rect 405 339 406 340
rect 404 339 405 340
rect 403 339 404 340
rect 402 339 403 340
rect 401 339 402 340
rect 400 339 401 340
rect 399 339 400 340
rect 398 339 399 340
rect 397 339 398 340
rect 396 339 397 340
rect 395 339 396 340
rect 394 339 395 340
rect 393 339 394 340
rect 168 339 169 340
rect 167 339 168 340
rect 166 339 167 340
rect 165 339 166 340
rect 164 339 165 340
rect 163 339 164 340
rect 162 339 163 340
rect 161 339 162 340
rect 160 339 161 340
rect 159 339 160 340
rect 158 339 159 340
rect 157 339 158 340
rect 156 339 157 340
rect 155 339 156 340
rect 154 339 155 340
rect 153 339 154 340
rect 152 339 153 340
rect 151 339 152 340
rect 150 339 151 340
rect 149 339 150 340
rect 148 339 149 340
rect 147 339 148 340
rect 146 339 147 340
rect 145 339 146 340
rect 144 339 145 340
rect 143 339 144 340
rect 142 339 143 340
rect 141 339 142 340
rect 140 339 141 340
rect 139 339 140 340
rect 138 339 139 340
rect 137 339 138 340
rect 136 339 137 340
rect 135 339 136 340
rect 134 339 135 340
rect 133 339 134 340
rect 132 339 133 340
rect 131 339 132 340
rect 130 339 131 340
rect 129 339 130 340
rect 128 339 129 340
rect 127 339 128 340
rect 126 339 127 340
rect 125 339 126 340
rect 124 339 125 340
rect 123 339 124 340
rect 122 339 123 340
rect 121 339 122 340
rect 120 339 121 340
rect 119 339 120 340
rect 118 339 119 340
rect 117 339 118 340
rect 116 339 117 340
rect 115 339 116 340
rect 114 339 115 340
rect 113 339 114 340
rect 112 339 113 340
rect 90 339 91 340
rect 89 339 90 340
rect 88 339 89 340
rect 87 339 88 340
rect 86 339 87 340
rect 85 339 86 340
rect 84 339 85 340
rect 83 339 84 340
rect 82 339 83 340
rect 81 339 82 340
rect 80 339 81 340
rect 79 339 80 340
rect 78 339 79 340
rect 77 339 78 340
rect 76 339 77 340
rect 75 339 76 340
rect 74 339 75 340
rect 73 339 74 340
rect 72 339 73 340
rect 71 339 72 340
rect 70 339 71 340
rect 69 339 70 340
rect 68 339 69 340
rect 67 339 68 340
rect 66 339 67 340
rect 65 339 66 340
rect 64 339 65 340
rect 63 339 64 340
rect 62 339 63 340
rect 61 339 62 340
rect 60 339 61 340
rect 59 339 60 340
rect 58 339 59 340
rect 57 339 58 340
rect 56 339 57 340
rect 55 339 56 340
rect 54 339 55 340
rect 53 339 54 340
rect 41 339 42 340
rect 40 339 41 340
rect 39 339 40 340
rect 38 339 39 340
rect 37 339 38 340
rect 36 339 37 340
rect 35 339 36 340
rect 437 340 438 341
rect 436 340 437 341
rect 435 340 436 341
rect 434 340 435 341
rect 433 340 434 341
rect 432 340 433 341
rect 431 340 432 341
rect 430 340 431 341
rect 429 340 430 341
rect 428 340 429 341
rect 427 340 428 341
rect 426 340 427 341
rect 425 340 426 341
rect 424 340 425 341
rect 423 340 424 341
rect 422 340 423 341
rect 421 340 422 341
rect 420 340 421 341
rect 419 340 420 341
rect 418 340 419 341
rect 417 340 418 341
rect 416 340 417 341
rect 415 340 416 341
rect 414 340 415 341
rect 413 340 414 341
rect 412 340 413 341
rect 411 340 412 341
rect 410 340 411 341
rect 409 340 410 341
rect 408 340 409 341
rect 407 340 408 341
rect 406 340 407 341
rect 405 340 406 341
rect 404 340 405 341
rect 403 340 404 341
rect 402 340 403 341
rect 401 340 402 341
rect 400 340 401 341
rect 399 340 400 341
rect 398 340 399 341
rect 397 340 398 341
rect 396 340 397 341
rect 395 340 396 341
rect 394 340 395 341
rect 393 340 394 341
rect 166 340 167 341
rect 165 340 166 341
rect 164 340 165 341
rect 163 340 164 341
rect 162 340 163 341
rect 161 340 162 341
rect 160 340 161 341
rect 159 340 160 341
rect 158 340 159 341
rect 157 340 158 341
rect 156 340 157 341
rect 155 340 156 341
rect 154 340 155 341
rect 153 340 154 341
rect 152 340 153 341
rect 151 340 152 341
rect 150 340 151 341
rect 149 340 150 341
rect 148 340 149 341
rect 147 340 148 341
rect 146 340 147 341
rect 145 340 146 341
rect 144 340 145 341
rect 143 340 144 341
rect 142 340 143 341
rect 141 340 142 341
rect 140 340 141 341
rect 139 340 140 341
rect 138 340 139 341
rect 137 340 138 341
rect 136 340 137 341
rect 135 340 136 341
rect 134 340 135 341
rect 133 340 134 341
rect 132 340 133 341
rect 131 340 132 341
rect 130 340 131 341
rect 129 340 130 341
rect 128 340 129 341
rect 127 340 128 341
rect 126 340 127 341
rect 125 340 126 341
rect 124 340 125 341
rect 123 340 124 341
rect 122 340 123 341
rect 121 340 122 341
rect 120 340 121 341
rect 119 340 120 341
rect 118 340 119 341
rect 117 340 118 341
rect 116 340 117 341
rect 115 340 116 341
rect 114 340 115 341
rect 113 340 114 341
rect 91 340 92 341
rect 90 340 91 341
rect 89 340 90 341
rect 88 340 89 341
rect 87 340 88 341
rect 86 340 87 341
rect 85 340 86 341
rect 84 340 85 341
rect 83 340 84 341
rect 82 340 83 341
rect 81 340 82 341
rect 80 340 81 341
rect 79 340 80 341
rect 78 340 79 341
rect 77 340 78 341
rect 76 340 77 341
rect 75 340 76 341
rect 74 340 75 341
rect 73 340 74 341
rect 72 340 73 341
rect 71 340 72 341
rect 70 340 71 341
rect 69 340 70 341
rect 68 340 69 341
rect 67 340 68 341
rect 66 340 67 341
rect 65 340 66 341
rect 64 340 65 341
rect 63 340 64 341
rect 62 340 63 341
rect 61 340 62 341
rect 60 340 61 341
rect 59 340 60 341
rect 58 340 59 341
rect 57 340 58 341
rect 56 340 57 341
rect 55 340 56 341
rect 54 340 55 341
rect 53 340 54 341
rect 42 340 43 341
rect 41 340 42 341
rect 40 340 41 341
rect 39 340 40 341
rect 38 340 39 341
rect 37 340 38 341
rect 36 340 37 341
rect 437 341 438 342
rect 436 341 437 342
rect 435 341 436 342
rect 434 341 435 342
rect 433 341 434 342
rect 432 341 433 342
rect 431 341 432 342
rect 430 341 431 342
rect 429 341 430 342
rect 428 341 429 342
rect 427 341 428 342
rect 426 341 427 342
rect 425 341 426 342
rect 424 341 425 342
rect 423 341 424 342
rect 422 341 423 342
rect 421 341 422 342
rect 420 341 421 342
rect 419 341 420 342
rect 418 341 419 342
rect 417 341 418 342
rect 416 341 417 342
rect 415 341 416 342
rect 414 341 415 342
rect 413 341 414 342
rect 412 341 413 342
rect 411 341 412 342
rect 410 341 411 342
rect 409 341 410 342
rect 408 341 409 342
rect 407 341 408 342
rect 406 341 407 342
rect 405 341 406 342
rect 404 341 405 342
rect 403 341 404 342
rect 402 341 403 342
rect 401 341 402 342
rect 400 341 401 342
rect 399 341 400 342
rect 398 341 399 342
rect 397 341 398 342
rect 396 341 397 342
rect 395 341 396 342
rect 394 341 395 342
rect 393 341 394 342
rect 164 341 165 342
rect 163 341 164 342
rect 162 341 163 342
rect 161 341 162 342
rect 160 341 161 342
rect 159 341 160 342
rect 158 341 159 342
rect 157 341 158 342
rect 156 341 157 342
rect 155 341 156 342
rect 154 341 155 342
rect 153 341 154 342
rect 152 341 153 342
rect 151 341 152 342
rect 150 341 151 342
rect 149 341 150 342
rect 148 341 149 342
rect 147 341 148 342
rect 146 341 147 342
rect 145 341 146 342
rect 144 341 145 342
rect 143 341 144 342
rect 142 341 143 342
rect 141 341 142 342
rect 140 341 141 342
rect 139 341 140 342
rect 138 341 139 342
rect 137 341 138 342
rect 136 341 137 342
rect 135 341 136 342
rect 134 341 135 342
rect 133 341 134 342
rect 132 341 133 342
rect 131 341 132 342
rect 130 341 131 342
rect 129 341 130 342
rect 128 341 129 342
rect 127 341 128 342
rect 126 341 127 342
rect 125 341 126 342
rect 124 341 125 342
rect 123 341 124 342
rect 122 341 123 342
rect 121 341 122 342
rect 120 341 121 342
rect 119 341 120 342
rect 118 341 119 342
rect 117 341 118 342
rect 116 341 117 342
rect 115 341 116 342
rect 92 341 93 342
rect 91 341 92 342
rect 90 341 91 342
rect 89 341 90 342
rect 88 341 89 342
rect 87 341 88 342
rect 86 341 87 342
rect 85 341 86 342
rect 84 341 85 342
rect 83 341 84 342
rect 82 341 83 342
rect 81 341 82 342
rect 80 341 81 342
rect 79 341 80 342
rect 78 341 79 342
rect 77 341 78 342
rect 76 341 77 342
rect 75 341 76 342
rect 74 341 75 342
rect 73 341 74 342
rect 72 341 73 342
rect 71 341 72 342
rect 70 341 71 342
rect 69 341 70 342
rect 68 341 69 342
rect 67 341 68 342
rect 66 341 67 342
rect 65 341 66 342
rect 64 341 65 342
rect 63 341 64 342
rect 62 341 63 342
rect 61 341 62 342
rect 60 341 61 342
rect 59 341 60 342
rect 58 341 59 342
rect 57 341 58 342
rect 56 341 57 342
rect 55 341 56 342
rect 54 341 55 342
rect 42 341 43 342
rect 41 341 42 342
rect 40 341 41 342
rect 39 341 40 342
rect 38 341 39 342
rect 437 342 438 343
rect 436 342 437 343
rect 435 342 436 343
rect 434 342 435 343
rect 433 342 434 343
rect 432 342 433 343
rect 431 342 432 343
rect 430 342 431 343
rect 429 342 430 343
rect 428 342 429 343
rect 427 342 428 343
rect 426 342 427 343
rect 425 342 426 343
rect 424 342 425 343
rect 423 342 424 343
rect 422 342 423 343
rect 421 342 422 343
rect 420 342 421 343
rect 419 342 420 343
rect 418 342 419 343
rect 417 342 418 343
rect 416 342 417 343
rect 415 342 416 343
rect 414 342 415 343
rect 413 342 414 343
rect 412 342 413 343
rect 411 342 412 343
rect 410 342 411 343
rect 409 342 410 343
rect 408 342 409 343
rect 407 342 408 343
rect 406 342 407 343
rect 405 342 406 343
rect 404 342 405 343
rect 403 342 404 343
rect 402 342 403 343
rect 401 342 402 343
rect 400 342 401 343
rect 399 342 400 343
rect 398 342 399 343
rect 397 342 398 343
rect 396 342 397 343
rect 395 342 396 343
rect 394 342 395 343
rect 393 342 394 343
rect 161 342 162 343
rect 160 342 161 343
rect 159 342 160 343
rect 158 342 159 343
rect 157 342 158 343
rect 156 342 157 343
rect 155 342 156 343
rect 154 342 155 343
rect 153 342 154 343
rect 152 342 153 343
rect 151 342 152 343
rect 150 342 151 343
rect 149 342 150 343
rect 148 342 149 343
rect 147 342 148 343
rect 146 342 147 343
rect 145 342 146 343
rect 144 342 145 343
rect 143 342 144 343
rect 142 342 143 343
rect 141 342 142 343
rect 140 342 141 343
rect 139 342 140 343
rect 138 342 139 343
rect 137 342 138 343
rect 136 342 137 343
rect 135 342 136 343
rect 134 342 135 343
rect 133 342 134 343
rect 132 342 133 343
rect 131 342 132 343
rect 130 342 131 343
rect 129 342 130 343
rect 128 342 129 343
rect 127 342 128 343
rect 126 342 127 343
rect 125 342 126 343
rect 124 342 125 343
rect 123 342 124 343
rect 122 342 123 343
rect 121 342 122 343
rect 120 342 121 343
rect 119 342 120 343
rect 118 342 119 343
rect 117 342 118 343
rect 116 342 117 343
rect 93 342 94 343
rect 92 342 93 343
rect 91 342 92 343
rect 90 342 91 343
rect 89 342 90 343
rect 88 342 89 343
rect 87 342 88 343
rect 86 342 87 343
rect 85 342 86 343
rect 84 342 85 343
rect 83 342 84 343
rect 82 342 83 343
rect 81 342 82 343
rect 80 342 81 343
rect 79 342 80 343
rect 78 342 79 343
rect 77 342 78 343
rect 76 342 77 343
rect 75 342 76 343
rect 74 342 75 343
rect 73 342 74 343
rect 72 342 73 343
rect 71 342 72 343
rect 70 342 71 343
rect 69 342 70 343
rect 68 342 69 343
rect 67 342 68 343
rect 66 342 67 343
rect 65 342 66 343
rect 64 342 65 343
rect 63 342 64 343
rect 62 342 63 343
rect 61 342 62 343
rect 60 342 61 343
rect 59 342 60 343
rect 58 342 59 343
rect 57 342 58 343
rect 56 342 57 343
rect 55 342 56 343
rect 54 342 55 343
rect 43 342 44 343
rect 42 342 43 343
rect 41 342 42 343
rect 437 343 438 344
rect 436 343 437 344
rect 435 343 436 344
rect 434 343 435 344
rect 433 343 434 344
rect 432 343 433 344
rect 431 343 432 344
rect 430 343 431 344
rect 429 343 430 344
rect 428 343 429 344
rect 427 343 428 344
rect 426 343 427 344
rect 425 343 426 344
rect 424 343 425 344
rect 423 343 424 344
rect 422 343 423 344
rect 421 343 422 344
rect 420 343 421 344
rect 419 343 420 344
rect 418 343 419 344
rect 417 343 418 344
rect 416 343 417 344
rect 415 343 416 344
rect 414 343 415 344
rect 413 343 414 344
rect 412 343 413 344
rect 411 343 412 344
rect 410 343 411 344
rect 409 343 410 344
rect 408 343 409 344
rect 407 343 408 344
rect 406 343 407 344
rect 405 343 406 344
rect 404 343 405 344
rect 403 343 404 344
rect 402 343 403 344
rect 401 343 402 344
rect 400 343 401 344
rect 399 343 400 344
rect 398 343 399 344
rect 397 343 398 344
rect 396 343 397 344
rect 395 343 396 344
rect 394 343 395 344
rect 393 343 394 344
rect 158 343 159 344
rect 157 343 158 344
rect 156 343 157 344
rect 155 343 156 344
rect 154 343 155 344
rect 153 343 154 344
rect 152 343 153 344
rect 151 343 152 344
rect 150 343 151 344
rect 149 343 150 344
rect 148 343 149 344
rect 147 343 148 344
rect 146 343 147 344
rect 145 343 146 344
rect 144 343 145 344
rect 143 343 144 344
rect 142 343 143 344
rect 141 343 142 344
rect 140 343 141 344
rect 139 343 140 344
rect 138 343 139 344
rect 137 343 138 344
rect 136 343 137 344
rect 135 343 136 344
rect 134 343 135 344
rect 133 343 134 344
rect 132 343 133 344
rect 131 343 132 344
rect 130 343 131 344
rect 129 343 130 344
rect 128 343 129 344
rect 127 343 128 344
rect 126 343 127 344
rect 125 343 126 344
rect 124 343 125 344
rect 123 343 124 344
rect 122 343 123 344
rect 121 343 122 344
rect 120 343 121 344
rect 119 343 120 344
rect 94 343 95 344
rect 93 343 94 344
rect 92 343 93 344
rect 91 343 92 344
rect 90 343 91 344
rect 89 343 90 344
rect 88 343 89 344
rect 87 343 88 344
rect 86 343 87 344
rect 85 343 86 344
rect 84 343 85 344
rect 83 343 84 344
rect 82 343 83 344
rect 81 343 82 344
rect 80 343 81 344
rect 79 343 80 344
rect 78 343 79 344
rect 77 343 78 344
rect 76 343 77 344
rect 75 343 76 344
rect 74 343 75 344
rect 73 343 74 344
rect 72 343 73 344
rect 71 343 72 344
rect 70 343 71 344
rect 69 343 70 344
rect 68 343 69 344
rect 67 343 68 344
rect 66 343 67 344
rect 65 343 66 344
rect 64 343 65 344
rect 63 343 64 344
rect 62 343 63 344
rect 61 343 62 344
rect 60 343 61 344
rect 59 343 60 344
rect 58 343 59 344
rect 57 343 58 344
rect 56 343 57 344
rect 55 343 56 344
rect 437 344 438 345
rect 436 344 437 345
rect 435 344 436 345
rect 434 344 435 345
rect 433 344 434 345
rect 432 344 433 345
rect 431 344 432 345
rect 430 344 431 345
rect 429 344 430 345
rect 428 344 429 345
rect 427 344 428 345
rect 426 344 427 345
rect 425 344 426 345
rect 424 344 425 345
rect 423 344 424 345
rect 422 344 423 345
rect 421 344 422 345
rect 420 344 421 345
rect 419 344 420 345
rect 418 344 419 345
rect 417 344 418 345
rect 416 344 417 345
rect 415 344 416 345
rect 414 344 415 345
rect 413 344 414 345
rect 412 344 413 345
rect 411 344 412 345
rect 410 344 411 345
rect 409 344 410 345
rect 408 344 409 345
rect 407 344 408 345
rect 406 344 407 345
rect 405 344 406 345
rect 404 344 405 345
rect 403 344 404 345
rect 402 344 403 345
rect 401 344 402 345
rect 400 344 401 345
rect 399 344 400 345
rect 398 344 399 345
rect 397 344 398 345
rect 396 344 397 345
rect 395 344 396 345
rect 394 344 395 345
rect 393 344 394 345
rect 154 344 155 345
rect 153 344 154 345
rect 152 344 153 345
rect 151 344 152 345
rect 150 344 151 345
rect 149 344 150 345
rect 148 344 149 345
rect 147 344 148 345
rect 146 344 147 345
rect 145 344 146 345
rect 144 344 145 345
rect 143 344 144 345
rect 142 344 143 345
rect 141 344 142 345
rect 140 344 141 345
rect 139 344 140 345
rect 138 344 139 345
rect 137 344 138 345
rect 136 344 137 345
rect 135 344 136 345
rect 134 344 135 345
rect 133 344 134 345
rect 132 344 133 345
rect 131 344 132 345
rect 130 344 131 345
rect 129 344 130 345
rect 128 344 129 345
rect 127 344 128 345
rect 126 344 127 345
rect 125 344 126 345
rect 124 344 125 345
rect 123 344 124 345
rect 122 344 123 345
rect 95 344 96 345
rect 94 344 95 345
rect 93 344 94 345
rect 92 344 93 345
rect 91 344 92 345
rect 90 344 91 345
rect 89 344 90 345
rect 88 344 89 345
rect 87 344 88 345
rect 86 344 87 345
rect 85 344 86 345
rect 84 344 85 345
rect 83 344 84 345
rect 82 344 83 345
rect 81 344 82 345
rect 80 344 81 345
rect 79 344 80 345
rect 78 344 79 345
rect 77 344 78 345
rect 76 344 77 345
rect 75 344 76 345
rect 74 344 75 345
rect 73 344 74 345
rect 72 344 73 345
rect 71 344 72 345
rect 70 344 71 345
rect 69 344 70 345
rect 68 344 69 345
rect 67 344 68 345
rect 66 344 67 345
rect 65 344 66 345
rect 64 344 65 345
rect 63 344 64 345
rect 62 344 63 345
rect 61 344 62 345
rect 60 344 61 345
rect 59 344 60 345
rect 58 344 59 345
rect 57 344 58 345
rect 56 344 57 345
rect 55 344 56 345
rect 437 345 438 346
rect 436 345 437 346
rect 435 345 436 346
rect 434 345 435 346
rect 416 345 417 346
rect 415 345 416 346
rect 414 345 415 346
rect 413 345 414 346
rect 395 345 396 346
rect 394 345 395 346
rect 393 345 394 346
rect 148 345 149 346
rect 147 345 148 346
rect 146 345 147 346
rect 145 345 146 346
rect 144 345 145 346
rect 143 345 144 346
rect 142 345 143 346
rect 141 345 142 346
rect 140 345 141 346
rect 139 345 140 346
rect 138 345 139 346
rect 137 345 138 346
rect 136 345 137 346
rect 135 345 136 346
rect 134 345 135 346
rect 133 345 134 346
rect 132 345 133 346
rect 131 345 132 346
rect 130 345 131 346
rect 129 345 130 346
rect 128 345 129 346
rect 127 345 128 346
rect 96 345 97 346
rect 95 345 96 346
rect 94 345 95 346
rect 93 345 94 346
rect 92 345 93 346
rect 91 345 92 346
rect 90 345 91 346
rect 89 345 90 346
rect 88 345 89 346
rect 87 345 88 346
rect 86 345 87 346
rect 85 345 86 346
rect 84 345 85 346
rect 83 345 84 346
rect 82 345 83 346
rect 81 345 82 346
rect 80 345 81 346
rect 79 345 80 346
rect 78 345 79 346
rect 77 345 78 346
rect 76 345 77 346
rect 75 345 76 346
rect 74 345 75 346
rect 73 345 74 346
rect 72 345 73 346
rect 71 345 72 346
rect 70 345 71 346
rect 69 345 70 346
rect 68 345 69 346
rect 67 345 68 346
rect 66 345 67 346
rect 65 345 66 346
rect 64 345 65 346
rect 63 345 64 346
rect 62 345 63 346
rect 61 345 62 346
rect 60 345 61 346
rect 59 345 60 346
rect 58 345 59 346
rect 57 345 58 346
rect 56 345 57 346
rect 437 346 438 347
rect 436 346 437 347
rect 435 346 436 347
rect 434 346 435 347
rect 416 346 417 347
rect 415 346 416 347
rect 414 346 415 347
rect 413 346 414 347
rect 395 346 396 347
rect 394 346 395 347
rect 393 346 394 347
rect 97 346 98 347
rect 96 346 97 347
rect 95 346 96 347
rect 94 346 95 347
rect 93 346 94 347
rect 92 346 93 347
rect 91 346 92 347
rect 90 346 91 347
rect 89 346 90 347
rect 88 346 89 347
rect 87 346 88 347
rect 86 346 87 347
rect 85 346 86 347
rect 84 346 85 347
rect 83 346 84 347
rect 82 346 83 347
rect 81 346 82 347
rect 80 346 81 347
rect 79 346 80 347
rect 78 346 79 347
rect 77 346 78 347
rect 76 346 77 347
rect 75 346 76 347
rect 74 346 75 347
rect 73 346 74 347
rect 72 346 73 347
rect 71 346 72 347
rect 70 346 71 347
rect 69 346 70 347
rect 68 346 69 347
rect 67 346 68 347
rect 66 346 67 347
rect 65 346 66 347
rect 64 346 65 347
rect 63 346 64 347
rect 62 346 63 347
rect 61 346 62 347
rect 60 346 61 347
rect 59 346 60 347
rect 58 346 59 347
rect 57 346 58 347
rect 56 346 57 347
rect 437 347 438 348
rect 436 347 437 348
rect 435 347 436 348
rect 416 347 417 348
rect 415 347 416 348
rect 414 347 415 348
rect 413 347 414 348
rect 395 347 396 348
rect 394 347 395 348
rect 393 347 394 348
rect 98 347 99 348
rect 97 347 98 348
rect 96 347 97 348
rect 95 347 96 348
rect 94 347 95 348
rect 93 347 94 348
rect 92 347 93 348
rect 91 347 92 348
rect 90 347 91 348
rect 89 347 90 348
rect 88 347 89 348
rect 87 347 88 348
rect 86 347 87 348
rect 85 347 86 348
rect 84 347 85 348
rect 83 347 84 348
rect 82 347 83 348
rect 81 347 82 348
rect 80 347 81 348
rect 79 347 80 348
rect 78 347 79 348
rect 77 347 78 348
rect 76 347 77 348
rect 75 347 76 348
rect 74 347 75 348
rect 73 347 74 348
rect 72 347 73 348
rect 71 347 72 348
rect 70 347 71 348
rect 69 347 70 348
rect 68 347 69 348
rect 67 347 68 348
rect 66 347 67 348
rect 65 347 66 348
rect 64 347 65 348
rect 63 347 64 348
rect 62 347 63 348
rect 61 347 62 348
rect 60 347 61 348
rect 59 347 60 348
rect 58 347 59 348
rect 57 347 58 348
rect 56 347 57 348
rect 437 348 438 349
rect 436 348 437 349
rect 435 348 436 349
rect 416 348 417 349
rect 415 348 416 349
rect 414 348 415 349
rect 413 348 414 349
rect 395 348 396 349
rect 394 348 395 349
rect 393 348 394 349
rect 99 348 100 349
rect 98 348 99 349
rect 97 348 98 349
rect 96 348 97 349
rect 95 348 96 349
rect 94 348 95 349
rect 93 348 94 349
rect 92 348 93 349
rect 91 348 92 349
rect 90 348 91 349
rect 89 348 90 349
rect 88 348 89 349
rect 87 348 88 349
rect 86 348 87 349
rect 85 348 86 349
rect 84 348 85 349
rect 83 348 84 349
rect 82 348 83 349
rect 81 348 82 349
rect 80 348 81 349
rect 79 348 80 349
rect 78 348 79 349
rect 77 348 78 349
rect 76 348 77 349
rect 75 348 76 349
rect 74 348 75 349
rect 73 348 74 349
rect 72 348 73 349
rect 71 348 72 349
rect 70 348 71 349
rect 69 348 70 349
rect 68 348 69 349
rect 67 348 68 349
rect 66 348 67 349
rect 65 348 66 349
rect 64 348 65 349
rect 63 348 64 349
rect 62 348 63 349
rect 61 348 62 349
rect 60 348 61 349
rect 59 348 60 349
rect 58 348 59 349
rect 57 348 58 349
rect 437 349 438 350
rect 436 349 437 350
rect 435 349 436 350
rect 416 349 417 350
rect 415 349 416 350
rect 414 349 415 350
rect 413 349 414 350
rect 395 349 396 350
rect 394 349 395 350
rect 393 349 394 350
rect 101 349 102 350
rect 100 349 101 350
rect 99 349 100 350
rect 98 349 99 350
rect 97 349 98 350
rect 96 349 97 350
rect 95 349 96 350
rect 94 349 95 350
rect 93 349 94 350
rect 92 349 93 350
rect 91 349 92 350
rect 90 349 91 350
rect 89 349 90 350
rect 88 349 89 350
rect 87 349 88 350
rect 86 349 87 350
rect 85 349 86 350
rect 84 349 85 350
rect 83 349 84 350
rect 82 349 83 350
rect 81 349 82 350
rect 80 349 81 350
rect 79 349 80 350
rect 78 349 79 350
rect 77 349 78 350
rect 76 349 77 350
rect 75 349 76 350
rect 74 349 75 350
rect 73 349 74 350
rect 72 349 73 350
rect 71 349 72 350
rect 70 349 71 350
rect 69 349 70 350
rect 68 349 69 350
rect 67 349 68 350
rect 66 349 67 350
rect 65 349 66 350
rect 64 349 65 350
rect 63 349 64 350
rect 62 349 63 350
rect 61 349 62 350
rect 60 349 61 350
rect 59 349 60 350
rect 58 349 59 350
rect 437 350 438 351
rect 436 350 437 351
rect 435 350 436 351
rect 416 350 417 351
rect 415 350 416 351
rect 414 350 415 351
rect 413 350 414 351
rect 395 350 396 351
rect 394 350 395 351
rect 393 350 394 351
rect 102 350 103 351
rect 101 350 102 351
rect 100 350 101 351
rect 99 350 100 351
rect 98 350 99 351
rect 97 350 98 351
rect 96 350 97 351
rect 95 350 96 351
rect 94 350 95 351
rect 93 350 94 351
rect 92 350 93 351
rect 91 350 92 351
rect 90 350 91 351
rect 89 350 90 351
rect 88 350 89 351
rect 87 350 88 351
rect 86 350 87 351
rect 85 350 86 351
rect 84 350 85 351
rect 83 350 84 351
rect 82 350 83 351
rect 81 350 82 351
rect 80 350 81 351
rect 79 350 80 351
rect 78 350 79 351
rect 77 350 78 351
rect 76 350 77 351
rect 75 350 76 351
rect 74 350 75 351
rect 73 350 74 351
rect 72 350 73 351
rect 71 350 72 351
rect 70 350 71 351
rect 69 350 70 351
rect 68 350 69 351
rect 67 350 68 351
rect 66 350 67 351
rect 65 350 66 351
rect 64 350 65 351
rect 63 350 64 351
rect 62 350 63 351
rect 61 350 62 351
rect 60 350 61 351
rect 59 350 60 351
rect 437 351 438 352
rect 436 351 437 352
rect 435 351 436 352
rect 416 351 417 352
rect 415 351 416 352
rect 414 351 415 352
rect 413 351 414 352
rect 395 351 396 352
rect 394 351 395 352
rect 393 351 394 352
rect 103 351 104 352
rect 102 351 103 352
rect 101 351 102 352
rect 100 351 101 352
rect 99 351 100 352
rect 98 351 99 352
rect 97 351 98 352
rect 96 351 97 352
rect 95 351 96 352
rect 94 351 95 352
rect 93 351 94 352
rect 92 351 93 352
rect 91 351 92 352
rect 90 351 91 352
rect 89 351 90 352
rect 88 351 89 352
rect 87 351 88 352
rect 86 351 87 352
rect 85 351 86 352
rect 84 351 85 352
rect 83 351 84 352
rect 82 351 83 352
rect 81 351 82 352
rect 80 351 81 352
rect 79 351 80 352
rect 78 351 79 352
rect 77 351 78 352
rect 76 351 77 352
rect 75 351 76 352
rect 74 351 75 352
rect 73 351 74 352
rect 72 351 73 352
rect 71 351 72 352
rect 70 351 71 352
rect 69 351 70 352
rect 68 351 69 352
rect 67 351 68 352
rect 66 351 67 352
rect 65 351 66 352
rect 64 351 65 352
rect 63 351 64 352
rect 62 351 63 352
rect 61 351 62 352
rect 60 351 61 352
rect 59 351 60 352
rect 437 352 438 353
rect 436 352 437 353
rect 435 352 436 353
rect 416 352 417 353
rect 415 352 416 353
rect 414 352 415 353
rect 413 352 414 353
rect 395 352 396 353
rect 394 352 395 353
rect 393 352 394 353
rect 105 352 106 353
rect 104 352 105 353
rect 103 352 104 353
rect 102 352 103 353
rect 101 352 102 353
rect 100 352 101 353
rect 99 352 100 353
rect 98 352 99 353
rect 97 352 98 353
rect 96 352 97 353
rect 95 352 96 353
rect 94 352 95 353
rect 93 352 94 353
rect 92 352 93 353
rect 91 352 92 353
rect 90 352 91 353
rect 89 352 90 353
rect 88 352 89 353
rect 87 352 88 353
rect 86 352 87 353
rect 85 352 86 353
rect 84 352 85 353
rect 83 352 84 353
rect 82 352 83 353
rect 81 352 82 353
rect 80 352 81 353
rect 79 352 80 353
rect 78 352 79 353
rect 77 352 78 353
rect 76 352 77 353
rect 75 352 76 353
rect 74 352 75 353
rect 73 352 74 353
rect 72 352 73 353
rect 71 352 72 353
rect 70 352 71 353
rect 69 352 70 353
rect 68 352 69 353
rect 67 352 68 353
rect 66 352 67 353
rect 65 352 66 353
rect 64 352 65 353
rect 63 352 64 353
rect 62 352 63 353
rect 61 352 62 353
rect 437 353 438 354
rect 436 353 437 354
rect 435 353 436 354
rect 416 353 417 354
rect 415 353 416 354
rect 414 353 415 354
rect 413 353 414 354
rect 395 353 396 354
rect 394 353 395 354
rect 393 353 394 354
rect 106 353 107 354
rect 105 353 106 354
rect 104 353 105 354
rect 103 353 104 354
rect 102 353 103 354
rect 101 353 102 354
rect 100 353 101 354
rect 99 353 100 354
rect 98 353 99 354
rect 97 353 98 354
rect 96 353 97 354
rect 95 353 96 354
rect 94 353 95 354
rect 93 353 94 354
rect 92 353 93 354
rect 91 353 92 354
rect 90 353 91 354
rect 89 353 90 354
rect 88 353 89 354
rect 87 353 88 354
rect 86 353 87 354
rect 85 353 86 354
rect 84 353 85 354
rect 83 353 84 354
rect 82 353 83 354
rect 81 353 82 354
rect 80 353 81 354
rect 79 353 80 354
rect 78 353 79 354
rect 77 353 78 354
rect 76 353 77 354
rect 75 353 76 354
rect 74 353 75 354
rect 73 353 74 354
rect 72 353 73 354
rect 71 353 72 354
rect 70 353 71 354
rect 69 353 70 354
rect 68 353 69 354
rect 67 353 68 354
rect 66 353 67 354
rect 65 353 66 354
rect 64 353 65 354
rect 63 353 64 354
rect 62 353 63 354
rect 437 354 438 355
rect 436 354 437 355
rect 435 354 436 355
rect 416 354 417 355
rect 415 354 416 355
rect 414 354 415 355
rect 413 354 414 355
rect 396 354 397 355
rect 395 354 396 355
rect 394 354 395 355
rect 393 354 394 355
rect 108 354 109 355
rect 107 354 108 355
rect 106 354 107 355
rect 105 354 106 355
rect 104 354 105 355
rect 103 354 104 355
rect 102 354 103 355
rect 101 354 102 355
rect 100 354 101 355
rect 99 354 100 355
rect 98 354 99 355
rect 97 354 98 355
rect 96 354 97 355
rect 95 354 96 355
rect 94 354 95 355
rect 93 354 94 355
rect 92 354 93 355
rect 91 354 92 355
rect 90 354 91 355
rect 89 354 90 355
rect 88 354 89 355
rect 87 354 88 355
rect 86 354 87 355
rect 85 354 86 355
rect 84 354 85 355
rect 83 354 84 355
rect 82 354 83 355
rect 81 354 82 355
rect 80 354 81 355
rect 79 354 80 355
rect 78 354 79 355
rect 77 354 78 355
rect 76 354 77 355
rect 75 354 76 355
rect 74 354 75 355
rect 73 354 74 355
rect 72 354 73 355
rect 71 354 72 355
rect 70 354 71 355
rect 69 354 70 355
rect 68 354 69 355
rect 67 354 68 355
rect 66 354 67 355
rect 65 354 66 355
rect 64 354 65 355
rect 63 354 64 355
rect 437 355 438 356
rect 436 355 437 356
rect 435 355 436 356
rect 417 355 418 356
rect 416 355 417 356
rect 415 355 416 356
rect 414 355 415 356
rect 413 355 414 356
rect 412 355 413 356
rect 396 355 397 356
rect 395 355 396 356
rect 394 355 395 356
rect 393 355 394 356
rect 109 355 110 356
rect 108 355 109 356
rect 107 355 108 356
rect 106 355 107 356
rect 105 355 106 356
rect 104 355 105 356
rect 103 355 104 356
rect 102 355 103 356
rect 101 355 102 356
rect 100 355 101 356
rect 99 355 100 356
rect 98 355 99 356
rect 97 355 98 356
rect 96 355 97 356
rect 95 355 96 356
rect 94 355 95 356
rect 93 355 94 356
rect 92 355 93 356
rect 91 355 92 356
rect 90 355 91 356
rect 89 355 90 356
rect 88 355 89 356
rect 87 355 88 356
rect 86 355 87 356
rect 85 355 86 356
rect 84 355 85 356
rect 83 355 84 356
rect 82 355 83 356
rect 81 355 82 356
rect 80 355 81 356
rect 79 355 80 356
rect 78 355 79 356
rect 77 355 78 356
rect 76 355 77 356
rect 75 355 76 356
rect 74 355 75 356
rect 73 355 74 356
rect 72 355 73 356
rect 71 355 72 356
rect 70 355 71 356
rect 69 355 70 356
rect 68 355 69 356
rect 67 355 68 356
rect 66 355 67 356
rect 65 355 66 356
rect 437 356 438 357
rect 436 356 437 357
rect 435 356 436 357
rect 420 356 421 357
rect 419 356 420 357
rect 418 356 419 357
rect 417 356 418 357
rect 416 356 417 357
rect 415 356 416 357
rect 414 356 415 357
rect 413 356 414 357
rect 412 356 413 357
rect 411 356 412 357
rect 410 356 411 357
rect 409 356 410 357
rect 396 356 397 357
rect 395 356 396 357
rect 394 356 395 357
rect 393 356 394 357
rect 111 356 112 357
rect 110 356 111 357
rect 109 356 110 357
rect 108 356 109 357
rect 107 356 108 357
rect 106 356 107 357
rect 105 356 106 357
rect 104 356 105 357
rect 103 356 104 357
rect 102 356 103 357
rect 101 356 102 357
rect 100 356 101 357
rect 99 356 100 357
rect 98 356 99 357
rect 97 356 98 357
rect 96 356 97 357
rect 95 356 96 357
rect 94 356 95 357
rect 93 356 94 357
rect 92 356 93 357
rect 91 356 92 357
rect 90 356 91 357
rect 89 356 90 357
rect 88 356 89 357
rect 87 356 88 357
rect 86 356 87 357
rect 85 356 86 357
rect 84 356 85 357
rect 83 356 84 357
rect 82 356 83 357
rect 81 356 82 357
rect 80 356 81 357
rect 79 356 80 357
rect 78 356 79 357
rect 77 356 78 357
rect 76 356 77 357
rect 75 356 76 357
rect 74 356 75 357
rect 73 356 74 357
rect 72 356 73 357
rect 71 356 72 357
rect 70 356 71 357
rect 69 356 70 357
rect 68 356 69 357
rect 67 356 68 357
rect 437 357 438 358
rect 436 357 437 358
rect 435 357 436 358
rect 434 357 435 358
rect 421 357 422 358
rect 420 357 421 358
rect 419 357 420 358
rect 418 357 419 358
rect 417 357 418 358
rect 416 357 417 358
rect 415 357 416 358
rect 414 357 415 358
rect 413 357 414 358
rect 412 357 413 358
rect 411 357 412 358
rect 410 357 411 358
rect 409 357 410 358
rect 408 357 409 358
rect 397 357 398 358
rect 396 357 397 358
rect 395 357 396 358
rect 394 357 395 358
rect 393 357 394 358
rect 113 357 114 358
rect 112 357 113 358
rect 111 357 112 358
rect 110 357 111 358
rect 109 357 110 358
rect 108 357 109 358
rect 107 357 108 358
rect 106 357 107 358
rect 105 357 106 358
rect 104 357 105 358
rect 103 357 104 358
rect 102 357 103 358
rect 101 357 102 358
rect 100 357 101 358
rect 99 357 100 358
rect 98 357 99 358
rect 97 357 98 358
rect 96 357 97 358
rect 95 357 96 358
rect 94 357 95 358
rect 93 357 94 358
rect 92 357 93 358
rect 91 357 92 358
rect 90 357 91 358
rect 89 357 90 358
rect 88 357 89 358
rect 87 357 88 358
rect 86 357 87 358
rect 85 357 86 358
rect 84 357 85 358
rect 83 357 84 358
rect 82 357 83 358
rect 81 357 82 358
rect 80 357 81 358
rect 79 357 80 358
rect 78 357 79 358
rect 77 357 78 358
rect 76 357 77 358
rect 75 357 76 358
rect 74 357 75 358
rect 73 357 74 358
rect 72 357 73 358
rect 71 357 72 358
rect 70 357 71 358
rect 69 357 70 358
rect 437 358 438 359
rect 436 358 437 359
rect 435 358 436 359
rect 434 358 435 359
rect 421 358 422 359
rect 420 358 421 359
rect 419 358 420 359
rect 418 358 419 359
rect 417 358 418 359
rect 416 358 417 359
rect 415 358 416 359
rect 414 358 415 359
rect 413 358 414 359
rect 412 358 413 359
rect 411 358 412 359
rect 410 358 411 359
rect 409 358 410 359
rect 408 358 409 359
rect 398 358 399 359
rect 397 358 398 359
rect 396 358 397 359
rect 395 358 396 359
rect 394 358 395 359
rect 393 358 394 359
rect 115 358 116 359
rect 114 358 115 359
rect 113 358 114 359
rect 112 358 113 359
rect 111 358 112 359
rect 110 358 111 359
rect 109 358 110 359
rect 108 358 109 359
rect 107 358 108 359
rect 106 358 107 359
rect 105 358 106 359
rect 104 358 105 359
rect 103 358 104 359
rect 102 358 103 359
rect 101 358 102 359
rect 100 358 101 359
rect 99 358 100 359
rect 98 358 99 359
rect 97 358 98 359
rect 96 358 97 359
rect 95 358 96 359
rect 94 358 95 359
rect 93 358 94 359
rect 92 358 93 359
rect 91 358 92 359
rect 90 358 91 359
rect 89 358 90 359
rect 88 358 89 359
rect 87 358 88 359
rect 86 358 87 359
rect 85 358 86 359
rect 84 358 85 359
rect 83 358 84 359
rect 82 358 83 359
rect 81 358 82 359
rect 80 358 81 359
rect 79 358 80 359
rect 78 358 79 359
rect 77 358 78 359
rect 76 358 77 359
rect 75 358 76 359
rect 74 358 75 359
rect 73 358 74 359
rect 72 358 73 359
rect 71 358 72 359
rect 437 359 438 360
rect 436 359 437 360
rect 435 359 436 360
rect 434 359 435 360
rect 433 359 434 360
rect 400 359 401 360
rect 399 359 400 360
rect 398 359 399 360
rect 397 359 398 360
rect 396 359 397 360
rect 395 359 396 360
rect 394 359 395 360
rect 393 359 394 360
rect 114 359 115 360
rect 113 359 114 360
rect 112 359 113 360
rect 111 359 112 360
rect 110 359 111 360
rect 109 359 110 360
rect 108 359 109 360
rect 107 359 108 360
rect 106 359 107 360
rect 105 359 106 360
rect 104 359 105 360
rect 103 359 104 360
rect 102 359 103 360
rect 101 359 102 360
rect 100 359 101 360
rect 99 359 100 360
rect 98 359 99 360
rect 97 359 98 360
rect 96 359 97 360
rect 95 359 96 360
rect 94 359 95 360
rect 93 359 94 360
rect 92 359 93 360
rect 91 359 92 360
rect 90 359 91 360
rect 89 359 90 360
rect 88 359 89 360
rect 87 359 88 360
rect 86 359 87 360
rect 85 359 86 360
rect 84 359 85 360
rect 83 359 84 360
rect 82 359 83 360
rect 81 359 82 360
rect 80 359 81 360
rect 79 359 80 360
rect 78 359 79 360
rect 77 359 78 360
rect 76 359 77 360
rect 75 359 76 360
rect 74 359 75 360
rect 437 360 438 361
rect 436 360 437 361
rect 435 360 436 361
rect 434 360 435 361
rect 433 360 434 361
rect 432 360 433 361
rect 403 360 404 361
rect 402 360 403 361
rect 401 360 402 361
rect 400 360 401 361
rect 399 360 400 361
rect 398 360 399 361
rect 397 360 398 361
rect 396 360 397 361
rect 395 360 396 361
rect 394 360 395 361
rect 393 360 394 361
rect 112 360 113 361
rect 111 360 112 361
rect 110 360 111 361
rect 109 360 110 361
rect 108 360 109 361
rect 107 360 108 361
rect 106 360 107 361
rect 105 360 106 361
rect 104 360 105 361
rect 103 360 104 361
rect 102 360 103 361
rect 101 360 102 361
rect 100 360 101 361
rect 99 360 100 361
rect 98 360 99 361
rect 97 360 98 361
rect 96 360 97 361
rect 95 360 96 361
rect 94 360 95 361
rect 93 360 94 361
rect 92 360 93 361
rect 91 360 92 361
rect 90 360 91 361
rect 89 360 90 361
rect 88 360 89 361
rect 87 360 88 361
rect 86 360 87 361
rect 85 360 86 361
rect 84 360 85 361
rect 83 360 84 361
rect 82 360 83 361
rect 81 360 82 361
rect 80 360 81 361
rect 79 360 80 361
rect 78 360 79 361
rect 437 361 438 362
rect 436 361 437 362
rect 435 361 436 362
rect 434 361 435 362
rect 433 361 434 362
rect 432 361 433 362
rect 431 361 432 362
rect 403 361 404 362
rect 402 361 403 362
rect 401 361 402 362
rect 400 361 401 362
rect 399 361 400 362
rect 398 361 399 362
rect 397 361 398 362
rect 396 361 397 362
rect 395 361 396 362
rect 394 361 395 362
rect 393 361 394 362
rect 109 361 110 362
rect 108 361 109 362
rect 107 361 108 362
rect 106 361 107 362
rect 105 361 106 362
rect 104 361 105 362
rect 103 361 104 362
rect 102 361 103 362
rect 101 361 102 362
rect 100 361 101 362
rect 99 361 100 362
rect 98 361 99 362
rect 97 361 98 362
rect 96 361 97 362
rect 95 361 96 362
rect 94 361 95 362
rect 93 361 94 362
rect 92 361 93 362
rect 91 361 92 362
rect 90 361 91 362
rect 89 361 90 362
rect 88 361 89 362
rect 87 361 88 362
rect 86 361 87 362
rect 85 361 86 362
rect 84 361 85 362
rect 83 361 84 362
rect 82 361 83 362
rect 437 362 438 363
rect 436 362 437 363
rect 435 362 436 363
rect 434 362 435 363
rect 433 362 434 363
rect 432 362 433 363
rect 431 362 432 363
rect 430 362 431 363
rect 429 362 430 363
rect 403 362 404 363
rect 402 362 403 363
rect 401 362 402 363
rect 400 362 401 363
rect 399 362 400 363
rect 398 362 399 363
rect 397 362 398 363
rect 396 362 397 363
rect 395 362 396 363
rect 103 362 104 363
rect 102 362 103 363
rect 101 362 102 363
rect 100 362 101 363
rect 99 362 100 363
rect 98 362 99 363
rect 97 362 98 363
rect 96 362 97 363
rect 95 362 96 363
rect 94 362 95 363
rect 93 362 94 363
rect 92 362 93 363
rect 91 362 92 363
rect 90 362 91 363
rect 89 362 90 363
rect 437 363 438 364
rect 436 363 437 364
rect 435 363 436 364
rect 434 363 435 364
rect 433 363 434 364
rect 432 363 433 364
rect 431 363 432 364
rect 430 363 431 364
rect 429 363 430 364
rect 428 363 429 364
rect 427 363 428 364
rect 436 364 437 365
rect 435 364 436 365
rect 434 364 435 365
rect 433 364 434 365
rect 432 364 433 365
rect 431 364 432 365
rect 430 364 431 365
rect 429 364 430 365
rect 428 364 429 365
rect 427 364 428 365
rect 426 364 427 365
rect 431 365 432 366
rect 430 365 431 366
rect 429 365 430 366
rect 428 365 429 366
rect 427 365 428 366
rect 426 365 427 366
rect 437 372 438 373
rect 436 372 437 373
rect 437 373 438 374
rect 436 373 437 374
rect 435 373 436 374
rect 395 373 396 374
rect 394 373 395 374
rect 393 373 394 374
rect 437 374 438 375
rect 436 374 437 375
rect 435 374 436 375
rect 395 374 396 375
rect 394 374 395 375
rect 393 374 394 375
rect 437 375 438 376
rect 436 375 437 376
rect 435 375 436 376
rect 395 375 396 376
rect 394 375 395 376
rect 393 375 394 376
rect 437 376 438 377
rect 436 376 437 377
rect 435 376 436 377
rect 395 376 396 377
rect 394 376 395 377
rect 393 376 394 377
rect 437 377 438 378
rect 436 377 437 378
rect 435 377 436 378
rect 434 377 435 378
rect 396 377 397 378
rect 395 377 396 378
rect 394 377 395 378
rect 393 377 394 378
rect 437 378 438 379
rect 436 378 437 379
rect 435 378 436 379
rect 434 378 435 379
rect 433 378 434 379
rect 432 378 433 379
rect 431 378 432 379
rect 430 378 431 379
rect 429 378 430 379
rect 428 378 429 379
rect 427 378 428 379
rect 426 378 427 379
rect 425 378 426 379
rect 424 378 425 379
rect 423 378 424 379
rect 422 378 423 379
rect 421 378 422 379
rect 420 378 421 379
rect 419 378 420 379
rect 418 378 419 379
rect 417 378 418 379
rect 416 378 417 379
rect 415 378 416 379
rect 414 378 415 379
rect 413 378 414 379
rect 412 378 413 379
rect 411 378 412 379
rect 410 378 411 379
rect 409 378 410 379
rect 408 378 409 379
rect 407 378 408 379
rect 406 378 407 379
rect 405 378 406 379
rect 404 378 405 379
rect 403 378 404 379
rect 402 378 403 379
rect 401 378 402 379
rect 400 378 401 379
rect 399 378 400 379
rect 398 378 399 379
rect 397 378 398 379
rect 396 378 397 379
rect 395 378 396 379
rect 394 378 395 379
rect 393 378 394 379
rect 437 379 438 380
rect 436 379 437 380
rect 435 379 436 380
rect 434 379 435 380
rect 433 379 434 380
rect 432 379 433 380
rect 431 379 432 380
rect 430 379 431 380
rect 429 379 430 380
rect 428 379 429 380
rect 427 379 428 380
rect 426 379 427 380
rect 425 379 426 380
rect 424 379 425 380
rect 423 379 424 380
rect 422 379 423 380
rect 421 379 422 380
rect 420 379 421 380
rect 419 379 420 380
rect 418 379 419 380
rect 417 379 418 380
rect 416 379 417 380
rect 415 379 416 380
rect 414 379 415 380
rect 413 379 414 380
rect 412 379 413 380
rect 411 379 412 380
rect 410 379 411 380
rect 409 379 410 380
rect 408 379 409 380
rect 407 379 408 380
rect 406 379 407 380
rect 405 379 406 380
rect 404 379 405 380
rect 403 379 404 380
rect 402 379 403 380
rect 401 379 402 380
rect 400 379 401 380
rect 399 379 400 380
rect 398 379 399 380
rect 397 379 398 380
rect 396 379 397 380
rect 395 379 396 380
rect 394 379 395 380
rect 393 379 394 380
rect 437 380 438 381
rect 436 380 437 381
rect 435 380 436 381
rect 434 380 435 381
rect 433 380 434 381
rect 432 380 433 381
rect 431 380 432 381
rect 430 380 431 381
rect 429 380 430 381
rect 428 380 429 381
rect 427 380 428 381
rect 426 380 427 381
rect 425 380 426 381
rect 424 380 425 381
rect 423 380 424 381
rect 422 380 423 381
rect 421 380 422 381
rect 420 380 421 381
rect 419 380 420 381
rect 418 380 419 381
rect 417 380 418 381
rect 416 380 417 381
rect 415 380 416 381
rect 414 380 415 381
rect 413 380 414 381
rect 412 380 413 381
rect 411 380 412 381
rect 410 380 411 381
rect 409 380 410 381
rect 408 380 409 381
rect 407 380 408 381
rect 406 380 407 381
rect 405 380 406 381
rect 404 380 405 381
rect 403 380 404 381
rect 402 380 403 381
rect 401 380 402 381
rect 400 380 401 381
rect 399 380 400 381
rect 398 380 399 381
rect 397 380 398 381
rect 396 380 397 381
rect 395 380 396 381
rect 394 380 395 381
rect 393 380 394 381
rect 437 381 438 382
rect 436 381 437 382
rect 435 381 436 382
rect 434 381 435 382
rect 433 381 434 382
rect 432 381 433 382
rect 431 381 432 382
rect 430 381 431 382
rect 429 381 430 382
rect 428 381 429 382
rect 427 381 428 382
rect 426 381 427 382
rect 425 381 426 382
rect 424 381 425 382
rect 423 381 424 382
rect 422 381 423 382
rect 421 381 422 382
rect 420 381 421 382
rect 419 381 420 382
rect 418 381 419 382
rect 417 381 418 382
rect 416 381 417 382
rect 415 381 416 382
rect 414 381 415 382
rect 413 381 414 382
rect 412 381 413 382
rect 411 381 412 382
rect 410 381 411 382
rect 409 381 410 382
rect 408 381 409 382
rect 407 381 408 382
rect 406 381 407 382
rect 405 381 406 382
rect 404 381 405 382
rect 403 381 404 382
rect 402 381 403 382
rect 401 381 402 382
rect 400 381 401 382
rect 399 381 400 382
rect 398 381 399 382
rect 397 381 398 382
rect 396 381 397 382
rect 395 381 396 382
rect 394 381 395 382
rect 393 381 394 382
rect 437 382 438 383
rect 436 382 437 383
rect 435 382 436 383
rect 434 382 435 383
rect 433 382 434 383
rect 432 382 433 383
rect 431 382 432 383
rect 430 382 431 383
rect 429 382 430 383
rect 428 382 429 383
rect 427 382 428 383
rect 426 382 427 383
rect 425 382 426 383
rect 424 382 425 383
rect 423 382 424 383
rect 422 382 423 383
rect 421 382 422 383
rect 420 382 421 383
rect 419 382 420 383
rect 418 382 419 383
rect 417 382 418 383
rect 416 382 417 383
rect 415 382 416 383
rect 414 382 415 383
rect 413 382 414 383
rect 412 382 413 383
rect 411 382 412 383
rect 410 382 411 383
rect 409 382 410 383
rect 408 382 409 383
rect 407 382 408 383
rect 406 382 407 383
rect 405 382 406 383
rect 404 382 405 383
rect 403 382 404 383
rect 402 382 403 383
rect 401 382 402 383
rect 400 382 401 383
rect 399 382 400 383
rect 398 382 399 383
rect 397 382 398 383
rect 396 382 397 383
rect 395 382 396 383
rect 394 382 395 383
rect 393 382 394 383
rect 437 383 438 384
rect 436 383 437 384
rect 435 383 436 384
rect 434 383 435 384
rect 433 383 434 384
rect 432 383 433 384
rect 431 383 432 384
rect 430 383 431 384
rect 429 383 430 384
rect 428 383 429 384
rect 427 383 428 384
rect 426 383 427 384
rect 425 383 426 384
rect 424 383 425 384
rect 423 383 424 384
rect 422 383 423 384
rect 421 383 422 384
rect 420 383 421 384
rect 419 383 420 384
rect 418 383 419 384
rect 417 383 418 384
rect 416 383 417 384
rect 415 383 416 384
rect 414 383 415 384
rect 413 383 414 384
rect 412 383 413 384
rect 411 383 412 384
rect 410 383 411 384
rect 409 383 410 384
rect 408 383 409 384
rect 407 383 408 384
rect 406 383 407 384
rect 405 383 406 384
rect 404 383 405 384
rect 403 383 404 384
rect 402 383 403 384
rect 401 383 402 384
rect 400 383 401 384
rect 399 383 400 384
rect 398 383 399 384
rect 397 383 398 384
rect 396 383 397 384
rect 395 383 396 384
rect 394 383 395 384
rect 393 383 394 384
rect 437 384 438 385
rect 436 384 437 385
rect 435 384 436 385
rect 434 384 435 385
rect 433 384 434 385
rect 432 384 433 385
rect 431 384 432 385
rect 430 384 431 385
rect 429 384 430 385
rect 428 384 429 385
rect 427 384 428 385
rect 426 384 427 385
rect 425 384 426 385
rect 424 384 425 385
rect 423 384 424 385
rect 422 384 423 385
rect 421 384 422 385
rect 420 384 421 385
rect 419 384 420 385
rect 418 384 419 385
rect 417 384 418 385
rect 416 384 417 385
rect 415 384 416 385
rect 414 384 415 385
rect 413 384 414 385
rect 412 384 413 385
rect 411 384 412 385
rect 410 384 411 385
rect 409 384 410 385
rect 408 384 409 385
rect 407 384 408 385
rect 406 384 407 385
rect 405 384 406 385
rect 404 384 405 385
rect 403 384 404 385
rect 402 384 403 385
rect 401 384 402 385
rect 400 384 401 385
rect 399 384 400 385
rect 398 384 399 385
rect 397 384 398 385
rect 396 384 397 385
rect 395 384 396 385
rect 394 384 395 385
rect 393 384 394 385
rect 437 385 438 386
rect 436 385 437 386
rect 435 385 436 386
rect 434 385 435 386
rect 433 385 434 386
rect 432 385 433 386
rect 431 385 432 386
rect 430 385 431 386
rect 429 385 430 386
rect 428 385 429 386
rect 427 385 428 386
rect 426 385 427 386
rect 425 385 426 386
rect 424 385 425 386
rect 423 385 424 386
rect 422 385 423 386
rect 421 385 422 386
rect 420 385 421 386
rect 419 385 420 386
rect 418 385 419 386
rect 417 385 418 386
rect 416 385 417 386
rect 415 385 416 386
rect 414 385 415 386
rect 413 385 414 386
rect 412 385 413 386
rect 411 385 412 386
rect 410 385 411 386
rect 409 385 410 386
rect 408 385 409 386
rect 407 385 408 386
rect 406 385 407 386
rect 405 385 406 386
rect 404 385 405 386
rect 403 385 404 386
rect 402 385 403 386
rect 401 385 402 386
rect 400 385 401 386
rect 399 385 400 386
rect 398 385 399 386
rect 397 385 398 386
rect 396 385 397 386
rect 395 385 396 386
rect 394 385 395 386
rect 393 385 394 386
rect 437 386 438 387
rect 436 386 437 387
rect 435 386 436 387
rect 434 386 435 387
rect 433 386 434 387
rect 432 386 433 387
rect 431 386 432 387
rect 430 386 431 387
rect 429 386 430 387
rect 428 386 429 387
rect 427 386 428 387
rect 426 386 427 387
rect 425 386 426 387
rect 424 386 425 387
rect 423 386 424 387
rect 422 386 423 387
rect 421 386 422 387
rect 420 386 421 387
rect 419 386 420 387
rect 418 386 419 387
rect 417 386 418 387
rect 416 386 417 387
rect 415 386 416 387
rect 414 386 415 387
rect 413 386 414 387
rect 412 386 413 387
rect 411 386 412 387
rect 410 386 411 387
rect 409 386 410 387
rect 408 386 409 387
rect 407 386 408 387
rect 406 386 407 387
rect 405 386 406 387
rect 404 386 405 387
rect 403 386 404 387
rect 402 386 403 387
rect 401 386 402 387
rect 400 386 401 387
rect 399 386 400 387
rect 398 386 399 387
rect 397 386 398 387
rect 396 386 397 387
rect 395 386 396 387
rect 394 386 395 387
rect 393 386 394 387
rect 437 387 438 388
rect 436 387 437 388
rect 435 387 436 388
rect 434 387 435 388
rect 433 387 434 388
rect 432 387 433 388
rect 431 387 432 388
rect 430 387 431 388
rect 429 387 430 388
rect 428 387 429 388
rect 427 387 428 388
rect 426 387 427 388
rect 425 387 426 388
rect 424 387 425 388
rect 423 387 424 388
rect 422 387 423 388
rect 421 387 422 388
rect 420 387 421 388
rect 419 387 420 388
rect 418 387 419 388
rect 417 387 418 388
rect 416 387 417 388
rect 415 387 416 388
rect 414 387 415 388
rect 413 387 414 388
rect 412 387 413 388
rect 411 387 412 388
rect 410 387 411 388
rect 409 387 410 388
rect 408 387 409 388
rect 407 387 408 388
rect 406 387 407 388
rect 405 387 406 388
rect 404 387 405 388
rect 403 387 404 388
rect 402 387 403 388
rect 401 387 402 388
rect 400 387 401 388
rect 399 387 400 388
rect 398 387 399 388
rect 397 387 398 388
rect 396 387 397 388
rect 395 387 396 388
rect 394 387 395 388
rect 393 387 394 388
rect 437 388 438 389
rect 436 388 437 389
rect 435 388 436 389
rect 434 388 435 389
rect 433 388 434 389
rect 416 388 417 389
rect 415 388 416 389
rect 414 388 415 389
rect 413 388 414 389
rect 396 388 397 389
rect 395 388 396 389
rect 394 388 395 389
rect 393 388 394 389
rect 437 389 438 390
rect 436 389 437 390
rect 435 389 436 390
rect 434 389 435 390
rect 416 389 417 390
rect 415 389 416 390
rect 414 389 415 390
rect 413 389 414 390
rect 395 389 396 390
rect 394 389 395 390
rect 393 389 394 390
rect 437 390 438 391
rect 436 390 437 391
rect 435 390 436 391
rect 416 390 417 391
rect 415 390 416 391
rect 414 390 415 391
rect 413 390 414 391
rect 395 390 396 391
rect 394 390 395 391
rect 393 390 394 391
rect 437 391 438 392
rect 436 391 437 392
rect 435 391 436 392
rect 416 391 417 392
rect 415 391 416 392
rect 414 391 415 392
rect 413 391 414 392
rect 395 391 396 392
rect 394 391 395 392
rect 393 391 394 392
rect 437 392 438 393
rect 436 392 437 393
rect 435 392 436 393
rect 416 392 417 393
rect 415 392 416 393
rect 414 392 415 393
rect 413 392 414 393
rect 395 392 396 393
rect 394 392 395 393
rect 393 392 394 393
rect 437 393 438 394
rect 436 393 437 394
rect 435 393 436 394
rect 416 393 417 394
rect 415 393 416 394
rect 414 393 415 394
rect 413 393 414 394
rect 395 393 396 394
rect 394 393 395 394
rect 393 393 394 394
rect 437 394 438 395
rect 436 394 437 395
rect 435 394 436 395
rect 416 394 417 395
rect 415 394 416 395
rect 414 394 415 395
rect 413 394 414 395
rect 395 394 396 395
rect 394 394 395 395
rect 393 394 394 395
rect 437 395 438 396
rect 436 395 437 396
rect 435 395 436 396
rect 416 395 417 396
rect 415 395 416 396
rect 414 395 415 396
rect 413 395 414 396
rect 395 395 396 396
rect 394 395 395 396
rect 393 395 394 396
rect 437 396 438 397
rect 436 396 437 397
rect 435 396 436 397
rect 416 396 417 397
rect 415 396 416 397
rect 414 396 415 397
rect 413 396 414 397
rect 395 396 396 397
rect 394 396 395 397
rect 393 396 394 397
rect 437 397 438 398
rect 436 397 437 398
rect 435 397 436 398
rect 416 397 417 398
rect 415 397 416 398
rect 414 397 415 398
rect 413 397 414 398
rect 396 397 397 398
rect 395 397 396 398
rect 394 397 395 398
rect 393 397 394 398
rect 437 398 438 399
rect 436 398 437 399
rect 435 398 436 399
rect 417 398 418 399
rect 416 398 417 399
rect 415 398 416 399
rect 414 398 415 399
rect 413 398 414 399
rect 412 398 413 399
rect 396 398 397 399
rect 395 398 396 399
rect 394 398 395 399
rect 393 398 394 399
rect 437 399 438 400
rect 436 399 437 400
rect 435 399 436 400
rect 419 399 420 400
rect 418 399 419 400
rect 417 399 418 400
rect 416 399 417 400
rect 415 399 416 400
rect 414 399 415 400
rect 413 399 414 400
rect 412 399 413 400
rect 411 399 412 400
rect 410 399 411 400
rect 396 399 397 400
rect 395 399 396 400
rect 394 399 395 400
rect 393 399 394 400
rect 437 400 438 401
rect 436 400 437 401
rect 435 400 436 401
rect 434 400 435 401
rect 421 400 422 401
rect 420 400 421 401
rect 419 400 420 401
rect 418 400 419 401
rect 417 400 418 401
rect 416 400 417 401
rect 415 400 416 401
rect 414 400 415 401
rect 413 400 414 401
rect 412 400 413 401
rect 411 400 412 401
rect 410 400 411 401
rect 409 400 410 401
rect 408 400 409 401
rect 397 400 398 401
rect 396 400 397 401
rect 395 400 396 401
rect 394 400 395 401
rect 393 400 394 401
rect 437 401 438 402
rect 436 401 437 402
rect 435 401 436 402
rect 434 401 435 402
rect 421 401 422 402
rect 420 401 421 402
rect 419 401 420 402
rect 418 401 419 402
rect 417 401 418 402
rect 416 401 417 402
rect 415 401 416 402
rect 414 401 415 402
rect 413 401 414 402
rect 412 401 413 402
rect 411 401 412 402
rect 410 401 411 402
rect 409 401 410 402
rect 408 401 409 402
rect 398 401 399 402
rect 397 401 398 402
rect 396 401 397 402
rect 395 401 396 402
rect 394 401 395 402
rect 393 401 394 402
rect 437 402 438 403
rect 436 402 437 403
rect 435 402 436 403
rect 434 402 435 403
rect 433 402 434 403
rect 421 402 422 403
rect 420 402 421 403
rect 419 402 420 403
rect 418 402 419 403
rect 417 402 418 403
rect 416 402 417 403
rect 415 402 416 403
rect 414 402 415 403
rect 413 402 414 403
rect 412 402 413 403
rect 411 402 412 403
rect 410 402 411 403
rect 409 402 410 403
rect 408 402 409 403
rect 400 402 401 403
rect 399 402 400 403
rect 398 402 399 403
rect 397 402 398 403
rect 396 402 397 403
rect 395 402 396 403
rect 394 402 395 403
rect 393 402 394 403
rect 437 403 438 404
rect 436 403 437 404
rect 435 403 436 404
rect 434 403 435 404
rect 433 403 434 404
rect 432 403 433 404
rect 403 403 404 404
rect 402 403 403 404
rect 401 403 402 404
rect 400 403 401 404
rect 399 403 400 404
rect 398 403 399 404
rect 397 403 398 404
rect 396 403 397 404
rect 395 403 396 404
rect 394 403 395 404
rect 393 403 394 404
rect 437 404 438 405
rect 436 404 437 405
rect 435 404 436 405
rect 434 404 435 405
rect 433 404 434 405
rect 432 404 433 405
rect 431 404 432 405
rect 403 404 404 405
rect 402 404 403 405
rect 401 404 402 405
rect 400 404 401 405
rect 399 404 400 405
rect 398 404 399 405
rect 397 404 398 405
rect 396 404 397 405
rect 395 404 396 405
rect 394 404 395 405
rect 393 404 394 405
rect 437 405 438 406
rect 436 405 437 406
rect 435 405 436 406
rect 434 405 435 406
rect 433 405 434 406
rect 432 405 433 406
rect 431 405 432 406
rect 430 405 431 406
rect 429 405 430 406
rect 403 405 404 406
rect 402 405 403 406
rect 401 405 402 406
rect 400 405 401 406
rect 399 405 400 406
rect 398 405 399 406
rect 397 405 398 406
rect 396 405 397 406
rect 395 405 396 406
rect 394 405 395 406
rect 393 405 394 406
rect 437 406 438 407
rect 436 406 437 407
rect 435 406 436 407
rect 434 406 435 407
rect 433 406 434 407
rect 432 406 433 407
rect 431 406 432 407
rect 430 406 431 407
rect 429 406 430 407
rect 428 406 429 407
rect 427 406 428 407
rect 436 407 437 408
rect 435 407 436 408
rect 434 407 435 408
rect 433 407 434 408
rect 432 407 433 408
rect 431 407 432 408
rect 430 407 431 408
rect 429 407 430 408
rect 428 407 429 408
rect 427 407 428 408
rect 426 407 427 408
rect 432 408 433 409
rect 431 408 432 409
rect 430 408 431 409
rect 429 408 430 409
rect 428 408 429 409
rect 427 408 428 409
rect 426 408 427 409
rect 427 409 428 410
rect 426 409 427 410
<< metal2 >>
rect 439 2 440 3
rect 438 2 439 3
rect 397 2 398 3
rect 396 2 397 3
rect 395 2 396 3
rect 439 3 440 4
rect 438 3 439 4
rect 437 3 438 4
rect 397 3 398 4
rect 396 3 397 4
rect 395 3 396 4
rect 439 4 440 5
rect 438 4 439 5
rect 437 4 438 5
rect 397 4 398 5
rect 396 4 397 5
rect 395 4 396 5
rect 439 5 440 6
rect 438 5 439 6
rect 437 5 438 6
rect 397 5 398 6
rect 396 5 397 6
rect 395 5 396 6
rect 439 6 440 7
rect 438 6 439 7
rect 437 6 438 7
rect 398 6 399 7
rect 397 6 398 7
rect 396 6 397 7
rect 395 6 396 7
rect 439 7 440 8
rect 438 7 439 8
rect 437 7 438 8
rect 436 7 437 8
rect 435 7 436 8
rect 399 7 400 8
rect 398 7 399 8
rect 397 7 398 8
rect 396 7 397 8
rect 395 7 396 8
rect 439 8 440 9
rect 438 8 439 9
rect 437 8 438 9
rect 436 8 437 9
rect 435 8 436 9
rect 434 8 435 9
rect 433 8 434 9
rect 432 8 433 9
rect 431 8 432 9
rect 430 8 431 9
rect 429 8 430 9
rect 428 8 429 9
rect 427 8 428 9
rect 426 8 427 9
rect 425 8 426 9
rect 424 8 425 9
rect 423 8 424 9
rect 422 8 423 9
rect 421 8 422 9
rect 420 8 421 9
rect 419 8 420 9
rect 418 8 419 9
rect 417 8 418 9
rect 416 8 417 9
rect 415 8 416 9
rect 414 8 415 9
rect 413 8 414 9
rect 412 8 413 9
rect 411 8 412 9
rect 410 8 411 9
rect 409 8 410 9
rect 408 8 409 9
rect 407 8 408 9
rect 406 8 407 9
rect 405 8 406 9
rect 404 8 405 9
rect 403 8 404 9
rect 402 8 403 9
rect 401 8 402 9
rect 400 8 401 9
rect 399 8 400 9
rect 398 8 399 9
rect 397 8 398 9
rect 396 8 397 9
rect 395 8 396 9
rect 439 9 440 10
rect 438 9 439 10
rect 437 9 438 10
rect 436 9 437 10
rect 435 9 436 10
rect 434 9 435 10
rect 433 9 434 10
rect 432 9 433 10
rect 431 9 432 10
rect 430 9 431 10
rect 429 9 430 10
rect 428 9 429 10
rect 427 9 428 10
rect 426 9 427 10
rect 425 9 426 10
rect 424 9 425 10
rect 423 9 424 10
rect 422 9 423 10
rect 421 9 422 10
rect 420 9 421 10
rect 419 9 420 10
rect 418 9 419 10
rect 417 9 418 10
rect 416 9 417 10
rect 415 9 416 10
rect 414 9 415 10
rect 413 9 414 10
rect 412 9 413 10
rect 411 9 412 10
rect 410 9 411 10
rect 409 9 410 10
rect 408 9 409 10
rect 407 9 408 10
rect 406 9 407 10
rect 405 9 406 10
rect 404 9 405 10
rect 403 9 404 10
rect 402 9 403 10
rect 401 9 402 10
rect 400 9 401 10
rect 399 9 400 10
rect 398 9 399 10
rect 397 9 398 10
rect 396 9 397 10
rect 395 9 396 10
rect 439 10 440 11
rect 438 10 439 11
rect 437 10 438 11
rect 436 10 437 11
rect 435 10 436 11
rect 434 10 435 11
rect 433 10 434 11
rect 432 10 433 11
rect 431 10 432 11
rect 430 10 431 11
rect 429 10 430 11
rect 428 10 429 11
rect 427 10 428 11
rect 426 10 427 11
rect 425 10 426 11
rect 424 10 425 11
rect 423 10 424 11
rect 422 10 423 11
rect 421 10 422 11
rect 420 10 421 11
rect 419 10 420 11
rect 418 10 419 11
rect 417 10 418 11
rect 416 10 417 11
rect 415 10 416 11
rect 414 10 415 11
rect 413 10 414 11
rect 412 10 413 11
rect 411 10 412 11
rect 410 10 411 11
rect 409 10 410 11
rect 408 10 409 11
rect 407 10 408 11
rect 406 10 407 11
rect 405 10 406 11
rect 404 10 405 11
rect 403 10 404 11
rect 402 10 403 11
rect 401 10 402 11
rect 400 10 401 11
rect 399 10 400 11
rect 398 10 399 11
rect 397 10 398 11
rect 396 10 397 11
rect 395 10 396 11
rect 439 11 440 12
rect 438 11 439 12
rect 437 11 438 12
rect 436 11 437 12
rect 435 11 436 12
rect 434 11 435 12
rect 433 11 434 12
rect 432 11 433 12
rect 431 11 432 12
rect 430 11 431 12
rect 429 11 430 12
rect 428 11 429 12
rect 427 11 428 12
rect 426 11 427 12
rect 425 11 426 12
rect 424 11 425 12
rect 423 11 424 12
rect 422 11 423 12
rect 421 11 422 12
rect 420 11 421 12
rect 419 11 420 12
rect 418 11 419 12
rect 417 11 418 12
rect 416 11 417 12
rect 415 11 416 12
rect 414 11 415 12
rect 413 11 414 12
rect 412 11 413 12
rect 411 11 412 12
rect 410 11 411 12
rect 409 11 410 12
rect 408 11 409 12
rect 407 11 408 12
rect 406 11 407 12
rect 405 11 406 12
rect 404 11 405 12
rect 403 11 404 12
rect 402 11 403 12
rect 401 11 402 12
rect 400 11 401 12
rect 399 11 400 12
rect 398 11 399 12
rect 397 11 398 12
rect 396 11 397 12
rect 395 11 396 12
rect 439 12 440 13
rect 438 12 439 13
rect 437 12 438 13
rect 436 12 437 13
rect 435 12 436 13
rect 434 12 435 13
rect 433 12 434 13
rect 432 12 433 13
rect 431 12 432 13
rect 430 12 431 13
rect 429 12 430 13
rect 428 12 429 13
rect 427 12 428 13
rect 426 12 427 13
rect 425 12 426 13
rect 424 12 425 13
rect 423 12 424 13
rect 422 12 423 13
rect 421 12 422 13
rect 420 12 421 13
rect 419 12 420 13
rect 418 12 419 13
rect 417 12 418 13
rect 416 12 417 13
rect 415 12 416 13
rect 414 12 415 13
rect 413 12 414 13
rect 412 12 413 13
rect 411 12 412 13
rect 410 12 411 13
rect 409 12 410 13
rect 408 12 409 13
rect 407 12 408 13
rect 406 12 407 13
rect 405 12 406 13
rect 404 12 405 13
rect 403 12 404 13
rect 402 12 403 13
rect 401 12 402 13
rect 400 12 401 13
rect 399 12 400 13
rect 398 12 399 13
rect 397 12 398 13
rect 396 12 397 13
rect 395 12 396 13
rect 439 13 440 14
rect 438 13 439 14
rect 437 13 438 14
rect 436 13 437 14
rect 435 13 436 14
rect 434 13 435 14
rect 433 13 434 14
rect 432 13 433 14
rect 431 13 432 14
rect 430 13 431 14
rect 429 13 430 14
rect 428 13 429 14
rect 427 13 428 14
rect 426 13 427 14
rect 425 13 426 14
rect 424 13 425 14
rect 423 13 424 14
rect 422 13 423 14
rect 421 13 422 14
rect 420 13 421 14
rect 419 13 420 14
rect 418 13 419 14
rect 417 13 418 14
rect 416 13 417 14
rect 415 13 416 14
rect 414 13 415 14
rect 413 13 414 14
rect 412 13 413 14
rect 411 13 412 14
rect 410 13 411 14
rect 409 13 410 14
rect 408 13 409 14
rect 407 13 408 14
rect 406 13 407 14
rect 405 13 406 14
rect 404 13 405 14
rect 403 13 404 14
rect 402 13 403 14
rect 401 13 402 14
rect 400 13 401 14
rect 399 13 400 14
rect 398 13 399 14
rect 397 13 398 14
rect 396 13 397 14
rect 395 13 396 14
rect 439 14 440 15
rect 438 14 439 15
rect 437 14 438 15
rect 436 14 437 15
rect 435 14 436 15
rect 434 14 435 15
rect 433 14 434 15
rect 432 14 433 15
rect 431 14 432 15
rect 430 14 431 15
rect 429 14 430 15
rect 428 14 429 15
rect 427 14 428 15
rect 426 14 427 15
rect 425 14 426 15
rect 424 14 425 15
rect 423 14 424 15
rect 422 14 423 15
rect 421 14 422 15
rect 420 14 421 15
rect 419 14 420 15
rect 418 14 419 15
rect 417 14 418 15
rect 416 14 417 15
rect 415 14 416 15
rect 414 14 415 15
rect 413 14 414 15
rect 412 14 413 15
rect 411 14 412 15
rect 410 14 411 15
rect 409 14 410 15
rect 408 14 409 15
rect 407 14 408 15
rect 406 14 407 15
rect 405 14 406 15
rect 404 14 405 15
rect 403 14 404 15
rect 402 14 403 15
rect 401 14 402 15
rect 400 14 401 15
rect 399 14 400 15
rect 398 14 399 15
rect 397 14 398 15
rect 396 14 397 15
rect 395 14 396 15
rect 439 15 440 16
rect 438 15 439 16
rect 437 15 438 16
rect 436 15 437 16
rect 435 15 436 16
rect 434 15 435 16
rect 433 15 434 16
rect 432 15 433 16
rect 431 15 432 16
rect 430 15 431 16
rect 429 15 430 16
rect 428 15 429 16
rect 427 15 428 16
rect 426 15 427 16
rect 425 15 426 16
rect 424 15 425 16
rect 423 15 424 16
rect 422 15 423 16
rect 421 15 422 16
rect 420 15 421 16
rect 419 15 420 16
rect 418 15 419 16
rect 417 15 418 16
rect 416 15 417 16
rect 415 15 416 16
rect 414 15 415 16
rect 413 15 414 16
rect 412 15 413 16
rect 411 15 412 16
rect 410 15 411 16
rect 409 15 410 16
rect 408 15 409 16
rect 407 15 408 16
rect 406 15 407 16
rect 405 15 406 16
rect 404 15 405 16
rect 403 15 404 16
rect 402 15 403 16
rect 401 15 402 16
rect 400 15 401 16
rect 399 15 400 16
rect 398 15 399 16
rect 397 15 398 16
rect 396 15 397 16
rect 395 15 396 16
rect 439 16 440 17
rect 438 16 439 17
rect 437 16 438 17
rect 436 16 437 17
rect 435 16 436 17
rect 434 16 435 17
rect 433 16 434 17
rect 432 16 433 17
rect 431 16 432 17
rect 430 16 431 17
rect 429 16 430 17
rect 428 16 429 17
rect 427 16 428 17
rect 426 16 427 17
rect 425 16 426 17
rect 424 16 425 17
rect 423 16 424 17
rect 422 16 423 17
rect 421 16 422 17
rect 420 16 421 17
rect 419 16 420 17
rect 418 16 419 17
rect 417 16 418 17
rect 416 16 417 17
rect 415 16 416 17
rect 414 16 415 17
rect 413 16 414 17
rect 412 16 413 17
rect 411 16 412 17
rect 410 16 411 17
rect 409 16 410 17
rect 408 16 409 17
rect 407 16 408 17
rect 406 16 407 17
rect 405 16 406 17
rect 404 16 405 17
rect 403 16 404 17
rect 402 16 403 17
rect 401 16 402 17
rect 400 16 401 17
rect 399 16 400 17
rect 398 16 399 17
rect 397 16 398 17
rect 396 16 397 17
rect 395 16 396 17
rect 439 17 440 18
rect 438 17 439 18
rect 437 17 438 18
rect 436 17 437 18
rect 435 17 436 18
rect 418 17 419 18
rect 417 17 418 18
rect 416 17 417 18
rect 399 17 400 18
rect 398 17 399 18
rect 397 17 398 18
rect 396 17 397 18
rect 395 17 396 18
rect 439 18 440 19
rect 438 18 439 19
rect 437 18 438 19
rect 436 18 437 19
rect 418 18 419 19
rect 417 18 418 19
rect 416 18 417 19
rect 415 18 416 19
rect 398 18 399 19
rect 397 18 398 19
rect 396 18 397 19
rect 395 18 396 19
rect 439 19 440 20
rect 438 19 439 20
rect 437 19 438 20
rect 419 19 420 20
rect 418 19 419 20
rect 417 19 418 20
rect 416 19 417 20
rect 415 19 416 20
rect 397 19 398 20
rect 396 19 397 20
rect 395 19 396 20
rect 439 20 440 21
rect 438 20 439 21
rect 437 20 438 21
rect 420 20 421 21
rect 419 20 420 21
rect 418 20 419 21
rect 417 20 418 21
rect 416 20 417 21
rect 415 20 416 21
rect 414 20 415 21
rect 397 20 398 21
rect 396 20 397 21
rect 395 20 396 21
rect 439 21 440 22
rect 438 21 439 22
rect 437 21 438 22
rect 421 21 422 22
rect 420 21 421 22
rect 419 21 420 22
rect 418 21 419 22
rect 417 21 418 22
rect 416 21 417 22
rect 415 21 416 22
rect 414 21 415 22
rect 413 21 414 22
rect 397 21 398 22
rect 396 21 397 22
rect 395 21 396 22
rect 439 22 440 23
rect 438 22 439 23
rect 437 22 438 23
rect 423 22 424 23
rect 422 22 423 23
rect 421 22 422 23
rect 420 22 421 23
rect 419 22 420 23
rect 418 22 419 23
rect 417 22 418 23
rect 416 22 417 23
rect 415 22 416 23
rect 414 22 415 23
rect 413 22 414 23
rect 412 22 413 23
rect 397 22 398 23
rect 396 22 397 23
rect 395 22 396 23
rect 424 23 425 24
rect 423 23 424 24
rect 422 23 423 24
rect 421 23 422 24
rect 420 23 421 24
rect 419 23 420 24
rect 418 23 419 24
rect 417 23 418 24
rect 416 23 417 24
rect 415 23 416 24
rect 414 23 415 24
rect 413 23 414 24
rect 412 23 413 24
rect 411 23 412 24
rect 426 24 427 25
rect 425 24 426 25
rect 424 24 425 25
rect 423 24 424 25
rect 422 24 423 25
rect 421 24 422 25
rect 420 24 421 25
rect 419 24 420 25
rect 418 24 419 25
rect 417 24 418 25
rect 416 24 417 25
rect 415 24 416 25
rect 414 24 415 25
rect 413 24 414 25
rect 412 24 413 25
rect 411 24 412 25
rect 410 24 411 25
rect 427 25 428 26
rect 426 25 427 26
rect 425 25 426 26
rect 424 25 425 26
rect 423 25 424 26
rect 422 25 423 26
rect 421 25 422 26
rect 420 25 421 26
rect 419 25 420 26
rect 418 25 419 26
rect 417 25 418 26
rect 416 25 417 26
rect 415 25 416 26
rect 414 25 415 26
rect 413 25 414 26
rect 412 25 413 26
rect 411 25 412 26
rect 410 25 411 26
rect 409 25 410 26
rect 429 26 430 27
rect 428 26 429 27
rect 427 26 428 27
rect 426 26 427 27
rect 425 26 426 27
rect 424 26 425 27
rect 423 26 424 27
rect 422 26 423 27
rect 421 26 422 27
rect 420 26 421 27
rect 419 26 420 27
rect 418 26 419 27
rect 417 26 418 27
rect 416 26 417 27
rect 415 26 416 27
rect 414 26 415 27
rect 413 26 414 27
rect 411 26 412 27
rect 410 26 411 27
rect 409 26 410 27
rect 408 26 409 27
rect 430 27 431 28
rect 429 27 430 28
rect 428 27 429 28
rect 427 27 428 28
rect 426 27 427 28
rect 425 27 426 28
rect 424 27 425 28
rect 423 27 424 28
rect 422 27 423 28
rect 421 27 422 28
rect 420 27 421 28
rect 419 27 420 28
rect 418 27 419 28
rect 417 27 418 28
rect 416 27 417 28
rect 415 27 416 28
rect 410 27 411 28
rect 409 27 410 28
rect 408 27 409 28
rect 407 27 408 28
rect 431 28 432 29
rect 430 28 431 29
rect 429 28 430 29
rect 428 28 429 29
rect 427 28 428 29
rect 426 28 427 29
rect 425 28 426 29
rect 424 28 425 29
rect 423 28 424 29
rect 422 28 423 29
rect 421 28 422 29
rect 420 28 421 29
rect 419 28 420 29
rect 418 28 419 29
rect 417 28 418 29
rect 416 28 417 29
rect 409 28 410 29
rect 408 28 409 29
rect 407 28 408 29
rect 406 28 407 29
rect 433 29 434 30
rect 432 29 433 30
rect 431 29 432 30
rect 430 29 431 30
rect 429 29 430 30
rect 428 29 429 30
rect 427 29 428 30
rect 426 29 427 30
rect 425 29 426 30
rect 424 29 425 30
rect 423 29 424 30
rect 422 29 423 30
rect 421 29 422 30
rect 420 29 421 30
rect 419 29 420 30
rect 418 29 419 30
rect 417 29 418 30
rect 408 29 409 30
rect 407 29 408 30
rect 406 29 407 30
rect 405 29 406 30
rect 404 29 405 30
rect 397 29 398 30
rect 396 29 397 30
rect 395 29 396 30
rect 434 30 435 31
rect 433 30 434 31
rect 432 30 433 31
rect 431 30 432 31
rect 430 30 431 31
rect 429 30 430 31
rect 428 30 429 31
rect 427 30 428 31
rect 426 30 427 31
rect 425 30 426 31
rect 424 30 425 31
rect 423 30 424 31
rect 422 30 423 31
rect 421 30 422 31
rect 420 30 421 31
rect 419 30 420 31
rect 407 30 408 31
rect 406 30 407 31
rect 405 30 406 31
rect 404 30 405 31
rect 403 30 404 31
rect 397 30 398 31
rect 396 30 397 31
rect 395 30 396 31
rect 436 31 437 32
rect 435 31 436 32
rect 434 31 435 32
rect 433 31 434 32
rect 432 31 433 32
rect 431 31 432 32
rect 430 31 431 32
rect 429 31 430 32
rect 428 31 429 32
rect 427 31 428 32
rect 426 31 427 32
rect 425 31 426 32
rect 424 31 425 32
rect 423 31 424 32
rect 422 31 423 32
rect 421 31 422 32
rect 420 31 421 32
rect 406 31 407 32
rect 405 31 406 32
rect 404 31 405 32
rect 403 31 404 32
rect 402 31 403 32
rect 397 31 398 32
rect 396 31 397 32
rect 395 31 396 32
rect 437 32 438 33
rect 436 32 437 33
rect 435 32 436 33
rect 434 32 435 33
rect 433 32 434 33
rect 432 32 433 33
rect 431 32 432 33
rect 430 32 431 33
rect 429 32 430 33
rect 428 32 429 33
rect 427 32 428 33
rect 426 32 427 33
rect 425 32 426 33
rect 424 32 425 33
rect 423 32 424 33
rect 422 32 423 33
rect 405 32 406 33
rect 404 32 405 33
rect 403 32 404 33
rect 402 32 403 33
rect 401 32 402 33
rect 400 32 401 33
rect 397 32 398 33
rect 396 32 397 33
rect 395 32 396 33
rect 439 33 440 34
rect 438 33 439 34
rect 437 33 438 34
rect 436 33 437 34
rect 435 33 436 34
rect 434 33 435 34
rect 433 33 434 34
rect 432 33 433 34
rect 431 33 432 34
rect 430 33 431 34
rect 429 33 430 34
rect 428 33 429 34
rect 427 33 428 34
rect 426 33 427 34
rect 425 33 426 34
rect 424 33 425 34
rect 423 33 424 34
rect 404 33 405 34
rect 403 33 404 34
rect 402 33 403 34
rect 401 33 402 34
rect 400 33 401 34
rect 399 33 400 34
rect 398 33 399 34
rect 397 33 398 34
rect 396 33 397 34
rect 395 33 396 34
rect 439 34 440 35
rect 438 34 439 35
rect 437 34 438 35
rect 436 34 437 35
rect 435 34 436 35
rect 434 34 435 35
rect 433 34 434 35
rect 432 34 433 35
rect 431 34 432 35
rect 430 34 431 35
rect 429 34 430 35
rect 428 34 429 35
rect 427 34 428 35
rect 426 34 427 35
rect 425 34 426 35
rect 424 34 425 35
rect 403 34 404 35
rect 402 34 403 35
rect 401 34 402 35
rect 400 34 401 35
rect 399 34 400 35
rect 398 34 399 35
rect 397 34 398 35
rect 396 34 397 35
rect 395 34 396 35
rect 439 35 440 36
rect 438 35 439 36
rect 437 35 438 36
rect 436 35 437 36
rect 435 35 436 36
rect 434 35 435 36
rect 433 35 434 36
rect 432 35 433 36
rect 431 35 432 36
rect 430 35 431 36
rect 429 35 430 36
rect 428 35 429 36
rect 427 35 428 36
rect 426 35 427 36
rect 402 35 403 36
rect 401 35 402 36
rect 400 35 401 36
rect 399 35 400 36
rect 398 35 399 36
rect 397 35 398 36
rect 396 35 397 36
rect 395 35 396 36
rect 439 36 440 37
rect 438 36 439 37
rect 437 36 438 37
rect 436 36 437 37
rect 435 36 436 37
rect 434 36 435 37
rect 433 36 434 37
rect 432 36 433 37
rect 431 36 432 37
rect 430 36 431 37
rect 429 36 430 37
rect 428 36 429 37
rect 427 36 428 37
rect 401 36 402 37
rect 400 36 401 37
rect 399 36 400 37
rect 398 36 399 37
rect 397 36 398 37
rect 396 36 397 37
rect 395 36 396 37
rect 439 37 440 38
rect 438 37 439 38
rect 437 37 438 38
rect 436 37 437 38
rect 435 37 436 38
rect 434 37 435 38
rect 433 37 434 38
rect 432 37 433 38
rect 431 37 432 38
rect 430 37 431 38
rect 429 37 430 38
rect 428 37 429 38
rect 400 37 401 38
rect 399 37 400 38
rect 398 37 399 38
rect 397 37 398 38
rect 396 37 397 38
rect 395 37 396 38
rect 439 38 440 39
rect 438 38 439 39
rect 437 38 438 39
rect 436 38 437 39
rect 435 38 436 39
rect 434 38 435 39
rect 433 38 434 39
rect 432 38 433 39
rect 431 38 432 39
rect 430 38 431 39
rect 400 38 401 39
rect 399 38 400 39
rect 398 38 399 39
rect 397 38 398 39
rect 396 38 397 39
rect 395 38 396 39
rect 439 39 440 40
rect 438 39 439 40
rect 437 39 438 40
rect 436 39 437 40
rect 435 39 436 40
rect 434 39 435 40
rect 433 39 434 40
rect 432 39 433 40
rect 431 39 432 40
rect 399 39 400 40
rect 398 39 399 40
rect 397 39 398 40
rect 396 39 397 40
rect 395 39 396 40
rect 439 40 440 41
rect 438 40 439 41
rect 437 40 438 41
rect 436 40 437 41
rect 435 40 436 41
rect 434 40 435 41
rect 433 40 434 41
rect 432 40 433 41
rect 398 40 399 41
rect 397 40 398 41
rect 396 40 397 41
rect 395 40 396 41
rect 439 41 440 42
rect 438 41 439 42
rect 437 41 438 42
rect 436 41 437 42
rect 435 41 436 42
rect 434 41 435 42
rect 433 41 434 42
rect 398 41 399 42
rect 397 41 398 42
rect 396 41 397 42
rect 395 41 396 42
rect 439 42 440 43
rect 438 42 439 43
rect 437 42 438 43
rect 436 42 437 43
rect 435 42 436 43
rect 398 42 399 43
rect 397 42 398 43
rect 396 42 397 43
rect 395 42 396 43
rect 439 43 440 44
rect 438 43 439 44
rect 437 43 438 44
rect 436 43 437 44
rect 435 43 436 44
rect 397 43 398 44
rect 396 43 397 44
rect 395 43 396 44
rect 439 44 440 45
rect 438 44 439 45
rect 437 44 438 45
rect 436 44 437 45
rect 397 44 398 45
rect 396 44 397 45
rect 395 44 396 45
rect 439 45 440 46
rect 438 45 439 46
rect 437 45 438 46
rect 397 45 398 46
rect 396 45 397 46
rect 395 45 396 46
rect 439 46 440 47
rect 438 46 439 47
rect 437 46 438 47
rect 397 46 398 47
rect 396 46 397 47
rect 395 46 396 47
rect 439 47 440 48
rect 438 47 439 48
rect 437 47 438 48
rect 91 49 92 50
rect 90 49 91 50
rect 89 49 90 50
rect 88 49 89 50
rect 87 49 88 50
rect 86 49 87 50
rect 93 50 94 51
rect 92 50 93 51
rect 91 50 92 51
rect 90 50 91 51
rect 89 50 90 51
rect 88 50 89 51
rect 87 50 88 51
rect 86 50 87 51
rect 85 50 86 51
rect 84 50 85 51
rect 94 51 95 52
rect 93 51 94 52
rect 92 51 93 52
rect 91 51 92 52
rect 90 51 91 52
rect 89 51 90 52
rect 88 51 89 52
rect 87 51 88 52
rect 86 51 87 52
rect 85 51 86 52
rect 84 51 85 52
rect 83 51 84 52
rect 396 52 397 53
rect 395 52 396 53
rect 94 52 95 53
rect 93 52 94 53
rect 92 52 93 53
rect 91 52 92 53
rect 90 52 91 53
rect 89 52 90 53
rect 88 52 89 53
rect 87 52 88 53
rect 86 52 87 53
rect 85 52 86 53
rect 84 52 85 53
rect 83 52 84 53
rect 82 52 83 53
rect 397 53 398 54
rect 396 53 397 54
rect 395 53 396 54
rect 95 53 96 54
rect 94 53 95 54
rect 93 53 94 54
rect 92 53 93 54
rect 91 53 92 54
rect 90 53 91 54
rect 89 53 90 54
rect 88 53 89 54
rect 87 53 88 54
rect 86 53 87 54
rect 85 53 86 54
rect 84 53 85 54
rect 83 53 84 54
rect 82 53 83 54
rect 81 53 82 54
rect 397 54 398 55
rect 396 54 397 55
rect 395 54 396 55
rect 95 54 96 55
rect 94 54 95 55
rect 93 54 94 55
rect 92 54 93 55
rect 91 54 92 55
rect 90 54 91 55
rect 89 54 90 55
rect 88 54 89 55
rect 87 54 88 55
rect 86 54 87 55
rect 85 54 86 55
rect 84 54 85 55
rect 83 54 84 55
rect 82 54 83 55
rect 81 54 82 55
rect 80 54 81 55
rect 397 55 398 56
rect 396 55 397 56
rect 395 55 396 56
rect 95 55 96 56
rect 94 55 95 56
rect 93 55 94 56
rect 92 55 93 56
rect 91 55 92 56
rect 90 55 91 56
rect 89 55 90 56
rect 88 55 89 56
rect 87 55 88 56
rect 86 55 87 56
rect 85 55 86 56
rect 84 55 85 56
rect 83 55 84 56
rect 82 55 83 56
rect 81 55 82 56
rect 80 55 81 56
rect 79 55 80 56
rect 398 56 399 57
rect 397 56 398 57
rect 396 56 397 57
rect 395 56 396 57
rect 107 56 108 57
rect 94 56 95 57
rect 93 56 94 57
rect 92 56 93 57
rect 91 56 92 57
rect 90 56 91 57
rect 89 56 90 57
rect 88 56 89 57
rect 87 56 88 57
rect 86 56 87 57
rect 85 56 86 57
rect 84 56 85 57
rect 83 56 84 57
rect 82 56 83 57
rect 81 56 82 57
rect 80 56 81 57
rect 79 56 80 57
rect 78 56 79 57
rect 399 57 400 58
rect 398 57 399 58
rect 397 57 398 58
rect 396 57 397 58
rect 395 57 396 58
rect 110 57 111 58
rect 109 57 110 58
rect 108 57 109 58
rect 107 57 108 58
rect 106 57 107 58
rect 105 57 106 58
rect 104 57 105 58
rect 94 57 95 58
rect 93 57 94 58
rect 92 57 93 58
rect 91 57 92 58
rect 90 57 91 58
rect 89 57 90 58
rect 88 57 89 58
rect 87 57 88 58
rect 86 57 87 58
rect 85 57 86 58
rect 84 57 85 58
rect 83 57 84 58
rect 82 57 83 58
rect 81 57 82 58
rect 80 57 81 58
rect 79 57 80 58
rect 78 57 79 58
rect 400 58 401 59
rect 399 58 400 59
rect 398 58 399 59
rect 397 58 398 59
rect 396 58 397 59
rect 395 58 396 59
rect 112 58 113 59
rect 111 58 112 59
rect 110 58 111 59
rect 109 58 110 59
rect 108 58 109 59
rect 107 58 108 59
rect 106 58 107 59
rect 105 58 106 59
rect 104 58 105 59
rect 103 58 104 59
rect 102 58 103 59
rect 94 58 95 59
rect 93 58 94 59
rect 92 58 93 59
rect 91 58 92 59
rect 90 58 91 59
rect 89 58 90 59
rect 88 58 89 59
rect 87 58 88 59
rect 86 58 87 59
rect 85 58 86 59
rect 84 58 85 59
rect 83 58 84 59
rect 82 58 83 59
rect 81 58 82 59
rect 80 58 81 59
rect 79 58 80 59
rect 78 58 79 59
rect 77 58 78 59
rect 402 59 403 60
rect 401 59 402 60
rect 400 59 401 60
rect 399 59 400 60
rect 398 59 399 60
rect 397 59 398 60
rect 396 59 397 60
rect 395 59 396 60
rect 114 59 115 60
rect 113 59 114 60
rect 112 59 113 60
rect 111 59 112 60
rect 110 59 111 60
rect 109 59 110 60
rect 108 59 109 60
rect 107 59 108 60
rect 106 59 107 60
rect 105 59 106 60
rect 104 59 105 60
rect 103 59 104 60
rect 102 59 103 60
rect 101 59 102 60
rect 94 59 95 60
rect 93 59 94 60
rect 92 59 93 60
rect 91 59 92 60
rect 90 59 91 60
rect 89 59 90 60
rect 88 59 89 60
rect 87 59 88 60
rect 86 59 87 60
rect 85 59 86 60
rect 84 59 85 60
rect 83 59 84 60
rect 82 59 83 60
rect 81 59 82 60
rect 80 59 81 60
rect 79 59 80 60
rect 78 59 79 60
rect 77 59 78 60
rect 76 59 77 60
rect 404 60 405 61
rect 403 60 404 61
rect 402 60 403 61
rect 401 60 402 61
rect 400 60 401 61
rect 399 60 400 61
rect 398 60 399 61
rect 397 60 398 61
rect 396 60 397 61
rect 395 60 396 61
rect 116 60 117 61
rect 115 60 116 61
rect 114 60 115 61
rect 113 60 114 61
rect 112 60 113 61
rect 111 60 112 61
rect 110 60 111 61
rect 109 60 110 61
rect 108 60 109 61
rect 107 60 108 61
rect 106 60 107 61
rect 105 60 106 61
rect 104 60 105 61
rect 103 60 104 61
rect 102 60 103 61
rect 101 60 102 61
rect 100 60 101 61
rect 93 60 94 61
rect 92 60 93 61
rect 91 60 92 61
rect 90 60 91 61
rect 89 60 90 61
rect 88 60 89 61
rect 87 60 88 61
rect 86 60 87 61
rect 85 60 86 61
rect 84 60 85 61
rect 83 60 84 61
rect 82 60 83 61
rect 81 60 82 61
rect 80 60 81 61
rect 79 60 80 61
rect 78 60 79 61
rect 77 60 78 61
rect 76 60 77 61
rect 405 61 406 62
rect 404 61 405 62
rect 403 61 404 62
rect 402 61 403 62
rect 401 61 402 62
rect 400 61 401 62
rect 399 61 400 62
rect 398 61 399 62
rect 397 61 398 62
rect 396 61 397 62
rect 395 61 396 62
rect 117 61 118 62
rect 116 61 117 62
rect 115 61 116 62
rect 114 61 115 62
rect 113 61 114 62
rect 112 61 113 62
rect 111 61 112 62
rect 110 61 111 62
rect 109 61 110 62
rect 108 61 109 62
rect 107 61 108 62
rect 106 61 107 62
rect 105 61 106 62
rect 104 61 105 62
rect 103 61 104 62
rect 102 61 103 62
rect 101 61 102 62
rect 100 61 101 62
rect 99 61 100 62
rect 93 61 94 62
rect 92 61 93 62
rect 91 61 92 62
rect 90 61 91 62
rect 89 61 90 62
rect 88 61 89 62
rect 87 61 88 62
rect 86 61 87 62
rect 85 61 86 62
rect 84 61 85 62
rect 83 61 84 62
rect 82 61 83 62
rect 81 61 82 62
rect 80 61 81 62
rect 79 61 80 62
rect 78 61 79 62
rect 77 61 78 62
rect 76 61 77 62
rect 75 61 76 62
rect 407 62 408 63
rect 406 62 407 63
rect 405 62 406 63
rect 404 62 405 63
rect 403 62 404 63
rect 402 62 403 63
rect 401 62 402 63
rect 400 62 401 63
rect 399 62 400 63
rect 398 62 399 63
rect 397 62 398 63
rect 396 62 397 63
rect 395 62 396 63
rect 118 62 119 63
rect 117 62 118 63
rect 116 62 117 63
rect 115 62 116 63
rect 114 62 115 63
rect 113 62 114 63
rect 112 62 113 63
rect 111 62 112 63
rect 110 62 111 63
rect 109 62 110 63
rect 108 62 109 63
rect 107 62 108 63
rect 106 62 107 63
rect 105 62 106 63
rect 104 62 105 63
rect 103 62 104 63
rect 102 62 103 63
rect 101 62 102 63
rect 100 62 101 63
rect 99 62 100 63
rect 98 62 99 63
rect 93 62 94 63
rect 92 62 93 63
rect 91 62 92 63
rect 90 62 91 63
rect 89 62 90 63
rect 88 62 89 63
rect 87 62 88 63
rect 86 62 87 63
rect 85 62 86 63
rect 84 62 85 63
rect 83 62 84 63
rect 82 62 83 63
rect 81 62 82 63
rect 80 62 81 63
rect 79 62 80 63
rect 78 62 79 63
rect 77 62 78 63
rect 76 62 77 63
rect 75 62 76 63
rect 439 63 440 64
rect 438 63 439 64
rect 409 63 410 64
rect 408 63 409 64
rect 407 63 408 64
rect 406 63 407 64
rect 405 63 406 64
rect 404 63 405 64
rect 403 63 404 64
rect 402 63 403 64
rect 401 63 402 64
rect 400 63 401 64
rect 399 63 400 64
rect 398 63 399 64
rect 397 63 398 64
rect 396 63 397 64
rect 395 63 396 64
rect 119 63 120 64
rect 118 63 119 64
rect 117 63 118 64
rect 116 63 117 64
rect 115 63 116 64
rect 114 63 115 64
rect 113 63 114 64
rect 112 63 113 64
rect 111 63 112 64
rect 110 63 111 64
rect 109 63 110 64
rect 108 63 109 64
rect 107 63 108 64
rect 106 63 107 64
rect 105 63 106 64
rect 104 63 105 64
rect 103 63 104 64
rect 102 63 103 64
rect 101 63 102 64
rect 100 63 101 64
rect 99 63 100 64
rect 98 63 99 64
rect 97 63 98 64
rect 92 63 93 64
rect 91 63 92 64
rect 90 63 91 64
rect 89 63 90 64
rect 88 63 89 64
rect 87 63 88 64
rect 86 63 87 64
rect 85 63 86 64
rect 84 63 85 64
rect 83 63 84 64
rect 82 63 83 64
rect 81 63 82 64
rect 80 63 81 64
rect 79 63 80 64
rect 78 63 79 64
rect 77 63 78 64
rect 76 63 77 64
rect 75 63 76 64
rect 74 63 75 64
rect 439 64 440 65
rect 438 64 439 65
rect 437 64 438 65
rect 411 64 412 65
rect 410 64 411 65
rect 409 64 410 65
rect 408 64 409 65
rect 407 64 408 65
rect 406 64 407 65
rect 405 64 406 65
rect 404 64 405 65
rect 403 64 404 65
rect 402 64 403 65
rect 401 64 402 65
rect 400 64 401 65
rect 399 64 400 65
rect 398 64 399 65
rect 397 64 398 65
rect 396 64 397 65
rect 395 64 396 65
rect 120 64 121 65
rect 119 64 120 65
rect 118 64 119 65
rect 117 64 118 65
rect 116 64 117 65
rect 115 64 116 65
rect 114 64 115 65
rect 113 64 114 65
rect 112 64 113 65
rect 111 64 112 65
rect 110 64 111 65
rect 109 64 110 65
rect 108 64 109 65
rect 107 64 108 65
rect 106 64 107 65
rect 105 64 106 65
rect 104 64 105 65
rect 103 64 104 65
rect 102 64 103 65
rect 101 64 102 65
rect 100 64 101 65
rect 99 64 100 65
rect 98 64 99 65
rect 97 64 98 65
rect 96 64 97 65
rect 92 64 93 65
rect 91 64 92 65
rect 90 64 91 65
rect 89 64 90 65
rect 88 64 89 65
rect 87 64 88 65
rect 86 64 87 65
rect 85 64 86 65
rect 84 64 85 65
rect 83 64 84 65
rect 82 64 83 65
rect 81 64 82 65
rect 80 64 81 65
rect 79 64 80 65
rect 78 64 79 65
rect 77 64 78 65
rect 76 64 77 65
rect 75 64 76 65
rect 74 64 75 65
rect 73 64 74 65
rect 439 65 440 66
rect 438 65 439 66
rect 437 65 438 66
rect 412 65 413 66
rect 411 65 412 66
rect 410 65 411 66
rect 409 65 410 66
rect 408 65 409 66
rect 407 65 408 66
rect 406 65 407 66
rect 405 65 406 66
rect 404 65 405 66
rect 403 65 404 66
rect 402 65 403 66
rect 401 65 402 66
rect 400 65 401 66
rect 399 65 400 66
rect 398 65 399 66
rect 397 65 398 66
rect 396 65 397 66
rect 395 65 396 66
rect 121 65 122 66
rect 120 65 121 66
rect 119 65 120 66
rect 118 65 119 66
rect 117 65 118 66
rect 116 65 117 66
rect 115 65 116 66
rect 114 65 115 66
rect 113 65 114 66
rect 112 65 113 66
rect 111 65 112 66
rect 110 65 111 66
rect 109 65 110 66
rect 108 65 109 66
rect 107 65 108 66
rect 106 65 107 66
rect 105 65 106 66
rect 104 65 105 66
rect 103 65 104 66
rect 102 65 103 66
rect 101 65 102 66
rect 100 65 101 66
rect 99 65 100 66
rect 98 65 99 66
rect 97 65 98 66
rect 96 65 97 66
rect 95 65 96 66
rect 91 65 92 66
rect 90 65 91 66
rect 89 65 90 66
rect 88 65 89 66
rect 87 65 88 66
rect 86 65 87 66
rect 85 65 86 66
rect 84 65 85 66
rect 83 65 84 66
rect 82 65 83 66
rect 81 65 82 66
rect 80 65 81 66
rect 79 65 80 66
rect 78 65 79 66
rect 77 65 78 66
rect 76 65 77 66
rect 75 65 76 66
rect 74 65 75 66
rect 73 65 74 66
rect 439 66 440 67
rect 438 66 439 67
rect 437 66 438 67
rect 414 66 415 67
rect 413 66 414 67
rect 412 66 413 67
rect 411 66 412 67
rect 410 66 411 67
rect 409 66 410 67
rect 408 66 409 67
rect 407 66 408 67
rect 406 66 407 67
rect 405 66 406 67
rect 404 66 405 67
rect 403 66 404 67
rect 402 66 403 67
rect 401 66 402 67
rect 400 66 401 67
rect 399 66 400 67
rect 398 66 399 67
rect 397 66 398 67
rect 396 66 397 67
rect 395 66 396 67
rect 122 66 123 67
rect 121 66 122 67
rect 120 66 121 67
rect 119 66 120 67
rect 118 66 119 67
rect 117 66 118 67
rect 116 66 117 67
rect 115 66 116 67
rect 114 66 115 67
rect 113 66 114 67
rect 112 66 113 67
rect 111 66 112 67
rect 110 66 111 67
rect 109 66 110 67
rect 108 66 109 67
rect 107 66 108 67
rect 106 66 107 67
rect 105 66 106 67
rect 104 66 105 67
rect 103 66 104 67
rect 102 66 103 67
rect 101 66 102 67
rect 100 66 101 67
rect 99 66 100 67
rect 98 66 99 67
rect 97 66 98 67
rect 96 66 97 67
rect 95 66 96 67
rect 94 66 95 67
rect 91 66 92 67
rect 90 66 91 67
rect 89 66 90 67
rect 88 66 89 67
rect 87 66 88 67
rect 86 66 87 67
rect 85 66 86 67
rect 84 66 85 67
rect 83 66 84 67
rect 82 66 83 67
rect 81 66 82 67
rect 80 66 81 67
rect 79 66 80 67
rect 78 66 79 67
rect 77 66 78 67
rect 76 66 77 67
rect 75 66 76 67
rect 74 66 75 67
rect 73 66 74 67
rect 72 66 73 67
rect 439 67 440 68
rect 438 67 439 68
rect 437 67 438 68
rect 416 67 417 68
rect 415 67 416 68
rect 414 67 415 68
rect 413 67 414 68
rect 412 67 413 68
rect 411 67 412 68
rect 410 67 411 68
rect 409 67 410 68
rect 408 67 409 68
rect 407 67 408 68
rect 406 67 407 68
rect 405 67 406 68
rect 404 67 405 68
rect 403 67 404 68
rect 402 67 403 68
rect 401 67 402 68
rect 400 67 401 68
rect 399 67 400 68
rect 398 67 399 68
rect 397 67 398 68
rect 396 67 397 68
rect 395 67 396 68
rect 123 67 124 68
rect 122 67 123 68
rect 121 67 122 68
rect 120 67 121 68
rect 119 67 120 68
rect 118 67 119 68
rect 117 67 118 68
rect 116 67 117 68
rect 115 67 116 68
rect 114 67 115 68
rect 113 67 114 68
rect 112 67 113 68
rect 111 67 112 68
rect 110 67 111 68
rect 109 67 110 68
rect 108 67 109 68
rect 107 67 108 68
rect 106 67 107 68
rect 105 67 106 68
rect 104 67 105 68
rect 103 67 104 68
rect 102 67 103 68
rect 101 67 102 68
rect 100 67 101 68
rect 99 67 100 68
rect 98 67 99 68
rect 97 67 98 68
rect 96 67 97 68
rect 95 67 96 68
rect 94 67 95 68
rect 93 67 94 68
rect 90 67 91 68
rect 89 67 90 68
rect 88 67 89 68
rect 87 67 88 68
rect 86 67 87 68
rect 85 67 86 68
rect 84 67 85 68
rect 83 67 84 68
rect 82 67 83 68
rect 81 67 82 68
rect 80 67 81 68
rect 79 67 80 68
rect 78 67 79 68
rect 77 67 78 68
rect 76 67 77 68
rect 75 67 76 68
rect 74 67 75 68
rect 73 67 74 68
rect 72 67 73 68
rect 439 68 440 69
rect 438 68 439 69
rect 437 68 438 69
rect 436 68 437 69
rect 418 68 419 69
rect 417 68 418 69
rect 416 68 417 69
rect 415 68 416 69
rect 414 68 415 69
rect 413 68 414 69
rect 412 68 413 69
rect 411 68 412 69
rect 410 68 411 69
rect 409 68 410 69
rect 408 68 409 69
rect 407 68 408 69
rect 406 68 407 69
rect 405 68 406 69
rect 404 68 405 69
rect 403 68 404 69
rect 402 68 403 69
rect 401 68 402 69
rect 400 68 401 69
rect 398 68 399 69
rect 397 68 398 69
rect 396 68 397 69
rect 395 68 396 69
rect 123 68 124 69
rect 122 68 123 69
rect 121 68 122 69
rect 120 68 121 69
rect 119 68 120 69
rect 118 68 119 69
rect 117 68 118 69
rect 116 68 117 69
rect 115 68 116 69
rect 114 68 115 69
rect 113 68 114 69
rect 112 68 113 69
rect 111 68 112 69
rect 110 68 111 69
rect 109 68 110 69
rect 108 68 109 69
rect 107 68 108 69
rect 106 68 107 69
rect 105 68 106 69
rect 104 68 105 69
rect 103 68 104 69
rect 102 68 103 69
rect 101 68 102 69
rect 100 68 101 69
rect 99 68 100 69
rect 98 68 99 69
rect 97 68 98 69
rect 96 68 97 69
rect 95 68 96 69
rect 94 68 95 69
rect 93 68 94 69
rect 92 68 93 69
rect 90 68 91 69
rect 89 68 90 69
rect 88 68 89 69
rect 87 68 88 69
rect 86 68 87 69
rect 85 68 86 69
rect 84 68 85 69
rect 83 68 84 69
rect 82 68 83 69
rect 81 68 82 69
rect 80 68 81 69
rect 79 68 80 69
rect 78 68 79 69
rect 77 68 78 69
rect 76 68 77 69
rect 75 68 76 69
rect 74 68 75 69
rect 73 68 74 69
rect 72 68 73 69
rect 439 69 440 70
rect 438 69 439 70
rect 437 69 438 70
rect 436 69 437 70
rect 435 69 436 70
rect 434 69 435 70
rect 433 69 434 70
rect 432 69 433 70
rect 431 69 432 70
rect 430 69 431 70
rect 429 69 430 70
rect 428 69 429 70
rect 427 69 428 70
rect 426 69 427 70
rect 425 69 426 70
rect 424 69 425 70
rect 423 69 424 70
rect 422 69 423 70
rect 421 69 422 70
rect 420 69 421 70
rect 419 69 420 70
rect 418 69 419 70
rect 417 69 418 70
rect 416 69 417 70
rect 415 69 416 70
rect 414 69 415 70
rect 413 69 414 70
rect 412 69 413 70
rect 411 69 412 70
rect 410 69 411 70
rect 409 69 410 70
rect 408 69 409 70
rect 407 69 408 70
rect 406 69 407 70
rect 405 69 406 70
rect 404 69 405 70
rect 403 69 404 70
rect 402 69 403 70
rect 397 69 398 70
rect 396 69 397 70
rect 395 69 396 70
rect 124 69 125 70
rect 123 69 124 70
rect 122 69 123 70
rect 121 69 122 70
rect 120 69 121 70
rect 119 69 120 70
rect 118 69 119 70
rect 117 69 118 70
rect 116 69 117 70
rect 115 69 116 70
rect 114 69 115 70
rect 113 69 114 70
rect 112 69 113 70
rect 111 69 112 70
rect 110 69 111 70
rect 109 69 110 70
rect 108 69 109 70
rect 107 69 108 70
rect 106 69 107 70
rect 105 69 106 70
rect 104 69 105 70
rect 103 69 104 70
rect 102 69 103 70
rect 101 69 102 70
rect 100 69 101 70
rect 99 69 100 70
rect 98 69 99 70
rect 97 69 98 70
rect 96 69 97 70
rect 95 69 96 70
rect 94 69 95 70
rect 93 69 94 70
rect 92 69 93 70
rect 91 69 92 70
rect 89 69 90 70
rect 88 69 89 70
rect 87 69 88 70
rect 86 69 87 70
rect 85 69 86 70
rect 84 69 85 70
rect 83 69 84 70
rect 82 69 83 70
rect 81 69 82 70
rect 80 69 81 70
rect 79 69 80 70
rect 78 69 79 70
rect 77 69 78 70
rect 76 69 77 70
rect 75 69 76 70
rect 74 69 75 70
rect 73 69 74 70
rect 72 69 73 70
rect 71 69 72 70
rect 439 70 440 71
rect 438 70 439 71
rect 437 70 438 71
rect 436 70 437 71
rect 435 70 436 71
rect 434 70 435 71
rect 433 70 434 71
rect 432 70 433 71
rect 431 70 432 71
rect 430 70 431 71
rect 429 70 430 71
rect 428 70 429 71
rect 427 70 428 71
rect 426 70 427 71
rect 425 70 426 71
rect 424 70 425 71
rect 423 70 424 71
rect 422 70 423 71
rect 421 70 422 71
rect 420 70 421 71
rect 419 70 420 71
rect 418 70 419 71
rect 417 70 418 71
rect 416 70 417 71
rect 415 70 416 71
rect 414 70 415 71
rect 413 70 414 71
rect 412 70 413 71
rect 411 70 412 71
rect 410 70 411 71
rect 409 70 410 71
rect 408 70 409 71
rect 407 70 408 71
rect 406 70 407 71
rect 405 70 406 71
rect 404 70 405 71
rect 397 70 398 71
rect 396 70 397 71
rect 395 70 396 71
rect 124 70 125 71
rect 123 70 124 71
rect 122 70 123 71
rect 121 70 122 71
rect 120 70 121 71
rect 119 70 120 71
rect 118 70 119 71
rect 117 70 118 71
rect 116 70 117 71
rect 115 70 116 71
rect 114 70 115 71
rect 113 70 114 71
rect 112 70 113 71
rect 111 70 112 71
rect 110 70 111 71
rect 109 70 110 71
rect 108 70 109 71
rect 107 70 108 71
rect 106 70 107 71
rect 105 70 106 71
rect 104 70 105 71
rect 103 70 104 71
rect 102 70 103 71
rect 101 70 102 71
rect 100 70 101 71
rect 99 70 100 71
rect 98 70 99 71
rect 97 70 98 71
rect 96 70 97 71
rect 95 70 96 71
rect 94 70 95 71
rect 93 70 94 71
rect 92 70 93 71
rect 91 70 92 71
rect 90 70 91 71
rect 89 70 90 71
rect 88 70 89 71
rect 87 70 88 71
rect 86 70 87 71
rect 85 70 86 71
rect 84 70 85 71
rect 83 70 84 71
rect 82 70 83 71
rect 81 70 82 71
rect 80 70 81 71
rect 79 70 80 71
rect 78 70 79 71
rect 77 70 78 71
rect 76 70 77 71
rect 75 70 76 71
rect 74 70 75 71
rect 73 70 74 71
rect 72 70 73 71
rect 71 70 72 71
rect 439 71 440 72
rect 438 71 439 72
rect 437 71 438 72
rect 436 71 437 72
rect 435 71 436 72
rect 434 71 435 72
rect 433 71 434 72
rect 432 71 433 72
rect 431 71 432 72
rect 430 71 431 72
rect 429 71 430 72
rect 428 71 429 72
rect 427 71 428 72
rect 426 71 427 72
rect 425 71 426 72
rect 424 71 425 72
rect 423 71 424 72
rect 422 71 423 72
rect 421 71 422 72
rect 420 71 421 72
rect 419 71 420 72
rect 418 71 419 72
rect 417 71 418 72
rect 416 71 417 72
rect 415 71 416 72
rect 414 71 415 72
rect 413 71 414 72
rect 412 71 413 72
rect 411 71 412 72
rect 410 71 411 72
rect 409 71 410 72
rect 408 71 409 72
rect 407 71 408 72
rect 406 71 407 72
rect 397 71 398 72
rect 396 71 397 72
rect 395 71 396 72
rect 139 71 140 72
rect 138 71 139 72
rect 137 71 138 72
rect 136 71 137 72
rect 135 71 136 72
rect 134 71 135 72
rect 124 71 125 72
rect 123 71 124 72
rect 122 71 123 72
rect 121 71 122 72
rect 120 71 121 72
rect 119 71 120 72
rect 118 71 119 72
rect 117 71 118 72
rect 116 71 117 72
rect 115 71 116 72
rect 114 71 115 72
rect 113 71 114 72
rect 112 71 113 72
rect 111 71 112 72
rect 110 71 111 72
rect 109 71 110 72
rect 108 71 109 72
rect 107 71 108 72
rect 106 71 107 72
rect 105 71 106 72
rect 104 71 105 72
rect 103 71 104 72
rect 102 71 103 72
rect 101 71 102 72
rect 100 71 101 72
rect 99 71 100 72
rect 98 71 99 72
rect 97 71 98 72
rect 96 71 97 72
rect 95 71 96 72
rect 94 71 95 72
rect 93 71 94 72
rect 92 71 93 72
rect 91 71 92 72
rect 90 71 91 72
rect 89 71 90 72
rect 88 71 89 72
rect 87 71 88 72
rect 86 71 87 72
rect 85 71 86 72
rect 84 71 85 72
rect 83 71 84 72
rect 82 71 83 72
rect 81 71 82 72
rect 80 71 81 72
rect 79 71 80 72
rect 78 71 79 72
rect 77 71 78 72
rect 76 71 77 72
rect 75 71 76 72
rect 74 71 75 72
rect 73 71 74 72
rect 72 71 73 72
rect 71 71 72 72
rect 70 71 71 72
rect 439 72 440 73
rect 438 72 439 73
rect 437 72 438 73
rect 436 72 437 73
rect 435 72 436 73
rect 434 72 435 73
rect 433 72 434 73
rect 432 72 433 73
rect 431 72 432 73
rect 430 72 431 73
rect 429 72 430 73
rect 428 72 429 73
rect 427 72 428 73
rect 426 72 427 73
rect 425 72 426 73
rect 424 72 425 73
rect 423 72 424 73
rect 422 72 423 73
rect 421 72 422 73
rect 420 72 421 73
rect 419 72 420 73
rect 418 72 419 73
rect 417 72 418 73
rect 416 72 417 73
rect 415 72 416 73
rect 414 72 415 73
rect 413 72 414 73
rect 412 72 413 73
rect 411 72 412 73
rect 410 72 411 73
rect 409 72 410 73
rect 408 72 409 73
rect 142 72 143 73
rect 141 72 142 73
rect 140 72 141 73
rect 139 72 140 73
rect 138 72 139 73
rect 137 72 138 73
rect 136 72 137 73
rect 135 72 136 73
rect 134 72 135 73
rect 133 72 134 73
rect 132 72 133 73
rect 124 72 125 73
rect 123 72 124 73
rect 122 72 123 73
rect 121 72 122 73
rect 120 72 121 73
rect 119 72 120 73
rect 118 72 119 73
rect 117 72 118 73
rect 116 72 117 73
rect 115 72 116 73
rect 114 72 115 73
rect 113 72 114 73
rect 112 72 113 73
rect 111 72 112 73
rect 110 72 111 73
rect 109 72 110 73
rect 108 72 109 73
rect 107 72 108 73
rect 106 72 107 73
rect 105 72 106 73
rect 104 72 105 73
rect 103 72 104 73
rect 102 72 103 73
rect 101 72 102 73
rect 100 72 101 73
rect 99 72 100 73
rect 98 72 99 73
rect 97 72 98 73
rect 96 72 97 73
rect 95 72 96 73
rect 94 72 95 73
rect 93 72 94 73
rect 92 72 93 73
rect 91 72 92 73
rect 90 72 91 73
rect 89 72 90 73
rect 88 72 89 73
rect 87 72 88 73
rect 86 72 87 73
rect 85 72 86 73
rect 84 72 85 73
rect 83 72 84 73
rect 82 72 83 73
rect 81 72 82 73
rect 80 72 81 73
rect 79 72 80 73
rect 78 72 79 73
rect 77 72 78 73
rect 76 72 77 73
rect 75 72 76 73
rect 74 72 75 73
rect 73 72 74 73
rect 72 72 73 73
rect 71 72 72 73
rect 70 72 71 73
rect 439 73 440 74
rect 438 73 439 74
rect 437 73 438 74
rect 436 73 437 74
rect 435 73 436 74
rect 434 73 435 74
rect 433 73 434 74
rect 432 73 433 74
rect 431 73 432 74
rect 430 73 431 74
rect 429 73 430 74
rect 428 73 429 74
rect 427 73 428 74
rect 426 73 427 74
rect 425 73 426 74
rect 424 73 425 74
rect 423 73 424 74
rect 422 73 423 74
rect 421 73 422 74
rect 420 73 421 74
rect 419 73 420 74
rect 418 73 419 74
rect 417 73 418 74
rect 416 73 417 74
rect 415 73 416 74
rect 414 73 415 74
rect 413 73 414 74
rect 412 73 413 74
rect 411 73 412 74
rect 410 73 411 74
rect 144 73 145 74
rect 143 73 144 74
rect 142 73 143 74
rect 141 73 142 74
rect 140 73 141 74
rect 139 73 140 74
rect 138 73 139 74
rect 137 73 138 74
rect 136 73 137 74
rect 135 73 136 74
rect 134 73 135 74
rect 133 73 134 74
rect 132 73 133 74
rect 124 73 125 74
rect 123 73 124 74
rect 122 73 123 74
rect 121 73 122 74
rect 120 73 121 74
rect 119 73 120 74
rect 118 73 119 74
rect 117 73 118 74
rect 116 73 117 74
rect 115 73 116 74
rect 114 73 115 74
rect 113 73 114 74
rect 112 73 113 74
rect 111 73 112 74
rect 110 73 111 74
rect 109 73 110 74
rect 108 73 109 74
rect 107 73 108 74
rect 106 73 107 74
rect 105 73 106 74
rect 104 73 105 74
rect 103 73 104 74
rect 102 73 103 74
rect 101 73 102 74
rect 100 73 101 74
rect 99 73 100 74
rect 98 73 99 74
rect 97 73 98 74
rect 96 73 97 74
rect 95 73 96 74
rect 94 73 95 74
rect 93 73 94 74
rect 92 73 93 74
rect 91 73 92 74
rect 90 73 91 74
rect 89 73 90 74
rect 88 73 89 74
rect 87 73 88 74
rect 86 73 87 74
rect 85 73 86 74
rect 84 73 85 74
rect 83 73 84 74
rect 82 73 83 74
rect 81 73 82 74
rect 80 73 81 74
rect 79 73 80 74
rect 78 73 79 74
rect 77 73 78 74
rect 76 73 77 74
rect 75 73 76 74
rect 74 73 75 74
rect 73 73 74 74
rect 72 73 73 74
rect 71 73 72 74
rect 70 73 71 74
rect 69 73 70 74
rect 439 74 440 75
rect 438 74 439 75
rect 437 74 438 75
rect 436 74 437 75
rect 435 74 436 75
rect 434 74 435 75
rect 433 74 434 75
rect 432 74 433 75
rect 431 74 432 75
rect 430 74 431 75
rect 429 74 430 75
rect 428 74 429 75
rect 427 74 428 75
rect 426 74 427 75
rect 425 74 426 75
rect 424 74 425 75
rect 423 74 424 75
rect 422 74 423 75
rect 421 74 422 75
rect 420 74 421 75
rect 419 74 420 75
rect 418 74 419 75
rect 417 74 418 75
rect 416 74 417 75
rect 415 74 416 75
rect 414 74 415 75
rect 413 74 414 75
rect 412 74 413 75
rect 146 74 147 75
rect 145 74 146 75
rect 144 74 145 75
rect 143 74 144 75
rect 142 74 143 75
rect 141 74 142 75
rect 140 74 141 75
rect 139 74 140 75
rect 138 74 139 75
rect 137 74 138 75
rect 136 74 137 75
rect 135 74 136 75
rect 134 74 135 75
rect 133 74 134 75
rect 132 74 133 75
rect 131 74 132 75
rect 125 74 126 75
rect 124 74 125 75
rect 123 74 124 75
rect 122 74 123 75
rect 121 74 122 75
rect 120 74 121 75
rect 119 74 120 75
rect 118 74 119 75
rect 117 74 118 75
rect 116 74 117 75
rect 115 74 116 75
rect 114 74 115 75
rect 113 74 114 75
rect 112 74 113 75
rect 111 74 112 75
rect 110 74 111 75
rect 109 74 110 75
rect 108 74 109 75
rect 107 74 108 75
rect 106 74 107 75
rect 105 74 106 75
rect 104 74 105 75
rect 103 74 104 75
rect 102 74 103 75
rect 101 74 102 75
rect 100 74 101 75
rect 99 74 100 75
rect 98 74 99 75
rect 97 74 98 75
rect 96 74 97 75
rect 95 74 96 75
rect 94 74 95 75
rect 93 74 94 75
rect 92 74 93 75
rect 91 74 92 75
rect 90 74 91 75
rect 89 74 90 75
rect 88 74 89 75
rect 87 74 88 75
rect 86 74 87 75
rect 85 74 86 75
rect 84 74 85 75
rect 83 74 84 75
rect 82 74 83 75
rect 81 74 82 75
rect 80 74 81 75
rect 79 74 80 75
rect 78 74 79 75
rect 77 74 78 75
rect 76 74 77 75
rect 75 74 76 75
rect 74 74 75 75
rect 73 74 74 75
rect 72 74 73 75
rect 71 74 72 75
rect 70 74 71 75
rect 69 74 70 75
rect 439 75 440 76
rect 438 75 439 76
rect 437 75 438 76
rect 436 75 437 76
rect 435 75 436 76
rect 434 75 435 76
rect 433 75 434 76
rect 432 75 433 76
rect 431 75 432 76
rect 430 75 431 76
rect 429 75 430 76
rect 428 75 429 76
rect 427 75 428 76
rect 426 75 427 76
rect 425 75 426 76
rect 424 75 425 76
rect 423 75 424 76
rect 422 75 423 76
rect 421 75 422 76
rect 420 75 421 76
rect 419 75 420 76
rect 418 75 419 76
rect 417 75 418 76
rect 416 75 417 76
rect 415 75 416 76
rect 414 75 415 76
rect 147 75 148 76
rect 146 75 147 76
rect 145 75 146 76
rect 144 75 145 76
rect 143 75 144 76
rect 142 75 143 76
rect 141 75 142 76
rect 140 75 141 76
rect 139 75 140 76
rect 138 75 139 76
rect 137 75 138 76
rect 136 75 137 76
rect 135 75 136 76
rect 134 75 135 76
rect 133 75 134 76
rect 132 75 133 76
rect 131 75 132 76
rect 124 75 125 76
rect 123 75 124 76
rect 122 75 123 76
rect 121 75 122 76
rect 120 75 121 76
rect 119 75 120 76
rect 118 75 119 76
rect 117 75 118 76
rect 116 75 117 76
rect 115 75 116 76
rect 114 75 115 76
rect 113 75 114 76
rect 112 75 113 76
rect 111 75 112 76
rect 110 75 111 76
rect 109 75 110 76
rect 108 75 109 76
rect 107 75 108 76
rect 106 75 107 76
rect 105 75 106 76
rect 104 75 105 76
rect 103 75 104 76
rect 102 75 103 76
rect 101 75 102 76
rect 100 75 101 76
rect 99 75 100 76
rect 98 75 99 76
rect 97 75 98 76
rect 96 75 97 76
rect 95 75 96 76
rect 94 75 95 76
rect 93 75 94 76
rect 92 75 93 76
rect 91 75 92 76
rect 90 75 91 76
rect 89 75 90 76
rect 88 75 89 76
rect 87 75 88 76
rect 86 75 87 76
rect 85 75 86 76
rect 84 75 85 76
rect 83 75 84 76
rect 82 75 83 76
rect 81 75 82 76
rect 80 75 81 76
rect 79 75 80 76
rect 78 75 79 76
rect 77 75 78 76
rect 76 75 77 76
rect 75 75 76 76
rect 74 75 75 76
rect 73 75 74 76
rect 72 75 73 76
rect 71 75 72 76
rect 70 75 71 76
rect 69 75 70 76
rect 68 75 69 76
rect 439 76 440 77
rect 438 76 439 77
rect 437 76 438 77
rect 436 76 437 77
rect 435 76 436 77
rect 434 76 435 77
rect 433 76 434 77
rect 432 76 433 77
rect 431 76 432 77
rect 430 76 431 77
rect 429 76 430 77
rect 428 76 429 77
rect 427 76 428 77
rect 426 76 427 77
rect 425 76 426 77
rect 424 76 425 77
rect 423 76 424 77
rect 422 76 423 77
rect 421 76 422 77
rect 420 76 421 77
rect 419 76 420 77
rect 418 76 419 77
rect 417 76 418 77
rect 416 76 417 77
rect 149 76 150 77
rect 148 76 149 77
rect 147 76 148 77
rect 146 76 147 77
rect 145 76 146 77
rect 144 76 145 77
rect 143 76 144 77
rect 142 76 143 77
rect 141 76 142 77
rect 140 76 141 77
rect 139 76 140 77
rect 138 76 139 77
rect 137 76 138 77
rect 136 76 137 77
rect 135 76 136 77
rect 134 76 135 77
rect 133 76 134 77
rect 132 76 133 77
rect 131 76 132 77
rect 124 76 125 77
rect 123 76 124 77
rect 122 76 123 77
rect 121 76 122 77
rect 120 76 121 77
rect 119 76 120 77
rect 118 76 119 77
rect 117 76 118 77
rect 116 76 117 77
rect 115 76 116 77
rect 114 76 115 77
rect 113 76 114 77
rect 112 76 113 77
rect 111 76 112 77
rect 110 76 111 77
rect 109 76 110 77
rect 108 76 109 77
rect 107 76 108 77
rect 106 76 107 77
rect 105 76 106 77
rect 104 76 105 77
rect 103 76 104 77
rect 102 76 103 77
rect 101 76 102 77
rect 100 76 101 77
rect 99 76 100 77
rect 98 76 99 77
rect 97 76 98 77
rect 96 76 97 77
rect 95 76 96 77
rect 94 76 95 77
rect 93 76 94 77
rect 92 76 93 77
rect 91 76 92 77
rect 90 76 91 77
rect 89 76 90 77
rect 88 76 89 77
rect 87 76 88 77
rect 86 76 87 77
rect 85 76 86 77
rect 84 76 85 77
rect 83 76 84 77
rect 82 76 83 77
rect 81 76 82 77
rect 80 76 81 77
rect 79 76 80 77
rect 78 76 79 77
rect 77 76 78 77
rect 76 76 77 77
rect 75 76 76 77
rect 74 76 75 77
rect 73 76 74 77
rect 72 76 73 77
rect 71 76 72 77
rect 70 76 71 77
rect 69 76 70 77
rect 68 76 69 77
rect 439 77 440 78
rect 438 77 439 78
rect 437 77 438 78
rect 436 77 437 78
rect 435 77 436 78
rect 434 77 435 78
rect 433 77 434 78
rect 432 77 433 78
rect 431 77 432 78
rect 430 77 431 78
rect 429 77 430 78
rect 428 77 429 78
rect 427 77 428 78
rect 426 77 427 78
rect 425 77 426 78
rect 424 77 425 78
rect 423 77 424 78
rect 422 77 423 78
rect 421 77 422 78
rect 420 77 421 78
rect 419 77 420 78
rect 418 77 419 78
rect 417 77 418 78
rect 416 77 417 78
rect 415 77 416 78
rect 150 77 151 78
rect 149 77 150 78
rect 148 77 149 78
rect 147 77 148 78
rect 146 77 147 78
rect 145 77 146 78
rect 144 77 145 78
rect 143 77 144 78
rect 142 77 143 78
rect 141 77 142 78
rect 140 77 141 78
rect 139 77 140 78
rect 138 77 139 78
rect 137 77 138 78
rect 136 77 137 78
rect 135 77 136 78
rect 134 77 135 78
rect 133 77 134 78
rect 132 77 133 78
rect 131 77 132 78
rect 124 77 125 78
rect 123 77 124 78
rect 122 77 123 78
rect 121 77 122 78
rect 120 77 121 78
rect 119 77 120 78
rect 118 77 119 78
rect 117 77 118 78
rect 116 77 117 78
rect 115 77 116 78
rect 114 77 115 78
rect 113 77 114 78
rect 112 77 113 78
rect 111 77 112 78
rect 110 77 111 78
rect 109 77 110 78
rect 108 77 109 78
rect 107 77 108 78
rect 106 77 107 78
rect 105 77 106 78
rect 104 77 105 78
rect 103 77 104 78
rect 102 77 103 78
rect 101 77 102 78
rect 100 77 101 78
rect 99 77 100 78
rect 98 77 99 78
rect 97 77 98 78
rect 96 77 97 78
rect 95 77 96 78
rect 94 77 95 78
rect 93 77 94 78
rect 92 77 93 78
rect 91 77 92 78
rect 90 77 91 78
rect 89 77 90 78
rect 88 77 89 78
rect 87 77 88 78
rect 86 77 87 78
rect 85 77 86 78
rect 84 77 85 78
rect 83 77 84 78
rect 82 77 83 78
rect 81 77 82 78
rect 80 77 81 78
rect 79 77 80 78
rect 78 77 79 78
rect 77 77 78 78
rect 76 77 77 78
rect 75 77 76 78
rect 74 77 75 78
rect 73 77 74 78
rect 72 77 73 78
rect 71 77 72 78
rect 70 77 71 78
rect 69 77 70 78
rect 68 77 69 78
rect 67 77 68 78
rect 439 78 440 79
rect 438 78 439 79
rect 437 78 438 79
rect 436 78 437 79
rect 435 78 436 79
rect 434 78 435 79
rect 433 78 434 79
rect 432 78 433 79
rect 431 78 432 79
rect 430 78 431 79
rect 429 78 430 79
rect 428 78 429 79
rect 427 78 428 79
rect 426 78 427 79
rect 425 78 426 79
rect 424 78 425 79
rect 423 78 424 79
rect 422 78 423 79
rect 421 78 422 79
rect 420 78 421 79
rect 419 78 420 79
rect 418 78 419 79
rect 417 78 418 79
rect 416 78 417 79
rect 415 78 416 79
rect 414 78 415 79
rect 413 78 414 79
rect 152 78 153 79
rect 151 78 152 79
rect 150 78 151 79
rect 149 78 150 79
rect 148 78 149 79
rect 147 78 148 79
rect 146 78 147 79
rect 145 78 146 79
rect 144 78 145 79
rect 143 78 144 79
rect 142 78 143 79
rect 141 78 142 79
rect 140 78 141 79
rect 139 78 140 79
rect 138 78 139 79
rect 137 78 138 79
rect 136 78 137 79
rect 135 78 136 79
rect 134 78 135 79
rect 133 78 134 79
rect 132 78 133 79
rect 131 78 132 79
rect 124 78 125 79
rect 123 78 124 79
rect 122 78 123 79
rect 121 78 122 79
rect 120 78 121 79
rect 119 78 120 79
rect 118 78 119 79
rect 117 78 118 79
rect 116 78 117 79
rect 115 78 116 79
rect 114 78 115 79
rect 113 78 114 79
rect 112 78 113 79
rect 111 78 112 79
rect 110 78 111 79
rect 109 78 110 79
rect 108 78 109 79
rect 107 78 108 79
rect 106 78 107 79
rect 105 78 106 79
rect 104 78 105 79
rect 103 78 104 79
rect 102 78 103 79
rect 101 78 102 79
rect 100 78 101 79
rect 99 78 100 79
rect 98 78 99 79
rect 97 78 98 79
rect 96 78 97 79
rect 95 78 96 79
rect 94 78 95 79
rect 93 78 94 79
rect 92 78 93 79
rect 91 78 92 79
rect 90 78 91 79
rect 89 78 90 79
rect 88 78 89 79
rect 87 78 88 79
rect 86 78 87 79
rect 85 78 86 79
rect 84 78 85 79
rect 83 78 84 79
rect 82 78 83 79
rect 81 78 82 79
rect 80 78 81 79
rect 79 78 80 79
rect 78 78 79 79
rect 77 78 78 79
rect 76 78 77 79
rect 75 78 76 79
rect 74 78 75 79
rect 73 78 74 79
rect 72 78 73 79
rect 71 78 72 79
rect 70 78 71 79
rect 69 78 70 79
rect 68 78 69 79
rect 67 78 68 79
rect 439 79 440 80
rect 438 79 439 80
rect 437 79 438 80
rect 436 79 437 80
rect 417 79 418 80
rect 416 79 417 80
rect 415 79 416 80
rect 414 79 415 80
rect 413 79 414 80
rect 412 79 413 80
rect 411 79 412 80
rect 154 79 155 80
rect 153 79 154 80
rect 152 79 153 80
rect 151 79 152 80
rect 150 79 151 80
rect 149 79 150 80
rect 148 79 149 80
rect 147 79 148 80
rect 146 79 147 80
rect 145 79 146 80
rect 144 79 145 80
rect 143 79 144 80
rect 142 79 143 80
rect 141 79 142 80
rect 140 79 141 80
rect 139 79 140 80
rect 138 79 139 80
rect 137 79 138 80
rect 136 79 137 80
rect 135 79 136 80
rect 134 79 135 80
rect 133 79 134 80
rect 132 79 133 80
rect 131 79 132 80
rect 124 79 125 80
rect 123 79 124 80
rect 122 79 123 80
rect 121 79 122 80
rect 120 79 121 80
rect 119 79 120 80
rect 118 79 119 80
rect 117 79 118 80
rect 116 79 117 80
rect 115 79 116 80
rect 114 79 115 80
rect 113 79 114 80
rect 112 79 113 80
rect 111 79 112 80
rect 110 79 111 80
rect 109 79 110 80
rect 108 79 109 80
rect 107 79 108 80
rect 106 79 107 80
rect 105 79 106 80
rect 104 79 105 80
rect 103 79 104 80
rect 102 79 103 80
rect 101 79 102 80
rect 100 79 101 80
rect 99 79 100 80
rect 98 79 99 80
rect 97 79 98 80
rect 96 79 97 80
rect 95 79 96 80
rect 94 79 95 80
rect 93 79 94 80
rect 92 79 93 80
rect 91 79 92 80
rect 90 79 91 80
rect 89 79 90 80
rect 88 79 89 80
rect 87 79 88 80
rect 86 79 87 80
rect 85 79 86 80
rect 84 79 85 80
rect 83 79 84 80
rect 82 79 83 80
rect 81 79 82 80
rect 80 79 81 80
rect 79 79 80 80
rect 78 79 79 80
rect 77 79 78 80
rect 76 79 77 80
rect 75 79 76 80
rect 74 79 75 80
rect 73 79 74 80
rect 72 79 73 80
rect 71 79 72 80
rect 70 79 71 80
rect 69 79 70 80
rect 68 79 69 80
rect 67 79 68 80
rect 66 79 67 80
rect 439 80 440 81
rect 438 80 439 81
rect 437 80 438 81
rect 415 80 416 81
rect 414 80 415 81
rect 413 80 414 81
rect 412 80 413 81
rect 411 80 412 81
rect 410 80 411 81
rect 409 80 410 81
rect 397 80 398 81
rect 396 80 397 81
rect 395 80 396 81
rect 157 80 158 81
rect 156 80 157 81
rect 155 80 156 81
rect 154 80 155 81
rect 153 80 154 81
rect 152 80 153 81
rect 151 80 152 81
rect 150 80 151 81
rect 149 80 150 81
rect 148 80 149 81
rect 147 80 148 81
rect 146 80 147 81
rect 145 80 146 81
rect 144 80 145 81
rect 143 80 144 81
rect 142 80 143 81
rect 141 80 142 81
rect 140 80 141 81
rect 139 80 140 81
rect 138 80 139 81
rect 137 80 138 81
rect 136 80 137 81
rect 135 80 136 81
rect 134 80 135 81
rect 133 80 134 81
rect 132 80 133 81
rect 131 80 132 81
rect 124 80 125 81
rect 123 80 124 81
rect 122 80 123 81
rect 121 80 122 81
rect 120 80 121 81
rect 119 80 120 81
rect 118 80 119 81
rect 117 80 118 81
rect 116 80 117 81
rect 115 80 116 81
rect 114 80 115 81
rect 113 80 114 81
rect 112 80 113 81
rect 111 80 112 81
rect 110 80 111 81
rect 109 80 110 81
rect 108 80 109 81
rect 107 80 108 81
rect 106 80 107 81
rect 105 80 106 81
rect 104 80 105 81
rect 103 80 104 81
rect 102 80 103 81
rect 101 80 102 81
rect 100 80 101 81
rect 99 80 100 81
rect 98 80 99 81
rect 97 80 98 81
rect 96 80 97 81
rect 95 80 96 81
rect 94 80 95 81
rect 93 80 94 81
rect 92 80 93 81
rect 91 80 92 81
rect 90 80 91 81
rect 89 80 90 81
rect 88 80 89 81
rect 87 80 88 81
rect 86 80 87 81
rect 85 80 86 81
rect 84 80 85 81
rect 83 80 84 81
rect 82 80 83 81
rect 81 80 82 81
rect 80 80 81 81
rect 79 80 80 81
rect 78 80 79 81
rect 77 80 78 81
rect 76 80 77 81
rect 75 80 76 81
rect 74 80 75 81
rect 73 80 74 81
rect 72 80 73 81
rect 71 80 72 81
rect 70 80 71 81
rect 69 80 70 81
rect 68 80 69 81
rect 67 80 68 81
rect 66 80 67 81
rect 65 80 66 81
rect 460 81 461 82
rect 439 81 440 82
rect 438 81 439 82
rect 437 81 438 82
rect 413 81 414 82
rect 412 81 413 82
rect 411 81 412 82
rect 410 81 411 82
rect 409 81 410 82
rect 408 81 409 82
rect 407 81 408 82
rect 397 81 398 82
rect 396 81 397 82
rect 395 81 396 82
rect 159 81 160 82
rect 158 81 159 82
rect 157 81 158 82
rect 156 81 157 82
rect 155 81 156 82
rect 154 81 155 82
rect 153 81 154 82
rect 152 81 153 82
rect 151 81 152 82
rect 150 81 151 82
rect 149 81 150 82
rect 148 81 149 82
rect 147 81 148 82
rect 146 81 147 82
rect 145 81 146 82
rect 144 81 145 82
rect 143 81 144 82
rect 142 81 143 82
rect 141 81 142 82
rect 140 81 141 82
rect 139 81 140 82
rect 138 81 139 82
rect 137 81 138 82
rect 136 81 137 82
rect 135 81 136 82
rect 134 81 135 82
rect 133 81 134 82
rect 132 81 133 82
rect 131 81 132 82
rect 124 81 125 82
rect 123 81 124 82
rect 122 81 123 82
rect 121 81 122 82
rect 120 81 121 82
rect 119 81 120 82
rect 118 81 119 82
rect 117 81 118 82
rect 116 81 117 82
rect 115 81 116 82
rect 114 81 115 82
rect 113 81 114 82
rect 112 81 113 82
rect 111 81 112 82
rect 110 81 111 82
rect 109 81 110 82
rect 108 81 109 82
rect 107 81 108 82
rect 106 81 107 82
rect 105 81 106 82
rect 104 81 105 82
rect 103 81 104 82
rect 102 81 103 82
rect 101 81 102 82
rect 100 81 101 82
rect 99 81 100 82
rect 98 81 99 82
rect 97 81 98 82
rect 96 81 97 82
rect 95 81 96 82
rect 94 81 95 82
rect 93 81 94 82
rect 92 81 93 82
rect 91 81 92 82
rect 90 81 91 82
rect 89 81 90 82
rect 88 81 89 82
rect 87 81 88 82
rect 86 81 87 82
rect 85 81 86 82
rect 84 81 85 82
rect 83 81 84 82
rect 82 81 83 82
rect 81 81 82 82
rect 80 81 81 82
rect 79 81 80 82
rect 78 81 79 82
rect 77 81 78 82
rect 76 81 77 82
rect 75 81 76 82
rect 74 81 75 82
rect 73 81 74 82
rect 72 81 73 82
rect 71 81 72 82
rect 70 81 71 82
rect 69 81 70 82
rect 68 81 69 82
rect 67 81 68 82
rect 66 81 67 82
rect 65 81 66 82
rect 460 82 461 83
rect 439 82 440 83
rect 438 82 439 83
rect 437 82 438 83
rect 411 82 412 83
rect 410 82 411 83
rect 409 82 410 83
rect 408 82 409 83
rect 407 82 408 83
rect 406 82 407 83
rect 405 82 406 83
rect 397 82 398 83
rect 396 82 397 83
rect 395 82 396 83
rect 161 82 162 83
rect 160 82 161 83
rect 159 82 160 83
rect 158 82 159 83
rect 157 82 158 83
rect 156 82 157 83
rect 155 82 156 83
rect 154 82 155 83
rect 153 82 154 83
rect 152 82 153 83
rect 151 82 152 83
rect 150 82 151 83
rect 149 82 150 83
rect 148 82 149 83
rect 147 82 148 83
rect 146 82 147 83
rect 145 82 146 83
rect 144 82 145 83
rect 143 82 144 83
rect 142 82 143 83
rect 141 82 142 83
rect 140 82 141 83
rect 139 82 140 83
rect 138 82 139 83
rect 137 82 138 83
rect 136 82 137 83
rect 135 82 136 83
rect 134 82 135 83
rect 133 82 134 83
rect 132 82 133 83
rect 131 82 132 83
rect 124 82 125 83
rect 123 82 124 83
rect 122 82 123 83
rect 121 82 122 83
rect 120 82 121 83
rect 119 82 120 83
rect 118 82 119 83
rect 117 82 118 83
rect 116 82 117 83
rect 115 82 116 83
rect 114 82 115 83
rect 113 82 114 83
rect 112 82 113 83
rect 111 82 112 83
rect 110 82 111 83
rect 109 82 110 83
rect 108 82 109 83
rect 107 82 108 83
rect 106 82 107 83
rect 105 82 106 83
rect 104 82 105 83
rect 103 82 104 83
rect 102 82 103 83
rect 101 82 102 83
rect 100 82 101 83
rect 99 82 100 83
rect 98 82 99 83
rect 97 82 98 83
rect 96 82 97 83
rect 95 82 96 83
rect 94 82 95 83
rect 93 82 94 83
rect 92 82 93 83
rect 91 82 92 83
rect 90 82 91 83
rect 89 82 90 83
rect 88 82 89 83
rect 87 82 88 83
rect 86 82 87 83
rect 85 82 86 83
rect 84 82 85 83
rect 83 82 84 83
rect 82 82 83 83
rect 81 82 82 83
rect 80 82 81 83
rect 79 82 80 83
rect 78 82 79 83
rect 77 82 78 83
rect 76 82 77 83
rect 75 82 76 83
rect 74 82 75 83
rect 73 82 74 83
rect 72 82 73 83
rect 71 82 72 83
rect 70 82 71 83
rect 69 82 70 83
rect 68 82 69 83
rect 67 82 68 83
rect 66 82 67 83
rect 65 82 66 83
rect 64 82 65 83
rect 461 83 462 84
rect 460 83 461 84
rect 439 83 440 84
rect 438 83 439 84
rect 437 83 438 84
rect 410 83 411 84
rect 409 83 410 84
rect 408 83 409 84
rect 407 83 408 84
rect 406 83 407 84
rect 405 83 406 84
rect 404 83 405 84
rect 403 83 404 84
rect 397 83 398 84
rect 396 83 397 84
rect 395 83 396 84
rect 225 83 226 84
rect 224 83 225 84
rect 223 83 224 84
rect 222 83 223 84
rect 221 83 222 84
rect 220 83 221 84
rect 219 83 220 84
rect 218 83 219 84
rect 217 83 218 84
rect 216 83 217 84
rect 215 83 216 84
rect 214 83 215 84
rect 213 83 214 84
rect 212 83 213 84
rect 211 83 212 84
rect 210 83 211 84
rect 209 83 210 84
rect 162 83 163 84
rect 161 83 162 84
rect 160 83 161 84
rect 159 83 160 84
rect 158 83 159 84
rect 157 83 158 84
rect 156 83 157 84
rect 155 83 156 84
rect 154 83 155 84
rect 153 83 154 84
rect 152 83 153 84
rect 151 83 152 84
rect 150 83 151 84
rect 149 83 150 84
rect 148 83 149 84
rect 147 83 148 84
rect 146 83 147 84
rect 145 83 146 84
rect 144 83 145 84
rect 143 83 144 84
rect 142 83 143 84
rect 141 83 142 84
rect 140 83 141 84
rect 139 83 140 84
rect 138 83 139 84
rect 137 83 138 84
rect 136 83 137 84
rect 135 83 136 84
rect 134 83 135 84
rect 133 83 134 84
rect 132 83 133 84
rect 131 83 132 84
rect 124 83 125 84
rect 123 83 124 84
rect 122 83 123 84
rect 121 83 122 84
rect 120 83 121 84
rect 119 83 120 84
rect 118 83 119 84
rect 117 83 118 84
rect 116 83 117 84
rect 115 83 116 84
rect 114 83 115 84
rect 113 83 114 84
rect 112 83 113 84
rect 111 83 112 84
rect 110 83 111 84
rect 109 83 110 84
rect 108 83 109 84
rect 107 83 108 84
rect 106 83 107 84
rect 105 83 106 84
rect 104 83 105 84
rect 103 83 104 84
rect 102 83 103 84
rect 101 83 102 84
rect 100 83 101 84
rect 99 83 100 84
rect 98 83 99 84
rect 97 83 98 84
rect 96 83 97 84
rect 95 83 96 84
rect 94 83 95 84
rect 93 83 94 84
rect 92 83 93 84
rect 91 83 92 84
rect 90 83 91 84
rect 89 83 90 84
rect 88 83 89 84
rect 87 83 88 84
rect 86 83 87 84
rect 85 83 86 84
rect 84 83 85 84
rect 83 83 84 84
rect 82 83 83 84
rect 81 83 82 84
rect 80 83 81 84
rect 79 83 80 84
rect 78 83 79 84
rect 77 83 78 84
rect 76 83 77 84
rect 75 83 76 84
rect 74 83 75 84
rect 73 83 74 84
rect 72 83 73 84
rect 71 83 72 84
rect 70 83 71 84
rect 69 83 70 84
rect 68 83 69 84
rect 67 83 68 84
rect 66 83 67 84
rect 65 83 66 84
rect 64 83 65 84
rect 476 84 477 85
rect 475 84 476 85
rect 474 84 475 85
rect 473 84 474 85
rect 472 84 473 85
rect 471 84 472 85
rect 470 84 471 85
rect 469 84 470 85
rect 468 84 469 85
rect 467 84 468 85
rect 466 84 467 85
rect 465 84 466 85
rect 464 84 465 85
rect 463 84 464 85
rect 462 84 463 85
rect 461 84 462 85
rect 460 84 461 85
rect 439 84 440 85
rect 438 84 439 85
rect 408 84 409 85
rect 407 84 408 85
rect 406 84 407 85
rect 405 84 406 85
rect 404 84 405 85
rect 403 84 404 85
rect 402 84 403 85
rect 401 84 402 85
rect 400 84 401 85
rect 399 84 400 85
rect 398 84 399 85
rect 397 84 398 85
rect 396 84 397 85
rect 395 84 396 85
rect 231 84 232 85
rect 230 84 231 85
rect 229 84 230 85
rect 228 84 229 85
rect 227 84 228 85
rect 226 84 227 85
rect 225 84 226 85
rect 224 84 225 85
rect 223 84 224 85
rect 222 84 223 85
rect 221 84 222 85
rect 220 84 221 85
rect 219 84 220 85
rect 218 84 219 85
rect 217 84 218 85
rect 216 84 217 85
rect 215 84 216 85
rect 214 84 215 85
rect 213 84 214 85
rect 212 84 213 85
rect 211 84 212 85
rect 210 84 211 85
rect 209 84 210 85
rect 208 84 209 85
rect 207 84 208 85
rect 206 84 207 85
rect 205 84 206 85
rect 204 84 205 85
rect 162 84 163 85
rect 161 84 162 85
rect 160 84 161 85
rect 159 84 160 85
rect 158 84 159 85
rect 157 84 158 85
rect 156 84 157 85
rect 155 84 156 85
rect 154 84 155 85
rect 153 84 154 85
rect 152 84 153 85
rect 151 84 152 85
rect 150 84 151 85
rect 149 84 150 85
rect 148 84 149 85
rect 147 84 148 85
rect 146 84 147 85
rect 145 84 146 85
rect 144 84 145 85
rect 143 84 144 85
rect 142 84 143 85
rect 141 84 142 85
rect 140 84 141 85
rect 139 84 140 85
rect 138 84 139 85
rect 137 84 138 85
rect 136 84 137 85
rect 135 84 136 85
rect 134 84 135 85
rect 133 84 134 85
rect 132 84 133 85
rect 131 84 132 85
rect 130 84 131 85
rect 123 84 124 85
rect 122 84 123 85
rect 121 84 122 85
rect 120 84 121 85
rect 119 84 120 85
rect 118 84 119 85
rect 117 84 118 85
rect 116 84 117 85
rect 115 84 116 85
rect 114 84 115 85
rect 113 84 114 85
rect 112 84 113 85
rect 111 84 112 85
rect 110 84 111 85
rect 109 84 110 85
rect 108 84 109 85
rect 107 84 108 85
rect 106 84 107 85
rect 105 84 106 85
rect 104 84 105 85
rect 103 84 104 85
rect 102 84 103 85
rect 101 84 102 85
rect 100 84 101 85
rect 99 84 100 85
rect 98 84 99 85
rect 97 84 98 85
rect 96 84 97 85
rect 95 84 96 85
rect 94 84 95 85
rect 93 84 94 85
rect 92 84 93 85
rect 91 84 92 85
rect 90 84 91 85
rect 89 84 90 85
rect 88 84 89 85
rect 87 84 88 85
rect 86 84 87 85
rect 85 84 86 85
rect 84 84 85 85
rect 83 84 84 85
rect 82 84 83 85
rect 81 84 82 85
rect 80 84 81 85
rect 79 84 80 85
rect 78 84 79 85
rect 77 84 78 85
rect 76 84 77 85
rect 75 84 76 85
rect 74 84 75 85
rect 73 84 74 85
rect 72 84 73 85
rect 71 84 72 85
rect 70 84 71 85
rect 69 84 70 85
rect 68 84 69 85
rect 67 84 68 85
rect 66 84 67 85
rect 65 84 66 85
rect 64 84 65 85
rect 63 84 64 85
rect 478 85 479 86
rect 477 85 478 86
rect 476 85 477 86
rect 475 85 476 86
rect 474 85 475 86
rect 473 85 474 86
rect 472 85 473 86
rect 471 85 472 86
rect 470 85 471 86
rect 469 85 470 86
rect 468 85 469 86
rect 467 85 468 86
rect 466 85 467 86
rect 465 85 466 86
rect 464 85 465 86
rect 463 85 464 86
rect 462 85 463 86
rect 461 85 462 86
rect 460 85 461 86
rect 439 85 440 86
rect 438 85 439 86
rect 406 85 407 86
rect 405 85 406 86
rect 404 85 405 86
rect 403 85 404 86
rect 402 85 403 86
rect 401 85 402 86
rect 400 85 401 86
rect 399 85 400 86
rect 398 85 399 86
rect 397 85 398 86
rect 396 85 397 86
rect 395 85 396 86
rect 235 85 236 86
rect 234 85 235 86
rect 233 85 234 86
rect 232 85 233 86
rect 231 85 232 86
rect 230 85 231 86
rect 229 85 230 86
rect 228 85 229 86
rect 227 85 228 86
rect 226 85 227 86
rect 225 85 226 86
rect 224 85 225 86
rect 223 85 224 86
rect 222 85 223 86
rect 221 85 222 86
rect 220 85 221 86
rect 219 85 220 86
rect 218 85 219 86
rect 217 85 218 86
rect 216 85 217 86
rect 215 85 216 86
rect 214 85 215 86
rect 213 85 214 86
rect 212 85 213 86
rect 211 85 212 86
rect 210 85 211 86
rect 209 85 210 86
rect 208 85 209 86
rect 207 85 208 86
rect 206 85 207 86
rect 205 85 206 86
rect 204 85 205 86
rect 203 85 204 86
rect 202 85 203 86
rect 201 85 202 86
rect 200 85 201 86
rect 162 85 163 86
rect 161 85 162 86
rect 160 85 161 86
rect 159 85 160 86
rect 158 85 159 86
rect 157 85 158 86
rect 156 85 157 86
rect 155 85 156 86
rect 154 85 155 86
rect 153 85 154 86
rect 152 85 153 86
rect 151 85 152 86
rect 150 85 151 86
rect 149 85 150 86
rect 148 85 149 86
rect 147 85 148 86
rect 146 85 147 86
rect 145 85 146 86
rect 144 85 145 86
rect 143 85 144 86
rect 142 85 143 86
rect 141 85 142 86
rect 140 85 141 86
rect 139 85 140 86
rect 138 85 139 86
rect 137 85 138 86
rect 136 85 137 86
rect 135 85 136 86
rect 134 85 135 86
rect 133 85 134 86
rect 132 85 133 86
rect 131 85 132 86
rect 130 85 131 86
rect 123 85 124 86
rect 122 85 123 86
rect 121 85 122 86
rect 120 85 121 86
rect 119 85 120 86
rect 118 85 119 86
rect 117 85 118 86
rect 116 85 117 86
rect 115 85 116 86
rect 114 85 115 86
rect 113 85 114 86
rect 112 85 113 86
rect 111 85 112 86
rect 110 85 111 86
rect 109 85 110 86
rect 108 85 109 86
rect 107 85 108 86
rect 106 85 107 86
rect 105 85 106 86
rect 104 85 105 86
rect 103 85 104 86
rect 102 85 103 86
rect 101 85 102 86
rect 100 85 101 86
rect 99 85 100 86
rect 98 85 99 86
rect 97 85 98 86
rect 96 85 97 86
rect 95 85 96 86
rect 94 85 95 86
rect 93 85 94 86
rect 92 85 93 86
rect 91 85 92 86
rect 90 85 91 86
rect 89 85 90 86
rect 88 85 89 86
rect 87 85 88 86
rect 86 85 87 86
rect 85 85 86 86
rect 84 85 85 86
rect 83 85 84 86
rect 82 85 83 86
rect 81 85 82 86
rect 80 85 81 86
rect 79 85 80 86
rect 78 85 79 86
rect 77 85 78 86
rect 76 85 77 86
rect 75 85 76 86
rect 74 85 75 86
rect 73 85 74 86
rect 72 85 73 86
rect 71 85 72 86
rect 70 85 71 86
rect 69 85 70 86
rect 68 85 69 86
rect 67 85 68 86
rect 66 85 67 86
rect 65 85 66 86
rect 64 85 65 86
rect 63 85 64 86
rect 62 85 63 86
rect 479 86 480 87
rect 478 86 479 87
rect 477 86 478 87
rect 476 86 477 87
rect 475 86 476 87
rect 474 86 475 87
rect 473 86 474 87
rect 472 86 473 87
rect 471 86 472 87
rect 470 86 471 87
rect 469 86 470 87
rect 468 86 469 87
rect 467 86 468 87
rect 466 86 467 87
rect 465 86 466 87
rect 464 86 465 87
rect 463 86 464 87
rect 462 86 463 87
rect 461 86 462 87
rect 460 86 461 87
rect 405 86 406 87
rect 404 86 405 87
rect 403 86 404 87
rect 402 86 403 87
rect 401 86 402 87
rect 400 86 401 87
rect 399 86 400 87
rect 398 86 399 87
rect 397 86 398 87
rect 396 86 397 87
rect 395 86 396 87
rect 238 86 239 87
rect 237 86 238 87
rect 236 86 237 87
rect 235 86 236 87
rect 234 86 235 87
rect 233 86 234 87
rect 232 86 233 87
rect 231 86 232 87
rect 230 86 231 87
rect 229 86 230 87
rect 228 86 229 87
rect 227 86 228 87
rect 226 86 227 87
rect 225 86 226 87
rect 224 86 225 87
rect 223 86 224 87
rect 222 86 223 87
rect 221 86 222 87
rect 220 86 221 87
rect 219 86 220 87
rect 218 86 219 87
rect 217 86 218 87
rect 216 86 217 87
rect 215 86 216 87
rect 214 86 215 87
rect 213 86 214 87
rect 212 86 213 87
rect 211 86 212 87
rect 210 86 211 87
rect 209 86 210 87
rect 208 86 209 87
rect 207 86 208 87
rect 206 86 207 87
rect 205 86 206 87
rect 204 86 205 87
rect 203 86 204 87
rect 202 86 203 87
rect 201 86 202 87
rect 200 86 201 87
rect 199 86 200 87
rect 198 86 199 87
rect 162 86 163 87
rect 161 86 162 87
rect 160 86 161 87
rect 159 86 160 87
rect 158 86 159 87
rect 157 86 158 87
rect 156 86 157 87
rect 155 86 156 87
rect 154 86 155 87
rect 153 86 154 87
rect 152 86 153 87
rect 151 86 152 87
rect 150 86 151 87
rect 149 86 150 87
rect 148 86 149 87
rect 147 86 148 87
rect 146 86 147 87
rect 145 86 146 87
rect 144 86 145 87
rect 143 86 144 87
rect 142 86 143 87
rect 141 86 142 87
rect 140 86 141 87
rect 139 86 140 87
rect 138 86 139 87
rect 137 86 138 87
rect 136 86 137 87
rect 135 86 136 87
rect 134 86 135 87
rect 133 86 134 87
rect 132 86 133 87
rect 131 86 132 87
rect 130 86 131 87
rect 123 86 124 87
rect 122 86 123 87
rect 121 86 122 87
rect 120 86 121 87
rect 119 86 120 87
rect 118 86 119 87
rect 117 86 118 87
rect 116 86 117 87
rect 115 86 116 87
rect 114 86 115 87
rect 113 86 114 87
rect 112 86 113 87
rect 111 86 112 87
rect 110 86 111 87
rect 109 86 110 87
rect 108 86 109 87
rect 107 86 108 87
rect 106 86 107 87
rect 105 86 106 87
rect 104 86 105 87
rect 103 86 104 87
rect 102 86 103 87
rect 101 86 102 87
rect 100 86 101 87
rect 99 86 100 87
rect 98 86 99 87
rect 97 86 98 87
rect 96 86 97 87
rect 95 86 96 87
rect 94 86 95 87
rect 93 86 94 87
rect 92 86 93 87
rect 91 86 92 87
rect 90 86 91 87
rect 89 86 90 87
rect 88 86 89 87
rect 87 86 88 87
rect 86 86 87 87
rect 85 86 86 87
rect 84 86 85 87
rect 83 86 84 87
rect 82 86 83 87
rect 81 86 82 87
rect 80 86 81 87
rect 79 86 80 87
rect 78 86 79 87
rect 77 86 78 87
rect 76 86 77 87
rect 75 86 76 87
rect 74 86 75 87
rect 73 86 74 87
rect 72 86 73 87
rect 71 86 72 87
rect 70 86 71 87
rect 69 86 70 87
rect 68 86 69 87
rect 67 86 68 87
rect 66 86 67 87
rect 65 86 66 87
rect 64 86 65 87
rect 63 86 64 87
rect 62 86 63 87
rect 480 87 481 88
rect 479 87 480 88
rect 478 87 479 88
rect 477 87 478 88
rect 476 87 477 88
rect 475 87 476 88
rect 474 87 475 88
rect 473 87 474 88
rect 472 87 473 88
rect 471 87 472 88
rect 470 87 471 88
rect 469 87 470 88
rect 468 87 469 88
rect 467 87 468 88
rect 466 87 467 88
rect 465 87 466 88
rect 464 87 465 88
rect 463 87 464 88
rect 462 87 463 88
rect 461 87 462 88
rect 460 87 461 88
rect 403 87 404 88
rect 402 87 403 88
rect 401 87 402 88
rect 400 87 401 88
rect 399 87 400 88
rect 398 87 399 88
rect 397 87 398 88
rect 396 87 397 88
rect 395 87 396 88
rect 241 87 242 88
rect 240 87 241 88
rect 239 87 240 88
rect 238 87 239 88
rect 237 87 238 88
rect 236 87 237 88
rect 235 87 236 88
rect 234 87 235 88
rect 233 87 234 88
rect 232 87 233 88
rect 231 87 232 88
rect 230 87 231 88
rect 229 87 230 88
rect 228 87 229 88
rect 227 87 228 88
rect 226 87 227 88
rect 225 87 226 88
rect 224 87 225 88
rect 223 87 224 88
rect 222 87 223 88
rect 221 87 222 88
rect 220 87 221 88
rect 219 87 220 88
rect 218 87 219 88
rect 217 87 218 88
rect 216 87 217 88
rect 215 87 216 88
rect 214 87 215 88
rect 213 87 214 88
rect 212 87 213 88
rect 211 87 212 88
rect 210 87 211 88
rect 209 87 210 88
rect 208 87 209 88
rect 207 87 208 88
rect 206 87 207 88
rect 205 87 206 88
rect 204 87 205 88
rect 203 87 204 88
rect 202 87 203 88
rect 201 87 202 88
rect 200 87 201 88
rect 199 87 200 88
rect 198 87 199 88
rect 197 87 198 88
rect 196 87 197 88
rect 162 87 163 88
rect 161 87 162 88
rect 160 87 161 88
rect 159 87 160 88
rect 158 87 159 88
rect 157 87 158 88
rect 156 87 157 88
rect 155 87 156 88
rect 154 87 155 88
rect 153 87 154 88
rect 152 87 153 88
rect 151 87 152 88
rect 150 87 151 88
rect 149 87 150 88
rect 148 87 149 88
rect 147 87 148 88
rect 146 87 147 88
rect 145 87 146 88
rect 144 87 145 88
rect 143 87 144 88
rect 142 87 143 88
rect 141 87 142 88
rect 140 87 141 88
rect 139 87 140 88
rect 138 87 139 88
rect 137 87 138 88
rect 136 87 137 88
rect 135 87 136 88
rect 134 87 135 88
rect 133 87 134 88
rect 132 87 133 88
rect 131 87 132 88
rect 130 87 131 88
rect 123 87 124 88
rect 122 87 123 88
rect 121 87 122 88
rect 120 87 121 88
rect 119 87 120 88
rect 118 87 119 88
rect 117 87 118 88
rect 116 87 117 88
rect 115 87 116 88
rect 114 87 115 88
rect 113 87 114 88
rect 112 87 113 88
rect 111 87 112 88
rect 110 87 111 88
rect 109 87 110 88
rect 108 87 109 88
rect 107 87 108 88
rect 106 87 107 88
rect 105 87 106 88
rect 104 87 105 88
rect 103 87 104 88
rect 102 87 103 88
rect 101 87 102 88
rect 100 87 101 88
rect 99 87 100 88
rect 98 87 99 88
rect 97 87 98 88
rect 96 87 97 88
rect 95 87 96 88
rect 94 87 95 88
rect 93 87 94 88
rect 92 87 93 88
rect 91 87 92 88
rect 90 87 91 88
rect 89 87 90 88
rect 88 87 89 88
rect 87 87 88 88
rect 86 87 87 88
rect 85 87 86 88
rect 84 87 85 88
rect 83 87 84 88
rect 82 87 83 88
rect 81 87 82 88
rect 80 87 81 88
rect 79 87 80 88
rect 78 87 79 88
rect 77 87 78 88
rect 76 87 77 88
rect 75 87 76 88
rect 74 87 75 88
rect 73 87 74 88
rect 72 87 73 88
rect 71 87 72 88
rect 70 87 71 88
rect 69 87 70 88
rect 68 87 69 88
rect 67 87 68 88
rect 66 87 67 88
rect 65 87 66 88
rect 64 87 65 88
rect 63 87 64 88
rect 62 87 63 88
rect 61 87 62 88
rect 481 88 482 89
rect 480 88 481 89
rect 479 88 480 89
rect 478 88 479 89
rect 477 88 478 89
rect 476 88 477 89
rect 475 88 476 89
rect 474 88 475 89
rect 473 88 474 89
rect 462 88 463 89
rect 461 88 462 89
rect 460 88 461 89
rect 401 88 402 89
rect 400 88 401 89
rect 399 88 400 89
rect 398 88 399 89
rect 397 88 398 89
rect 396 88 397 89
rect 395 88 396 89
rect 243 88 244 89
rect 242 88 243 89
rect 241 88 242 89
rect 240 88 241 89
rect 239 88 240 89
rect 238 88 239 89
rect 237 88 238 89
rect 236 88 237 89
rect 235 88 236 89
rect 234 88 235 89
rect 233 88 234 89
rect 232 88 233 89
rect 231 88 232 89
rect 230 88 231 89
rect 229 88 230 89
rect 228 88 229 89
rect 227 88 228 89
rect 226 88 227 89
rect 225 88 226 89
rect 224 88 225 89
rect 223 88 224 89
rect 222 88 223 89
rect 221 88 222 89
rect 220 88 221 89
rect 219 88 220 89
rect 218 88 219 89
rect 217 88 218 89
rect 216 88 217 89
rect 215 88 216 89
rect 214 88 215 89
rect 213 88 214 89
rect 212 88 213 89
rect 211 88 212 89
rect 210 88 211 89
rect 209 88 210 89
rect 208 88 209 89
rect 207 88 208 89
rect 206 88 207 89
rect 205 88 206 89
rect 204 88 205 89
rect 203 88 204 89
rect 202 88 203 89
rect 201 88 202 89
rect 200 88 201 89
rect 199 88 200 89
rect 198 88 199 89
rect 197 88 198 89
rect 196 88 197 89
rect 195 88 196 89
rect 194 88 195 89
rect 162 88 163 89
rect 161 88 162 89
rect 160 88 161 89
rect 159 88 160 89
rect 158 88 159 89
rect 157 88 158 89
rect 156 88 157 89
rect 155 88 156 89
rect 154 88 155 89
rect 153 88 154 89
rect 152 88 153 89
rect 151 88 152 89
rect 150 88 151 89
rect 149 88 150 89
rect 148 88 149 89
rect 147 88 148 89
rect 146 88 147 89
rect 145 88 146 89
rect 144 88 145 89
rect 143 88 144 89
rect 142 88 143 89
rect 141 88 142 89
rect 140 88 141 89
rect 139 88 140 89
rect 138 88 139 89
rect 137 88 138 89
rect 136 88 137 89
rect 135 88 136 89
rect 134 88 135 89
rect 133 88 134 89
rect 132 88 133 89
rect 131 88 132 89
rect 130 88 131 89
rect 123 88 124 89
rect 122 88 123 89
rect 121 88 122 89
rect 120 88 121 89
rect 119 88 120 89
rect 118 88 119 89
rect 117 88 118 89
rect 116 88 117 89
rect 115 88 116 89
rect 114 88 115 89
rect 113 88 114 89
rect 112 88 113 89
rect 111 88 112 89
rect 110 88 111 89
rect 109 88 110 89
rect 108 88 109 89
rect 107 88 108 89
rect 106 88 107 89
rect 105 88 106 89
rect 104 88 105 89
rect 103 88 104 89
rect 102 88 103 89
rect 101 88 102 89
rect 100 88 101 89
rect 99 88 100 89
rect 98 88 99 89
rect 97 88 98 89
rect 96 88 97 89
rect 95 88 96 89
rect 94 88 95 89
rect 93 88 94 89
rect 92 88 93 89
rect 91 88 92 89
rect 90 88 91 89
rect 89 88 90 89
rect 88 88 89 89
rect 87 88 88 89
rect 86 88 87 89
rect 85 88 86 89
rect 84 88 85 89
rect 83 88 84 89
rect 82 88 83 89
rect 81 88 82 89
rect 80 88 81 89
rect 79 88 80 89
rect 78 88 79 89
rect 77 88 78 89
rect 76 88 77 89
rect 75 88 76 89
rect 74 88 75 89
rect 73 88 74 89
rect 72 88 73 89
rect 71 88 72 89
rect 70 88 71 89
rect 69 88 70 89
rect 68 88 69 89
rect 67 88 68 89
rect 66 88 67 89
rect 65 88 66 89
rect 64 88 65 89
rect 63 88 64 89
rect 62 88 63 89
rect 61 88 62 89
rect 60 88 61 89
rect 481 89 482 90
rect 480 89 481 90
rect 479 89 480 90
rect 478 89 479 90
rect 477 89 478 90
rect 460 89 461 90
rect 400 89 401 90
rect 399 89 400 90
rect 398 89 399 90
rect 397 89 398 90
rect 396 89 397 90
rect 395 89 396 90
rect 246 89 247 90
rect 245 89 246 90
rect 244 89 245 90
rect 243 89 244 90
rect 242 89 243 90
rect 241 89 242 90
rect 240 89 241 90
rect 239 89 240 90
rect 238 89 239 90
rect 237 89 238 90
rect 236 89 237 90
rect 235 89 236 90
rect 234 89 235 90
rect 233 89 234 90
rect 232 89 233 90
rect 231 89 232 90
rect 230 89 231 90
rect 229 89 230 90
rect 228 89 229 90
rect 227 89 228 90
rect 226 89 227 90
rect 225 89 226 90
rect 224 89 225 90
rect 223 89 224 90
rect 222 89 223 90
rect 221 89 222 90
rect 220 89 221 90
rect 219 89 220 90
rect 218 89 219 90
rect 217 89 218 90
rect 216 89 217 90
rect 215 89 216 90
rect 214 89 215 90
rect 213 89 214 90
rect 212 89 213 90
rect 211 89 212 90
rect 210 89 211 90
rect 209 89 210 90
rect 208 89 209 90
rect 207 89 208 90
rect 206 89 207 90
rect 205 89 206 90
rect 204 89 205 90
rect 203 89 204 90
rect 202 89 203 90
rect 201 89 202 90
rect 200 89 201 90
rect 199 89 200 90
rect 198 89 199 90
rect 197 89 198 90
rect 196 89 197 90
rect 195 89 196 90
rect 194 89 195 90
rect 193 89 194 90
rect 192 89 193 90
rect 162 89 163 90
rect 161 89 162 90
rect 160 89 161 90
rect 159 89 160 90
rect 158 89 159 90
rect 157 89 158 90
rect 156 89 157 90
rect 155 89 156 90
rect 154 89 155 90
rect 153 89 154 90
rect 152 89 153 90
rect 151 89 152 90
rect 150 89 151 90
rect 149 89 150 90
rect 148 89 149 90
rect 147 89 148 90
rect 146 89 147 90
rect 145 89 146 90
rect 144 89 145 90
rect 143 89 144 90
rect 142 89 143 90
rect 141 89 142 90
rect 140 89 141 90
rect 139 89 140 90
rect 138 89 139 90
rect 137 89 138 90
rect 136 89 137 90
rect 135 89 136 90
rect 134 89 135 90
rect 133 89 134 90
rect 132 89 133 90
rect 131 89 132 90
rect 130 89 131 90
rect 123 89 124 90
rect 122 89 123 90
rect 121 89 122 90
rect 120 89 121 90
rect 119 89 120 90
rect 118 89 119 90
rect 117 89 118 90
rect 116 89 117 90
rect 115 89 116 90
rect 114 89 115 90
rect 113 89 114 90
rect 112 89 113 90
rect 111 89 112 90
rect 110 89 111 90
rect 109 89 110 90
rect 108 89 109 90
rect 107 89 108 90
rect 106 89 107 90
rect 105 89 106 90
rect 104 89 105 90
rect 103 89 104 90
rect 102 89 103 90
rect 101 89 102 90
rect 100 89 101 90
rect 99 89 100 90
rect 98 89 99 90
rect 97 89 98 90
rect 96 89 97 90
rect 95 89 96 90
rect 94 89 95 90
rect 93 89 94 90
rect 92 89 93 90
rect 91 89 92 90
rect 90 89 91 90
rect 89 89 90 90
rect 88 89 89 90
rect 87 89 88 90
rect 86 89 87 90
rect 85 89 86 90
rect 84 89 85 90
rect 83 89 84 90
rect 82 89 83 90
rect 81 89 82 90
rect 80 89 81 90
rect 79 89 80 90
rect 78 89 79 90
rect 77 89 78 90
rect 76 89 77 90
rect 75 89 76 90
rect 74 89 75 90
rect 73 89 74 90
rect 72 89 73 90
rect 71 89 72 90
rect 70 89 71 90
rect 69 89 70 90
rect 68 89 69 90
rect 67 89 68 90
rect 66 89 67 90
rect 65 89 66 90
rect 64 89 65 90
rect 63 89 64 90
rect 62 89 63 90
rect 61 89 62 90
rect 60 89 61 90
rect 481 90 482 91
rect 480 90 481 91
rect 479 90 480 91
rect 478 90 479 91
rect 460 90 461 91
rect 399 90 400 91
rect 398 90 399 91
rect 397 90 398 91
rect 396 90 397 91
rect 395 90 396 91
rect 248 90 249 91
rect 247 90 248 91
rect 246 90 247 91
rect 245 90 246 91
rect 244 90 245 91
rect 243 90 244 91
rect 242 90 243 91
rect 241 90 242 91
rect 240 90 241 91
rect 239 90 240 91
rect 238 90 239 91
rect 237 90 238 91
rect 236 90 237 91
rect 235 90 236 91
rect 234 90 235 91
rect 233 90 234 91
rect 232 90 233 91
rect 231 90 232 91
rect 230 90 231 91
rect 229 90 230 91
rect 228 90 229 91
rect 227 90 228 91
rect 226 90 227 91
rect 225 90 226 91
rect 224 90 225 91
rect 223 90 224 91
rect 222 90 223 91
rect 221 90 222 91
rect 220 90 221 91
rect 219 90 220 91
rect 218 90 219 91
rect 217 90 218 91
rect 216 90 217 91
rect 215 90 216 91
rect 214 90 215 91
rect 213 90 214 91
rect 212 90 213 91
rect 211 90 212 91
rect 210 90 211 91
rect 209 90 210 91
rect 208 90 209 91
rect 207 90 208 91
rect 206 90 207 91
rect 205 90 206 91
rect 204 90 205 91
rect 203 90 204 91
rect 202 90 203 91
rect 201 90 202 91
rect 200 90 201 91
rect 199 90 200 91
rect 198 90 199 91
rect 197 90 198 91
rect 196 90 197 91
rect 195 90 196 91
rect 194 90 195 91
rect 193 90 194 91
rect 192 90 193 91
rect 191 90 192 91
rect 190 90 191 91
rect 161 90 162 91
rect 160 90 161 91
rect 159 90 160 91
rect 158 90 159 91
rect 157 90 158 91
rect 156 90 157 91
rect 155 90 156 91
rect 154 90 155 91
rect 153 90 154 91
rect 152 90 153 91
rect 151 90 152 91
rect 150 90 151 91
rect 149 90 150 91
rect 148 90 149 91
rect 147 90 148 91
rect 146 90 147 91
rect 145 90 146 91
rect 144 90 145 91
rect 143 90 144 91
rect 142 90 143 91
rect 141 90 142 91
rect 140 90 141 91
rect 139 90 140 91
rect 138 90 139 91
rect 137 90 138 91
rect 136 90 137 91
rect 135 90 136 91
rect 134 90 135 91
rect 133 90 134 91
rect 132 90 133 91
rect 131 90 132 91
rect 130 90 131 91
rect 123 90 124 91
rect 122 90 123 91
rect 121 90 122 91
rect 120 90 121 91
rect 119 90 120 91
rect 118 90 119 91
rect 117 90 118 91
rect 116 90 117 91
rect 115 90 116 91
rect 114 90 115 91
rect 113 90 114 91
rect 112 90 113 91
rect 111 90 112 91
rect 110 90 111 91
rect 109 90 110 91
rect 108 90 109 91
rect 107 90 108 91
rect 106 90 107 91
rect 105 90 106 91
rect 104 90 105 91
rect 103 90 104 91
rect 102 90 103 91
rect 101 90 102 91
rect 100 90 101 91
rect 99 90 100 91
rect 98 90 99 91
rect 97 90 98 91
rect 96 90 97 91
rect 95 90 96 91
rect 94 90 95 91
rect 93 90 94 91
rect 92 90 93 91
rect 91 90 92 91
rect 90 90 91 91
rect 89 90 90 91
rect 88 90 89 91
rect 87 90 88 91
rect 86 90 87 91
rect 85 90 86 91
rect 84 90 85 91
rect 83 90 84 91
rect 82 90 83 91
rect 81 90 82 91
rect 80 90 81 91
rect 79 90 80 91
rect 78 90 79 91
rect 77 90 78 91
rect 76 90 77 91
rect 75 90 76 91
rect 74 90 75 91
rect 73 90 74 91
rect 72 90 73 91
rect 71 90 72 91
rect 70 90 71 91
rect 69 90 70 91
rect 68 90 69 91
rect 67 90 68 91
rect 66 90 67 91
rect 65 90 66 91
rect 64 90 65 91
rect 63 90 64 91
rect 62 90 63 91
rect 61 90 62 91
rect 60 90 61 91
rect 59 90 60 91
rect 481 91 482 92
rect 480 91 481 92
rect 479 91 480 92
rect 398 91 399 92
rect 397 91 398 92
rect 396 91 397 92
rect 395 91 396 92
rect 250 91 251 92
rect 249 91 250 92
rect 248 91 249 92
rect 247 91 248 92
rect 246 91 247 92
rect 245 91 246 92
rect 244 91 245 92
rect 243 91 244 92
rect 242 91 243 92
rect 241 91 242 92
rect 240 91 241 92
rect 239 91 240 92
rect 238 91 239 92
rect 237 91 238 92
rect 236 91 237 92
rect 235 91 236 92
rect 234 91 235 92
rect 233 91 234 92
rect 232 91 233 92
rect 231 91 232 92
rect 230 91 231 92
rect 229 91 230 92
rect 228 91 229 92
rect 227 91 228 92
rect 226 91 227 92
rect 225 91 226 92
rect 224 91 225 92
rect 223 91 224 92
rect 222 91 223 92
rect 221 91 222 92
rect 220 91 221 92
rect 219 91 220 92
rect 218 91 219 92
rect 217 91 218 92
rect 216 91 217 92
rect 215 91 216 92
rect 214 91 215 92
rect 213 91 214 92
rect 212 91 213 92
rect 211 91 212 92
rect 210 91 211 92
rect 209 91 210 92
rect 208 91 209 92
rect 207 91 208 92
rect 206 91 207 92
rect 205 91 206 92
rect 204 91 205 92
rect 203 91 204 92
rect 202 91 203 92
rect 201 91 202 92
rect 200 91 201 92
rect 199 91 200 92
rect 198 91 199 92
rect 197 91 198 92
rect 196 91 197 92
rect 195 91 196 92
rect 194 91 195 92
rect 193 91 194 92
rect 192 91 193 92
rect 191 91 192 92
rect 190 91 191 92
rect 189 91 190 92
rect 161 91 162 92
rect 160 91 161 92
rect 159 91 160 92
rect 158 91 159 92
rect 157 91 158 92
rect 156 91 157 92
rect 155 91 156 92
rect 154 91 155 92
rect 153 91 154 92
rect 152 91 153 92
rect 151 91 152 92
rect 150 91 151 92
rect 149 91 150 92
rect 148 91 149 92
rect 147 91 148 92
rect 146 91 147 92
rect 145 91 146 92
rect 144 91 145 92
rect 143 91 144 92
rect 142 91 143 92
rect 141 91 142 92
rect 140 91 141 92
rect 139 91 140 92
rect 138 91 139 92
rect 137 91 138 92
rect 136 91 137 92
rect 135 91 136 92
rect 134 91 135 92
rect 133 91 134 92
rect 132 91 133 92
rect 131 91 132 92
rect 130 91 131 92
rect 123 91 124 92
rect 122 91 123 92
rect 121 91 122 92
rect 120 91 121 92
rect 119 91 120 92
rect 118 91 119 92
rect 117 91 118 92
rect 116 91 117 92
rect 115 91 116 92
rect 114 91 115 92
rect 113 91 114 92
rect 112 91 113 92
rect 111 91 112 92
rect 110 91 111 92
rect 109 91 110 92
rect 108 91 109 92
rect 107 91 108 92
rect 106 91 107 92
rect 105 91 106 92
rect 104 91 105 92
rect 103 91 104 92
rect 102 91 103 92
rect 101 91 102 92
rect 100 91 101 92
rect 99 91 100 92
rect 98 91 99 92
rect 97 91 98 92
rect 96 91 97 92
rect 95 91 96 92
rect 94 91 95 92
rect 93 91 94 92
rect 92 91 93 92
rect 91 91 92 92
rect 90 91 91 92
rect 89 91 90 92
rect 88 91 89 92
rect 87 91 88 92
rect 86 91 87 92
rect 85 91 86 92
rect 84 91 85 92
rect 83 91 84 92
rect 82 91 83 92
rect 81 91 82 92
rect 80 91 81 92
rect 79 91 80 92
rect 78 91 79 92
rect 77 91 78 92
rect 76 91 77 92
rect 75 91 76 92
rect 74 91 75 92
rect 73 91 74 92
rect 72 91 73 92
rect 71 91 72 92
rect 70 91 71 92
rect 69 91 70 92
rect 68 91 69 92
rect 67 91 68 92
rect 66 91 67 92
rect 65 91 66 92
rect 64 91 65 92
rect 63 91 64 92
rect 62 91 63 92
rect 61 91 62 92
rect 60 91 61 92
rect 59 91 60 92
rect 58 91 59 92
rect 481 92 482 93
rect 480 92 481 93
rect 479 92 480 93
rect 398 92 399 93
rect 397 92 398 93
rect 396 92 397 93
rect 395 92 396 93
rect 252 92 253 93
rect 251 92 252 93
rect 250 92 251 93
rect 249 92 250 93
rect 248 92 249 93
rect 247 92 248 93
rect 246 92 247 93
rect 245 92 246 93
rect 244 92 245 93
rect 243 92 244 93
rect 242 92 243 93
rect 241 92 242 93
rect 240 92 241 93
rect 239 92 240 93
rect 238 92 239 93
rect 237 92 238 93
rect 236 92 237 93
rect 235 92 236 93
rect 234 92 235 93
rect 233 92 234 93
rect 232 92 233 93
rect 231 92 232 93
rect 230 92 231 93
rect 229 92 230 93
rect 228 92 229 93
rect 227 92 228 93
rect 226 92 227 93
rect 225 92 226 93
rect 224 92 225 93
rect 223 92 224 93
rect 222 92 223 93
rect 221 92 222 93
rect 220 92 221 93
rect 219 92 220 93
rect 218 92 219 93
rect 217 92 218 93
rect 216 92 217 93
rect 215 92 216 93
rect 214 92 215 93
rect 213 92 214 93
rect 212 92 213 93
rect 211 92 212 93
rect 210 92 211 93
rect 209 92 210 93
rect 208 92 209 93
rect 207 92 208 93
rect 206 92 207 93
rect 205 92 206 93
rect 204 92 205 93
rect 203 92 204 93
rect 202 92 203 93
rect 201 92 202 93
rect 200 92 201 93
rect 199 92 200 93
rect 198 92 199 93
rect 197 92 198 93
rect 196 92 197 93
rect 195 92 196 93
rect 194 92 195 93
rect 193 92 194 93
rect 192 92 193 93
rect 191 92 192 93
rect 190 92 191 93
rect 189 92 190 93
rect 188 92 189 93
rect 187 92 188 93
rect 161 92 162 93
rect 160 92 161 93
rect 159 92 160 93
rect 158 92 159 93
rect 157 92 158 93
rect 156 92 157 93
rect 155 92 156 93
rect 154 92 155 93
rect 153 92 154 93
rect 152 92 153 93
rect 151 92 152 93
rect 150 92 151 93
rect 149 92 150 93
rect 148 92 149 93
rect 147 92 148 93
rect 146 92 147 93
rect 145 92 146 93
rect 144 92 145 93
rect 143 92 144 93
rect 142 92 143 93
rect 141 92 142 93
rect 140 92 141 93
rect 139 92 140 93
rect 138 92 139 93
rect 137 92 138 93
rect 136 92 137 93
rect 135 92 136 93
rect 134 92 135 93
rect 133 92 134 93
rect 132 92 133 93
rect 131 92 132 93
rect 130 92 131 93
rect 122 92 123 93
rect 121 92 122 93
rect 120 92 121 93
rect 119 92 120 93
rect 118 92 119 93
rect 117 92 118 93
rect 116 92 117 93
rect 115 92 116 93
rect 114 92 115 93
rect 113 92 114 93
rect 112 92 113 93
rect 111 92 112 93
rect 110 92 111 93
rect 109 92 110 93
rect 108 92 109 93
rect 107 92 108 93
rect 106 92 107 93
rect 105 92 106 93
rect 104 92 105 93
rect 103 92 104 93
rect 102 92 103 93
rect 101 92 102 93
rect 100 92 101 93
rect 99 92 100 93
rect 98 92 99 93
rect 97 92 98 93
rect 96 92 97 93
rect 95 92 96 93
rect 94 92 95 93
rect 93 92 94 93
rect 92 92 93 93
rect 91 92 92 93
rect 90 92 91 93
rect 89 92 90 93
rect 88 92 89 93
rect 87 92 88 93
rect 86 92 87 93
rect 85 92 86 93
rect 84 92 85 93
rect 83 92 84 93
rect 82 92 83 93
rect 81 92 82 93
rect 80 92 81 93
rect 79 92 80 93
rect 78 92 79 93
rect 77 92 78 93
rect 76 92 77 93
rect 75 92 76 93
rect 74 92 75 93
rect 73 92 74 93
rect 72 92 73 93
rect 71 92 72 93
rect 70 92 71 93
rect 69 92 70 93
rect 68 92 69 93
rect 67 92 68 93
rect 66 92 67 93
rect 65 92 66 93
rect 64 92 65 93
rect 63 92 64 93
rect 62 92 63 93
rect 61 92 62 93
rect 60 92 61 93
rect 59 92 60 93
rect 58 92 59 93
rect 481 93 482 94
rect 480 93 481 94
rect 397 93 398 94
rect 396 93 397 94
rect 395 93 396 94
rect 254 93 255 94
rect 253 93 254 94
rect 252 93 253 94
rect 251 93 252 94
rect 250 93 251 94
rect 249 93 250 94
rect 248 93 249 94
rect 247 93 248 94
rect 246 93 247 94
rect 245 93 246 94
rect 244 93 245 94
rect 243 93 244 94
rect 242 93 243 94
rect 241 93 242 94
rect 240 93 241 94
rect 239 93 240 94
rect 238 93 239 94
rect 237 93 238 94
rect 236 93 237 94
rect 235 93 236 94
rect 234 93 235 94
rect 233 93 234 94
rect 232 93 233 94
rect 231 93 232 94
rect 230 93 231 94
rect 229 93 230 94
rect 228 93 229 94
rect 227 93 228 94
rect 226 93 227 94
rect 225 93 226 94
rect 224 93 225 94
rect 223 93 224 94
rect 222 93 223 94
rect 221 93 222 94
rect 220 93 221 94
rect 219 93 220 94
rect 218 93 219 94
rect 217 93 218 94
rect 216 93 217 94
rect 215 93 216 94
rect 214 93 215 94
rect 213 93 214 94
rect 212 93 213 94
rect 211 93 212 94
rect 210 93 211 94
rect 209 93 210 94
rect 208 93 209 94
rect 207 93 208 94
rect 206 93 207 94
rect 205 93 206 94
rect 204 93 205 94
rect 203 93 204 94
rect 202 93 203 94
rect 201 93 202 94
rect 200 93 201 94
rect 199 93 200 94
rect 198 93 199 94
rect 197 93 198 94
rect 196 93 197 94
rect 195 93 196 94
rect 194 93 195 94
rect 193 93 194 94
rect 192 93 193 94
rect 191 93 192 94
rect 190 93 191 94
rect 189 93 190 94
rect 188 93 189 94
rect 187 93 188 94
rect 186 93 187 94
rect 160 93 161 94
rect 159 93 160 94
rect 158 93 159 94
rect 157 93 158 94
rect 156 93 157 94
rect 155 93 156 94
rect 154 93 155 94
rect 153 93 154 94
rect 152 93 153 94
rect 151 93 152 94
rect 150 93 151 94
rect 149 93 150 94
rect 148 93 149 94
rect 147 93 148 94
rect 146 93 147 94
rect 145 93 146 94
rect 144 93 145 94
rect 143 93 144 94
rect 142 93 143 94
rect 141 93 142 94
rect 140 93 141 94
rect 139 93 140 94
rect 138 93 139 94
rect 137 93 138 94
rect 136 93 137 94
rect 135 93 136 94
rect 134 93 135 94
rect 133 93 134 94
rect 132 93 133 94
rect 131 93 132 94
rect 130 93 131 94
rect 129 93 130 94
rect 122 93 123 94
rect 121 93 122 94
rect 120 93 121 94
rect 119 93 120 94
rect 118 93 119 94
rect 117 93 118 94
rect 116 93 117 94
rect 115 93 116 94
rect 114 93 115 94
rect 113 93 114 94
rect 112 93 113 94
rect 111 93 112 94
rect 110 93 111 94
rect 109 93 110 94
rect 108 93 109 94
rect 107 93 108 94
rect 106 93 107 94
rect 105 93 106 94
rect 104 93 105 94
rect 103 93 104 94
rect 102 93 103 94
rect 101 93 102 94
rect 100 93 101 94
rect 99 93 100 94
rect 98 93 99 94
rect 97 93 98 94
rect 96 93 97 94
rect 95 93 96 94
rect 94 93 95 94
rect 93 93 94 94
rect 92 93 93 94
rect 91 93 92 94
rect 90 93 91 94
rect 89 93 90 94
rect 88 93 89 94
rect 87 93 88 94
rect 86 93 87 94
rect 85 93 86 94
rect 84 93 85 94
rect 83 93 84 94
rect 82 93 83 94
rect 81 93 82 94
rect 80 93 81 94
rect 79 93 80 94
rect 78 93 79 94
rect 77 93 78 94
rect 76 93 77 94
rect 75 93 76 94
rect 74 93 75 94
rect 73 93 74 94
rect 72 93 73 94
rect 71 93 72 94
rect 70 93 71 94
rect 69 93 70 94
rect 68 93 69 94
rect 67 93 68 94
rect 66 93 67 94
rect 65 93 66 94
rect 64 93 65 94
rect 63 93 64 94
rect 62 93 63 94
rect 61 93 62 94
rect 60 93 61 94
rect 59 93 60 94
rect 58 93 59 94
rect 57 93 58 94
rect 481 94 482 95
rect 480 94 481 95
rect 397 94 398 95
rect 396 94 397 95
rect 395 94 396 95
rect 255 94 256 95
rect 254 94 255 95
rect 253 94 254 95
rect 252 94 253 95
rect 251 94 252 95
rect 250 94 251 95
rect 249 94 250 95
rect 248 94 249 95
rect 247 94 248 95
rect 246 94 247 95
rect 245 94 246 95
rect 244 94 245 95
rect 243 94 244 95
rect 242 94 243 95
rect 241 94 242 95
rect 240 94 241 95
rect 239 94 240 95
rect 238 94 239 95
rect 237 94 238 95
rect 236 94 237 95
rect 235 94 236 95
rect 234 94 235 95
rect 233 94 234 95
rect 232 94 233 95
rect 231 94 232 95
rect 230 94 231 95
rect 229 94 230 95
rect 228 94 229 95
rect 227 94 228 95
rect 226 94 227 95
rect 225 94 226 95
rect 224 94 225 95
rect 223 94 224 95
rect 222 94 223 95
rect 221 94 222 95
rect 220 94 221 95
rect 219 94 220 95
rect 218 94 219 95
rect 217 94 218 95
rect 216 94 217 95
rect 215 94 216 95
rect 214 94 215 95
rect 213 94 214 95
rect 212 94 213 95
rect 211 94 212 95
rect 210 94 211 95
rect 209 94 210 95
rect 208 94 209 95
rect 207 94 208 95
rect 206 94 207 95
rect 205 94 206 95
rect 204 94 205 95
rect 203 94 204 95
rect 202 94 203 95
rect 201 94 202 95
rect 200 94 201 95
rect 199 94 200 95
rect 198 94 199 95
rect 197 94 198 95
rect 196 94 197 95
rect 195 94 196 95
rect 194 94 195 95
rect 193 94 194 95
rect 192 94 193 95
rect 191 94 192 95
rect 190 94 191 95
rect 189 94 190 95
rect 188 94 189 95
rect 187 94 188 95
rect 186 94 187 95
rect 185 94 186 95
rect 160 94 161 95
rect 159 94 160 95
rect 158 94 159 95
rect 157 94 158 95
rect 156 94 157 95
rect 155 94 156 95
rect 154 94 155 95
rect 153 94 154 95
rect 152 94 153 95
rect 151 94 152 95
rect 150 94 151 95
rect 149 94 150 95
rect 148 94 149 95
rect 147 94 148 95
rect 146 94 147 95
rect 145 94 146 95
rect 144 94 145 95
rect 143 94 144 95
rect 142 94 143 95
rect 141 94 142 95
rect 140 94 141 95
rect 139 94 140 95
rect 138 94 139 95
rect 137 94 138 95
rect 136 94 137 95
rect 135 94 136 95
rect 134 94 135 95
rect 133 94 134 95
rect 132 94 133 95
rect 131 94 132 95
rect 130 94 131 95
rect 129 94 130 95
rect 122 94 123 95
rect 121 94 122 95
rect 120 94 121 95
rect 119 94 120 95
rect 118 94 119 95
rect 117 94 118 95
rect 116 94 117 95
rect 115 94 116 95
rect 114 94 115 95
rect 113 94 114 95
rect 112 94 113 95
rect 111 94 112 95
rect 110 94 111 95
rect 109 94 110 95
rect 108 94 109 95
rect 107 94 108 95
rect 106 94 107 95
rect 105 94 106 95
rect 104 94 105 95
rect 103 94 104 95
rect 102 94 103 95
rect 101 94 102 95
rect 100 94 101 95
rect 99 94 100 95
rect 98 94 99 95
rect 97 94 98 95
rect 96 94 97 95
rect 95 94 96 95
rect 94 94 95 95
rect 93 94 94 95
rect 92 94 93 95
rect 91 94 92 95
rect 90 94 91 95
rect 89 94 90 95
rect 88 94 89 95
rect 87 94 88 95
rect 86 94 87 95
rect 85 94 86 95
rect 84 94 85 95
rect 83 94 84 95
rect 82 94 83 95
rect 81 94 82 95
rect 80 94 81 95
rect 79 94 80 95
rect 78 94 79 95
rect 77 94 78 95
rect 76 94 77 95
rect 75 94 76 95
rect 74 94 75 95
rect 73 94 74 95
rect 72 94 73 95
rect 71 94 72 95
rect 70 94 71 95
rect 69 94 70 95
rect 68 94 69 95
rect 67 94 68 95
rect 66 94 67 95
rect 65 94 66 95
rect 64 94 65 95
rect 63 94 64 95
rect 62 94 63 95
rect 61 94 62 95
rect 60 94 61 95
rect 59 94 60 95
rect 58 94 59 95
rect 57 94 58 95
rect 56 94 57 95
rect 481 95 482 96
rect 480 95 481 96
rect 479 95 480 96
rect 397 95 398 96
rect 396 95 397 96
rect 395 95 396 96
rect 257 95 258 96
rect 256 95 257 96
rect 255 95 256 96
rect 254 95 255 96
rect 253 95 254 96
rect 252 95 253 96
rect 251 95 252 96
rect 250 95 251 96
rect 249 95 250 96
rect 248 95 249 96
rect 247 95 248 96
rect 246 95 247 96
rect 245 95 246 96
rect 244 95 245 96
rect 243 95 244 96
rect 242 95 243 96
rect 241 95 242 96
rect 240 95 241 96
rect 239 95 240 96
rect 238 95 239 96
rect 237 95 238 96
rect 236 95 237 96
rect 235 95 236 96
rect 234 95 235 96
rect 233 95 234 96
rect 232 95 233 96
rect 231 95 232 96
rect 230 95 231 96
rect 229 95 230 96
rect 228 95 229 96
rect 227 95 228 96
rect 226 95 227 96
rect 225 95 226 96
rect 224 95 225 96
rect 223 95 224 96
rect 222 95 223 96
rect 221 95 222 96
rect 220 95 221 96
rect 219 95 220 96
rect 218 95 219 96
rect 217 95 218 96
rect 216 95 217 96
rect 215 95 216 96
rect 214 95 215 96
rect 213 95 214 96
rect 212 95 213 96
rect 211 95 212 96
rect 210 95 211 96
rect 209 95 210 96
rect 208 95 209 96
rect 207 95 208 96
rect 206 95 207 96
rect 205 95 206 96
rect 204 95 205 96
rect 203 95 204 96
rect 202 95 203 96
rect 201 95 202 96
rect 200 95 201 96
rect 199 95 200 96
rect 198 95 199 96
rect 197 95 198 96
rect 196 95 197 96
rect 195 95 196 96
rect 194 95 195 96
rect 193 95 194 96
rect 192 95 193 96
rect 191 95 192 96
rect 190 95 191 96
rect 189 95 190 96
rect 188 95 189 96
rect 187 95 188 96
rect 186 95 187 96
rect 185 95 186 96
rect 184 95 185 96
rect 160 95 161 96
rect 159 95 160 96
rect 158 95 159 96
rect 157 95 158 96
rect 156 95 157 96
rect 155 95 156 96
rect 154 95 155 96
rect 153 95 154 96
rect 152 95 153 96
rect 151 95 152 96
rect 150 95 151 96
rect 149 95 150 96
rect 148 95 149 96
rect 147 95 148 96
rect 146 95 147 96
rect 145 95 146 96
rect 144 95 145 96
rect 143 95 144 96
rect 142 95 143 96
rect 141 95 142 96
rect 140 95 141 96
rect 139 95 140 96
rect 138 95 139 96
rect 137 95 138 96
rect 136 95 137 96
rect 135 95 136 96
rect 134 95 135 96
rect 133 95 134 96
rect 132 95 133 96
rect 131 95 132 96
rect 130 95 131 96
rect 129 95 130 96
rect 122 95 123 96
rect 121 95 122 96
rect 120 95 121 96
rect 119 95 120 96
rect 118 95 119 96
rect 117 95 118 96
rect 116 95 117 96
rect 115 95 116 96
rect 114 95 115 96
rect 113 95 114 96
rect 112 95 113 96
rect 111 95 112 96
rect 110 95 111 96
rect 109 95 110 96
rect 108 95 109 96
rect 107 95 108 96
rect 106 95 107 96
rect 105 95 106 96
rect 104 95 105 96
rect 103 95 104 96
rect 102 95 103 96
rect 101 95 102 96
rect 100 95 101 96
rect 99 95 100 96
rect 98 95 99 96
rect 97 95 98 96
rect 96 95 97 96
rect 95 95 96 96
rect 94 95 95 96
rect 93 95 94 96
rect 92 95 93 96
rect 91 95 92 96
rect 90 95 91 96
rect 89 95 90 96
rect 88 95 89 96
rect 87 95 88 96
rect 86 95 87 96
rect 85 95 86 96
rect 84 95 85 96
rect 83 95 84 96
rect 82 95 83 96
rect 81 95 82 96
rect 80 95 81 96
rect 79 95 80 96
rect 78 95 79 96
rect 77 95 78 96
rect 76 95 77 96
rect 75 95 76 96
rect 74 95 75 96
rect 73 95 74 96
rect 72 95 73 96
rect 71 95 72 96
rect 70 95 71 96
rect 69 95 70 96
rect 68 95 69 96
rect 67 95 68 96
rect 66 95 67 96
rect 65 95 66 96
rect 64 95 65 96
rect 63 95 64 96
rect 62 95 63 96
rect 61 95 62 96
rect 60 95 61 96
rect 59 95 60 96
rect 58 95 59 96
rect 57 95 58 96
rect 56 95 57 96
rect 55 95 56 96
rect 480 96 481 97
rect 479 96 480 97
rect 460 96 461 97
rect 259 96 260 97
rect 258 96 259 97
rect 257 96 258 97
rect 256 96 257 97
rect 255 96 256 97
rect 254 96 255 97
rect 253 96 254 97
rect 252 96 253 97
rect 251 96 252 97
rect 250 96 251 97
rect 249 96 250 97
rect 248 96 249 97
rect 247 96 248 97
rect 246 96 247 97
rect 245 96 246 97
rect 244 96 245 97
rect 243 96 244 97
rect 242 96 243 97
rect 241 96 242 97
rect 240 96 241 97
rect 239 96 240 97
rect 238 96 239 97
rect 237 96 238 97
rect 236 96 237 97
rect 235 96 236 97
rect 234 96 235 97
rect 233 96 234 97
rect 232 96 233 97
rect 231 96 232 97
rect 230 96 231 97
rect 229 96 230 97
rect 228 96 229 97
rect 227 96 228 97
rect 226 96 227 97
rect 225 96 226 97
rect 224 96 225 97
rect 223 96 224 97
rect 222 96 223 97
rect 221 96 222 97
rect 220 96 221 97
rect 219 96 220 97
rect 218 96 219 97
rect 217 96 218 97
rect 216 96 217 97
rect 215 96 216 97
rect 214 96 215 97
rect 213 96 214 97
rect 212 96 213 97
rect 211 96 212 97
rect 210 96 211 97
rect 209 96 210 97
rect 208 96 209 97
rect 207 96 208 97
rect 206 96 207 97
rect 205 96 206 97
rect 204 96 205 97
rect 203 96 204 97
rect 202 96 203 97
rect 201 96 202 97
rect 200 96 201 97
rect 199 96 200 97
rect 198 96 199 97
rect 197 96 198 97
rect 196 96 197 97
rect 195 96 196 97
rect 194 96 195 97
rect 193 96 194 97
rect 192 96 193 97
rect 191 96 192 97
rect 190 96 191 97
rect 189 96 190 97
rect 188 96 189 97
rect 187 96 188 97
rect 186 96 187 97
rect 185 96 186 97
rect 184 96 185 97
rect 183 96 184 97
rect 159 96 160 97
rect 158 96 159 97
rect 157 96 158 97
rect 156 96 157 97
rect 155 96 156 97
rect 154 96 155 97
rect 153 96 154 97
rect 152 96 153 97
rect 151 96 152 97
rect 150 96 151 97
rect 149 96 150 97
rect 148 96 149 97
rect 147 96 148 97
rect 146 96 147 97
rect 145 96 146 97
rect 144 96 145 97
rect 143 96 144 97
rect 142 96 143 97
rect 141 96 142 97
rect 140 96 141 97
rect 139 96 140 97
rect 138 96 139 97
rect 137 96 138 97
rect 136 96 137 97
rect 135 96 136 97
rect 134 96 135 97
rect 133 96 134 97
rect 132 96 133 97
rect 131 96 132 97
rect 130 96 131 97
rect 129 96 130 97
rect 121 96 122 97
rect 120 96 121 97
rect 119 96 120 97
rect 118 96 119 97
rect 117 96 118 97
rect 116 96 117 97
rect 115 96 116 97
rect 114 96 115 97
rect 113 96 114 97
rect 112 96 113 97
rect 111 96 112 97
rect 110 96 111 97
rect 109 96 110 97
rect 108 96 109 97
rect 107 96 108 97
rect 106 96 107 97
rect 105 96 106 97
rect 104 96 105 97
rect 103 96 104 97
rect 102 96 103 97
rect 101 96 102 97
rect 100 96 101 97
rect 99 96 100 97
rect 98 96 99 97
rect 97 96 98 97
rect 96 96 97 97
rect 95 96 96 97
rect 94 96 95 97
rect 93 96 94 97
rect 92 96 93 97
rect 91 96 92 97
rect 90 96 91 97
rect 89 96 90 97
rect 88 96 89 97
rect 87 96 88 97
rect 86 96 87 97
rect 85 96 86 97
rect 84 96 85 97
rect 83 96 84 97
rect 82 96 83 97
rect 81 96 82 97
rect 80 96 81 97
rect 79 96 80 97
rect 78 96 79 97
rect 77 96 78 97
rect 76 96 77 97
rect 75 96 76 97
rect 74 96 75 97
rect 73 96 74 97
rect 72 96 73 97
rect 71 96 72 97
rect 70 96 71 97
rect 69 96 70 97
rect 68 96 69 97
rect 67 96 68 97
rect 66 96 67 97
rect 65 96 66 97
rect 64 96 65 97
rect 63 96 64 97
rect 62 96 63 97
rect 61 96 62 97
rect 60 96 61 97
rect 59 96 60 97
rect 58 96 59 97
rect 57 96 58 97
rect 56 96 57 97
rect 55 96 56 97
rect 54 96 55 97
rect 480 97 481 98
rect 479 97 480 98
rect 478 97 479 98
rect 460 97 461 98
rect 260 97 261 98
rect 259 97 260 98
rect 258 97 259 98
rect 257 97 258 98
rect 256 97 257 98
rect 255 97 256 98
rect 254 97 255 98
rect 253 97 254 98
rect 252 97 253 98
rect 251 97 252 98
rect 250 97 251 98
rect 249 97 250 98
rect 248 97 249 98
rect 247 97 248 98
rect 246 97 247 98
rect 245 97 246 98
rect 244 97 245 98
rect 243 97 244 98
rect 242 97 243 98
rect 241 97 242 98
rect 240 97 241 98
rect 239 97 240 98
rect 238 97 239 98
rect 237 97 238 98
rect 236 97 237 98
rect 235 97 236 98
rect 234 97 235 98
rect 233 97 234 98
rect 232 97 233 98
rect 231 97 232 98
rect 230 97 231 98
rect 229 97 230 98
rect 228 97 229 98
rect 227 97 228 98
rect 226 97 227 98
rect 225 97 226 98
rect 224 97 225 98
rect 223 97 224 98
rect 222 97 223 98
rect 221 97 222 98
rect 220 97 221 98
rect 219 97 220 98
rect 218 97 219 98
rect 217 97 218 98
rect 216 97 217 98
rect 215 97 216 98
rect 214 97 215 98
rect 213 97 214 98
rect 212 97 213 98
rect 211 97 212 98
rect 210 97 211 98
rect 209 97 210 98
rect 208 97 209 98
rect 207 97 208 98
rect 206 97 207 98
rect 205 97 206 98
rect 204 97 205 98
rect 203 97 204 98
rect 202 97 203 98
rect 201 97 202 98
rect 200 97 201 98
rect 199 97 200 98
rect 198 97 199 98
rect 197 97 198 98
rect 196 97 197 98
rect 195 97 196 98
rect 194 97 195 98
rect 193 97 194 98
rect 192 97 193 98
rect 191 97 192 98
rect 190 97 191 98
rect 189 97 190 98
rect 188 97 189 98
rect 187 97 188 98
rect 186 97 187 98
rect 185 97 186 98
rect 184 97 185 98
rect 183 97 184 98
rect 182 97 183 98
rect 159 97 160 98
rect 158 97 159 98
rect 157 97 158 98
rect 156 97 157 98
rect 155 97 156 98
rect 154 97 155 98
rect 153 97 154 98
rect 152 97 153 98
rect 151 97 152 98
rect 150 97 151 98
rect 149 97 150 98
rect 148 97 149 98
rect 147 97 148 98
rect 146 97 147 98
rect 145 97 146 98
rect 144 97 145 98
rect 143 97 144 98
rect 142 97 143 98
rect 141 97 142 98
rect 140 97 141 98
rect 139 97 140 98
rect 138 97 139 98
rect 137 97 138 98
rect 136 97 137 98
rect 135 97 136 98
rect 134 97 135 98
rect 133 97 134 98
rect 132 97 133 98
rect 131 97 132 98
rect 130 97 131 98
rect 129 97 130 98
rect 121 97 122 98
rect 120 97 121 98
rect 119 97 120 98
rect 118 97 119 98
rect 117 97 118 98
rect 116 97 117 98
rect 115 97 116 98
rect 114 97 115 98
rect 113 97 114 98
rect 112 97 113 98
rect 111 97 112 98
rect 110 97 111 98
rect 109 97 110 98
rect 108 97 109 98
rect 107 97 108 98
rect 106 97 107 98
rect 105 97 106 98
rect 104 97 105 98
rect 103 97 104 98
rect 102 97 103 98
rect 101 97 102 98
rect 100 97 101 98
rect 99 97 100 98
rect 98 97 99 98
rect 97 97 98 98
rect 96 97 97 98
rect 95 97 96 98
rect 94 97 95 98
rect 93 97 94 98
rect 92 97 93 98
rect 91 97 92 98
rect 90 97 91 98
rect 89 97 90 98
rect 88 97 89 98
rect 87 97 88 98
rect 86 97 87 98
rect 85 97 86 98
rect 84 97 85 98
rect 83 97 84 98
rect 82 97 83 98
rect 81 97 82 98
rect 80 97 81 98
rect 79 97 80 98
rect 78 97 79 98
rect 77 97 78 98
rect 76 97 77 98
rect 75 97 76 98
rect 72 97 73 98
rect 71 97 72 98
rect 70 97 71 98
rect 69 97 70 98
rect 68 97 69 98
rect 67 97 68 98
rect 66 97 67 98
rect 65 97 66 98
rect 64 97 65 98
rect 63 97 64 98
rect 62 97 63 98
rect 61 97 62 98
rect 60 97 61 98
rect 59 97 60 98
rect 58 97 59 98
rect 57 97 58 98
rect 56 97 57 98
rect 55 97 56 98
rect 54 97 55 98
rect 53 97 54 98
rect 479 98 480 99
rect 478 98 479 99
rect 477 98 478 99
rect 461 98 462 99
rect 460 98 461 99
rect 262 98 263 99
rect 261 98 262 99
rect 260 98 261 99
rect 259 98 260 99
rect 258 98 259 99
rect 257 98 258 99
rect 256 98 257 99
rect 255 98 256 99
rect 254 98 255 99
rect 253 98 254 99
rect 252 98 253 99
rect 251 98 252 99
rect 250 98 251 99
rect 249 98 250 99
rect 248 98 249 99
rect 247 98 248 99
rect 246 98 247 99
rect 245 98 246 99
rect 244 98 245 99
rect 243 98 244 99
rect 242 98 243 99
rect 241 98 242 99
rect 240 98 241 99
rect 239 98 240 99
rect 238 98 239 99
rect 237 98 238 99
rect 236 98 237 99
rect 235 98 236 99
rect 234 98 235 99
rect 233 98 234 99
rect 232 98 233 99
rect 231 98 232 99
rect 230 98 231 99
rect 229 98 230 99
rect 228 98 229 99
rect 227 98 228 99
rect 226 98 227 99
rect 225 98 226 99
rect 224 98 225 99
rect 223 98 224 99
rect 222 98 223 99
rect 221 98 222 99
rect 220 98 221 99
rect 219 98 220 99
rect 218 98 219 99
rect 217 98 218 99
rect 216 98 217 99
rect 215 98 216 99
rect 214 98 215 99
rect 213 98 214 99
rect 212 98 213 99
rect 211 98 212 99
rect 210 98 211 99
rect 209 98 210 99
rect 208 98 209 99
rect 207 98 208 99
rect 206 98 207 99
rect 205 98 206 99
rect 204 98 205 99
rect 203 98 204 99
rect 202 98 203 99
rect 201 98 202 99
rect 200 98 201 99
rect 199 98 200 99
rect 198 98 199 99
rect 197 98 198 99
rect 196 98 197 99
rect 195 98 196 99
rect 194 98 195 99
rect 193 98 194 99
rect 192 98 193 99
rect 191 98 192 99
rect 190 98 191 99
rect 189 98 190 99
rect 188 98 189 99
rect 187 98 188 99
rect 186 98 187 99
rect 185 98 186 99
rect 184 98 185 99
rect 183 98 184 99
rect 182 98 183 99
rect 181 98 182 99
rect 159 98 160 99
rect 158 98 159 99
rect 157 98 158 99
rect 156 98 157 99
rect 155 98 156 99
rect 154 98 155 99
rect 153 98 154 99
rect 152 98 153 99
rect 151 98 152 99
rect 150 98 151 99
rect 149 98 150 99
rect 148 98 149 99
rect 147 98 148 99
rect 146 98 147 99
rect 145 98 146 99
rect 144 98 145 99
rect 143 98 144 99
rect 142 98 143 99
rect 141 98 142 99
rect 140 98 141 99
rect 139 98 140 99
rect 138 98 139 99
rect 137 98 138 99
rect 136 98 137 99
rect 135 98 136 99
rect 134 98 135 99
rect 133 98 134 99
rect 132 98 133 99
rect 131 98 132 99
rect 130 98 131 99
rect 129 98 130 99
rect 121 98 122 99
rect 120 98 121 99
rect 119 98 120 99
rect 118 98 119 99
rect 117 98 118 99
rect 116 98 117 99
rect 115 98 116 99
rect 114 98 115 99
rect 113 98 114 99
rect 112 98 113 99
rect 111 98 112 99
rect 110 98 111 99
rect 109 98 110 99
rect 108 98 109 99
rect 107 98 108 99
rect 106 98 107 99
rect 105 98 106 99
rect 104 98 105 99
rect 103 98 104 99
rect 102 98 103 99
rect 101 98 102 99
rect 100 98 101 99
rect 99 98 100 99
rect 98 98 99 99
rect 97 98 98 99
rect 96 98 97 99
rect 95 98 96 99
rect 94 98 95 99
rect 93 98 94 99
rect 92 98 93 99
rect 91 98 92 99
rect 90 98 91 99
rect 89 98 90 99
rect 88 98 89 99
rect 87 98 88 99
rect 86 98 87 99
rect 85 98 86 99
rect 84 98 85 99
rect 83 98 84 99
rect 82 98 83 99
rect 81 98 82 99
rect 80 98 81 99
rect 79 98 80 99
rect 78 98 79 99
rect 77 98 78 99
rect 76 98 77 99
rect 75 98 76 99
rect 71 98 72 99
rect 70 98 71 99
rect 69 98 70 99
rect 68 98 69 99
rect 67 98 68 99
rect 66 98 67 99
rect 65 98 66 99
rect 64 98 65 99
rect 63 98 64 99
rect 62 98 63 99
rect 61 98 62 99
rect 60 98 61 99
rect 59 98 60 99
rect 58 98 59 99
rect 57 98 58 99
rect 56 98 57 99
rect 55 98 56 99
rect 54 98 55 99
rect 53 98 54 99
rect 52 98 53 99
rect 478 99 479 100
rect 477 99 478 100
rect 476 99 477 100
rect 475 99 476 100
rect 474 99 475 100
rect 473 99 474 100
rect 472 99 473 100
rect 471 99 472 100
rect 470 99 471 100
rect 469 99 470 100
rect 468 99 469 100
rect 467 99 468 100
rect 466 99 467 100
rect 465 99 466 100
rect 464 99 465 100
rect 463 99 464 100
rect 462 99 463 100
rect 461 99 462 100
rect 460 99 461 100
rect 263 99 264 100
rect 262 99 263 100
rect 261 99 262 100
rect 260 99 261 100
rect 259 99 260 100
rect 258 99 259 100
rect 257 99 258 100
rect 256 99 257 100
rect 255 99 256 100
rect 254 99 255 100
rect 253 99 254 100
rect 252 99 253 100
rect 251 99 252 100
rect 250 99 251 100
rect 249 99 250 100
rect 248 99 249 100
rect 247 99 248 100
rect 246 99 247 100
rect 245 99 246 100
rect 244 99 245 100
rect 243 99 244 100
rect 242 99 243 100
rect 241 99 242 100
rect 240 99 241 100
rect 239 99 240 100
rect 238 99 239 100
rect 237 99 238 100
rect 236 99 237 100
rect 235 99 236 100
rect 234 99 235 100
rect 233 99 234 100
rect 232 99 233 100
rect 231 99 232 100
rect 230 99 231 100
rect 229 99 230 100
rect 228 99 229 100
rect 227 99 228 100
rect 226 99 227 100
rect 225 99 226 100
rect 224 99 225 100
rect 223 99 224 100
rect 222 99 223 100
rect 221 99 222 100
rect 220 99 221 100
rect 219 99 220 100
rect 218 99 219 100
rect 217 99 218 100
rect 216 99 217 100
rect 215 99 216 100
rect 214 99 215 100
rect 213 99 214 100
rect 212 99 213 100
rect 211 99 212 100
rect 210 99 211 100
rect 209 99 210 100
rect 208 99 209 100
rect 207 99 208 100
rect 206 99 207 100
rect 205 99 206 100
rect 204 99 205 100
rect 203 99 204 100
rect 202 99 203 100
rect 201 99 202 100
rect 200 99 201 100
rect 199 99 200 100
rect 198 99 199 100
rect 197 99 198 100
rect 196 99 197 100
rect 195 99 196 100
rect 194 99 195 100
rect 193 99 194 100
rect 192 99 193 100
rect 191 99 192 100
rect 190 99 191 100
rect 189 99 190 100
rect 188 99 189 100
rect 187 99 188 100
rect 186 99 187 100
rect 185 99 186 100
rect 184 99 185 100
rect 183 99 184 100
rect 182 99 183 100
rect 181 99 182 100
rect 180 99 181 100
rect 158 99 159 100
rect 157 99 158 100
rect 156 99 157 100
rect 155 99 156 100
rect 154 99 155 100
rect 153 99 154 100
rect 152 99 153 100
rect 151 99 152 100
rect 150 99 151 100
rect 149 99 150 100
rect 148 99 149 100
rect 147 99 148 100
rect 146 99 147 100
rect 145 99 146 100
rect 144 99 145 100
rect 143 99 144 100
rect 142 99 143 100
rect 141 99 142 100
rect 140 99 141 100
rect 139 99 140 100
rect 138 99 139 100
rect 137 99 138 100
rect 136 99 137 100
rect 135 99 136 100
rect 134 99 135 100
rect 133 99 134 100
rect 132 99 133 100
rect 131 99 132 100
rect 130 99 131 100
rect 129 99 130 100
rect 128 99 129 100
rect 120 99 121 100
rect 119 99 120 100
rect 118 99 119 100
rect 117 99 118 100
rect 116 99 117 100
rect 115 99 116 100
rect 114 99 115 100
rect 113 99 114 100
rect 112 99 113 100
rect 111 99 112 100
rect 110 99 111 100
rect 109 99 110 100
rect 108 99 109 100
rect 107 99 108 100
rect 106 99 107 100
rect 105 99 106 100
rect 104 99 105 100
rect 103 99 104 100
rect 102 99 103 100
rect 101 99 102 100
rect 100 99 101 100
rect 99 99 100 100
rect 98 99 99 100
rect 97 99 98 100
rect 96 99 97 100
rect 95 99 96 100
rect 94 99 95 100
rect 93 99 94 100
rect 92 99 93 100
rect 91 99 92 100
rect 90 99 91 100
rect 89 99 90 100
rect 88 99 89 100
rect 87 99 88 100
rect 86 99 87 100
rect 85 99 86 100
rect 84 99 85 100
rect 83 99 84 100
rect 82 99 83 100
rect 81 99 82 100
rect 80 99 81 100
rect 79 99 80 100
rect 78 99 79 100
rect 77 99 78 100
rect 76 99 77 100
rect 75 99 76 100
rect 74 99 75 100
rect 70 99 71 100
rect 69 99 70 100
rect 68 99 69 100
rect 67 99 68 100
rect 66 99 67 100
rect 65 99 66 100
rect 64 99 65 100
rect 63 99 64 100
rect 62 99 63 100
rect 61 99 62 100
rect 60 99 61 100
rect 59 99 60 100
rect 58 99 59 100
rect 57 99 58 100
rect 56 99 57 100
rect 55 99 56 100
rect 54 99 55 100
rect 53 99 54 100
rect 52 99 53 100
rect 51 99 52 100
rect 476 100 477 101
rect 475 100 476 101
rect 474 100 475 101
rect 473 100 474 101
rect 472 100 473 101
rect 471 100 472 101
rect 470 100 471 101
rect 469 100 470 101
rect 468 100 469 101
rect 467 100 468 101
rect 466 100 467 101
rect 465 100 466 101
rect 464 100 465 101
rect 463 100 464 101
rect 462 100 463 101
rect 461 100 462 101
rect 460 100 461 101
rect 264 100 265 101
rect 263 100 264 101
rect 262 100 263 101
rect 261 100 262 101
rect 260 100 261 101
rect 259 100 260 101
rect 258 100 259 101
rect 257 100 258 101
rect 256 100 257 101
rect 255 100 256 101
rect 254 100 255 101
rect 253 100 254 101
rect 252 100 253 101
rect 251 100 252 101
rect 250 100 251 101
rect 249 100 250 101
rect 248 100 249 101
rect 247 100 248 101
rect 246 100 247 101
rect 245 100 246 101
rect 244 100 245 101
rect 243 100 244 101
rect 242 100 243 101
rect 241 100 242 101
rect 240 100 241 101
rect 239 100 240 101
rect 238 100 239 101
rect 237 100 238 101
rect 236 100 237 101
rect 235 100 236 101
rect 234 100 235 101
rect 233 100 234 101
rect 232 100 233 101
rect 231 100 232 101
rect 230 100 231 101
rect 229 100 230 101
rect 228 100 229 101
rect 227 100 228 101
rect 226 100 227 101
rect 225 100 226 101
rect 224 100 225 101
rect 223 100 224 101
rect 222 100 223 101
rect 221 100 222 101
rect 220 100 221 101
rect 219 100 220 101
rect 218 100 219 101
rect 217 100 218 101
rect 216 100 217 101
rect 215 100 216 101
rect 214 100 215 101
rect 213 100 214 101
rect 212 100 213 101
rect 211 100 212 101
rect 210 100 211 101
rect 209 100 210 101
rect 208 100 209 101
rect 207 100 208 101
rect 206 100 207 101
rect 205 100 206 101
rect 204 100 205 101
rect 203 100 204 101
rect 202 100 203 101
rect 201 100 202 101
rect 200 100 201 101
rect 199 100 200 101
rect 198 100 199 101
rect 197 100 198 101
rect 196 100 197 101
rect 195 100 196 101
rect 194 100 195 101
rect 193 100 194 101
rect 192 100 193 101
rect 191 100 192 101
rect 190 100 191 101
rect 189 100 190 101
rect 188 100 189 101
rect 187 100 188 101
rect 186 100 187 101
rect 185 100 186 101
rect 184 100 185 101
rect 183 100 184 101
rect 182 100 183 101
rect 181 100 182 101
rect 180 100 181 101
rect 179 100 180 101
rect 158 100 159 101
rect 157 100 158 101
rect 156 100 157 101
rect 155 100 156 101
rect 154 100 155 101
rect 153 100 154 101
rect 152 100 153 101
rect 151 100 152 101
rect 150 100 151 101
rect 149 100 150 101
rect 148 100 149 101
rect 147 100 148 101
rect 146 100 147 101
rect 145 100 146 101
rect 144 100 145 101
rect 143 100 144 101
rect 142 100 143 101
rect 141 100 142 101
rect 140 100 141 101
rect 139 100 140 101
rect 138 100 139 101
rect 137 100 138 101
rect 136 100 137 101
rect 135 100 136 101
rect 134 100 135 101
rect 133 100 134 101
rect 132 100 133 101
rect 131 100 132 101
rect 130 100 131 101
rect 129 100 130 101
rect 128 100 129 101
rect 119 100 120 101
rect 118 100 119 101
rect 117 100 118 101
rect 116 100 117 101
rect 115 100 116 101
rect 114 100 115 101
rect 113 100 114 101
rect 112 100 113 101
rect 111 100 112 101
rect 110 100 111 101
rect 109 100 110 101
rect 108 100 109 101
rect 107 100 108 101
rect 106 100 107 101
rect 105 100 106 101
rect 104 100 105 101
rect 103 100 104 101
rect 102 100 103 101
rect 101 100 102 101
rect 100 100 101 101
rect 99 100 100 101
rect 98 100 99 101
rect 97 100 98 101
rect 96 100 97 101
rect 95 100 96 101
rect 94 100 95 101
rect 93 100 94 101
rect 92 100 93 101
rect 91 100 92 101
rect 90 100 91 101
rect 89 100 90 101
rect 88 100 89 101
rect 87 100 88 101
rect 86 100 87 101
rect 85 100 86 101
rect 84 100 85 101
rect 83 100 84 101
rect 82 100 83 101
rect 81 100 82 101
rect 80 100 81 101
rect 79 100 80 101
rect 78 100 79 101
rect 77 100 78 101
rect 76 100 77 101
rect 75 100 76 101
rect 74 100 75 101
rect 69 100 70 101
rect 68 100 69 101
rect 67 100 68 101
rect 66 100 67 101
rect 65 100 66 101
rect 64 100 65 101
rect 63 100 64 101
rect 62 100 63 101
rect 61 100 62 101
rect 60 100 61 101
rect 59 100 60 101
rect 58 100 59 101
rect 57 100 58 101
rect 56 100 57 101
rect 55 100 56 101
rect 54 100 55 101
rect 53 100 54 101
rect 52 100 53 101
rect 51 100 52 101
rect 50 100 51 101
rect 463 101 464 102
rect 462 101 463 102
rect 461 101 462 102
rect 460 101 461 102
rect 265 101 266 102
rect 264 101 265 102
rect 263 101 264 102
rect 262 101 263 102
rect 261 101 262 102
rect 260 101 261 102
rect 259 101 260 102
rect 258 101 259 102
rect 257 101 258 102
rect 256 101 257 102
rect 255 101 256 102
rect 254 101 255 102
rect 253 101 254 102
rect 252 101 253 102
rect 251 101 252 102
rect 250 101 251 102
rect 249 101 250 102
rect 248 101 249 102
rect 247 101 248 102
rect 246 101 247 102
rect 245 101 246 102
rect 244 101 245 102
rect 243 101 244 102
rect 242 101 243 102
rect 241 101 242 102
rect 240 101 241 102
rect 239 101 240 102
rect 238 101 239 102
rect 237 101 238 102
rect 236 101 237 102
rect 235 101 236 102
rect 234 101 235 102
rect 233 101 234 102
rect 232 101 233 102
rect 231 101 232 102
rect 230 101 231 102
rect 229 101 230 102
rect 228 101 229 102
rect 227 101 228 102
rect 226 101 227 102
rect 225 101 226 102
rect 224 101 225 102
rect 223 101 224 102
rect 222 101 223 102
rect 221 101 222 102
rect 220 101 221 102
rect 219 101 220 102
rect 218 101 219 102
rect 217 101 218 102
rect 216 101 217 102
rect 215 101 216 102
rect 214 101 215 102
rect 213 101 214 102
rect 212 101 213 102
rect 211 101 212 102
rect 210 101 211 102
rect 209 101 210 102
rect 208 101 209 102
rect 207 101 208 102
rect 206 101 207 102
rect 205 101 206 102
rect 204 101 205 102
rect 203 101 204 102
rect 202 101 203 102
rect 201 101 202 102
rect 200 101 201 102
rect 199 101 200 102
rect 198 101 199 102
rect 197 101 198 102
rect 196 101 197 102
rect 195 101 196 102
rect 194 101 195 102
rect 193 101 194 102
rect 192 101 193 102
rect 191 101 192 102
rect 190 101 191 102
rect 189 101 190 102
rect 188 101 189 102
rect 187 101 188 102
rect 186 101 187 102
rect 185 101 186 102
rect 184 101 185 102
rect 183 101 184 102
rect 182 101 183 102
rect 181 101 182 102
rect 180 101 181 102
rect 179 101 180 102
rect 158 101 159 102
rect 157 101 158 102
rect 156 101 157 102
rect 155 101 156 102
rect 154 101 155 102
rect 153 101 154 102
rect 152 101 153 102
rect 151 101 152 102
rect 150 101 151 102
rect 149 101 150 102
rect 148 101 149 102
rect 147 101 148 102
rect 146 101 147 102
rect 145 101 146 102
rect 144 101 145 102
rect 143 101 144 102
rect 142 101 143 102
rect 141 101 142 102
rect 140 101 141 102
rect 139 101 140 102
rect 138 101 139 102
rect 137 101 138 102
rect 136 101 137 102
rect 135 101 136 102
rect 134 101 135 102
rect 133 101 134 102
rect 132 101 133 102
rect 131 101 132 102
rect 130 101 131 102
rect 129 101 130 102
rect 128 101 129 102
rect 118 101 119 102
rect 117 101 118 102
rect 116 101 117 102
rect 115 101 116 102
rect 114 101 115 102
rect 113 101 114 102
rect 112 101 113 102
rect 111 101 112 102
rect 110 101 111 102
rect 109 101 110 102
rect 108 101 109 102
rect 107 101 108 102
rect 106 101 107 102
rect 105 101 106 102
rect 104 101 105 102
rect 103 101 104 102
rect 102 101 103 102
rect 101 101 102 102
rect 100 101 101 102
rect 99 101 100 102
rect 98 101 99 102
rect 97 101 98 102
rect 96 101 97 102
rect 95 101 96 102
rect 94 101 95 102
rect 93 101 94 102
rect 92 101 93 102
rect 91 101 92 102
rect 90 101 91 102
rect 89 101 90 102
rect 88 101 89 102
rect 87 101 88 102
rect 86 101 87 102
rect 85 101 86 102
rect 84 101 85 102
rect 83 101 84 102
rect 82 101 83 102
rect 81 101 82 102
rect 80 101 81 102
rect 79 101 80 102
rect 78 101 79 102
rect 77 101 78 102
rect 76 101 77 102
rect 75 101 76 102
rect 74 101 75 102
rect 69 101 70 102
rect 68 101 69 102
rect 67 101 68 102
rect 66 101 67 102
rect 65 101 66 102
rect 64 101 65 102
rect 63 101 64 102
rect 62 101 63 102
rect 61 101 62 102
rect 60 101 61 102
rect 59 101 60 102
rect 58 101 59 102
rect 57 101 58 102
rect 56 101 57 102
rect 55 101 56 102
rect 54 101 55 102
rect 53 101 54 102
rect 52 101 53 102
rect 51 101 52 102
rect 50 101 51 102
rect 49 101 50 102
rect 461 102 462 103
rect 460 102 461 103
rect 397 102 398 103
rect 396 102 397 103
rect 395 102 396 103
rect 267 102 268 103
rect 266 102 267 103
rect 265 102 266 103
rect 264 102 265 103
rect 263 102 264 103
rect 262 102 263 103
rect 261 102 262 103
rect 260 102 261 103
rect 259 102 260 103
rect 258 102 259 103
rect 257 102 258 103
rect 256 102 257 103
rect 255 102 256 103
rect 254 102 255 103
rect 253 102 254 103
rect 252 102 253 103
rect 251 102 252 103
rect 250 102 251 103
rect 249 102 250 103
rect 248 102 249 103
rect 247 102 248 103
rect 246 102 247 103
rect 245 102 246 103
rect 244 102 245 103
rect 243 102 244 103
rect 242 102 243 103
rect 241 102 242 103
rect 240 102 241 103
rect 239 102 240 103
rect 238 102 239 103
rect 237 102 238 103
rect 236 102 237 103
rect 235 102 236 103
rect 234 102 235 103
rect 233 102 234 103
rect 232 102 233 103
rect 231 102 232 103
rect 230 102 231 103
rect 229 102 230 103
rect 228 102 229 103
rect 227 102 228 103
rect 226 102 227 103
rect 225 102 226 103
rect 224 102 225 103
rect 223 102 224 103
rect 222 102 223 103
rect 221 102 222 103
rect 220 102 221 103
rect 219 102 220 103
rect 218 102 219 103
rect 217 102 218 103
rect 216 102 217 103
rect 215 102 216 103
rect 214 102 215 103
rect 213 102 214 103
rect 212 102 213 103
rect 211 102 212 103
rect 210 102 211 103
rect 209 102 210 103
rect 208 102 209 103
rect 207 102 208 103
rect 206 102 207 103
rect 205 102 206 103
rect 204 102 205 103
rect 203 102 204 103
rect 202 102 203 103
rect 201 102 202 103
rect 200 102 201 103
rect 199 102 200 103
rect 198 102 199 103
rect 197 102 198 103
rect 196 102 197 103
rect 195 102 196 103
rect 194 102 195 103
rect 193 102 194 103
rect 192 102 193 103
rect 191 102 192 103
rect 190 102 191 103
rect 189 102 190 103
rect 188 102 189 103
rect 187 102 188 103
rect 186 102 187 103
rect 185 102 186 103
rect 184 102 185 103
rect 183 102 184 103
rect 182 102 183 103
rect 181 102 182 103
rect 180 102 181 103
rect 179 102 180 103
rect 178 102 179 103
rect 157 102 158 103
rect 156 102 157 103
rect 155 102 156 103
rect 154 102 155 103
rect 153 102 154 103
rect 152 102 153 103
rect 151 102 152 103
rect 150 102 151 103
rect 149 102 150 103
rect 148 102 149 103
rect 147 102 148 103
rect 146 102 147 103
rect 145 102 146 103
rect 144 102 145 103
rect 143 102 144 103
rect 142 102 143 103
rect 141 102 142 103
rect 140 102 141 103
rect 139 102 140 103
rect 138 102 139 103
rect 137 102 138 103
rect 136 102 137 103
rect 135 102 136 103
rect 134 102 135 103
rect 133 102 134 103
rect 132 102 133 103
rect 131 102 132 103
rect 130 102 131 103
rect 129 102 130 103
rect 128 102 129 103
rect 117 102 118 103
rect 116 102 117 103
rect 115 102 116 103
rect 114 102 115 103
rect 113 102 114 103
rect 112 102 113 103
rect 111 102 112 103
rect 110 102 111 103
rect 109 102 110 103
rect 108 102 109 103
rect 107 102 108 103
rect 106 102 107 103
rect 105 102 106 103
rect 104 102 105 103
rect 103 102 104 103
rect 102 102 103 103
rect 101 102 102 103
rect 100 102 101 103
rect 99 102 100 103
rect 98 102 99 103
rect 97 102 98 103
rect 96 102 97 103
rect 95 102 96 103
rect 94 102 95 103
rect 93 102 94 103
rect 92 102 93 103
rect 91 102 92 103
rect 90 102 91 103
rect 89 102 90 103
rect 88 102 89 103
rect 87 102 88 103
rect 86 102 87 103
rect 85 102 86 103
rect 84 102 85 103
rect 83 102 84 103
rect 82 102 83 103
rect 81 102 82 103
rect 80 102 81 103
rect 79 102 80 103
rect 78 102 79 103
rect 77 102 78 103
rect 76 102 77 103
rect 75 102 76 103
rect 74 102 75 103
rect 68 102 69 103
rect 67 102 68 103
rect 66 102 67 103
rect 65 102 66 103
rect 64 102 65 103
rect 63 102 64 103
rect 62 102 63 103
rect 61 102 62 103
rect 60 102 61 103
rect 59 102 60 103
rect 58 102 59 103
rect 57 102 58 103
rect 56 102 57 103
rect 55 102 56 103
rect 54 102 55 103
rect 53 102 54 103
rect 52 102 53 103
rect 51 102 52 103
rect 50 102 51 103
rect 49 102 50 103
rect 48 102 49 103
rect 460 103 461 104
rect 397 103 398 104
rect 396 103 397 104
rect 395 103 396 104
rect 268 103 269 104
rect 267 103 268 104
rect 266 103 267 104
rect 265 103 266 104
rect 264 103 265 104
rect 263 103 264 104
rect 262 103 263 104
rect 261 103 262 104
rect 260 103 261 104
rect 259 103 260 104
rect 258 103 259 104
rect 257 103 258 104
rect 256 103 257 104
rect 255 103 256 104
rect 254 103 255 104
rect 253 103 254 104
rect 252 103 253 104
rect 251 103 252 104
rect 250 103 251 104
rect 249 103 250 104
rect 248 103 249 104
rect 247 103 248 104
rect 246 103 247 104
rect 245 103 246 104
rect 244 103 245 104
rect 243 103 244 104
rect 242 103 243 104
rect 241 103 242 104
rect 240 103 241 104
rect 239 103 240 104
rect 238 103 239 104
rect 237 103 238 104
rect 236 103 237 104
rect 235 103 236 104
rect 234 103 235 104
rect 233 103 234 104
rect 232 103 233 104
rect 231 103 232 104
rect 230 103 231 104
rect 229 103 230 104
rect 228 103 229 104
rect 227 103 228 104
rect 226 103 227 104
rect 225 103 226 104
rect 224 103 225 104
rect 223 103 224 104
rect 222 103 223 104
rect 221 103 222 104
rect 220 103 221 104
rect 219 103 220 104
rect 218 103 219 104
rect 217 103 218 104
rect 216 103 217 104
rect 215 103 216 104
rect 214 103 215 104
rect 213 103 214 104
rect 212 103 213 104
rect 211 103 212 104
rect 210 103 211 104
rect 209 103 210 104
rect 208 103 209 104
rect 207 103 208 104
rect 206 103 207 104
rect 205 103 206 104
rect 204 103 205 104
rect 203 103 204 104
rect 202 103 203 104
rect 201 103 202 104
rect 200 103 201 104
rect 199 103 200 104
rect 198 103 199 104
rect 197 103 198 104
rect 196 103 197 104
rect 195 103 196 104
rect 194 103 195 104
rect 193 103 194 104
rect 192 103 193 104
rect 191 103 192 104
rect 190 103 191 104
rect 189 103 190 104
rect 188 103 189 104
rect 187 103 188 104
rect 186 103 187 104
rect 185 103 186 104
rect 184 103 185 104
rect 183 103 184 104
rect 182 103 183 104
rect 181 103 182 104
rect 180 103 181 104
rect 179 103 180 104
rect 178 103 179 104
rect 177 103 178 104
rect 157 103 158 104
rect 156 103 157 104
rect 155 103 156 104
rect 154 103 155 104
rect 153 103 154 104
rect 152 103 153 104
rect 151 103 152 104
rect 150 103 151 104
rect 149 103 150 104
rect 148 103 149 104
rect 147 103 148 104
rect 146 103 147 104
rect 145 103 146 104
rect 144 103 145 104
rect 143 103 144 104
rect 142 103 143 104
rect 141 103 142 104
rect 140 103 141 104
rect 139 103 140 104
rect 138 103 139 104
rect 137 103 138 104
rect 136 103 137 104
rect 135 103 136 104
rect 134 103 135 104
rect 133 103 134 104
rect 132 103 133 104
rect 131 103 132 104
rect 130 103 131 104
rect 129 103 130 104
rect 128 103 129 104
rect 127 103 128 104
rect 116 103 117 104
rect 115 103 116 104
rect 114 103 115 104
rect 113 103 114 104
rect 112 103 113 104
rect 111 103 112 104
rect 110 103 111 104
rect 109 103 110 104
rect 108 103 109 104
rect 107 103 108 104
rect 106 103 107 104
rect 105 103 106 104
rect 104 103 105 104
rect 103 103 104 104
rect 102 103 103 104
rect 101 103 102 104
rect 100 103 101 104
rect 99 103 100 104
rect 98 103 99 104
rect 97 103 98 104
rect 96 103 97 104
rect 95 103 96 104
rect 94 103 95 104
rect 93 103 94 104
rect 92 103 93 104
rect 91 103 92 104
rect 90 103 91 104
rect 89 103 90 104
rect 88 103 89 104
rect 87 103 88 104
rect 86 103 87 104
rect 85 103 86 104
rect 84 103 85 104
rect 83 103 84 104
rect 82 103 83 104
rect 81 103 82 104
rect 80 103 81 104
rect 79 103 80 104
rect 78 103 79 104
rect 77 103 78 104
rect 76 103 77 104
rect 75 103 76 104
rect 74 103 75 104
rect 68 103 69 104
rect 67 103 68 104
rect 66 103 67 104
rect 65 103 66 104
rect 64 103 65 104
rect 63 103 64 104
rect 62 103 63 104
rect 61 103 62 104
rect 60 103 61 104
rect 59 103 60 104
rect 58 103 59 104
rect 57 103 58 104
rect 56 103 57 104
rect 55 103 56 104
rect 54 103 55 104
rect 53 103 54 104
rect 52 103 53 104
rect 51 103 52 104
rect 50 103 51 104
rect 49 103 50 104
rect 48 103 49 104
rect 47 103 48 104
rect 397 104 398 105
rect 396 104 397 105
rect 395 104 396 105
rect 269 104 270 105
rect 268 104 269 105
rect 267 104 268 105
rect 266 104 267 105
rect 265 104 266 105
rect 264 104 265 105
rect 263 104 264 105
rect 262 104 263 105
rect 261 104 262 105
rect 260 104 261 105
rect 259 104 260 105
rect 258 104 259 105
rect 257 104 258 105
rect 256 104 257 105
rect 255 104 256 105
rect 254 104 255 105
rect 253 104 254 105
rect 252 104 253 105
rect 251 104 252 105
rect 250 104 251 105
rect 249 104 250 105
rect 248 104 249 105
rect 247 104 248 105
rect 246 104 247 105
rect 245 104 246 105
rect 244 104 245 105
rect 243 104 244 105
rect 242 104 243 105
rect 241 104 242 105
rect 240 104 241 105
rect 239 104 240 105
rect 238 104 239 105
rect 237 104 238 105
rect 236 104 237 105
rect 235 104 236 105
rect 234 104 235 105
rect 233 104 234 105
rect 232 104 233 105
rect 231 104 232 105
rect 230 104 231 105
rect 229 104 230 105
rect 228 104 229 105
rect 227 104 228 105
rect 226 104 227 105
rect 225 104 226 105
rect 224 104 225 105
rect 223 104 224 105
rect 222 104 223 105
rect 221 104 222 105
rect 220 104 221 105
rect 219 104 220 105
rect 218 104 219 105
rect 217 104 218 105
rect 216 104 217 105
rect 215 104 216 105
rect 214 104 215 105
rect 213 104 214 105
rect 212 104 213 105
rect 211 104 212 105
rect 210 104 211 105
rect 209 104 210 105
rect 208 104 209 105
rect 207 104 208 105
rect 206 104 207 105
rect 205 104 206 105
rect 204 104 205 105
rect 203 104 204 105
rect 202 104 203 105
rect 201 104 202 105
rect 200 104 201 105
rect 199 104 200 105
rect 198 104 199 105
rect 197 104 198 105
rect 196 104 197 105
rect 195 104 196 105
rect 194 104 195 105
rect 193 104 194 105
rect 192 104 193 105
rect 191 104 192 105
rect 190 104 191 105
rect 189 104 190 105
rect 188 104 189 105
rect 187 104 188 105
rect 186 104 187 105
rect 185 104 186 105
rect 184 104 185 105
rect 183 104 184 105
rect 182 104 183 105
rect 181 104 182 105
rect 180 104 181 105
rect 179 104 180 105
rect 178 104 179 105
rect 177 104 178 105
rect 157 104 158 105
rect 156 104 157 105
rect 155 104 156 105
rect 154 104 155 105
rect 153 104 154 105
rect 152 104 153 105
rect 151 104 152 105
rect 150 104 151 105
rect 149 104 150 105
rect 148 104 149 105
rect 147 104 148 105
rect 146 104 147 105
rect 145 104 146 105
rect 144 104 145 105
rect 143 104 144 105
rect 142 104 143 105
rect 141 104 142 105
rect 140 104 141 105
rect 139 104 140 105
rect 138 104 139 105
rect 137 104 138 105
rect 136 104 137 105
rect 135 104 136 105
rect 134 104 135 105
rect 133 104 134 105
rect 132 104 133 105
rect 131 104 132 105
rect 130 104 131 105
rect 129 104 130 105
rect 128 104 129 105
rect 127 104 128 105
rect 116 104 117 105
rect 115 104 116 105
rect 114 104 115 105
rect 113 104 114 105
rect 112 104 113 105
rect 111 104 112 105
rect 110 104 111 105
rect 109 104 110 105
rect 108 104 109 105
rect 107 104 108 105
rect 106 104 107 105
rect 105 104 106 105
rect 104 104 105 105
rect 103 104 104 105
rect 102 104 103 105
rect 101 104 102 105
rect 100 104 101 105
rect 99 104 100 105
rect 98 104 99 105
rect 97 104 98 105
rect 96 104 97 105
rect 95 104 96 105
rect 94 104 95 105
rect 93 104 94 105
rect 92 104 93 105
rect 91 104 92 105
rect 90 104 91 105
rect 89 104 90 105
rect 88 104 89 105
rect 87 104 88 105
rect 86 104 87 105
rect 85 104 86 105
rect 84 104 85 105
rect 83 104 84 105
rect 82 104 83 105
rect 81 104 82 105
rect 80 104 81 105
rect 79 104 80 105
rect 78 104 79 105
rect 77 104 78 105
rect 76 104 77 105
rect 75 104 76 105
rect 74 104 75 105
rect 73 104 74 105
rect 67 104 68 105
rect 66 104 67 105
rect 65 104 66 105
rect 64 104 65 105
rect 63 104 64 105
rect 62 104 63 105
rect 61 104 62 105
rect 60 104 61 105
rect 59 104 60 105
rect 58 104 59 105
rect 57 104 58 105
rect 56 104 57 105
rect 55 104 56 105
rect 54 104 55 105
rect 53 104 54 105
rect 52 104 53 105
rect 51 104 52 105
rect 50 104 51 105
rect 49 104 50 105
rect 48 104 49 105
rect 47 104 48 105
rect 46 104 47 105
rect 397 105 398 106
rect 396 105 397 106
rect 395 105 396 106
rect 270 105 271 106
rect 269 105 270 106
rect 268 105 269 106
rect 267 105 268 106
rect 266 105 267 106
rect 265 105 266 106
rect 264 105 265 106
rect 263 105 264 106
rect 262 105 263 106
rect 261 105 262 106
rect 260 105 261 106
rect 259 105 260 106
rect 258 105 259 106
rect 257 105 258 106
rect 256 105 257 106
rect 255 105 256 106
rect 254 105 255 106
rect 253 105 254 106
rect 252 105 253 106
rect 251 105 252 106
rect 250 105 251 106
rect 249 105 250 106
rect 248 105 249 106
rect 247 105 248 106
rect 246 105 247 106
rect 245 105 246 106
rect 244 105 245 106
rect 243 105 244 106
rect 242 105 243 106
rect 241 105 242 106
rect 240 105 241 106
rect 239 105 240 106
rect 238 105 239 106
rect 237 105 238 106
rect 236 105 237 106
rect 235 105 236 106
rect 234 105 235 106
rect 233 105 234 106
rect 232 105 233 106
rect 231 105 232 106
rect 230 105 231 106
rect 229 105 230 106
rect 228 105 229 106
rect 227 105 228 106
rect 226 105 227 106
rect 225 105 226 106
rect 224 105 225 106
rect 223 105 224 106
rect 222 105 223 106
rect 221 105 222 106
rect 220 105 221 106
rect 219 105 220 106
rect 218 105 219 106
rect 217 105 218 106
rect 216 105 217 106
rect 215 105 216 106
rect 214 105 215 106
rect 213 105 214 106
rect 212 105 213 106
rect 211 105 212 106
rect 210 105 211 106
rect 209 105 210 106
rect 208 105 209 106
rect 207 105 208 106
rect 206 105 207 106
rect 205 105 206 106
rect 204 105 205 106
rect 203 105 204 106
rect 202 105 203 106
rect 201 105 202 106
rect 200 105 201 106
rect 199 105 200 106
rect 198 105 199 106
rect 197 105 198 106
rect 196 105 197 106
rect 195 105 196 106
rect 194 105 195 106
rect 193 105 194 106
rect 192 105 193 106
rect 191 105 192 106
rect 190 105 191 106
rect 189 105 190 106
rect 188 105 189 106
rect 187 105 188 106
rect 186 105 187 106
rect 185 105 186 106
rect 184 105 185 106
rect 183 105 184 106
rect 182 105 183 106
rect 181 105 182 106
rect 180 105 181 106
rect 179 105 180 106
rect 178 105 179 106
rect 177 105 178 106
rect 176 105 177 106
rect 156 105 157 106
rect 155 105 156 106
rect 154 105 155 106
rect 153 105 154 106
rect 152 105 153 106
rect 151 105 152 106
rect 150 105 151 106
rect 149 105 150 106
rect 148 105 149 106
rect 147 105 148 106
rect 146 105 147 106
rect 145 105 146 106
rect 144 105 145 106
rect 143 105 144 106
rect 142 105 143 106
rect 141 105 142 106
rect 140 105 141 106
rect 139 105 140 106
rect 138 105 139 106
rect 137 105 138 106
rect 136 105 137 106
rect 135 105 136 106
rect 134 105 135 106
rect 133 105 134 106
rect 132 105 133 106
rect 131 105 132 106
rect 130 105 131 106
rect 129 105 130 106
rect 128 105 129 106
rect 127 105 128 106
rect 115 105 116 106
rect 114 105 115 106
rect 113 105 114 106
rect 112 105 113 106
rect 111 105 112 106
rect 110 105 111 106
rect 109 105 110 106
rect 108 105 109 106
rect 107 105 108 106
rect 106 105 107 106
rect 105 105 106 106
rect 104 105 105 106
rect 103 105 104 106
rect 102 105 103 106
rect 101 105 102 106
rect 100 105 101 106
rect 99 105 100 106
rect 98 105 99 106
rect 97 105 98 106
rect 96 105 97 106
rect 95 105 96 106
rect 94 105 95 106
rect 93 105 94 106
rect 92 105 93 106
rect 91 105 92 106
rect 90 105 91 106
rect 89 105 90 106
rect 88 105 89 106
rect 87 105 88 106
rect 86 105 87 106
rect 85 105 86 106
rect 84 105 85 106
rect 83 105 84 106
rect 82 105 83 106
rect 81 105 82 106
rect 80 105 81 106
rect 79 105 80 106
rect 78 105 79 106
rect 77 105 78 106
rect 76 105 77 106
rect 75 105 76 106
rect 74 105 75 106
rect 73 105 74 106
rect 67 105 68 106
rect 66 105 67 106
rect 65 105 66 106
rect 64 105 65 106
rect 63 105 64 106
rect 62 105 63 106
rect 61 105 62 106
rect 60 105 61 106
rect 59 105 60 106
rect 58 105 59 106
rect 57 105 58 106
rect 56 105 57 106
rect 55 105 56 106
rect 54 105 55 106
rect 53 105 54 106
rect 52 105 53 106
rect 51 105 52 106
rect 50 105 51 106
rect 49 105 50 106
rect 48 105 49 106
rect 47 105 48 106
rect 46 105 47 106
rect 45 105 46 106
rect 44 105 45 106
rect 398 106 399 107
rect 397 106 398 107
rect 396 106 397 107
rect 395 106 396 107
rect 271 106 272 107
rect 270 106 271 107
rect 269 106 270 107
rect 268 106 269 107
rect 267 106 268 107
rect 266 106 267 107
rect 265 106 266 107
rect 264 106 265 107
rect 263 106 264 107
rect 262 106 263 107
rect 261 106 262 107
rect 260 106 261 107
rect 259 106 260 107
rect 258 106 259 107
rect 257 106 258 107
rect 256 106 257 107
rect 255 106 256 107
rect 254 106 255 107
rect 253 106 254 107
rect 252 106 253 107
rect 251 106 252 107
rect 250 106 251 107
rect 249 106 250 107
rect 248 106 249 107
rect 247 106 248 107
rect 246 106 247 107
rect 245 106 246 107
rect 244 106 245 107
rect 243 106 244 107
rect 242 106 243 107
rect 241 106 242 107
rect 240 106 241 107
rect 239 106 240 107
rect 238 106 239 107
rect 237 106 238 107
rect 236 106 237 107
rect 235 106 236 107
rect 234 106 235 107
rect 233 106 234 107
rect 232 106 233 107
rect 231 106 232 107
rect 230 106 231 107
rect 229 106 230 107
rect 228 106 229 107
rect 227 106 228 107
rect 226 106 227 107
rect 225 106 226 107
rect 224 106 225 107
rect 223 106 224 107
rect 222 106 223 107
rect 221 106 222 107
rect 220 106 221 107
rect 219 106 220 107
rect 218 106 219 107
rect 217 106 218 107
rect 216 106 217 107
rect 215 106 216 107
rect 214 106 215 107
rect 213 106 214 107
rect 212 106 213 107
rect 211 106 212 107
rect 210 106 211 107
rect 209 106 210 107
rect 208 106 209 107
rect 207 106 208 107
rect 206 106 207 107
rect 205 106 206 107
rect 204 106 205 107
rect 203 106 204 107
rect 202 106 203 107
rect 201 106 202 107
rect 200 106 201 107
rect 199 106 200 107
rect 198 106 199 107
rect 197 106 198 107
rect 196 106 197 107
rect 195 106 196 107
rect 194 106 195 107
rect 193 106 194 107
rect 192 106 193 107
rect 191 106 192 107
rect 190 106 191 107
rect 189 106 190 107
rect 188 106 189 107
rect 187 106 188 107
rect 186 106 187 107
rect 185 106 186 107
rect 184 106 185 107
rect 183 106 184 107
rect 182 106 183 107
rect 181 106 182 107
rect 180 106 181 107
rect 179 106 180 107
rect 178 106 179 107
rect 177 106 178 107
rect 176 106 177 107
rect 175 106 176 107
rect 156 106 157 107
rect 155 106 156 107
rect 154 106 155 107
rect 153 106 154 107
rect 152 106 153 107
rect 151 106 152 107
rect 150 106 151 107
rect 149 106 150 107
rect 148 106 149 107
rect 147 106 148 107
rect 146 106 147 107
rect 145 106 146 107
rect 144 106 145 107
rect 143 106 144 107
rect 142 106 143 107
rect 141 106 142 107
rect 140 106 141 107
rect 139 106 140 107
rect 138 106 139 107
rect 137 106 138 107
rect 136 106 137 107
rect 135 106 136 107
rect 134 106 135 107
rect 133 106 134 107
rect 132 106 133 107
rect 131 106 132 107
rect 130 106 131 107
rect 129 106 130 107
rect 128 106 129 107
rect 127 106 128 107
rect 126 106 127 107
rect 115 106 116 107
rect 114 106 115 107
rect 113 106 114 107
rect 112 106 113 107
rect 111 106 112 107
rect 110 106 111 107
rect 109 106 110 107
rect 108 106 109 107
rect 107 106 108 107
rect 106 106 107 107
rect 105 106 106 107
rect 104 106 105 107
rect 103 106 104 107
rect 102 106 103 107
rect 101 106 102 107
rect 100 106 101 107
rect 99 106 100 107
rect 98 106 99 107
rect 97 106 98 107
rect 96 106 97 107
rect 95 106 96 107
rect 94 106 95 107
rect 93 106 94 107
rect 92 106 93 107
rect 91 106 92 107
rect 90 106 91 107
rect 89 106 90 107
rect 88 106 89 107
rect 87 106 88 107
rect 86 106 87 107
rect 85 106 86 107
rect 84 106 85 107
rect 83 106 84 107
rect 82 106 83 107
rect 81 106 82 107
rect 80 106 81 107
rect 79 106 80 107
rect 78 106 79 107
rect 77 106 78 107
rect 66 106 67 107
rect 65 106 66 107
rect 64 106 65 107
rect 63 106 64 107
rect 62 106 63 107
rect 61 106 62 107
rect 60 106 61 107
rect 59 106 60 107
rect 58 106 59 107
rect 57 106 58 107
rect 56 106 57 107
rect 55 106 56 107
rect 54 106 55 107
rect 53 106 54 107
rect 52 106 53 107
rect 51 106 52 107
rect 50 106 51 107
rect 49 106 50 107
rect 48 106 49 107
rect 47 106 48 107
rect 46 106 47 107
rect 45 106 46 107
rect 44 106 45 107
rect 43 106 44 107
rect 423 107 424 108
rect 422 107 423 108
rect 421 107 422 108
rect 420 107 421 108
rect 419 107 420 108
rect 418 107 419 108
rect 417 107 418 108
rect 416 107 417 108
rect 415 107 416 108
rect 414 107 415 108
rect 413 107 414 108
rect 412 107 413 108
rect 411 107 412 108
rect 410 107 411 108
rect 409 107 410 108
rect 408 107 409 108
rect 407 107 408 108
rect 406 107 407 108
rect 405 107 406 108
rect 404 107 405 108
rect 403 107 404 108
rect 402 107 403 108
rect 401 107 402 108
rect 400 107 401 108
rect 399 107 400 108
rect 398 107 399 108
rect 397 107 398 108
rect 396 107 397 108
rect 395 107 396 108
rect 272 107 273 108
rect 271 107 272 108
rect 270 107 271 108
rect 269 107 270 108
rect 268 107 269 108
rect 267 107 268 108
rect 266 107 267 108
rect 265 107 266 108
rect 264 107 265 108
rect 263 107 264 108
rect 262 107 263 108
rect 261 107 262 108
rect 260 107 261 108
rect 259 107 260 108
rect 258 107 259 108
rect 257 107 258 108
rect 256 107 257 108
rect 255 107 256 108
rect 254 107 255 108
rect 253 107 254 108
rect 252 107 253 108
rect 251 107 252 108
rect 250 107 251 108
rect 249 107 250 108
rect 248 107 249 108
rect 247 107 248 108
rect 246 107 247 108
rect 245 107 246 108
rect 244 107 245 108
rect 243 107 244 108
rect 242 107 243 108
rect 241 107 242 108
rect 240 107 241 108
rect 239 107 240 108
rect 238 107 239 108
rect 237 107 238 108
rect 236 107 237 108
rect 235 107 236 108
rect 234 107 235 108
rect 233 107 234 108
rect 232 107 233 108
rect 231 107 232 108
rect 230 107 231 108
rect 229 107 230 108
rect 228 107 229 108
rect 227 107 228 108
rect 226 107 227 108
rect 225 107 226 108
rect 224 107 225 108
rect 223 107 224 108
rect 222 107 223 108
rect 221 107 222 108
rect 220 107 221 108
rect 219 107 220 108
rect 218 107 219 108
rect 217 107 218 108
rect 216 107 217 108
rect 215 107 216 108
rect 214 107 215 108
rect 213 107 214 108
rect 212 107 213 108
rect 211 107 212 108
rect 210 107 211 108
rect 209 107 210 108
rect 208 107 209 108
rect 207 107 208 108
rect 206 107 207 108
rect 205 107 206 108
rect 204 107 205 108
rect 203 107 204 108
rect 202 107 203 108
rect 201 107 202 108
rect 200 107 201 108
rect 199 107 200 108
rect 198 107 199 108
rect 197 107 198 108
rect 196 107 197 108
rect 195 107 196 108
rect 194 107 195 108
rect 193 107 194 108
rect 192 107 193 108
rect 191 107 192 108
rect 190 107 191 108
rect 189 107 190 108
rect 188 107 189 108
rect 187 107 188 108
rect 186 107 187 108
rect 185 107 186 108
rect 184 107 185 108
rect 183 107 184 108
rect 182 107 183 108
rect 181 107 182 108
rect 180 107 181 108
rect 179 107 180 108
rect 178 107 179 108
rect 177 107 178 108
rect 176 107 177 108
rect 175 107 176 108
rect 156 107 157 108
rect 155 107 156 108
rect 154 107 155 108
rect 153 107 154 108
rect 152 107 153 108
rect 151 107 152 108
rect 150 107 151 108
rect 149 107 150 108
rect 148 107 149 108
rect 147 107 148 108
rect 146 107 147 108
rect 145 107 146 108
rect 144 107 145 108
rect 143 107 144 108
rect 142 107 143 108
rect 141 107 142 108
rect 140 107 141 108
rect 139 107 140 108
rect 138 107 139 108
rect 137 107 138 108
rect 136 107 137 108
rect 135 107 136 108
rect 134 107 135 108
rect 133 107 134 108
rect 132 107 133 108
rect 131 107 132 108
rect 130 107 131 108
rect 129 107 130 108
rect 128 107 129 108
rect 127 107 128 108
rect 126 107 127 108
rect 116 107 117 108
rect 115 107 116 108
rect 114 107 115 108
rect 113 107 114 108
rect 112 107 113 108
rect 111 107 112 108
rect 110 107 111 108
rect 109 107 110 108
rect 108 107 109 108
rect 107 107 108 108
rect 106 107 107 108
rect 105 107 106 108
rect 104 107 105 108
rect 103 107 104 108
rect 102 107 103 108
rect 101 107 102 108
rect 100 107 101 108
rect 99 107 100 108
rect 98 107 99 108
rect 97 107 98 108
rect 96 107 97 108
rect 95 107 96 108
rect 94 107 95 108
rect 93 107 94 108
rect 92 107 93 108
rect 91 107 92 108
rect 90 107 91 108
rect 89 107 90 108
rect 88 107 89 108
rect 87 107 88 108
rect 86 107 87 108
rect 85 107 86 108
rect 84 107 85 108
rect 83 107 84 108
rect 82 107 83 108
rect 81 107 82 108
rect 80 107 81 108
rect 65 107 66 108
rect 64 107 65 108
rect 63 107 64 108
rect 62 107 63 108
rect 61 107 62 108
rect 60 107 61 108
rect 59 107 60 108
rect 58 107 59 108
rect 57 107 58 108
rect 56 107 57 108
rect 55 107 56 108
rect 54 107 55 108
rect 53 107 54 108
rect 52 107 53 108
rect 51 107 52 108
rect 50 107 51 108
rect 49 107 50 108
rect 48 107 49 108
rect 47 107 48 108
rect 46 107 47 108
rect 45 107 46 108
rect 44 107 45 108
rect 43 107 44 108
rect 42 107 43 108
rect 41 107 42 108
rect 429 108 430 109
rect 428 108 429 109
rect 427 108 428 109
rect 426 108 427 109
rect 425 108 426 109
rect 424 108 425 109
rect 423 108 424 109
rect 422 108 423 109
rect 421 108 422 109
rect 420 108 421 109
rect 419 108 420 109
rect 418 108 419 109
rect 417 108 418 109
rect 416 108 417 109
rect 415 108 416 109
rect 414 108 415 109
rect 413 108 414 109
rect 412 108 413 109
rect 411 108 412 109
rect 410 108 411 109
rect 409 108 410 109
rect 408 108 409 109
rect 407 108 408 109
rect 406 108 407 109
rect 405 108 406 109
rect 404 108 405 109
rect 403 108 404 109
rect 402 108 403 109
rect 401 108 402 109
rect 400 108 401 109
rect 399 108 400 109
rect 398 108 399 109
rect 397 108 398 109
rect 396 108 397 109
rect 395 108 396 109
rect 273 108 274 109
rect 272 108 273 109
rect 271 108 272 109
rect 270 108 271 109
rect 269 108 270 109
rect 268 108 269 109
rect 267 108 268 109
rect 266 108 267 109
rect 265 108 266 109
rect 264 108 265 109
rect 263 108 264 109
rect 262 108 263 109
rect 261 108 262 109
rect 260 108 261 109
rect 259 108 260 109
rect 258 108 259 109
rect 257 108 258 109
rect 256 108 257 109
rect 255 108 256 109
rect 254 108 255 109
rect 253 108 254 109
rect 252 108 253 109
rect 251 108 252 109
rect 250 108 251 109
rect 249 108 250 109
rect 248 108 249 109
rect 247 108 248 109
rect 246 108 247 109
rect 245 108 246 109
rect 244 108 245 109
rect 243 108 244 109
rect 242 108 243 109
rect 241 108 242 109
rect 240 108 241 109
rect 239 108 240 109
rect 238 108 239 109
rect 237 108 238 109
rect 236 108 237 109
rect 235 108 236 109
rect 234 108 235 109
rect 233 108 234 109
rect 232 108 233 109
rect 231 108 232 109
rect 230 108 231 109
rect 229 108 230 109
rect 228 108 229 109
rect 227 108 228 109
rect 226 108 227 109
rect 225 108 226 109
rect 224 108 225 109
rect 223 108 224 109
rect 222 108 223 109
rect 221 108 222 109
rect 220 108 221 109
rect 219 108 220 109
rect 218 108 219 109
rect 217 108 218 109
rect 216 108 217 109
rect 215 108 216 109
rect 214 108 215 109
rect 213 108 214 109
rect 212 108 213 109
rect 211 108 212 109
rect 210 108 211 109
rect 209 108 210 109
rect 208 108 209 109
rect 207 108 208 109
rect 206 108 207 109
rect 205 108 206 109
rect 204 108 205 109
rect 203 108 204 109
rect 202 108 203 109
rect 201 108 202 109
rect 200 108 201 109
rect 199 108 200 109
rect 198 108 199 109
rect 197 108 198 109
rect 196 108 197 109
rect 195 108 196 109
rect 194 108 195 109
rect 193 108 194 109
rect 192 108 193 109
rect 191 108 192 109
rect 190 108 191 109
rect 189 108 190 109
rect 188 108 189 109
rect 187 108 188 109
rect 186 108 187 109
rect 185 108 186 109
rect 184 108 185 109
rect 183 108 184 109
rect 182 108 183 109
rect 181 108 182 109
rect 180 108 181 109
rect 179 108 180 109
rect 178 108 179 109
rect 177 108 178 109
rect 176 108 177 109
rect 175 108 176 109
rect 174 108 175 109
rect 155 108 156 109
rect 154 108 155 109
rect 153 108 154 109
rect 152 108 153 109
rect 151 108 152 109
rect 150 108 151 109
rect 149 108 150 109
rect 148 108 149 109
rect 147 108 148 109
rect 146 108 147 109
rect 145 108 146 109
rect 144 108 145 109
rect 143 108 144 109
rect 142 108 143 109
rect 141 108 142 109
rect 140 108 141 109
rect 139 108 140 109
rect 138 108 139 109
rect 137 108 138 109
rect 136 108 137 109
rect 135 108 136 109
rect 134 108 135 109
rect 133 108 134 109
rect 132 108 133 109
rect 131 108 132 109
rect 130 108 131 109
rect 129 108 130 109
rect 128 108 129 109
rect 127 108 128 109
rect 126 108 127 109
rect 116 108 117 109
rect 115 108 116 109
rect 114 108 115 109
rect 113 108 114 109
rect 112 108 113 109
rect 111 108 112 109
rect 110 108 111 109
rect 109 108 110 109
rect 108 108 109 109
rect 107 108 108 109
rect 106 108 107 109
rect 105 108 106 109
rect 104 108 105 109
rect 103 108 104 109
rect 102 108 103 109
rect 101 108 102 109
rect 100 108 101 109
rect 99 108 100 109
rect 98 108 99 109
rect 97 108 98 109
rect 96 108 97 109
rect 95 108 96 109
rect 94 108 95 109
rect 93 108 94 109
rect 92 108 93 109
rect 91 108 92 109
rect 90 108 91 109
rect 89 108 90 109
rect 88 108 89 109
rect 87 108 88 109
rect 86 108 87 109
rect 85 108 86 109
rect 84 108 85 109
rect 83 108 84 109
rect 82 108 83 109
rect 81 108 82 109
rect 65 108 66 109
rect 64 108 65 109
rect 63 108 64 109
rect 62 108 63 109
rect 61 108 62 109
rect 60 108 61 109
rect 59 108 60 109
rect 58 108 59 109
rect 57 108 58 109
rect 56 108 57 109
rect 55 108 56 109
rect 54 108 55 109
rect 53 108 54 109
rect 52 108 53 109
rect 51 108 52 109
rect 50 108 51 109
rect 49 108 50 109
rect 48 108 49 109
rect 47 108 48 109
rect 46 108 47 109
rect 45 108 46 109
rect 44 108 45 109
rect 43 108 44 109
rect 42 108 43 109
rect 41 108 42 109
rect 40 108 41 109
rect 432 109 433 110
rect 431 109 432 110
rect 430 109 431 110
rect 429 109 430 110
rect 428 109 429 110
rect 427 109 428 110
rect 426 109 427 110
rect 425 109 426 110
rect 424 109 425 110
rect 423 109 424 110
rect 422 109 423 110
rect 421 109 422 110
rect 420 109 421 110
rect 419 109 420 110
rect 418 109 419 110
rect 417 109 418 110
rect 416 109 417 110
rect 415 109 416 110
rect 414 109 415 110
rect 413 109 414 110
rect 412 109 413 110
rect 411 109 412 110
rect 410 109 411 110
rect 409 109 410 110
rect 408 109 409 110
rect 407 109 408 110
rect 406 109 407 110
rect 405 109 406 110
rect 404 109 405 110
rect 403 109 404 110
rect 402 109 403 110
rect 401 109 402 110
rect 400 109 401 110
rect 399 109 400 110
rect 398 109 399 110
rect 397 109 398 110
rect 396 109 397 110
rect 395 109 396 110
rect 274 109 275 110
rect 273 109 274 110
rect 272 109 273 110
rect 271 109 272 110
rect 270 109 271 110
rect 269 109 270 110
rect 268 109 269 110
rect 267 109 268 110
rect 266 109 267 110
rect 265 109 266 110
rect 264 109 265 110
rect 263 109 264 110
rect 262 109 263 110
rect 261 109 262 110
rect 260 109 261 110
rect 259 109 260 110
rect 258 109 259 110
rect 257 109 258 110
rect 256 109 257 110
rect 255 109 256 110
rect 254 109 255 110
rect 253 109 254 110
rect 252 109 253 110
rect 251 109 252 110
rect 250 109 251 110
rect 249 109 250 110
rect 248 109 249 110
rect 247 109 248 110
rect 246 109 247 110
rect 245 109 246 110
rect 244 109 245 110
rect 243 109 244 110
rect 242 109 243 110
rect 241 109 242 110
rect 240 109 241 110
rect 239 109 240 110
rect 238 109 239 110
rect 237 109 238 110
rect 236 109 237 110
rect 235 109 236 110
rect 234 109 235 110
rect 233 109 234 110
rect 232 109 233 110
rect 231 109 232 110
rect 230 109 231 110
rect 229 109 230 110
rect 228 109 229 110
rect 227 109 228 110
rect 226 109 227 110
rect 225 109 226 110
rect 224 109 225 110
rect 223 109 224 110
rect 222 109 223 110
rect 221 109 222 110
rect 220 109 221 110
rect 219 109 220 110
rect 218 109 219 110
rect 217 109 218 110
rect 216 109 217 110
rect 215 109 216 110
rect 214 109 215 110
rect 213 109 214 110
rect 212 109 213 110
rect 211 109 212 110
rect 210 109 211 110
rect 209 109 210 110
rect 208 109 209 110
rect 207 109 208 110
rect 206 109 207 110
rect 205 109 206 110
rect 204 109 205 110
rect 203 109 204 110
rect 202 109 203 110
rect 201 109 202 110
rect 200 109 201 110
rect 199 109 200 110
rect 198 109 199 110
rect 197 109 198 110
rect 196 109 197 110
rect 195 109 196 110
rect 194 109 195 110
rect 193 109 194 110
rect 192 109 193 110
rect 191 109 192 110
rect 190 109 191 110
rect 189 109 190 110
rect 188 109 189 110
rect 187 109 188 110
rect 186 109 187 110
rect 185 109 186 110
rect 184 109 185 110
rect 183 109 184 110
rect 182 109 183 110
rect 181 109 182 110
rect 180 109 181 110
rect 179 109 180 110
rect 178 109 179 110
rect 177 109 178 110
rect 176 109 177 110
rect 175 109 176 110
rect 174 109 175 110
rect 155 109 156 110
rect 154 109 155 110
rect 153 109 154 110
rect 152 109 153 110
rect 151 109 152 110
rect 150 109 151 110
rect 149 109 150 110
rect 148 109 149 110
rect 147 109 148 110
rect 146 109 147 110
rect 145 109 146 110
rect 144 109 145 110
rect 143 109 144 110
rect 142 109 143 110
rect 141 109 142 110
rect 140 109 141 110
rect 139 109 140 110
rect 138 109 139 110
rect 137 109 138 110
rect 136 109 137 110
rect 135 109 136 110
rect 134 109 135 110
rect 133 109 134 110
rect 132 109 133 110
rect 131 109 132 110
rect 130 109 131 110
rect 129 109 130 110
rect 128 109 129 110
rect 127 109 128 110
rect 126 109 127 110
rect 125 109 126 110
rect 117 109 118 110
rect 116 109 117 110
rect 115 109 116 110
rect 114 109 115 110
rect 113 109 114 110
rect 112 109 113 110
rect 111 109 112 110
rect 110 109 111 110
rect 109 109 110 110
rect 108 109 109 110
rect 107 109 108 110
rect 106 109 107 110
rect 105 109 106 110
rect 104 109 105 110
rect 103 109 104 110
rect 102 109 103 110
rect 101 109 102 110
rect 100 109 101 110
rect 99 109 100 110
rect 98 109 99 110
rect 97 109 98 110
rect 96 109 97 110
rect 95 109 96 110
rect 94 109 95 110
rect 93 109 94 110
rect 92 109 93 110
rect 91 109 92 110
rect 90 109 91 110
rect 89 109 90 110
rect 88 109 89 110
rect 87 109 88 110
rect 86 109 87 110
rect 85 109 86 110
rect 84 109 85 110
rect 83 109 84 110
rect 82 109 83 110
rect 64 109 65 110
rect 63 109 64 110
rect 62 109 63 110
rect 61 109 62 110
rect 60 109 61 110
rect 59 109 60 110
rect 58 109 59 110
rect 57 109 58 110
rect 56 109 57 110
rect 55 109 56 110
rect 54 109 55 110
rect 53 109 54 110
rect 52 109 53 110
rect 51 109 52 110
rect 50 109 51 110
rect 49 109 50 110
rect 48 109 49 110
rect 47 109 48 110
rect 46 109 47 110
rect 45 109 46 110
rect 44 109 45 110
rect 43 109 44 110
rect 42 109 43 110
rect 41 109 42 110
rect 40 109 41 110
rect 39 109 40 110
rect 38 109 39 110
rect 434 110 435 111
rect 433 110 434 111
rect 432 110 433 111
rect 431 110 432 111
rect 430 110 431 111
rect 429 110 430 111
rect 428 110 429 111
rect 427 110 428 111
rect 426 110 427 111
rect 425 110 426 111
rect 424 110 425 111
rect 423 110 424 111
rect 422 110 423 111
rect 421 110 422 111
rect 420 110 421 111
rect 419 110 420 111
rect 418 110 419 111
rect 417 110 418 111
rect 416 110 417 111
rect 415 110 416 111
rect 414 110 415 111
rect 413 110 414 111
rect 412 110 413 111
rect 411 110 412 111
rect 410 110 411 111
rect 409 110 410 111
rect 408 110 409 111
rect 407 110 408 111
rect 406 110 407 111
rect 405 110 406 111
rect 404 110 405 111
rect 403 110 404 111
rect 402 110 403 111
rect 401 110 402 111
rect 400 110 401 111
rect 399 110 400 111
rect 398 110 399 111
rect 397 110 398 111
rect 396 110 397 111
rect 395 110 396 111
rect 275 110 276 111
rect 274 110 275 111
rect 273 110 274 111
rect 272 110 273 111
rect 271 110 272 111
rect 270 110 271 111
rect 269 110 270 111
rect 268 110 269 111
rect 267 110 268 111
rect 266 110 267 111
rect 265 110 266 111
rect 264 110 265 111
rect 263 110 264 111
rect 262 110 263 111
rect 261 110 262 111
rect 260 110 261 111
rect 259 110 260 111
rect 258 110 259 111
rect 257 110 258 111
rect 256 110 257 111
rect 255 110 256 111
rect 254 110 255 111
rect 253 110 254 111
rect 252 110 253 111
rect 251 110 252 111
rect 250 110 251 111
rect 249 110 250 111
rect 248 110 249 111
rect 247 110 248 111
rect 246 110 247 111
rect 245 110 246 111
rect 244 110 245 111
rect 243 110 244 111
rect 242 110 243 111
rect 241 110 242 111
rect 240 110 241 111
rect 239 110 240 111
rect 238 110 239 111
rect 237 110 238 111
rect 236 110 237 111
rect 235 110 236 111
rect 234 110 235 111
rect 233 110 234 111
rect 232 110 233 111
rect 231 110 232 111
rect 230 110 231 111
rect 229 110 230 111
rect 228 110 229 111
rect 227 110 228 111
rect 226 110 227 111
rect 225 110 226 111
rect 224 110 225 111
rect 223 110 224 111
rect 222 110 223 111
rect 221 110 222 111
rect 220 110 221 111
rect 219 110 220 111
rect 218 110 219 111
rect 217 110 218 111
rect 216 110 217 111
rect 215 110 216 111
rect 214 110 215 111
rect 213 110 214 111
rect 212 110 213 111
rect 211 110 212 111
rect 210 110 211 111
rect 209 110 210 111
rect 208 110 209 111
rect 207 110 208 111
rect 206 110 207 111
rect 205 110 206 111
rect 204 110 205 111
rect 203 110 204 111
rect 202 110 203 111
rect 201 110 202 111
rect 200 110 201 111
rect 199 110 200 111
rect 198 110 199 111
rect 197 110 198 111
rect 196 110 197 111
rect 195 110 196 111
rect 194 110 195 111
rect 193 110 194 111
rect 192 110 193 111
rect 191 110 192 111
rect 190 110 191 111
rect 189 110 190 111
rect 188 110 189 111
rect 187 110 188 111
rect 186 110 187 111
rect 185 110 186 111
rect 184 110 185 111
rect 183 110 184 111
rect 182 110 183 111
rect 181 110 182 111
rect 180 110 181 111
rect 179 110 180 111
rect 178 110 179 111
rect 177 110 178 111
rect 176 110 177 111
rect 175 110 176 111
rect 174 110 175 111
rect 173 110 174 111
rect 155 110 156 111
rect 154 110 155 111
rect 153 110 154 111
rect 152 110 153 111
rect 151 110 152 111
rect 150 110 151 111
rect 149 110 150 111
rect 148 110 149 111
rect 147 110 148 111
rect 146 110 147 111
rect 145 110 146 111
rect 144 110 145 111
rect 143 110 144 111
rect 142 110 143 111
rect 141 110 142 111
rect 140 110 141 111
rect 139 110 140 111
rect 138 110 139 111
rect 137 110 138 111
rect 136 110 137 111
rect 135 110 136 111
rect 134 110 135 111
rect 133 110 134 111
rect 132 110 133 111
rect 131 110 132 111
rect 130 110 131 111
rect 129 110 130 111
rect 128 110 129 111
rect 127 110 128 111
rect 126 110 127 111
rect 125 110 126 111
rect 118 110 119 111
rect 117 110 118 111
rect 116 110 117 111
rect 115 110 116 111
rect 114 110 115 111
rect 113 110 114 111
rect 112 110 113 111
rect 111 110 112 111
rect 110 110 111 111
rect 109 110 110 111
rect 108 110 109 111
rect 107 110 108 111
rect 106 110 107 111
rect 105 110 106 111
rect 104 110 105 111
rect 103 110 104 111
rect 102 110 103 111
rect 101 110 102 111
rect 100 110 101 111
rect 99 110 100 111
rect 98 110 99 111
rect 97 110 98 111
rect 96 110 97 111
rect 95 110 96 111
rect 94 110 95 111
rect 93 110 94 111
rect 92 110 93 111
rect 91 110 92 111
rect 90 110 91 111
rect 89 110 90 111
rect 88 110 89 111
rect 87 110 88 111
rect 86 110 87 111
rect 85 110 86 111
rect 84 110 85 111
rect 83 110 84 111
rect 82 110 83 111
rect 64 110 65 111
rect 63 110 64 111
rect 62 110 63 111
rect 61 110 62 111
rect 60 110 61 111
rect 59 110 60 111
rect 58 110 59 111
rect 57 110 58 111
rect 56 110 57 111
rect 55 110 56 111
rect 54 110 55 111
rect 53 110 54 111
rect 52 110 53 111
rect 51 110 52 111
rect 50 110 51 111
rect 49 110 50 111
rect 48 110 49 111
rect 47 110 48 111
rect 46 110 47 111
rect 45 110 46 111
rect 44 110 45 111
rect 43 110 44 111
rect 42 110 43 111
rect 41 110 42 111
rect 40 110 41 111
rect 39 110 40 111
rect 38 110 39 111
rect 37 110 38 111
rect 480 111 481 112
rect 460 111 461 112
rect 435 111 436 112
rect 434 111 435 112
rect 433 111 434 112
rect 432 111 433 112
rect 431 111 432 112
rect 430 111 431 112
rect 429 111 430 112
rect 428 111 429 112
rect 427 111 428 112
rect 426 111 427 112
rect 425 111 426 112
rect 424 111 425 112
rect 423 111 424 112
rect 422 111 423 112
rect 421 111 422 112
rect 420 111 421 112
rect 419 111 420 112
rect 418 111 419 112
rect 417 111 418 112
rect 416 111 417 112
rect 415 111 416 112
rect 414 111 415 112
rect 413 111 414 112
rect 412 111 413 112
rect 411 111 412 112
rect 410 111 411 112
rect 409 111 410 112
rect 408 111 409 112
rect 407 111 408 112
rect 406 111 407 112
rect 405 111 406 112
rect 404 111 405 112
rect 403 111 404 112
rect 402 111 403 112
rect 401 111 402 112
rect 400 111 401 112
rect 399 111 400 112
rect 398 111 399 112
rect 397 111 398 112
rect 396 111 397 112
rect 395 111 396 112
rect 276 111 277 112
rect 275 111 276 112
rect 274 111 275 112
rect 273 111 274 112
rect 272 111 273 112
rect 271 111 272 112
rect 270 111 271 112
rect 269 111 270 112
rect 268 111 269 112
rect 267 111 268 112
rect 266 111 267 112
rect 265 111 266 112
rect 264 111 265 112
rect 263 111 264 112
rect 262 111 263 112
rect 261 111 262 112
rect 260 111 261 112
rect 259 111 260 112
rect 258 111 259 112
rect 257 111 258 112
rect 256 111 257 112
rect 255 111 256 112
rect 254 111 255 112
rect 253 111 254 112
rect 252 111 253 112
rect 251 111 252 112
rect 250 111 251 112
rect 249 111 250 112
rect 248 111 249 112
rect 247 111 248 112
rect 246 111 247 112
rect 245 111 246 112
rect 244 111 245 112
rect 243 111 244 112
rect 242 111 243 112
rect 241 111 242 112
rect 240 111 241 112
rect 239 111 240 112
rect 238 111 239 112
rect 237 111 238 112
rect 236 111 237 112
rect 235 111 236 112
rect 234 111 235 112
rect 233 111 234 112
rect 232 111 233 112
rect 231 111 232 112
rect 230 111 231 112
rect 229 111 230 112
rect 228 111 229 112
rect 227 111 228 112
rect 226 111 227 112
rect 225 111 226 112
rect 224 111 225 112
rect 223 111 224 112
rect 222 111 223 112
rect 221 111 222 112
rect 220 111 221 112
rect 219 111 220 112
rect 218 111 219 112
rect 217 111 218 112
rect 216 111 217 112
rect 215 111 216 112
rect 214 111 215 112
rect 213 111 214 112
rect 212 111 213 112
rect 211 111 212 112
rect 210 111 211 112
rect 209 111 210 112
rect 208 111 209 112
rect 207 111 208 112
rect 206 111 207 112
rect 205 111 206 112
rect 204 111 205 112
rect 203 111 204 112
rect 202 111 203 112
rect 201 111 202 112
rect 200 111 201 112
rect 199 111 200 112
rect 198 111 199 112
rect 197 111 198 112
rect 196 111 197 112
rect 195 111 196 112
rect 194 111 195 112
rect 193 111 194 112
rect 192 111 193 112
rect 191 111 192 112
rect 190 111 191 112
rect 189 111 190 112
rect 188 111 189 112
rect 187 111 188 112
rect 186 111 187 112
rect 185 111 186 112
rect 184 111 185 112
rect 183 111 184 112
rect 182 111 183 112
rect 181 111 182 112
rect 180 111 181 112
rect 179 111 180 112
rect 178 111 179 112
rect 177 111 178 112
rect 176 111 177 112
rect 175 111 176 112
rect 174 111 175 112
rect 173 111 174 112
rect 155 111 156 112
rect 154 111 155 112
rect 153 111 154 112
rect 152 111 153 112
rect 151 111 152 112
rect 150 111 151 112
rect 149 111 150 112
rect 148 111 149 112
rect 147 111 148 112
rect 146 111 147 112
rect 145 111 146 112
rect 144 111 145 112
rect 143 111 144 112
rect 142 111 143 112
rect 141 111 142 112
rect 140 111 141 112
rect 139 111 140 112
rect 138 111 139 112
rect 137 111 138 112
rect 136 111 137 112
rect 135 111 136 112
rect 134 111 135 112
rect 133 111 134 112
rect 132 111 133 112
rect 131 111 132 112
rect 130 111 131 112
rect 129 111 130 112
rect 128 111 129 112
rect 127 111 128 112
rect 126 111 127 112
rect 125 111 126 112
rect 124 111 125 112
rect 123 111 124 112
rect 120 111 121 112
rect 119 111 120 112
rect 118 111 119 112
rect 117 111 118 112
rect 116 111 117 112
rect 115 111 116 112
rect 114 111 115 112
rect 113 111 114 112
rect 112 111 113 112
rect 111 111 112 112
rect 110 111 111 112
rect 109 111 110 112
rect 108 111 109 112
rect 107 111 108 112
rect 106 111 107 112
rect 105 111 106 112
rect 104 111 105 112
rect 103 111 104 112
rect 102 111 103 112
rect 101 111 102 112
rect 100 111 101 112
rect 99 111 100 112
rect 98 111 99 112
rect 97 111 98 112
rect 96 111 97 112
rect 95 111 96 112
rect 94 111 95 112
rect 93 111 94 112
rect 92 111 93 112
rect 91 111 92 112
rect 90 111 91 112
rect 89 111 90 112
rect 88 111 89 112
rect 87 111 88 112
rect 86 111 87 112
rect 85 111 86 112
rect 84 111 85 112
rect 83 111 84 112
rect 82 111 83 112
rect 81 111 82 112
rect 63 111 64 112
rect 62 111 63 112
rect 61 111 62 112
rect 60 111 61 112
rect 59 111 60 112
rect 58 111 59 112
rect 57 111 58 112
rect 56 111 57 112
rect 55 111 56 112
rect 54 111 55 112
rect 53 111 54 112
rect 52 111 53 112
rect 51 111 52 112
rect 50 111 51 112
rect 49 111 50 112
rect 48 111 49 112
rect 47 111 48 112
rect 46 111 47 112
rect 45 111 46 112
rect 44 111 45 112
rect 43 111 44 112
rect 42 111 43 112
rect 41 111 42 112
rect 40 111 41 112
rect 39 111 40 112
rect 38 111 39 112
rect 37 111 38 112
rect 36 111 37 112
rect 480 112 481 113
rect 460 112 461 113
rect 436 112 437 113
rect 435 112 436 113
rect 434 112 435 113
rect 433 112 434 113
rect 432 112 433 113
rect 431 112 432 113
rect 430 112 431 113
rect 429 112 430 113
rect 428 112 429 113
rect 427 112 428 113
rect 426 112 427 113
rect 425 112 426 113
rect 424 112 425 113
rect 423 112 424 113
rect 422 112 423 113
rect 421 112 422 113
rect 420 112 421 113
rect 419 112 420 113
rect 418 112 419 113
rect 417 112 418 113
rect 416 112 417 113
rect 415 112 416 113
rect 414 112 415 113
rect 413 112 414 113
rect 412 112 413 113
rect 411 112 412 113
rect 410 112 411 113
rect 409 112 410 113
rect 408 112 409 113
rect 407 112 408 113
rect 406 112 407 113
rect 405 112 406 113
rect 404 112 405 113
rect 403 112 404 113
rect 402 112 403 113
rect 401 112 402 113
rect 400 112 401 113
rect 399 112 400 113
rect 398 112 399 113
rect 397 112 398 113
rect 396 112 397 113
rect 395 112 396 113
rect 277 112 278 113
rect 276 112 277 113
rect 275 112 276 113
rect 274 112 275 113
rect 273 112 274 113
rect 272 112 273 113
rect 271 112 272 113
rect 270 112 271 113
rect 269 112 270 113
rect 268 112 269 113
rect 267 112 268 113
rect 266 112 267 113
rect 265 112 266 113
rect 264 112 265 113
rect 263 112 264 113
rect 262 112 263 113
rect 261 112 262 113
rect 260 112 261 113
rect 259 112 260 113
rect 258 112 259 113
rect 257 112 258 113
rect 256 112 257 113
rect 255 112 256 113
rect 254 112 255 113
rect 253 112 254 113
rect 252 112 253 113
rect 251 112 252 113
rect 250 112 251 113
rect 249 112 250 113
rect 248 112 249 113
rect 247 112 248 113
rect 246 112 247 113
rect 245 112 246 113
rect 244 112 245 113
rect 243 112 244 113
rect 242 112 243 113
rect 241 112 242 113
rect 240 112 241 113
rect 239 112 240 113
rect 238 112 239 113
rect 237 112 238 113
rect 236 112 237 113
rect 235 112 236 113
rect 234 112 235 113
rect 233 112 234 113
rect 232 112 233 113
rect 231 112 232 113
rect 230 112 231 113
rect 229 112 230 113
rect 228 112 229 113
rect 227 112 228 113
rect 226 112 227 113
rect 225 112 226 113
rect 224 112 225 113
rect 223 112 224 113
rect 222 112 223 113
rect 221 112 222 113
rect 220 112 221 113
rect 219 112 220 113
rect 218 112 219 113
rect 217 112 218 113
rect 216 112 217 113
rect 215 112 216 113
rect 214 112 215 113
rect 213 112 214 113
rect 212 112 213 113
rect 211 112 212 113
rect 210 112 211 113
rect 209 112 210 113
rect 208 112 209 113
rect 207 112 208 113
rect 206 112 207 113
rect 205 112 206 113
rect 204 112 205 113
rect 203 112 204 113
rect 202 112 203 113
rect 201 112 202 113
rect 200 112 201 113
rect 199 112 200 113
rect 198 112 199 113
rect 197 112 198 113
rect 196 112 197 113
rect 195 112 196 113
rect 194 112 195 113
rect 193 112 194 113
rect 192 112 193 113
rect 191 112 192 113
rect 190 112 191 113
rect 189 112 190 113
rect 188 112 189 113
rect 187 112 188 113
rect 186 112 187 113
rect 185 112 186 113
rect 184 112 185 113
rect 183 112 184 113
rect 182 112 183 113
rect 181 112 182 113
rect 180 112 181 113
rect 179 112 180 113
rect 178 112 179 113
rect 177 112 178 113
rect 176 112 177 113
rect 175 112 176 113
rect 174 112 175 113
rect 173 112 174 113
rect 172 112 173 113
rect 154 112 155 113
rect 153 112 154 113
rect 152 112 153 113
rect 151 112 152 113
rect 150 112 151 113
rect 149 112 150 113
rect 148 112 149 113
rect 147 112 148 113
rect 146 112 147 113
rect 145 112 146 113
rect 144 112 145 113
rect 143 112 144 113
rect 142 112 143 113
rect 141 112 142 113
rect 140 112 141 113
rect 139 112 140 113
rect 138 112 139 113
rect 137 112 138 113
rect 136 112 137 113
rect 135 112 136 113
rect 134 112 135 113
rect 133 112 134 113
rect 132 112 133 113
rect 131 112 132 113
rect 130 112 131 113
rect 129 112 130 113
rect 128 112 129 113
rect 127 112 128 113
rect 126 112 127 113
rect 125 112 126 113
rect 124 112 125 113
rect 123 112 124 113
rect 122 112 123 113
rect 121 112 122 113
rect 120 112 121 113
rect 119 112 120 113
rect 118 112 119 113
rect 117 112 118 113
rect 116 112 117 113
rect 115 112 116 113
rect 114 112 115 113
rect 113 112 114 113
rect 112 112 113 113
rect 111 112 112 113
rect 110 112 111 113
rect 109 112 110 113
rect 108 112 109 113
rect 107 112 108 113
rect 106 112 107 113
rect 105 112 106 113
rect 104 112 105 113
rect 103 112 104 113
rect 102 112 103 113
rect 101 112 102 113
rect 100 112 101 113
rect 99 112 100 113
rect 98 112 99 113
rect 97 112 98 113
rect 96 112 97 113
rect 95 112 96 113
rect 94 112 95 113
rect 93 112 94 113
rect 92 112 93 113
rect 91 112 92 113
rect 90 112 91 113
rect 89 112 90 113
rect 88 112 89 113
rect 87 112 88 113
rect 86 112 87 113
rect 85 112 86 113
rect 84 112 85 113
rect 83 112 84 113
rect 82 112 83 113
rect 81 112 82 113
rect 80 112 81 113
rect 79 112 80 113
rect 63 112 64 113
rect 62 112 63 113
rect 61 112 62 113
rect 60 112 61 113
rect 59 112 60 113
rect 58 112 59 113
rect 57 112 58 113
rect 56 112 57 113
rect 55 112 56 113
rect 54 112 55 113
rect 53 112 54 113
rect 52 112 53 113
rect 51 112 52 113
rect 50 112 51 113
rect 49 112 50 113
rect 48 112 49 113
rect 47 112 48 113
rect 46 112 47 113
rect 45 112 46 113
rect 44 112 45 113
rect 43 112 44 113
rect 42 112 43 113
rect 41 112 42 113
rect 40 112 41 113
rect 39 112 40 113
rect 38 112 39 113
rect 37 112 38 113
rect 36 112 37 113
rect 35 112 36 113
rect 480 113 481 114
rect 479 113 480 114
rect 461 113 462 114
rect 460 113 461 114
rect 437 113 438 114
rect 436 113 437 114
rect 435 113 436 114
rect 434 113 435 114
rect 433 113 434 114
rect 432 113 433 114
rect 431 113 432 114
rect 430 113 431 114
rect 429 113 430 114
rect 428 113 429 114
rect 427 113 428 114
rect 426 113 427 114
rect 425 113 426 114
rect 424 113 425 114
rect 423 113 424 114
rect 422 113 423 114
rect 421 113 422 114
rect 420 113 421 114
rect 419 113 420 114
rect 418 113 419 114
rect 417 113 418 114
rect 416 113 417 114
rect 415 113 416 114
rect 414 113 415 114
rect 413 113 414 114
rect 412 113 413 114
rect 411 113 412 114
rect 410 113 411 114
rect 409 113 410 114
rect 408 113 409 114
rect 407 113 408 114
rect 406 113 407 114
rect 405 113 406 114
rect 404 113 405 114
rect 403 113 404 114
rect 402 113 403 114
rect 401 113 402 114
rect 400 113 401 114
rect 399 113 400 114
rect 398 113 399 114
rect 397 113 398 114
rect 396 113 397 114
rect 395 113 396 114
rect 265 113 266 114
rect 264 113 265 114
rect 263 113 264 114
rect 262 113 263 114
rect 261 113 262 114
rect 260 113 261 114
rect 259 113 260 114
rect 258 113 259 114
rect 257 113 258 114
rect 256 113 257 114
rect 255 113 256 114
rect 254 113 255 114
rect 253 113 254 114
rect 252 113 253 114
rect 251 113 252 114
rect 250 113 251 114
rect 249 113 250 114
rect 248 113 249 114
rect 247 113 248 114
rect 246 113 247 114
rect 245 113 246 114
rect 244 113 245 114
rect 243 113 244 114
rect 242 113 243 114
rect 241 113 242 114
rect 240 113 241 114
rect 239 113 240 114
rect 238 113 239 114
rect 237 113 238 114
rect 236 113 237 114
rect 235 113 236 114
rect 234 113 235 114
rect 233 113 234 114
rect 232 113 233 114
rect 231 113 232 114
rect 230 113 231 114
rect 229 113 230 114
rect 228 113 229 114
rect 227 113 228 114
rect 226 113 227 114
rect 225 113 226 114
rect 224 113 225 114
rect 223 113 224 114
rect 222 113 223 114
rect 221 113 222 114
rect 220 113 221 114
rect 219 113 220 114
rect 218 113 219 114
rect 217 113 218 114
rect 216 113 217 114
rect 215 113 216 114
rect 214 113 215 114
rect 213 113 214 114
rect 212 113 213 114
rect 211 113 212 114
rect 210 113 211 114
rect 209 113 210 114
rect 208 113 209 114
rect 207 113 208 114
rect 206 113 207 114
rect 205 113 206 114
rect 204 113 205 114
rect 203 113 204 114
rect 202 113 203 114
rect 201 113 202 114
rect 200 113 201 114
rect 199 113 200 114
rect 198 113 199 114
rect 197 113 198 114
rect 196 113 197 114
rect 195 113 196 114
rect 194 113 195 114
rect 193 113 194 114
rect 192 113 193 114
rect 191 113 192 114
rect 190 113 191 114
rect 189 113 190 114
rect 188 113 189 114
rect 187 113 188 114
rect 186 113 187 114
rect 185 113 186 114
rect 184 113 185 114
rect 183 113 184 114
rect 182 113 183 114
rect 181 113 182 114
rect 180 113 181 114
rect 179 113 180 114
rect 178 113 179 114
rect 177 113 178 114
rect 176 113 177 114
rect 175 113 176 114
rect 174 113 175 114
rect 173 113 174 114
rect 172 113 173 114
rect 154 113 155 114
rect 153 113 154 114
rect 152 113 153 114
rect 151 113 152 114
rect 150 113 151 114
rect 149 113 150 114
rect 148 113 149 114
rect 147 113 148 114
rect 146 113 147 114
rect 145 113 146 114
rect 144 113 145 114
rect 143 113 144 114
rect 142 113 143 114
rect 141 113 142 114
rect 140 113 141 114
rect 139 113 140 114
rect 138 113 139 114
rect 137 113 138 114
rect 136 113 137 114
rect 135 113 136 114
rect 134 113 135 114
rect 133 113 134 114
rect 132 113 133 114
rect 131 113 132 114
rect 130 113 131 114
rect 129 113 130 114
rect 128 113 129 114
rect 127 113 128 114
rect 126 113 127 114
rect 125 113 126 114
rect 124 113 125 114
rect 123 113 124 114
rect 122 113 123 114
rect 121 113 122 114
rect 120 113 121 114
rect 119 113 120 114
rect 118 113 119 114
rect 117 113 118 114
rect 116 113 117 114
rect 115 113 116 114
rect 114 113 115 114
rect 113 113 114 114
rect 112 113 113 114
rect 111 113 112 114
rect 110 113 111 114
rect 109 113 110 114
rect 108 113 109 114
rect 107 113 108 114
rect 106 113 107 114
rect 105 113 106 114
rect 104 113 105 114
rect 103 113 104 114
rect 102 113 103 114
rect 101 113 102 114
rect 100 113 101 114
rect 99 113 100 114
rect 98 113 99 114
rect 97 113 98 114
rect 96 113 97 114
rect 95 113 96 114
rect 94 113 95 114
rect 93 113 94 114
rect 92 113 93 114
rect 91 113 92 114
rect 90 113 91 114
rect 89 113 90 114
rect 88 113 89 114
rect 87 113 88 114
rect 86 113 87 114
rect 85 113 86 114
rect 84 113 85 114
rect 83 113 84 114
rect 82 113 83 114
rect 81 113 82 114
rect 80 113 81 114
rect 79 113 80 114
rect 78 113 79 114
rect 77 113 78 114
rect 63 113 64 114
rect 62 113 63 114
rect 61 113 62 114
rect 60 113 61 114
rect 59 113 60 114
rect 58 113 59 114
rect 57 113 58 114
rect 56 113 57 114
rect 55 113 56 114
rect 54 113 55 114
rect 53 113 54 114
rect 52 113 53 114
rect 51 113 52 114
rect 50 113 51 114
rect 49 113 50 114
rect 48 113 49 114
rect 47 113 48 114
rect 46 113 47 114
rect 45 113 46 114
rect 44 113 45 114
rect 43 113 44 114
rect 42 113 43 114
rect 41 113 42 114
rect 40 113 41 114
rect 39 113 40 114
rect 38 113 39 114
rect 37 113 38 114
rect 36 113 37 114
rect 35 113 36 114
rect 34 113 35 114
rect 480 114 481 115
rect 479 114 480 115
rect 478 114 479 115
rect 477 114 478 115
rect 476 114 477 115
rect 475 114 476 115
rect 474 114 475 115
rect 473 114 474 115
rect 472 114 473 115
rect 471 114 472 115
rect 470 114 471 115
rect 469 114 470 115
rect 468 114 469 115
rect 467 114 468 115
rect 466 114 467 115
rect 465 114 466 115
rect 464 114 465 115
rect 463 114 464 115
rect 462 114 463 115
rect 461 114 462 115
rect 460 114 461 115
rect 438 114 439 115
rect 437 114 438 115
rect 436 114 437 115
rect 435 114 436 115
rect 434 114 435 115
rect 433 114 434 115
rect 432 114 433 115
rect 431 114 432 115
rect 430 114 431 115
rect 429 114 430 115
rect 428 114 429 115
rect 427 114 428 115
rect 426 114 427 115
rect 425 114 426 115
rect 424 114 425 115
rect 423 114 424 115
rect 422 114 423 115
rect 421 114 422 115
rect 420 114 421 115
rect 419 114 420 115
rect 418 114 419 115
rect 417 114 418 115
rect 416 114 417 115
rect 415 114 416 115
rect 414 114 415 115
rect 413 114 414 115
rect 412 114 413 115
rect 411 114 412 115
rect 410 114 411 115
rect 409 114 410 115
rect 408 114 409 115
rect 407 114 408 115
rect 406 114 407 115
rect 405 114 406 115
rect 404 114 405 115
rect 403 114 404 115
rect 402 114 403 115
rect 401 114 402 115
rect 400 114 401 115
rect 399 114 400 115
rect 398 114 399 115
rect 397 114 398 115
rect 396 114 397 115
rect 395 114 396 115
rect 257 114 258 115
rect 256 114 257 115
rect 255 114 256 115
rect 254 114 255 115
rect 253 114 254 115
rect 252 114 253 115
rect 251 114 252 115
rect 250 114 251 115
rect 249 114 250 115
rect 248 114 249 115
rect 247 114 248 115
rect 246 114 247 115
rect 245 114 246 115
rect 244 114 245 115
rect 243 114 244 115
rect 242 114 243 115
rect 241 114 242 115
rect 240 114 241 115
rect 239 114 240 115
rect 238 114 239 115
rect 237 114 238 115
rect 236 114 237 115
rect 235 114 236 115
rect 234 114 235 115
rect 233 114 234 115
rect 232 114 233 115
rect 231 114 232 115
rect 230 114 231 115
rect 229 114 230 115
rect 228 114 229 115
rect 227 114 228 115
rect 226 114 227 115
rect 225 114 226 115
rect 224 114 225 115
rect 223 114 224 115
rect 222 114 223 115
rect 221 114 222 115
rect 220 114 221 115
rect 219 114 220 115
rect 218 114 219 115
rect 217 114 218 115
rect 216 114 217 115
rect 215 114 216 115
rect 214 114 215 115
rect 213 114 214 115
rect 212 114 213 115
rect 211 114 212 115
rect 210 114 211 115
rect 209 114 210 115
rect 208 114 209 115
rect 207 114 208 115
rect 206 114 207 115
rect 205 114 206 115
rect 204 114 205 115
rect 203 114 204 115
rect 202 114 203 115
rect 201 114 202 115
rect 200 114 201 115
rect 199 114 200 115
rect 198 114 199 115
rect 197 114 198 115
rect 196 114 197 115
rect 195 114 196 115
rect 194 114 195 115
rect 193 114 194 115
rect 192 114 193 115
rect 191 114 192 115
rect 190 114 191 115
rect 189 114 190 115
rect 188 114 189 115
rect 187 114 188 115
rect 186 114 187 115
rect 185 114 186 115
rect 184 114 185 115
rect 183 114 184 115
rect 182 114 183 115
rect 181 114 182 115
rect 180 114 181 115
rect 179 114 180 115
rect 178 114 179 115
rect 177 114 178 115
rect 176 114 177 115
rect 175 114 176 115
rect 174 114 175 115
rect 173 114 174 115
rect 172 114 173 115
rect 171 114 172 115
rect 153 114 154 115
rect 152 114 153 115
rect 151 114 152 115
rect 150 114 151 115
rect 149 114 150 115
rect 148 114 149 115
rect 147 114 148 115
rect 146 114 147 115
rect 145 114 146 115
rect 144 114 145 115
rect 143 114 144 115
rect 142 114 143 115
rect 141 114 142 115
rect 140 114 141 115
rect 139 114 140 115
rect 138 114 139 115
rect 137 114 138 115
rect 136 114 137 115
rect 135 114 136 115
rect 134 114 135 115
rect 133 114 134 115
rect 132 114 133 115
rect 131 114 132 115
rect 130 114 131 115
rect 129 114 130 115
rect 128 114 129 115
rect 127 114 128 115
rect 126 114 127 115
rect 125 114 126 115
rect 124 114 125 115
rect 123 114 124 115
rect 122 114 123 115
rect 121 114 122 115
rect 120 114 121 115
rect 119 114 120 115
rect 118 114 119 115
rect 117 114 118 115
rect 116 114 117 115
rect 115 114 116 115
rect 114 114 115 115
rect 113 114 114 115
rect 112 114 113 115
rect 111 114 112 115
rect 110 114 111 115
rect 109 114 110 115
rect 108 114 109 115
rect 107 114 108 115
rect 106 114 107 115
rect 105 114 106 115
rect 104 114 105 115
rect 103 114 104 115
rect 102 114 103 115
rect 101 114 102 115
rect 100 114 101 115
rect 99 114 100 115
rect 98 114 99 115
rect 97 114 98 115
rect 96 114 97 115
rect 95 114 96 115
rect 94 114 95 115
rect 93 114 94 115
rect 92 114 93 115
rect 91 114 92 115
rect 90 114 91 115
rect 89 114 90 115
rect 88 114 89 115
rect 87 114 88 115
rect 86 114 87 115
rect 85 114 86 115
rect 84 114 85 115
rect 83 114 84 115
rect 82 114 83 115
rect 81 114 82 115
rect 80 114 81 115
rect 79 114 80 115
rect 78 114 79 115
rect 77 114 78 115
rect 76 114 77 115
rect 75 114 76 115
rect 62 114 63 115
rect 61 114 62 115
rect 60 114 61 115
rect 59 114 60 115
rect 58 114 59 115
rect 57 114 58 115
rect 56 114 57 115
rect 55 114 56 115
rect 54 114 55 115
rect 53 114 54 115
rect 52 114 53 115
rect 51 114 52 115
rect 50 114 51 115
rect 49 114 50 115
rect 48 114 49 115
rect 47 114 48 115
rect 46 114 47 115
rect 45 114 46 115
rect 44 114 45 115
rect 43 114 44 115
rect 42 114 43 115
rect 41 114 42 115
rect 40 114 41 115
rect 39 114 40 115
rect 38 114 39 115
rect 37 114 38 115
rect 36 114 37 115
rect 35 114 36 115
rect 34 114 35 115
rect 33 114 34 115
rect 480 115 481 116
rect 479 115 480 116
rect 478 115 479 116
rect 477 115 478 116
rect 476 115 477 116
rect 475 115 476 116
rect 474 115 475 116
rect 473 115 474 116
rect 472 115 473 116
rect 471 115 472 116
rect 470 115 471 116
rect 469 115 470 116
rect 468 115 469 116
rect 467 115 468 116
rect 466 115 467 116
rect 465 115 466 116
rect 464 115 465 116
rect 463 115 464 116
rect 462 115 463 116
rect 461 115 462 116
rect 460 115 461 116
rect 438 115 439 116
rect 437 115 438 116
rect 436 115 437 116
rect 435 115 436 116
rect 434 115 435 116
rect 433 115 434 116
rect 432 115 433 116
rect 431 115 432 116
rect 430 115 431 116
rect 429 115 430 116
rect 428 115 429 116
rect 427 115 428 116
rect 426 115 427 116
rect 425 115 426 116
rect 424 115 425 116
rect 423 115 424 116
rect 422 115 423 116
rect 421 115 422 116
rect 420 115 421 116
rect 419 115 420 116
rect 418 115 419 116
rect 417 115 418 116
rect 416 115 417 116
rect 415 115 416 116
rect 414 115 415 116
rect 413 115 414 116
rect 412 115 413 116
rect 411 115 412 116
rect 410 115 411 116
rect 409 115 410 116
rect 408 115 409 116
rect 407 115 408 116
rect 406 115 407 116
rect 405 115 406 116
rect 404 115 405 116
rect 403 115 404 116
rect 402 115 403 116
rect 401 115 402 116
rect 400 115 401 116
rect 399 115 400 116
rect 398 115 399 116
rect 397 115 398 116
rect 396 115 397 116
rect 395 115 396 116
rect 253 115 254 116
rect 252 115 253 116
rect 251 115 252 116
rect 250 115 251 116
rect 249 115 250 116
rect 248 115 249 116
rect 247 115 248 116
rect 246 115 247 116
rect 245 115 246 116
rect 244 115 245 116
rect 243 115 244 116
rect 242 115 243 116
rect 241 115 242 116
rect 240 115 241 116
rect 239 115 240 116
rect 238 115 239 116
rect 237 115 238 116
rect 236 115 237 116
rect 235 115 236 116
rect 234 115 235 116
rect 233 115 234 116
rect 232 115 233 116
rect 231 115 232 116
rect 230 115 231 116
rect 229 115 230 116
rect 228 115 229 116
rect 227 115 228 116
rect 226 115 227 116
rect 225 115 226 116
rect 224 115 225 116
rect 223 115 224 116
rect 222 115 223 116
rect 221 115 222 116
rect 220 115 221 116
rect 219 115 220 116
rect 218 115 219 116
rect 217 115 218 116
rect 216 115 217 116
rect 215 115 216 116
rect 214 115 215 116
rect 213 115 214 116
rect 212 115 213 116
rect 211 115 212 116
rect 210 115 211 116
rect 209 115 210 116
rect 208 115 209 116
rect 207 115 208 116
rect 206 115 207 116
rect 205 115 206 116
rect 204 115 205 116
rect 203 115 204 116
rect 202 115 203 116
rect 201 115 202 116
rect 200 115 201 116
rect 199 115 200 116
rect 198 115 199 116
rect 197 115 198 116
rect 196 115 197 116
rect 195 115 196 116
rect 194 115 195 116
rect 193 115 194 116
rect 192 115 193 116
rect 191 115 192 116
rect 190 115 191 116
rect 189 115 190 116
rect 188 115 189 116
rect 187 115 188 116
rect 186 115 187 116
rect 185 115 186 116
rect 184 115 185 116
rect 183 115 184 116
rect 182 115 183 116
rect 181 115 182 116
rect 180 115 181 116
rect 179 115 180 116
rect 178 115 179 116
rect 177 115 178 116
rect 176 115 177 116
rect 175 115 176 116
rect 174 115 175 116
rect 173 115 174 116
rect 172 115 173 116
rect 171 115 172 116
rect 153 115 154 116
rect 152 115 153 116
rect 151 115 152 116
rect 150 115 151 116
rect 149 115 150 116
rect 148 115 149 116
rect 147 115 148 116
rect 146 115 147 116
rect 145 115 146 116
rect 144 115 145 116
rect 143 115 144 116
rect 142 115 143 116
rect 141 115 142 116
rect 140 115 141 116
rect 139 115 140 116
rect 138 115 139 116
rect 137 115 138 116
rect 136 115 137 116
rect 135 115 136 116
rect 134 115 135 116
rect 133 115 134 116
rect 132 115 133 116
rect 131 115 132 116
rect 130 115 131 116
rect 129 115 130 116
rect 128 115 129 116
rect 127 115 128 116
rect 126 115 127 116
rect 125 115 126 116
rect 124 115 125 116
rect 123 115 124 116
rect 122 115 123 116
rect 121 115 122 116
rect 120 115 121 116
rect 119 115 120 116
rect 118 115 119 116
rect 117 115 118 116
rect 116 115 117 116
rect 115 115 116 116
rect 114 115 115 116
rect 113 115 114 116
rect 112 115 113 116
rect 111 115 112 116
rect 110 115 111 116
rect 109 115 110 116
rect 108 115 109 116
rect 107 115 108 116
rect 106 115 107 116
rect 105 115 106 116
rect 104 115 105 116
rect 103 115 104 116
rect 102 115 103 116
rect 101 115 102 116
rect 100 115 101 116
rect 99 115 100 116
rect 98 115 99 116
rect 97 115 98 116
rect 96 115 97 116
rect 95 115 96 116
rect 94 115 95 116
rect 93 115 94 116
rect 92 115 93 116
rect 91 115 92 116
rect 90 115 91 116
rect 89 115 90 116
rect 88 115 89 116
rect 87 115 88 116
rect 86 115 87 116
rect 85 115 86 116
rect 84 115 85 116
rect 83 115 84 116
rect 82 115 83 116
rect 81 115 82 116
rect 80 115 81 116
rect 79 115 80 116
rect 78 115 79 116
rect 77 115 78 116
rect 76 115 77 116
rect 75 115 76 116
rect 74 115 75 116
rect 62 115 63 116
rect 61 115 62 116
rect 60 115 61 116
rect 59 115 60 116
rect 58 115 59 116
rect 57 115 58 116
rect 56 115 57 116
rect 55 115 56 116
rect 54 115 55 116
rect 53 115 54 116
rect 52 115 53 116
rect 51 115 52 116
rect 50 115 51 116
rect 49 115 50 116
rect 48 115 49 116
rect 47 115 48 116
rect 46 115 47 116
rect 45 115 46 116
rect 44 115 45 116
rect 43 115 44 116
rect 42 115 43 116
rect 41 115 42 116
rect 40 115 41 116
rect 39 115 40 116
rect 38 115 39 116
rect 37 115 38 116
rect 36 115 37 116
rect 35 115 36 116
rect 34 115 35 116
rect 33 115 34 116
rect 32 115 33 116
rect 480 116 481 117
rect 479 116 480 117
rect 478 116 479 117
rect 465 116 466 117
rect 464 116 465 117
rect 463 116 464 117
rect 462 116 463 117
rect 461 116 462 117
rect 460 116 461 117
rect 439 116 440 117
rect 438 116 439 117
rect 437 116 438 117
rect 436 116 437 117
rect 435 116 436 117
rect 434 116 435 117
rect 433 116 434 117
rect 432 116 433 117
rect 431 116 432 117
rect 430 116 431 117
rect 429 116 430 117
rect 428 116 429 117
rect 427 116 428 117
rect 426 116 427 117
rect 425 116 426 117
rect 424 116 425 117
rect 423 116 424 117
rect 422 116 423 117
rect 421 116 422 117
rect 420 116 421 117
rect 419 116 420 117
rect 418 116 419 117
rect 417 116 418 117
rect 416 116 417 117
rect 415 116 416 117
rect 414 116 415 117
rect 413 116 414 117
rect 412 116 413 117
rect 411 116 412 117
rect 410 116 411 117
rect 409 116 410 117
rect 408 116 409 117
rect 407 116 408 117
rect 406 116 407 117
rect 405 116 406 117
rect 404 116 405 117
rect 403 116 404 117
rect 402 116 403 117
rect 401 116 402 117
rect 400 116 401 117
rect 399 116 400 117
rect 398 116 399 117
rect 397 116 398 117
rect 396 116 397 117
rect 395 116 396 117
rect 249 116 250 117
rect 248 116 249 117
rect 247 116 248 117
rect 246 116 247 117
rect 245 116 246 117
rect 244 116 245 117
rect 243 116 244 117
rect 242 116 243 117
rect 241 116 242 117
rect 240 116 241 117
rect 239 116 240 117
rect 238 116 239 117
rect 237 116 238 117
rect 236 116 237 117
rect 235 116 236 117
rect 234 116 235 117
rect 233 116 234 117
rect 232 116 233 117
rect 231 116 232 117
rect 230 116 231 117
rect 229 116 230 117
rect 228 116 229 117
rect 227 116 228 117
rect 226 116 227 117
rect 225 116 226 117
rect 224 116 225 117
rect 223 116 224 117
rect 222 116 223 117
rect 221 116 222 117
rect 220 116 221 117
rect 219 116 220 117
rect 218 116 219 117
rect 217 116 218 117
rect 216 116 217 117
rect 215 116 216 117
rect 214 116 215 117
rect 213 116 214 117
rect 212 116 213 117
rect 211 116 212 117
rect 210 116 211 117
rect 209 116 210 117
rect 208 116 209 117
rect 207 116 208 117
rect 206 116 207 117
rect 205 116 206 117
rect 204 116 205 117
rect 203 116 204 117
rect 202 116 203 117
rect 201 116 202 117
rect 200 116 201 117
rect 199 116 200 117
rect 198 116 199 117
rect 197 116 198 117
rect 196 116 197 117
rect 195 116 196 117
rect 194 116 195 117
rect 193 116 194 117
rect 192 116 193 117
rect 191 116 192 117
rect 190 116 191 117
rect 189 116 190 117
rect 188 116 189 117
rect 187 116 188 117
rect 186 116 187 117
rect 185 116 186 117
rect 184 116 185 117
rect 183 116 184 117
rect 182 116 183 117
rect 181 116 182 117
rect 180 116 181 117
rect 179 116 180 117
rect 178 116 179 117
rect 177 116 178 117
rect 176 116 177 117
rect 175 116 176 117
rect 174 116 175 117
rect 173 116 174 117
rect 172 116 173 117
rect 171 116 172 117
rect 170 116 171 117
rect 153 116 154 117
rect 152 116 153 117
rect 151 116 152 117
rect 150 116 151 117
rect 149 116 150 117
rect 148 116 149 117
rect 147 116 148 117
rect 146 116 147 117
rect 145 116 146 117
rect 144 116 145 117
rect 143 116 144 117
rect 142 116 143 117
rect 141 116 142 117
rect 140 116 141 117
rect 139 116 140 117
rect 138 116 139 117
rect 137 116 138 117
rect 136 116 137 117
rect 135 116 136 117
rect 134 116 135 117
rect 133 116 134 117
rect 132 116 133 117
rect 131 116 132 117
rect 130 116 131 117
rect 129 116 130 117
rect 128 116 129 117
rect 127 116 128 117
rect 126 116 127 117
rect 125 116 126 117
rect 124 116 125 117
rect 123 116 124 117
rect 122 116 123 117
rect 121 116 122 117
rect 120 116 121 117
rect 119 116 120 117
rect 118 116 119 117
rect 117 116 118 117
rect 116 116 117 117
rect 115 116 116 117
rect 114 116 115 117
rect 113 116 114 117
rect 112 116 113 117
rect 111 116 112 117
rect 110 116 111 117
rect 109 116 110 117
rect 108 116 109 117
rect 107 116 108 117
rect 106 116 107 117
rect 105 116 106 117
rect 104 116 105 117
rect 103 116 104 117
rect 102 116 103 117
rect 101 116 102 117
rect 100 116 101 117
rect 99 116 100 117
rect 98 116 99 117
rect 97 116 98 117
rect 96 116 97 117
rect 95 116 96 117
rect 94 116 95 117
rect 93 116 94 117
rect 92 116 93 117
rect 91 116 92 117
rect 90 116 91 117
rect 89 116 90 117
rect 88 116 89 117
rect 87 116 88 117
rect 86 116 87 117
rect 85 116 86 117
rect 84 116 85 117
rect 83 116 84 117
rect 82 116 83 117
rect 81 116 82 117
rect 80 116 81 117
rect 79 116 80 117
rect 78 116 79 117
rect 77 116 78 117
rect 76 116 77 117
rect 75 116 76 117
rect 74 116 75 117
rect 73 116 74 117
rect 62 116 63 117
rect 61 116 62 117
rect 60 116 61 117
rect 59 116 60 117
rect 58 116 59 117
rect 57 116 58 117
rect 56 116 57 117
rect 55 116 56 117
rect 54 116 55 117
rect 53 116 54 117
rect 52 116 53 117
rect 51 116 52 117
rect 50 116 51 117
rect 49 116 50 117
rect 48 116 49 117
rect 47 116 48 117
rect 46 116 47 117
rect 45 116 46 117
rect 44 116 45 117
rect 43 116 44 117
rect 42 116 43 117
rect 41 116 42 117
rect 40 116 41 117
rect 39 116 40 117
rect 38 116 39 117
rect 37 116 38 117
rect 36 116 37 117
rect 35 116 36 117
rect 34 116 35 117
rect 33 116 34 117
rect 32 116 33 117
rect 480 117 481 118
rect 466 117 467 118
rect 465 117 466 118
rect 464 117 465 118
rect 463 117 464 118
rect 462 117 463 118
rect 461 117 462 118
rect 460 117 461 118
rect 439 117 440 118
rect 438 117 439 118
rect 437 117 438 118
rect 436 117 437 118
rect 435 117 436 118
rect 434 117 435 118
rect 433 117 434 118
rect 432 117 433 118
rect 431 117 432 118
rect 430 117 431 118
rect 429 117 430 118
rect 428 117 429 118
rect 427 117 428 118
rect 426 117 427 118
rect 399 117 400 118
rect 398 117 399 118
rect 397 117 398 118
rect 396 117 397 118
rect 395 117 396 118
rect 246 117 247 118
rect 245 117 246 118
rect 244 117 245 118
rect 243 117 244 118
rect 242 117 243 118
rect 241 117 242 118
rect 240 117 241 118
rect 239 117 240 118
rect 238 117 239 118
rect 237 117 238 118
rect 236 117 237 118
rect 235 117 236 118
rect 234 117 235 118
rect 233 117 234 118
rect 232 117 233 118
rect 231 117 232 118
rect 230 117 231 118
rect 229 117 230 118
rect 228 117 229 118
rect 227 117 228 118
rect 226 117 227 118
rect 225 117 226 118
rect 224 117 225 118
rect 223 117 224 118
rect 222 117 223 118
rect 221 117 222 118
rect 220 117 221 118
rect 219 117 220 118
rect 218 117 219 118
rect 217 117 218 118
rect 216 117 217 118
rect 215 117 216 118
rect 214 117 215 118
rect 213 117 214 118
rect 212 117 213 118
rect 211 117 212 118
rect 210 117 211 118
rect 209 117 210 118
rect 208 117 209 118
rect 207 117 208 118
rect 206 117 207 118
rect 205 117 206 118
rect 204 117 205 118
rect 203 117 204 118
rect 202 117 203 118
rect 201 117 202 118
rect 200 117 201 118
rect 199 117 200 118
rect 198 117 199 118
rect 197 117 198 118
rect 196 117 197 118
rect 195 117 196 118
rect 194 117 195 118
rect 193 117 194 118
rect 192 117 193 118
rect 191 117 192 118
rect 190 117 191 118
rect 189 117 190 118
rect 188 117 189 118
rect 187 117 188 118
rect 186 117 187 118
rect 185 117 186 118
rect 184 117 185 118
rect 183 117 184 118
rect 182 117 183 118
rect 181 117 182 118
rect 180 117 181 118
rect 179 117 180 118
rect 178 117 179 118
rect 177 117 178 118
rect 176 117 177 118
rect 175 117 176 118
rect 174 117 175 118
rect 173 117 174 118
rect 172 117 173 118
rect 171 117 172 118
rect 170 117 171 118
rect 152 117 153 118
rect 151 117 152 118
rect 150 117 151 118
rect 149 117 150 118
rect 148 117 149 118
rect 147 117 148 118
rect 146 117 147 118
rect 145 117 146 118
rect 144 117 145 118
rect 143 117 144 118
rect 142 117 143 118
rect 141 117 142 118
rect 140 117 141 118
rect 139 117 140 118
rect 138 117 139 118
rect 137 117 138 118
rect 136 117 137 118
rect 135 117 136 118
rect 134 117 135 118
rect 133 117 134 118
rect 132 117 133 118
rect 131 117 132 118
rect 130 117 131 118
rect 129 117 130 118
rect 128 117 129 118
rect 127 117 128 118
rect 126 117 127 118
rect 125 117 126 118
rect 124 117 125 118
rect 123 117 124 118
rect 122 117 123 118
rect 121 117 122 118
rect 120 117 121 118
rect 119 117 120 118
rect 118 117 119 118
rect 117 117 118 118
rect 116 117 117 118
rect 115 117 116 118
rect 114 117 115 118
rect 113 117 114 118
rect 112 117 113 118
rect 111 117 112 118
rect 110 117 111 118
rect 109 117 110 118
rect 108 117 109 118
rect 107 117 108 118
rect 106 117 107 118
rect 105 117 106 118
rect 104 117 105 118
rect 103 117 104 118
rect 102 117 103 118
rect 101 117 102 118
rect 100 117 101 118
rect 99 117 100 118
rect 98 117 99 118
rect 97 117 98 118
rect 96 117 97 118
rect 95 117 96 118
rect 94 117 95 118
rect 93 117 94 118
rect 92 117 93 118
rect 91 117 92 118
rect 90 117 91 118
rect 89 117 90 118
rect 88 117 89 118
rect 87 117 88 118
rect 86 117 87 118
rect 85 117 86 118
rect 84 117 85 118
rect 83 117 84 118
rect 82 117 83 118
rect 81 117 82 118
rect 80 117 81 118
rect 79 117 80 118
rect 78 117 79 118
rect 77 117 78 118
rect 76 117 77 118
rect 75 117 76 118
rect 74 117 75 118
rect 73 117 74 118
rect 72 117 73 118
rect 71 117 72 118
rect 62 117 63 118
rect 61 117 62 118
rect 60 117 61 118
rect 59 117 60 118
rect 58 117 59 118
rect 57 117 58 118
rect 56 117 57 118
rect 55 117 56 118
rect 54 117 55 118
rect 53 117 54 118
rect 52 117 53 118
rect 51 117 52 118
rect 50 117 51 118
rect 49 117 50 118
rect 48 117 49 118
rect 47 117 48 118
rect 46 117 47 118
rect 45 117 46 118
rect 44 117 45 118
rect 43 117 44 118
rect 42 117 43 118
rect 41 117 42 118
rect 40 117 41 118
rect 39 117 40 118
rect 38 117 39 118
rect 37 117 38 118
rect 36 117 37 118
rect 35 117 36 118
rect 34 117 35 118
rect 33 117 34 118
rect 32 117 33 118
rect 31 117 32 118
rect 480 118 481 119
rect 467 118 468 119
rect 466 118 467 119
rect 465 118 466 119
rect 464 118 465 119
rect 463 118 464 119
rect 462 118 463 119
rect 461 118 462 119
rect 439 118 440 119
rect 438 118 439 119
rect 437 118 438 119
rect 436 118 437 119
rect 435 118 436 119
rect 434 118 435 119
rect 433 118 434 119
rect 432 118 433 119
rect 431 118 432 119
rect 430 118 431 119
rect 398 118 399 119
rect 397 118 398 119
rect 396 118 397 119
rect 395 118 396 119
rect 244 118 245 119
rect 243 118 244 119
rect 242 118 243 119
rect 241 118 242 119
rect 240 118 241 119
rect 239 118 240 119
rect 238 118 239 119
rect 237 118 238 119
rect 236 118 237 119
rect 235 118 236 119
rect 234 118 235 119
rect 233 118 234 119
rect 232 118 233 119
rect 231 118 232 119
rect 230 118 231 119
rect 229 118 230 119
rect 228 118 229 119
rect 227 118 228 119
rect 226 118 227 119
rect 225 118 226 119
rect 224 118 225 119
rect 223 118 224 119
rect 222 118 223 119
rect 221 118 222 119
rect 220 118 221 119
rect 219 118 220 119
rect 218 118 219 119
rect 217 118 218 119
rect 216 118 217 119
rect 215 118 216 119
rect 214 118 215 119
rect 213 118 214 119
rect 212 118 213 119
rect 211 118 212 119
rect 210 118 211 119
rect 209 118 210 119
rect 208 118 209 119
rect 207 118 208 119
rect 206 118 207 119
rect 205 118 206 119
rect 204 118 205 119
rect 203 118 204 119
rect 202 118 203 119
rect 201 118 202 119
rect 200 118 201 119
rect 199 118 200 119
rect 198 118 199 119
rect 197 118 198 119
rect 196 118 197 119
rect 195 118 196 119
rect 194 118 195 119
rect 193 118 194 119
rect 192 118 193 119
rect 191 118 192 119
rect 190 118 191 119
rect 189 118 190 119
rect 188 118 189 119
rect 187 118 188 119
rect 186 118 187 119
rect 185 118 186 119
rect 184 118 185 119
rect 183 118 184 119
rect 182 118 183 119
rect 181 118 182 119
rect 180 118 181 119
rect 179 118 180 119
rect 178 118 179 119
rect 177 118 178 119
rect 176 118 177 119
rect 175 118 176 119
rect 174 118 175 119
rect 173 118 174 119
rect 172 118 173 119
rect 171 118 172 119
rect 170 118 171 119
rect 152 118 153 119
rect 151 118 152 119
rect 150 118 151 119
rect 149 118 150 119
rect 148 118 149 119
rect 147 118 148 119
rect 146 118 147 119
rect 145 118 146 119
rect 144 118 145 119
rect 143 118 144 119
rect 142 118 143 119
rect 141 118 142 119
rect 140 118 141 119
rect 139 118 140 119
rect 138 118 139 119
rect 137 118 138 119
rect 136 118 137 119
rect 135 118 136 119
rect 134 118 135 119
rect 133 118 134 119
rect 132 118 133 119
rect 131 118 132 119
rect 130 118 131 119
rect 129 118 130 119
rect 128 118 129 119
rect 127 118 128 119
rect 126 118 127 119
rect 125 118 126 119
rect 124 118 125 119
rect 123 118 124 119
rect 122 118 123 119
rect 121 118 122 119
rect 120 118 121 119
rect 119 118 120 119
rect 118 118 119 119
rect 117 118 118 119
rect 116 118 117 119
rect 115 118 116 119
rect 114 118 115 119
rect 113 118 114 119
rect 112 118 113 119
rect 111 118 112 119
rect 110 118 111 119
rect 109 118 110 119
rect 108 118 109 119
rect 107 118 108 119
rect 106 118 107 119
rect 105 118 106 119
rect 104 118 105 119
rect 103 118 104 119
rect 102 118 103 119
rect 101 118 102 119
rect 100 118 101 119
rect 99 118 100 119
rect 98 118 99 119
rect 97 118 98 119
rect 96 118 97 119
rect 95 118 96 119
rect 94 118 95 119
rect 93 118 94 119
rect 92 118 93 119
rect 91 118 92 119
rect 90 118 91 119
rect 89 118 90 119
rect 88 118 89 119
rect 87 118 88 119
rect 86 118 87 119
rect 85 118 86 119
rect 84 118 85 119
rect 83 118 84 119
rect 82 118 83 119
rect 81 118 82 119
rect 80 118 81 119
rect 79 118 80 119
rect 78 118 79 119
rect 77 118 78 119
rect 76 118 77 119
rect 75 118 76 119
rect 74 118 75 119
rect 73 118 74 119
rect 72 118 73 119
rect 71 118 72 119
rect 70 118 71 119
rect 61 118 62 119
rect 60 118 61 119
rect 59 118 60 119
rect 58 118 59 119
rect 57 118 58 119
rect 56 118 57 119
rect 55 118 56 119
rect 54 118 55 119
rect 53 118 54 119
rect 52 118 53 119
rect 51 118 52 119
rect 50 118 51 119
rect 49 118 50 119
rect 48 118 49 119
rect 47 118 48 119
rect 46 118 47 119
rect 45 118 46 119
rect 44 118 45 119
rect 43 118 44 119
rect 42 118 43 119
rect 41 118 42 119
rect 40 118 41 119
rect 39 118 40 119
rect 38 118 39 119
rect 37 118 38 119
rect 36 118 37 119
rect 35 118 36 119
rect 34 118 35 119
rect 33 118 34 119
rect 32 118 33 119
rect 31 118 32 119
rect 480 119 481 120
rect 468 119 469 120
rect 467 119 468 120
rect 466 119 467 120
rect 465 119 466 120
rect 464 119 465 120
rect 463 119 464 120
rect 462 119 463 120
rect 440 119 441 120
rect 439 119 440 120
rect 438 119 439 120
rect 437 119 438 120
rect 436 119 437 120
rect 435 119 436 120
rect 434 119 435 120
rect 433 119 434 120
rect 432 119 433 120
rect 397 119 398 120
rect 396 119 397 120
rect 395 119 396 120
rect 242 119 243 120
rect 241 119 242 120
rect 240 119 241 120
rect 239 119 240 120
rect 238 119 239 120
rect 237 119 238 120
rect 236 119 237 120
rect 235 119 236 120
rect 234 119 235 120
rect 233 119 234 120
rect 232 119 233 120
rect 231 119 232 120
rect 230 119 231 120
rect 229 119 230 120
rect 228 119 229 120
rect 227 119 228 120
rect 226 119 227 120
rect 225 119 226 120
rect 224 119 225 120
rect 223 119 224 120
rect 222 119 223 120
rect 221 119 222 120
rect 220 119 221 120
rect 219 119 220 120
rect 218 119 219 120
rect 217 119 218 120
rect 216 119 217 120
rect 215 119 216 120
rect 214 119 215 120
rect 213 119 214 120
rect 212 119 213 120
rect 211 119 212 120
rect 210 119 211 120
rect 209 119 210 120
rect 208 119 209 120
rect 207 119 208 120
rect 206 119 207 120
rect 205 119 206 120
rect 204 119 205 120
rect 203 119 204 120
rect 202 119 203 120
rect 201 119 202 120
rect 200 119 201 120
rect 199 119 200 120
rect 198 119 199 120
rect 197 119 198 120
rect 196 119 197 120
rect 195 119 196 120
rect 194 119 195 120
rect 193 119 194 120
rect 192 119 193 120
rect 191 119 192 120
rect 190 119 191 120
rect 189 119 190 120
rect 188 119 189 120
rect 187 119 188 120
rect 186 119 187 120
rect 185 119 186 120
rect 184 119 185 120
rect 183 119 184 120
rect 182 119 183 120
rect 181 119 182 120
rect 180 119 181 120
rect 179 119 180 120
rect 178 119 179 120
rect 177 119 178 120
rect 176 119 177 120
rect 175 119 176 120
rect 174 119 175 120
rect 173 119 174 120
rect 172 119 173 120
rect 171 119 172 120
rect 170 119 171 120
rect 169 119 170 120
rect 152 119 153 120
rect 151 119 152 120
rect 150 119 151 120
rect 149 119 150 120
rect 148 119 149 120
rect 147 119 148 120
rect 146 119 147 120
rect 145 119 146 120
rect 144 119 145 120
rect 143 119 144 120
rect 142 119 143 120
rect 141 119 142 120
rect 140 119 141 120
rect 139 119 140 120
rect 138 119 139 120
rect 137 119 138 120
rect 136 119 137 120
rect 135 119 136 120
rect 134 119 135 120
rect 133 119 134 120
rect 132 119 133 120
rect 131 119 132 120
rect 130 119 131 120
rect 129 119 130 120
rect 128 119 129 120
rect 127 119 128 120
rect 126 119 127 120
rect 125 119 126 120
rect 124 119 125 120
rect 123 119 124 120
rect 122 119 123 120
rect 121 119 122 120
rect 120 119 121 120
rect 119 119 120 120
rect 118 119 119 120
rect 117 119 118 120
rect 116 119 117 120
rect 115 119 116 120
rect 114 119 115 120
rect 113 119 114 120
rect 112 119 113 120
rect 111 119 112 120
rect 110 119 111 120
rect 109 119 110 120
rect 108 119 109 120
rect 107 119 108 120
rect 106 119 107 120
rect 105 119 106 120
rect 104 119 105 120
rect 103 119 104 120
rect 102 119 103 120
rect 101 119 102 120
rect 100 119 101 120
rect 99 119 100 120
rect 98 119 99 120
rect 97 119 98 120
rect 96 119 97 120
rect 95 119 96 120
rect 94 119 95 120
rect 93 119 94 120
rect 92 119 93 120
rect 91 119 92 120
rect 90 119 91 120
rect 89 119 90 120
rect 88 119 89 120
rect 87 119 88 120
rect 86 119 87 120
rect 85 119 86 120
rect 84 119 85 120
rect 83 119 84 120
rect 82 119 83 120
rect 81 119 82 120
rect 80 119 81 120
rect 79 119 80 120
rect 78 119 79 120
rect 77 119 78 120
rect 76 119 77 120
rect 75 119 76 120
rect 74 119 75 120
rect 73 119 74 120
rect 72 119 73 120
rect 71 119 72 120
rect 70 119 71 120
rect 69 119 70 120
rect 61 119 62 120
rect 60 119 61 120
rect 59 119 60 120
rect 58 119 59 120
rect 57 119 58 120
rect 56 119 57 120
rect 55 119 56 120
rect 54 119 55 120
rect 53 119 54 120
rect 52 119 53 120
rect 51 119 52 120
rect 50 119 51 120
rect 49 119 50 120
rect 48 119 49 120
rect 47 119 48 120
rect 46 119 47 120
rect 45 119 46 120
rect 44 119 45 120
rect 43 119 44 120
rect 42 119 43 120
rect 41 119 42 120
rect 40 119 41 120
rect 39 119 40 120
rect 38 119 39 120
rect 37 119 38 120
rect 36 119 37 120
rect 35 119 36 120
rect 34 119 35 120
rect 33 119 34 120
rect 32 119 33 120
rect 31 119 32 120
rect 30 119 31 120
rect 469 120 470 121
rect 468 120 469 121
rect 467 120 468 121
rect 466 120 467 121
rect 465 120 466 121
rect 464 120 465 121
rect 463 120 464 121
rect 440 120 441 121
rect 439 120 440 121
rect 438 120 439 121
rect 437 120 438 121
rect 436 120 437 121
rect 435 120 436 121
rect 434 120 435 121
rect 433 120 434 121
rect 397 120 398 121
rect 396 120 397 121
rect 395 120 396 121
rect 240 120 241 121
rect 239 120 240 121
rect 238 120 239 121
rect 237 120 238 121
rect 236 120 237 121
rect 235 120 236 121
rect 234 120 235 121
rect 233 120 234 121
rect 232 120 233 121
rect 231 120 232 121
rect 230 120 231 121
rect 229 120 230 121
rect 228 120 229 121
rect 227 120 228 121
rect 226 120 227 121
rect 225 120 226 121
rect 224 120 225 121
rect 223 120 224 121
rect 222 120 223 121
rect 221 120 222 121
rect 220 120 221 121
rect 219 120 220 121
rect 218 120 219 121
rect 217 120 218 121
rect 216 120 217 121
rect 215 120 216 121
rect 214 120 215 121
rect 213 120 214 121
rect 212 120 213 121
rect 211 120 212 121
rect 210 120 211 121
rect 209 120 210 121
rect 208 120 209 121
rect 207 120 208 121
rect 206 120 207 121
rect 205 120 206 121
rect 204 120 205 121
rect 203 120 204 121
rect 202 120 203 121
rect 201 120 202 121
rect 200 120 201 121
rect 199 120 200 121
rect 198 120 199 121
rect 197 120 198 121
rect 196 120 197 121
rect 195 120 196 121
rect 194 120 195 121
rect 193 120 194 121
rect 192 120 193 121
rect 191 120 192 121
rect 190 120 191 121
rect 189 120 190 121
rect 188 120 189 121
rect 187 120 188 121
rect 186 120 187 121
rect 185 120 186 121
rect 184 120 185 121
rect 183 120 184 121
rect 182 120 183 121
rect 181 120 182 121
rect 180 120 181 121
rect 179 120 180 121
rect 178 120 179 121
rect 177 120 178 121
rect 176 120 177 121
rect 175 120 176 121
rect 174 120 175 121
rect 173 120 174 121
rect 172 120 173 121
rect 171 120 172 121
rect 170 120 171 121
rect 169 120 170 121
rect 151 120 152 121
rect 150 120 151 121
rect 149 120 150 121
rect 148 120 149 121
rect 147 120 148 121
rect 146 120 147 121
rect 145 120 146 121
rect 144 120 145 121
rect 143 120 144 121
rect 142 120 143 121
rect 141 120 142 121
rect 140 120 141 121
rect 139 120 140 121
rect 138 120 139 121
rect 137 120 138 121
rect 136 120 137 121
rect 135 120 136 121
rect 134 120 135 121
rect 133 120 134 121
rect 132 120 133 121
rect 131 120 132 121
rect 130 120 131 121
rect 129 120 130 121
rect 128 120 129 121
rect 127 120 128 121
rect 126 120 127 121
rect 125 120 126 121
rect 124 120 125 121
rect 123 120 124 121
rect 122 120 123 121
rect 121 120 122 121
rect 120 120 121 121
rect 119 120 120 121
rect 118 120 119 121
rect 117 120 118 121
rect 116 120 117 121
rect 115 120 116 121
rect 114 120 115 121
rect 113 120 114 121
rect 112 120 113 121
rect 111 120 112 121
rect 110 120 111 121
rect 109 120 110 121
rect 108 120 109 121
rect 107 120 108 121
rect 106 120 107 121
rect 105 120 106 121
rect 104 120 105 121
rect 103 120 104 121
rect 102 120 103 121
rect 101 120 102 121
rect 100 120 101 121
rect 99 120 100 121
rect 98 120 99 121
rect 97 120 98 121
rect 96 120 97 121
rect 95 120 96 121
rect 94 120 95 121
rect 93 120 94 121
rect 92 120 93 121
rect 91 120 92 121
rect 90 120 91 121
rect 89 120 90 121
rect 88 120 89 121
rect 87 120 88 121
rect 86 120 87 121
rect 85 120 86 121
rect 84 120 85 121
rect 83 120 84 121
rect 82 120 83 121
rect 81 120 82 121
rect 80 120 81 121
rect 79 120 80 121
rect 78 120 79 121
rect 77 120 78 121
rect 76 120 77 121
rect 75 120 76 121
rect 74 120 75 121
rect 73 120 74 121
rect 72 120 73 121
rect 71 120 72 121
rect 70 120 71 121
rect 69 120 70 121
rect 61 120 62 121
rect 60 120 61 121
rect 59 120 60 121
rect 58 120 59 121
rect 57 120 58 121
rect 56 120 57 121
rect 55 120 56 121
rect 54 120 55 121
rect 53 120 54 121
rect 52 120 53 121
rect 51 120 52 121
rect 50 120 51 121
rect 49 120 50 121
rect 48 120 49 121
rect 47 120 48 121
rect 46 120 47 121
rect 45 120 46 121
rect 44 120 45 121
rect 43 120 44 121
rect 42 120 43 121
rect 41 120 42 121
rect 40 120 41 121
rect 39 120 40 121
rect 38 120 39 121
rect 37 120 38 121
rect 36 120 37 121
rect 35 120 36 121
rect 34 120 35 121
rect 33 120 34 121
rect 32 120 33 121
rect 31 120 32 121
rect 30 120 31 121
rect 471 121 472 122
rect 470 121 471 122
rect 469 121 470 122
rect 468 121 469 122
rect 467 121 468 122
rect 466 121 467 122
rect 465 121 466 122
rect 464 121 465 122
rect 440 121 441 122
rect 439 121 440 122
rect 438 121 439 122
rect 437 121 438 122
rect 436 121 437 122
rect 435 121 436 122
rect 434 121 435 122
rect 397 121 398 122
rect 396 121 397 122
rect 395 121 396 122
rect 238 121 239 122
rect 237 121 238 122
rect 236 121 237 122
rect 235 121 236 122
rect 234 121 235 122
rect 233 121 234 122
rect 232 121 233 122
rect 231 121 232 122
rect 230 121 231 122
rect 229 121 230 122
rect 228 121 229 122
rect 227 121 228 122
rect 226 121 227 122
rect 225 121 226 122
rect 224 121 225 122
rect 223 121 224 122
rect 222 121 223 122
rect 221 121 222 122
rect 220 121 221 122
rect 219 121 220 122
rect 218 121 219 122
rect 217 121 218 122
rect 216 121 217 122
rect 215 121 216 122
rect 214 121 215 122
rect 213 121 214 122
rect 212 121 213 122
rect 211 121 212 122
rect 210 121 211 122
rect 209 121 210 122
rect 208 121 209 122
rect 207 121 208 122
rect 206 121 207 122
rect 205 121 206 122
rect 204 121 205 122
rect 203 121 204 122
rect 202 121 203 122
rect 201 121 202 122
rect 200 121 201 122
rect 199 121 200 122
rect 198 121 199 122
rect 197 121 198 122
rect 196 121 197 122
rect 195 121 196 122
rect 194 121 195 122
rect 193 121 194 122
rect 192 121 193 122
rect 191 121 192 122
rect 190 121 191 122
rect 189 121 190 122
rect 188 121 189 122
rect 187 121 188 122
rect 186 121 187 122
rect 185 121 186 122
rect 184 121 185 122
rect 183 121 184 122
rect 182 121 183 122
rect 181 121 182 122
rect 180 121 181 122
rect 179 121 180 122
rect 178 121 179 122
rect 177 121 178 122
rect 176 121 177 122
rect 175 121 176 122
rect 174 121 175 122
rect 173 121 174 122
rect 172 121 173 122
rect 171 121 172 122
rect 170 121 171 122
rect 169 121 170 122
rect 168 121 169 122
rect 151 121 152 122
rect 150 121 151 122
rect 149 121 150 122
rect 148 121 149 122
rect 147 121 148 122
rect 146 121 147 122
rect 145 121 146 122
rect 144 121 145 122
rect 143 121 144 122
rect 142 121 143 122
rect 141 121 142 122
rect 140 121 141 122
rect 139 121 140 122
rect 138 121 139 122
rect 137 121 138 122
rect 136 121 137 122
rect 135 121 136 122
rect 134 121 135 122
rect 133 121 134 122
rect 132 121 133 122
rect 131 121 132 122
rect 130 121 131 122
rect 129 121 130 122
rect 128 121 129 122
rect 127 121 128 122
rect 126 121 127 122
rect 125 121 126 122
rect 124 121 125 122
rect 123 121 124 122
rect 122 121 123 122
rect 121 121 122 122
rect 120 121 121 122
rect 119 121 120 122
rect 118 121 119 122
rect 117 121 118 122
rect 116 121 117 122
rect 115 121 116 122
rect 114 121 115 122
rect 113 121 114 122
rect 112 121 113 122
rect 111 121 112 122
rect 110 121 111 122
rect 109 121 110 122
rect 108 121 109 122
rect 107 121 108 122
rect 106 121 107 122
rect 105 121 106 122
rect 104 121 105 122
rect 103 121 104 122
rect 102 121 103 122
rect 101 121 102 122
rect 100 121 101 122
rect 99 121 100 122
rect 98 121 99 122
rect 97 121 98 122
rect 96 121 97 122
rect 95 121 96 122
rect 94 121 95 122
rect 93 121 94 122
rect 92 121 93 122
rect 91 121 92 122
rect 90 121 91 122
rect 89 121 90 122
rect 88 121 89 122
rect 87 121 88 122
rect 86 121 87 122
rect 85 121 86 122
rect 84 121 85 122
rect 83 121 84 122
rect 82 121 83 122
rect 81 121 82 122
rect 80 121 81 122
rect 79 121 80 122
rect 78 121 79 122
rect 77 121 78 122
rect 76 121 77 122
rect 75 121 76 122
rect 74 121 75 122
rect 73 121 74 122
rect 72 121 73 122
rect 71 121 72 122
rect 70 121 71 122
rect 69 121 70 122
rect 68 121 69 122
rect 60 121 61 122
rect 59 121 60 122
rect 58 121 59 122
rect 57 121 58 122
rect 56 121 57 122
rect 55 121 56 122
rect 54 121 55 122
rect 53 121 54 122
rect 52 121 53 122
rect 51 121 52 122
rect 50 121 51 122
rect 49 121 50 122
rect 48 121 49 122
rect 47 121 48 122
rect 46 121 47 122
rect 45 121 46 122
rect 44 121 45 122
rect 43 121 44 122
rect 42 121 43 122
rect 41 121 42 122
rect 40 121 41 122
rect 39 121 40 122
rect 38 121 39 122
rect 37 121 38 122
rect 36 121 37 122
rect 35 121 36 122
rect 34 121 35 122
rect 33 121 34 122
rect 32 121 33 122
rect 31 121 32 122
rect 30 121 31 122
rect 472 122 473 123
rect 471 122 472 123
rect 470 122 471 123
rect 469 122 470 123
rect 468 122 469 123
rect 467 122 468 123
rect 466 122 467 123
rect 440 122 441 123
rect 439 122 440 123
rect 438 122 439 123
rect 437 122 438 123
rect 436 122 437 123
rect 435 122 436 123
rect 396 122 397 123
rect 395 122 396 123
rect 237 122 238 123
rect 236 122 237 123
rect 235 122 236 123
rect 234 122 235 123
rect 233 122 234 123
rect 232 122 233 123
rect 231 122 232 123
rect 230 122 231 123
rect 229 122 230 123
rect 228 122 229 123
rect 227 122 228 123
rect 226 122 227 123
rect 225 122 226 123
rect 224 122 225 123
rect 223 122 224 123
rect 222 122 223 123
rect 221 122 222 123
rect 220 122 221 123
rect 219 122 220 123
rect 218 122 219 123
rect 217 122 218 123
rect 216 122 217 123
rect 215 122 216 123
rect 214 122 215 123
rect 213 122 214 123
rect 212 122 213 123
rect 211 122 212 123
rect 210 122 211 123
rect 209 122 210 123
rect 208 122 209 123
rect 207 122 208 123
rect 206 122 207 123
rect 205 122 206 123
rect 204 122 205 123
rect 203 122 204 123
rect 202 122 203 123
rect 201 122 202 123
rect 200 122 201 123
rect 199 122 200 123
rect 198 122 199 123
rect 197 122 198 123
rect 196 122 197 123
rect 195 122 196 123
rect 194 122 195 123
rect 193 122 194 123
rect 192 122 193 123
rect 191 122 192 123
rect 190 122 191 123
rect 189 122 190 123
rect 188 122 189 123
rect 187 122 188 123
rect 186 122 187 123
rect 185 122 186 123
rect 184 122 185 123
rect 183 122 184 123
rect 182 122 183 123
rect 181 122 182 123
rect 180 122 181 123
rect 179 122 180 123
rect 178 122 179 123
rect 177 122 178 123
rect 176 122 177 123
rect 175 122 176 123
rect 174 122 175 123
rect 173 122 174 123
rect 172 122 173 123
rect 171 122 172 123
rect 170 122 171 123
rect 169 122 170 123
rect 168 122 169 123
rect 151 122 152 123
rect 150 122 151 123
rect 149 122 150 123
rect 148 122 149 123
rect 147 122 148 123
rect 146 122 147 123
rect 145 122 146 123
rect 144 122 145 123
rect 143 122 144 123
rect 142 122 143 123
rect 141 122 142 123
rect 140 122 141 123
rect 139 122 140 123
rect 138 122 139 123
rect 137 122 138 123
rect 136 122 137 123
rect 135 122 136 123
rect 134 122 135 123
rect 133 122 134 123
rect 132 122 133 123
rect 131 122 132 123
rect 130 122 131 123
rect 129 122 130 123
rect 128 122 129 123
rect 127 122 128 123
rect 126 122 127 123
rect 125 122 126 123
rect 124 122 125 123
rect 123 122 124 123
rect 122 122 123 123
rect 121 122 122 123
rect 120 122 121 123
rect 119 122 120 123
rect 118 122 119 123
rect 117 122 118 123
rect 116 122 117 123
rect 115 122 116 123
rect 114 122 115 123
rect 113 122 114 123
rect 112 122 113 123
rect 111 122 112 123
rect 110 122 111 123
rect 109 122 110 123
rect 108 122 109 123
rect 107 122 108 123
rect 106 122 107 123
rect 105 122 106 123
rect 104 122 105 123
rect 103 122 104 123
rect 102 122 103 123
rect 101 122 102 123
rect 100 122 101 123
rect 99 122 100 123
rect 98 122 99 123
rect 97 122 98 123
rect 96 122 97 123
rect 95 122 96 123
rect 94 122 95 123
rect 93 122 94 123
rect 92 122 93 123
rect 91 122 92 123
rect 90 122 91 123
rect 89 122 90 123
rect 88 122 89 123
rect 87 122 88 123
rect 86 122 87 123
rect 85 122 86 123
rect 84 122 85 123
rect 83 122 84 123
rect 82 122 83 123
rect 81 122 82 123
rect 80 122 81 123
rect 79 122 80 123
rect 78 122 79 123
rect 77 122 78 123
rect 76 122 77 123
rect 75 122 76 123
rect 74 122 75 123
rect 73 122 74 123
rect 72 122 73 123
rect 71 122 72 123
rect 70 122 71 123
rect 69 122 70 123
rect 68 122 69 123
rect 67 122 68 123
rect 60 122 61 123
rect 59 122 60 123
rect 58 122 59 123
rect 57 122 58 123
rect 56 122 57 123
rect 55 122 56 123
rect 54 122 55 123
rect 53 122 54 123
rect 52 122 53 123
rect 51 122 52 123
rect 50 122 51 123
rect 49 122 50 123
rect 48 122 49 123
rect 47 122 48 123
rect 46 122 47 123
rect 45 122 46 123
rect 44 122 45 123
rect 43 122 44 123
rect 42 122 43 123
rect 41 122 42 123
rect 40 122 41 123
rect 39 122 40 123
rect 38 122 39 123
rect 37 122 38 123
rect 36 122 37 123
rect 35 122 36 123
rect 34 122 35 123
rect 33 122 34 123
rect 32 122 33 123
rect 31 122 32 123
rect 30 122 31 123
rect 29 122 30 123
rect 473 123 474 124
rect 472 123 473 124
rect 471 123 472 124
rect 470 123 471 124
rect 469 123 470 124
rect 468 123 469 124
rect 467 123 468 124
rect 440 123 441 124
rect 439 123 440 124
rect 438 123 439 124
rect 437 123 438 124
rect 436 123 437 124
rect 435 123 436 124
rect 290 123 291 124
rect 289 123 290 124
rect 288 123 289 124
rect 287 123 288 124
rect 286 123 287 124
rect 285 123 286 124
rect 284 123 285 124
rect 283 123 284 124
rect 282 123 283 124
rect 281 123 282 124
rect 235 123 236 124
rect 234 123 235 124
rect 233 123 234 124
rect 232 123 233 124
rect 231 123 232 124
rect 230 123 231 124
rect 229 123 230 124
rect 228 123 229 124
rect 227 123 228 124
rect 226 123 227 124
rect 225 123 226 124
rect 224 123 225 124
rect 223 123 224 124
rect 222 123 223 124
rect 221 123 222 124
rect 220 123 221 124
rect 219 123 220 124
rect 218 123 219 124
rect 217 123 218 124
rect 216 123 217 124
rect 215 123 216 124
rect 214 123 215 124
rect 213 123 214 124
rect 212 123 213 124
rect 211 123 212 124
rect 210 123 211 124
rect 209 123 210 124
rect 208 123 209 124
rect 207 123 208 124
rect 206 123 207 124
rect 205 123 206 124
rect 204 123 205 124
rect 203 123 204 124
rect 202 123 203 124
rect 201 123 202 124
rect 200 123 201 124
rect 199 123 200 124
rect 198 123 199 124
rect 197 123 198 124
rect 196 123 197 124
rect 195 123 196 124
rect 194 123 195 124
rect 193 123 194 124
rect 192 123 193 124
rect 191 123 192 124
rect 190 123 191 124
rect 189 123 190 124
rect 188 123 189 124
rect 187 123 188 124
rect 186 123 187 124
rect 185 123 186 124
rect 184 123 185 124
rect 183 123 184 124
rect 182 123 183 124
rect 181 123 182 124
rect 180 123 181 124
rect 179 123 180 124
rect 178 123 179 124
rect 177 123 178 124
rect 176 123 177 124
rect 175 123 176 124
rect 174 123 175 124
rect 173 123 174 124
rect 172 123 173 124
rect 171 123 172 124
rect 170 123 171 124
rect 169 123 170 124
rect 168 123 169 124
rect 167 123 168 124
rect 150 123 151 124
rect 149 123 150 124
rect 148 123 149 124
rect 147 123 148 124
rect 146 123 147 124
rect 145 123 146 124
rect 144 123 145 124
rect 143 123 144 124
rect 142 123 143 124
rect 141 123 142 124
rect 140 123 141 124
rect 139 123 140 124
rect 138 123 139 124
rect 137 123 138 124
rect 136 123 137 124
rect 135 123 136 124
rect 134 123 135 124
rect 133 123 134 124
rect 132 123 133 124
rect 131 123 132 124
rect 130 123 131 124
rect 129 123 130 124
rect 128 123 129 124
rect 127 123 128 124
rect 126 123 127 124
rect 125 123 126 124
rect 124 123 125 124
rect 123 123 124 124
rect 122 123 123 124
rect 121 123 122 124
rect 120 123 121 124
rect 119 123 120 124
rect 118 123 119 124
rect 117 123 118 124
rect 116 123 117 124
rect 115 123 116 124
rect 114 123 115 124
rect 113 123 114 124
rect 112 123 113 124
rect 111 123 112 124
rect 110 123 111 124
rect 109 123 110 124
rect 108 123 109 124
rect 107 123 108 124
rect 106 123 107 124
rect 105 123 106 124
rect 104 123 105 124
rect 103 123 104 124
rect 102 123 103 124
rect 101 123 102 124
rect 100 123 101 124
rect 99 123 100 124
rect 98 123 99 124
rect 97 123 98 124
rect 96 123 97 124
rect 95 123 96 124
rect 94 123 95 124
rect 93 123 94 124
rect 92 123 93 124
rect 91 123 92 124
rect 90 123 91 124
rect 89 123 90 124
rect 88 123 89 124
rect 87 123 88 124
rect 86 123 87 124
rect 85 123 86 124
rect 84 123 85 124
rect 83 123 84 124
rect 82 123 83 124
rect 81 123 82 124
rect 80 123 81 124
rect 79 123 80 124
rect 78 123 79 124
rect 77 123 78 124
rect 76 123 77 124
rect 75 123 76 124
rect 74 123 75 124
rect 73 123 74 124
rect 72 123 73 124
rect 71 123 72 124
rect 70 123 71 124
rect 69 123 70 124
rect 68 123 69 124
rect 67 123 68 124
rect 60 123 61 124
rect 59 123 60 124
rect 58 123 59 124
rect 57 123 58 124
rect 56 123 57 124
rect 55 123 56 124
rect 54 123 55 124
rect 53 123 54 124
rect 52 123 53 124
rect 51 123 52 124
rect 50 123 51 124
rect 49 123 50 124
rect 48 123 49 124
rect 47 123 48 124
rect 46 123 47 124
rect 45 123 46 124
rect 44 123 45 124
rect 43 123 44 124
rect 42 123 43 124
rect 41 123 42 124
rect 40 123 41 124
rect 39 123 40 124
rect 38 123 39 124
rect 37 123 38 124
rect 36 123 37 124
rect 35 123 36 124
rect 34 123 35 124
rect 33 123 34 124
rect 32 123 33 124
rect 31 123 32 124
rect 30 123 31 124
rect 29 123 30 124
rect 474 124 475 125
rect 473 124 474 125
rect 472 124 473 125
rect 471 124 472 125
rect 470 124 471 125
rect 469 124 470 125
rect 468 124 469 125
rect 440 124 441 125
rect 439 124 440 125
rect 438 124 439 125
rect 437 124 438 125
rect 436 124 437 125
rect 293 124 294 125
rect 292 124 293 125
rect 291 124 292 125
rect 290 124 291 125
rect 289 124 290 125
rect 288 124 289 125
rect 287 124 288 125
rect 286 124 287 125
rect 285 124 286 125
rect 284 124 285 125
rect 283 124 284 125
rect 282 124 283 125
rect 281 124 282 125
rect 280 124 281 125
rect 279 124 280 125
rect 278 124 279 125
rect 277 124 278 125
rect 276 124 277 125
rect 234 124 235 125
rect 233 124 234 125
rect 232 124 233 125
rect 231 124 232 125
rect 230 124 231 125
rect 229 124 230 125
rect 228 124 229 125
rect 227 124 228 125
rect 226 124 227 125
rect 225 124 226 125
rect 224 124 225 125
rect 223 124 224 125
rect 222 124 223 125
rect 221 124 222 125
rect 220 124 221 125
rect 219 124 220 125
rect 218 124 219 125
rect 217 124 218 125
rect 216 124 217 125
rect 215 124 216 125
rect 214 124 215 125
rect 213 124 214 125
rect 212 124 213 125
rect 211 124 212 125
rect 210 124 211 125
rect 209 124 210 125
rect 208 124 209 125
rect 207 124 208 125
rect 206 124 207 125
rect 205 124 206 125
rect 204 124 205 125
rect 203 124 204 125
rect 202 124 203 125
rect 201 124 202 125
rect 200 124 201 125
rect 199 124 200 125
rect 198 124 199 125
rect 197 124 198 125
rect 196 124 197 125
rect 195 124 196 125
rect 194 124 195 125
rect 193 124 194 125
rect 192 124 193 125
rect 191 124 192 125
rect 190 124 191 125
rect 189 124 190 125
rect 188 124 189 125
rect 187 124 188 125
rect 186 124 187 125
rect 185 124 186 125
rect 184 124 185 125
rect 183 124 184 125
rect 182 124 183 125
rect 181 124 182 125
rect 180 124 181 125
rect 179 124 180 125
rect 178 124 179 125
rect 177 124 178 125
rect 176 124 177 125
rect 175 124 176 125
rect 174 124 175 125
rect 173 124 174 125
rect 172 124 173 125
rect 171 124 172 125
rect 170 124 171 125
rect 169 124 170 125
rect 168 124 169 125
rect 167 124 168 125
rect 150 124 151 125
rect 149 124 150 125
rect 148 124 149 125
rect 147 124 148 125
rect 146 124 147 125
rect 145 124 146 125
rect 144 124 145 125
rect 143 124 144 125
rect 142 124 143 125
rect 141 124 142 125
rect 140 124 141 125
rect 139 124 140 125
rect 138 124 139 125
rect 137 124 138 125
rect 136 124 137 125
rect 135 124 136 125
rect 134 124 135 125
rect 133 124 134 125
rect 132 124 133 125
rect 131 124 132 125
rect 130 124 131 125
rect 129 124 130 125
rect 128 124 129 125
rect 127 124 128 125
rect 126 124 127 125
rect 125 124 126 125
rect 124 124 125 125
rect 123 124 124 125
rect 122 124 123 125
rect 121 124 122 125
rect 120 124 121 125
rect 119 124 120 125
rect 118 124 119 125
rect 117 124 118 125
rect 116 124 117 125
rect 115 124 116 125
rect 114 124 115 125
rect 113 124 114 125
rect 112 124 113 125
rect 111 124 112 125
rect 110 124 111 125
rect 109 124 110 125
rect 108 124 109 125
rect 107 124 108 125
rect 106 124 107 125
rect 105 124 106 125
rect 104 124 105 125
rect 103 124 104 125
rect 102 124 103 125
rect 101 124 102 125
rect 100 124 101 125
rect 99 124 100 125
rect 98 124 99 125
rect 97 124 98 125
rect 96 124 97 125
rect 95 124 96 125
rect 94 124 95 125
rect 93 124 94 125
rect 92 124 93 125
rect 91 124 92 125
rect 90 124 91 125
rect 89 124 90 125
rect 88 124 89 125
rect 87 124 88 125
rect 86 124 87 125
rect 85 124 86 125
rect 84 124 85 125
rect 83 124 84 125
rect 82 124 83 125
rect 81 124 82 125
rect 80 124 81 125
rect 79 124 80 125
rect 78 124 79 125
rect 77 124 78 125
rect 76 124 77 125
rect 75 124 76 125
rect 74 124 75 125
rect 73 124 74 125
rect 72 124 73 125
rect 71 124 72 125
rect 70 124 71 125
rect 69 124 70 125
rect 68 124 69 125
rect 67 124 68 125
rect 66 124 67 125
rect 60 124 61 125
rect 59 124 60 125
rect 58 124 59 125
rect 57 124 58 125
rect 56 124 57 125
rect 55 124 56 125
rect 54 124 55 125
rect 53 124 54 125
rect 52 124 53 125
rect 51 124 52 125
rect 50 124 51 125
rect 49 124 50 125
rect 48 124 49 125
rect 47 124 48 125
rect 46 124 47 125
rect 45 124 46 125
rect 44 124 45 125
rect 43 124 44 125
rect 42 124 43 125
rect 41 124 42 125
rect 40 124 41 125
rect 39 124 40 125
rect 38 124 39 125
rect 37 124 38 125
rect 36 124 37 125
rect 35 124 36 125
rect 34 124 35 125
rect 33 124 34 125
rect 32 124 33 125
rect 31 124 32 125
rect 30 124 31 125
rect 29 124 30 125
rect 475 125 476 126
rect 474 125 475 126
rect 473 125 474 126
rect 472 125 473 126
rect 471 125 472 126
rect 470 125 471 126
rect 469 125 470 126
rect 440 125 441 126
rect 439 125 440 126
rect 438 125 439 126
rect 437 125 438 126
rect 436 125 437 126
rect 295 125 296 126
rect 294 125 295 126
rect 293 125 294 126
rect 292 125 293 126
rect 291 125 292 126
rect 290 125 291 126
rect 289 125 290 126
rect 288 125 289 126
rect 287 125 288 126
rect 286 125 287 126
rect 285 125 286 126
rect 284 125 285 126
rect 283 125 284 126
rect 282 125 283 126
rect 281 125 282 126
rect 280 125 281 126
rect 279 125 280 126
rect 278 125 279 126
rect 277 125 278 126
rect 276 125 277 126
rect 275 125 276 126
rect 274 125 275 126
rect 273 125 274 126
rect 272 125 273 126
rect 233 125 234 126
rect 232 125 233 126
rect 231 125 232 126
rect 230 125 231 126
rect 229 125 230 126
rect 228 125 229 126
rect 227 125 228 126
rect 226 125 227 126
rect 225 125 226 126
rect 224 125 225 126
rect 223 125 224 126
rect 222 125 223 126
rect 221 125 222 126
rect 220 125 221 126
rect 219 125 220 126
rect 218 125 219 126
rect 217 125 218 126
rect 216 125 217 126
rect 215 125 216 126
rect 214 125 215 126
rect 213 125 214 126
rect 212 125 213 126
rect 211 125 212 126
rect 210 125 211 126
rect 209 125 210 126
rect 208 125 209 126
rect 207 125 208 126
rect 206 125 207 126
rect 205 125 206 126
rect 204 125 205 126
rect 203 125 204 126
rect 202 125 203 126
rect 201 125 202 126
rect 200 125 201 126
rect 199 125 200 126
rect 198 125 199 126
rect 197 125 198 126
rect 196 125 197 126
rect 195 125 196 126
rect 194 125 195 126
rect 193 125 194 126
rect 192 125 193 126
rect 191 125 192 126
rect 190 125 191 126
rect 189 125 190 126
rect 188 125 189 126
rect 187 125 188 126
rect 186 125 187 126
rect 185 125 186 126
rect 184 125 185 126
rect 183 125 184 126
rect 182 125 183 126
rect 181 125 182 126
rect 180 125 181 126
rect 179 125 180 126
rect 178 125 179 126
rect 177 125 178 126
rect 176 125 177 126
rect 175 125 176 126
rect 174 125 175 126
rect 173 125 174 126
rect 172 125 173 126
rect 171 125 172 126
rect 170 125 171 126
rect 169 125 170 126
rect 168 125 169 126
rect 167 125 168 126
rect 149 125 150 126
rect 148 125 149 126
rect 147 125 148 126
rect 146 125 147 126
rect 145 125 146 126
rect 144 125 145 126
rect 143 125 144 126
rect 142 125 143 126
rect 141 125 142 126
rect 140 125 141 126
rect 139 125 140 126
rect 138 125 139 126
rect 137 125 138 126
rect 136 125 137 126
rect 135 125 136 126
rect 134 125 135 126
rect 133 125 134 126
rect 132 125 133 126
rect 131 125 132 126
rect 130 125 131 126
rect 129 125 130 126
rect 128 125 129 126
rect 127 125 128 126
rect 126 125 127 126
rect 125 125 126 126
rect 124 125 125 126
rect 123 125 124 126
rect 122 125 123 126
rect 121 125 122 126
rect 120 125 121 126
rect 119 125 120 126
rect 118 125 119 126
rect 117 125 118 126
rect 116 125 117 126
rect 115 125 116 126
rect 114 125 115 126
rect 113 125 114 126
rect 112 125 113 126
rect 111 125 112 126
rect 110 125 111 126
rect 109 125 110 126
rect 108 125 109 126
rect 107 125 108 126
rect 106 125 107 126
rect 105 125 106 126
rect 104 125 105 126
rect 103 125 104 126
rect 102 125 103 126
rect 101 125 102 126
rect 100 125 101 126
rect 99 125 100 126
rect 98 125 99 126
rect 97 125 98 126
rect 96 125 97 126
rect 95 125 96 126
rect 94 125 95 126
rect 93 125 94 126
rect 92 125 93 126
rect 91 125 92 126
rect 90 125 91 126
rect 89 125 90 126
rect 88 125 89 126
rect 87 125 88 126
rect 86 125 87 126
rect 85 125 86 126
rect 84 125 85 126
rect 83 125 84 126
rect 82 125 83 126
rect 81 125 82 126
rect 80 125 81 126
rect 79 125 80 126
rect 78 125 79 126
rect 77 125 78 126
rect 76 125 77 126
rect 75 125 76 126
rect 74 125 75 126
rect 73 125 74 126
rect 72 125 73 126
rect 71 125 72 126
rect 70 125 71 126
rect 69 125 70 126
rect 68 125 69 126
rect 67 125 68 126
rect 66 125 67 126
rect 59 125 60 126
rect 58 125 59 126
rect 57 125 58 126
rect 56 125 57 126
rect 55 125 56 126
rect 54 125 55 126
rect 53 125 54 126
rect 52 125 53 126
rect 51 125 52 126
rect 50 125 51 126
rect 49 125 50 126
rect 48 125 49 126
rect 47 125 48 126
rect 46 125 47 126
rect 45 125 46 126
rect 44 125 45 126
rect 43 125 44 126
rect 42 125 43 126
rect 41 125 42 126
rect 40 125 41 126
rect 39 125 40 126
rect 38 125 39 126
rect 37 125 38 126
rect 36 125 37 126
rect 35 125 36 126
rect 34 125 35 126
rect 33 125 34 126
rect 32 125 33 126
rect 31 125 32 126
rect 30 125 31 126
rect 29 125 30 126
rect 477 126 478 127
rect 476 126 477 127
rect 475 126 476 127
rect 474 126 475 127
rect 473 126 474 127
rect 472 126 473 127
rect 471 126 472 127
rect 470 126 471 127
rect 460 126 461 127
rect 440 126 441 127
rect 439 126 440 127
rect 438 126 439 127
rect 437 126 438 127
rect 436 126 437 127
rect 297 126 298 127
rect 296 126 297 127
rect 295 126 296 127
rect 294 126 295 127
rect 293 126 294 127
rect 292 126 293 127
rect 291 126 292 127
rect 290 126 291 127
rect 289 126 290 127
rect 288 126 289 127
rect 287 126 288 127
rect 286 126 287 127
rect 285 126 286 127
rect 284 126 285 127
rect 283 126 284 127
rect 282 126 283 127
rect 281 126 282 127
rect 280 126 281 127
rect 279 126 280 127
rect 278 126 279 127
rect 277 126 278 127
rect 276 126 277 127
rect 275 126 276 127
rect 274 126 275 127
rect 273 126 274 127
rect 272 126 273 127
rect 271 126 272 127
rect 270 126 271 127
rect 269 126 270 127
rect 232 126 233 127
rect 231 126 232 127
rect 230 126 231 127
rect 229 126 230 127
rect 228 126 229 127
rect 227 126 228 127
rect 226 126 227 127
rect 225 126 226 127
rect 224 126 225 127
rect 223 126 224 127
rect 222 126 223 127
rect 221 126 222 127
rect 220 126 221 127
rect 219 126 220 127
rect 218 126 219 127
rect 217 126 218 127
rect 216 126 217 127
rect 215 126 216 127
rect 214 126 215 127
rect 213 126 214 127
rect 212 126 213 127
rect 211 126 212 127
rect 210 126 211 127
rect 209 126 210 127
rect 208 126 209 127
rect 207 126 208 127
rect 206 126 207 127
rect 205 126 206 127
rect 204 126 205 127
rect 203 126 204 127
rect 202 126 203 127
rect 201 126 202 127
rect 200 126 201 127
rect 199 126 200 127
rect 198 126 199 127
rect 197 126 198 127
rect 196 126 197 127
rect 195 126 196 127
rect 194 126 195 127
rect 193 126 194 127
rect 192 126 193 127
rect 191 126 192 127
rect 190 126 191 127
rect 189 126 190 127
rect 188 126 189 127
rect 187 126 188 127
rect 186 126 187 127
rect 185 126 186 127
rect 184 126 185 127
rect 183 126 184 127
rect 182 126 183 127
rect 181 126 182 127
rect 180 126 181 127
rect 179 126 180 127
rect 178 126 179 127
rect 177 126 178 127
rect 176 126 177 127
rect 175 126 176 127
rect 174 126 175 127
rect 173 126 174 127
rect 172 126 173 127
rect 171 126 172 127
rect 170 126 171 127
rect 169 126 170 127
rect 168 126 169 127
rect 167 126 168 127
rect 166 126 167 127
rect 149 126 150 127
rect 148 126 149 127
rect 147 126 148 127
rect 146 126 147 127
rect 145 126 146 127
rect 144 126 145 127
rect 143 126 144 127
rect 142 126 143 127
rect 141 126 142 127
rect 140 126 141 127
rect 139 126 140 127
rect 138 126 139 127
rect 137 126 138 127
rect 136 126 137 127
rect 135 126 136 127
rect 134 126 135 127
rect 133 126 134 127
rect 132 126 133 127
rect 131 126 132 127
rect 130 126 131 127
rect 129 126 130 127
rect 128 126 129 127
rect 127 126 128 127
rect 126 126 127 127
rect 125 126 126 127
rect 124 126 125 127
rect 123 126 124 127
rect 122 126 123 127
rect 121 126 122 127
rect 120 126 121 127
rect 119 126 120 127
rect 118 126 119 127
rect 117 126 118 127
rect 116 126 117 127
rect 115 126 116 127
rect 114 126 115 127
rect 113 126 114 127
rect 112 126 113 127
rect 111 126 112 127
rect 110 126 111 127
rect 109 126 110 127
rect 108 126 109 127
rect 107 126 108 127
rect 106 126 107 127
rect 105 126 106 127
rect 104 126 105 127
rect 103 126 104 127
rect 102 126 103 127
rect 101 126 102 127
rect 100 126 101 127
rect 99 126 100 127
rect 98 126 99 127
rect 97 126 98 127
rect 96 126 97 127
rect 95 126 96 127
rect 94 126 95 127
rect 93 126 94 127
rect 92 126 93 127
rect 91 126 92 127
rect 90 126 91 127
rect 89 126 90 127
rect 88 126 89 127
rect 87 126 88 127
rect 86 126 87 127
rect 85 126 86 127
rect 84 126 85 127
rect 83 126 84 127
rect 82 126 83 127
rect 81 126 82 127
rect 80 126 81 127
rect 79 126 80 127
rect 78 126 79 127
rect 77 126 78 127
rect 76 126 77 127
rect 75 126 76 127
rect 74 126 75 127
rect 73 126 74 127
rect 72 126 73 127
rect 71 126 72 127
rect 70 126 71 127
rect 69 126 70 127
rect 68 126 69 127
rect 67 126 68 127
rect 66 126 67 127
rect 65 126 66 127
rect 59 126 60 127
rect 58 126 59 127
rect 57 126 58 127
rect 56 126 57 127
rect 55 126 56 127
rect 54 126 55 127
rect 53 126 54 127
rect 52 126 53 127
rect 51 126 52 127
rect 50 126 51 127
rect 49 126 50 127
rect 48 126 49 127
rect 47 126 48 127
rect 46 126 47 127
rect 45 126 46 127
rect 44 126 45 127
rect 43 126 44 127
rect 42 126 43 127
rect 41 126 42 127
rect 40 126 41 127
rect 39 126 40 127
rect 38 126 39 127
rect 37 126 38 127
rect 36 126 37 127
rect 35 126 36 127
rect 34 126 35 127
rect 33 126 34 127
rect 32 126 33 127
rect 31 126 32 127
rect 30 126 31 127
rect 29 126 30 127
rect 478 127 479 128
rect 477 127 478 128
rect 476 127 477 128
rect 475 127 476 128
rect 474 127 475 128
rect 473 127 474 128
rect 472 127 473 128
rect 471 127 472 128
rect 460 127 461 128
rect 440 127 441 128
rect 439 127 440 128
rect 438 127 439 128
rect 437 127 438 128
rect 436 127 437 128
rect 299 127 300 128
rect 298 127 299 128
rect 297 127 298 128
rect 296 127 297 128
rect 295 127 296 128
rect 294 127 295 128
rect 293 127 294 128
rect 292 127 293 128
rect 291 127 292 128
rect 290 127 291 128
rect 289 127 290 128
rect 288 127 289 128
rect 287 127 288 128
rect 286 127 287 128
rect 285 127 286 128
rect 284 127 285 128
rect 283 127 284 128
rect 282 127 283 128
rect 281 127 282 128
rect 280 127 281 128
rect 279 127 280 128
rect 278 127 279 128
rect 277 127 278 128
rect 276 127 277 128
rect 275 127 276 128
rect 274 127 275 128
rect 273 127 274 128
rect 272 127 273 128
rect 271 127 272 128
rect 270 127 271 128
rect 269 127 270 128
rect 268 127 269 128
rect 267 127 268 128
rect 266 127 267 128
rect 231 127 232 128
rect 230 127 231 128
rect 229 127 230 128
rect 228 127 229 128
rect 227 127 228 128
rect 226 127 227 128
rect 225 127 226 128
rect 224 127 225 128
rect 223 127 224 128
rect 222 127 223 128
rect 221 127 222 128
rect 220 127 221 128
rect 219 127 220 128
rect 218 127 219 128
rect 217 127 218 128
rect 216 127 217 128
rect 215 127 216 128
rect 214 127 215 128
rect 213 127 214 128
rect 212 127 213 128
rect 211 127 212 128
rect 210 127 211 128
rect 209 127 210 128
rect 208 127 209 128
rect 207 127 208 128
rect 206 127 207 128
rect 205 127 206 128
rect 204 127 205 128
rect 203 127 204 128
rect 202 127 203 128
rect 201 127 202 128
rect 200 127 201 128
rect 199 127 200 128
rect 198 127 199 128
rect 197 127 198 128
rect 196 127 197 128
rect 195 127 196 128
rect 194 127 195 128
rect 193 127 194 128
rect 192 127 193 128
rect 191 127 192 128
rect 190 127 191 128
rect 189 127 190 128
rect 188 127 189 128
rect 187 127 188 128
rect 186 127 187 128
rect 185 127 186 128
rect 184 127 185 128
rect 183 127 184 128
rect 182 127 183 128
rect 181 127 182 128
rect 180 127 181 128
rect 179 127 180 128
rect 178 127 179 128
rect 177 127 178 128
rect 176 127 177 128
rect 175 127 176 128
rect 174 127 175 128
rect 173 127 174 128
rect 172 127 173 128
rect 171 127 172 128
rect 170 127 171 128
rect 169 127 170 128
rect 168 127 169 128
rect 167 127 168 128
rect 166 127 167 128
rect 148 127 149 128
rect 147 127 148 128
rect 146 127 147 128
rect 145 127 146 128
rect 144 127 145 128
rect 143 127 144 128
rect 142 127 143 128
rect 141 127 142 128
rect 140 127 141 128
rect 139 127 140 128
rect 138 127 139 128
rect 137 127 138 128
rect 136 127 137 128
rect 135 127 136 128
rect 134 127 135 128
rect 133 127 134 128
rect 132 127 133 128
rect 131 127 132 128
rect 130 127 131 128
rect 129 127 130 128
rect 128 127 129 128
rect 127 127 128 128
rect 126 127 127 128
rect 125 127 126 128
rect 124 127 125 128
rect 123 127 124 128
rect 122 127 123 128
rect 121 127 122 128
rect 120 127 121 128
rect 119 127 120 128
rect 118 127 119 128
rect 117 127 118 128
rect 116 127 117 128
rect 115 127 116 128
rect 114 127 115 128
rect 113 127 114 128
rect 112 127 113 128
rect 111 127 112 128
rect 110 127 111 128
rect 109 127 110 128
rect 108 127 109 128
rect 107 127 108 128
rect 106 127 107 128
rect 105 127 106 128
rect 104 127 105 128
rect 103 127 104 128
rect 102 127 103 128
rect 101 127 102 128
rect 100 127 101 128
rect 99 127 100 128
rect 98 127 99 128
rect 97 127 98 128
rect 96 127 97 128
rect 95 127 96 128
rect 94 127 95 128
rect 93 127 94 128
rect 92 127 93 128
rect 91 127 92 128
rect 90 127 91 128
rect 89 127 90 128
rect 88 127 89 128
rect 87 127 88 128
rect 86 127 87 128
rect 85 127 86 128
rect 84 127 85 128
rect 83 127 84 128
rect 82 127 83 128
rect 81 127 82 128
rect 80 127 81 128
rect 79 127 80 128
rect 78 127 79 128
rect 77 127 78 128
rect 76 127 77 128
rect 75 127 76 128
rect 74 127 75 128
rect 73 127 74 128
rect 72 127 73 128
rect 71 127 72 128
rect 70 127 71 128
rect 69 127 70 128
rect 68 127 69 128
rect 67 127 68 128
rect 66 127 67 128
rect 65 127 66 128
rect 59 127 60 128
rect 58 127 59 128
rect 57 127 58 128
rect 56 127 57 128
rect 55 127 56 128
rect 54 127 55 128
rect 53 127 54 128
rect 52 127 53 128
rect 51 127 52 128
rect 50 127 51 128
rect 49 127 50 128
rect 48 127 49 128
rect 47 127 48 128
rect 46 127 47 128
rect 45 127 46 128
rect 44 127 45 128
rect 43 127 44 128
rect 42 127 43 128
rect 41 127 42 128
rect 40 127 41 128
rect 39 127 40 128
rect 38 127 39 128
rect 37 127 38 128
rect 36 127 37 128
rect 35 127 36 128
rect 34 127 35 128
rect 33 127 34 128
rect 32 127 33 128
rect 31 127 32 128
rect 30 127 31 128
rect 479 128 480 129
rect 478 128 479 129
rect 477 128 478 129
rect 476 128 477 129
rect 475 128 476 129
rect 474 128 475 129
rect 473 128 474 129
rect 472 128 473 129
rect 460 128 461 129
rect 440 128 441 129
rect 439 128 440 129
rect 438 128 439 129
rect 437 128 438 129
rect 436 128 437 129
rect 300 128 301 129
rect 299 128 300 129
rect 298 128 299 129
rect 297 128 298 129
rect 296 128 297 129
rect 295 128 296 129
rect 294 128 295 129
rect 293 128 294 129
rect 292 128 293 129
rect 291 128 292 129
rect 290 128 291 129
rect 289 128 290 129
rect 288 128 289 129
rect 287 128 288 129
rect 286 128 287 129
rect 285 128 286 129
rect 284 128 285 129
rect 283 128 284 129
rect 282 128 283 129
rect 281 128 282 129
rect 280 128 281 129
rect 279 128 280 129
rect 278 128 279 129
rect 277 128 278 129
rect 276 128 277 129
rect 275 128 276 129
rect 274 128 275 129
rect 273 128 274 129
rect 272 128 273 129
rect 271 128 272 129
rect 270 128 271 129
rect 269 128 270 129
rect 268 128 269 129
rect 267 128 268 129
rect 266 128 267 129
rect 265 128 266 129
rect 264 128 265 129
rect 230 128 231 129
rect 229 128 230 129
rect 228 128 229 129
rect 227 128 228 129
rect 226 128 227 129
rect 225 128 226 129
rect 224 128 225 129
rect 223 128 224 129
rect 222 128 223 129
rect 221 128 222 129
rect 220 128 221 129
rect 219 128 220 129
rect 218 128 219 129
rect 217 128 218 129
rect 216 128 217 129
rect 215 128 216 129
rect 214 128 215 129
rect 213 128 214 129
rect 212 128 213 129
rect 211 128 212 129
rect 210 128 211 129
rect 209 128 210 129
rect 208 128 209 129
rect 207 128 208 129
rect 206 128 207 129
rect 205 128 206 129
rect 204 128 205 129
rect 203 128 204 129
rect 202 128 203 129
rect 201 128 202 129
rect 200 128 201 129
rect 199 128 200 129
rect 198 128 199 129
rect 197 128 198 129
rect 196 128 197 129
rect 195 128 196 129
rect 194 128 195 129
rect 193 128 194 129
rect 192 128 193 129
rect 191 128 192 129
rect 190 128 191 129
rect 189 128 190 129
rect 188 128 189 129
rect 187 128 188 129
rect 186 128 187 129
rect 185 128 186 129
rect 184 128 185 129
rect 183 128 184 129
rect 182 128 183 129
rect 181 128 182 129
rect 180 128 181 129
rect 179 128 180 129
rect 178 128 179 129
rect 177 128 178 129
rect 176 128 177 129
rect 175 128 176 129
rect 174 128 175 129
rect 173 128 174 129
rect 172 128 173 129
rect 171 128 172 129
rect 170 128 171 129
rect 169 128 170 129
rect 168 128 169 129
rect 167 128 168 129
rect 166 128 167 129
rect 165 128 166 129
rect 148 128 149 129
rect 147 128 148 129
rect 146 128 147 129
rect 145 128 146 129
rect 144 128 145 129
rect 143 128 144 129
rect 142 128 143 129
rect 141 128 142 129
rect 140 128 141 129
rect 139 128 140 129
rect 138 128 139 129
rect 137 128 138 129
rect 136 128 137 129
rect 135 128 136 129
rect 134 128 135 129
rect 133 128 134 129
rect 132 128 133 129
rect 131 128 132 129
rect 130 128 131 129
rect 129 128 130 129
rect 128 128 129 129
rect 127 128 128 129
rect 126 128 127 129
rect 125 128 126 129
rect 124 128 125 129
rect 123 128 124 129
rect 122 128 123 129
rect 121 128 122 129
rect 120 128 121 129
rect 119 128 120 129
rect 118 128 119 129
rect 117 128 118 129
rect 116 128 117 129
rect 115 128 116 129
rect 114 128 115 129
rect 113 128 114 129
rect 112 128 113 129
rect 111 128 112 129
rect 110 128 111 129
rect 109 128 110 129
rect 108 128 109 129
rect 107 128 108 129
rect 106 128 107 129
rect 105 128 106 129
rect 104 128 105 129
rect 103 128 104 129
rect 102 128 103 129
rect 101 128 102 129
rect 100 128 101 129
rect 99 128 100 129
rect 98 128 99 129
rect 97 128 98 129
rect 96 128 97 129
rect 95 128 96 129
rect 94 128 95 129
rect 93 128 94 129
rect 92 128 93 129
rect 91 128 92 129
rect 90 128 91 129
rect 89 128 90 129
rect 88 128 89 129
rect 87 128 88 129
rect 86 128 87 129
rect 85 128 86 129
rect 84 128 85 129
rect 83 128 84 129
rect 82 128 83 129
rect 81 128 82 129
rect 80 128 81 129
rect 79 128 80 129
rect 78 128 79 129
rect 77 128 78 129
rect 76 128 77 129
rect 75 128 76 129
rect 74 128 75 129
rect 73 128 74 129
rect 72 128 73 129
rect 71 128 72 129
rect 70 128 71 129
rect 69 128 70 129
rect 68 128 69 129
rect 67 128 68 129
rect 66 128 67 129
rect 65 128 66 129
rect 64 128 65 129
rect 59 128 60 129
rect 58 128 59 129
rect 57 128 58 129
rect 56 128 57 129
rect 55 128 56 129
rect 54 128 55 129
rect 53 128 54 129
rect 52 128 53 129
rect 51 128 52 129
rect 50 128 51 129
rect 49 128 50 129
rect 48 128 49 129
rect 47 128 48 129
rect 46 128 47 129
rect 45 128 46 129
rect 44 128 45 129
rect 43 128 44 129
rect 42 128 43 129
rect 41 128 42 129
rect 40 128 41 129
rect 39 128 40 129
rect 38 128 39 129
rect 37 128 38 129
rect 36 128 37 129
rect 35 128 36 129
rect 34 128 35 129
rect 33 128 34 129
rect 32 128 33 129
rect 31 128 32 129
rect 30 128 31 129
rect 480 129 481 130
rect 479 129 480 130
rect 478 129 479 130
rect 477 129 478 130
rect 476 129 477 130
rect 475 129 476 130
rect 474 129 475 130
rect 473 129 474 130
rect 462 129 463 130
rect 461 129 462 130
rect 460 129 461 130
rect 440 129 441 130
rect 439 129 440 130
rect 438 129 439 130
rect 437 129 438 130
rect 436 129 437 130
rect 302 129 303 130
rect 301 129 302 130
rect 300 129 301 130
rect 299 129 300 130
rect 298 129 299 130
rect 297 129 298 130
rect 296 129 297 130
rect 295 129 296 130
rect 294 129 295 130
rect 293 129 294 130
rect 292 129 293 130
rect 291 129 292 130
rect 290 129 291 130
rect 289 129 290 130
rect 288 129 289 130
rect 287 129 288 130
rect 286 129 287 130
rect 285 129 286 130
rect 284 129 285 130
rect 283 129 284 130
rect 282 129 283 130
rect 281 129 282 130
rect 280 129 281 130
rect 279 129 280 130
rect 278 129 279 130
rect 277 129 278 130
rect 276 129 277 130
rect 275 129 276 130
rect 274 129 275 130
rect 273 129 274 130
rect 272 129 273 130
rect 271 129 272 130
rect 270 129 271 130
rect 269 129 270 130
rect 268 129 269 130
rect 267 129 268 130
rect 266 129 267 130
rect 265 129 266 130
rect 264 129 265 130
rect 263 129 264 130
rect 262 129 263 130
rect 230 129 231 130
rect 229 129 230 130
rect 228 129 229 130
rect 227 129 228 130
rect 226 129 227 130
rect 225 129 226 130
rect 224 129 225 130
rect 223 129 224 130
rect 222 129 223 130
rect 221 129 222 130
rect 220 129 221 130
rect 219 129 220 130
rect 218 129 219 130
rect 217 129 218 130
rect 216 129 217 130
rect 215 129 216 130
rect 214 129 215 130
rect 213 129 214 130
rect 212 129 213 130
rect 211 129 212 130
rect 210 129 211 130
rect 209 129 210 130
rect 208 129 209 130
rect 207 129 208 130
rect 206 129 207 130
rect 205 129 206 130
rect 204 129 205 130
rect 203 129 204 130
rect 202 129 203 130
rect 201 129 202 130
rect 200 129 201 130
rect 199 129 200 130
rect 198 129 199 130
rect 197 129 198 130
rect 196 129 197 130
rect 195 129 196 130
rect 194 129 195 130
rect 193 129 194 130
rect 192 129 193 130
rect 191 129 192 130
rect 190 129 191 130
rect 189 129 190 130
rect 188 129 189 130
rect 187 129 188 130
rect 186 129 187 130
rect 185 129 186 130
rect 184 129 185 130
rect 183 129 184 130
rect 182 129 183 130
rect 181 129 182 130
rect 180 129 181 130
rect 179 129 180 130
rect 178 129 179 130
rect 177 129 178 130
rect 176 129 177 130
rect 175 129 176 130
rect 174 129 175 130
rect 173 129 174 130
rect 172 129 173 130
rect 171 129 172 130
rect 170 129 171 130
rect 169 129 170 130
rect 168 129 169 130
rect 167 129 168 130
rect 166 129 167 130
rect 165 129 166 130
rect 147 129 148 130
rect 146 129 147 130
rect 145 129 146 130
rect 144 129 145 130
rect 143 129 144 130
rect 142 129 143 130
rect 141 129 142 130
rect 140 129 141 130
rect 139 129 140 130
rect 138 129 139 130
rect 137 129 138 130
rect 136 129 137 130
rect 135 129 136 130
rect 134 129 135 130
rect 133 129 134 130
rect 132 129 133 130
rect 131 129 132 130
rect 130 129 131 130
rect 129 129 130 130
rect 128 129 129 130
rect 127 129 128 130
rect 126 129 127 130
rect 125 129 126 130
rect 124 129 125 130
rect 123 129 124 130
rect 122 129 123 130
rect 121 129 122 130
rect 120 129 121 130
rect 119 129 120 130
rect 118 129 119 130
rect 117 129 118 130
rect 116 129 117 130
rect 115 129 116 130
rect 114 129 115 130
rect 113 129 114 130
rect 112 129 113 130
rect 111 129 112 130
rect 110 129 111 130
rect 109 129 110 130
rect 108 129 109 130
rect 107 129 108 130
rect 106 129 107 130
rect 105 129 106 130
rect 104 129 105 130
rect 103 129 104 130
rect 102 129 103 130
rect 101 129 102 130
rect 100 129 101 130
rect 99 129 100 130
rect 98 129 99 130
rect 97 129 98 130
rect 96 129 97 130
rect 95 129 96 130
rect 94 129 95 130
rect 93 129 94 130
rect 92 129 93 130
rect 91 129 92 130
rect 90 129 91 130
rect 89 129 90 130
rect 88 129 89 130
rect 87 129 88 130
rect 86 129 87 130
rect 85 129 86 130
rect 84 129 85 130
rect 83 129 84 130
rect 82 129 83 130
rect 81 129 82 130
rect 80 129 81 130
rect 79 129 80 130
rect 78 129 79 130
rect 77 129 78 130
rect 76 129 77 130
rect 75 129 76 130
rect 74 129 75 130
rect 73 129 74 130
rect 72 129 73 130
rect 71 129 72 130
rect 70 129 71 130
rect 69 129 70 130
rect 68 129 69 130
rect 67 129 68 130
rect 66 129 67 130
rect 65 129 66 130
rect 64 129 65 130
rect 63 129 64 130
rect 59 129 60 130
rect 58 129 59 130
rect 57 129 58 130
rect 56 129 57 130
rect 55 129 56 130
rect 54 129 55 130
rect 53 129 54 130
rect 52 129 53 130
rect 51 129 52 130
rect 50 129 51 130
rect 49 129 50 130
rect 48 129 49 130
rect 47 129 48 130
rect 46 129 47 130
rect 45 129 46 130
rect 44 129 45 130
rect 43 129 44 130
rect 42 129 43 130
rect 41 129 42 130
rect 40 129 41 130
rect 39 129 40 130
rect 38 129 39 130
rect 37 129 38 130
rect 36 129 37 130
rect 35 129 36 130
rect 34 129 35 130
rect 33 129 34 130
rect 32 129 33 130
rect 31 129 32 130
rect 30 129 31 130
rect 481 130 482 131
rect 480 130 481 131
rect 479 130 480 131
rect 478 130 479 131
rect 477 130 478 131
rect 476 130 477 131
rect 475 130 476 131
rect 474 130 475 131
rect 473 130 474 131
rect 472 130 473 131
rect 471 130 472 131
rect 470 130 471 131
rect 469 130 470 131
rect 468 130 469 131
rect 467 130 468 131
rect 466 130 467 131
rect 465 130 466 131
rect 464 130 465 131
rect 463 130 464 131
rect 462 130 463 131
rect 461 130 462 131
rect 460 130 461 131
rect 440 130 441 131
rect 439 130 440 131
rect 438 130 439 131
rect 437 130 438 131
rect 436 130 437 131
rect 303 130 304 131
rect 302 130 303 131
rect 301 130 302 131
rect 300 130 301 131
rect 299 130 300 131
rect 298 130 299 131
rect 297 130 298 131
rect 296 130 297 131
rect 295 130 296 131
rect 294 130 295 131
rect 293 130 294 131
rect 292 130 293 131
rect 291 130 292 131
rect 290 130 291 131
rect 289 130 290 131
rect 288 130 289 131
rect 287 130 288 131
rect 286 130 287 131
rect 285 130 286 131
rect 284 130 285 131
rect 283 130 284 131
rect 282 130 283 131
rect 281 130 282 131
rect 280 130 281 131
rect 279 130 280 131
rect 278 130 279 131
rect 277 130 278 131
rect 276 130 277 131
rect 275 130 276 131
rect 274 130 275 131
rect 273 130 274 131
rect 272 130 273 131
rect 271 130 272 131
rect 270 130 271 131
rect 269 130 270 131
rect 268 130 269 131
rect 267 130 268 131
rect 266 130 267 131
rect 265 130 266 131
rect 264 130 265 131
rect 263 130 264 131
rect 262 130 263 131
rect 261 130 262 131
rect 260 130 261 131
rect 229 130 230 131
rect 228 130 229 131
rect 227 130 228 131
rect 226 130 227 131
rect 225 130 226 131
rect 224 130 225 131
rect 223 130 224 131
rect 222 130 223 131
rect 221 130 222 131
rect 220 130 221 131
rect 219 130 220 131
rect 218 130 219 131
rect 217 130 218 131
rect 216 130 217 131
rect 215 130 216 131
rect 214 130 215 131
rect 213 130 214 131
rect 212 130 213 131
rect 211 130 212 131
rect 210 130 211 131
rect 209 130 210 131
rect 208 130 209 131
rect 207 130 208 131
rect 206 130 207 131
rect 205 130 206 131
rect 204 130 205 131
rect 203 130 204 131
rect 202 130 203 131
rect 201 130 202 131
rect 200 130 201 131
rect 199 130 200 131
rect 198 130 199 131
rect 197 130 198 131
rect 196 130 197 131
rect 195 130 196 131
rect 194 130 195 131
rect 193 130 194 131
rect 192 130 193 131
rect 191 130 192 131
rect 190 130 191 131
rect 189 130 190 131
rect 188 130 189 131
rect 187 130 188 131
rect 186 130 187 131
rect 185 130 186 131
rect 184 130 185 131
rect 183 130 184 131
rect 182 130 183 131
rect 181 130 182 131
rect 180 130 181 131
rect 179 130 180 131
rect 178 130 179 131
rect 177 130 178 131
rect 176 130 177 131
rect 175 130 176 131
rect 174 130 175 131
rect 173 130 174 131
rect 172 130 173 131
rect 171 130 172 131
rect 170 130 171 131
rect 169 130 170 131
rect 168 130 169 131
rect 167 130 168 131
rect 166 130 167 131
rect 165 130 166 131
rect 164 130 165 131
rect 147 130 148 131
rect 146 130 147 131
rect 145 130 146 131
rect 144 130 145 131
rect 143 130 144 131
rect 142 130 143 131
rect 141 130 142 131
rect 140 130 141 131
rect 139 130 140 131
rect 138 130 139 131
rect 137 130 138 131
rect 136 130 137 131
rect 135 130 136 131
rect 134 130 135 131
rect 133 130 134 131
rect 132 130 133 131
rect 131 130 132 131
rect 130 130 131 131
rect 129 130 130 131
rect 128 130 129 131
rect 127 130 128 131
rect 126 130 127 131
rect 125 130 126 131
rect 124 130 125 131
rect 123 130 124 131
rect 122 130 123 131
rect 121 130 122 131
rect 120 130 121 131
rect 119 130 120 131
rect 118 130 119 131
rect 117 130 118 131
rect 116 130 117 131
rect 115 130 116 131
rect 114 130 115 131
rect 113 130 114 131
rect 112 130 113 131
rect 111 130 112 131
rect 110 130 111 131
rect 109 130 110 131
rect 108 130 109 131
rect 107 130 108 131
rect 106 130 107 131
rect 105 130 106 131
rect 104 130 105 131
rect 103 130 104 131
rect 102 130 103 131
rect 101 130 102 131
rect 100 130 101 131
rect 99 130 100 131
rect 98 130 99 131
rect 97 130 98 131
rect 96 130 97 131
rect 95 130 96 131
rect 94 130 95 131
rect 93 130 94 131
rect 92 130 93 131
rect 91 130 92 131
rect 90 130 91 131
rect 89 130 90 131
rect 88 130 89 131
rect 87 130 88 131
rect 86 130 87 131
rect 85 130 86 131
rect 84 130 85 131
rect 83 130 84 131
rect 82 130 83 131
rect 81 130 82 131
rect 80 130 81 131
rect 79 130 80 131
rect 78 130 79 131
rect 77 130 78 131
rect 76 130 77 131
rect 75 130 76 131
rect 74 130 75 131
rect 73 130 74 131
rect 72 130 73 131
rect 71 130 72 131
rect 70 130 71 131
rect 69 130 70 131
rect 68 130 69 131
rect 67 130 68 131
rect 66 130 67 131
rect 65 130 66 131
rect 64 130 65 131
rect 63 130 64 131
rect 58 130 59 131
rect 57 130 58 131
rect 56 130 57 131
rect 55 130 56 131
rect 54 130 55 131
rect 53 130 54 131
rect 52 130 53 131
rect 51 130 52 131
rect 50 130 51 131
rect 49 130 50 131
rect 48 130 49 131
rect 47 130 48 131
rect 46 130 47 131
rect 45 130 46 131
rect 44 130 45 131
rect 43 130 44 131
rect 42 130 43 131
rect 41 130 42 131
rect 40 130 41 131
rect 39 130 40 131
rect 38 130 39 131
rect 37 130 38 131
rect 36 130 37 131
rect 35 130 36 131
rect 34 130 35 131
rect 33 130 34 131
rect 32 130 33 131
rect 31 130 32 131
rect 481 131 482 132
rect 480 131 481 132
rect 479 131 480 132
rect 478 131 479 132
rect 477 131 478 132
rect 476 131 477 132
rect 475 131 476 132
rect 474 131 475 132
rect 473 131 474 132
rect 472 131 473 132
rect 471 131 472 132
rect 470 131 471 132
rect 469 131 470 132
rect 468 131 469 132
rect 467 131 468 132
rect 466 131 467 132
rect 465 131 466 132
rect 464 131 465 132
rect 463 131 464 132
rect 462 131 463 132
rect 461 131 462 132
rect 460 131 461 132
rect 440 131 441 132
rect 439 131 440 132
rect 438 131 439 132
rect 437 131 438 132
rect 436 131 437 132
rect 304 131 305 132
rect 303 131 304 132
rect 302 131 303 132
rect 301 131 302 132
rect 300 131 301 132
rect 299 131 300 132
rect 298 131 299 132
rect 297 131 298 132
rect 296 131 297 132
rect 295 131 296 132
rect 294 131 295 132
rect 293 131 294 132
rect 292 131 293 132
rect 291 131 292 132
rect 290 131 291 132
rect 289 131 290 132
rect 288 131 289 132
rect 287 131 288 132
rect 286 131 287 132
rect 285 131 286 132
rect 284 131 285 132
rect 283 131 284 132
rect 282 131 283 132
rect 281 131 282 132
rect 280 131 281 132
rect 279 131 280 132
rect 278 131 279 132
rect 277 131 278 132
rect 276 131 277 132
rect 275 131 276 132
rect 274 131 275 132
rect 273 131 274 132
rect 272 131 273 132
rect 271 131 272 132
rect 270 131 271 132
rect 269 131 270 132
rect 268 131 269 132
rect 267 131 268 132
rect 266 131 267 132
rect 265 131 266 132
rect 264 131 265 132
rect 263 131 264 132
rect 262 131 263 132
rect 261 131 262 132
rect 260 131 261 132
rect 259 131 260 132
rect 258 131 259 132
rect 228 131 229 132
rect 227 131 228 132
rect 226 131 227 132
rect 225 131 226 132
rect 224 131 225 132
rect 223 131 224 132
rect 222 131 223 132
rect 221 131 222 132
rect 220 131 221 132
rect 219 131 220 132
rect 218 131 219 132
rect 217 131 218 132
rect 216 131 217 132
rect 215 131 216 132
rect 214 131 215 132
rect 213 131 214 132
rect 212 131 213 132
rect 211 131 212 132
rect 210 131 211 132
rect 209 131 210 132
rect 208 131 209 132
rect 207 131 208 132
rect 206 131 207 132
rect 205 131 206 132
rect 204 131 205 132
rect 203 131 204 132
rect 202 131 203 132
rect 201 131 202 132
rect 200 131 201 132
rect 199 131 200 132
rect 198 131 199 132
rect 197 131 198 132
rect 196 131 197 132
rect 195 131 196 132
rect 194 131 195 132
rect 193 131 194 132
rect 192 131 193 132
rect 191 131 192 132
rect 190 131 191 132
rect 189 131 190 132
rect 188 131 189 132
rect 187 131 188 132
rect 186 131 187 132
rect 185 131 186 132
rect 184 131 185 132
rect 183 131 184 132
rect 182 131 183 132
rect 181 131 182 132
rect 180 131 181 132
rect 179 131 180 132
rect 178 131 179 132
rect 177 131 178 132
rect 176 131 177 132
rect 175 131 176 132
rect 174 131 175 132
rect 173 131 174 132
rect 172 131 173 132
rect 171 131 172 132
rect 170 131 171 132
rect 169 131 170 132
rect 168 131 169 132
rect 167 131 168 132
rect 166 131 167 132
rect 165 131 166 132
rect 164 131 165 132
rect 146 131 147 132
rect 145 131 146 132
rect 144 131 145 132
rect 143 131 144 132
rect 142 131 143 132
rect 141 131 142 132
rect 140 131 141 132
rect 139 131 140 132
rect 138 131 139 132
rect 137 131 138 132
rect 136 131 137 132
rect 135 131 136 132
rect 134 131 135 132
rect 133 131 134 132
rect 132 131 133 132
rect 131 131 132 132
rect 130 131 131 132
rect 129 131 130 132
rect 128 131 129 132
rect 127 131 128 132
rect 126 131 127 132
rect 125 131 126 132
rect 124 131 125 132
rect 123 131 124 132
rect 122 131 123 132
rect 121 131 122 132
rect 120 131 121 132
rect 119 131 120 132
rect 118 131 119 132
rect 117 131 118 132
rect 116 131 117 132
rect 115 131 116 132
rect 114 131 115 132
rect 113 131 114 132
rect 112 131 113 132
rect 111 131 112 132
rect 110 131 111 132
rect 109 131 110 132
rect 108 131 109 132
rect 107 131 108 132
rect 106 131 107 132
rect 105 131 106 132
rect 104 131 105 132
rect 103 131 104 132
rect 102 131 103 132
rect 101 131 102 132
rect 100 131 101 132
rect 99 131 100 132
rect 98 131 99 132
rect 97 131 98 132
rect 96 131 97 132
rect 95 131 96 132
rect 94 131 95 132
rect 93 131 94 132
rect 92 131 93 132
rect 91 131 92 132
rect 90 131 91 132
rect 89 131 90 132
rect 88 131 89 132
rect 87 131 88 132
rect 86 131 87 132
rect 85 131 86 132
rect 84 131 85 132
rect 83 131 84 132
rect 82 131 83 132
rect 81 131 82 132
rect 80 131 81 132
rect 79 131 80 132
rect 78 131 79 132
rect 77 131 78 132
rect 76 131 77 132
rect 75 131 76 132
rect 74 131 75 132
rect 73 131 74 132
rect 72 131 73 132
rect 71 131 72 132
rect 70 131 71 132
rect 69 131 70 132
rect 68 131 69 132
rect 67 131 68 132
rect 66 131 67 132
rect 65 131 66 132
rect 64 131 65 132
rect 63 131 64 132
rect 62 131 63 132
rect 58 131 59 132
rect 57 131 58 132
rect 56 131 57 132
rect 55 131 56 132
rect 54 131 55 132
rect 53 131 54 132
rect 52 131 53 132
rect 51 131 52 132
rect 50 131 51 132
rect 49 131 50 132
rect 48 131 49 132
rect 47 131 48 132
rect 46 131 47 132
rect 45 131 46 132
rect 44 131 45 132
rect 43 131 44 132
rect 42 131 43 132
rect 41 131 42 132
rect 40 131 41 132
rect 39 131 40 132
rect 38 131 39 132
rect 37 131 38 132
rect 36 131 37 132
rect 35 131 36 132
rect 34 131 35 132
rect 33 131 34 132
rect 32 131 33 132
rect 31 131 32 132
rect 461 132 462 133
rect 460 132 461 133
rect 440 132 441 133
rect 439 132 440 133
rect 438 132 439 133
rect 437 132 438 133
rect 436 132 437 133
rect 435 132 436 133
rect 396 132 397 133
rect 395 132 396 133
rect 306 132 307 133
rect 305 132 306 133
rect 304 132 305 133
rect 303 132 304 133
rect 302 132 303 133
rect 301 132 302 133
rect 300 132 301 133
rect 299 132 300 133
rect 298 132 299 133
rect 297 132 298 133
rect 296 132 297 133
rect 295 132 296 133
rect 294 132 295 133
rect 293 132 294 133
rect 292 132 293 133
rect 291 132 292 133
rect 290 132 291 133
rect 289 132 290 133
rect 288 132 289 133
rect 287 132 288 133
rect 286 132 287 133
rect 285 132 286 133
rect 284 132 285 133
rect 283 132 284 133
rect 282 132 283 133
rect 281 132 282 133
rect 280 132 281 133
rect 279 132 280 133
rect 278 132 279 133
rect 277 132 278 133
rect 276 132 277 133
rect 275 132 276 133
rect 274 132 275 133
rect 273 132 274 133
rect 272 132 273 133
rect 271 132 272 133
rect 270 132 271 133
rect 269 132 270 133
rect 268 132 269 133
rect 267 132 268 133
rect 266 132 267 133
rect 265 132 266 133
rect 264 132 265 133
rect 263 132 264 133
rect 262 132 263 133
rect 261 132 262 133
rect 260 132 261 133
rect 259 132 260 133
rect 258 132 259 133
rect 257 132 258 133
rect 227 132 228 133
rect 226 132 227 133
rect 225 132 226 133
rect 224 132 225 133
rect 223 132 224 133
rect 222 132 223 133
rect 221 132 222 133
rect 220 132 221 133
rect 219 132 220 133
rect 218 132 219 133
rect 217 132 218 133
rect 216 132 217 133
rect 215 132 216 133
rect 214 132 215 133
rect 213 132 214 133
rect 212 132 213 133
rect 211 132 212 133
rect 210 132 211 133
rect 209 132 210 133
rect 208 132 209 133
rect 207 132 208 133
rect 206 132 207 133
rect 205 132 206 133
rect 204 132 205 133
rect 203 132 204 133
rect 202 132 203 133
rect 201 132 202 133
rect 200 132 201 133
rect 199 132 200 133
rect 198 132 199 133
rect 197 132 198 133
rect 196 132 197 133
rect 195 132 196 133
rect 194 132 195 133
rect 193 132 194 133
rect 192 132 193 133
rect 191 132 192 133
rect 190 132 191 133
rect 189 132 190 133
rect 188 132 189 133
rect 187 132 188 133
rect 186 132 187 133
rect 185 132 186 133
rect 184 132 185 133
rect 183 132 184 133
rect 182 132 183 133
rect 181 132 182 133
rect 180 132 181 133
rect 179 132 180 133
rect 178 132 179 133
rect 177 132 178 133
rect 176 132 177 133
rect 175 132 176 133
rect 174 132 175 133
rect 173 132 174 133
rect 172 132 173 133
rect 171 132 172 133
rect 170 132 171 133
rect 169 132 170 133
rect 168 132 169 133
rect 167 132 168 133
rect 166 132 167 133
rect 165 132 166 133
rect 164 132 165 133
rect 146 132 147 133
rect 145 132 146 133
rect 144 132 145 133
rect 143 132 144 133
rect 142 132 143 133
rect 141 132 142 133
rect 140 132 141 133
rect 139 132 140 133
rect 138 132 139 133
rect 137 132 138 133
rect 136 132 137 133
rect 135 132 136 133
rect 134 132 135 133
rect 133 132 134 133
rect 132 132 133 133
rect 131 132 132 133
rect 130 132 131 133
rect 129 132 130 133
rect 128 132 129 133
rect 127 132 128 133
rect 126 132 127 133
rect 125 132 126 133
rect 124 132 125 133
rect 123 132 124 133
rect 122 132 123 133
rect 121 132 122 133
rect 120 132 121 133
rect 119 132 120 133
rect 118 132 119 133
rect 117 132 118 133
rect 116 132 117 133
rect 115 132 116 133
rect 114 132 115 133
rect 113 132 114 133
rect 112 132 113 133
rect 111 132 112 133
rect 110 132 111 133
rect 109 132 110 133
rect 108 132 109 133
rect 107 132 108 133
rect 106 132 107 133
rect 105 132 106 133
rect 104 132 105 133
rect 103 132 104 133
rect 102 132 103 133
rect 101 132 102 133
rect 100 132 101 133
rect 99 132 100 133
rect 98 132 99 133
rect 97 132 98 133
rect 96 132 97 133
rect 95 132 96 133
rect 94 132 95 133
rect 93 132 94 133
rect 92 132 93 133
rect 91 132 92 133
rect 90 132 91 133
rect 89 132 90 133
rect 88 132 89 133
rect 87 132 88 133
rect 86 132 87 133
rect 85 132 86 133
rect 84 132 85 133
rect 83 132 84 133
rect 82 132 83 133
rect 81 132 82 133
rect 80 132 81 133
rect 79 132 80 133
rect 78 132 79 133
rect 77 132 78 133
rect 76 132 77 133
rect 75 132 76 133
rect 74 132 75 133
rect 73 132 74 133
rect 72 132 73 133
rect 71 132 72 133
rect 70 132 71 133
rect 69 132 70 133
rect 68 132 69 133
rect 67 132 68 133
rect 66 132 67 133
rect 65 132 66 133
rect 64 132 65 133
rect 63 132 64 133
rect 62 132 63 133
rect 61 132 62 133
rect 58 132 59 133
rect 57 132 58 133
rect 56 132 57 133
rect 55 132 56 133
rect 54 132 55 133
rect 53 132 54 133
rect 52 132 53 133
rect 51 132 52 133
rect 50 132 51 133
rect 49 132 50 133
rect 48 132 49 133
rect 47 132 48 133
rect 46 132 47 133
rect 45 132 46 133
rect 44 132 45 133
rect 43 132 44 133
rect 42 132 43 133
rect 41 132 42 133
rect 40 132 41 133
rect 39 132 40 133
rect 38 132 39 133
rect 37 132 38 133
rect 36 132 37 133
rect 35 132 36 133
rect 34 132 35 133
rect 33 132 34 133
rect 32 132 33 133
rect 31 132 32 133
rect 460 133 461 134
rect 439 133 440 134
rect 438 133 439 134
rect 437 133 438 134
rect 436 133 437 134
rect 435 133 436 134
rect 397 133 398 134
rect 396 133 397 134
rect 395 133 396 134
rect 307 133 308 134
rect 306 133 307 134
rect 305 133 306 134
rect 304 133 305 134
rect 303 133 304 134
rect 302 133 303 134
rect 301 133 302 134
rect 300 133 301 134
rect 299 133 300 134
rect 298 133 299 134
rect 297 133 298 134
rect 296 133 297 134
rect 295 133 296 134
rect 294 133 295 134
rect 293 133 294 134
rect 292 133 293 134
rect 291 133 292 134
rect 290 133 291 134
rect 289 133 290 134
rect 288 133 289 134
rect 287 133 288 134
rect 286 133 287 134
rect 285 133 286 134
rect 284 133 285 134
rect 283 133 284 134
rect 282 133 283 134
rect 281 133 282 134
rect 280 133 281 134
rect 279 133 280 134
rect 278 133 279 134
rect 277 133 278 134
rect 276 133 277 134
rect 275 133 276 134
rect 274 133 275 134
rect 273 133 274 134
rect 272 133 273 134
rect 271 133 272 134
rect 270 133 271 134
rect 269 133 270 134
rect 268 133 269 134
rect 267 133 268 134
rect 266 133 267 134
rect 265 133 266 134
rect 264 133 265 134
rect 263 133 264 134
rect 262 133 263 134
rect 261 133 262 134
rect 260 133 261 134
rect 259 133 260 134
rect 258 133 259 134
rect 257 133 258 134
rect 256 133 257 134
rect 255 133 256 134
rect 227 133 228 134
rect 226 133 227 134
rect 225 133 226 134
rect 224 133 225 134
rect 223 133 224 134
rect 222 133 223 134
rect 221 133 222 134
rect 220 133 221 134
rect 219 133 220 134
rect 218 133 219 134
rect 217 133 218 134
rect 216 133 217 134
rect 215 133 216 134
rect 214 133 215 134
rect 213 133 214 134
rect 212 133 213 134
rect 211 133 212 134
rect 210 133 211 134
rect 209 133 210 134
rect 208 133 209 134
rect 207 133 208 134
rect 206 133 207 134
rect 205 133 206 134
rect 204 133 205 134
rect 203 133 204 134
rect 202 133 203 134
rect 201 133 202 134
rect 200 133 201 134
rect 199 133 200 134
rect 198 133 199 134
rect 197 133 198 134
rect 196 133 197 134
rect 195 133 196 134
rect 194 133 195 134
rect 193 133 194 134
rect 192 133 193 134
rect 191 133 192 134
rect 190 133 191 134
rect 189 133 190 134
rect 188 133 189 134
rect 187 133 188 134
rect 186 133 187 134
rect 185 133 186 134
rect 184 133 185 134
rect 183 133 184 134
rect 182 133 183 134
rect 181 133 182 134
rect 180 133 181 134
rect 179 133 180 134
rect 178 133 179 134
rect 177 133 178 134
rect 176 133 177 134
rect 175 133 176 134
rect 174 133 175 134
rect 173 133 174 134
rect 172 133 173 134
rect 171 133 172 134
rect 170 133 171 134
rect 169 133 170 134
rect 168 133 169 134
rect 167 133 168 134
rect 166 133 167 134
rect 165 133 166 134
rect 164 133 165 134
rect 163 133 164 134
rect 145 133 146 134
rect 144 133 145 134
rect 143 133 144 134
rect 142 133 143 134
rect 141 133 142 134
rect 140 133 141 134
rect 139 133 140 134
rect 138 133 139 134
rect 137 133 138 134
rect 136 133 137 134
rect 135 133 136 134
rect 134 133 135 134
rect 133 133 134 134
rect 132 133 133 134
rect 131 133 132 134
rect 130 133 131 134
rect 129 133 130 134
rect 128 133 129 134
rect 127 133 128 134
rect 126 133 127 134
rect 125 133 126 134
rect 124 133 125 134
rect 123 133 124 134
rect 122 133 123 134
rect 121 133 122 134
rect 120 133 121 134
rect 119 133 120 134
rect 118 133 119 134
rect 117 133 118 134
rect 116 133 117 134
rect 115 133 116 134
rect 114 133 115 134
rect 113 133 114 134
rect 112 133 113 134
rect 111 133 112 134
rect 110 133 111 134
rect 109 133 110 134
rect 108 133 109 134
rect 107 133 108 134
rect 106 133 107 134
rect 105 133 106 134
rect 104 133 105 134
rect 103 133 104 134
rect 102 133 103 134
rect 101 133 102 134
rect 100 133 101 134
rect 99 133 100 134
rect 98 133 99 134
rect 97 133 98 134
rect 96 133 97 134
rect 95 133 96 134
rect 94 133 95 134
rect 93 133 94 134
rect 92 133 93 134
rect 91 133 92 134
rect 90 133 91 134
rect 89 133 90 134
rect 88 133 89 134
rect 87 133 88 134
rect 86 133 87 134
rect 85 133 86 134
rect 84 133 85 134
rect 83 133 84 134
rect 82 133 83 134
rect 81 133 82 134
rect 80 133 81 134
rect 79 133 80 134
rect 78 133 79 134
rect 77 133 78 134
rect 76 133 77 134
rect 75 133 76 134
rect 74 133 75 134
rect 73 133 74 134
rect 72 133 73 134
rect 71 133 72 134
rect 70 133 71 134
rect 69 133 70 134
rect 68 133 69 134
rect 67 133 68 134
rect 66 133 67 134
rect 65 133 66 134
rect 64 133 65 134
rect 63 133 64 134
rect 62 133 63 134
rect 61 133 62 134
rect 58 133 59 134
rect 57 133 58 134
rect 56 133 57 134
rect 55 133 56 134
rect 54 133 55 134
rect 53 133 54 134
rect 52 133 53 134
rect 51 133 52 134
rect 50 133 51 134
rect 49 133 50 134
rect 48 133 49 134
rect 47 133 48 134
rect 46 133 47 134
rect 45 133 46 134
rect 44 133 45 134
rect 43 133 44 134
rect 42 133 43 134
rect 41 133 42 134
rect 40 133 41 134
rect 39 133 40 134
rect 38 133 39 134
rect 37 133 38 134
rect 36 133 37 134
rect 35 133 36 134
rect 34 133 35 134
rect 33 133 34 134
rect 32 133 33 134
rect 460 134 461 135
rect 439 134 440 135
rect 438 134 439 135
rect 437 134 438 135
rect 436 134 437 135
rect 435 134 436 135
rect 434 134 435 135
rect 397 134 398 135
rect 396 134 397 135
rect 395 134 396 135
rect 308 134 309 135
rect 307 134 308 135
rect 306 134 307 135
rect 305 134 306 135
rect 304 134 305 135
rect 303 134 304 135
rect 302 134 303 135
rect 301 134 302 135
rect 300 134 301 135
rect 299 134 300 135
rect 298 134 299 135
rect 297 134 298 135
rect 296 134 297 135
rect 295 134 296 135
rect 294 134 295 135
rect 293 134 294 135
rect 292 134 293 135
rect 291 134 292 135
rect 290 134 291 135
rect 289 134 290 135
rect 288 134 289 135
rect 287 134 288 135
rect 286 134 287 135
rect 285 134 286 135
rect 284 134 285 135
rect 283 134 284 135
rect 282 134 283 135
rect 281 134 282 135
rect 280 134 281 135
rect 279 134 280 135
rect 278 134 279 135
rect 277 134 278 135
rect 276 134 277 135
rect 275 134 276 135
rect 274 134 275 135
rect 273 134 274 135
rect 272 134 273 135
rect 271 134 272 135
rect 270 134 271 135
rect 269 134 270 135
rect 268 134 269 135
rect 267 134 268 135
rect 266 134 267 135
rect 265 134 266 135
rect 264 134 265 135
rect 263 134 264 135
rect 262 134 263 135
rect 261 134 262 135
rect 260 134 261 135
rect 259 134 260 135
rect 258 134 259 135
rect 257 134 258 135
rect 256 134 257 135
rect 255 134 256 135
rect 254 134 255 135
rect 226 134 227 135
rect 225 134 226 135
rect 224 134 225 135
rect 223 134 224 135
rect 222 134 223 135
rect 221 134 222 135
rect 220 134 221 135
rect 219 134 220 135
rect 218 134 219 135
rect 217 134 218 135
rect 216 134 217 135
rect 215 134 216 135
rect 214 134 215 135
rect 213 134 214 135
rect 212 134 213 135
rect 211 134 212 135
rect 210 134 211 135
rect 209 134 210 135
rect 208 134 209 135
rect 207 134 208 135
rect 206 134 207 135
rect 205 134 206 135
rect 204 134 205 135
rect 203 134 204 135
rect 202 134 203 135
rect 201 134 202 135
rect 200 134 201 135
rect 199 134 200 135
rect 198 134 199 135
rect 197 134 198 135
rect 196 134 197 135
rect 195 134 196 135
rect 194 134 195 135
rect 193 134 194 135
rect 192 134 193 135
rect 191 134 192 135
rect 190 134 191 135
rect 189 134 190 135
rect 188 134 189 135
rect 187 134 188 135
rect 186 134 187 135
rect 185 134 186 135
rect 184 134 185 135
rect 183 134 184 135
rect 182 134 183 135
rect 181 134 182 135
rect 180 134 181 135
rect 179 134 180 135
rect 178 134 179 135
rect 177 134 178 135
rect 176 134 177 135
rect 175 134 176 135
rect 174 134 175 135
rect 173 134 174 135
rect 172 134 173 135
rect 171 134 172 135
rect 170 134 171 135
rect 169 134 170 135
rect 168 134 169 135
rect 167 134 168 135
rect 166 134 167 135
rect 165 134 166 135
rect 164 134 165 135
rect 163 134 164 135
rect 145 134 146 135
rect 144 134 145 135
rect 143 134 144 135
rect 142 134 143 135
rect 141 134 142 135
rect 140 134 141 135
rect 139 134 140 135
rect 138 134 139 135
rect 137 134 138 135
rect 136 134 137 135
rect 135 134 136 135
rect 134 134 135 135
rect 133 134 134 135
rect 132 134 133 135
rect 131 134 132 135
rect 130 134 131 135
rect 129 134 130 135
rect 128 134 129 135
rect 127 134 128 135
rect 126 134 127 135
rect 125 134 126 135
rect 124 134 125 135
rect 123 134 124 135
rect 122 134 123 135
rect 121 134 122 135
rect 120 134 121 135
rect 119 134 120 135
rect 118 134 119 135
rect 117 134 118 135
rect 116 134 117 135
rect 115 134 116 135
rect 114 134 115 135
rect 113 134 114 135
rect 112 134 113 135
rect 111 134 112 135
rect 110 134 111 135
rect 109 134 110 135
rect 108 134 109 135
rect 107 134 108 135
rect 106 134 107 135
rect 105 134 106 135
rect 104 134 105 135
rect 103 134 104 135
rect 102 134 103 135
rect 101 134 102 135
rect 100 134 101 135
rect 99 134 100 135
rect 98 134 99 135
rect 97 134 98 135
rect 96 134 97 135
rect 95 134 96 135
rect 94 134 95 135
rect 93 134 94 135
rect 92 134 93 135
rect 91 134 92 135
rect 90 134 91 135
rect 89 134 90 135
rect 88 134 89 135
rect 87 134 88 135
rect 86 134 87 135
rect 85 134 86 135
rect 84 134 85 135
rect 83 134 84 135
rect 82 134 83 135
rect 81 134 82 135
rect 80 134 81 135
rect 79 134 80 135
rect 78 134 79 135
rect 77 134 78 135
rect 76 134 77 135
rect 75 134 76 135
rect 74 134 75 135
rect 73 134 74 135
rect 72 134 73 135
rect 71 134 72 135
rect 70 134 71 135
rect 69 134 70 135
rect 68 134 69 135
rect 67 134 68 135
rect 66 134 67 135
rect 65 134 66 135
rect 64 134 65 135
rect 63 134 64 135
rect 62 134 63 135
rect 61 134 62 135
rect 60 134 61 135
rect 58 134 59 135
rect 57 134 58 135
rect 56 134 57 135
rect 55 134 56 135
rect 54 134 55 135
rect 53 134 54 135
rect 52 134 53 135
rect 51 134 52 135
rect 50 134 51 135
rect 49 134 50 135
rect 48 134 49 135
rect 47 134 48 135
rect 46 134 47 135
rect 45 134 46 135
rect 44 134 45 135
rect 43 134 44 135
rect 42 134 43 135
rect 41 134 42 135
rect 40 134 41 135
rect 39 134 40 135
rect 38 134 39 135
rect 37 134 38 135
rect 36 134 37 135
rect 35 134 36 135
rect 34 134 35 135
rect 33 134 34 135
rect 439 135 440 136
rect 438 135 439 136
rect 437 135 438 136
rect 436 135 437 136
rect 435 135 436 136
rect 434 135 435 136
rect 433 135 434 136
rect 397 135 398 136
rect 396 135 397 136
rect 395 135 396 136
rect 309 135 310 136
rect 308 135 309 136
rect 307 135 308 136
rect 306 135 307 136
rect 305 135 306 136
rect 304 135 305 136
rect 303 135 304 136
rect 302 135 303 136
rect 301 135 302 136
rect 300 135 301 136
rect 299 135 300 136
rect 298 135 299 136
rect 297 135 298 136
rect 296 135 297 136
rect 295 135 296 136
rect 294 135 295 136
rect 293 135 294 136
rect 292 135 293 136
rect 291 135 292 136
rect 290 135 291 136
rect 289 135 290 136
rect 288 135 289 136
rect 287 135 288 136
rect 286 135 287 136
rect 285 135 286 136
rect 284 135 285 136
rect 283 135 284 136
rect 282 135 283 136
rect 281 135 282 136
rect 280 135 281 136
rect 279 135 280 136
rect 278 135 279 136
rect 277 135 278 136
rect 276 135 277 136
rect 275 135 276 136
rect 274 135 275 136
rect 273 135 274 136
rect 272 135 273 136
rect 271 135 272 136
rect 270 135 271 136
rect 269 135 270 136
rect 268 135 269 136
rect 267 135 268 136
rect 266 135 267 136
rect 265 135 266 136
rect 264 135 265 136
rect 263 135 264 136
rect 262 135 263 136
rect 261 135 262 136
rect 260 135 261 136
rect 259 135 260 136
rect 258 135 259 136
rect 257 135 258 136
rect 256 135 257 136
rect 255 135 256 136
rect 254 135 255 136
rect 253 135 254 136
rect 225 135 226 136
rect 224 135 225 136
rect 223 135 224 136
rect 222 135 223 136
rect 221 135 222 136
rect 220 135 221 136
rect 219 135 220 136
rect 218 135 219 136
rect 217 135 218 136
rect 216 135 217 136
rect 215 135 216 136
rect 214 135 215 136
rect 213 135 214 136
rect 212 135 213 136
rect 211 135 212 136
rect 210 135 211 136
rect 209 135 210 136
rect 208 135 209 136
rect 207 135 208 136
rect 206 135 207 136
rect 205 135 206 136
rect 204 135 205 136
rect 203 135 204 136
rect 202 135 203 136
rect 201 135 202 136
rect 200 135 201 136
rect 199 135 200 136
rect 198 135 199 136
rect 197 135 198 136
rect 196 135 197 136
rect 195 135 196 136
rect 194 135 195 136
rect 193 135 194 136
rect 192 135 193 136
rect 191 135 192 136
rect 190 135 191 136
rect 189 135 190 136
rect 188 135 189 136
rect 187 135 188 136
rect 186 135 187 136
rect 185 135 186 136
rect 184 135 185 136
rect 183 135 184 136
rect 182 135 183 136
rect 181 135 182 136
rect 180 135 181 136
rect 179 135 180 136
rect 178 135 179 136
rect 177 135 178 136
rect 176 135 177 136
rect 175 135 176 136
rect 174 135 175 136
rect 173 135 174 136
rect 172 135 173 136
rect 171 135 172 136
rect 170 135 171 136
rect 169 135 170 136
rect 168 135 169 136
rect 167 135 168 136
rect 166 135 167 136
rect 165 135 166 136
rect 164 135 165 136
rect 163 135 164 136
rect 162 135 163 136
rect 144 135 145 136
rect 143 135 144 136
rect 142 135 143 136
rect 141 135 142 136
rect 140 135 141 136
rect 139 135 140 136
rect 138 135 139 136
rect 137 135 138 136
rect 136 135 137 136
rect 135 135 136 136
rect 134 135 135 136
rect 133 135 134 136
rect 132 135 133 136
rect 131 135 132 136
rect 130 135 131 136
rect 129 135 130 136
rect 128 135 129 136
rect 127 135 128 136
rect 126 135 127 136
rect 125 135 126 136
rect 124 135 125 136
rect 123 135 124 136
rect 122 135 123 136
rect 121 135 122 136
rect 120 135 121 136
rect 119 135 120 136
rect 118 135 119 136
rect 117 135 118 136
rect 116 135 117 136
rect 115 135 116 136
rect 114 135 115 136
rect 113 135 114 136
rect 112 135 113 136
rect 111 135 112 136
rect 110 135 111 136
rect 109 135 110 136
rect 108 135 109 136
rect 107 135 108 136
rect 106 135 107 136
rect 105 135 106 136
rect 104 135 105 136
rect 103 135 104 136
rect 102 135 103 136
rect 101 135 102 136
rect 100 135 101 136
rect 99 135 100 136
rect 98 135 99 136
rect 97 135 98 136
rect 96 135 97 136
rect 95 135 96 136
rect 94 135 95 136
rect 93 135 94 136
rect 92 135 93 136
rect 91 135 92 136
rect 90 135 91 136
rect 89 135 90 136
rect 88 135 89 136
rect 87 135 88 136
rect 86 135 87 136
rect 85 135 86 136
rect 84 135 85 136
rect 83 135 84 136
rect 82 135 83 136
rect 81 135 82 136
rect 80 135 81 136
rect 79 135 80 136
rect 78 135 79 136
rect 77 135 78 136
rect 76 135 77 136
rect 75 135 76 136
rect 74 135 75 136
rect 73 135 74 136
rect 72 135 73 136
rect 71 135 72 136
rect 70 135 71 136
rect 69 135 70 136
rect 68 135 69 136
rect 67 135 68 136
rect 66 135 67 136
rect 65 135 66 136
rect 64 135 65 136
rect 63 135 64 136
rect 62 135 63 136
rect 61 135 62 136
rect 60 135 61 136
rect 59 135 60 136
rect 58 135 59 136
rect 57 135 58 136
rect 56 135 57 136
rect 55 135 56 136
rect 54 135 55 136
rect 53 135 54 136
rect 52 135 53 136
rect 51 135 52 136
rect 50 135 51 136
rect 49 135 50 136
rect 48 135 49 136
rect 47 135 48 136
rect 46 135 47 136
rect 45 135 46 136
rect 44 135 45 136
rect 43 135 44 136
rect 42 135 43 136
rect 41 135 42 136
rect 40 135 41 136
rect 39 135 40 136
rect 38 135 39 136
rect 37 135 38 136
rect 36 135 37 136
rect 35 135 36 136
rect 34 135 35 136
rect 33 135 34 136
rect 438 136 439 137
rect 437 136 438 137
rect 436 136 437 137
rect 435 136 436 137
rect 434 136 435 137
rect 433 136 434 137
rect 432 136 433 137
rect 398 136 399 137
rect 397 136 398 137
rect 396 136 397 137
rect 395 136 396 137
rect 310 136 311 137
rect 309 136 310 137
rect 308 136 309 137
rect 307 136 308 137
rect 306 136 307 137
rect 305 136 306 137
rect 304 136 305 137
rect 303 136 304 137
rect 302 136 303 137
rect 301 136 302 137
rect 300 136 301 137
rect 299 136 300 137
rect 298 136 299 137
rect 297 136 298 137
rect 296 136 297 137
rect 295 136 296 137
rect 294 136 295 137
rect 293 136 294 137
rect 292 136 293 137
rect 291 136 292 137
rect 290 136 291 137
rect 289 136 290 137
rect 288 136 289 137
rect 287 136 288 137
rect 286 136 287 137
rect 285 136 286 137
rect 284 136 285 137
rect 283 136 284 137
rect 282 136 283 137
rect 281 136 282 137
rect 280 136 281 137
rect 279 136 280 137
rect 278 136 279 137
rect 277 136 278 137
rect 276 136 277 137
rect 275 136 276 137
rect 274 136 275 137
rect 273 136 274 137
rect 272 136 273 137
rect 271 136 272 137
rect 270 136 271 137
rect 269 136 270 137
rect 268 136 269 137
rect 267 136 268 137
rect 266 136 267 137
rect 265 136 266 137
rect 264 136 265 137
rect 263 136 264 137
rect 262 136 263 137
rect 261 136 262 137
rect 260 136 261 137
rect 259 136 260 137
rect 258 136 259 137
rect 257 136 258 137
rect 256 136 257 137
rect 255 136 256 137
rect 254 136 255 137
rect 253 136 254 137
rect 252 136 253 137
rect 251 136 252 137
rect 225 136 226 137
rect 224 136 225 137
rect 223 136 224 137
rect 222 136 223 137
rect 221 136 222 137
rect 220 136 221 137
rect 219 136 220 137
rect 218 136 219 137
rect 217 136 218 137
rect 216 136 217 137
rect 215 136 216 137
rect 214 136 215 137
rect 213 136 214 137
rect 212 136 213 137
rect 211 136 212 137
rect 210 136 211 137
rect 209 136 210 137
rect 208 136 209 137
rect 207 136 208 137
rect 206 136 207 137
rect 205 136 206 137
rect 204 136 205 137
rect 203 136 204 137
rect 202 136 203 137
rect 201 136 202 137
rect 200 136 201 137
rect 199 136 200 137
rect 198 136 199 137
rect 197 136 198 137
rect 196 136 197 137
rect 195 136 196 137
rect 194 136 195 137
rect 193 136 194 137
rect 192 136 193 137
rect 191 136 192 137
rect 190 136 191 137
rect 189 136 190 137
rect 188 136 189 137
rect 187 136 188 137
rect 186 136 187 137
rect 185 136 186 137
rect 184 136 185 137
rect 183 136 184 137
rect 182 136 183 137
rect 181 136 182 137
rect 180 136 181 137
rect 179 136 180 137
rect 178 136 179 137
rect 177 136 178 137
rect 176 136 177 137
rect 175 136 176 137
rect 174 136 175 137
rect 173 136 174 137
rect 172 136 173 137
rect 171 136 172 137
rect 170 136 171 137
rect 169 136 170 137
rect 168 136 169 137
rect 167 136 168 137
rect 166 136 167 137
rect 165 136 166 137
rect 164 136 165 137
rect 163 136 164 137
rect 162 136 163 137
rect 143 136 144 137
rect 142 136 143 137
rect 141 136 142 137
rect 140 136 141 137
rect 139 136 140 137
rect 138 136 139 137
rect 137 136 138 137
rect 136 136 137 137
rect 135 136 136 137
rect 134 136 135 137
rect 133 136 134 137
rect 132 136 133 137
rect 131 136 132 137
rect 130 136 131 137
rect 129 136 130 137
rect 128 136 129 137
rect 127 136 128 137
rect 126 136 127 137
rect 125 136 126 137
rect 124 136 125 137
rect 123 136 124 137
rect 122 136 123 137
rect 121 136 122 137
rect 120 136 121 137
rect 119 136 120 137
rect 118 136 119 137
rect 117 136 118 137
rect 116 136 117 137
rect 115 136 116 137
rect 114 136 115 137
rect 113 136 114 137
rect 112 136 113 137
rect 111 136 112 137
rect 110 136 111 137
rect 109 136 110 137
rect 108 136 109 137
rect 107 136 108 137
rect 106 136 107 137
rect 105 136 106 137
rect 104 136 105 137
rect 103 136 104 137
rect 102 136 103 137
rect 101 136 102 137
rect 100 136 101 137
rect 99 136 100 137
rect 98 136 99 137
rect 97 136 98 137
rect 96 136 97 137
rect 95 136 96 137
rect 94 136 95 137
rect 93 136 94 137
rect 92 136 93 137
rect 91 136 92 137
rect 90 136 91 137
rect 89 136 90 137
rect 88 136 89 137
rect 87 136 88 137
rect 86 136 87 137
rect 85 136 86 137
rect 84 136 85 137
rect 83 136 84 137
rect 82 136 83 137
rect 81 136 82 137
rect 80 136 81 137
rect 79 136 80 137
rect 78 136 79 137
rect 77 136 78 137
rect 76 136 77 137
rect 75 136 76 137
rect 74 136 75 137
rect 73 136 74 137
rect 72 136 73 137
rect 71 136 72 137
rect 70 136 71 137
rect 69 136 70 137
rect 68 136 69 137
rect 67 136 68 137
rect 66 136 67 137
rect 65 136 66 137
rect 64 136 65 137
rect 63 136 64 137
rect 62 136 63 137
rect 61 136 62 137
rect 60 136 61 137
rect 59 136 60 137
rect 58 136 59 137
rect 57 136 58 137
rect 56 136 57 137
rect 55 136 56 137
rect 54 136 55 137
rect 53 136 54 137
rect 52 136 53 137
rect 51 136 52 137
rect 50 136 51 137
rect 49 136 50 137
rect 48 136 49 137
rect 47 136 48 137
rect 46 136 47 137
rect 45 136 46 137
rect 44 136 45 137
rect 43 136 44 137
rect 42 136 43 137
rect 41 136 42 137
rect 40 136 41 137
rect 39 136 40 137
rect 38 136 39 137
rect 37 136 38 137
rect 36 136 37 137
rect 35 136 36 137
rect 34 136 35 137
rect 438 137 439 138
rect 437 137 438 138
rect 436 137 437 138
rect 435 137 436 138
rect 434 137 435 138
rect 433 137 434 138
rect 432 137 433 138
rect 431 137 432 138
rect 430 137 431 138
rect 429 137 430 138
rect 399 137 400 138
rect 398 137 399 138
rect 397 137 398 138
rect 396 137 397 138
rect 395 137 396 138
rect 310 137 311 138
rect 309 137 310 138
rect 308 137 309 138
rect 307 137 308 138
rect 306 137 307 138
rect 305 137 306 138
rect 304 137 305 138
rect 303 137 304 138
rect 302 137 303 138
rect 301 137 302 138
rect 300 137 301 138
rect 299 137 300 138
rect 298 137 299 138
rect 297 137 298 138
rect 296 137 297 138
rect 295 137 296 138
rect 294 137 295 138
rect 293 137 294 138
rect 292 137 293 138
rect 291 137 292 138
rect 290 137 291 138
rect 289 137 290 138
rect 288 137 289 138
rect 287 137 288 138
rect 286 137 287 138
rect 285 137 286 138
rect 284 137 285 138
rect 283 137 284 138
rect 282 137 283 138
rect 281 137 282 138
rect 280 137 281 138
rect 279 137 280 138
rect 278 137 279 138
rect 277 137 278 138
rect 276 137 277 138
rect 275 137 276 138
rect 274 137 275 138
rect 273 137 274 138
rect 272 137 273 138
rect 271 137 272 138
rect 270 137 271 138
rect 269 137 270 138
rect 268 137 269 138
rect 267 137 268 138
rect 266 137 267 138
rect 265 137 266 138
rect 264 137 265 138
rect 263 137 264 138
rect 262 137 263 138
rect 261 137 262 138
rect 260 137 261 138
rect 259 137 260 138
rect 258 137 259 138
rect 257 137 258 138
rect 256 137 257 138
rect 255 137 256 138
rect 254 137 255 138
rect 253 137 254 138
rect 252 137 253 138
rect 251 137 252 138
rect 250 137 251 138
rect 224 137 225 138
rect 223 137 224 138
rect 222 137 223 138
rect 221 137 222 138
rect 220 137 221 138
rect 219 137 220 138
rect 218 137 219 138
rect 217 137 218 138
rect 216 137 217 138
rect 215 137 216 138
rect 214 137 215 138
rect 213 137 214 138
rect 212 137 213 138
rect 211 137 212 138
rect 210 137 211 138
rect 209 137 210 138
rect 208 137 209 138
rect 207 137 208 138
rect 206 137 207 138
rect 205 137 206 138
rect 204 137 205 138
rect 203 137 204 138
rect 202 137 203 138
rect 201 137 202 138
rect 200 137 201 138
rect 199 137 200 138
rect 198 137 199 138
rect 197 137 198 138
rect 196 137 197 138
rect 195 137 196 138
rect 194 137 195 138
rect 193 137 194 138
rect 192 137 193 138
rect 191 137 192 138
rect 190 137 191 138
rect 189 137 190 138
rect 188 137 189 138
rect 187 137 188 138
rect 186 137 187 138
rect 185 137 186 138
rect 184 137 185 138
rect 183 137 184 138
rect 182 137 183 138
rect 181 137 182 138
rect 180 137 181 138
rect 179 137 180 138
rect 178 137 179 138
rect 177 137 178 138
rect 176 137 177 138
rect 175 137 176 138
rect 174 137 175 138
rect 173 137 174 138
rect 172 137 173 138
rect 171 137 172 138
rect 170 137 171 138
rect 169 137 170 138
rect 168 137 169 138
rect 167 137 168 138
rect 166 137 167 138
rect 165 137 166 138
rect 164 137 165 138
rect 163 137 164 138
rect 162 137 163 138
rect 161 137 162 138
rect 143 137 144 138
rect 142 137 143 138
rect 141 137 142 138
rect 140 137 141 138
rect 139 137 140 138
rect 138 137 139 138
rect 137 137 138 138
rect 136 137 137 138
rect 135 137 136 138
rect 134 137 135 138
rect 133 137 134 138
rect 132 137 133 138
rect 131 137 132 138
rect 130 137 131 138
rect 129 137 130 138
rect 128 137 129 138
rect 127 137 128 138
rect 126 137 127 138
rect 125 137 126 138
rect 124 137 125 138
rect 123 137 124 138
rect 122 137 123 138
rect 121 137 122 138
rect 120 137 121 138
rect 119 137 120 138
rect 118 137 119 138
rect 117 137 118 138
rect 116 137 117 138
rect 115 137 116 138
rect 114 137 115 138
rect 113 137 114 138
rect 112 137 113 138
rect 111 137 112 138
rect 110 137 111 138
rect 109 137 110 138
rect 108 137 109 138
rect 107 137 108 138
rect 106 137 107 138
rect 105 137 106 138
rect 104 137 105 138
rect 103 137 104 138
rect 102 137 103 138
rect 101 137 102 138
rect 100 137 101 138
rect 99 137 100 138
rect 98 137 99 138
rect 97 137 98 138
rect 96 137 97 138
rect 95 137 96 138
rect 94 137 95 138
rect 93 137 94 138
rect 92 137 93 138
rect 91 137 92 138
rect 90 137 91 138
rect 89 137 90 138
rect 88 137 89 138
rect 87 137 88 138
rect 86 137 87 138
rect 85 137 86 138
rect 84 137 85 138
rect 83 137 84 138
rect 82 137 83 138
rect 81 137 82 138
rect 80 137 81 138
rect 79 137 80 138
rect 78 137 79 138
rect 77 137 78 138
rect 76 137 77 138
rect 75 137 76 138
rect 74 137 75 138
rect 73 137 74 138
rect 72 137 73 138
rect 71 137 72 138
rect 70 137 71 138
rect 69 137 70 138
rect 68 137 69 138
rect 67 137 68 138
rect 66 137 67 138
rect 65 137 66 138
rect 64 137 65 138
rect 63 137 64 138
rect 62 137 63 138
rect 61 137 62 138
rect 60 137 61 138
rect 59 137 60 138
rect 58 137 59 138
rect 57 137 58 138
rect 56 137 57 138
rect 55 137 56 138
rect 54 137 55 138
rect 53 137 54 138
rect 52 137 53 138
rect 51 137 52 138
rect 50 137 51 138
rect 49 137 50 138
rect 48 137 49 138
rect 47 137 48 138
rect 46 137 47 138
rect 45 137 46 138
rect 44 137 45 138
rect 43 137 44 138
rect 42 137 43 138
rect 41 137 42 138
rect 40 137 41 138
rect 39 137 40 138
rect 38 137 39 138
rect 37 137 38 138
rect 36 137 37 138
rect 35 137 36 138
rect 437 138 438 139
rect 436 138 437 139
rect 435 138 436 139
rect 434 138 435 139
rect 433 138 434 139
rect 432 138 433 139
rect 431 138 432 139
rect 430 138 431 139
rect 429 138 430 139
rect 428 138 429 139
rect 427 138 428 139
rect 426 138 427 139
rect 425 138 426 139
rect 424 138 425 139
rect 405 138 406 139
rect 404 138 405 139
rect 403 138 404 139
rect 402 138 403 139
rect 401 138 402 139
rect 400 138 401 139
rect 399 138 400 139
rect 398 138 399 139
rect 397 138 398 139
rect 396 138 397 139
rect 395 138 396 139
rect 311 138 312 139
rect 310 138 311 139
rect 309 138 310 139
rect 308 138 309 139
rect 307 138 308 139
rect 306 138 307 139
rect 305 138 306 139
rect 304 138 305 139
rect 303 138 304 139
rect 302 138 303 139
rect 301 138 302 139
rect 300 138 301 139
rect 299 138 300 139
rect 298 138 299 139
rect 297 138 298 139
rect 296 138 297 139
rect 295 138 296 139
rect 294 138 295 139
rect 293 138 294 139
rect 292 138 293 139
rect 291 138 292 139
rect 290 138 291 139
rect 289 138 290 139
rect 288 138 289 139
rect 287 138 288 139
rect 286 138 287 139
rect 285 138 286 139
rect 284 138 285 139
rect 283 138 284 139
rect 282 138 283 139
rect 281 138 282 139
rect 280 138 281 139
rect 279 138 280 139
rect 278 138 279 139
rect 277 138 278 139
rect 276 138 277 139
rect 275 138 276 139
rect 274 138 275 139
rect 273 138 274 139
rect 272 138 273 139
rect 271 138 272 139
rect 270 138 271 139
rect 269 138 270 139
rect 268 138 269 139
rect 267 138 268 139
rect 266 138 267 139
rect 265 138 266 139
rect 264 138 265 139
rect 263 138 264 139
rect 262 138 263 139
rect 261 138 262 139
rect 260 138 261 139
rect 259 138 260 139
rect 258 138 259 139
rect 257 138 258 139
rect 256 138 257 139
rect 255 138 256 139
rect 254 138 255 139
rect 253 138 254 139
rect 252 138 253 139
rect 251 138 252 139
rect 250 138 251 139
rect 249 138 250 139
rect 224 138 225 139
rect 223 138 224 139
rect 222 138 223 139
rect 221 138 222 139
rect 220 138 221 139
rect 219 138 220 139
rect 218 138 219 139
rect 217 138 218 139
rect 216 138 217 139
rect 215 138 216 139
rect 214 138 215 139
rect 213 138 214 139
rect 212 138 213 139
rect 211 138 212 139
rect 210 138 211 139
rect 209 138 210 139
rect 208 138 209 139
rect 207 138 208 139
rect 206 138 207 139
rect 205 138 206 139
rect 204 138 205 139
rect 203 138 204 139
rect 202 138 203 139
rect 201 138 202 139
rect 200 138 201 139
rect 199 138 200 139
rect 198 138 199 139
rect 197 138 198 139
rect 196 138 197 139
rect 195 138 196 139
rect 194 138 195 139
rect 193 138 194 139
rect 192 138 193 139
rect 191 138 192 139
rect 190 138 191 139
rect 189 138 190 139
rect 188 138 189 139
rect 187 138 188 139
rect 186 138 187 139
rect 185 138 186 139
rect 184 138 185 139
rect 183 138 184 139
rect 182 138 183 139
rect 181 138 182 139
rect 180 138 181 139
rect 179 138 180 139
rect 178 138 179 139
rect 177 138 178 139
rect 176 138 177 139
rect 175 138 176 139
rect 174 138 175 139
rect 173 138 174 139
rect 172 138 173 139
rect 171 138 172 139
rect 170 138 171 139
rect 169 138 170 139
rect 168 138 169 139
rect 167 138 168 139
rect 166 138 167 139
rect 165 138 166 139
rect 164 138 165 139
rect 163 138 164 139
rect 162 138 163 139
rect 161 138 162 139
rect 142 138 143 139
rect 141 138 142 139
rect 140 138 141 139
rect 139 138 140 139
rect 138 138 139 139
rect 137 138 138 139
rect 136 138 137 139
rect 135 138 136 139
rect 134 138 135 139
rect 133 138 134 139
rect 132 138 133 139
rect 131 138 132 139
rect 130 138 131 139
rect 129 138 130 139
rect 128 138 129 139
rect 127 138 128 139
rect 126 138 127 139
rect 125 138 126 139
rect 124 138 125 139
rect 123 138 124 139
rect 122 138 123 139
rect 121 138 122 139
rect 120 138 121 139
rect 119 138 120 139
rect 118 138 119 139
rect 117 138 118 139
rect 116 138 117 139
rect 115 138 116 139
rect 114 138 115 139
rect 113 138 114 139
rect 112 138 113 139
rect 111 138 112 139
rect 110 138 111 139
rect 109 138 110 139
rect 108 138 109 139
rect 107 138 108 139
rect 106 138 107 139
rect 105 138 106 139
rect 104 138 105 139
rect 103 138 104 139
rect 102 138 103 139
rect 101 138 102 139
rect 100 138 101 139
rect 99 138 100 139
rect 98 138 99 139
rect 97 138 98 139
rect 96 138 97 139
rect 95 138 96 139
rect 94 138 95 139
rect 93 138 94 139
rect 92 138 93 139
rect 91 138 92 139
rect 90 138 91 139
rect 89 138 90 139
rect 88 138 89 139
rect 87 138 88 139
rect 86 138 87 139
rect 85 138 86 139
rect 84 138 85 139
rect 83 138 84 139
rect 82 138 83 139
rect 81 138 82 139
rect 80 138 81 139
rect 79 138 80 139
rect 78 138 79 139
rect 77 138 78 139
rect 76 138 77 139
rect 75 138 76 139
rect 74 138 75 139
rect 73 138 74 139
rect 72 138 73 139
rect 71 138 72 139
rect 70 138 71 139
rect 69 138 70 139
rect 68 138 69 139
rect 67 138 68 139
rect 66 138 67 139
rect 65 138 66 139
rect 64 138 65 139
rect 63 138 64 139
rect 62 138 63 139
rect 61 138 62 139
rect 60 138 61 139
rect 59 138 60 139
rect 58 138 59 139
rect 57 138 58 139
rect 56 138 57 139
rect 55 138 56 139
rect 54 138 55 139
rect 53 138 54 139
rect 52 138 53 139
rect 51 138 52 139
rect 50 138 51 139
rect 49 138 50 139
rect 48 138 49 139
rect 47 138 48 139
rect 46 138 47 139
rect 45 138 46 139
rect 44 138 45 139
rect 43 138 44 139
rect 42 138 43 139
rect 41 138 42 139
rect 40 138 41 139
rect 39 138 40 139
rect 38 138 39 139
rect 37 138 38 139
rect 36 138 37 139
rect 436 139 437 140
rect 435 139 436 140
rect 434 139 435 140
rect 433 139 434 140
rect 432 139 433 140
rect 431 139 432 140
rect 430 139 431 140
rect 429 139 430 140
rect 428 139 429 140
rect 427 139 428 140
rect 426 139 427 140
rect 425 139 426 140
rect 424 139 425 140
rect 423 139 424 140
rect 422 139 423 140
rect 421 139 422 140
rect 420 139 421 140
rect 419 139 420 140
rect 418 139 419 140
rect 417 139 418 140
rect 416 139 417 140
rect 415 139 416 140
rect 414 139 415 140
rect 413 139 414 140
rect 412 139 413 140
rect 411 139 412 140
rect 410 139 411 140
rect 409 139 410 140
rect 408 139 409 140
rect 407 139 408 140
rect 406 139 407 140
rect 405 139 406 140
rect 404 139 405 140
rect 403 139 404 140
rect 402 139 403 140
rect 401 139 402 140
rect 400 139 401 140
rect 399 139 400 140
rect 398 139 399 140
rect 397 139 398 140
rect 396 139 397 140
rect 395 139 396 140
rect 312 139 313 140
rect 311 139 312 140
rect 310 139 311 140
rect 309 139 310 140
rect 308 139 309 140
rect 307 139 308 140
rect 306 139 307 140
rect 305 139 306 140
rect 304 139 305 140
rect 303 139 304 140
rect 302 139 303 140
rect 301 139 302 140
rect 300 139 301 140
rect 299 139 300 140
rect 298 139 299 140
rect 297 139 298 140
rect 296 139 297 140
rect 295 139 296 140
rect 294 139 295 140
rect 293 139 294 140
rect 292 139 293 140
rect 291 139 292 140
rect 290 139 291 140
rect 289 139 290 140
rect 288 139 289 140
rect 287 139 288 140
rect 286 139 287 140
rect 285 139 286 140
rect 284 139 285 140
rect 283 139 284 140
rect 282 139 283 140
rect 281 139 282 140
rect 280 139 281 140
rect 279 139 280 140
rect 278 139 279 140
rect 277 139 278 140
rect 276 139 277 140
rect 275 139 276 140
rect 274 139 275 140
rect 273 139 274 140
rect 272 139 273 140
rect 271 139 272 140
rect 270 139 271 140
rect 269 139 270 140
rect 268 139 269 140
rect 267 139 268 140
rect 266 139 267 140
rect 265 139 266 140
rect 264 139 265 140
rect 263 139 264 140
rect 262 139 263 140
rect 261 139 262 140
rect 260 139 261 140
rect 259 139 260 140
rect 258 139 259 140
rect 257 139 258 140
rect 256 139 257 140
rect 255 139 256 140
rect 254 139 255 140
rect 253 139 254 140
rect 252 139 253 140
rect 251 139 252 140
rect 250 139 251 140
rect 249 139 250 140
rect 248 139 249 140
rect 223 139 224 140
rect 222 139 223 140
rect 221 139 222 140
rect 220 139 221 140
rect 219 139 220 140
rect 218 139 219 140
rect 217 139 218 140
rect 216 139 217 140
rect 215 139 216 140
rect 214 139 215 140
rect 213 139 214 140
rect 212 139 213 140
rect 211 139 212 140
rect 210 139 211 140
rect 209 139 210 140
rect 208 139 209 140
rect 207 139 208 140
rect 206 139 207 140
rect 205 139 206 140
rect 204 139 205 140
rect 203 139 204 140
rect 202 139 203 140
rect 201 139 202 140
rect 200 139 201 140
rect 199 139 200 140
rect 198 139 199 140
rect 197 139 198 140
rect 196 139 197 140
rect 195 139 196 140
rect 194 139 195 140
rect 193 139 194 140
rect 192 139 193 140
rect 191 139 192 140
rect 190 139 191 140
rect 189 139 190 140
rect 188 139 189 140
rect 187 139 188 140
rect 186 139 187 140
rect 185 139 186 140
rect 184 139 185 140
rect 183 139 184 140
rect 182 139 183 140
rect 181 139 182 140
rect 180 139 181 140
rect 179 139 180 140
rect 178 139 179 140
rect 177 139 178 140
rect 176 139 177 140
rect 175 139 176 140
rect 174 139 175 140
rect 173 139 174 140
rect 172 139 173 140
rect 171 139 172 140
rect 170 139 171 140
rect 169 139 170 140
rect 168 139 169 140
rect 167 139 168 140
rect 166 139 167 140
rect 165 139 166 140
rect 164 139 165 140
rect 163 139 164 140
rect 162 139 163 140
rect 161 139 162 140
rect 160 139 161 140
rect 141 139 142 140
rect 140 139 141 140
rect 139 139 140 140
rect 138 139 139 140
rect 137 139 138 140
rect 136 139 137 140
rect 135 139 136 140
rect 134 139 135 140
rect 133 139 134 140
rect 132 139 133 140
rect 131 139 132 140
rect 130 139 131 140
rect 129 139 130 140
rect 128 139 129 140
rect 127 139 128 140
rect 126 139 127 140
rect 125 139 126 140
rect 124 139 125 140
rect 123 139 124 140
rect 122 139 123 140
rect 121 139 122 140
rect 120 139 121 140
rect 119 139 120 140
rect 118 139 119 140
rect 117 139 118 140
rect 116 139 117 140
rect 115 139 116 140
rect 114 139 115 140
rect 113 139 114 140
rect 112 139 113 140
rect 111 139 112 140
rect 110 139 111 140
rect 109 139 110 140
rect 108 139 109 140
rect 107 139 108 140
rect 106 139 107 140
rect 105 139 106 140
rect 104 139 105 140
rect 103 139 104 140
rect 102 139 103 140
rect 101 139 102 140
rect 100 139 101 140
rect 99 139 100 140
rect 98 139 99 140
rect 97 139 98 140
rect 96 139 97 140
rect 95 139 96 140
rect 94 139 95 140
rect 93 139 94 140
rect 92 139 93 140
rect 91 139 92 140
rect 90 139 91 140
rect 89 139 90 140
rect 88 139 89 140
rect 87 139 88 140
rect 86 139 87 140
rect 85 139 86 140
rect 84 139 85 140
rect 83 139 84 140
rect 82 139 83 140
rect 81 139 82 140
rect 80 139 81 140
rect 79 139 80 140
rect 78 139 79 140
rect 77 139 78 140
rect 76 139 77 140
rect 75 139 76 140
rect 74 139 75 140
rect 73 139 74 140
rect 72 139 73 140
rect 71 139 72 140
rect 70 139 71 140
rect 69 139 70 140
rect 68 139 69 140
rect 67 139 68 140
rect 66 139 67 140
rect 65 139 66 140
rect 64 139 65 140
rect 63 139 64 140
rect 62 139 63 140
rect 61 139 62 140
rect 60 139 61 140
rect 59 139 60 140
rect 58 139 59 140
rect 57 139 58 140
rect 56 139 57 140
rect 55 139 56 140
rect 54 139 55 140
rect 53 139 54 140
rect 52 139 53 140
rect 51 139 52 140
rect 50 139 51 140
rect 49 139 50 140
rect 48 139 49 140
rect 47 139 48 140
rect 46 139 47 140
rect 45 139 46 140
rect 44 139 45 140
rect 43 139 44 140
rect 42 139 43 140
rect 41 139 42 140
rect 40 139 41 140
rect 39 139 40 140
rect 38 139 39 140
rect 37 139 38 140
rect 435 140 436 141
rect 434 140 435 141
rect 433 140 434 141
rect 432 140 433 141
rect 431 140 432 141
rect 430 140 431 141
rect 429 140 430 141
rect 428 140 429 141
rect 427 140 428 141
rect 426 140 427 141
rect 425 140 426 141
rect 424 140 425 141
rect 423 140 424 141
rect 422 140 423 141
rect 421 140 422 141
rect 420 140 421 141
rect 419 140 420 141
rect 418 140 419 141
rect 417 140 418 141
rect 416 140 417 141
rect 415 140 416 141
rect 414 140 415 141
rect 413 140 414 141
rect 412 140 413 141
rect 411 140 412 141
rect 410 140 411 141
rect 409 140 410 141
rect 408 140 409 141
rect 407 140 408 141
rect 406 140 407 141
rect 405 140 406 141
rect 404 140 405 141
rect 403 140 404 141
rect 402 140 403 141
rect 401 140 402 141
rect 400 140 401 141
rect 399 140 400 141
rect 398 140 399 141
rect 397 140 398 141
rect 396 140 397 141
rect 395 140 396 141
rect 313 140 314 141
rect 312 140 313 141
rect 311 140 312 141
rect 310 140 311 141
rect 309 140 310 141
rect 308 140 309 141
rect 307 140 308 141
rect 306 140 307 141
rect 305 140 306 141
rect 304 140 305 141
rect 303 140 304 141
rect 302 140 303 141
rect 301 140 302 141
rect 300 140 301 141
rect 299 140 300 141
rect 298 140 299 141
rect 297 140 298 141
rect 296 140 297 141
rect 295 140 296 141
rect 294 140 295 141
rect 293 140 294 141
rect 292 140 293 141
rect 291 140 292 141
rect 290 140 291 141
rect 289 140 290 141
rect 288 140 289 141
rect 287 140 288 141
rect 286 140 287 141
rect 285 140 286 141
rect 284 140 285 141
rect 283 140 284 141
rect 282 140 283 141
rect 281 140 282 141
rect 280 140 281 141
rect 279 140 280 141
rect 278 140 279 141
rect 277 140 278 141
rect 276 140 277 141
rect 275 140 276 141
rect 274 140 275 141
rect 273 140 274 141
rect 272 140 273 141
rect 271 140 272 141
rect 270 140 271 141
rect 269 140 270 141
rect 268 140 269 141
rect 267 140 268 141
rect 266 140 267 141
rect 265 140 266 141
rect 264 140 265 141
rect 263 140 264 141
rect 262 140 263 141
rect 261 140 262 141
rect 260 140 261 141
rect 259 140 260 141
rect 258 140 259 141
rect 257 140 258 141
rect 256 140 257 141
rect 255 140 256 141
rect 254 140 255 141
rect 253 140 254 141
rect 252 140 253 141
rect 251 140 252 141
rect 250 140 251 141
rect 249 140 250 141
rect 248 140 249 141
rect 247 140 248 141
rect 223 140 224 141
rect 222 140 223 141
rect 221 140 222 141
rect 220 140 221 141
rect 219 140 220 141
rect 218 140 219 141
rect 217 140 218 141
rect 216 140 217 141
rect 215 140 216 141
rect 214 140 215 141
rect 213 140 214 141
rect 212 140 213 141
rect 211 140 212 141
rect 210 140 211 141
rect 209 140 210 141
rect 208 140 209 141
rect 207 140 208 141
rect 206 140 207 141
rect 205 140 206 141
rect 204 140 205 141
rect 203 140 204 141
rect 202 140 203 141
rect 201 140 202 141
rect 200 140 201 141
rect 199 140 200 141
rect 198 140 199 141
rect 197 140 198 141
rect 196 140 197 141
rect 195 140 196 141
rect 194 140 195 141
rect 193 140 194 141
rect 192 140 193 141
rect 191 140 192 141
rect 190 140 191 141
rect 189 140 190 141
rect 188 140 189 141
rect 187 140 188 141
rect 186 140 187 141
rect 185 140 186 141
rect 184 140 185 141
rect 183 140 184 141
rect 182 140 183 141
rect 181 140 182 141
rect 180 140 181 141
rect 179 140 180 141
rect 178 140 179 141
rect 177 140 178 141
rect 176 140 177 141
rect 175 140 176 141
rect 174 140 175 141
rect 173 140 174 141
rect 172 140 173 141
rect 171 140 172 141
rect 170 140 171 141
rect 169 140 170 141
rect 168 140 169 141
rect 167 140 168 141
rect 166 140 167 141
rect 165 140 166 141
rect 164 140 165 141
rect 163 140 164 141
rect 162 140 163 141
rect 161 140 162 141
rect 160 140 161 141
rect 140 140 141 141
rect 139 140 140 141
rect 138 140 139 141
rect 137 140 138 141
rect 136 140 137 141
rect 135 140 136 141
rect 134 140 135 141
rect 133 140 134 141
rect 132 140 133 141
rect 131 140 132 141
rect 130 140 131 141
rect 129 140 130 141
rect 128 140 129 141
rect 127 140 128 141
rect 126 140 127 141
rect 125 140 126 141
rect 124 140 125 141
rect 123 140 124 141
rect 122 140 123 141
rect 121 140 122 141
rect 120 140 121 141
rect 119 140 120 141
rect 118 140 119 141
rect 117 140 118 141
rect 116 140 117 141
rect 115 140 116 141
rect 114 140 115 141
rect 113 140 114 141
rect 112 140 113 141
rect 111 140 112 141
rect 110 140 111 141
rect 109 140 110 141
rect 108 140 109 141
rect 107 140 108 141
rect 106 140 107 141
rect 105 140 106 141
rect 104 140 105 141
rect 103 140 104 141
rect 102 140 103 141
rect 101 140 102 141
rect 100 140 101 141
rect 99 140 100 141
rect 98 140 99 141
rect 97 140 98 141
rect 96 140 97 141
rect 95 140 96 141
rect 94 140 95 141
rect 93 140 94 141
rect 92 140 93 141
rect 91 140 92 141
rect 90 140 91 141
rect 89 140 90 141
rect 88 140 89 141
rect 87 140 88 141
rect 86 140 87 141
rect 85 140 86 141
rect 84 140 85 141
rect 83 140 84 141
rect 82 140 83 141
rect 81 140 82 141
rect 80 140 81 141
rect 79 140 80 141
rect 78 140 79 141
rect 77 140 78 141
rect 76 140 77 141
rect 75 140 76 141
rect 74 140 75 141
rect 73 140 74 141
rect 72 140 73 141
rect 71 140 72 141
rect 70 140 71 141
rect 69 140 70 141
rect 68 140 69 141
rect 67 140 68 141
rect 66 140 67 141
rect 65 140 66 141
rect 64 140 65 141
rect 63 140 64 141
rect 62 140 63 141
rect 61 140 62 141
rect 60 140 61 141
rect 59 140 60 141
rect 58 140 59 141
rect 57 140 58 141
rect 56 140 57 141
rect 55 140 56 141
rect 54 140 55 141
rect 53 140 54 141
rect 52 140 53 141
rect 51 140 52 141
rect 50 140 51 141
rect 49 140 50 141
rect 48 140 49 141
rect 47 140 48 141
rect 46 140 47 141
rect 45 140 46 141
rect 44 140 45 141
rect 43 140 44 141
rect 42 140 43 141
rect 41 140 42 141
rect 40 140 41 141
rect 39 140 40 141
rect 38 140 39 141
rect 433 141 434 142
rect 432 141 433 142
rect 431 141 432 142
rect 430 141 431 142
rect 429 141 430 142
rect 428 141 429 142
rect 427 141 428 142
rect 426 141 427 142
rect 425 141 426 142
rect 424 141 425 142
rect 423 141 424 142
rect 422 141 423 142
rect 421 141 422 142
rect 420 141 421 142
rect 419 141 420 142
rect 418 141 419 142
rect 417 141 418 142
rect 416 141 417 142
rect 415 141 416 142
rect 414 141 415 142
rect 413 141 414 142
rect 412 141 413 142
rect 411 141 412 142
rect 410 141 411 142
rect 409 141 410 142
rect 408 141 409 142
rect 407 141 408 142
rect 406 141 407 142
rect 405 141 406 142
rect 404 141 405 142
rect 403 141 404 142
rect 402 141 403 142
rect 401 141 402 142
rect 400 141 401 142
rect 399 141 400 142
rect 398 141 399 142
rect 397 141 398 142
rect 396 141 397 142
rect 395 141 396 142
rect 313 141 314 142
rect 312 141 313 142
rect 311 141 312 142
rect 310 141 311 142
rect 309 141 310 142
rect 308 141 309 142
rect 307 141 308 142
rect 306 141 307 142
rect 305 141 306 142
rect 304 141 305 142
rect 303 141 304 142
rect 302 141 303 142
rect 301 141 302 142
rect 300 141 301 142
rect 299 141 300 142
rect 298 141 299 142
rect 297 141 298 142
rect 296 141 297 142
rect 295 141 296 142
rect 294 141 295 142
rect 293 141 294 142
rect 292 141 293 142
rect 291 141 292 142
rect 290 141 291 142
rect 289 141 290 142
rect 288 141 289 142
rect 287 141 288 142
rect 286 141 287 142
rect 285 141 286 142
rect 284 141 285 142
rect 283 141 284 142
rect 282 141 283 142
rect 281 141 282 142
rect 280 141 281 142
rect 279 141 280 142
rect 278 141 279 142
rect 277 141 278 142
rect 276 141 277 142
rect 275 141 276 142
rect 274 141 275 142
rect 273 141 274 142
rect 272 141 273 142
rect 271 141 272 142
rect 270 141 271 142
rect 269 141 270 142
rect 268 141 269 142
rect 267 141 268 142
rect 266 141 267 142
rect 265 141 266 142
rect 264 141 265 142
rect 263 141 264 142
rect 262 141 263 142
rect 261 141 262 142
rect 260 141 261 142
rect 259 141 260 142
rect 258 141 259 142
rect 257 141 258 142
rect 256 141 257 142
rect 255 141 256 142
rect 254 141 255 142
rect 253 141 254 142
rect 252 141 253 142
rect 251 141 252 142
rect 250 141 251 142
rect 249 141 250 142
rect 248 141 249 142
rect 247 141 248 142
rect 246 141 247 142
rect 222 141 223 142
rect 221 141 222 142
rect 220 141 221 142
rect 219 141 220 142
rect 218 141 219 142
rect 217 141 218 142
rect 216 141 217 142
rect 215 141 216 142
rect 214 141 215 142
rect 213 141 214 142
rect 212 141 213 142
rect 211 141 212 142
rect 210 141 211 142
rect 209 141 210 142
rect 208 141 209 142
rect 207 141 208 142
rect 206 141 207 142
rect 205 141 206 142
rect 204 141 205 142
rect 203 141 204 142
rect 202 141 203 142
rect 201 141 202 142
rect 200 141 201 142
rect 199 141 200 142
rect 198 141 199 142
rect 197 141 198 142
rect 196 141 197 142
rect 195 141 196 142
rect 194 141 195 142
rect 193 141 194 142
rect 192 141 193 142
rect 191 141 192 142
rect 190 141 191 142
rect 189 141 190 142
rect 188 141 189 142
rect 187 141 188 142
rect 186 141 187 142
rect 185 141 186 142
rect 184 141 185 142
rect 183 141 184 142
rect 182 141 183 142
rect 181 141 182 142
rect 180 141 181 142
rect 179 141 180 142
rect 178 141 179 142
rect 177 141 178 142
rect 176 141 177 142
rect 175 141 176 142
rect 174 141 175 142
rect 173 141 174 142
rect 172 141 173 142
rect 171 141 172 142
rect 170 141 171 142
rect 169 141 170 142
rect 168 141 169 142
rect 167 141 168 142
rect 166 141 167 142
rect 165 141 166 142
rect 164 141 165 142
rect 163 141 164 142
rect 162 141 163 142
rect 161 141 162 142
rect 160 141 161 142
rect 159 141 160 142
rect 139 141 140 142
rect 138 141 139 142
rect 137 141 138 142
rect 136 141 137 142
rect 135 141 136 142
rect 134 141 135 142
rect 133 141 134 142
rect 132 141 133 142
rect 131 141 132 142
rect 130 141 131 142
rect 129 141 130 142
rect 128 141 129 142
rect 127 141 128 142
rect 126 141 127 142
rect 125 141 126 142
rect 124 141 125 142
rect 123 141 124 142
rect 122 141 123 142
rect 121 141 122 142
rect 120 141 121 142
rect 119 141 120 142
rect 118 141 119 142
rect 117 141 118 142
rect 116 141 117 142
rect 115 141 116 142
rect 114 141 115 142
rect 113 141 114 142
rect 112 141 113 142
rect 111 141 112 142
rect 110 141 111 142
rect 109 141 110 142
rect 108 141 109 142
rect 107 141 108 142
rect 106 141 107 142
rect 105 141 106 142
rect 104 141 105 142
rect 103 141 104 142
rect 102 141 103 142
rect 101 141 102 142
rect 100 141 101 142
rect 99 141 100 142
rect 98 141 99 142
rect 97 141 98 142
rect 96 141 97 142
rect 95 141 96 142
rect 94 141 95 142
rect 93 141 94 142
rect 92 141 93 142
rect 91 141 92 142
rect 90 141 91 142
rect 89 141 90 142
rect 88 141 89 142
rect 87 141 88 142
rect 86 141 87 142
rect 85 141 86 142
rect 84 141 85 142
rect 83 141 84 142
rect 82 141 83 142
rect 81 141 82 142
rect 80 141 81 142
rect 79 141 80 142
rect 78 141 79 142
rect 77 141 78 142
rect 76 141 77 142
rect 75 141 76 142
rect 74 141 75 142
rect 73 141 74 142
rect 72 141 73 142
rect 71 141 72 142
rect 70 141 71 142
rect 69 141 70 142
rect 68 141 69 142
rect 67 141 68 142
rect 66 141 67 142
rect 65 141 66 142
rect 64 141 65 142
rect 63 141 64 142
rect 62 141 63 142
rect 61 141 62 142
rect 60 141 61 142
rect 59 141 60 142
rect 58 141 59 142
rect 57 141 58 142
rect 56 141 57 142
rect 55 141 56 142
rect 54 141 55 142
rect 53 141 54 142
rect 52 141 53 142
rect 51 141 52 142
rect 50 141 51 142
rect 49 141 50 142
rect 48 141 49 142
rect 47 141 48 142
rect 46 141 47 142
rect 45 141 46 142
rect 44 141 45 142
rect 43 141 44 142
rect 42 141 43 142
rect 41 141 42 142
rect 40 141 41 142
rect 39 141 40 142
rect 480 142 481 143
rect 460 142 461 143
rect 431 142 432 143
rect 430 142 431 143
rect 429 142 430 143
rect 428 142 429 143
rect 427 142 428 143
rect 426 142 427 143
rect 425 142 426 143
rect 424 142 425 143
rect 423 142 424 143
rect 422 142 423 143
rect 421 142 422 143
rect 420 142 421 143
rect 419 142 420 143
rect 418 142 419 143
rect 417 142 418 143
rect 416 142 417 143
rect 415 142 416 143
rect 414 142 415 143
rect 413 142 414 143
rect 412 142 413 143
rect 411 142 412 143
rect 410 142 411 143
rect 409 142 410 143
rect 408 142 409 143
rect 407 142 408 143
rect 406 142 407 143
rect 405 142 406 143
rect 404 142 405 143
rect 403 142 404 143
rect 402 142 403 143
rect 401 142 402 143
rect 400 142 401 143
rect 399 142 400 143
rect 398 142 399 143
rect 397 142 398 143
rect 396 142 397 143
rect 395 142 396 143
rect 314 142 315 143
rect 313 142 314 143
rect 312 142 313 143
rect 311 142 312 143
rect 310 142 311 143
rect 309 142 310 143
rect 308 142 309 143
rect 307 142 308 143
rect 306 142 307 143
rect 305 142 306 143
rect 304 142 305 143
rect 303 142 304 143
rect 302 142 303 143
rect 301 142 302 143
rect 300 142 301 143
rect 299 142 300 143
rect 298 142 299 143
rect 297 142 298 143
rect 296 142 297 143
rect 295 142 296 143
rect 294 142 295 143
rect 293 142 294 143
rect 292 142 293 143
rect 291 142 292 143
rect 290 142 291 143
rect 289 142 290 143
rect 288 142 289 143
rect 287 142 288 143
rect 286 142 287 143
rect 285 142 286 143
rect 284 142 285 143
rect 283 142 284 143
rect 282 142 283 143
rect 281 142 282 143
rect 280 142 281 143
rect 279 142 280 143
rect 278 142 279 143
rect 277 142 278 143
rect 276 142 277 143
rect 275 142 276 143
rect 274 142 275 143
rect 273 142 274 143
rect 272 142 273 143
rect 271 142 272 143
rect 270 142 271 143
rect 269 142 270 143
rect 268 142 269 143
rect 267 142 268 143
rect 266 142 267 143
rect 265 142 266 143
rect 264 142 265 143
rect 263 142 264 143
rect 262 142 263 143
rect 261 142 262 143
rect 260 142 261 143
rect 259 142 260 143
rect 258 142 259 143
rect 257 142 258 143
rect 256 142 257 143
rect 255 142 256 143
rect 254 142 255 143
rect 253 142 254 143
rect 252 142 253 143
rect 251 142 252 143
rect 250 142 251 143
rect 249 142 250 143
rect 248 142 249 143
rect 247 142 248 143
rect 246 142 247 143
rect 245 142 246 143
rect 222 142 223 143
rect 221 142 222 143
rect 220 142 221 143
rect 219 142 220 143
rect 218 142 219 143
rect 217 142 218 143
rect 216 142 217 143
rect 215 142 216 143
rect 214 142 215 143
rect 213 142 214 143
rect 212 142 213 143
rect 211 142 212 143
rect 210 142 211 143
rect 209 142 210 143
rect 208 142 209 143
rect 207 142 208 143
rect 206 142 207 143
rect 205 142 206 143
rect 204 142 205 143
rect 203 142 204 143
rect 202 142 203 143
rect 201 142 202 143
rect 200 142 201 143
rect 199 142 200 143
rect 198 142 199 143
rect 197 142 198 143
rect 196 142 197 143
rect 195 142 196 143
rect 194 142 195 143
rect 193 142 194 143
rect 192 142 193 143
rect 191 142 192 143
rect 190 142 191 143
rect 189 142 190 143
rect 188 142 189 143
rect 187 142 188 143
rect 186 142 187 143
rect 185 142 186 143
rect 184 142 185 143
rect 183 142 184 143
rect 182 142 183 143
rect 181 142 182 143
rect 180 142 181 143
rect 179 142 180 143
rect 178 142 179 143
rect 177 142 178 143
rect 176 142 177 143
rect 175 142 176 143
rect 174 142 175 143
rect 173 142 174 143
rect 172 142 173 143
rect 171 142 172 143
rect 170 142 171 143
rect 169 142 170 143
rect 168 142 169 143
rect 167 142 168 143
rect 166 142 167 143
rect 165 142 166 143
rect 164 142 165 143
rect 163 142 164 143
rect 162 142 163 143
rect 161 142 162 143
rect 160 142 161 143
rect 159 142 160 143
rect 138 142 139 143
rect 137 142 138 143
rect 136 142 137 143
rect 135 142 136 143
rect 134 142 135 143
rect 133 142 134 143
rect 132 142 133 143
rect 131 142 132 143
rect 130 142 131 143
rect 129 142 130 143
rect 128 142 129 143
rect 127 142 128 143
rect 126 142 127 143
rect 125 142 126 143
rect 124 142 125 143
rect 123 142 124 143
rect 122 142 123 143
rect 121 142 122 143
rect 120 142 121 143
rect 119 142 120 143
rect 118 142 119 143
rect 117 142 118 143
rect 116 142 117 143
rect 115 142 116 143
rect 114 142 115 143
rect 113 142 114 143
rect 112 142 113 143
rect 111 142 112 143
rect 110 142 111 143
rect 109 142 110 143
rect 108 142 109 143
rect 107 142 108 143
rect 106 142 107 143
rect 105 142 106 143
rect 104 142 105 143
rect 103 142 104 143
rect 102 142 103 143
rect 101 142 102 143
rect 100 142 101 143
rect 99 142 100 143
rect 98 142 99 143
rect 97 142 98 143
rect 96 142 97 143
rect 95 142 96 143
rect 94 142 95 143
rect 93 142 94 143
rect 92 142 93 143
rect 91 142 92 143
rect 90 142 91 143
rect 89 142 90 143
rect 88 142 89 143
rect 87 142 88 143
rect 86 142 87 143
rect 85 142 86 143
rect 84 142 85 143
rect 83 142 84 143
rect 82 142 83 143
rect 81 142 82 143
rect 80 142 81 143
rect 79 142 80 143
rect 78 142 79 143
rect 77 142 78 143
rect 76 142 77 143
rect 75 142 76 143
rect 74 142 75 143
rect 73 142 74 143
rect 72 142 73 143
rect 71 142 72 143
rect 70 142 71 143
rect 69 142 70 143
rect 68 142 69 143
rect 67 142 68 143
rect 66 142 67 143
rect 65 142 66 143
rect 64 142 65 143
rect 63 142 64 143
rect 62 142 63 143
rect 61 142 62 143
rect 60 142 61 143
rect 59 142 60 143
rect 58 142 59 143
rect 57 142 58 143
rect 56 142 57 143
rect 55 142 56 143
rect 54 142 55 143
rect 53 142 54 143
rect 52 142 53 143
rect 51 142 52 143
rect 50 142 51 143
rect 49 142 50 143
rect 48 142 49 143
rect 47 142 48 143
rect 46 142 47 143
rect 45 142 46 143
rect 44 142 45 143
rect 43 142 44 143
rect 42 142 43 143
rect 41 142 42 143
rect 40 142 41 143
rect 39 142 40 143
rect 24 142 25 143
rect 23 142 24 143
rect 22 142 23 143
rect 21 142 22 143
rect 20 142 21 143
rect 480 143 481 144
rect 460 143 461 144
rect 427 143 428 144
rect 426 143 427 144
rect 425 143 426 144
rect 424 143 425 144
rect 423 143 424 144
rect 422 143 423 144
rect 421 143 422 144
rect 420 143 421 144
rect 419 143 420 144
rect 418 143 419 144
rect 417 143 418 144
rect 416 143 417 144
rect 415 143 416 144
rect 414 143 415 144
rect 413 143 414 144
rect 412 143 413 144
rect 411 143 412 144
rect 410 143 411 144
rect 409 143 410 144
rect 408 143 409 144
rect 407 143 408 144
rect 406 143 407 144
rect 405 143 406 144
rect 404 143 405 144
rect 403 143 404 144
rect 402 143 403 144
rect 401 143 402 144
rect 400 143 401 144
rect 399 143 400 144
rect 398 143 399 144
rect 397 143 398 144
rect 396 143 397 144
rect 395 143 396 144
rect 315 143 316 144
rect 314 143 315 144
rect 313 143 314 144
rect 312 143 313 144
rect 311 143 312 144
rect 310 143 311 144
rect 309 143 310 144
rect 308 143 309 144
rect 307 143 308 144
rect 306 143 307 144
rect 305 143 306 144
rect 304 143 305 144
rect 303 143 304 144
rect 302 143 303 144
rect 301 143 302 144
rect 300 143 301 144
rect 299 143 300 144
rect 298 143 299 144
rect 297 143 298 144
rect 296 143 297 144
rect 295 143 296 144
rect 294 143 295 144
rect 293 143 294 144
rect 292 143 293 144
rect 291 143 292 144
rect 290 143 291 144
rect 289 143 290 144
rect 288 143 289 144
rect 287 143 288 144
rect 286 143 287 144
rect 285 143 286 144
rect 284 143 285 144
rect 283 143 284 144
rect 282 143 283 144
rect 281 143 282 144
rect 280 143 281 144
rect 279 143 280 144
rect 278 143 279 144
rect 277 143 278 144
rect 276 143 277 144
rect 275 143 276 144
rect 274 143 275 144
rect 273 143 274 144
rect 272 143 273 144
rect 271 143 272 144
rect 270 143 271 144
rect 269 143 270 144
rect 268 143 269 144
rect 267 143 268 144
rect 266 143 267 144
rect 265 143 266 144
rect 264 143 265 144
rect 263 143 264 144
rect 262 143 263 144
rect 261 143 262 144
rect 260 143 261 144
rect 259 143 260 144
rect 258 143 259 144
rect 257 143 258 144
rect 256 143 257 144
rect 255 143 256 144
rect 254 143 255 144
rect 253 143 254 144
rect 252 143 253 144
rect 251 143 252 144
rect 250 143 251 144
rect 249 143 250 144
rect 248 143 249 144
rect 247 143 248 144
rect 246 143 247 144
rect 245 143 246 144
rect 244 143 245 144
rect 221 143 222 144
rect 220 143 221 144
rect 219 143 220 144
rect 218 143 219 144
rect 217 143 218 144
rect 216 143 217 144
rect 215 143 216 144
rect 214 143 215 144
rect 213 143 214 144
rect 212 143 213 144
rect 211 143 212 144
rect 210 143 211 144
rect 209 143 210 144
rect 208 143 209 144
rect 207 143 208 144
rect 206 143 207 144
rect 205 143 206 144
rect 204 143 205 144
rect 203 143 204 144
rect 202 143 203 144
rect 201 143 202 144
rect 200 143 201 144
rect 199 143 200 144
rect 198 143 199 144
rect 197 143 198 144
rect 196 143 197 144
rect 195 143 196 144
rect 194 143 195 144
rect 193 143 194 144
rect 192 143 193 144
rect 191 143 192 144
rect 190 143 191 144
rect 189 143 190 144
rect 188 143 189 144
rect 187 143 188 144
rect 186 143 187 144
rect 185 143 186 144
rect 184 143 185 144
rect 183 143 184 144
rect 182 143 183 144
rect 181 143 182 144
rect 180 143 181 144
rect 179 143 180 144
rect 178 143 179 144
rect 177 143 178 144
rect 176 143 177 144
rect 175 143 176 144
rect 174 143 175 144
rect 173 143 174 144
rect 172 143 173 144
rect 171 143 172 144
rect 170 143 171 144
rect 169 143 170 144
rect 168 143 169 144
rect 167 143 168 144
rect 166 143 167 144
rect 165 143 166 144
rect 164 143 165 144
rect 163 143 164 144
rect 162 143 163 144
rect 161 143 162 144
rect 160 143 161 144
rect 159 143 160 144
rect 158 143 159 144
rect 137 143 138 144
rect 136 143 137 144
rect 135 143 136 144
rect 134 143 135 144
rect 133 143 134 144
rect 132 143 133 144
rect 131 143 132 144
rect 130 143 131 144
rect 129 143 130 144
rect 128 143 129 144
rect 127 143 128 144
rect 126 143 127 144
rect 125 143 126 144
rect 124 143 125 144
rect 123 143 124 144
rect 122 143 123 144
rect 121 143 122 144
rect 120 143 121 144
rect 119 143 120 144
rect 118 143 119 144
rect 117 143 118 144
rect 116 143 117 144
rect 115 143 116 144
rect 114 143 115 144
rect 113 143 114 144
rect 112 143 113 144
rect 111 143 112 144
rect 110 143 111 144
rect 109 143 110 144
rect 108 143 109 144
rect 107 143 108 144
rect 106 143 107 144
rect 105 143 106 144
rect 104 143 105 144
rect 103 143 104 144
rect 102 143 103 144
rect 101 143 102 144
rect 100 143 101 144
rect 99 143 100 144
rect 98 143 99 144
rect 97 143 98 144
rect 96 143 97 144
rect 95 143 96 144
rect 94 143 95 144
rect 93 143 94 144
rect 92 143 93 144
rect 91 143 92 144
rect 90 143 91 144
rect 89 143 90 144
rect 88 143 89 144
rect 87 143 88 144
rect 86 143 87 144
rect 85 143 86 144
rect 84 143 85 144
rect 83 143 84 144
rect 82 143 83 144
rect 81 143 82 144
rect 80 143 81 144
rect 79 143 80 144
rect 78 143 79 144
rect 77 143 78 144
rect 76 143 77 144
rect 75 143 76 144
rect 74 143 75 144
rect 73 143 74 144
rect 72 143 73 144
rect 71 143 72 144
rect 70 143 71 144
rect 69 143 70 144
rect 68 143 69 144
rect 67 143 68 144
rect 66 143 67 144
rect 65 143 66 144
rect 64 143 65 144
rect 63 143 64 144
rect 62 143 63 144
rect 61 143 62 144
rect 60 143 61 144
rect 59 143 60 144
rect 58 143 59 144
rect 57 143 58 144
rect 56 143 57 144
rect 55 143 56 144
rect 54 143 55 144
rect 53 143 54 144
rect 52 143 53 144
rect 51 143 52 144
rect 50 143 51 144
rect 49 143 50 144
rect 48 143 49 144
rect 47 143 48 144
rect 46 143 47 144
rect 45 143 46 144
rect 44 143 45 144
rect 43 143 44 144
rect 42 143 43 144
rect 41 143 42 144
rect 40 143 41 144
rect 26 143 27 144
rect 25 143 26 144
rect 24 143 25 144
rect 23 143 24 144
rect 22 143 23 144
rect 21 143 22 144
rect 20 143 21 144
rect 19 143 20 144
rect 18 143 19 144
rect 17 143 18 144
rect 480 144 481 145
rect 479 144 480 145
rect 461 144 462 145
rect 460 144 461 145
rect 404 144 405 145
rect 403 144 404 145
rect 402 144 403 145
rect 401 144 402 145
rect 400 144 401 145
rect 399 144 400 145
rect 398 144 399 145
rect 397 144 398 145
rect 396 144 397 145
rect 395 144 396 145
rect 316 144 317 145
rect 315 144 316 145
rect 314 144 315 145
rect 313 144 314 145
rect 312 144 313 145
rect 311 144 312 145
rect 310 144 311 145
rect 309 144 310 145
rect 308 144 309 145
rect 307 144 308 145
rect 306 144 307 145
rect 305 144 306 145
rect 304 144 305 145
rect 303 144 304 145
rect 302 144 303 145
rect 301 144 302 145
rect 300 144 301 145
rect 299 144 300 145
rect 298 144 299 145
rect 297 144 298 145
rect 296 144 297 145
rect 295 144 296 145
rect 294 144 295 145
rect 293 144 294 145
rect 292 144 293 145
rect 291 144 292 145
rect 290 144 291 145
rect 289 144 290 145
rect 288 144 289 145
rect 287 144 288 145
rect 286 144 287 145
rect 285 144 286 145
rect 284 144 285 145
rect 283 144 284 145
rect 282 144 283 145
rect 281 144 282 145
rect 280 144 281 145
rect 279 144 280 145
rect 278 144 279 145
rect 277 144 278 145
rect 276 144 277 145
rect 275 144 276 145
rect 274 144 275 145
rect 273 144 274 145
rect 272 144 273 145
rect 271 144 272 145
rect 270 144 271 145
rect 269 144 270 145
rect 268 144 269 145
rect 267 144 268 145
rect 266 144 267 145
rect 265 144 266 145
rect 264 144 265 145
rect 263 144 264 145
rect 262 144 263 145
rect 261 144 262 145
rect 260 144 261 145
rect 259 144 260 145
rect 258 144 259 145
rect 257 144 258 145
rect 256 144 257 145
rect 255 144 256 145
rect 254 144 255 145
rect 253 144 254 145
rect 252 144 253 145
rect 251 144 252 145
rect 250 144 251 145
rect 249 144 250 145
rect 248 144 249 145
rect 247 144 248 145
rect 246 144 247 145
rect 245 144 246 145
rect 244 144 245 145
rect 243 144 244 145
rect 221 144 222 145
rect 220 144 221 145
rect 219 144 220 145
rect 218 144 219 145
rect 217 144 218 145
rect 216 144 217 145
rect 215 144 216 145
rect 214 144 215 145
rect 213 144 214 145
rect 212 144 213 145
rect 211 144 212 145
rect 210 144 211 145
rect 209 144 210 145
rect 208 144 209 145
rect 207 144 208 145
rect 206 144 207 145
rect 205 144 206 145
rect 204 144 205 145
rect 203 144 204 145
rect 202 144 203 145
rect 201 144 202 145
rect 200 144 201 145
rect 199 144 200 145
rect 198 144 199 145
rect 197 144 198 145
rect 196 144 197 145
rect 195 144 196 145
rect 194 144 195 145
rect 193 144 194 145
rect 192 144 193 145
rect 191 144 192 145
rect 190 144 191 145
rect 189 144 190 145
rect 188 144 189 145
rect 187 144 188 145
rect 186 144 187 145
rect 185 144 186 145
rect 184 144 185 145
rect 183 144 184 145
rect 182 144 183 145
rect 181 144 182 145
rect 180 144 181 145
rect 179 144 180 145
rect 178 144 179 145
rect 177 144 178 145
rect 176 144 177 145
rect 175 144 176 145
rect 174 144 175 145
rect 173 144 174 145
rect 172 144 173 145
rect 171 144 172 145
rect 170 144 171 145
rect 169 144 170 145
rect 168 144 169 145
rect 167 144 168 145
rect 166 144 167 145
rect 165 144 166 145
rect 164 144 165 145
rect 163 144 164 145
rect 162 144 163 145
rect 161 144 162 145
rect 160 144 161 145
rect 159 144 160 145
rect 158 144 159 145
rect 136 144 137 145
rect 135 144 136 145
rect 134 144 135 145
rect 133 144 134 145
rect 132 144 133 145
rect 131 144 132 145
rect 130 144 131 145
rect 129 144 130 145
rect 128 144 129 145
rect 127 144 128 145
rect 126 144 127 145
rect 125 144 126 145
rect 124 144 125 145
rect 123 144 124 145
rect 122 144 123 145
rect 121 144 122 145
rect 120 144 121 145
rect 119 144 120 145
rect 118 144 119 145
rect 117 144 118 145
rect 116 144 117 145
rect 115 144 116 145
rect 114 144 115 145
rect 113 144 114 145
rect 112 144 113 145
rect 111 144 112 145
rect 110 144 111 145
rect 109 144 110 145
rect 108 144 109 145
rect 107 144 108 145
rect 106 144 107 145
rect 105 144 106 145
rect 104 144 105 145
rect 103 144 104 145
rect 102 144 103 145
rect 101 144 102 145
rect 100 144 101 145
rect 99 144 100 145
rect 98 144 99 145
rect 97 144 98 145
rect 96 144 97 145
rect 95 144 96 145
rect 94 144 95 145
rect 93 144 94 145
rect 92 144 93 145
rect 91 144 92 145
rect 90 144 91 145
rect 89 144 90 145
rect 88 144 89 145
rect 87 144 88 145
rect 86 144 87 145
rect 85 144 86 145
rect 84 144 85 145
rect 83 144 84 145
rect 82 144 83 145
rect 81 144 82 145
rect 80 144 81 145
rect 79 144 80 145
rect 78 144 79 145
rect 77 144 78 145
rect 76 144 77 145
rect 75 144 76 145
rect 74 144 75 145
rect 73 144 74 145
rect 72 144 73 145
rect 71 144 72 145
rect 70 144 71 145
rect 69 144 70 145
rect 68 144 69 145
rect 67 144 68 145
rect 66 144 67 145
rect 65 144 66 145
rect 64 144 65 145
rect 63 144 64 145
rect 62 144 63 145
rect 61 144 62 145
rect 60 144 61 145
rect 59 144 60 145
rect 58 144 59 145
rect 57 144 58 145
rect 56 144 57 145
rect 55 144 56 145
rect 54 144 55 145
rect 53 144 54 145
rect 52 144 53 145
rect 51 144 52 145
rect 50 144 51 145
rect 49 144 50 145
rect 48 144 49 145
rect 47 144 48 145
rect 46 144 47 145
rect 45 144 46 145
rect 44 144 45 145
rect 43 144 44 145
rect 42 144 43 145
rect 41 144 42 145
rect 40 144 41 145
rect 27 144 28 145
rect 26 144 27 145
rect 25 144 26 145
rect 24 144 25 145
rect 23 144 24 145
rect 22 144 23 145
rect 21 144 22 145
rect 20 144 21 145
rect 19 144 20 145
rect 18 144 19 145
rect 17 144 18 145
rect 16 144 17 145
rect 480 145 481 146
rect 479 145 480 146
rect 478 145 479 146
rect 477 145 478 146
rect 476 145 477 146
rect 475 145 476 146
rect 474 145 475 146
rect 473 145 474 146
rect 472 145 473 146
rect 471 145 472 146
rect 470 145 471 146
rect 469 145 470 146
rect 468 145 469 146
rect 467 145 468 146
rect 466 145 467 146
rect 465 145 466 146
rect 464 145 465 146
rect 463 145 464 146
rect 462 145 463 146
rect 461 145 462 146
rect 460 145 461 146
rect 399 145 400 146
rect 398 145 399 146
rect 397 145 398 146
rect 396 145 397 146
rect 395 145 396 146
rect 316 145 317 146
rect 315 145 316 146
rect 314 145 315 146
rect 313 145 314 146
rect 312 145 313 146
rect 311 145 312 146
rect 310 145 311 146
rect 309 145 310 146
rect 308 145 309 146
rect 307 145 308 146
rect 306 145 307 146
rect 305 145 306 146
rect 304 145 305 146
rect 303 145 304 146
rect 302 145 303 146
rect 301 145 302 146
rect 300 145 301 146
rect 299 145 300 146
rect 298 145 299 146
rect 297 145 298 146
rect 296 145 297 146
rect 295 145 296 146
rect 294 145 295 146
rect 293 145 294 146
rect 292 145 293 146
rect 291 145 292 146
rect 290 145 291 146
rect 289 145 290 146
rect 288 145 289 146
rect 287 145 288 146
rect 286 145 287 146
rect 285 145 286 146
rect 284 145 285 146
rect 283 145 284 146
rect 282 145 283 146
rect 281 145 282 146
rect 280 145 281 146
rect 279 145 280 146
rect 278 145 279 146
rect 277 145 278 146
rect 276 145 277 146
rect 275 145 276 146
rect 274 145 275 146
rect 273 145 274 146
rect 272 145 273 146
rect 271 145 272 146
rect 270 145 271 146
rect 269 145 270 146
rect 268 145 269 146
rect 267 145 268 146
rect 266 145 267 146
rect 265 145 266 146
rect 264 145 265 146
rect 263 145 264 146
rect 262 145 263 146
rect 261 145 262 146
rect 260 145 261 146
rect 259 145 260 146
rect 258 145 259 146
rect 257 145 258 146
rect 256 145 257 146
rect 255 145 256 146
rect 254 145 255 146
rect 253 145 254 146
rect 252 145 253 146
rect 251 145 252 146
rect 250 145 251 146
rect 249 145 250 146
rect 248 145 249 146
rect 247 145 248 146
rect 246 145 247 146
rect 245 145 246 146
rect 244 145 245 146
rect 243 145 244 146
rect 221 145 222 146
rect 220 145 221 146
rect 219 145 220 146
rect 218 145 219 146
rect 217 145 218 146
rect 216 145 217 146
rect 215 145 216 146
rect 214 145 215 146
rect 213 145 214 146
rect 212 145 213 146
rect 211 145 212 146
rect 210 145 211 146
rect 209 145 210 146
rect 208 145 209 146
rect 207 145 208 146
rect 206 145 207 146
rect 205 145 206 146
rect 204 145 205 146
rect 203 145 204 146
rect 202 145 203 146
rect 201 145 202 146
rect 200 145 201 146
rect 199 145 200 146
rect 198 145 199 146
rect 197 145 198 146
rect 196 145 197 146
rect 195 145 196 146
rect 194 145 195 146
rect 193 145 194 146
rect 192 145 193 146
rect 191 145 192 146
rect 190 145 191 146
rect 189 145 190 146
rect 188 145 189 146
rect 187 145 188 146
rect 186 145 187 146
rect 185 145 186 146
rect 184 145 185 146
rect 183 145 184 146
rect 182 145 183 146
rect 181 145 182 146
rect 180 145 181 146
rect 179 145 180 146
rect 178 145 179 146
rect 177 145 178 146
rect 176 145 177 146
rect 175 145 176 146
rect 174 145 175 146
rect 173 145 174 146
rect 172 145 173 146
rect 171 145 172 146
rect 170 145 171 146
rect 169 145 170 146
rect 168 145 169 146
rect 167 145 168 146
rect 166 145 167 146
rect 165 145 166 146
rect 164 145 165 146
rect 163 145 164 146
rect 162 145 163 146
rect 161 145 162 146
rect 160 145 161 146
rect 159 145 160 146
rect 158 145 159 146
rect 157 145 158 146
rect 135 145 136 146
rect 134 145 135 146
rect 133 145 134 146
rect 132 145 133 146
rect 131 145 132 146
rect 130 145 131 146
rect 129 145 130 146
rect 128 145 129 146
rect 127 145 128 146
rect 126 145 127 146
rect 125 145 126 146
rect 124 145 125 146
rect 123 145 124 146
rect 122 145 123 146
rect 121 145 122 146
rect 120 145 121 146
rect 119 145 120 146
rect 118 145 119 146
rect 117 145 118 146
rect 116 145 117 146
rect 115 145 116 146
rect 114 145 115 146
rect 113 145 114 146
rect 112 145 113 146
rect 111 145 112 146
rect 110 145 111 146
rect 109 145 110 146
rect 108 145 109 146
rect 107 145 108 146
rect 106 145 107 146
rect 105 145 106 146
rect 104 145 105 146
rect 103 145 104 146
rect 102 145 103 146
rect 101 145 102 146
rect 100 145 101 146
rect 99 145 100 146
rect 98 145 99 146
rect 97 145 98 146
rect 96 145 97 146
rect 95 145 96 146
rect 94 145 95 146
rect 93 145 94 146
rect 92 145 93 146
rect 91 145 92 146
rect 90 145 91 146
rect 89 145 90 146
rect 88 145 89 146
rect 87 145 88 146
rect 86 145 87 146
rect 85 145 86 146
rect 84 145 85 146
rect 83 145 84 146
rect 82 145 83 146
rect 81 145 82 146
rect 80 145 81 146
rect 79 145 80 146
rect 78 145 79 146
rect 77 145 78 146
rect 76 145 77 146
rect 75 145 76 146
rect 74 145 75 146
rect 73 145 74 146
rect 72 145 73 146
rect 71 145 72 146
rect 70 145 71 146
rect 69 145 70 146
rect 68 145 69 146
rect 67 145 68 146
rect 66 145 67 146
rect 65 145 66 146
rect 64 145 65 146
rect 63 145 64 146
rect 62 145 63 146
rect 61 145 62 146
rect 60 145 61 146
rect 59 145 60 146
rect 58 145 59 146
rect 57 145 58 146
rect 56 145 57 146
rect 55 145 56 146
rect 54 145 55 146
rect 53 145 54 146
rect 52 145 53 146
rect 51 145 52 146
rect 50 145 51 146
rect 49 145 50 146
rect 48 145 49 146
rect 47 145 48 146
rect 46 145 47 146
rect 45 145 46 146
rect 44 145 45 146
rect 43 145 44 146
rect 42 145 43 146
rect 41 145 42 146
rect 40 145 41 146
rect 28 145 29 146
rect 27 145 28 146
rect 26 145 27 146
rect 25 145 26 146
rect 24 145 25 146
rect 23 145 24 146
rect 22 145 23 146
rect 21 145 22 146
rect 20 145 21 146
rect 19 145 20 146
rect 18 145 19 146
rect 17 145 18 146
rect 16 145 17 146
rect 15 145 16 146
rect 14 145 15 146
rect 480 146 481 147
rect 479 146 480 147
rect 478 146 479 147
rect 477 146 478 147
rect 476 146 477 147
rect 475 146 476 147
rect 474 146 475 147
rect 473 146 474 147
rect 472 146 473 147
rect 471 146 472 147
rect 470 146 471 147
rect 469 146 470 147
rect 468 146 469 147
rect 467 146 468 147
rect 466 146 467 147
rect 465 146 466 147
rect 464 146 465 147
rect 463 146 464 147
rect 462 146 463 147
rect 461 146 462 147
rect 460 146 461 147
rect 398 146 399 147
rect 397 146 398 147
rect 396 146 397 147
rect 395 146 396 147
rect 317 146 318 147
rect 316 146 317 147
rect 315 146 316 147
rect 314 146 315 147
rect 313 146 314 147
rect 312 146 313 147
rect 311 146 312 147
rect 310 146 311 147
rect 309 146 310 147
rect 308 146 309 147
rect 307 146 308 147
rect 306 146 307 147
rect 305 146 306 147
rect 304 146 305 147
rect 303 146 304 147
rect 302 146 303 147
rect 301 146 302 147
rect 300 146 301 147
rect 299 146 300 147
rect 298 146 299 147
rect 297 146 298 147
rect 296 146 297 147
rect 295 146 296 147
rect 294 146 295 147
rect 293 146 294 147
rect 292 146 293 147
rect 291 146 292 147
rect 290 146 291 147
rect 289 146 290 147
rect 288 146 289 147
rect 287 146 288 147
rect 286 146 287 147
rect 285 146 286 147
rect 284 146 285 147
rect 283 146 284 147
rect 282 146 283 147
rect 281 146 282 147
rect 280 146 281 147
rect 279 146 280 147
rect 278 146 279 147
rect 277 146 278 147
rect 276 146 277 147
rect 275 146 276 147
rect 274 146 275 147
rect 273 146 274 147
rect 272 146 273 147
rect 271 146 272 147
rect 270 146 271 147
rect 269 146 270 147
rect 268 146 269 147
rect 267 146 268 147
rect 266 146 267 147
rect 265 146 266 147
rect 264 146 265 147
rect 263 146 264 147
rect 262 146 263 147
rect 261 146 262 147
rect 260 146 261 147
rect 259 146 260 147
rect 258 146 259 147
rect 257 146 258 147
rect 256 146 257 147
rect 255 146 256 147
rect 254 146 255 147
rect 253 146 254 147
rect 252 146 253 147
rect 251 146 252 147
rect 250 146 251 147
rect 249 146 250 147
rect 248 146 249 147
rect 247 146 248 147
rect 246 146 247 147
rect 245 146 246 147
rect 244 146 245 147
rect 243 146 244 147
rect 242 146 243 147
rect 220 146 221 147
rect 219 146 220 147
rect 218 146 219 147
rect 217 146 218 147
rect 216 146 217 147
rect 215 146 216 147
rect 214 146 215 147
rect 213 146 214 147
rect 212 146 213 147
rect 211 146 212 147
rect 210 146 211 147
rect 209 146 210 147
rect 208 146 209 147
rect 207 146 208 147
rect 206 146 207 147
rect 205 146 206 147
rect 204 146 205 147
rect 203 146 204 147
rect 202 146 203 147
rect 201 146 202 147
rect 200 146 201 147
rect 199 146 200 147
rect 198 146 199 147
rect 197 146 198 147
rect 196 146 197 147
rect 195 146 196 147
rect 194 146 195 147
rect 193 146 194 147
rect 192 146 193 147
rect 191 146 192 147
rect 190 146 191 147
rect 189 146 190 147
rect 188 146 189 147
rect 187 146 188 147
rect 186 146 187 147
rect 185 146 186 147
rect 184 146 185 147
rect 183 146 184 147
rect 182 146 183 147
rect 181 146 182 147
rect 180 146 181 147
rect 179 146 180 147
rect 178 146 179 147
rect 177 146 178 147
rect 176 146 177 147
rect 175 146 176 147
rect 174 146 175 147
rect 173 146 174 147
rect 172 146 173 147
rect 171 146 172 147
rect 170 146 171 147
rect 169 146 170 147
rect 168 146 169 147
rect 167 146 168 147
rect 166 146 167 147
rect 165 146 166 147
rect 164 146 165 147
rect 163 146 164 147
rect 162 146 163 147
rect 161 146 162 147
rect 160 146 161 147
rect 159 146 160 147
rect 158 146 159 147
rect 157 146 158 147
rect 156 146 157 147
rect 134 146 135 147
rect 133 146 134 147
rect 132 146 133 147
rect 131 146 132 147
rect 130 146 131 147
rect 129 146 130 147
rect 128 146 129 147
rect 127 146 128 147
rect 126 146 127 147
rect 125 146 126 147
rect 124 146 125 147
rect 123 146 124 147
rect 122 146 123 147
rect 121 146 122 147
rect 120 146 121 147
rect 119 146 120 147
rect 118 146 119 147
rect 117 146 118 147
rect 116 146 117 147
rect 115 146 116 147
rect 114 146 115 147
rect 113 146 114 147
rect 112 146 113 147
rect 111 146 112 147
rect 110 146 111 147
rect 109 146 110 147
rect 108 146 109 147
rect 107 146 108 147
rect 106 146 107 147
rect 105 146 106 147
rect 104 146 105 147
rect 103 146 104 147
rect 102 146 103 147
rect 101 146 102 147
rect 100 146 101 147
rect 99 146 100 147
rect 98 146 99 147
rect 97 146 98 147
rect 96 146 97 147
rect 95 146 96 147
rect 94 146 95 147
rect 93 146 94 147
rect 92 146 93 147
rect 91 146 92 147
rect 90 146 91 147
rect 89 146 90 147
rect 88 146 89 147
rect 87 146 88 147
rect 86 146 87 147
rect 85 146 86 147
rect 84 146 85 147
rect 83 146 84 147
rect 82 146 83 147
rect 81 146 82 147
rect 80 146 81 147
rect 79 146 80 147
rect 78 146 79 147
rect 77 146 78 147
rect 76 146 77 147
rect 75 146 76 147
rect 74 146 75 147
rect 73 146 74 147
rect 72 146 73 147
rect 71 146 72 147
rect 70 146 71 147
rect 69 146 70 147
rect 68 146 69 147
rect 67 146 68 147
rect 66 146 67 147
rect 65 146 66 147
rect 64 146 65 147
rect 63 146 64 147
rect 62 146 63 147
rect 61 146 62 147
rect 60 146 61 147
rect 59 146 60 147
rect 58 146 59 147
rect 57 146 58 147
rect 56 146 57 147
rect 55 146 56 147
rect 54 146 55 147
rect 53 146 54 147
rect 52 146 53 147
rect 51 146 52 147
rect 50 146 51 147
rect 49 146 50 147
rect 48 146 49 147
rect 47 146 48 147
rect 46 146 47 147
rect 45 146 46 147
rect 44 146 45 147
rect 43 146 44 147
rect 42 146 43 147
rect 41 146 42 147
rect 40 146 41 147
rect 28 146 29 147
rect 27 146 28 147
rect 26 146 27 147
rect 25 146 26 147
rect 24 146 25 147
rect 23 146 24 147
rect 22 146 23 147
rect 21 146 22 147
rect 20 146 21 147
rect 19 146 20 147
rect 18 146 19 147
rect 17 146 18 147
rect 16 146 17 147
rect 15 146 16 147
rect 14 146 15 147
rect 13 146 14 147
rect 480 147 481 148
rect 479 147 480 148
rect 478 147 479 148
rect 477 147 478 148
rect 476 147 477 148
rect 475 147 476 148
rect 474 147 475 148
rect 473 147 474 148
rect 472 147 473 148
rect 471 147 472 148
rect 470 147 471 148
rect 469 147 470 148
rect 468 147 469 148
rect 467 147 468 148
rect 466 147 467 148
rect 465 147 466 148
rect 464 147 465 148
rect 463 147 464 148
rect 462 147 463 148
rect 461 147 462 148
rect 460 147 461 148
rect 397 147 398 148
rect 396 147 397 148
rect 395 147 396 148
rect 318 147 319 148
rect 317 147 318 148
rect 316 147 317 148
rect 315 147 316 148
rect 314 147 315 148
rect 313 147 314 148
rect 312 147 313 148
rect 311 147 312 148
rect 310 147 311 148
rect 309 147 310 148
rect 308 147 309 148
rect 307 147 308 148
rect 306 147 307 148
rect 305 147 306 148
rect 304 147 305 148
rect 303 147 304 148
rect 302 147 303 148
rect 301 147 302 148
rect 300 147 301 148
rect 299 147 300 148
rect 298 147 299 148
rect 297 147 298 148
rect 296 147 297 148
rect 295 147 296 148
rect 294 147 295 148
rect 293 147 294 148
rect 292 147 293 148
rect 291 147 292 148
rect 290 147 291 148
rect 289 147 290 148
rect 288 147 289 148
rect 287 147 288 148
rect 286 147 287 148
rect 285 147 286 148
rect 284 147 285 148
rect 283 147 284 148
rect 282 147 283 148
rect 281 147 282 148
rect 280 147 281 148
rect 279 147 280 148
rect 278 147 279 148
rect 277 147 278 148
rect 276 147 277 148
rect 275 147 276 148
rect 274 147 275 148
rect 273 147 274 148
rect 272 147 273 148
rect 271 147 272 148
rect 270 147 271 148
rect 269 147 270 148
rect 268 147 269 148
rect 267 147 268 148
rect 266 147 267 148
rect 265 147 266 148
rect 264 147 265 148
rect 263 147 264 148
rect 262 147 263 148
rect 261 147 262 148
rect 260 147 261 148
rect 259 147 260 148
rect 258 147 259 148
rect 257 147 258 148
rect 256 147 257 148
rect 255 147 256 148
rect 254 147 255 148
rect 253 147 254 148
rect 252 147 253 148
rect 251 147 252 148
rect 250 147 251 148
rect 249 147 250 148
rect 248 147 249 148
rect 247 147 248 148
rect 246 147 247 148
rect 245 147 246 148
rect 244 147 245 148
rect 243 147 244 148
rect 242 147 243 148
rect 241 147 242 148
rect 220 147 221 148
rect 219 147 220 148
rect 218 147 219 148
rect 217 147 218 148
rect 216 147 217 148
rect 215 147 216 148
rect 214 147 215 148
rect 213 147 214 148
rect 212 147 213 148
rect 211 147 212 148
rect 210 147 211 148
rect 209 147 210 148
rect 208 147 209 148
rect 207 147 208 148
rect 206 147 207 148
rect 205 147 206 148
rect 204 147 205 148
rect 203 147 204 148
rect 202 147 203 148
rect 201 147 202 148
rect 200 147 201 148
rect 199 147 200 148
rect 198 147 199 148
rect 197 147 198 148
rect 196 147 197 148
rect 195 147 196 148
rect 194 147 195 148
rect 193 147 194 148
rect 192 147 193 148
rect 191 147 192 148
rect 190 147 191 148
rect 189 147 190 148
rect 188 147 189 148
rect 187 147 188 148
rect 186 147 187 148
rect 185 147 186 148
rect 184 147 185 148
rect 183 147 184 148
rect 182 147 183 148
rect 181 147 182 148
rect 180 147 181 148
rect 179 147 180 148
rect 178 147 179 148
rect 177 147 178 148
rect 176 147 177 148
rect 175 147 176 148
rect 174 147 175 148
rect 173 147 174 148
rect 172 147 173 148
rect 171 147 172 148
rect 170 147 171 148
rect 169 147 170 148
rect 168 147 169 148
rect 167 147 168 148
rect 166 147 167 148
rect 165 147 166 148
rect 164 147 165 148
rect 163 147 164 148
rect 162 147 163 148
rect 161 147 162 148
rect 160 147 161 148
rect 159 147 160 148
rect 158 147 159 148
rect 157 147 158 148
rect 156 147 157 148
rect 132 147 133 148
rect 131 147 132 148
rect 130 147 131 148
rect 129 147 130 148
rect 128 147 129 148
rect 127 147 128 148
rect 126 147 127 148
rect 125 147 126 148
rect 124 147 125 148
rect 123 147 124 148
rect 122 147 123 148
rect 121 147 122 148
rect 120 147 121 148
rect 119 147 120 148
rect 118 147 119 148
rect 117 147 118 148
rect 116 147 117 148
rect 115 147 116 148
rect 114 147 115 148
rect 113 147 114 148
rect 112 147 113 148
rect 111 147 112 148
rect 110 147 111 148
rect 109 147 110 148
rect 108 147 109 148
rect 107 147 108 148
rect 106 147 107 148
rect 105 147 106 148
rect 104 147 105 148
rect 103 147 104 148
rect 102 147 103 148
rect 101 147 102 148
rect 100 147 101 148
rect 99 147 100 148
rect 98 147 99 148
rect 97 147 98 148
rect 96 147 97 148
rect 95 147 96 148
rect 94 147 95 148
rect 93 147 94 148
rect 92 147 93 148
rect 91 147 92 148
rect 90 147 91 148
rect 89 147 90 148
rect 88 147 89 148
rect 87 147 88 148
rect 86 147 87 148
rect 85 147 86 148
rect 84 147 85 148
rect 83 147 84 148
rect 82 147 83 148
rect 81 147 82 148
rect 80 147 81 148
rect 79 147 80 148
rect 78 147 79 148
rect 77 147 78 148
rect 76 147 77 148
rect 75 147 76 148
rect 74 147 75 148
rect 73 147 74 148
rect 72 147 73 148
rect 71 147 72 148
rect 70 147 71 148
rect 69 147 70 148
rect 68 147 69 148
rect 67 147 68 148
rect 66 147 67 148
rect 65 147 66 148
rect 64 147 65 148
rect 63 147 64 148
rect 62 147 63 148
rect 61 147 62 148
rect 60 147 61 148
rect 59 147 60 148
rect 58 147 59 148
rect 57 147 58 148
rect 56 147 57 148
rect 55 147 56 148
rect 54 147 55 148
rect 53 147 54 148
rect 52 147 53 148
rect 51 147 52 148
rect 50 147 51 148
rect 49 147 50 148
rect 48 147 49 148
rect 47 147 48 148
rect 46 147 47 148
rect 45 147 46 148
rect 44 147 45 148
rect 43 147 44 148
rect 42 147 43 148
rect 41 147 42 148
rect 40 147 41 148
rect 29 147 30 148
rect 28 147 29 148
rect 27 147 28 148
rect 26 147 27 148
rect 25 147 26 148
rect 24 147 25 148
rect 23 147 24 148
rect 22 147 23 148
rect 21 147 22 148
rect 20 147 21 148
rect 19 147 20 148
rect 18 147 19 148
rect 17 147 18 148
rect 16 147 17 148
rect 15 147 16 148
rect 14 147 15 148
rect 13 147 14 148
rect 12 147 13 148
rect 480 148 481 149
rect 479 148 480 149
rect 478 148 479 149
rect 477 148 478 149
rect 476 148 477 149
rect 475 148 476 149
rect 474 148 475 149
rect 473 148 474 149
rect 472 148 473 149
rect 471 148 472 149
rect 470 148 471 149
rect 469 148 470 149
rect 468 148 469 149
rect 467 148 468 149
rect 466 148 467 149
rect 465 148 466 149
rect 464 148 465 149
rect 463 148 464 149
rect 462 148 463 149
rect 461 148 462 149
rect 460 148 461 149
rect 397 148 398 149
rect 396 148 397 149
rect 395 148 396 149
rect 319 148 320 149
rect 318 148 319 149
rect 317 148 318 149
rect 316 148 317 149
rect 315 148 316 149
rect 314 148 315 149
rect 313 148 314 149
rect 312 148 313 149
rect 311 148 312 149
rect 310 148 311 149
rect 309 148 310 149
rect 308 148 309 149
rect 307 148 308 149
rect 306 148 307 149
rect 305 148 306 149
rect 304 148 305 149
rect 303 148 304 149
rect 302 148 303 149
rect 301 148 302 149
rect 300 148 301 149
rect 299 148 300 149
rect 298 148 299 149
rect 297 148 298 149
rect 296 148 297 149
rect 295 148 296 149
rect 294 148 295 149
rect 293 148 294 149
rect 292 148 293 149
rect 291 148 292 149
rect 290 148 291 149
rect 289 148 290 149
rect 288 148 289 149
rect 287 148 288 149
rect 286 148 287 149
rect 285 148 286 149
rect 284 148 285 149
rect 283 148 284 149
rect 282 148 283 149
rect 281 148 282 149
rect 280 148 281 149
rect 279 148 280 149
rect 278 148 279 149
rect 277 148 278 149
rect 276 148 277 149
rect 275 148 276 149
rect 274 148 275 149
rect 273 148 274 149
rect 272 148 273 149
rect 271 148 272 149
rect 270 148 271 149
rect 269 148 270 149
rect 268 148 269 149
rect 267 148 268 149
rect 266 148 267 149
rect 265 148 266 149
rect 264 148 265 149
rect 263 148 264 149
rect 262 148 263 149
rect 261 148 262 149
rect 260 148 261 149
rect 259 148 260 149
rect 258 148 259 149
rect 257 148 258 149
rect 256 148 257 149
rect 255 148 256 149
rect 254 148 255 149
rect 253 148 254 149
rect 252 148 253 149
rect 251 148 252 149
rect 250 148 251 149
rect 249 148 250 149
rect 248 148 249 149
rect 247 148 248 149
rect 246 148 247 149
rect 245 148 246 149
rect 244 148 245 149
rect 243 148 244 149
rect 242 148 243 149
rect 241 148 242 149
rect 240 148 241 149
rect 219 148 220 149
rect 218 148 219 149
rect 217 148 218 149
rect 216 148 217 149
rect 215 148 216 149
rect 214 148 215 149
rect 213 148 214 149
rect 212 148 213 149
rect 211 148 212 149
rect 210 148 211 149
rect 209 148 210 149
rect 208 148 209 149
rect 207 148 208 149
rect 206 148 207 149
rect 205 148 206 149
rect 204 148 205 149
rect 203 148 204 149
rect 202 148 203 149
rect 201 148 202 149
rect 200 148 201 149
rect 199 148 200 149
rect 198 148 199 149
rect 197 148 198 149
rect 196 148 197 149
rect 195 148 196 149
rect 194 148 195 149
rect 193 148 194 149
rect 192 148 193 149
rect 191 148 192 149
rect 190 148 191 149
rect 189 148 190 149
rect 188 148 189 149
rect 187 148 188 149
rect 186 148 187 149
rect 185 148 186 149
rect 184 148 185 149
rect 183 148 184 149
rect 182 148 183 149
rect 181 148 182 149
rect 180 148 181 149
rect 179 148 180 149
rect 178 148 179 149
rect 177 148 178 149
rect 176 148 177 149
rect 175 148 176 149
rect 174 148 175 149
rect 173 148 174 149
rect 172 148 173 149
rect 171 148 172 149
rect 170 148 171 149
rect 169 148 170 149
rect 168 148 169 149
rect 167 148 168 149
rect 166 148 167 149
rect 165 148 166 149
rect 164 148 165 149
rect 163 148 164 149
rect 162 148 163 149
rect 161 148 162 149
rect 160 148 161 149
rect 159 148 160 149
rect 158 148 159 149
rect 157 148 158 149
rect 156 148 157 149
rect 155 148 156 149
rect 131 148 132 149
rect 130 148 131 149
rect 129 148 130 149
rect 128 148 129 149
rect 127 148 128 149
rect 126 148 127 149
rect 125 148 126 149
rect 124 148 125 149
rect 123 148 124 149
rect 122 148 123 149
rect 121 148 122 149
rect 120 148 121 149
rect 119 148 120 149
rect 118 148 119 149
rect 117 148 118 149
rect 116 148 117 149
rect 115 148 116 149
rect 114 148 115 149
rect 113 148 114 149
rect 112 148 113 149
rect 111 148 112 149
rect 110 148 111 149
rect 109 148 110 149
rect 108 148 109 149
rect 107 148 108 149
rect 106 148 107 149
rect 105 148 106 149
rect 104 148 105 149
rect 103 148 104 149
rect 102 148 103 149
rect 101 148 102 149
rect 100 148 101 149
rect 99 148 100 149
rect 98 148 99 149
rect 97 148 98 149
rect 96 148 97 149
rect 95 148 96 149
rect 94 148 95 149
rect 93 148 94 149
rect 92 148 93 149
rect 91 148 92 149
rect 90 148 91 149
rect 89 148 90 149
rect 88 148 89 149
rect 87 148 88 149
rect 86 148 87 149
rect 85 148 86 149
rect 84 148 85 149
rect 83 148 84 149
rect 82 148 83 149
rect 81 148 82 149
rect 80 148 81 149
rect 79 148 80 149
rect 78 148 79 149
rect 77 148 78 149
rect 76 148 77 149
rect 75 148 76 149
rect 74 148 75 149
rect 73 148 74 149
rect 72 148 73 149
rect 71 148 72 149
rect 70 148 71 149
rect 69 148 70 149
rect 68 148 69 149
rect 67 148 68 149
rect 66 148 67 149
rect 65 148 66 149
rect 64 148 65 149
rect 63 148 64 149
rect 62 148 63 149
rect 61 148 62 149
rect 60 148 61 149
rect 59 148 60 149
rect 58 148 59 149
rect 57 148 58 149
rect 56 148 57 149
rect 55 148 56 149
rect 54 148 55 149
rect 53 148 54 149
rect 52 148 53 149
rect 51 148 52 149
rect 50 148 51 149
rect 49 148 50 149
rect 48 148 49 149
rect 47 148 48 149
rect 46 148 47 149
rect 45 148 46 149
rect 44 148 45 149
rect 43 148 44 149
rect 42 148 43 149
rect 41 148 42 149
rect 40 148 41 149
rect 29 148 30 149
rect 28 148 29 149
rect 27 148 28 149
rect 26 148 27 149
rect 25 148 26 149
rect 24 148 25 149
rect 23 148 24 149
rect 22 148 23 149
rect 21 148 22 149
rect 20 148 21 149
rect 19 148 20 149
rect 18 148 19 149
rect 17 148 18 149
rect 16 148 17 149
rect 15 148 16 149
rect 14 148 15 149
rect 13 148 14 149
rect 12 148 13 149
rect 11 148 12 149
rect 480 149 481 150
rect 479 149 480 150
rect 478 149 479 150
rect 477 149 478 150
rect 476 149 477 150
rect 475 149 476 150
rect 474 149 475 150
rect 473 149 474 150
rect 472 149 473 150
rect 471 149 472 150
rect 470 149 471 150
rect 469 149 470 150
rect 468 149 469 150
rect 467 149 468 150
rect 466 149 467 150
rect 465 149 466 150
rect 464 149 465 150
rect 463 149 464 150
rect 462 149 463 150
rect 461 149 462 150
rect 460 149 461 150
rect 397 149 398 150
rect 396 149 397 150
rect 395 149 396 150
rect 319 149 320 150
rect 318 149 319 150
rect 317 149 318 150
rect 316 149 317 150
rect 315 149 316 150
rect 314 149 315 150
rect 313 149 314 150
rect 312 149 313 150
rect 311 149 312 150
rect 310 149 311 150
rect 309 149 310 150
rect 308 149 309 150
rect 307 149 308 150
rect 306 149 307 150
rect 305 149 306 150
rect 304 149 305 150
rect 303 149 304 150
rect 302 149 303 150
rect 301 149 302 150
rect 300 149 301 150
rect 299 149 300 150
rect 298 149 299 150
rect 297 149 298 150
rect 296 149 297 150
rect 295 149 296 150
rect 294 149 295 150
rect 293 149 294 150
rect 292 149 293 150
rect 291 149 292 150
rect 290 149 291 150
rect 289 149 290 150
rect 288 149 289 150
rect 287 149 288 150
rect 286 149 287 150
rect 285 149 286 150
rect 284 149 285 150
rect 283 149 284 150
rect 282 149 283 150
rect 281 149 282 150
rect 280 149 281 150
rect 279 149 280 150
rect 278 149 279 150
rect 277 149 278 150
rect 276 149 277 150
rect 275 149 276 150
rect 274 149 275 150
rect 273 149 274 150
rect 272 149 273 150
rect 271 149 272 150
rect 270 149 271 150
rect 269 149 270 150
rect 268 149 269 150
rect 267 149 268 150
rect 266 149 267 150
rect 265 149 266 150
rect 264 149 265 150
rect 263 149 264 150
rect 262 149 263 150
rect 261 149 262 150
rect 260 149 261 150
rect 259 149 260 150
rect 258 149 259 150
rect 257 149 258 150
rect 256 149 257 150
rect 255 149 256 150
rect 254 149 255 150
rect 253 149 254 150
rect 252 149 253 150
rect 251 149 252 150
rect 250 149 251 150
rect 249 149 250 150
rect 248 149 249 150
rect 247 149 248 150
rect 246 149 247 150
rect 245 149 246 150
rect 244 149 245 150
rect 243 149 244 150
rect 242 149 243 150
rect 241 149 242 150
rect 240 149 241 150
rect 219 149 220 150
rect 218 149 219 150
rect 217 149 218 150
rect 216 149 217 150
rect 215 149 216 150
rect 214 149 215 150
rect 213 149 214 150
rect 212 149 213 150
rect 211 149 212 150
rect 210 149 211 150
rect 209 149 210 150
rect 208 149 209 150
rect 207 149 208 150
rect 206 149 207 150
rect 205 149 206 150
rect 204 149 205 150
rect 203 149 204 150
rect 202 149 203 150
rect 201 149 202 150
rect 200 149 201 150
rect 199 149 200 150
rect 198 149 199 150
rect 197 149 198 150
rect 196 149 197 150
rect 195 149 196 150
rect 194 149 195 150
rect 193 149 194 150
rect 192 149 193 150
rect 191 149 192 150
rect 190 149 191 150
rect 189 149 190 150
rect 188 149 189 150
rect 187 149 188 150
rect 186 149 187 150
rect 185 149 186 150
rect 184 149 185 150
rect 183 149 184 150
rect 182 149 183 150
rect 181 149 182 150
rect 180 149 181 150
rect 179 149 180 150
rect 178 149 179 150
rect 177 149 178 150
rect 176 149 177 150
rect 175 149 176 150
rect 174 149 175 150
rect 173 149 174 150
rect 172 149 173 150
rect 171 149 172 150
rect 170 149 171 150
rect 169 149 170 150
rect 168 149 169 150
rect 167 149 168 150
rect 166 149 167 150
rect 165 149 166 150
rect 164 149 165 150
rect 163 149 164 150
rect 162 149 163 150
rect 161 149 162 150
rect 160 149 161 150
rect 159 149 160 150
rect 158 149 159 150
rect 157 149 158 150
rect 156 149 157 150
rect 155 149 156 150
rect 129 149 130 150
rect 128 149 129 150
rect 127 149 128 150
rect 126 149 127 150
rect 125 149 126 150
rect 124 149 125 150
rect 123 149 124 150
rect 122 149 123 150
rect 121 149 122 150
rect 120 149 121 150
rect 119 149 120 150
rect 118 149 119 150
rect 117 149 118 150
rect 116 149 117 150
rect 115 149 116 150
rect 114 149 115 150
rect 113 149 114 150
rect 112 149 113 150
rect 111 149 112 150
rect 110 149 111 150
rect 109 149 110 150
rect 108 149 109 150
rect 107 149 108 150
rect 106 149 107 150
rect 105 149 106 150
rect 104 149 105 150
rect 103 149 104 150
rect 102 149 103 150
rect 101 149 102 150
rect 100 149 101 150
rect 99 149 100 150
rect 98 149 99 150
rect 97 149 98 150
rect 96 149 97 150
rect 95 149 96 150
rect 94 149 95 150
rect 93 149 94 150
rect 92 149 93 150
rect 91 149 92 150
rect 90 149 91 150
rect 89 149 90 150
rect 88 149 89 150
rect 87 149 88 150
rect 86 149 87 150
rect 85 149 86 150
rect 84 149 85 150
rect 83 149 84 150
rect 82 149 83 150
rect 81 149 82 150
rect 80 149 81 150
rect 79 149 80 150
rect 78 149 79 150
rect 77 149 78 150
rect 76 149 77 150
rect 75 149 76 150
rect 74 149 75 150
rect 73 149 74 150
rect 72 149 73 150
rect 71 149 72 150
rect 70 149 71 150
rect 69 149 70 150
rect 68 149 69 150
rect 67 149 68 150
rect 66 149 67 150
rect 65 149 66 150
rect 64 149 65 150
rect 63 149 64 150
rect 62 149 63 150
rect 61 149 62 150
rect 60 149 61 150
rect 59 149 60 150
rect 58 149 59 150
rect 57 149 58 150
rect 56 149 57 150
rect 55 149 56 150
rect 54 149 55 150
rect 53 149 54 150
rect 52 149 53 150
rect 51 149 52 150
rect 50 149 51 150
rect 49 149 50 150
rect 48 149 49 150
rect 47 149 48 150
rect 46 149 47 150
rect 45 149 46 150
rect 44 149 45 150
rect 43 149 44 150
rect 42 149 43 150
rect 41 149 42 150
rect 40 149 41 150
rect 39 149 40 150
rect 29 149 30 150
rect 28 149 29 150
rect 27 149 28 150
rect 26 149 27 150
rect 25 149 26 150
rect 24 149 25 150
rect 23 149 24 150
rect 22 149 23 150
rect 21 149 22 150
rect 20 149 21 150
rect 19 149 20 150
rect 18 149 19 150
rect 17 149 18 150
rect 16 149 17 150
rect 15 149 16 150
rect 14 149 15 150
rect 13 149 14 150
rect 12 149 13 150
rect 11 149 12 150
rect 480 150 481 151
rect 460 150 461 151
rect 320 150 321 151
rect 319 150 320 151
rect 318 150 319 151
rect 317 150 318 151
rect 316 150 317 151
rect 315 150 316 151
rect 314 150 315 151
rect 313 150 314 151
rect 312 150 313 151
rect 311 150 312 151
rect 310 150 311 151
rect 309 150 310 151
rect 308 150 309 151
rect 307 150 308 151
rect 306 150 307 151
rect 305 150 306 151
rect 304 150 305 151
rect 303 150 304 151
rect 302 150 303 151
rect 301 150 302 151
rect 300 150 301 151
rect 299 150 300 151
rect 298 150 299 151
rect 297 150 298 151
rect 296 150 297 151
rect 295 150 296 151
rect 294 150 295 151
rect 293 150 294 151
rect 292 150 293 151
rect 291 150 292 151
rect 290 150 291 151
rect 289 150 290 151
rect 288 150 289 151
rect 287 150 288 151
rect 286 150 287 151
rect 285 150 286 151
rect 284 150 285 151
rect 283 150 284 151
rect 282 150 283 151
rect 281 150 282 151
rect 280 150 281 151
rect 279 150 280 151
rect 278 150 279 151
rect 277 150 278 151
rect 276 150 277 151
rect 275 150 276 151
rect 274 150 275 151
rect 273 150 274 151
rect 272 150 273 151
rect 271 150 272 151
rect 270 150 271 151
rect 269 150 270 151
rect 268 150 269 151
rect 267 150 268 151
rect 266 150 267 151
rect 265 150 266 151
rect 264 150 265 151
rect 263 150 264 151
rect 262 150 263 151
rect 261 150 262 151
rect 260 150 261 151
rect 259 150 260 151
rect 258 150 259 151
rect 257 150 258 151
rect 256 150 257 151
rect 255 150 256 151
rect 254 150 255 151
rect 253 150 254 151
rect 252 150 253 151
rect 251 150 252 151
rect 250 150 251 151
rect 249 150 250 151
rect 248 150 249 151
rect 247 150 248 151
rect 246 150 247 151
rect 245 150 246 151
rect 244 150 245 151
rect 243 150 244 151
rect 242 150 243 151
rect 241 150 242 151
rect 240 150 241 151
rect 239 150 240 151
rect 218 150 219 151
rect 217 150 218 151
rect 216 150 217 151
rect 215 150 216 151
rect 214 150 215 151
rect 213 150 214 151
rect 212 150 213 151
rect 211 150 212 151
rect 210 150 211 151
rect 209 150 210 151
rect 208 150 209 151
rect 207 150 208 151
rect 206 150 207 151
rect 205 150 206 151
rect 204 150 205 151
rect 203 150 204 151
rect 202 150 203 151
rect 201 150 202 151
rect 200 150 201 151
rect 199 150 200 151
rect 198 150 199 151
rect 197 150 198 151
rect 196 150 197 151
rect 195 150 196 151
rect 194 150 195 151
rect 193 150 194 151
rect 192 150 193 151
rect 191 150 192 151
rect 190 150 191 151
rect 189 150 190 151
rect 188 150 189 151
rect 187 150 188 151
rect 186 150 187 151
rect 185 150 186 151
rect 184 150 185 151
rect 183 150 184 151
rect 182 150 183 151
rect 181 150 182 151
rect 180 150 181 151
rect 179 150 180 151
rect 178 150 179 151
rect 177 150 178 151
rect 176 150 177 151
rect 175 150 176 151
rect 174 150 175 151
rect 173 150 174 151
rect 172 150 173 151
rect 171 150 172 151
rect 170 150 171 151
rect 169 150 170 151
rect 168 150 169 151
rect 167 150 168 151
rect 166 150 167 151
rect 165 150 166 151
rect 164 150 165 151
rect 163 150 164 151
rect 162 150 163 151
rect 161 150 162 151
rect 160 150 161 151
rect 159 150 160 151
rect 158 150 159 151
rect 157 150 158 151
rect 156 150 157 151
rect 155 150 156 151
rect 154 150 155 151
rect 128 150 129 151
rect 127 150 128 151
rect 126 150 127 151
rect 125 150 126 151
rect 124 150 125 151
rect 123 150 124 151
rect 122 150 123 151
rect 121 150 122 151
rect 120 150 121 151
rect 119 150 120 151
rect 118 150 119 151
rect 117 150 118 151
rect 116 150 117 151
rect 115 150 116 151
rect 114 150 115 151
rect 113 150 114 151
rect 112 150 113 151
rect 111 150 112 151
rect 110 150 111 151
rect 109 150 110 151
rect 108 150 109 151
rect 107 150 108 151
rect 106 150 107 151
rect 105 150 106 151
rect 104 150 105 151
rect 103 150 104 151
rect 102 150 103 151
rect 101 150 102 151
rect 100 150 101 151
rect 99 150 100 151
rect 98 150 99 151
rect 97 150 98 151
rect 96 150 97 151
rect 95 150 96 151
rect 94 150 95 151
rect 93 150 94 151
rect 92 150 93 151
rect 91 150 92 151
rect 90 150 91 151
rect 89 150 90 151
rect 88 150 89 151
rect 87 150 88 151
rect 86 150 87 151
rect 85 150 86 151
rect 84 150 85 151
rect 83 150 84 151
rect 82 150 83 151
rect 81 150 82 151
rect 80 150 81 151
rect 79 150 80 151
rect 78 150 79 151
rect 77 150 78 151
rect 76 150 77 151
rect 75 150 76 151
rect 74 150 75 151
rect 73 150 74 151
rect 72 150 73 151
rect 71 150 72 151
rect 70 150 71 151
rect 69 150 70 151
rect 68 150 69 151
rect 67 150 68 151
rect 66 150 67 151
rect 65 150 66 151
rect 64 150 65 151
rect 63 150 64 151
rect 62 150 63 151
rect 61 150 62 151
rect 60 150 61 151
rect 59 150 60 151
rect 58 150 59 151
rect 57 150 58 151
rect 56 150 57 151
rect 55 150 56 151
rect 54 150 55 151
rect 53 150 54 151
rect 52 150 53 151
rect 51 150 52 151
rect 50 150 51 151
rect 49 150 50 151
rect 48 150 49 151
rect 47 150 48 151
rect 46 150 47 151
rect 45 150 46 151
rect 44 150 45 151
rect 43 150 44 151
rect 42 150 43 151
rect 41 150 42 151
rect 40 150 41 151
rect 39 150 40 151
rect 29 150 30 151
rect 28 150 29 151
rect 27 150 28 151
rect 26 150 27 151
rect 25 150 26 151
rect 24 150 25 151
rect 23 150 24 151
rect 22 150 23 151
rect 21 150 22 151
rect 20 150 21 151
rect 19 150 20 151
rect 18 150 19 151
rect 17 150 18 151
rect 16 150 17 151
rect 15 150 16 151
rect 14 150 15 151
rect 13 150 14 151
rect 12 150 13 151
rect 11 150 12 151
rect 10 150 11 151
rect 480 151 481 152
rect 460 151 461 152
rect 321 151 322 152
rect 320 151 321 152
rect 319 151 320 152
rect 318 151 319 152
rect 317 151 318 152
rect 316 151 317 152
rect 315 151 316 152
rect 314 151 315 152
rect 313 151 314 152
rect 312 151 313 152
rect 311 151 312 152
rect 310 151 311 152
rect 309 151 310 152
rect 308 151 309 152
rect 307 151 308 152
rect 306 151 307 152
rect 305 151 306 152
rect 304 151 305 152
rect 303 151 304 152
rect 302 151 303 152
rect 301 151 302 152
rect 300 151 301 152
rect 299 151 300 152
rect 298 151 299 152
rect 297 151 298 152
rect 296 151 297 152
rect 295 151 296 152
rect 294 151 295 152
rect 293 151 294 152
rect 292 151 293 152
rect 291 151 292 152
rect 290 151 291 152
rect 289 151 290 152
rect 288 151 289 152
rect 287 151 288 152
rect 286 151 287 152
rect 285 151 286 152
rect 284 151 285 152
rect 283 151 284 152
rect 282 151 283 152
rect 281 151 282 152
rect 280 151 281 152
rect 279 151 280 152
rect 278 151 279 152
rect 277 151 278 152
rect 276 151 277 152
rect 275 151 276 152
rect 274 151 275 152
rect 273 151 274 152
rect 272 151 273 152
rect 271 151 272 152
rect 270 151 271 152
rect 269 151 270 152
rect 268 151 269 152
rect 267 151 268 152
rect 266 151 267 152
rect 265 151 266 152
rect 264 151 265 152
rect 263 151 264 152
rect 262 151 263 152
rect 261 151 262 152
rect 260 151 261 152
rect 259 151 260 152
rect 258 151 259 152
rect 257 151 258 152
rect 256 151 257 152
rect 255 151 256 152
rect 254 151 255 152
rect 253 151 254 152
rect 252 151 253 152
rect 251 151 252 152
rect 250 151 251 152
rect 249 151 250 152
rect 248 151 249 152
rect 247 151 248 152
rect 246 151 247 152
rect 245 151 246 152
rect 244 151 245 152
rect 243 151 244 152
rect 242 151 243 152
rect 241 151 242 152
rect 240 151 241 152
rect 239 151 240 152
rect 238 151 239 152
rect 218 151 219 152
rect 217 151 218 152
rect 216 151 217 152
rect 215 151 216 152
rect 214 151 215 152
rect 213 151 214 152
rect 212 151 213 152
rect 211 151 212 152
rect 210 151 211 152
rect 209 151 210 152
rect 208 151 209 152
rect 207 151 208 152
rect 206 151 207 152
rect 205 151 206 152
rect 204 151 205 152
rect 203 151 204 152
rect 202 151 203 152
rect 201 151 202 152
rect 200 151 201 152
rect 199 151 200 152
rect 198 151 199 152
rect 197 151 198 152
rect 196 151 197 152
rect 195 151 196 152
rect 194 151 195 152
rect 193 151 194 152
rect 192 151 193 152
rect 191 151 192 152
rect 190 151 191 152
rect 189 151 190 152
rect 188 151 189 152
rect 187 151 188 152
rect 186 151 187 152
rect 185 151 186 152
rect 184 151 185 152
rect 183 151 184 152
rect 182 151 183 152
rect 181 151 182 152
rect 180 151 181 152
rect 179 151 180 152
rect 178 151 179 152
rect 177 151 178 152
rect 176 151 177 152
rect 175 151 176 152
rect 174 151 175 152
rect 173 151 174 152
rect 172 151 173 152
rect 171 151 172 152
rect 170 151 171 152
rect 169 151 170 152
rect 168 151 169 152
rect 167 151 168 152
rect 166 151 167 152
rect 165 151 166 152
rect 164 151 165 152
rect 163 151 164 152
rect 162 151 163 152
rect 161 151 162 152
rect 160 151 161 152
rect 159 151 160 152
rect 158 151 159 152
rect 157 151 158 152
rect 156 151 157 152
rect 155 151 156 152
rect 154 151 155 152
rect 153 151 154 152
rect 126 151 127 152
rect 125 151 126 152
rect 124 151 125 152
rect 123 151 124 152
rect 122 151 123 152
rect 121 151 122 152
rect 120 151 121 152
rect 119 151 120 152
rect 118 151 119 152
rect 117 151 118 152
rect 116 151 117 152
rect 115 151 116 152
rect 114 151 115 152
rect 113 151 114 152
rect 112 151 113 152
rect 111 151 112 152
rect 110 151 111 152
rect 109 151 110 152
rect 108 151 109 152
rect 107 151 108 152
rect 106 151 107 152
rect 105 151 106 152
rect 104 151 105 152
rect 103 151 104 152
rect 102 151 103 152
rect 101 151 102 152
rect 100 151 101 152
rect 99 151 100 152
rect 98 151 99 152
rect 97 151 98 152
rect 96 151 97 152
rect 95 151 96 152
rect 94 151 95 152
rect 93 151 94 152
rect 92 151 93 152
rect 91 151 92 152
rect 90 151 91 152
rect 89 151 90 152
rect 88 151 89 152
rect 87 151 88 152
rect 86 151 87 152
rect 85 151 86 152
rect 84 151 85 152
rect 83 151 84 152
rect 82 151 83 152
rect 81 151 82 152
rect 80 151 81 152
rect 79 151 80 152
rect 78 151 79 152
rect 77 151 78 152
rect 76 151 77 152
rect 75 151 76 152
rect 74 151 75 152
rect 73 151 74 152
rect 72 151 73 152
rect 71 151 72 152
rect 70 151 71 152
rect 69 151 70 152
rect 68 151 69 152
rect 67 151 68 152
rect 66 151 67 152
rect 65 151 66 152
rect 64 151 65 152
rect 63 151 64 152
rect 62 151 63 152
rect 61 151 62 152
rect 60 151 61 152
rect 59 151 60 152
rect 58 151 59 152
rect 57 151 58 152
rect 56 151 57 152
rect 55 151 56 152
rect 54 151 55 152
rect 53 151 54 152
rect 52 151 53 152
rect 51 151 52 152
rect 50 151 51 152
rect 49 151 50 152
rect 48 151 49 152
rect 47 151 48 152
rect 46 151 47 152
rect 45 151 46 152
rect 44 151 45 152
rect 43 151 44 152
rect 42 151 43 152
rect 41 151 42 152
rect 40 151 41 152
rect 39 151 40 152
rect 38 151 39 152
rect 29 151 30 152
rect 28 151 29 152
rect 27 151 28 152
rect 26 151 27 152
rect 25 151 26 152
rect 24 151 25 152
rect 23 151 24 152
rect 22 151 23 152
rect 21 151 22 152
rect 20 151 21 152
rect 19 151 20 152
rect 18 151 19 152
rect 17 151 18 152
rect 16 151 17 152
rect 15 151 16 152
rect 14 151 15 152
rect 13 151 14 152
rect 12 151 13 152
rect 11 151 12 152
rect 10 151 11 152
rect 9 151 10 152
rect 322 152 323 153
rect 321 152 322 153
rect 320 152 321 153
rect 319 152 320 153
rect 318 152 319 153
rect 317 152 318 153
rect 316 152 317 153
rect 315 152 316 153
rect 314 152 315 153
rect 313 152 314 153
rect 312 152 313 153
rect 311 152 312 153
rect 310 152 311 153
rect 309 152 310 153
rect 308 152 309 153
rect 307 152 308 153
rect 306 152 307 153
rect 305 152 306 153
rect 304 152 305 153
rect 303 152 304 153
rect 302 152 303 153
rect 301 152 302 153
rect 300 152 301 153
rect 299 152 300 153
rect 298 152 299 153
rect 297 152 298 153
rect 296 152 297 153
rect 295 152 296 153
rect 294 152 295 153
rect 293 152 294 153
rect 292 152 293 153
rect 291 152 292 153
rect 290 152 291 153
rect 289 152 290 153
rect 288 152 289 153
rect 287 152 288 153
rect 286 152 287 153
rect 285 152 286 153
rect 284 152 285 153
rect 283 152 284 153
rect 282 152 283 153
rect 281 152 282 153
rect 280 152 281 153
rect 279 152 280 153
rect 278 152 279 153
rect 277 152 278 153
rect 276 152 277 153
rect 275 152 276 153
rect 274 152 275 153
rect 273 152 274 153
rect 272 152 273 153
rect 271 152 272 153
rect 270 152 271 153
rect 269 152 270 153
rect 268 152 269 153
rect 267 152 268 153
rect 266 152 267 153
rect 265 152 266 153
rect 264 152 265 153
rect 263 152 264 153
rect 262 152 263 153
rect 261 152 262 153
rect 260 152 261 153
rect 259 152 260 153
rect 258 152 259 153
rect 257 152 258 153
rect 256 152 257 153
rect 255 152 256 153
rect 254 152 255 153
rect 253 152 254 153
rect 252 152 253 153
rect 251 152 252 153
rect 250 152 251 153
rect 249 152 250 153
rect 248 152 249 153
rect 247 152 248 153
rect 246 152 247 153
rect 245 152 246 153
rect 244 152 245 153
rect 243 152 244 153
rect 242 152 243 153
rect 241 152 242 153
rect 240 152 241 153
rect 239 152 240 153
rect 238 152 239 153
rect 218 152 219 153
rect 217 152 218 153
rect 216 152 217 153
rect 215 152 216 153
rect 214 152 215 153
rect 213 152 214 153
rect 212 152 213 153
rect 211 152 212 153
rect 210 152 211 153
rect 209 152 210 153
rect 208 152 209 153
rect 207 152 208 153
rect 206 152 207 153
rect 205 152 206 153
rect 204 152 205 153
rect 203 152 204 153
rect 202 152 203 153
rect 201 152 202 153
rect 200 152 201 153
rect 199 152 200 153
rect 198 152 199 153
rect 197 152 198 153
rect 196 152 197 153
rect 195 152 196 153
rect 194 152 195 153
rect 193 152 194 153
rect 192 152 193 153
rect 191 152 192 153
rect 190 152 191 153
rect 189 152 190 153
rect 188 152 189 153
rect 187 152 188 153
rect 186 152 187 153
rect 185 152 186 153
rect 184 152 185 153
rect 183 152 184 153
rect 182 152 183 153
rect 181 152 182 153
rect 180 152 181 153
rect 179 152 180 153
rect 178 152 179 153
rect 177 152 178 153
rect 176 152 177 153
rect 175 152 176 153
rect 174 152 175 153
rect 173 152 174 153
rect 172 152 173 153
rect 171 152 172 153
rect 170 152 171 153
rect 169 152 170 153
rect 168 152 169 153
rect 167 152 168 153
rect 166 152 167 153
rect 165 152 166 153
rect 164 152 165 153
rect 163 152 164 153
rect 162 152 163 153
rect 161 152 162 153
rect 160 152 161 153
rect 159 152 160 153
rect 158 152 159 153
rect 157 152 158 153
rect 156 152 157 153
rect 155 152 156 153
rect 154 152 155 153
rect 153 152 154 153
rect 152 152 153 153
rect 124 152 125 153
rect 123 152 124 153
rect 122 152 123 153
rect 121 152 122 153
rect 120 152 121 153
rect 119 152 120 153
rect 118 152 119 153
rect 117 152 118 153
rect 116 152 117 153
rect 115 152 116 153
rect 114 152 115 153
rect 113 152 114 153
rect 112 152 113 153
rect 111 152 112 153
rect 110 152 111 153
rect 109 152 110 153
rect 108 152 109 153
rect 107 152 108 153
rect 106 152 107 153
rect 105 152 106 153
rect 104 152 105 153
rect 103 152 104 153
rect 102 152 103 153
rect 101 152 102 153
rect 100 152 101 153
rect 99 152 100 153
rect 98 152 99 153
rect 97 152 98 153
rect 96 152 97 153
rect 95 152 96 153
rect 94 152 95 153
rect 93 152 94 153
rect 92 152 93 153
rect 91 152 92 153
rect 90 152 91 153
rect 89 152 90 153
rect 88 152 89 153
rect 87 152 88 153
rect 86 152 87 153
rect 85 152 86 153
rect 84 152 85 153
rect 83 152 84 153
rect 82 152 83 153
rect 81 152 82 153
rect 80 152 81 153
rect 79 152 80 153
rect 78 152 79 153
rect 77 152 78 153
rect 76 152 77 153
rect 75 152 76 153
rect 74 152 75 153
rect 73 152 74 153
rect 72 152 73 153
rect 71 152 72 153
rect 70 152 71 153
rect 69 152 70 153
rect 68 152 69 153
rect 67 152 68 153
rect 66 152 67 153
rect 65 152 66 153
rect 64 152 65 153
rect 63 152 64 153
rect 62 152 63 153
rect 61 152 62 153
rect 60 152 61 153
rect 59 152 60 153
rect 58 152 59 153
rect 57 152 58 153
rect 56 152 57 153
rect 55 152 56 153
rect 54 152 55 153
rect 53 152 54 153
rect 52 152 53 153
rect 51 152 52 153
rect 50 152 51 153
rect 49 152 50 153
rect 48 152 49 153
rect 47 152 48 153
rect 46 152 47 153
rect 45 152 46 153
rect 44 152 45 153
rect 43 152 44 153
rect 42 152 43 153
rect 41 152 42 153
rect 40 152 41 153
rect 39 152 40 153
rect 38 152 39 153
rect 28 152 29 153
rect 27 152 28 153
rect 26 152 27 153
rect 25 152 26 153
rect 24 152 25 153
rect 23 152 24 153
rect 22 152 23 153
rect 21 152 22 153
rect 20 152 21 153
rect 19 152 20 153
rect 18 152 19 153
rect 17 152 18 153
rect 16 152 17 153
rect 15 152 16 153
rect 14 152 15 153
rect 13 152 14 153
rect 12 152 13 153
rect 11 152 12 153
rect 10 152 11 153
rect 9 152 10 153
rect 323 153 324 154
rect 322 153 323 154
rect 321 153 322 154
rect 320 153 321 154
rect 319 153 320 154
rect 318 153 319 154
rect 317 153 318 154
rect 316 153 317 154
rect 315 153 316 154
rect 314 153 315 154
rect 313 153 314 154
rect 312 153 313 154
rect 311 153 312 154
rect 310 153 311 154
rect 309 153 310 154
rect 308 153 309 154
rect 307 153 308 154
rect 306 153 307 154
rect 305 153 306 154
rect 304 153 305 154
rect 303 153 304 154
rect 302 153 303 154
rect 301 153 302 154
rect 300 153 301 154
rect 299 153 300 154
rect 298 153 299 154
rect 297 153 298 154
rect 296 153 297 154
rect 295 153 296 154
rect 294 153 295 154
rect 293 153 294 154
rect 292 153 293 154
rect 291 153 292 154
rect 290 153 291 154
rect 289 153 290 154
rect 288 153 289 154
rect 287 153 288 154
rect 286 153 287 154
rect 285 153 286 154
rect 284 153 285 154
rect 283 153 284 154
rect 282 153 283 154
rect 281 153 282 154
rect 280 153 281 154
rect 279 153 280 154
rect 278 153 279 154
rect 277 153 278 154
rect 276 153 277 154
rect 275 153 276 154
rect 274 153 275 154
rect 273 153 274 154
rect 272 153 273 154
rect 271 153 272 154
rect 270 153 271 154
rect 269 153 270 154
rect 268 153 269 154
rect 267 153 268 154
rect 266 153 267 154
rect 265 153 266 154
rect 264 153 265 154
rect 263 153 264 154
rect 262 153 263 154
rect 261 153 262 154
rect 260 153 261 154
rect 259 153 260 154
rect 258 153 259 154
rect 257 153 258 154
rect 256 153 257 154
rect 255 153 256 154
rect 254 153 255 154
rect 253 153 254 154
rect 252 153 253 154
rect 251 153 252 154
rect 250 153 251 154
rect 249 153 250 154
rect 248 153 249 154
rect 247 153 248 154
rect 246 153 247 154
rect 245 153 246 154
rect 244 153 245 154
rect 243 153 244 154
rect 242 153 243 154
rect 241 153 242 154
rect 240 153 241 154
rect 239 153 240 154
rect 238 153 239 154
rect 237 153 238 154
rect 217 153 218 154
rect 216 153 217 154
rect 215 153 216 154
rect 214 153 215 154
rect 213 153 214 154
rect 212 153 213 154
rect 211 153 212 154
rect 210 153 211 154
rect 209 153 210 154
rect 208 153 209 154
rect 207 153 208 154
rect 206 153 207 154
rect 205 153 206 154
rect 204 153 205 154
rect 203 153 204 154
rect 202 153 203 154
rect 201 153 202 154
rect 200 153 201 154
rect 199 153 200 154
rect 198 153 199 154
rect 197 153 198 154
rect 196 153 197 154
rect 195 153 196 154
rect 194 153 195 154
rect 193 153 194 154
rect 192 153 193 154
rect 191 153 192 154
rect 190 153 191 154
rect 189 153 190 154
rect 188 153 189 154
rect 187 153 188 154
rect 186 153 187 154
rect 185 153 186 154
rect 184 153 185 154
rect 183 153 184 154
rect 182 153 183 154
rect 181 153 182 154
rect 180 153 181 154
rect 179 153 180 154
rect 178 153 179 154
rect 177 153 178 154
rect 176 153 177 154
rect 175 153 176 154
rect 174 153 175 154
rect 173 153 174 154
rect 172 153 173 154
rect 171 153 172 154
rect 170 153 171 154
rect 169 153 170 154
rect 168 153 169 154
rect 167 153 168 154
rect 166 153 167 154
rect 165 153 166 154
rect 164 153 165 154
rect 163 153 164 154
rect 162 153 163 154
rect 161 153 162 154
rect 160 153 161 154
rect 159 153 160 154
rect 158 153 159 154
rect 157 153 158 154
rect 156 153 157 154
rect 155 153 156 154
rect 154 153 155 154
rect 153 153 154 154
rect 152 153 153 154
rect 123 153 124 154
rect 122 153 123 154
rect 121 153 122 154
rect 120 153 121 154
rect 119 153 120 154
rect 118 153 119 154
rect 117 153 118 154
rect 116 153 117 154
rect 115 153 116 154
rect 114 153 115 154
rect 113 153 114 154
rect 112 153 113 154
rect 111 153 112 154
rect 110 153 111 154
rect 109 153 110 154
rect 108 153 109 154
rect 107 153 108 154
rect 106 153 107 154
rect 105 153 106 154
rect 104 153 105 154
rect 103 153 104 154
rect 102 153 103 154
rect 101 153 102 154
rect 100 153 101 154
rect 99 153 100 154
rect 98 153 99 154
rect 97 153 98 154
rect 96 153 97 154
rect 95 153 96 154
rect 94 153 95 154
rect 93 153 94 154
rect 92 153 93 154
rect 91 153 92 154
rect 90 153 91 154
rect 89 153 90 154
rect 88 153 89 154
rect 87 153 88 154
rect 86 153 87 154
rect 85 153 86 154
rect 84 153 85 154
rect 83 153 84 154
rect 82 153 83 154
rect 81 153 82 154
rect 80 153 81 154
rect 79 153 80 154
rect 78 153 79 154
rect 77 153 78 154
rect 76 153 77 154
rect 75 153 76 154
rect 74 153 75 154
rect 73 153 74 154
rect 72 153 73 154
rect 71 153 72 154
rect 70 153 71 154
rect 69 153 70 154
rect 68 153 69 154
rect 67 153 68 154
rect 66 153 67 154
rect 65 153 66 154
rect 64 153 65 154
rect 63 153 64 154
rect 62 153 63 154
rect 61 153 62 154
rect 60 153 61 154
rect 59 153 60 154
rect 58 153 59 154
rect 57 153 58 154
rect 56 153 57 154
rect 55 153 56 154
rect 54 153 55 154
rect 53 153 54 154
rect 52 153 53 154
rect 51 153 52 154
rect 50 153 51 154
rect 49 153 50 154
rect 48 153 49 154
rect 47 153 48 154
rect 46 153 47 154
rect 45 153 46 154
rect 44 153 45 154
rect 43 153 44 154
rect 42 153 43 154
rect 41 153 42 154
rect 40 153 41 154
rect 39 153 40 154
rect 38 153 39 154
rect 37 153 38 154
rect 28 153 29 154
rect 27 153 28 154
rect 26 153 27 154
rect 25 153 26 154
rect 24 153 25 154
rect 23 153 24 154
rect 22 153 23 154
rect 21 153 22 154
rect 20 153 21 154
rect 19 153 20 154
rect 18 153 19 154
rect 17 153 18 154
rect 16 153 17 154
rect 15 153 16 154
rect 14 153 15 154
rect 13 153 14 154
rect 12 153 13 154
rect 11 153 12 154
rect 10 153 11 154
rect 9 153 10 154
rect 8 153 9 154
rect 396 154 397 155
rect 395 154 396 155
rect 323 154 324 155
rect 322 154 323 155
rect 321 154 322 155
rect 320 154 321 155
rect 319 154 320 155
rect 318 154 319 155
rect 317 154 318 155
rect 316 154 317 155
rect 315 154 316 155
rect 314 154 315 155
rect 313 154 314 155
rect 312 154 313 155
rect 311 154 312 155
rect 310 154 311 155
rect 309 154 310 155
rect 308 154 309 155
rect 307 154 308 155
rect 306 154 307 155
rect 305 154 306 155
rect 304 154 305 155
rect 303 154 304 155
rect 302 154 303 155
rect 301 154 302 155
rect 300 154 301 155
rect 299 154 300 155
rect 298 154 299 155
rect 297 154 298 155
rect 296 154 297 155
rect 295 154 296 155
rect 294 154 295 155
rect 293 154 294 155
rect 292 154 293 155
rect 291 154 292 155
rect 290 154 291 155
rect 289 154 290 155
rect 288 154 289 155
rect 287 154 288 155
rect 286 154 287 155
rect 285 154 286 155
rect 284 154 285 155
rect 283 154 284 155
rect 282 154 283 155
rect 281 154 282 155
rect 280 154 281 155
rect 279 154 280 155
rect 278 154 279 155
rect 277 154 278 155
rect 276 154 277 155
rect 275 154 276 155
rect 274 154 275 155
rect 273 154 274 155
rect 272 154 273 155
rect 271 154 272 155
rect 270 154 271 155
rect 269 154 270 155
rect 268 154 269 155
rect 267 154 268 155
rect 266 154 267 155
rect 265 154 266 155
rect 264 154 265 155
rect 263 154 264 155
rect 262 154 263 155
rect 261 154 262 155
rect 260 154 261 155
rect 259 154 260 155
rect 258 154 259 155
rect 257 154 258 155
rect 256 154 257 155
rect 255 154 256 155
rect 254 154 255 155
rect 253 154 254 155
rect 252 154 253 155
rect 251 154 252 155
rect 250 154 251 155
rect 249 154 250 155
rect 248 154 249 155
rect 247 154 248 155
rect 246 154 247 155
rect 245 154 246 155
rect 244 154 245 155
rect 243 154 244 155
rect 242 154 243 155
rect 241 154 242 155
rect 240 154 241 155
rect 239 154 240 155
rect 238 154 239 155
rect 237 154 238 155
rect 236 154 237 155
rect 217 154 218 155
rect 216 154 217 155
rect 215 154 216 155
rect 214 154 215 155
rect 213 154 214 155
rect 212 154 213 155
rect 211 154 212 155
rect 210 154 211 155
rect 209 154 210 155
rect 208 154 209 155
rect 207 154 208 155
rect 206 154 207 155
rect 205 154 206 155
rect 204 154 205 155
rect 203 154 204 155
rect 202 154 203 155
rect 201 154 202 155
rect 200 154 201 155
rect 199 154 200 155
rect 198 154 199 155
rect 197 154 198 155
rect 196 154 197 155
rect 195 154 196 155
rect 194 154 195 155
rect 193 154 194 155
rect 192 154 193 155
rect 191 154 192 155
rect 190 154 191 155
rect 189 154 190 155
rect 188 154 189 155
rect 187 154 188 155
rect 186 154 187 155
rect 185 154 186 155
rect 184 154 185 155
rect 183 154 184 155
rect 182 154 183 155
rect 181 154 182 155
rect 180 154 181 155
rect 179 154 180 155
rect 178 154 179 155
rect 177 154 178 155
rect 176 154 177 155
rect 175 154 176 155
rect 174 154 175 155
rect 173 154 174 155
rect 172 154 173 155
rect 171 154 172 155
rect 170 154 171 155
rect 169 154 170 155
rect 168 154 169 155
rect 167 154 168 155
rect 166 154 167 155
rect 165 154 166 155
rect 164 154 165 155
rect 163 154 164 155
rect 162 154 163 155
rect 161 154 162 155
rect 160 154 161 155
rect 159 154 160 155
rect 158 154 159 155
rect 157 154 158 155
rect 156 154 157 155
rect 155 154 156 155
rect 154 154 155 155
rect 153 154 154 155
rect 152 154 153 155
rect 151 154 152 155
rect 121 154 122 155
rect 120 154 121 155
rect 119 154 120 155
rect 118 154 119 155
rect 117 154 118 155
rect 116 154 117 155
rect 115 154 116 155
rect 114 154 115 155
rect 113 154 114 155
rect 112 154 113 155
rect 111 154 112 155
rect 110 154 111 155
rect 109 154 110 155
rect 108 154 109 155
rect 107 154 108 155
rect 106 154 107 155
rect 105 154 106 155
rect 104 154 105 155
rect 103 154 104 155
rect 102 154 103 155
rect 101 154 102 155
rect 100 154 101 155
rect 99 154 100 155
rect 98 154 99 155
rect 97 154 98 155
rect 96 154 97 155
rect 95 154 96 155
rect 94 154 95 155
rect 93 154 94 155
rect 92 154 93 155
rect 91 154 92 155
rect 90 154 91 155
rect 89 154 90 155
rect 88 154 89 155
rect 87 154 88 155
rect 86 154 87 155
rect 85 154 86 155
rect 84 154 85 155
rect 83 154 84 155
rect 82 154 83 155
rect 81 154 82 155
rect 80 154 81 155
rect 79 154 80 155
rect 78 154 79 155
rect 77 154 78 155
rect 76 154 77 155
rect 75 154 76 155
rect 74 154 75 155
rect 73 154 74 155
rect 72 154 73 155
rect 71 154 72 155
rect 70 154 71 155
rect 69 154 70 155
rect 68 154 69 155
rect 67 154 68 155
rect 66 154 67 155
rect 65 154 66 155
rect 64 154 65 155
rect 63 154 64 155
rect 62 154 63 155
rect 61 154 62 155
rect 60 154 61 155
rect 59 154 60 155
rect 58 154 59 155
rect 57 154 58 155
rect 56 154 57 155
rect 55 154 56 155
rect 54 154 55 155
rect 53 154 54 155
rect 52 154 53 155
rect 51 154 52 155
rect 50 154 51 155
rect 49 154 50 155
rect 48 154 49 155
rect 47 154 48 155
rect 46 154 47 155
rect 45 154 46 155
rect 44 154 45 155
rect 43 154 44 155
rect 42 154 43 155
rect 41 154 42 155
rect 40 154 41 155
rect 39 154 40 155
rect 38 154 39 155
rect 37 154 38 155
rect 28 154 29 155
rect 27 154 28 155
rect 26 154 27 155
rect 25 154 26 155
rect 24 154 25 155
rect 23 154 24 155
rect 22 154 23 155
rect 21 154 22 155
rect 20 154 21 155
rect 19 154 20 155
rect 18 154 19 155
rect 17 154 18 155
rect 16 154 17 155
rect 15 154 16 155
rect 14 154 15 155
rect 13 154 14 155
rect 12 154 13 155
rect 11 154 12 155
rect 10 154 11 155
rect 9 154 10 155
rect 8 154 9 155
rect 439 155 440 156
rect 438 155 439 156
rect 397 155 398 156
rect 396 155 397 156
rect 395 155 396 156
rect 324 155 325 156
rect 323 155 324 156
rect 322 155 323 156
rect 321 155 322 156
rect 320 155 321 156
rect 319 155 320 156
rect 318 155 319 156
rect 317 155 318 156
rect 316 155 317 156
rect 315 155 316 156
rect 314 155 315 156
rect 313 155 314 156
rect 312 155 313 156
rect 311 155 312 156
rect 310 155 311 156
rect 309 155 310 156
rect 308 155 309 156
rect 307 155 308 156
rect 306 155 307 156
rect 305 155 306 156
rect 304 155 305 156
rect 303 155 304 156
rect 302 155 303 156
rect 301 155 302 156
rect 300 155 301 156
rect 299 155 300 156
rect 298 155 299 156
rect 297 155 298 156
rect 296 155 297 156
rect 295 155 296 156
rect 294 155 295 156
rect 293 155 294 156
rect 292 155 293 156
rect 291 155 292 156
rect 290 155 291 156
rect 289 155 290 156
rect 288 155 289 156
rect 287 155 288 156
rect 286 155 287 156
rect 285 155 286 156
rect 284 155 285 156
rect 283 155 284 156
rect 282 155 283 156
rect 281 155 282 156
rect 280 155 281 156
rect 279 155 280 156
rect 278 155 279 156
rect 277 155 278 156
rect 276 155 277 156
rect 275 155 276 156
rect 274 155 275 156
rect 273 155 274 156
rect 272 155 273 156
rect 271 155 272 156
rect 270 155 271 156
rect 269 155 270 156
rect 268 155 269 156
rect 267 155 268 156
rect 266 155 267 156
rect 265 155 266 156
rect 264 155 265 156
rect 263 155 264 156
rect 262 155 263 156
rect 261 155 262 156
rect 260 155 261 156
rect 259 155 260 156
rect 258 155 259 156
rect 257 155 258 156
rect 256 155 257 156
rect 255 155 256 156
rect 254 155 255 156
rect 253 155 254 156
rect 252 155 253 156
rect 251 155 252 156
rect 250 155 251 156
rect 249 155 250 156
rect 248 155 249 156
rect 247 155 248 156
rect 246 155 247 156
rect 245 155 246 156
rect 244 155 245 156
rect 243 155 244 156
rect 242 155 243 156
rect 241 155 242 156
rect 240 155 241 156
rect 239 155 240 156
rect 238 155 239 156
rect 237 155 238 156
rect 236 155 237 156
rect 216 155 217 156
rect 215 155 216 156
rect 214 155 215 156
rect 213 155 214 156
rect 212 155 213 156
rect 211 155 212 156
rect 210 155 211 156
rect 209 155 210 156
rect 208 155 209 156
rect 207 155 208 156
rect 206 155 207 156
rect 205 155 206 156
rect 204 155 205 156
rect 203 155 204 156
rect 202 155 203 156
rect 201 155 202 156
rect 200 155 201 156
rect 199 155 200 156
rect 198 155 199 156
rect 197 155 198 156
rect 196 155 197 156
rect 195 155 196 156
rect 194 155 195 156
rect 193 155 194 156
rect 192 155 193 156
rect 191 155 192 156
rect 190 155 191 156
rect 189 155 190 156
rect 188 155 189 156
rect 187 155 188 156
rect 186 155 187 156
rect 185 155 186 156
rect 184 155 185 156
rect 183 155 184 156
rect 182 155 183 156
rect 181 155 182 156
rect 180 155 181 156
rect 179 155 180 156
rect 178 155 179 156
rect 177 155 178 156
rect 176 155 177 156
rect 175 155 176 156
rect 174 155 175 156
rect 173 155 174 156
rect 172 155 173 156
rect 171 155 172 156
rect 170 155 171 156
rect 169 155 170 156
rect 168 155 169 156
rect 167 155 168 156
rect 166 155 167 156
rect 165 155 166 156
rect 164 155 165 156
rect 163 155 164 156
rect 162 155 163 156
rect 161 155 162 156
rect 160 155 161 156
rect 159 155 160 156
rect 158 155 159 156
rect 157 155 158 156
rect 156 155 157 156
rect 155 155 156 156
rect 154 155 155 156
rect 153 155 154 156
rect 152 155 153 156
rect 151 155 152 156
rect 150 155 151 156
rect 119 155 120 156
rect 118 155 119 156
rect 117 155 118 156
rect 116 155 117 156
rect 115 155 116 156
rect 114 155 115 156
rect 113 155 114 156
rect 112 155 113 156
rect 111 155 112 156
rect 110 155 111 156
rect 109 155 110 156
rect 108 155 109 156
rect 107 155 108 156
rect 106 155 107 156
rect 105 155 106 156
rect 104 155 105 156
rect 103 155 104 156
rect 102 155 103 156
rect 101 155 102 156
rect 100 155 101 156
rect 99 155 100 156
rect 98 155 99 156
rect 97 155 98 156
rect 96 155 97 156
rect 95 155 96 156
rect 94 155 95 156
rect 93 155 94 156
rect 92 155 93 156
rect 91 155 92 156
rect 90 155 91 156
rect 89 155 90 156
rect 88 155 89 156
rect 87 155 88 156
rect 86 155 87 156
rect 85 155 86 156
rect 84 155 85 156
rect 83 155 84 156
rect 82 155 83 156
rect 81 155 82 156
rect 80 155 81 156
rect 79 155 80 156
rect 78 155 79 156
rect 77 155 78 156
rect 76 155 77 156
rect 75 155 76 156
rect 74 155 75 156
rect 73 155 74 156
rect 72 155 73 156
rect 71 155 72 156
rect 70 155 71 156
rect 69 155 70 156
rect 68 155 69 156
rect 67 155 68 156
rect 66 155 67 156
rect 65 155 66 156
rect 64 155 65 156
rect 63 155 64 156
rect 62 155 63 156
rect 61 155 62 156
rect 60 155 61 156
rect 59 155 60 156
rect 58 155 59 156
rect 57 155 58 156
rect 56 155 57 156
rect 55 155 56 156
rect 54 155 55 156
rect 53 155 54 156
rect 52 155 53 156
rect 51 155 52 156
rect 50 155 51 156
rect 49 155 50 156
rect 48 155 49 156
rect 47 155 48 156
rect 46 155 47 156
rect 45 155 46 156
rect 44 155 45 156
rect 43 155 44 156
rect 42 155 43 156
rect 41 155 42 156
rect 40 155 41 156
rect 39 155 40 156
rect 38 155 39 156
rect 37 155 38 156
rect 36 155 37 156
rect 28 155 29 156
rect 27 155 28 156
rect 26 155 27 156
rect 25 155 26 156
rect 24 155 25 156
rect 23 155 24 156
rect 22 155 23 156
rect 21 155 22 156
rect 20 155 21 156
rect 19 155 20 156
rect 18 155 19 156
rect 17 155 18 156
rect 16 155 17 156
rect 15 155 16 156
rect 14 155 15 156
rect 13 155 14 156
rect 12 155 13 156
rect 11 155 12 156
rect 10 155 11 156
rect 9 155 10 156
rect 8 155 9 156
rect 439 156 440 157
rect 438 156 439 157
rect 437 156 438 157
rect 397 156 398 157
rect 396 156 397 157
rect 395 156 396 157
rect 325 156 326 157
rect 324 156 325 157
rect 323 156 324 157
rect 322 156 323 157
rect 321 156 322 157
rect 320 156 321 157
rect 319 156 320 157
rect 318 156 319 157
rect 317 156 318 157
rect 316 156 317 157
rect 315 156 316 157
rect 314 156 315 157
rect 313 156 314 157
rect 312 156 313 157
rect 311 156 312 157
rect 310 156 311 157
rect 309 156 310 157
rect 308 156 309 157
rect 307 156 308 157
rect 306 156 307 157
rect 305 156 306 157
rect 304 156 305 157
rect 303 156 304 157
rect 302 156 303 157
rect 301 156 302 157
rect 300 156 301 157
rect 299 156 300 157
rect 298 156 299 157
rect 297 156 298 157
rect 296 156 297 157
rect 295 156 296 157
rect 294 156 295 157
rect 293 156 294 157
rect 292 156 293 157
rect 291 156 292 157
rect 290 156 291 157
rect 289 156 290 157
rect 288 156 289 157
rect 287 156 288 157
rect 286 156 287 157
rect 285 156 286 157
rect 284 156 285 157
rect 283 156 284 157
rect 282 156 283 157
rect 281 156 282 157
rect 280 156 281 157
rect 279 156 280 157
rect 278 156 279 157
rect 277 156 278 157
rect 276 156 277 157
rect 275 156 276 157
rect 274 156 275 157
rect 273 156 274 157
rect 272 156 273 157
rect 271 156 272 157
rect 270 156 271 157
rect 269 156 270 157
rect 268 156 269 157
rect 267 156 268 157
rect 266 156 267 157
rect 265 156 266 157
rect 264 156 265 157
rect 263 156 264 157
rect 262 156 263 157
rect 261 156 262 157
rect 260 156 261 157
rect 259 156 260 157
rect 258 156 259 157
rect 257 156 258 157
rect 256 156 257 157
rect 255 156 256 157
rect 254 156 255 157
rect 253 156 254 157
rect 252 156 253 157
rect 251 156 252 157
rect 250 156 251 157
rect 249 156 250 157
rect 248 156 249 157
rect 247 156 248 157
rect 246 156 247 157
rect 245 156 246 157
rect 244 156 245 157
rect 243 156 244 157
rect 242 156 243 157
rect 241 156 242 157
rect 240 156 241 157
rect 239 156 240 157
rect 238 156 239 157
rect 237 156 238 157
rect 236 156 237 157
rect 235 156 236 157
rect 216 156 217 157
rect 215 156 216 157
rect 214 156 215 157
rect 213 156 214 157
rect 212 156 213 157
rect 211 156 212 157
rect 210 156 211 157
rect 209 156 210 157
rect 208 156 209 157
rect 207 156 208 157
rect 206 156 207 157
rect 205 156 206 157
rect 204 156 205 157
rect 203 156 204 157
rect 202 156 203 157
rect 201 156 202 157
rect 200 156 201 157
rect 199 156 200 157
rect 198 156 199 157
rect 197 156 198 157
rect 196 156 197 157
rect 195 156 196 157
rect 194 156 195 157
rect 193 156 194 157
rect 192 156 193 157
rect 191 156 192 157
rect 190 156 191 157
rect 189 156 190 157
rect 188 156 189 157
rect 187 156 188 157
rect 186 156 187 157
rect 185 156 186 157
rect 184 156 185 157
rect 183 156 184 157
rect 182 156 183 157
rect 181 156 182 157
rect 180 156 181 157
rect 179 156 180 157
rect 178 156 179 157
rect 177 156 178 157
rect 176 156 177 157
rect 175 156 176 157
rect 174 156 175 157
rect 173 156 174 157
rect 172 156 173 157
rect 171 156 172 157
rect 170 156 171 157
rect 169 156 170 157
rect 168 156 169 157
rect 167 156 168 157
rect 166 156 167 157
rect 165 156 166 157
rect 164 156 165 157
rect 163 156 164 157
rect 162 156 163 157
rect 161 156 162 157
rect 160 156 161 157
rect 159 156 160 157
rect 158 156 159 157
rect 157 156 158 157
rect 156 156 157 157
rect 155 156 156 157
rect 154 156 155 157
rect 153 156 154 157
rect 152 156 153 157
rect 151 156 152 157
rect 150 156 151 157
rect 149 156 150 157
rect 118 156 119 157
rect 117 156 118 157
rect 116 156 117 157
rect 115 156 116 157
rect 114 156 115 157
rect 113 156 114 157
rect 112 156 113 157
rect 111 156 112 157
rect 110 156 111 157
rect 109 156 110 157
rect 108 156 109 157
rect 107 156 108 157
rect 106 156 107 157
rect 105 156 106 157
rect 104 156 105 157
rect 103 156 104 157
rect 102 156 103 157
rect 101 156 102 157
rect 100 156 101 157
rect 99 156 100 157
rect 98 156 99 157
rect 97 156 98 157
rect 96 156 97 157
rect 95 156 96 157
rect 94 156 95 157
rect 93 156 94 157
rect 92 156 93 157
rect 91 156 92 157
rect 90 156 91 157
rect 89 156 90 157
rect 88 156 89 157
rect 87 156 88 157
rect 86 156 87 157
rect 85 156 86 157
rect 84 156 85 157
rect 83 156 84 157
rect 82 156 83 157
rect 81 156 82 157
rect 80 156 81 157
rect 79 156 80 157
rect 78 156 79 157
rect 77 156 78 157
rect 76 156 77 157
rect 75 156 76 157
rect 74 156 75 157
rect 73 156 74 157
rect 72 156 73 157
rect 71 156 72 157
rect 70 156 71 157
rect 69 156 70 157
rect 68 156 69 157
rect 67 156 68 157
rect 66 156 67 157
rect 65 156 66 157
rect 64 156 65 157
rect 63 156 64 157
rect 62 156 63 157
rect 61 156 62 157
rect 60 156 61 157
rect 59 156 60 157
rect 58 156 59 157
rect 57 156 58 157
rect 56 156 57 157
rect 55 156 56 157
rect 54 156 55 157
rect 53 156 54 157
rect 52 156 53 157
rect 51 156 52 157
rect 50 156 51 157
rect 49 156 50 157
rect 48 156 49 157
rect 47 156 48 157
rect 46 156 47 157
rect 45 156 46 157
rect 44 156 45 157
rect 43 156 44 157
rect 42 156 43 157
rect 41 156 42 157
rect 40 156 41 157
rect 39 156 40 157
rect 38 156 39 157
rect 37 156 38 157
rect 36 156 37 157
rect 27 156 28 157
rect 26 156 27 157
rect 25 156 26 157
rect 24 156 25 157
rect 23 156 24 157
rect 22 156 23 157
rect 21 156 22 157
rect 20 156 21 157
rect 19 156 20 157
rect 18 156 19 157
rect 17 156 18 157
rect 16 156 17 157
rect 15 156 16 157
rect 14 156 15 157
rect 13 156 14 157
rect 12 156 13 157
rect 11 156 12 157
rect 10 156 11 157
rect 9 156 10 157
rect 8 156 9 157
rect 439 157 440 158
rect 438 157 439 158
rect 437 157 438 158
rect 397 157 398 158
rect 396 157 397 158
rect 395 157 396 158
rect 326 157 327 158
rect 325 157 326 158
rect 324 157 325 158
rect 323 157 324 158
rect 322 157 323 158
rect 321 157 322 158
rect 320 157 321 158
rect 319 157 320 158
rect 318 157 319 158
rect 317 157 318 158
rect 316 157 317 158
rect 315 157 316 158
rect 314 157 315 158
rect 313 157 314 158
rect 312 157 313 158
rect 311 157 312 158
rect 310 157 311 158
rect 309 157 310 158
rect 308 157 309 158
rect 307 157 308 158
rect 306 157 307 158
rect 305 157 306 158
rect 304 157 305 158
rect 303 157 304 158
rect 302 157 303 158
rect 301 157 302 158
rect 300 157 301 158
rect 299 157 300 158
rect 298 157 299 158
rect 297 157 298 158
rect 296 157 297 158
rect 295 157 296 158
rect 294 157 295 158
rect 293 157 294 158
rect 292 157 293 158
rect 291 157 292 158
rect 290 157 291 158
rect 289 157 290 158
rect 288 157 289 158
rect 287 157 288 158
rect 286 157 287 158
rect 285 157 286 158
rect 284 157 285 158
rect 283 157 284 158
rect 282 157 283 158
rect 281 157 282 158
rect 280 157 281 158
rect 279 157 280 158
rect 278 157 279 158
rect 277 157 278 158
rect 276 157 277 158
rect 275 157 276 158
rect 274 157 275 158
rect 273 157 274 158
rect 272 157 273 158
rect 271 157 272 158
rect 270 157 271 158
rect 269 157 270 158
rect 268 157 269 158
rect 267 157 268 158
rect 266 157 267 158
rect 265 157 266 158
rect 264 157 265 158
rect 263 157 264 158
rect 262 157 263 158
rect 261 157 262 158
rect 260 157 261 158
rect 259 157 260 158
rect 258 157 259 158
rect 257 157 258 158
rect 256 157 257 158
rect 255 157 256 158
rect 254 157 255 158
rect 253 157 254 158
rect 252 157 253 158
rect 251 157 252 158
rect 250 157 251 158
rect 249 157 250 158
rect 248 157 249 158
rect 247 157 248 158
rect 246 157 247 158
rect 245 157 246 158
rect 244 157 245 158
rect 243 157 244 158
rect 242 157 243 158
rect 241 157 242 158
rect 240 157 241 158
rect 239 157 240 158
rect 238 157 239 158
rect 237 157 238 158
rect 236 157 237 158
rect 235 157 236 158
rect 215 157 216 158
rect 214 157 215 158
rect 213 157 214 158
rect 212 157 213 158
rect 211 157 212 158
rect 210 157 211 158
rect 209 157 210 158
rect 208 157 209 158
rect 207 157 208 158
rect 206 157 207 158
rect 205 157 206 158
rect 204 157 205 158
rect 203 157 204 158
rect 202 157 203 158
rect 201 157 202 158
rect 200 157 201 158
rect 199 157 200 158
rect 198 157 199 158
rect 197 157 198 158
rect 196 157 197 158
rect 195 157 196 158
rect 194 157 195 158
rect 193 157 194 158
rect 192 157 193 158
rect 191 157 192 158
rect 190 157 191 158
rect 189 157 190 158
rect 188 157 189 158
rect 187 157 188 158
rect 186 157 187 158
rect 185 157 186 158
rect 184 157 185 158
rect 183 157 184 158
rect 182 157 183 158
rect 181 157 182 158
rect 180 157 181 158
rect 179 157 180 158
rect 178 157 179 158
rect 177 157 178 158
rect 176 157 177 158
rect 175 157 176 158
rect 174 157 175 158
rect 173 157 174 158
rect 172 157 173 158
rect 171 157 172 158
rect 170 157 171 158
rect 169 157 170 158
rect 168 157 169 158
rect 167 157 168 158
rect 166 157 167 158
rect 165 157 166 158
rect 164 157 165 158
rect 163 157 164 158
rect 162 157 163 158
rect 161 157 162 158
rect 160 157 161 158
rect 159 157 160 158
rect 158 157 159 158
rect 157 157 158 158
rect 156 157 157 158
rect 155 157 156 158
rect 154 157 155 158
rect 153 157 154 158
rect 152 157 153 158
rect 151 157 152 158
rect 150 157 151 158
rect 149 157 150 158
rect 148 157 149 158
rect 117 157 118 158
rect 116 157 117 158
rect 115 157 116 158
rect 114 157 115 158
rect 113 157 114 158
rect 112 157 113 158
rect 111 157 112 158
rect 110 157 111 158
rect 109 157 110 158
rect 108 157 109 158
rect 107 157 108 158
rect 106 157 107 158
rect 105 157 106 158
rect 104 157 105 158
rect 103 157 104 158
rect 102 157 103 158
rect 101 157 102 158
rect 100 157 101 158
rect 99 157 100 158
rect 98 157 99 158
rect 97 157 98 158
rect 96 157 97 158
rect 95 157 96 158
rect 94 157 95 158
rect 93 157 94 158
rect 92 157 93 158
rect 91 157 92 158
rect 90 157 91 158
rect 89 157 90 158
rect 88 157 89 158
rect 87 157 88 158
rect 86 157 87 158
rect 85 157 86 158
rect 84 157 85 158
rect 83 157 84 158
rect 82 157 83 158
rect 81 157 82 158
rect 80 157 81 158
rect 79 157 80 158
rect 78 157 79 158
rect 77 157 78 158
rect 76 157 77 158
rect 75 157 76 158
rect 74 157 75 158
rect 73 157 74 158
rect 72 157 73 158
rect 71 157 72 158
rect 70 157 71 158
rect 69 157 70 158
rect 68 157 69 158
rect 67 157 68 158
rect 66 157 67 158
rect 65 157 66 158
rect 64 157 65 158
rect 63 157 64 158
rect 62 157 63 158
rect 61 157 62 158
rect 60 157 61 158
rect 59 157 60 158
rect 58 157 59 158
rect 57 157 58 158
rect 56 157 57 158
rect 55 157 56 158
rect 54 157 55 158
rect 53 157 54 158
rect 52 157 53 158
rect 51 157 52 158
rect 50 157 51 158
rect 49 157 50 158
rect 48 157 49 158
rect 47 157 48 158
rect 46 157 47 158
rect 45 157 46 158
rect 44 157 45 158
rect 43 157 44 158
rect 42 157 43 158
rect 41 157 42 158
rect 40 157 41 158
rect 39 157 40 158
rect 38 157 39 158
rect 37 157 38 158
rect 36 157 37 158
rect 35 157 36 158
rect 27 157 28 158
rect 26 157 27 158
rect 25 157 26 158
rect 24 157 25 158
rect 23 157 24 158
rect 22 157 23 158
rect 21 157 22 158
rect 20 157 21 158
rect 19 157 20 158
rect 18 157 19 158
rect 17 157 18 158
rect 16 157 17 158
rect 15 157 16 158
rect 14 157 15 158
rect 13 157 14 158
rect 12 157 13 158
rect 11 157 12 158
rect 10 157 11 158
rect 9 157 10 158
rect 8 157 9 158
rect 7 157 8 158
rect 439 158 440 159
rect 438 158 439 159
rect 437 158 438 159
rect 398 158 399 159
rect 397 158 398 159
rect 396 158 397 159
rect 395 158 396 159
rect 326 158 327 159
rect 325 158 326 159
rect 324 158 325 159
rect 323 158 324 159
rect 322 158 323 159
rect 321 158 322 159
rect 320 158 321 159
rect 319 158 320 159
rect 318 158 319 159
rect 317 158 318 159
rect 316 158 317 159
rect 315 158 316 159
rect 296 158 297 159
rect 295 158 296 159
rect 294 158 295 159
rect 293 158 294 159
rect 292 158 293 159
rect 291 158 292 159
rect 290 158 291 159
rect 289 158 290 159
rect 288 158 289 159
rect 287 158 288 159
rect 286 158 287 159
rect 285 158 286 159
rect 284 158 285 159
rect 283 158 284 159
rect 282 158 283 159
rect 281 158 282 159
rect 280 158 281 159
rect 279 158 280 159
rect 278 158 279 159
rect 277 158 278 159
rect 276 158 277 159
rect 275 158 276 159
rect 274 158 275 159
rect 273 158 274 159
rect 272 158 273 159
rect 271 158 272 159
rect 270 158 271 159
rect 269 158 270 159
rect 268 158 269 159
rect 267 158 268 159
rect 266 158 267 159
rect 265 158 266 159
rect 264 158 265 159
rect 263 158 264 159
rect 262 158 263 159
rect 261 158 262 159
rect 260 158 261 159
rect 259 158 260 159
rect 258 158 259 159
rect 257 158 258 159
rect 256 158 257 159
rect 255 158 256 159
rect 254 158 255 159
rect 253 158 254 159
rect 252 158 253 159
rect 251 158 252 159
rect 250 158 251 159
rect 249 158 250 159
rect 248 158 249 159
rect 247 158 248 159
rect 246 158 247 159
rect 245 158 246 159
rect 244 158 245 159
rect 243 158 244 159
rect 242 158 243 159
rect 241 158 242 159
rect 240 158 241 159
rect 239 158 240 159
rect 238 158 239 159
rect 237 158 238 159
rect 236 158 237 159
rect 235 158 236 159
rect 234 158 235 159
rect 215 158 216 159
rect 214 158 215 159
rect 213 158 214 159
rect 212 158 213 159
rect 211 158 212 159
rect 210 158 211 159
rect 209 158 210 159
rect 208 158 209 159
rect 207 158 208 159
rect 206 158 207 159
rect 205 158 206 159
rect 204 158 205 159
rect 203 158 204 159
rect 202 158 203 159
rect 201 158 202 159
rect 200 158 201 159
rect 199 158 200 159
rect 198 158 199 159
rect 197 158 198 159
rect 196 158 197 159
rect 195 158 196 159
rect 194 158 195 159
rect 193 158 194 159
rect 192 158 193 159
rect 191 158 192 159
rect 190 158 191 159
rect 189 158 190 159
rect 188 158 189 159
rect 187 158 188 159
rect 186 158 187 159
rect 185 158 186 159
rect 184 158 185 159
rect 183 158 184 159
rect 182 158 183 159
rect 181 158 182 159
rect 180 158 181 159
rect 179 158 180 159
rect 178 158 179 159
rect 177 158 178 159
rect 176 158 177 159
rect 175 158 176 159
rect 174 158 175 159
rect 173 158 174 159
rect 172 158 173 159
rect 171 158 172 159
rect 170 158 171 159
rect 169 158 170 159
rect 168 158 169 159
rect 167 158 168 159
rect 166 158 167 159
rect 165 158 166 159
rect 164 158 165 159
rect 163 158 164 159
rect 162 158 163 159
rect 161 158 162 159
rect 160 158 161 159
rect 159 158 160 159
rect 158 158 159 159
rect 157 158 158 159
rect 156 158 157 159
rect 155 158 156 159
rect 154 158 155 159
rect 153 158 154 159
rect 152 158 153 159
rect 151 158 152 159
rect 150 158 151 159
rect 149 158 150 159
rect 148 158 149 159
rect 147 158 148 159
rect 115 158 116 159
rect 114 158 115 159
rect 113 158 114 159
rect 112 158 113 159
rect 111 158 112 159
rect 110 158 111 159
rect 109 158 110 159
rect 108 158 109 159
rect 107 158 108 159
rect 106 158 107 159
rect 105 158 106 159
rect 104 158 105 159
rect 103 158 104 159
rect 102 158 103 159
rect 101 158 102 159
rect 100 158 101 159
rect 99 158 100 159
rect 98 158 99 159
rect 97 158 98 159
rect 96 158 97 159
rect 95 158 96 159
rect 94 158 95 159
rect 93 158 94 159
rect 92 158 93 159
rect 91 158 92 159
rect 90 158 91 159
rect 89 158 90 159
rect 88 158 89 159
rect 87 158 88 159
rect 86 158 87 159
rect 85 158 86 159
rect 84 158 85 159
rect 83 158 84 159
rect 82 158 83 159
rect 81 158 82 159
rect 80 158 81 159
rect 79 158 80 159
rect 78 158 79 159
rect 77 158 78 159
rect 76 158 77 159
rect 75 158 76 159
rect 74 158 75 159
rect 73 158 74 159
rect 72 158 73 159
rect 71 158 72 159
rect 70 158 71 159
rect 69 158 70 159
rect 68 158 69 159
rect 67 158 68 159
rect 66 158 67 159
rect 65 158 66 159
rect 64 158 65 159
rect 63 158 64 159
rect 62 158 63 159
rect 61 158 62 159
rect 60 158 61 159
rect 59 158 60 159
rect 58 158 59 159
rect 57 158 58 159
rect 56 158 57 159
rect 55 158 56 159
rect 54 158 55 159
rect 53 158 54 159
rect 52 158 53 159
rect 51 158 52 159
rect 50 158 51 159
rect 49 158 50 159
rect 48 158 49 159
rect 47 158 48 159
rect 46 158 47 159
rect 45 158 46 159
rect 44 158 45 159
rect 43 158 44 159
rect 42 158 43 159
rect 41 158 42 159
rect 40 158 41 159
rect 39 158 40 159
rect 38 158 39 159
rect 37 158 38 159
rect 36 158 37 159
rect 35 158 36 159
rect 26 158 27 159
rect 25 158 26 159
rect 24 158 25 159
rect 23 158 24 159
rect 22 158 23 159
rect 21 158 22 159
rect 20 158 21 159
rect 19 158 20 159
rect 18 158 19 159
rect 17 158 18 159
rect 16 158 17 159
rect 15 158 16 159
rect 14 158 15 159
rect 13 158 14 159
rect 12 158 13 159
rect 11 158 12 159
rect 10 158 11 159
rect 9 158 10 159
rect 8 158 9 159
rect 7 158 8 159
rect 439 159 440 160
rect 438 159 439 160
rect 437 159 438 160
rect 436 159 437 160
rect 398 159 399 160
rect 397 159 398 160
rect 396 159 397 160
rect 395 159 396 160
rect 327 159 328 160
rect 326 159 327 160
rect 325 159 326 160
rect 324 159 325 160
rect 323 159 324 160
rect 322 159 323 160
rect 321 159 322 160
rect 292 159 293 160
rect 291 159 292 160
rect 290 159 291 160
rect 289 159 290 160
rect 288 159 289 160
rect 287 159 288 160
rect 286 159 287 160
rect 285 159 286 160
rect 284 159 285 160
rect 283 159 284 160
rect 282 159 283 160
rect 281 159 282 160
rect 280 159 281 160
rect 279 159 280 160
rect 278 159 279 160
rect 277 159 278 160
rect 276 159 277 160
rect 275 159 276 160
rect 274 159 275 160
rect 273 159 274 160
rect 272 159 273 160
rect 271 159 272 160
rect 270 159 271 160
rect 269 159 270 160
rect 268 159 269 160
rect 267 159 268 160
rect 266 159 267 160
rect 265 159 266 160
rect 264 159 265 160
rect 263 159 264 160
rect 262 159 263 160
rect 261 159 262 160
rect 260 159 261 160
rect 259 159 260 160
rect 258 159 259 160
rect 257 159 258 160
rect 256 159 257 160
rect 255 159 256 160
rect 254 159 255 160
rect 253 159 254 160
rect 252 159 253 160
rect 251 159 252 160
rect 250 159 251 160
rect 249 159 250 160
rect 248 159 249 160
rect 247 159 248 160
rect 246 159 247 160
rect 245 159 246 160
rect 244 159 245 160
rect 243 159 244 160
rect 242 159 243 160
rect 241 159 242 160
rect 240 159 241 160
rect 239 159 240 160
rect 238 159 239 160
rect 237 159 238 160
rect 236 159 237 160
rect 235 159 236 160
rect 234 159 235 160
rect 233 159 234 160
rect 214 159 215 160
rect 213 159 214 160
rect 212 159 213 160
rect 211 159 212 160
rect 210 159 211 160
rect 209 159 210 160
rect 208 159 209 160
rect 207 159 208 160
rect 206 159 207 160
rect 205 159 206 160
rect 204 159 205 160
rect 203 159 204 160
rect 202 159 203 160
rect 201 159 202 160
rect 200 159 201 160
rect 199 159 200 160
rect 198 159 199 160
rect 197 159 198 160
rect 196 159 197 160
rect 195 159 196 160
rect 194 159 195 160
rect 193 159 194 160
rect 192 159 193 160
rect 191 159 192 160
rect 190 159 191 160
rect 189 159 190 160
rect 188 159 189 160
rect 187 159 188 160
rect 186 159 187 160
rect 185 159 186 160
rect 184 159 185 160
rect 183 159 184 160
rect 182 159 183 160
rect 181 159 182 160
rect 180 159 181 160
rect 179 159 180 160
rect 178 159 179 160
rect 177 159 178 160
rect 176 159 177 160
rect 175 159 176 160
rect 174 159 175 160
rect 173 159 174 160
rect 172 159 173 160
rect 171 159 172 160
rect 170 159 171 160
rect 169 159 170 160
rect 168 159 169 160
rect 167 159 168 160
rect 166 159 167 160
rect 165 159 166 160
rect 164 159 165 160
rect 163 159 164 160
rect 162 159 163 160
rect 161 159 162 160
rect 160 159 161 160
rect 159 159 160 160
rect 158 159 159 160
rect 157 159 158 160
rect 156 159 157 160
rect 155 159 156 160
rect 154 159 155 160
rect 153 159 154 160
rect 152 159 153 160
rect 151 159 152 160
rect 150 159 151 160
rect 149 159 150 160
rect 148 159 149 160
rect 147 159 148 160
rect 114 159 115 160
rect 113 159 114 160
rect 112 159 113 160
rect 111 159 112 160
rect 110 159 111 160
rect 109 159 110 160
rect 108 159 109 160
rect 107 159 108 160
rect 106 159 107 160
rect 105 159 106 160
rect 104 159 105 160
rect 103 159 104 160
rect 102 159 103 160
rect 101 159 102 160
rect 100 159 101 160
rect 99 159 100 160
rect 98 159 99 160
rect 97 159 98 160
rect 96 159 97 160
rect 95 159 96 160
rect 94 159 95 160
rect 93 159 94 160
rect 92 159 93 160
rect 91 159 92 160
rect 90 159 91 160
rect 89 159 90 160
rect 88 159 89 160
rect 87 159 88 160
rect 86 159 87 160
rect 85 159 86 160
rect 84 159 85 160
rect 83 159 84 160
rect 82 159 83 160
rect 81 159 82 160
rect 80 159 81 160
rect 79 159 80 160
rect 78 159 79 160
rect 77 159 78 160
rect 76 159 77 160
rect 75 159 76 160
rect 74 159 75 160
rect 73 159 74 160
rect 72 159 73 160
rect 71 159 72 160
rect 70 159 71 160
rect 69 159 70 160
rect 68 159 69 160
rect 67 159 68 160
rect 66 159 67 160
rect 65 159 66 160
rect 64 159 65 160
rect 63 159 64 160
rect 62 159 63 160
rect 61 159 62 160
rect 60 159 61 160
rect 59 159 60 160
rect 58 159 59 160
rect 57 159 58 160
rect 56 159 57 160
rect 55 159 56 160
rect 54 159 55 160
rect 53 159 54 160
rect 52 159 53 160
rect 51 159 52 160
rect 50 159 51 160
rect 49 159 50 160
rect 48 159 49 160
rect 47 159 48 160
rect 46 159 47 160
rect 45 159 46 160
rect 44 159 45 160
rect 43 159 44 160
rect 42 159 43 160
rect 41 159 42 160
rect 40 159 41 160
rect 39 159 40 160
rect 38 159 39 160
rect 37 159 38 160
rect 36 159 37 160
rect 35 159 36 160
rect 34 159 35 160
rect 25 159 26 160
rect 24 159 25 160
rect 23 159 24 160
rect 22 159 23 160
rect 21 159 22 160
rect 20 159 21 160
rect 19 159 20 160
rect 18 159 19 160
rect 17 159 18 160
rect 16 159 17 160
rect 15 159 16 160
rect 14 159 15 160
rect 13 159 14 160
rect 12 159 13 160
rect 11 159 12 160
rect 10 159 11 160
rect 9 159 10 160
rect 8 159 9 160
rect 7 159 8 160
rect 460 160 461 161
rect 439 160 440 161
rect 438 160 439 161
rect 437 160 438 161
rect 436 160 437 161
rect 435 160 436 161
rect 434 160 435 161
rect 400 160 401 161
rect 399 160 400 161
rect 398 160 399 161
rect 397 160 398 161
rect 396 160 397 161
rect 395 160 396 161
rect 328 160 329 161
rect 327 160 328 161
rect 326 160 327 161
rect 325 160 326 161
rect 289 160 290 161
rect 288 160 289 161
rect 287 160 288 161
rect 286 160 287 161
rect 285 160 286 161
rect 284 160 285 161
rect 283 160 284 161
rect 282 160 283 161
rect 281 160 282 161
rect 280 160 281 161
rect 279 160 280 161
rect 278 160 279 161
rect 277 160 278 161
rect 276 160 277 161
rect 275 160 276 161
rect 274 160 275 161
rect 273 160 274 161
rect 272 160 273 161
rect 271 160 272 161
rect 270 160 271 161
rect 269 160 270 161
rect 268 160 269 161
rect 267 160 268 161
rect 266 160 267 161
rect 265 160 266 161
rect 264 160 265 161
rect 263 160 264 161
rect 262 160 263 161
rect 261 160 262 161
rect 260 160 261 161
rect 259 160 260 161
rect 258 160 259 161
rect 257 160 258 161
rect 256 160 257 161
rect 255 160 256 161
rect 254 160 255 161
rect 253 160 254 161
rect 252 160 253 161
rect 251 160 252 161
rect 250 160 251 161
rect 249 160 250 161
rect 248 160 249 161
rect 247 160 248 161
rect 246 160 247 161
rect 245 160 246 161
rect 244 160 245 161
rect 243 160 244 161
rect 242 160 243 161
rect 241 160 242 161
rect 240 160 241 161
rect 239 160 240 161
rect 238 160 239 161
rect 237 160 238 161
rect 236 160 237 161
rect 235 160 236 161
rect 234 160 235 161
rect 233 160 234 161
rect 214 160 215 161
rect 213 160 214 161
rect 212 160 213 161
rect 211 160 212 161
rect 210 160 211 161
rect 209 160 210 161
rect 208 160 209 161
rect 207 160 208 161
rect 206 160 207 161
rect 205 160 206 161
rect 204 160 205 161
rect 203 160 204 161
rect 202 160 203 161
rect 201 160 202 161
rect 200 160 201 161
rect 199 160 200 161
rect 198 160 199 161
rect 197 160 198 161
rect 196 160 197 161
rect 195 160 196 161
rect 194 160 195 161
rect 193 160 194 161
rect 192 160 193 161
rect 191 160 192 161
rect 190 160 191 161
rect 189 160 190 161
rect 188 160 189 161
rect 187 160 188 161
rect 186 160 187 161
rect 185 160 186 161
rect 184 160 185 161
rect 183 160 184 161
rect 182 160 183 161
rect 181 160 182 161
rect 180 160 181 161
rect 179 160 180 161
rect 178 160 179 161
rect 177 160 178 161
rect 176 160 177 161
rect 175 160 176 161
rect 174 160 175 161
rect 173 160 174 161
rect 172 160 173 161
rect 171 160 172 161
rect 170 160 171 161
rect 169 160 170 161
rect 168 160 169 161
rect 167 160 168 161
rect 166 160 167 161
rect 165 160 166 161
rect 164 160 165 161
rect 163 160 164 161
rect 162 160 163 161
rect 161 160 162 161
rect 160 160 161 161
rect 159 160 160 161
rect 158 160 159 161
rect 157 160 158 161
rect 156 160 157 161
rect 155 160 156 161
rect 154 160 155 161
rect 153 160 154 161
rect 152 160 153 161
rect 151 160 152 161
rect 150 160 151 161
rect 149 160 150 161
rect 148 160 149 161
rect 147 160 148 161
rect 146 160 147 161
rect 112 160 113 161
rect 111 160 112 161
rect 110 160 111 161
rect 109 160 110 161
rect 108 160 109 161
rect 107 160 108 161
rect 106 160 107 161
rect 105 160 106 161
rect 104 160 105 161
rect 103 160 104 161
rect 102 160 103 161
rect 101 160 102 161
rect 100 160 101 161
rect 99 160 100 161
rect 98 160 99 161
rect 97 160 98 161
rect 96 160 97 161
rect 95 160 96 161
rect 94 160 95 161
rect 93 160 94 161
rect 92 160 93 161
rect 91 160 92 161
rect 90 160 91 161
rect 89 160 90 161
rect 88 160 89 161
rect 87 160 88 161
rect 86 160 87 161
rect 85 160 86 161
rect 84 160 85 161
rect 83 160 84 161
rect 82 160 83 161
rect 81 160 82 161
rect 80 160 81 161
rect 79 160 80 161
rect 78 160 79 161
rect 77 160 78 161
rect 76 160 77 161
rect 75 160 76 161
rect 74 160 75 161
rect 73 160 74 161
rect 72 160 73 161
rect 71 160 72 161
rect 70 160 71 161
rect 69 160 70 161
rect 68 160 69 161
rect 67 160 68 161
rect 66 160 67 161
rect 65 160 66 161
rect 64 160 65 161
rect 63 160 64 161
rect 62 160 63 161
rect 61 160 62 161
rect 60 160 61 161
rect 59 160 60 161
rect 58 160 59 161
rect 57 160 58 161
rect 56 160 57 161
rect 55 160 56 161
rect 54 160 55 161
rect 53 160 54 161
rect 52 160 53 161
rect 51 160 52 161
rect 50 160 51 161
rect 49 160 50 161
rect 48 160 49 161
rect 47 160 48 161
rect 46 160 47 161
rect 45 160 46 161
rect 44 160 45 161
rect 43 160 44 161
rect 42 160 43 161
rect 41 160 42 161
rect 40 160 41 161
rect 39 160 40 161
rect 38 160 39 161
rect 37 160 38 161
rect 36 160 37 161
rect 35 160 36 161
rect 34 160 35 161
rect 25 160 26 161
rect 24 160 25 161
rect 23 160 24 161
rect 22 160 23 161
rect 21 160 22 161
rect 20 160 21 161
rect 19 160 20 161
rect 18 160 19 161
rect 17 160 18 161
rect 16 160 17 161
rect 15 160 16 161
rect 14 160 15 161
rect 13 160 14 161
rect 12 160 13 161
rect 11 160 12 161
rect 10 160 11 161
rect 9 160 10 161
rect 8 160 9 161
rect 7 160 8 161
rect 460 161 461 162
rect 439 161 440 162
rect 438 161 439 162
rect 437 161 438 162
rect 436 161 437 162
rect 435 161 436 162
rect 434 161 435 162
rect 433 161 434 162
rect 432 161 433 162
rect 431 161 432 162
rect 430 161 431 162
rect 429 161 430 162
rect 428 161 429 162
rect 427 161 428 162
rect 426 161 427 162
rect 425 161 426 162
rect 424 161 425 162
rect 423 161 424 162
rect 422 161 423 162
rect 421 161 422 162
rect 420 161 421 162
rect 419 161 420 162
rect 418 161 419 162
rect 417 161 418 162
rect 416 161 417 162
rect 415 161 416 162
rect 414 161 415 162
rect 413 161 414 162
rect 412 161 413 162
rect 411 161 412 162
rect 410 161 411 162
rect 409 161 410 162
rect 408 161 409 162
rect 407 161 408 162
rect 406 161 407 162
rect 405 161 406 162
rect 404 161 405 162
rect 403 161 404 162
rect 402 161 403 162
rect 401 161 402 162
rect 400 161 401 162
rect 399 161 400 162
rect 398 161 399 162
rect 397 161 398 162
rect 396 161 397 162
rect 395 161 396 162
rect 286 161 287 162
rect 285 161 286 162
rect 284 161 285 162
rect 283 161 284 162
rect 282 161 283 162
rect 281 161 282 162
rect 280 161 281 162
rect 279 161 280 162
rect 278 161 279 162
rect 277 161 278 162
rect 276 161 277 162
rect 275 161 276 162
rect 274 161 275 162
rect 273 161 274 162
rect 272 161 273 162
rect 271 161 272 162
rect 270 161 271 162
rect 269 161 270 162
rect 268 161 269 162
rect 267 161 268 162
rect 266 161 267 162
rect 265 161 266 162
rect 264 161 265 162
rect 263 161 264 162
rect 262 161 263 162
rect 261 161 262 162
rect 260 161 261 162
rect 259 161 260 162
rect 258 161 259 162
rect 257 161 258 162
rect 256 161 257 162
rect 255 161 256 162
rect 254 161 255 162
rect 253 161 254 162
rect 252 161 253 162
rect 251 161 252 162
rect 250 161 251 162
rect 249 161 250 162
rect 248 161 249 162
rect 247 161 248 162
rect 246 161 247 162
rect 245 161 246 162
rect 244 161 245 162
rect 243 161 244 162
rect 242 161 243 162
rect 241 161 242 162
rect 240 161 241 162
rect 239 161 240 162
rect 238 161 239 162
rect 237 161 238 162
rect 236 161 237 162
rect 235 161 236 162
rect 234 161 235 162
rect 233 161 234 162
rect 232 161 233 162
rect 213 161 214 162
rect 212 161 213 162
rect 211 161 212 162
rect 210 161 211 162
rect 209 161 210 162
rect 208 161 209 162
rect 207 161 208 162
rect 206 161 207 162
rect 205 161 206 162
rect 204 161 205 162
rect 203 161 204 162
rect 202 161 203 162
rect 201 161 202 162
rect 200 161 201 162
rect 199 161 200 162
rect 198 161 199 162
rect 197 161 198 162
rect 196 161 197 162
rect 195 161 196 162
rect 194 161 195 162
rect 193 161 194 162
rect 192 161 193 162
rect 191 161 192 162
rect 190 161 191 162
rect 189 161 190 162
rect 188 161 189 162
rect 187 161 188 162
rect 186 161 187 162
rect 185 161 186 162
rect 184 161 185 162
rect 183 161 184 162
rect 182 161 183 162
rect 181 161 182 162
rect 180 161 181 162
rect 179 161 180 162
rect 178 161 179 162
rect 177 161 178 162
rect 176 161 177 162
rect 175 161 176 162
rect 174 161 175 162
rect 173 161 174 162
rect 172 161 173 162
rect 171 161 172 162
rect 170 161 171 162
rect 169 161 170 162
rect 168 161 169 162
rect 167 161 168 162
rect 166 161 167 162
rect 165 161 166 162
rect 164 161 165 162
rect 163 161 164 162
rect 162 161 163 162
rect 161 161 162 162
rect 160 161 161 162
rect 159 161 160 162
rect 158 161 159 162
rect 157 161 158 162
rect 156 161 157 162
rect 155 161 156 162
rect 154 161 155 162
rect 153 161 154 162
rect 152 161 153 162
rect 151 161 152 162
rect 150 161 151 162
rect 149 161 150 162
rect 148 161 149 162
rect 147 161 148 162
rect 146 161 147 162
rect 145 161 146 162
rect 111 161 112 162
rect 110 161 111 162
rect 109 161 110 162
rect 108 161 109 162
rect 107 161 108 162
rect 106 161 107 162
rect 105 161 106 162
rect 104 161 105 162
rect 103 161 104 162
rect 102 161 103 162
rect 101 161 102 162
rect 100 161 101 162
rect 99 161 100 162
rect 98 161 99 162
rect 97 161 98 162
rect 96 161 97 162
rect 95 161 96 162
rect 94 161 95 162
rect 93 161 94 162
rect 92 161 93 162
rect 91 161 92 162
rect 90 161 91 162
rect 89 161 90 162
rect 88 161 89 162
rect 87 161 88 162
rect 86 161 87 162
rect 85 161 86 162
rect 84 161 85 162
rect 83 161 84 162
rect 82 161 83 162
rect 81 161 82 162
rect 80 161 81 162
rect 79 161 80 162
rect 78 161 79 162
rect 77 161 78 162
rect 76 161 77 162
rect 75 161 76 162
rect 74 161 75 162
rect 73 161 74 162
rect 72 161 73 162
rect 71 161 72 162
rect 70 161 71 162
rect 69 161 70 162
rect 68 161 69 162
rect 67 161 68 162
rect 66 161 67 162
rect 65 161 66 162
rect 64 161 65 162
rect 63 161 64 162
rect 62 161 63 162
rect 61 161 62 162
rect 60 161 61 162
rect 59 161 60 162
rect 58 161 59 162
rect 57 161 58 162
rect 56 161 57 162
rect 55 161 56 162
rect 54 161 55 162
rect 53 161 54 162
rect 52 161 53 162
rect 51 161 52 162
rect 50 161 51 162
rect 49 161 50 162
rect 48 161 49 162
rect 47 161 48 162
rect 46 161 47 162
rect 45 161 46 162
rect 44 161 45 162
rect 43 161 44 162
rect 42 161 43 162
rect 41 161 42 162
rect 40 161 41 162
rect 39 161 40 162
rect 38 161 39 162
rect 37 161 38 162
rect 36 161 37 162
rect 35 161 36 162
rect 34 161 35 162
rect 24 161 25 162
rect 23 161 24 162
rect 22 161 23 162
rect 21 161 22 162
rect 20 161 21 162
rect 19 161 20 162
rect 18 161 19 162
rect 17 161 18 162
rect 16 161 17 162
rect 15 161 16 162
rect 14 161 15 162
rect 13 161 14 162
rect 12 161 13 162
rect 11 161 12 162
rect 10 161 11 162
rect 9 161 10 162
rect 8 161 9 162
rect 461 162 462 163
rect 460 162 461 163
rect 439 162 440 163
rect 438 162 439 163
rect 437 162 438 163
rect 436 162 437 163
rect 435 162 436 163
rect 434 162 435 163
rect 433 162 434 163
rect 432 162 433 163
rect 431 162 432 163
rect 430 162 431 163
rect 429 162 430 163
rect 428 162 429 163
rect 427 162 428 163
rect 426 162 427 163
rect 425 162 426 163
rect 424 162 425 163
rect 423 162 424 163
rect 422 162 423 163
rect 421 162 422 163
rect 420 162 421 163
rect 419 162 420 163
rect 418 162 419 163
rect 417 162 418 163
rect 416 162 417 163
rect 415 162 416 163
rect 414 162 415 163
rect 413 162 414 163
rect 412 162 413 163
rect 411 162 412 163
rect 410 162 411 163
rect 409 162 410 163
rect 408 162 409 163
rect 407 162 408 163
rect 406 162 407 163
rect 405 162 406 163
rect 404 162 405 163
rect 403 162 404 163
rect 402 162 403 163
rect 401 162 402 163
rect 400 162 401 163
rect 399 162 400 163
rect 398 162 399 163
rect 397 162 398 163
rect 396 162 397 163
rect 395 162 396 163
rect 284 162 285 163
rect 283 162 284 163
rect 282 162 283 163
rect 281 162 282 163
rect 280 162 281 163
rect 279 162 280 163
rect 278 162 279 163
rect 277 162 278 163
rect 276 162 277 163
rect 275 162 276 163
rect 274 162 275 163
rect 273 162 274 163
rect 272 162 273 163
rect 271 162 272 163
rect 270 162 271 163
rect 269 162 270 163
rect 268 162 269 163
rect 267 162 268 163
rect 266 162 267 163
rect 265 162 266 163
rect 264 162 265 163
rect 263 162 264 163
rect 262 162 263 163
rect 261 162 262 163
rect 260 162 261 163
rect 259 162 260 163
rect 258 162 259 163
rect 257 162 258 163
rect 256 162 257 163
rect 255 162 256 163
rect 254 162 255 163
rect 253 162 254 163
rect 252 162 253 163
rect 251 162 252 163
rect 250 162 251 163
rect 249 162 250 163
rect 248 162 249 163
rect 247 162 248 163
rect 246 162 247 163
rect 245 162 246 163
rect 244 162 245 163
rect 243 162 244 163
rect 242 162 243 163
rect 241 162 242 163
rect 240 162 241 163
rect 239 162 240 163
rect 238 162 239 163
rect 237 162 238 163
rect 236 162 237 163
rect 235 162 236 163
rect 234 162 235 163
rect 233 162 234 163
rect 232 162 233 163
rect 213 162 214 163
rect 212 162 213 163
rect 211 162 212 163
rect 210 162 211 163
rect 209 162 210 163
rect 208 162 209 163
rect 207 162 208 163
rect 206 162 207 163
rect 205 162 206 163
rect 204 162 205 163
rect 203 162 204 163
rect 202 162 203 163
rect 201 162 202 163
rect 200 162 201 163
rect 199 162 200 163
rect 198 162 199 163
rect 197 162 198 163
rect 196 162 197 163
rect 195 162 196 163
rect 194 162 195 163
rect 193 162 194 163
rect 192 162 193 163
rect 191 162 192 163
rect 190 162 191 163
rect 189 162 190 163
rect 188 162 189 163
rect 187 162 188 163
rect 186 162 187 163
rect 185 162 186 163
rect 184 162 185 163
rect 183 162 184 163
rect 182 162 183 163
rect 181 162 182 163
rect 180 162 181 163
rect 179 162 180 163
rect 178 162 179 163
rect 177 162 178 163
rect 176 162 177 163
rect 175 162 176 163
rect 174 162 175 163
rect 173 162 174 163
rect 172 162 173 163
rect 171 162 172 163
rect 170 162 171 163
rect 169 162 170 163
rect 168 162 169 163
rect 167 162 168 163
rect 166 162 167 163
rect 165 162 166 163
rect 164 162 165 163
rect 163 162 164 163
rect 162 162 163 163
rect 161 162 162 163
rect 160 162 161 163
rect 159 162 160 163
rect 158 162 159 163
rect 157 162 158 163
rect 156 162 157 163
rect 155 162 156 163
rect 154 162 155 163
rect 153 162 154 163
rect 152 162 153 163
rect 151 162 152 163
rect 150 162 151 163
rect 149 162 150 163
rect 148 162 149 163
rect 147 162 148 163
rect 146 162 147 163
rect 145 162 146 163
rect 144 162 145 163
rect 143 162 144 163
rect 109 162 110 163
rect 108 162 109 163
rect 107 162 108 163
rect 106 162 107 163
rect 105 162 106 163
rect 104 162 105 163
rect 103 162 104 163
rect 102 162 103 163
rect 101 162 102 163
rect 100 162 101 163
rect 99 162 100 163
rect 98 162 99 163
rect 97 162 98 163
rect 96 162 97 163
rect 95 162 96 163
rect 94 162 95 163
rect 93 162 94 163
rect 92 162 93 163
rect 91 162 92 163
rect 90 162 91 163
rect 89 162 90 163
rect 88 162 89 163
rect 87 162 88 163
rect 86 162 87 163
rect 85 162 86 163
rect 84 162 85 163
rect 83 162 84 163
rect 82 162 83 163
rect 81 162 82 163
rect 80 162 81 163
rect 79 162 80 163
rect 78 162 79 163
rect 77 162 78 163
rect 76 162 77 163
rect 75 162 76 163
rect 74 162 75 163
rect 73 162 74 163
rect 72 162 73 163
rect 71 162 72 163
rect 70 162 71 163
rect 69 162 70 163
rect 68 162 69 163
rect 67 162 68 163
rect 66 162 67 163
rect 65 162 66 163
rect 64 162 65 163
rect 63 162 64 163
rect 62 162 63 163
rect 61 162 62 163
rect 60 162 61 163
rect 59 162 60 163
rect 58 162 59 163
rect 57 162 58 163
rect 56 162 57 163
rect 55 162 56 163
rect 54 162 55 163
rect 53 162 54 163
rect 52 162 53 163
rect 51 162 52 163
rect 50 162 51 163
rect 49 162 50 163
rect 48 162 49 163
rect 47 162 48 163
rect 46 162 47 163
rect 45 162 46 163
rect 44 162 45 163
rect 43 162 44 163
rect 42 162 43 163
rect 41 162 42 163
rect 40 162 41 163
rect 39 162 40 163
rect 38 162 39 163
rect 37 162 38 163
rect 36 162 37 163
rect 35 162 36 163
rect 34 162 35 163
rect 24 162 25 163
rect 23 162 24 163
rect 22 162 23 163
rect 21 162 22 163
rect 20 162 21 163
rect 19 162 20 163
rect 18 162 19 163
rect 17 162 18 163
rect 16 162 17 163
rect 15 162 16 163
rect 14 162 15 163
rect 13 162 14 163
rect 12 162 13 163
rect 11 162 12 163
rect 10 162 11 163
rect 9 162 10 163
rect 8 162 9 163
rect 463 163 464 164
rect 462 163 463 164
rect 461 163 462 164
rect 460 163 461 164
rect 439 163 440 164
rect 438 163 439 164
rect 437 163 438 164
rect 436 163 437 164
rect 435 163 436 164
rect 434 163 435 164
rect 433 163 434 164
rect 432 163 433 164
rect 431 163 432 164
rect 430 163 431 164
rect 429 163 430 164
rect 428 163 429 164
rect 427 163 428 164
rect 426 163 427 164
rect 425 163 426 164
rect 424 163 425 164
rect 423 163 424 164
rect 422 163 423 164
rect 421 163 422 164
rect 420 163 421 164
rect 419 163 420 164
rect 418 163 419 164
rect 417 163 418 164
rect 416 163 417 164
rect 415 163 416 164
rect 414 163 415 164
rect 413 163 414 164
rect 412 163 413 164
rect 411 163 412 164
rect 410 163 411 164
rect 409 163 410 164
rect 408 163 409 164
rect 407 163 408 164
rect 406 163 407 164
rect 405 163 406 164
rect 404 163 405 164
rect 403 163 404 164
rect 402 163 403 164
rect 401 163 402 164
rect 400 163 401 164
rect 399 163 400 164
rect 398 163 399 164
rect 397 163 398 164
rect 396 163 397 164
rect 395 163 396 164
rect 282 163 283 164
rect 281 163 282 164
rect 280 163 281 164
rect 279 163 280 164
rect 278 163 279 164
rect 277 163 278 164
rect 276 163 277 164
rect 275 163 276 164
rect 274 163 275 164
rect 273 163 274 164
rect 272 163 273 164
rect 271 163 272 164
rect 270 163 271 164
rect 269 163 270 164
rect 268 163 269 164
rect 267 163 268 164
rect 266 163 267 164
rect 265 163 266 164
rect 264 163 265 164
rect 263 163 264 164
rect 262 163 263 164
rect 261 163 262 164
rect 260 163 261 164
rect 259 163 260 164
rect 258 163 259 164
rect 257 163 258 164
rect 256 163 257 164
rect 255 163 256 164
rect 254 163 255 164
rect 253 163 254 164
rect 252 163 253 164
rect 251 163 252 164
rect 250 163 251 164
rect 249 163 250 164
rect 248 163 249 164
rect 247 163 248 164
rect 246 163 247 164
rect 245 163 246 164
rect 244 163 245 164
rect 243 163 244 164
rect 242 163 243 164
rect 241 163 242 164
rect 240 163 241 164
rect 239 163 240 164
rect 238 163 239 164
rect 237 163 238 164
rect 236 163 237 164
rect 235 163 236 164
rect 234 163 235 164
rect 233 163 234 164
rect 232 163 233 164
rect 231 163 232 164
rect 213 163 214 164
rect 212 163 213 164
rect 211 163 212 164
rect 210 163 211 164
rect 209 163 210 164
rect 208 163 209 164
rect 207 163 208 164
rect 206 163 207 164
rect 205 163 206 164
rect 204 163 205 164
rect 203 163 204 164
rect 202 163 203 164
rect 201 163 202 164
rect 200 163 201 164
rect 199 163 200 164
rect 198 163 199 164
rect 197 163 198 164
rect 196 163 197 164
rect 195 163 196 164
rect 194 163 195 164
rect 193 163 194 164
rect 192 163 193 164
rect 191 163 192 164
rect 190 163 191 164
rect 189 163 190 164
rect 188 163 189 164
rect 187 163 188 164
rect 186 163 187 164
rect 185 163 186 164
rect 184 163 185 164
rect 183 163 184 164
rect 182 163 183 164
rect 181 163 182 164
rect 180 163 181 164
rect 179 163 180 164
rect 178 163 179 164
rect 177 163 178 164
rect 176 163 177 164
rect 175 163 176 164
rect 174 163 175 164
rect 173 163 174 164
rect 172 163 173 164
rect 171 163 172 164
rect 170 163 171 164
rect 169 163 170 164
rect 168 163 169 164
rect 167 163 168 164
rect 166 163 167 164
rect 165 163 166 164
rect 164 163 165 164
rect 163 163 164 164
rect 162 163 163 164
rect 161 163 162 164
rect 160 163 161 164
rect 159 163 160 164
rect 158 163 159 164
rect 157 163 158 164
rect 156 163 157 164
rect 155 163 156 164
rect 154 163 155 164
rect 153 163 154 164
rect 152 163 153 164
rect 151 163 152 164
rect 150 163 151 164
rect 149 163 150 164
rect 148 163 149 164
rect 147 163 148 164
rect 146 163 147 164
rect 145 163 146 164
rect 144 163 145 164
rect 143 163 144 164
rect 142 163 143 164
rect 108 163 109 164
rect 107 163 108 164
rect 106 163 107 164
rect 105 163 106 164
rect 104 163 105 164
rect 103 163 104 164
rect 102 163 103 164
rect 101 163 102 164
rect 100 163 101 164
rect 99 163 100 164
rect 98 163 99 164
rect 97 163 98 164
rect 96 163 97 164
rect 95 163 96 164
rect 94 163 95 164
rect 93 163 94 164
rect 92 163 93 164
rect 91 163 92 164
rect 90 163 91 164
rect 89 163 90 164
rect 88 163 89 164
rect 87 163 88 164
rect 86 163 87 164
rect 85 163 86 164
rect 84 163 85 164
rect 83 163 84 164
rect 82 163 83 164
rect 81 163 82 164
rect 80 163 81 164
rect 79 163 80 164
rect 78 163 79 164
rect 77 163 78 164
rect 76 163 77 164
rect 75 163 76 164
rect 74 163 75 164
rect 73 163 74 164
rect 72 163 73 164
rect 71 163 72 164
rect 70 163 71 164
rect 69 163 70 164
rect 68 163 69 164
rect 67 163 68 164
rect 66 163 67 164
rect 65 163 66 164
rect 64 163 65 164
rect 63 163 64 164
rect 62 163 63 164
rect 61 163 62 164
rect 60 163 61 164
rect 59 163 60 164
rect 58 163 59 164
rect 57 163 58 164
rect 56 163 57 164
rect 55 163 56 164
rect 54 163 55 164
rect 53 163 54 164
rect 52 163 53 164
rect 51 163 52 164
rect 50 163 51 164
rect 49 163 50 164
rect 48 163 49 164
rect 47 163 48 164
rect 46 163 47 164
rect 45 163 46 164
rect 44 163 45 164
rect 43 163 44 164
rect 42 163 43 164
rect 41 163 42 164
rect 40 163 41 164
rect 39 163 40 164
rect 38 163 39 164
rect 37 163 38 164
rect 36 163 37 164
rect 35 163 36 164
rect 34 163 35 164
rect 33 163 34 164
rect 24 163 25 164
rect 23 163 24 164
rect 22 163 23 164
rect 21 163 22 164
rect 20 163 21 164
rect 19 163 20 164
rect 18 163 19 164
rect 17 163 18 164
rect 16 163 17 164
rect 15 163 16 164
rect 14 163 15 164
rect 13 163 14 164
rect 12 163 13 164
rect 11 163 12 164
rect 10 163 11 164
rect 9 163 10 164
rect 8 163 9 164
rect 465 164 466 165
rect 464 164 465 165
rect 463 164 464 165
rect 462 164 463 165
rect 461 164 462 165
rect 460 164 461 165
rect 439 164 440 165
rect 438 164 439 165
rect 437 164 438 165
rect 436 164 437 165
rect 435 164 436 165
rect 434 164 435 165
rect 433 164 434 165
rect 432 164 433 165
rect 431 164 432 165
rect 430 164 431 165
rect 429 164 430 165
rect 428 164 429 165
rect 427 164 428 165
rect 426 164 427 165
rect 425 164 426 165
rect 424 164 425 165
rect 423 164 424 165
rect 422 164 423 165
rect 421 164 422 165
rect 420 164 421 165
rect 419 164 420 165
rect 418 164 419 165
rect 417 164 418 165
rect 416 164 417 165
rect 415 164 416 165
rect 414 164 415 165
rect 413 164 414 165
rect 412 164 413 165
rect 411 164 412 165
rect 410 164 411 165
rect 409 164 410 165
rect 408 164 409 165
rect 407 164 408 165
rect 406 164 407 165
rect 405 164 406 165
rect 404 164 405 165
rect 403 164 404 165
rect 402 164 403 165
rect 401 164 402 165
rect 400 164 401 165
rect 399 164 400 165
rect 398 164 399 165
rect 397 164 398 165
rect 396 164 397 165
rect 395 164 396 165
rect 280 164 281 165
rect 279 164 280 165
rect 278 164 279 165
rect 277 164 278 165
rect 276 164 277 165
rect 275 164 276 165
rect 274 164 275 165
rect 273 164 274 165
rect 272 164 273 165
rect 271 164 272 165
rect 270 164 271 165
rect 269 164 270 165
rect 268 164 269 165
rect 267 164 268 165
rect 266 164 267 165
rect 265 164 266 165
rect 264 164 265 165
rect 263 164 264 165
rect 262 164 263 165
rect 261 164 262 165
rect 260 164 261 165
rect 259 164 260 165
rect 258 164 259 165
rect 257 164 258 165
rect 256 164 257 165
rect 255 164 256 165
rect 254 164 255 165
rect 253 164 254 165
rect 252 164 253 165
rect 251 164 252 165
rect 250 164 251 165
rect 249 164 250 165
rect 248 164 249 165
rect 247 164 248 165
rect 246 164 247 165
rect 245 164 246 165
rect 244 164 245 165
rect 243 164 244 165
rect 242 164 243 165
rect 241 164 242 165
rect 240 164 241 165
rect 239 164 240 165
rect 238 164 239 165
rect 237 164 238 165
rect 236 164 237 165
rect 235 164 236 165
rect 234 164 235 165
rect 233 164 234 165
rect 232 164 233 165
rect 231 164 232 165
rect 212 164 213 165
rect 211 164 212 165
rect 210 164 211 165
rect 209 164 210 165
rect 208 164 209 165
rect 207 164 208 165
rect 206 164 207 165
rect 205 164 206 165
rect 204 164 205 165
rect 203 164 204 165
rect 202 164 203 165
rect 201 164 202 165
rect 200 164 201 165
rect 199 164 200 165
rect 198 164 199 165
rect 197 164 198 165
rect 196 164 197 165
rect 195 164 196 165
rect 194 164 195 165
rect 193 164 194 165
rect 192 164 193 165
rect 191 164 192 165
rect 190 164 191 165
rect 189 164 190 165
rect 188 164 189 165
rect 187 164 188 165
rect 186 164 187 165
rect 185 164 186 165
rect 184 164 185 165
rect 183 164 184 165
rect 182 164 183 165
rect 181 164 182 165
rect 180 164 181 165
rect 179 164 180 165
rect 178 164 179 165
rect 177 164 178 165
rect 176 164 177 165
rect 175 164 176 165
rect 174 164 175 165
rect 173 164 174 165
rect 172 164 173 165
rect 171 164 172 165
rect 170 164 171 165
rect 169 164 170 165
rect 168 164 169 165
rect 167 164 168 165
rect 166 164 167 165
rect 165 164 166 165
rect 164 164 165 165
rect 163 164 164 165
rect 162 164 163 165
rect 161 164 162 165
rect 160 164 161 165
rect 159 164 160 165
rect 158 164 159 165
rect 157 164 158 165
rect 156 164 157 165
rect 155 164 156 165
rect 154 164 155 165
rect 153 164 154 165
rect 152 164 153 165
rect 151 164 152 165
rect 150 164 151 165
rect 149 164 150 165
rect 148 164 149 165
rect 147 164 148 165
rect 146 164 147 165
rect 145 164 146 165
rect 144 164 145 165
rect 143 164 144 165
rect 142 164 143 165
rect 141 164 142 165
rect 106 164 107 165
rect 105 164 106 165
rect 104 164 105 165
rect 103 164 104 165
rect 102 164 103 165
rect 101 164 102 165
rect 100 164 101 165
rect 99 164 100 165
rect 98 164 99 165
rect 97 164 98 165
rect 96 164 97 165
rect 95 164 96 165
rect 94 164 95 165
rect 93 164 94 165
rect 92 164 93 165
rect 91 164 92 165
rect 90 164 91 165
rect 89 164 90 165
rect 88 164 89 165
rect 87 164 88 165
rect 86 164 87 165
rect 85 164 86 165
rect 84 164 85 165
rect 83 164 84 165
rect 82 164 83 165
rect 81 164 82 165
rect 80 164 81 165
rect 79 164 80 165
rect 78 164 79 165
rect 77 164 78 165
rect 76 164 77 165
rect 75 164 76 165
rect 74 164 75 165
rect 73 164 74 165
rect 68 164 69 165
rect 67 164 68 165
rect 66 164 67 165
rect 65 164 66 165
rect 64 164 65 165
rect 63 164 64 165
rect 62 164 63 165
rect 61 164 62 165
rect 60 164 61 165
rect 59 164 60 165
rect 58 164 59 165
rect 57 164 58 165
rect 56 164 57 165
rect 55 164 56 165
rect 54 164 55 165
rect 53 164 54 165
rect 52 164 53 165
rect 51 164 52 165
rect 50 164 51 165
rect 49 164 50 165
rect 48 164 49 165
rect 47 164 48 165
rect 46 164 47 165
rect 45 164 46 165
rect 44 164 45 165
rect 43 164 44 165
rect 42 164 43 165
rect 41 164 42 165
rect 40 164 41 165
rect 39 164 40 165
rect 38 164 39 165
rect 37 164 38 165
rect 36 164 37 165
rect 35 164 36 165
rect 34 164 35 165
rect 33 164 34 165
rect 23 164 24 165
rect 22 164 23 165
rect 21 164 22 165
rect 20 164 21 165
rect 19 164 20 165
rect 18 164 19 165
rect 17 164 18 165
rect 16 164 17 165
rect 15 164 16 165
rect 14 164 15 165
rect 13 164 14 165
rect 12 164 13 165
rect 11 164 12 165
rect 10 164 11 165
rect 9 164 10 165
rect 8 164 9 165
rect 468 165 469 166
rect 467 165 468 166
rect 466 165 467 166
rect 465 165 466 166
rect 464 165 465 166
rect 463 165 464 166
rect 462 165 463 166
rect 461 165 462 166
rect 460 165 461 166
rect 439 165 440 166
rect 438 165 439 166
rect 437 165 438 166
rect 436 165 437 166
rect 435 165 436 166
rect 434 165 435 166
rect 433 165 434 166
rect 406 165 407 166
rect 405 165 406 166
rect 404 165 405 166
rect 403 165 404 166
rect 402 165 403 166
rect 401 165 402 166
rect 400 165 401 166
rect 399 165 400 166
rect 398 165 399 166
rect 397 165 398 166
rect 396 165 397 166
rect 395 165 396 166
rect 279 165 280 166
rect 278 165 279 166
rect 277 165 278 166
rect 276 165 277 166
rect 275 165 276 166
rect 274 165 275 166
rect 273 165 274 166
rect 272 165 273 166
rect 271 165 272 166
rect 270 165 271 166
rect 269 165 270 166
rect 268 165 269 166
rect 267 165 268 166
rect 266 165 267 166
rect 265 165 266 166
rect 264 165 265 166
rect 263 165 264 166
rect 262 165 263 166
rect 261 165 262 166
rect 260 165 261 166
rect 259 165 260 166
rect 258 165 259 166
rect 257 165 258 166
rect 256 165 257 166
rect 255 165 256 166
rect 254 165 255 166
rect 253 165 254 166
rect 252 165 253 166
rect 251 165 252 166
rect 250 165 251 166
rect 249 165 250 166
rect 248 165 249 166
rect 247 165 248 166
rect 246 165 247 166
rect 245 165 246 166
rect 244 165 245 166
rect 243 165 244 166
rect 242 165 243 166
rect 241 165 242 166
rect 240 165 241 166
rect 239 165 240 166
rect 238 165 239 166
rect 237 165 238 166
rect 236 165 237 166
rect 235 165 236 166
rect 234 165 235 166
rect 233 165 234 166
rect 232 165 233 166
rect 231 165 232 166
rect 230 165 231 166
rect 211 165 212 166
rect 210 165 211 166
rect 209 165 210 166
rect 208 165 209 166
rect 207 165 208 166
rect 206 165 207 166
rect 205 165 206 166
rect 204 165 205 166
rect 203 165 204 166
rect 202 165 203 166
rect 201 165 202 166
rect 200 165 201 166
rect 199 165 200 166
rect 198 165 199 166
rect 197 165 198 166
rect 196 165 197 166
rect 195 165 196 166
rect 194 165 195 166
rect 193 165 194 166
rect 192 165 193 166
rect 191 165 192 166
rect 190 165 191 166
rect 189 165 190 166
rect 188 165 189 166
rect 187 165 188 166
rect 186 165 187 166
rect 185 165 186 166
rect 184 165 185 166
rect 183 165 184 166
rect 182 165 183 166
rect 181 165 182 166
rect 180 165 181 166
rect 179 165 180 166
rect 178 165 179 166
rect 177 165 178 166
rect 176 165 177 166
rect 175 165 176 166
rect 174 165 175 166
rect 173 165 174 166
rect 172 165 173 166
rect 171 165 172 166
rect 170 165 171 166
rect 169 165 170 166
rect 168 165 169 166
rect 167 165 168 166
rect 166 165 167 166
rect 165 165 166 166
rect 164 165 165 166
rect 163 165 164 166
rect 162 165 163 166
rect 161 165 162 166
rect 160 165 161 166
rect 159 165 160 166
rect 158 165 159 166
rect 157 165 158 166
rect 156 165 157 166
rect 155 165 156 166
rect 154 165 155 166
rect 153 165 154 166
rect 152 165 153 166
rect 151 165 152 166
rect 150 165 151 166
rect 149 165 150 166
rect 148 165 149 166
rect 147 165 148 166
rect 146 165 147 166
rect 145 165 146 166
rect 144 165 145 166
rect 143 165 144 166
rect 142 165 143 166
rect 141 165 142 166
rect 140 165 141 166
rect 104 165 105 166
rect 103 165 104 166
rect 102 165 103 166
rect 101 165 102 166
rect 100 165 101 166
rect 99 165 100 166
rect 98 165 99 166
rect 97 165 98 166
rect 96 165 97 166
rect 95 165 96 166
rect 94 165 95 166
rect 93 165 94 166
rect 92 165 93 166
rect 91 165 92 166
rect 90 165 91 166
rect 89 165 90 166
rect 88 165 89 166
rect 87 165 88 166
rect 86 165 87 166
rect 85 165 86 166
rect 84 165 85 166
rect 83 165 84 166
rect 82 165 83 166
rect 81 165 82 166
rect 80 165 81 166
rect 79 165 80 166
rect 78 165 79 166
rect 66 165 67 166
rect 65 165 66 166
rect 64 165 65 166
rect 63 165 64 166
rect 62 165 63 166
rect 61 165 62 166
rect 60 165 61 166
rect 59 165 60 166
rect 58 165 59 166
rect 57 165 58 166
rect 56 165 57 166
rect 55 165 56 166
rect 54 165 55 166
rect 53 165 54 166
rect 52 165 53 166
rect 51 165 52 166
rect 50 165 51 166
rect 49 165 50 166
rect 48 165 49 166
rect 47 165 48 166
rect 46 165 47 166
rect 45 165 46 166
rect 44 165 45 166
rect 43 165 44 166
rect 42 165 43 166
rect 41 165 42 166
rect 40 165 41 166
rect 39 165 40 166
rect 38 165 39 166
rect 37 165 38 166
rect 36 165 37 166
rect 35 165 36 166
rect 34 165 35 166
rect 33 165 34 166
rect 23 165 24 166
rect 22 165 23 166
rect 21 165 22 166
rect 20 165 21 166
rect 19 165 20 166
rect 18 165 19 166
rect 17 165 18 166
rect 16 165 17 166
rect 15 165 16 166
rect 14 165 15 166
rect 13 165 14 166
rect 12 165 13 166
rect 11 165 12 166
rect 10 165 11 166
rect 9 165 10 166
rect 8 165 9 166
rect 470 166 471 167
rect 469 166 470 167
rect 468 166 469 167
rect 467 166 468 167
rect 466 166 467 167
rect 465 166 466 167
rect 464 166 465 167
rect 463 166 464 167
rect 462 166 463 167
rect 461 166 462 167
rect 460 166 461 167
rect 439 166 440 167
rect 438 166 439 167
rect 437 166 438 167
rect 436 166 437 167
rect 407 166 408 167
rect 406 166 407 167
rect 405 166 406 167
rect 404 166 405 167
rect 403 166 404 167
rect 402 166 403 167
rect 401 166 402 167
rect 400 166 401 167
rect 399 166 400 167
rect 398 166 399 167
rect 397 166 398 167
rect 396 166 397 167
rect 395 166 396 167
rect 277 166 278 167
rect 276 166 277 167
rect 275 166 276 167
rect 274 166 275 167
rect 273 166 274 167
rect 272 166 273 167
rect 271 166 272 167
rect 270 166 271 167
rect 269 166 270 167
rect 268 166 269 167
rect 267 166 268 167
rect 266 166 267 167
rect 265 166 266 167
rect 264 166 265 167
rect 263 166 264 167
rect 262 166 263 167
rect 261 166 262 167
rect 260 166 261 167
rect 259 166 260 167
rect 258 166 259 167
rect 257 166 258 167
rect 256 166 257 167
rect 255 166 256 167
rect 254 166 255 167
rect 253 166 254 167
rect 252 166 253 167
rect 251 166 252 167
rect 250 166 251 167
rect 249 166 250 167
rect 248 166 249 167
rect 247 166 248 167
rect 246 166 247 167
rect 245 166 246 167
rect 244 166 245 167
rect 243 166 244 167
rect 242 166 243 167
rect 241 166 242 167
rect 240 166 241 167
rect 239 166 240 167
rect 238 166 239 167
rect 237 166 238 167
rect 236 166 237 167
rect 235 166 236 167
rect 234 166 235 167
rect 233 166 234 167
rect 232 166 233 167
rect 231 166 232 167
rect 230 166 231 167
rect 211 166 212 167
rect 210 166 211 167
rect 209 166 210 167
rect 208 166 209 167
rect 207 166 208 167
rect 206 166 207 167
rect 205 166 206 167
rect 204 166 205 167
rect 203 166 204 167
rect 202 166 203 167
rect 201 166 202 167
rect 200 166 201 167
rect 199 166 200 167
rect 198 166 199 167
rect 197 166 198 167
rect 196 166 197 167
rect 195 166 196 167
rect 194 166 195 167
rect 193 166 194 167
rect 192 166 193 167
rect 191 166 192 167
rect 190 166 191 167
rect 189 166 190 167
rect 188 166 189 167
rect 187 166 188 167
rect 186 166 187 167
rect 185 166 186 167
rect 184 166 185 167
rect 183 166 184 167
rect 182 166 183 167
rect 181 166 182 167
rect 180 166 181 167
rect 179 166 180 167
rect 178 166 179 167
rect 177 166 178 167
rect 176 166 177 167
rect 175 166 176 167
rect 174 166 175 167
rect 173 166 174 167
rect 172 166 173 167
rect 171 166 172 167
rect 170 166 171 167
rect 169 166 170 167
rect 168 166 169 167
rect 167 166 168 167
rect 166 166 167 167
rect 165 166 166 167
rect 164 166 165 167
rect 163 166 164 167
rect 162 166 163 167
rect 161 166 162 167
rect 160 166 161 167
rect 159 166 160 167
rect 158 166 159 167
rect 157 166 158 167
rect 156 166 157 167
rect 155 166 156 167
rect 154 166 155 167
rect 153 166 154 167
rect 152 166 153 167
rect 151 166 152 167
rect 150 166 151 167
rect 149 166 150 167
rect 148 166 149 167
rect 147 166 148 167
rect 146 166 147 167
rect 145 166 146 167
rect 144 166 145 167
rect 143 166 144 167
rect 142 166 143 167
rect 141 166 142 167
rect 140 166 141 167
rect 139 166 140 167
rect 101 166 102 167
rect 100 166 101 167
rect 99 166 100 167
rect 98 166 99 167
rect 97 166 98 167
rect 96 166 97 167
rect 95 166 96 167
rect 94 166 95 167
rect 93 166 94 167
rect 92 166 93 167
rect 91 166 92 167
rect 90 166 91 167
rect 89 166 90 167
rect 88 166 89 167
rect 87 166 88 167
rect 86 166 87 167
rect 85 166 86 167
rect 84 166 85 167
rect 83 166 84 167
rect 82 166 83 167
rect 64 166 65 167
rect 63 166 64 167
rect 62 166 63 167
rect 61 166 62 167
rect 60 166 61 167
rect 59 166 60 167
rect 58 166 59 167
rect 57 166 58 167
rect 56 166 57 167
rect 55 166 56 167
rect 54 166 55 167
rect 53 166 54 167
rect 52 166 53 167
rect 51 166 52 167
rect 50 166 51 167
rect 49 166 50 167
rect 48 166 49 167
rect 47 166 48 167
rect 46 166 47 167
rect 45 166 46 167
rect 44 166 45 167
rect 43 166 44 167
rect 42 166 43 167
rect 41 166 42 167
rect 40 166 41 167
rect 39 166 40 167
rect 38 166 39 167
rect 37 166 38 167
rect 36 166 37 167
rect 35 166 36 167
rect 34 166 35 167
rect 33 166 34 167
rect 23 166 24 167
rect 22 166 23 167
rect 21 166 22 167
rect 20 166 21 167
rect 19 166 20 167
rect 18 166 19 167
rect 17 166 18 167
rect 16 166 17 167
rect 15 166 16 167
rect 14 166 15 167
rect 13 166 14 167
rect 12 166 13 167
rect 11 166 12 167
rect 10 166 11 167
rect 9 166 10 167
rect 8 166 9 167
rect 473 167 474 168
rect 472 167 473 168
rect 471 167 472 168
rect 470 167 471 168
rect 469 167 470 168
rect 468 167 469 168
rect 467 167 468 168
rect 466 167 467 168
rect 465 167 466 168
rect 464 167 465 168
rect 463 167 464 168
rect 462 167 463 168
rect 461 167 462 168
rect 460 167 461 168
rect 439 167 440 168
rect 438 167 439 168
rect 437 167 438 168
rect 409 167 410 168
rect 408 167 409 168
rect 407 167 408 168
rect 406 167 407 168
rect 405 167 406 168
rect 404 167 405 168
rect 403 167 404 168
rect 402 167 403 168
rect 401 167 402 168
rect 400 167 401 168
rect 399 167 400 168
rect 398 167 399 168
rect 397 167 398 168
rect 396 167 397 168
rect 395 167 396 168
rect 276 167 277 168
rect 275 167 276 168
rect 274 167 275 168
rect 273 167 274 168
rect 272 167 273 168
rect 271 167 272 168
rect 270 167 271 168
rect 269 167 270 168
rect 268 167 269 168
rect 267 167 268 168
rect 266 167 267 168
rect 265 167 266 168
rect 264 167 265 168
rect 263 167 264 168
rect 262 167 263 168
rect 261 167 262 168
rect 260 167 261 168
rect 259 167 260 168
rect 258 167 259 168
rect 257 167 258 168
rect 256 167 257 168
rect 255 167 256 168
rect 254 167 255 168
rect 253 167 254 168
rect 252 167 253 168
rect 251 167 252 168
rect 250 167 251 168
rect 249 167 250 168
rect 248 167 249 168
rect 247 167 248 168
rect 246 167 247 168
rect 245 167 246 168
rect 244 167 245 168
rect 243 167 244 168
rect 242 167 243 168
rect 241 167 242 168
rect 240 167 241 168
rect 239 167 240 168
rect 238 167 239 168
rect 237 167 238 168
rect 236 167 237 168
rect 235 167 236 168
rect 234 167 235 168
rect 233 167 234 168
rect 232 167 233 168
rect 231 167 232 168
rect 230 167 231 168
rect 229 167 230 168
rect 210 167 211 168
rect 209 167 210 168
rect 208 167 209 168
rect 207 167 208 168
rect 206 167 207 168
rect 205 167 206 168
rect 204 167 205 168
rect 203 167 204 168
rect 202 167 203 168
rect 201 167 202 168
rect 200 167 201 168
rect 199 167 200 168
rect 198 167 199 168
rect 197 167 198 168
rect 196 167 197 168
rect 195 167 196 168
rect 194 167 195 168
rect 193 167 194 168
rect 192 167 193 168
rect 191 167 192 168
rect 190 167 191 168
rect 189 167 190 168
rect 188 167 189 168
rect 187 167 188 168
rect 186 167 187 168
rect 185 167 186 168
rect 184 167 185 168
rect 183 167 184 168
rect 182 167 183 168
rect 181 167 182 168
rect 180 167 181 168
rect 179 167 180 168
rect 178 167 179 168
rect 177 167 178 168
rect 176 167 177 168
rect 175 167 176 168
rect 174 167 175 168
rect 173 167 174 168
rect 172 167 173 168
rect 171 167 172 168
rect 170 167 171 168
rect 169 167 170 168
rect 168 167 169 168
rect 167 167 168 168
rect 166 167 167 168
rect 165 167 166 168
rect 164 167 165 168
rect 163 167 164 168
rect 162 167 163 168
rect 161 167 162 168
rect 160 167 161 168
rect 159 167 160 168
rect 158 167 159 168
rect 157 167 158 168
rect 156 167 157 168
rect 155 167 156 168
rect 154 167 155 168
rect 153 167 154 168
rect 152 167 153 168
rect 151 167 152 168
rect 150 167 151 168
rect 149 167 150 168
rect 148 167 149 168
rect 147 167 148 168
rect 146 167 147 168
rect 145 167 146 168
rect 144 167 145 168
rect 143 167 144 168
rect 142 167 143 168
rect 141 167 142 168
rect 140 167 141 168
rect 139 167 140 168
rect 138 167 139 168
rect 137 167 138 168
rect 97 167 98 168
rect 96 167 97 168
rect 95 167 96 168
rect 94 167 95 168
rect 93 167 94 168
rect 92 167 93 168
rect 91 167 92 168
rect 90 167 91 168
rect 89 167 90 168
rect 88 167 89 168
rect 63 167 64 168
rect 62 167 63 168
rect 61 167 62 168
rect 60 167 61 168
rect 59 167 60 168
rect 58 167 59 168
rect 57 167 58 168
rect 56 167 57 168
rect 55 167 56 168
rect 54 167 55 168
rect 53 167 54 168
rect 52 167 53 168
rect 51 167 52 168
rect 50 167 51 168
rect 49 167 50 168
rect 48 167 49 168
rect 47 167 48 168
rect 46 167 47 168
rect 45 167 46 168
rect 44 167 45 168
rect 43 167 44 168
rect 42 167 43 168
rect 41 167 42 168
rect 40 167 41 168
rect 39 167 40 168
rect 38 167 39 168
rect 37 167 38 168
rect 36 167 37 168
rect 35 167 36 168
rect 34 167 35 168
rect 33 167 34 168
rect 23 167 24 168
rect 22 167 23 168
rect 21 167 22 168
rect 20 167 21 168
rect 19 167 20 168
rect 18 167 19 168
rect 17 167 18 168
rect 16 167 17 168
rect 15 167 16 168
rect 14 167 15 168
rect 13 167 14 168
rect 12 167 13 168
rect 11 167 12 168
rect 10 167 11 168
rect 9 167 10 168
rect 475 168 476 169
rect 474 168 475 169
rect 473 168 474 169
rect 472 168 473 169
rect 471 168 472 169
rect 470 168 471 169
rect 469 168 470 169
rect 468 168 469 169
rect 467 168 468 169
rect 466 168 467 169
rect 465 168 466 169
rect 464 168 465 169
rect 463 168 464 169
rect 461 168 462 169
rect 460 168 461 169
rect 439 168 440 169
rect 438 168 439 169
rect 437 168 438 169
rect 410 168 411 169
rect 409 168 410 169
rect 408 168 409 169
rect 407 168 408 169
rect 406 168 407 169
rect 405 168 406 169
rect 404 168 405 169
rect 403 168 404 169
rect 402 168 403 169
rect 401 168 402 169
rect 400 168 401 169
rect 399 168 400 169
rect 398 168 399 169
rect 397 168 398 169
rect 396 168 397 169
rect 275 168 276 169
rect 274 168 275 169
rect 273 168 274 169
rect 272 168 273 169
rect 271 168 272 169
rect 270 168 271 169
rect 269 168 270 169
rect 268 168 269 169
rect 267 168 268 169
rect 266 168 267 169
rect 265 168 266 169
rect 264 168 265 169
rect 263 168 264 169
rect 262 168 263 169
rect 261 168 262 169
rect 260 168 261 169
rect 259 168 260 169
rect 258 168 259 169
rect 257 168 258 169
rect 256 168 257 169
rect 255 168 256 169
rect 254 168 255 169
rect 253 168 254 169
rect 252 168 253 169
rect 251 168 252 169
rect 250 168 251 169
rect 249 168 250 169
rect 248 168 249 169
rect 247 168 248 169
rect 246 168 247 169
rect 245 168 246 169
rect 244 168 245 169
rect 243 168 244 169
rect 242 168 243 169
rect 241 168 242 169
rect 240 168 241 169
rect 239 168 240 169
rect 238 168 239 169
rect 237 168 238 169
rect 236 168 237 169
rect 235 168 236 169
rect 234 168 235 169
rect 233 168 234 169
rect 232 168 233 169
rect 231 168 232 169
rect 230 168 231 169
rect 229 168 230 169
rect 210 168 211 169
rect 209 168 210 169
rect 208 168 209 169
rect 207 168 208 169
rect 206 168 207 169
rect 205 168 206 169
rect 204 168 205 169
rect 203 168 204 169
rect 202 168 203 169
rect 201 168 202 169
rect 200 168 201 169
rect 199 168 200 169
rect 198 168 199 169
rect 197 168 198 169
rect 196 168 197 169
rect 195 168 196 169
rect 194 168 195 169
rect 193 168 194 169
rect 192 168 193 169
rect 191 168 192 169
rect 190 168 191 169
rect 189 168 190 169
rect 188 168 189 169
rect 187 168 188 169
rect 186 168 187 169
rect 185 168 186 169
rect 184 168 185 169
rect 183 168 184 169
rect 182 168 183 169
rect 181 168 182 169
rect 180 168 181 169
rect 179 168 180 169
rect 178 168 179 169
rect 177 168 178 169
rect 176 168 177 169
rect 175 168 176 169
rect 174 168 175 169
rect 173 168 174 169
rect 172 168 173 169
rect 171 168 172 169
rect 170 168 171 169
rect 169 168 170 169
rect 168 168 169 169
rect 167 168 168 169
rect 166 168 167 169
rect 165 168 166 169
rect 164 168 165 169
rect 163 168 164 169
rect 162 168 163 169
rect 161 168 162 169
rect 160 168 161 169
rect 159 168 160 169
rect 158 168 159 169
rect 157 168 158 169
rect 156 168 157 169
rect 155 168 156 169
rect 154 168 155 169
rect 153 168 154 169
rect 152 168 153 169
rect 151 168 152 169
rect 150 168 151 169
rect 149 168 150 169
rect 148 168 149 169
rect 147 168 148 169
rect 146 168 147 169
rect 145 168 146 169
rect 144 168 145 169
rect 143 168 144 169
rect 142 168 143 169
rect 141 168 142 169
rect 140 168 141 169
rect 139 168 140 169
rect 138 168 139 169
rect 137 168 138 169
rect 136 168 137 169
rect 62 168 63 169
rect 61 168 62 169
rect 60 168 61 169
rect 59 168 60 169
rect 58 168 59 169
rect 57 168 58 169
rect 56 168 57 169
rect 55 168 56 169
rect 54 168 55 169
rect 53 168 54 169
rect 52 168 53 169
rect 51 168 52 169
rect 50 168 51 169
rect 49 168 50 169
rect 48 168 49 169
rect 47 168 48 169
rect 46 168 47 169
rect 45 168 46 169
rect 44 168 45 169
rect 43 168 44 169
rect 42 168 43 169
rect 41 168 42 169
rect 40 168 41 169
rect 39 168 40 169
rect 38 168 39 169
rect 37 168 38 169
rect 36 168 37 169
rect 35 168 36 169
rect 34 168 35 169
rect 33 168 34 169
rect 23 168 24 169
rect 22 168 23 169
rect 21 168 22 169
rect 20 168 21 169
rect 19 168 20 169
rect 18 168 19 169
rect 17 168 18 169
rect 16 168 17 169
rect 15 168 16 169
rect 14 168 15 169
rect 13 168 14 169
rect 12 168 13 169
rect 11 168 12 169
rect 10 168 11 169
rect 9 168 10 169
rect 478 169 479 170
rect 477 169 478 170
rect 476 169 477 170
rect 475 169 476 170
rect 474 169 475 170
rect 473 169 474 170
rect 472 169 473 170
rect 471 169 472 170
rect 470 169 471 170
rect 469 169 470 170
rect 468 169 469 170
rect 467 169 468 170
rect 466 169 467 170
rect 460 169 461 170
rect 439 169 440 170
rect 438 169 439 170
rect 437 169 438 170
rect 411 169 412 170
rect 410 169 411 170
rect 409 169 410 170
rect 408 169 409 170
rect 407 169 408 170
rect 406 169 407 170
rect 405 169 406 170
rect 404 169 405 170
rect 403 169 404 170
rect 402 169 403 170
rect 401 169 402 170
rect 400 169 401 170
rect 399 169 400 170
rect 398 169 399 170
rect 274 169 275 170
rect 273 169 274 170
rect 272 169 273 170
rect 271 169 272 170
rect 270 169 271 170
rect 269 169 270 170
rect 268 169 269 170
rect 267 169 268 170
rect 266 169 267 170
rect 265 169 266 170
rect 264 169 265 170
rect 263 169 264 170
rect 262 169 263 170
rect 261 169 262 170
rect 260 169 261 170
rect 259 169 260 170
rect 258 169 259 170
rect 257 169 258 170
rect 256 169 257 170
rect 255 169 256 170
rect 254 169 255 170
rect 253 169 254 170
rect 252 169 253 170
rect 251 169 252 170
rect 250 169 251 170
rect 249 169 250 170
rect 248 169 249 170
rect 247 169 248 170
rect 246 169 247 170
rect 245 169 246 170
rect 244 169 245 170
rect 243 169 244 170
rect 242 169 243 170
rect 241 169 242 170
rect 240 169 241 170
rect 239 169 240 170
rect 238 169 239 170
rect 237 169 238 170
rect 236 169 237 170
rect 235 169 236 170
rect 234 169 235 170
rect 233 169 234 170
rect 232 169 233 170
rect 231 169 232 170
rect 230 169 231 170
rect 229 169 230 170
rect 228 169 229 170
rect 209 169 210 170
rect 208 169 209 170
rect 207 169 208 170
rect 206 169 207 170
rect 205 169 206 170
rect 204 169 205 170
rect 203 169 204 170
rect 202 169 203 170
rect 201 169 202 170
rect 200 169 201 170
rect 199 169 200 170
rect 198 169 199 170
rect 197 169 198 170
rect 196 169 197 170
rect 195 169 196 170
rect 194 169 195 170
rect 193 169 194 170
rect 192 169 193 170
rect 191 169 192 170
rect 190 169 191 170
rect 189 169 190 170
rect 188 169 189 170
rect 187 169 188 170
rect 186 169 187 170
rect 185 169 186 170
rect 184 169 185 170
rect 183 169 184 170
rect 182 169 183 170
rect 181 169 182 170
rect 180 169 181 170
rect 179 169 180 170
rect 178 169 179 170
rect 177 169 178 170
rect 176 169 177 170
rect 175 169 176 170
rect 174 169 175 170
rect 173 169 174 170
rect 172 169 173 170
rect 171 169 172 170
rect 170 169 171 170
rect 169 169 170 170
rect 168 169 169 170
rect 167 169 168 170
rect 166 169 167 170
rect 165 169 166 170
rect 164 169 165 170
rect 163 169 164 170
rect 162 169 163 170
rect 161 169 162 170
rect 160 169 161 170
rect 159 169 160 170
rect 158 169 159 170
rect 157 169 158 170
rect 156 169 157 170
rect 155 169 156 170
rect 154 169 155 170
rect 153 169 154 170
rect 152 169 153 170
rect 151 169 152 170
rect 150 169 151 170
rect 149 169 150 170
rect 148 169 149 170
rect 147 169 148 170
rect 146 169 147 170
rect 145 169 146 170
rect 144 169 145 170
rect 143 169 144 170
rect 142 169 143 170
rect 141 169 142 170
rect 140 169 141 170
rect 139 169 140 170
rect 138 169 139 170
rect 137 169 138 170
rect 136 169 137 170
rect 135 169 136 170
rect 61 169 62 170
rect 60 169 61 170
rect 59 169 60 170
rect 58 169 59 170
rect 57 169 58 170
rect 56 169 57 170
rect 55 169 56 170
rect 54 169 55 170
rect 53 169 54 170
rect 52 169 53 170
rect 51 169 52 170
rect 50 169 51 170
rect 49 169 50 170
rect 48 169 49 170
rect 47 169 48 170
rect 46 169 47 170
rect 45 169 46 170
rect 44 169 45 170
rect 43 169 44 170
rect 42 169 43 170
rect 41 169 42 170
rect 40 169 41 170
rect 39 169 40 170
rect 38 169 39 170
rect 37 169 38 170
rect 36 169 37 170
rect 35 169 36 170
rect 34 169 35 170
rect 33 169 34 170
rect 23 169 24 170
rect 22 169 23 170
rect 21 169 22 170
rect 20 169 21 170
rect 19 169 20 170
rect 18 169 19 170
rect 17 169 18 170
rect 16 169 17 170
rect 15 169 16 170
rect 14 169 15 170
rect 13 169 14 170
rect 12 169 13 170
rect 11 169 12 170
rect 10 169 11 170
rect 9 169 10 170
rect 481 170 482 171
rect 480 170 481 171
rect 479 170 480 171
rect 478 170 479 171
rect 477 170 478 171
rect 476 170 477 171
rect 475 170 476 171
rect 474 170 475 171
rect 473 170 474 171
rect 472 170 473 171
rect 471 170 472 171
rect 470 170 471 171
rect 469 170 470 171
rect 439 170 440 171
rect 438 170 439 171
rect 437 170 438 171
rect 412 170 413 171
rect 411 170 412 171
rect 410 170 411 171
rect 409 170 410 171
rect 408 170 409 171
rect 407 170 408 171
rect 406 170 407 171
rect 405 170 406 171
rect 404 170 405 171
rect 403 170 404 171
rect 402 170 403 171
rect 401 170 402 171
rect 400 170 401 171
rect 399 170 400 171
rect 272 170 273 171
rect 271 170 272 171
rect 270 170 271 171
rect 269 170 270 171
rect 268 170 269 171
rect 267 170 268 171
rect 266 170 267 171
rect 265 170 266 171
rect 264 170 265 171
rect 263 170 264 171
rect 262 170 263 171
rect 261 170 262 171
rect 260 170 261 171
rect 259 170 260 171
rect 258 170 259 171
rect 257 170 258 171
rect 256 170 257 171
rect 255 170 256 171
rect 254 170 255 171
rect 253 170 254 171
rect 252 170 253 171
rect 251 170 252 171
rect 250 170 251 171
rect 249 170 250 171
rect 248 170 249 171
rect 247 170 248 171
rect 246 170 247 171
rect 245 170 246 171
rect 244 170 245 171
rect 243 170 244 171
rect 242 170 243 171
rect 241 170 242 171
rect 240 170 241 171
rect 239 170 240 171
rect 238 170 239 171
rect 237 170 238 171
rect 236 170 237 171
rect 235 170 236 171
rect 234 170 235 171
rect 233 170 234 171
rect 232 170 233 171
rect 231 170 232 171
rect 230 170 231 171
rect 229 170 230 171
rect 228 170 229 171
rect 209 170 210 171
rect 208 170 209 171
rect 207 170 208 171
rect 206 170 207 171
rect 205 170 206 171
rect 204 170 205 171
rect 203 170 204 171
rect 202 170 203 171
rect 201 170 202 171
rect 200 170 201 171
rect 199 170 200 171
rect 198 170 199 171
rect 197 170 198 171
rect 196 170 197 171
rect 195 170 196 171
rect 194 170 195 171
rect 193 170 194 171
rect 192 170 193 171
rect 191 170 192 171
rect 190 170 191 171
rect 189 170 190 171
rect 188 170 189 171
rect 187 170 188 171
rect 186 170 187 171
rect 185 170 186 171
rect 184 170 185 171
rect 183 170 184 171
rect 182 170 183 171
rect 181 170 182 171
rect 180 170 181 171
rect 179 170 180 171
rect 178 170 179 171
rect 177 170 178 171
rect 176 170 177 171
rect 175 170 176 171
rect 174 170 175 171
rect 173 170 174 171
rect 172 170 173 171
rect 171 170 172 171
rect 170 170 171 171
rect 169 170 170 171
rect 168 170 169 171
rect 167 170 168 171
rect 166 170 167 171
rect 165 170 166 171
rect 164 170 165 171
rect 163 170 164 171
rect 162 170 163 171
rect 161 170 162 171
rect 160 170 161 171
rect 159 170 160 171
rect 158 170 159 171
rect 157 170 158 171
rect 156 170 157 171
rect 155 170 156 171
rect 154 170 155 171
rect 153 170 154 171
rect 152 170 153 171
rect 151 170 152 171
rect 150 170 151 171
rect 149 170 150 171
rect 148 170 149 171
rect 147 170 148 171
rect 146 170 147 171
rect 145 170 146 171
rect 144 170 145 171
rect 143 170 144 171
rect 142 170 143 171
rect 141 170 142 171
rect 140 170 141 171
rect 139 170 140 171
rect 138 170 139 171
rect 137 170 138 171
rect 136 170 137 171
rect 135 170 136 171
rect 134 170 135 171
rect 133 170 134 171
rect 60 170 61 171
rect 59 170 60 171
rect 58 170 59 171
rect 57 170 58 171
rect 56 170 57 171
rect 55 170 56 171
rect 54 170 55 171
rect 53 170 54 171
rect 52 170 53 171
rect 51 170 52 171
rect 50 170 51 171
rect 49 170 50 171
rect 48 170 49 171
rect 47 170 48 171
rect 46 170 47 171
rect 45 170 46 171
rect 44 170 45 171
rect 43 170 44 171
rect 42 170 43 171
rect 41 170 42 171
rect 40 170 41 171
rect 39 170 40 171
rect 38 170 39 171
rect 37 170 38 171
rect 36 170 37 171
rect 35 170 36 171
rect 34 170 35 171
rect 33 170 34 171
rect 23 170 24 171
rect 22 170 23 171
rect 21 170 22 171
rect 20 170 21 171
rect 19 170 20 171
rect 18 170 19 171
rect 17 170 18 171
rect 16 170 17 171
rect 15 170 16 171
rect 14 170 15 171
rect 13 170 14 171
rect 12 170 13 171
rect 11 170 12 171
rect 10 170 11 171
rect 9 170 10 171
rect 481 171 482 172
rect 480 171 481 172
rect 479 171 480 172
rect 478 171 479 172
rect 477 171 478 172
rect 476 171 477 172
rect 475 171 476 172
rect 474 171 475 172
rect 473 171 474 172
rect 472 171 473 172
rect 471 171 472 172
rect 439 171 440 172
rect 438 171 439 172
rect 413 171 414 172
rect 412 171 413 172
rect 411 171 412 172
rect 410 171 411 172
rect 409 171 410 172
rect 408 171 409 172
rect 407 171 408 172
rect 406 171 407 172
rect 405 171 406 172
rect 404 171 405 172
rect 403 171 404 172
rect 402 171 403 172
rect 401 171 402 172
rect 400 171 401 172
rect 271 171 272 172
rect 270 171 271 172
rect 269 171 270 172
rect 268 171 269 172
rect 267 171 268 172
rect 266 171 267 172
rect 265 171 266 172
rect 264 171 265 172
rect 263 171 264 172
rect 262 171 263 172
rect 261 171 262 172
rect 260 171 261 172
rect 259 171 260 172
rect 258 171 259 172
rect 257 171 258 172
rect 256 171 257 172
rect 255 171 256 172
rect 254 171 255 172
rect 253 171 254 172
rect 252 171 253 172
rect 251 171 252 172
rect 250 171 251 172
rect 249 171 250 172
rect 248 171 249 172
rect 247 171 248 172
rect 246 171 247 172
rect 245 171 246 172
rect 244 171 245 172
rect 243 171 244 172
rect 242 171 243 172
rect 241 171 242 172
rect 240 171 241 172
rect 239 171 240 172
rect 238 171 239 172
rect 237 171 238 172
rect 236 171 237 172
rect 235 171 236 172
rect 234 171 235 172
rect 233 171 234 172
rect 232 171 233 172
rect 231 171 232 172
rect 230 171 231 172
rect 229 171 230 172
rect 228 171 229 172
rect 227 171 228 172
rect 208 171 209 172
rect 207 171 208 172
rect 206 171 207 172
rect 205 171 206 172
rect 204 171 205 172
rect 203 171 204 172
rect 202 171 203 172
rect 201 171 202 172
rect 200 171 201 172
rect 199 171 200 172
rect 198 171 199 172
rect 197 171 198 172
rect 196 171 197 172
rect 195 171 196 172
rect 194 171 195 172
rect 193 171 194 172
rect 192 171 193 172
rect 191 171 192 172
rect 190 171 191 172
rect 189 171 190 172
rect 188 171 189 172
rect 187 171 188 172
rect 186 171 187 172
rect 185 171 186 172
rect 184 171 185 172
rect 183 171 184 172
rect 182 171 183 172
rect 181 171 182 172
rect 180 171 181 172
rect 179 171 180 172
rect 178 171 179 172
rect 177 171 178 172
rect 176 171 177 172
rect 175 171 176 172
rect 174 171 175 172
rect 173 171 174 172
rect 172 171 173 172
rect 171 171 172 172
rect 170 171 171 172
rect 169 171 170 172
rect 168 171 169 172
rect 167 171 168 172
rect 166 171 167 172
rect 165 171 166 172
rect 164 171 165 172
rect 163 171 164 172
rect 162 171 163 172
rect 161 171 162 172
rect 160 171 161 172
rect 159 171 160 172
rect 158 171 159 172
rect 157 171 158 172
rect 156 171 157 172
rect 155 171 156 172
rect 154 171 155 172
rect 153 171 154 172
rect 152 171 153 172
rect 151 171 152 172
rect 150 171 151 172
rect 149 171 150 172
rect 148 171 149 172
rect 147 171 148 172
rect 146 171 147 172
rect 145 171 146 172
rect 144 171 145 172
rect 143 171 144 172
rect 142 171 143 172
rect 141 171 142 172
rect 140 171 141 172
rect 139 171 140 172
rect 138 171 139 172
rect 137 171 138 172
rect 136 171 137 172
rect 135 171 136 172
rect 134 171 135 172
rect 133 171 134 172
rect 132 171 133 172
rect 59 171 60 172
rect 58 171 59 172
rect 57 171 58 172
rect 56 171 57 172
rect 55 171 56 172
rect 54 171 55 172
rect 53 171 54 172
rect 52 171 53 172
rect 51 171 52 172
rect 50 171 51 172
rect 49 171 50 172
rect 48 171 49 172
rect 47 171 48 172
rect 46 171 47 172
rect 45 171 46 172
rect 44 171 45 172
rect 43 171 44 172
rect 42 171 43 172
rect 41 171 42 172
rect 40 171 41 172
rect 39 171 40 172
rect 38 171 39 172
rect 37 171 38 172
rect 36 171 37 172
rect 35 171 36 172
rect 34 171 35 172
rect 22 171 23 172
rect 21 171 22 172
rect 20 171 21 172
rect 19 171 20 172
rect 18 171 19 172
rect 17 171 18 172
rect 16 171 17 172
rect 15 171 16 172
rect 14 171 15 172
rect 13 171 14 172
rect 12 171 13 172
rect 11 171 12 172
rect 10 171 11 172
rect 480 172 481 173
rect 479 172 480 173
rect 478 172 479 173
rect 477 172 478 173
rect 476 172 477 173
rect 475 172 476 173
rect 474 172 475 173
rect 414 172 415 173
rect 413 172 414 173
rect 412 172 413 173
rect 411 172 412 173
rect 410 172 411 173
rect 409 172 410 173
rect 408 172 409 173
rect 407 172 408 173
rect 406 172 407 173
rect 405 172 406 173
rect 404 172 405 173
rect 403 172 404 173
rect 402 172 403 173
rect 401 172 402 173
rect 270 172 271 173
rect 269 172 270 173
rect 268 172 269 173
rect 267 172 268 173
rect 266 172 267 173
rect 265 172 266 173
rect 264 172 265 173
rect 263 172 264 173
rect 262 172 263 173
rect 261 172 262 173
rect 260 172 261 173
rect 259 172 260 173
rect 258 172 259 173
rect 257 172 258 173
rect 256 172 257 173
rect 255 172 256 173
rect 254 172 255 173
rect 253 172 254 173
rect 252 172 253 173
rect 251 172 252 173
rect 250 172 251 173
rect 249 172 250 173
rect 248 172 249 173
rect 247 172 248 173
rect 246 172 247 173
rect 245 172 246 173
rect 244 172 245 173
rect 243 172 244 173
rect 242 172 243 173
rect 241 172 242 173
rect 240 172 241 173
rect 239 172 240 173
rect 238 172 239 173
rect 237 172 238 173
rect 236 172 237 173
rect 235 172 236 173
rect 234 172 235 173
rect 233 172 234 173
rect 232 172 233 173
rect 231 172 232 173
rect 230 172 231 173
rect 229 172 230 173
rect 228 172 229 173
rect 227 172 228 173
rect 226 172 227 173
rect 208 172 209 173
rect 207 172 208 173
rect 206 172 207 173
rect 205 172 206 173
rect 204 172 205 173
rect 203 172 204 173
rect 202 172 203 173
rect 201 172 202 173
rect 200 172 201 173
rect 199 172 200 173
rect 198 172 199 173
rect 197 172 198 173
rect 196 172 197 173
rect 195 172 196 173
rect 194 172 195 173
rect 193 172 194 173
rect 192 172 193 173
rect 191 172 192 173
rect 190 172 191 173
rect 189 172 190 173
rect 188 172 189 173
rect 187 172 188 173
rect 186 172 187 173
rect 185 172 186 173
rect 184 172 185 173
rect 183 172 184 173
rect 182 172 183 173
rect 181 172 182 173
rect 180 172 181 173
rect 179 172 180 173
rect 178 172 179 173
rect 177 172 178 173
rect 176 172 177 173
rect 175 172 176 173
rect 174 172 175 173
rect 173 172 174 173
rect 172 172 173 173
rect 171 172 172 173
rect 170 172 171 173
rect 169 172 170 173
rect 168 172 169 173
rect 167 172 168 173
rect 166 172 167 173
rect 165 172 166 173
rect 164 172 165 173
rect 163 172 164 173
rect 162 172 163 173
rect 161 172 162 173
rect 160 172 161 173
rect 159 172 160 173
rect 158 172 159 173
rect 157 172 158 173
rect 156 172 157 173
rect 155 172 156 173
rect 154 172 155 173
rect 153 172 154 173
rect 152 172 153 173
rect 151 172 152 173
rect 150 172 151 173
rect 149 172 150 173
rect 148 172 149 173
rect 147 172 148 173
rect 146 172 147 173
rect 145 172 146 173
rect 144 172 145 173
rect 143 172 144 173
rect 142 172 143 173
rect 141 172 142 173
rect 140 172 141 173
rect 139 172 140 173
rect 138 172 139 173
rect 137 172 138 173
rect 136 172 137 173
rect 135 172 136 173
rect 134 172 135 173
rect 133 172 134 173
rect 132 172 133 173
rect 131 172 132 173
rect 130 172 131 173
rect 58 172 59 173
rect 57 172 58 173
rect 56 172 57 173
rect 55 172 56 173
rect 54 172 55 173
rect 53 172 54 173
rect 52 172 53 173
rect 51 172 52 173
rect 50 172 51 173
rect 49 172 50 173
rect 48 172 49 173
rect 47 172 48 173
rect 46 172 47 173
rect 45 172 46 173
rect 44 172 45 173
rect 43 172 44 173
rect 42 172 43 173
rect 41 172 42 173
rect 40 172 41 173
rect 39 172 40 173
rect 38 172 39 173
rect 37 172 38 173
rect 36 172 37 173
rect 35 172 36 173
rect 34 172 35 173
rect 22 172 23 173
rect 21 172 22 173
rect 20 172 21 173
rect 19 172 20 173
rect 18 172 19 173
rect 17 172 18 173
rect 16 172 17 173
rect 15 172 16 173
rect 14 172 15 173
rect 13 172 14 173
rect 12 172 13 173
rect 11 172 12 173
rect 10 172 11 173
rect 478 173 479 174
rect 477 173 478 174
rect 476 173 477 174
rect 475 173 476 174
rect 474 173 475 174
rect 416 173 417 174
rect 415 173 416 174
rect 414 173 415 174
rect 413 173 414 174
rect 412 173 413 174
rect 411 173 412 174
rect 410 173 411 174
rect 409 173 410 174
rect 408 173 409 174
rect 407 173 408 174
rect 406 173 407 174
rect 405 173 406 174
rect 404 173 405 174
rect 403 173 404 174
rect 402 173 403 174
rect 269 173 270 174
rect 268 173 269 174
rect 267 173 268 174
rect 266 173 267 174
rect 265 173 266 174
rect 264 173 265 174
rect 263 173 264 174
rect 262 173 263 174
rect 261 173 262 174
rect 260 173 261 174
rect 259 173 260 174
rect 258 173 259 174
rect 257 173 258 174
rect 256 173 257 174
rect 255 173 256 174
rect 254 173 255 174
rect 253 173 254 174
rect 252 173 253 174
rect 251 173 252 174
rect 250 173 251 174
rect 249 173 250 174
rect 248 173 249 174
rect 247 173 248 174
rect 246 173 247 174
rect 245 173 246 174
rect 244 173 245 174
rect 243 173 244 174
rect 242 173 243 174
rect 241 173 242 174
rect 240 173 241 174
rect 239 173 240 174
rect 238 173 239 174
rect 237 173 238 174
rect 236 173 237 174
rect 235 173 236 174
rect 234 173 235 174
rect 233 173 234 174
rect 232 173 233 174
rect 231 173 232 174
rect 230 173 231 174
rect 229 173 230 174
rect 228 173 229 174
rect 227 173 228 174
rect 226 173 227 174
rect 207 173 208 174
rect 206 173 207 174
rect 205 173 206 174
rect 204 173 205 174
rect 203 173 204 174
rect 202 173 203 174
rect 201 173 202 174
rect 200 173 201 174
rect 199 173 200 174
rect 198 173 199 174
rect 197 173 198 174
rect 196 173 197 174
rect 195 173 196 174
rect 194 173 195 174
rect 193 173 194 174
rect 192 173 193 174
rect 191 173 192 174
rect 190 173 191 174
rect 189 173 190 174
rect 188 173 189 174
rect 187 173 188 174
rect 186 173 187 174
rect 185 173 186 174
rect 184 173 185 174
rect 183 173 184 174
rect 182 173 183 174
rect 181 173 182 174
rect 180 173 181 174
rect 179 173 180 174
rect 178 173 179 174
rect 177 173 178 174
rect 176 173 177 174
rect 175 173 176 174
rect 174 173 175 174
rect 173 173 174 174
rect 172 173 173 174
rect 171 173 172 174
rect 170 173 171 174
rect 169 173 170 174
rect 168 173 169 174
rect 167 173 168 174
rect 166 173 167 174
rect 165 173 166 174
rect 164 173 165 174
rect 163 173 164 174
rect 162 173 163 174
rect 161 173 162 174
rect 160 173 161 174
rect 159 173 160 174
rect 158 173 159 174
rect 157 173 158 174
rect 156 173 157 174
rect 155 173 156 174
rect 154 173 155 174
rect 153 173 154 174
rect 152 173 153 174
rect 151 173 152 174
rect 150 173 151 174
rect 149 173 150 174
rect 148 173 149 174
rect 147 173 148 174
rect 146 173 147 174
rect 145 173 146 174
rect 144 173 145 174
rect 143 173 144 174
rect 142 173 143 174
rect 141 173 142 174
rect 140 173 141 174
rect 139 173 140 174
rect 138 173 139 174
rect 137 173 138 174
rect 136 173 137 174
rect 135 173 136 174
rect 134 173 135 174
rect 133 173 134 174
rect 132 173 133 174
rect 131 173 132 174
rect 130 173 131 174
rect 129 173 130 174
rect 128 173 129 174
rect 57 173 58 174
rect 56 173 57 174
rect 55 173 56 174
rect 54 173 55 174
rect 53 173 54 174
rect 52 173 53 174
rect 51 173 52 174
rect 50 173 51 174
rect 49 173 50 174
rect 48 173 49 174
rect 47 173 48 174
rect 46 173 47 174
rect 45 173 46 174
rect 44 173 45 174
rect 43 173 44 174
rect 42 173 43 174
rect 41 173 42 174
rect 40 173 41 174
rect 39 173 40 174
rect 38 173 39 174
rect 37 173 38 174
rect 36 173 37 174
rect 35 173 36 174
rect 34 173 35 174
rect 22 173 23 174
rect 21 173 22 174
rect 20 173 21 174
rect 19 173 20 174
rect 18 173 19 174
rect 17 173 18 174
rect 16 173 17 174
rect 15 173 16 174
rect 14 173 15 174
rect 13 173 14 174
rect 12 173 13 174
rect 11 173 12 174
rect 10 173 11 174
rect 475 174 476 175
rect 474 174 475 175
rect 473 174 474 175
rect 472 174 473 175
rect 471 174 472 175
rect 417 174 418 175
rect 416 174 417 175
rect 415 174 416 175
rect 414 174 415 175
rect 413 174 414 175
rect 412 174 413 175
rect 411 174 412 175
rect 410 174 411 175
rect 409 174 410 175
rect 408 174 409 175
rect 407 174 408 175
rect 406 174 407 175
rect 405 174 406 175
rect 404 174 405 175
rect 403 174 404 175
rect 268 174 269 175
rect 267 174 268 175
rect 266 174 267 175
rect 265 174 266 175
rect 264 174 265 175
rect 263 174 264 175
rect 262 174 263 175
rect 261 174 262 175
rect 260 174 261 175
rect 259 174 260 175
rect 258 174 259 175
rect 257 174 258 175
rect 256 174 257 175
rect 255 174 256 175
rect 254 174 255 175
rect 253 174 254 175
rect 252 174 253 175
rect 251 174 252 175
rect 250 174 251 175
rect 249 174 250 175
rect 248 174 249 175
rect 247 174 248 175
rect 246 174 247 175
rect 245 174 246 175
rect 244 174 245 175
rect 243 174 244 175
rect 242 174 243 175
rect 241 174 242 175
rect 240 174 241 175
rect 239 174 240 175
rect 238 174 239 175
rect 237 174 238 175
rect 236 174 237 175
rect 235 174 236 175
rect 234 174 235 175
rect 233 174 234 175
rect 232 174 233 175
rect 231 174 232 175
rect 230 174 231 175
rect 229 174 230 175
rect 228 174 229 175
rect 227 174 228 175
rect 226 174 227 175
rect 225 174 226 175
rect 206 174 207 175
rect 205 174 206 175
rect 204 174 205 175
rect 203 174 204 175
rect 202 174 203 175
rect 201 174 202 175
rect 200 174 201 175
rect 199 174 200 175
rect 198 174 199 175
rect 197 174 198 175
rect 196 174 197 175
rect 195 174 196 175
rect 194 174 195 175
rect 193 174 194 175
rect 192 174 193 175
rect 191 174 192 175
rect 190 174 191 175
rect 189 174 190 175
rect 188 174 189 175
rect 187 174 188 175
rect 186 174 187 175
rect 185 174 186 175
rect 184 174 185 175
rect 183 174 184 175
rect 182 174 183 175
rect 181 174 182 175
rect 180 174 181 175
rect 179 174 180 175
rect 178 174 179 175
rect 177 174 178 175
rect 176 174 177 175
rect 175 174 176 175
rect 174 174 175 175
rect 173 174 174 175
rect 172 174 173 175
rect 171 174 172 175
rect 170 174 171 175
rect 169 174 170 175
rect 168 174 169 175
rect 167 174 168 175
rect 166 174 167 175
rect 165 174 166 175
rect 164 174 165 175
rect 163 174 164 175
rect 162 174 163 175
rect 161 174 162 175
rect 160 174 161 175
rect 159 174 160 175
rect 158 174 159 175
rect 157 174 158 175
rect 156 174 157 175
rect 155 174 156 175
rect 154 174 155 175
rect 153 174 154 175
rect 152 174 153 175
rect 151 174 152 175
rect 150 174 151 175
rect 149 174 150 175
rect 148 174 149 175
rect 147 174 148 175
rect 146 174 147 175
rect 145 174 146 175
rect 144 174 145 175
rect 143 174 144 175
rect 142 174 143 175
rect 141 174 142 175
rect 140 174 141 175
rect 139 174 140 175
rect 138 174 139 175
rect 137 174 138 175
rect 136 174 137 175
rect 135 174 136 175
rect 134 174 135 175
rect 133 174 134 175
rect 132 174 133 175
rect 131 174 132 175
rect 130 174 131 175
rect 129 174 130 175
rect 128 174 129 175
rect 127 174 128 175
rect 57 174 58 175
rect 56 174 57 175
rect 55 174 56 175
rect 54 174 55 175
rect 53 174 54 175
rect 52 174 53 175
rect 51 174 52 175
rect 50 174 51 175
rect 49 174 50 175
rect 48 174 49 175
rect 47 174 48 175
rect 46 174 47 175
rect 45 174 46 175
rect 44 174 45 175
rect 43 174 44 175
rect 42 174 43 175
rect 41 174 42 175
rect 40 174 41 175
rect 39 174 40 175
rect 38 174 39 175
rect 37 174 38 175
rect 36 174 37 175
rect 35 174 36 175
rect 22 174 23 175
rect 21 174 22 175
rect 20 174 21 175
rect 19 174 20 175
rect 18 174 19 175
rect 17 174 18 175
rect 16 174 17 175
rect 15 174 16 175
rect 14 174 15 175
rect 13 174 14 175
rect 12 174 13 175
rect 11 174 12 175
rect 473 175 474 176
rect 472 175 473 176
rect 471 175 472 176
rect 470 175 471 176
rect 469 175 470 176
rect 460 175 461 176
rect 418 175 419 176
rect 417 175 418 176
rect 416 175 417 176
rect 415 175 416 176
rect 414 175 415 176
rect 413 175 414 176
rect 412 175 413 176
rect 411 175 412 176
rect 410 175 411 176
rect 409 175 410 176
rect 408 175 409 176
rect 407 175 408 176
rect 406 175 407 176
rect 405 175 406 176
rect 267 175 268 176
rect 266 175 267 176
rect 265 175 266 176
rect 264 175 265 176
rect 263 175 264 176
rect 262 175 263 176
rect 261 175 262 176
rect 260 175 261 176
rect 259 175 260 176
rect 258 175 259 176
rect 257 175 258 176
rect 256 175 257 176
rect 255 175 256 176
rect 254 175 255 176
rect 253 175 254 176
rect 252 175 253 176
rect 251 175 252 176
rect 250 175 251 176
rect 249 175 250 176
rect 248 175 249 176
rect 247 175 248 176
rect 246 175 247 176
rect 245 175 246 176
rect 244 175 245 176
rect 243 175 244 176
rect 242 175 243 176
rect 241 175 242 176
rect 240 175 241 176
rect 239 175 240 176
rect 238 175 239 176
rect 237 175 238 176
rect 236 175 237 176
rect 235 175 236 176
rect 234 175 235 176
rect 233 175 234 176
rect 232 175 233 176
rect 231 175 232 176
rect 230 175 231 176
rect 229 175 230 176
rect 228 175 229 176
rect 227 175 228 176
rect 226 175 227 176
rect 225 175 226 176
rect 206 175 207 176
rect 205 175 206 176
rect 204 175 205 176
rect 203 175 204 176
rect 202 175 203 176
rect 201 175 202 176
rect 200 175 201 176
rect 199 175 200 176
rect 198 175 199 176
rect 197 175 198 176
rect 196 175 197 176
rect 195 175 196 176
rect 194 175 195 176
rect 193 175 194 176
rect 192 175 193 176
rect 191 175 192 176
rect 190 175 191 176
rect 189 175 190 176
rect 188 175 189 176
rect 187 175 188 176
rect 186 175 187 176
rect 185 175 186 176
rect 184 175 185 176
rect 183 175 184 176
rect 182 175 183 176
rect 181 175 182 176
rect 180 175 181 176
rect 179 175 180 176
rect 178 175 179 176
rect 177 175 178 176
rect 176 175 177 176
rect 175 175 176 176
rect 174 175 175 176
rect 173 175 174 176
rect 172 175 173 176
rect 171 175 172 176
rect 170 175 171 176
rect 169 175 170 176
rect 168 175 169 176
rect 167 175 168 176
rect 166 175 167 176
rect 165 175 166 176
rect 164 175 165 176
rect 163 175 164 176
rect 162 175 163 176
rect 161 175 162 176
rect 160 175 161 176
rect 159 175 160 176
rect 158 175 159 176
rect 157 175 158 176
rect 156 175 157 176
rect 155 175 156 176
rect 154 175 155 176
rect 153 175 154 176
rect 152 175 153 176
rect 151 175 152 176
rect 150 175 151 176
rect 149 175 150 176
rect 148 175 149 176
rect 147 175 148 176
rect 146 175 147 176
rect 145 175 146 176
rect 144 175 145 176
rect 143 175 144 176
rect 142 175 143 176
rect 141 175 142 176
rect 140 175 141 176
rect 139 175 140 176
rect 138 175 139 176
rect 137 175 138 176
rect 136 175 137 176
rect 135 175 136 176
rect 134 175 135 176
rect 133 175 134 176
rect 132 175 133 176
rect 131 175 132 176
rect 130 175 131 176
rect 129 175 130 176
rect 128 175 129 176
rect 127 175 128 176
rect 126 175 127 176
rect 125 175 126 176
rect 56 175 57 176
rect 55 175 56 176
rect 54 175 55 176
rect 53 175 54 176
rect 52 175 53 176
rect 51 175 52 176
rect 50 175 51 176
rect 49 175 50 176
rect 48 175 49 176
rect 47 175 48 176
rect 46 175 47 176
rect 45 175 46 176
rect 44 175 45 176
rect 43 175 44 176
rect 42 175 43 176
rect 41 175 42 176
rect 40 175 41 176
rect 39 175 40 176
rect 38 175 39 176
rect 37 175 38 176
rect 36 175 37 176
rect 35 175 36 176
rect 23 175 24 176
rect 22 175 23 176
rect 21 175 22 176
rect 20 175 21 176
rect 19 175 20 176
rect 18 175 19 176
rect 17 175 18 176
rect 16 175 17 176
rect 15 175 16 176
rect 14 175 15 176
rect 13 175 14 176
rect 12 175 13 176
rect 11 175 12 176
rect 470 176 471 177
rect 469 176 470 177
rect 468 176 469 177
rect 467 176 468 177
rect 466 176 467 177
rect 460 176 461 177
rect 419 176 420 177
rect 418 176 419 177
rect 417 176 418 177
rect 416 176 417 177
rect 415 176 416 177
rect 414 176 415 177
rect 413 176 414 177
rect 412 176 413 177
rect 411 176 412 177
rect 410 176 411 177
rect 409 176 410 177
rect 408 176 409 177
rect 407 176 408 177
rect 406 176 407 177
rect 266 176 267 177
rect 265 176 266 177
rect 264 176 265 177
rect 263 176 264 177
rect 262 176 263 177
rect 261 176 262 177
rect 260 176 261 177
rect 259 176 260 177
rect 258 176 259 177
rect 257 176 258 177
rect 256 176 257 177
rect 255 176 256 177
rect 254 176 255 177
rect 253 176 254 177
rect 252 176 253 177
rect 251 176 252 177
rect 250 176 251 177
rect 249 176 250 177
rect 248 176 249 177
rect 247 176 248 177
rect 246 176 247 177
rect 245 176 246 177
rect 244 176 245 177
rect 243 176 244 177
rect 242 176 243 177
rect 241 176 242 177
rect 240 176 241 177
rect 239 176 240 177
rect 238 176 239 177
rect 237 176 238 177
rect 236 176 237 177
rect 235 176 236 177
rect 234 176 235 177
rect 233 176 234 177
rect 232 176 233 177
rect 231 176 232 177
rect 230 176 231 177
rect 229 176 230 177
rect 228 176 229 177
rect 227 176 228 177
rect 226 176 227 177
rect 225 176 226 177
rect 224 176 225 177
rect 205 176 206 177
rect 204 176 205 177
rect 203 176 204 177
rect 202 176 203 177
rect 201 176 202 177
rect 200 176 201 177
rect 199 176 200 177
rect 198 176 199 177
rect 197 176 198 177
rect 196 176 197 177
rect 195 176 196 177
rect 194 176 195 177
rect 193 176 194 177
rect 192 176 193 177
rect 191 176 192 177
rect 190 176 191 177
rect 189 176 190 177
rect 188 176 189 177
rect 187 176 188 177
rect 186 176 187 177
rect 185 176 186 177
rect 184 176 185 177
rect 183 176 184 177
rect 182 176 183 177
rect 181 176 182 177
rect 180 176 181 177
rect 179 176 180 177
rect 178 176 179 177
rect 177 176 178 177
rect 176 176 177 177
rect 175 176 176 177
rect 174 176 175 177
rect 173 176 174 177
rect 172 176 173 177
rect 171 176 172 177
rect 170 176 171 177
rect 169 176 170 177
rect 168 176 169 177
rect 167 176 168 177
rect 166 176 167 177
rect 165 176 166 177
rect 164 176 165 177
rect 163 176 164 177
rect 162 176 163 177
rect 161 176 162 177
rect 160 176 161 177
rect 159 176 160 177
rect 158 176 159 177
rect 157 176 158 177
rect 156 176 157 177
rect 155 176 156 177
rect 154 176 155 177
rect 153 176 154 177
rect 152 176 153 177
rect 151 176 152 177
rect 150 176 151 177
rect 149 176 150 177
rect 148 176 149 177
rect 147 176 148 177
rect 146 176 147 177
rect 145 176 146 177
rect 144 176 145 177
rect 143 176 144 177
rect 142 176 143 177
rect 141 176 142 177
rect 140 176 141 177
rect 139 176 140 177
rect 138 176 139 177
rect 137 176 138 177
rect 136 176 137 177
rect 135 176 136 177
rect 134 176 135 177
rect 133 176 134 177
rect 132 176 133 177
rect 131 176 132 177
rect 130 176 131 177
rect 129 176 130 177
rect 128 176 129 177
rect 127 176 128 177
rect 126 176 127 177
rect 125 176 126 177
rect 124 176 125 177
rect 123 176 124 177
rect 55 176 56 177
rect 54 176 55 177
rect 53 176 54 177
rect 52 176 53 177
rect 51 176 52 177
rect 50 176 51 177
rect 49 176 50 177
rect 48 176 49 177
rect 47 176 48 177
rect 46 176 47 177
rect 45 176 46 177
rect 44 176 45 177
rect 43 176 44 177
rect 42 176 43 177
rect 41 176 42 177
rect 40 176 41 177
rect 39 176 40 177
rect 38 176 39 177
rect 37 176 38 177
rect 36 176 37 177
rect 23 176 24 177
rect 22 176 23 177
rect 21 176 22 177
rect 20 176 21 177
rect 19 176 20 177
rect 18 176 19 177
rect 17 176 18 177
rect 16 176 17 177
rect 15 176 16 177
rect 14 176 15 177
rect 13 176 14 177
rect 12 176 13 177
rect 11 176 12 177
rect 467 177 468 178
rect 466 177 467 178
rect 465 177 466 178
rect 464 177 465 178
rect 463 177 464 178
rect 462 177 463 178
rect 461 177 462 178
rect 460 177 461 178
rect 420 177 421 178
rect 419 177 420 178
rect 418 177 419 178
rect 417 177 418 178
rect 416 177 417 178
rect 415 177 416 178
rect 414 177 415 178
rect 413 177 414 178
rect 412 177 413 178
rect 411 177 412 178
rect 410 177 411 178
rect 409 177 410 178
rect 408 177 409 178
rect 407 177 408 178
rect 265 177 266 178
rect 264 177 265 178
rect 263 177 264 178
rect 262 177 263 178
rect 261 177 262 178
rect 260 177 261 178
rect 259 177 260 178
rect 258 177 259 178
rect 257 177 258 178
rect 256 177 257 178
rect 255 177 256 178
rect 254 177 255 178
rect 253 177 254 178
rect 252 177 253 178
rect 251 177 252 178
rect 250 177 251 178
rect 249 177 250 178
rect 248 177 249 178
rect 247 177 248 178
rect 246 177 247 178
rect 245 177 246 178
rect 244 177 245 178
rect 243 177 244 178
rect 242 177 243 178
rect 241 177 242 178
rect 240 177 241 178
rect 239 177 240 178
rect 238 177 239 178
rect 237 177 238 178
rect 236 177 237 178
rect 235 177 236 178
rect 234 177 235 178
rect 233 177 234 178
rect 232 177 233 178
rect 231 177 232 178
rect 230 177 231 178
rect 229 177 230 178
rect 228 177 229 178
rect 227 177 228 178
rect 226 177 227 178
rect 225 177 226 178
rect 224 177 225 178
rect 204 177 205 178
rect 203 177 204 178
rect 202 177 203 178
rect 201 177 202 178
rect 200 177 201 178
rect 199 177 200 178
rect 198 177 199 178
rect 197 177 198 178
rect 196 177 197 178
rect 195 177 196 178
rect 194 177 195 178
rect 193 177 194 178
rect 192 177 193 178
rect 191 177 192 178
rect 190 177 191 178
rect 189 177 190 178
rect 188 177 189 178
rect 187 177 188 178
rect 186 177 187 178
rect 185 177 186 178
rect 184 177 185 178
rect 183 177 184 178
rect 182 177 183 178
rect 181 177 182 178
rect 180 177 181 178
rect 179 177 180 178
rect 178 177 179 178
rect 177 177 178 178
rect 176 177 177 178
rect 175 177 176 178
rect 174 177 175 178
rect 173 177 174 178
rect 172 177 173 178
rect 171 177 172 178
rect 170 177 171 178
rect 169 177 170 178
rect 168 177 169 178
rect 167 177 168 178
rect 166 177 167 178
rect 165 177 166 178
rect 164 177 165 178
rect 163 177 164 178
rect 162 177 163 178
rect 161 177 162 178
rect 160 177 161 178
rect 159 177 160 178
rect 158 177 159 178
rect 157 177 158 178
rect 156 177 157 178
rect 155 177 156 178
rect 154 177 155 178
rect 153 177 154 178
rect 152 177 153 178
rect 151 177 152 178
rect 150 177 151 178
rect 149 177 150 178
rect 148 177 149 178
rect 147 177 148 178
rect 146 177 147 178
rect 145 177 146 178
rect 144 177 145 178
rect 143 177 144 178
rect 142 177 143 178
rect 141 177 142 178
rect 140 177 141 178
rect 139 177 140 178
rect 138 177 139 178
rect 137 177 138 178
rect 136 177 137 178
rect 135 177 136 178
rect 134 177 135 178
rect 133 177 134 178
rect 132 177 133 178
rect 131 177 132 178
rect 130 177 131 178
rect 129 177 130 178
rect 128 177 129 178
rect 127 177 128 178
rect 126 177 127 178
rect 125 177 126 178
rect 124 177 125 178
rect 123 177 124 178
rect 122 177 123 178
rect 121 177 122 178
rect 54 177 55 178
rect 53 177 54 178
rect 52 177 53 178
rect 51 177 52 178
rect 50 177 51 178
rect 49 177 50 178
rect 48 177 49 178
rect 47 177 48 178
rect 46 177 47 178
rect 45 177 46 178
rect 44 177 45 178
rect 43 177 44 178
rect 42 177 43 178
rect 41 177 42 178
rect 40 177 41 178
rect 39 177 40 178
rect 38 177 39 178
rect 37 177 38 178
rect 36 177 37 178
rect 23 177 24 178
rect 22 177 23 178
rect 21 177 22 178
rect 20 177 21 178
rect 19 177 20 178
rect 18 177 19 178
rect 17 177 18 178
rect 16 177 17 178
rect 15 177 16 178
rect 14 177 15 178
rect 13 177 14 178
rect 12 177 13 178
rect 11 177 12 178
rect 465 178 466 179
rect 464 178 465 179
rect 463 178 464 179
rect 462 178 463 179
rect 461 178 462 179
rect 460 178 461 179
rect 422 178 423 179
rect 421 178 422 179
rect 420 178 421 179
rect 419 178 420 179
rect 418 178 419 179
rect 417 178 418 179
rect 416 178 417 179
rect 415 178 416 179
rect 414 178 415 179
rect 413 178 414 179
rect 412 178 413 179
rect 411 178 412 179
rect 410 178 411 179
rect 409 178 410 179
rect 408 178 409 179
rect 265 178 266 179
rect 264 178 265 179
rect 263 178 264 179
rect 262 178 263 179
rect 261 178 262 179
rect 260 178 261 179
rect 259 178 260 179
rect 258 178 259 179
rect 257 178 258 179
rect 256 178 257 179
rect 255 178 256 179
rect 254 178 255 179
rect 253 178 254 179
rect 252 178 253 179
rect 251 178 252 179
rect 250 178 251 179
rect 249 178 250 179
rect 248 178 249 179
rect 247 178 248 179
rect 246 178 247 179
rect 245 178 246 179
rect 244 178 245 179
rect 243 178 244 179
rect 242 178 243 179
rect 241 178 242 179
rect 240 178 241 179
rect 239 178 240 179
rect 238 178 239 179
rect 237 178 238 179
rect 236 178 237 179
rect 235 178 236 179
rect 234 178 235 179
rect 233 178 234 179
rect 232 178 233 179
rect 231 178 232 179
rect 230 178 231 179
rect 229 178 230 179
rect 228 178 229 179
rect 227 178 228 179
rect 226 178 227 179
rect 225 178 226 179
rect 224 178 225 179
rect 223 178 224 179
rect 204 178 205 179
rect 203 178 204 179
rect 202 178 203 179
rect 201 178 202 179
rect 200 178 201 179
rect 199 178 200 179
rect 198 178 199 179
rect 197 178 198 179
rect 196 178 197 179
rect 195 178 196 179
rect 194 178 195 179
rect 193 178 194 179
rect 192 178 193 179
rect 191 178 192 179
rect 190 178 191 179
rect 189 178 190 179
rect 188 178 189 179
rect 187 178 188 179
rect 186 178 187 179
rect 185 178 186 179
rect 184 178 185 179
rect 183 178 184 179
rect 182 178 183 179
rect 181 178 182 179
rect 180 178 181 179
rect 179 178 180 179
rect 178 178 179 179
rect 177 178 178 179
rect 176 178 177 179
rect 175 178 176 179
rect 174 178 175 179
rect 173 178 174 179
rect 172 178 173 179
rect 171 178 172 179
rect 170 178 171 179
rect 169 178 170 179
rect 168 178 169 179
rect 167 178 168 179
rect 166 178 167 179
rect 165 178 166 179
rect 164 178 165 179
rect 163 178 164 179
rect 162 178 163 179
rect 161 178 162 179
rect 160 178 161 179
rect 159 178 160 179
rect 158 178 159 179
rect 157 178 158 179
rect 156 178 157 179
rect 155 178 156 179
rect 154 178 155 179
rect 153 178 154 179
rect 152 178 153 179
rect 151 178 152 179
rect 150 178 151 179
rect 149 178 150 179
rect 148 178 149 179
rect 147 178 148 179
rect 146 178 147 179
rect 145 178 146 179
rect 144 178 145 179
rect 143 178 144 179
rect 142 178 143 179
rect 141 178 142 179
rect 140 178 141 179
rect 139 178 140 179
rect 138 178 139 179
rect 137 178 138 179
rect 136 178 137 179
rect 135 178 136 179
rect 134 178 135 179
rect 133 178 134 179
rect 132 178 133 179
rect 131 178 132 179
rect 130 178 131 179
rect 129 178 130 179
rect 128 178 129 179
rect 127 178 128 179
rect 126 178 127 179
rect 125 178 126 179
rect 124 178 125 179
rect 123 178 124 179
rect 122 178 123 179
rect 121 178 122 179
rect 120 178 121 179
rect 119 178 120 179
rect 118 178 119 179
rect 53 178 54 179
rect 52 178 53 179
rect 51 178 52 179
rect 50 178 51 179
rect 49 178 50 179
rect 48 178 49 179
rect 47 178 48 179
rect 46 178 47 179
rect 45 178 46 179
rect 44 178 45 179
rect 43 178 44 179
rect 42 178 43 179
rect 41 178 42 179
rect 40 178 41 179
rect 39 178 40 179
rect 38 178 39 179
rect 37 178 38 179
rect 23 178 24 179
rect 22 178 23 179
rect 21 178 22 179
rect 20 178 21 179
rect 19 178 20 179
rect 18 178 19 179
rect 17 178 18 179
rect 16 178 17 179
rect 15 178 16 179
rect 14 178 15 179
rect 13 178 14 179
rect 12 178 13 179
rect 11 178 12 179
rect 463 179 464 180
rect 462 179 463 180
rect 461 179 462 180
rect 460 179 461 180
rect 423 179 424 180
rect 422 179 423 180
rect 421 179 422 180
rect 420 179 421 180
rect 419 179 420 180
rect 418 179 419 180
rect 417 179 418 180
rect 416 179 417 180
rect 415 179 416 180
rect 414 179 415 180
rect 413 179 414 180
rect 412 179 413 180
rect 411 179 412 180
rect 410 179 411 180
rect 409 179 410 180
rect 264 179 265 180
rect 263 179 264 180
rect 262 179 263 180
rect 261 179 262 180
rect 260 179 261 180
rect 259 179 260 180
rect 258 179 259 180
rect 257 179 258 180
rect 256 179 257 180
rect 255 179 256 180
rect 254 179 255 180
rect 253 179 254 180
rect 252 179 253 180
rect 251 179 252 180
rect 250 179 251 180
rect 249 179 250 180
rect 248 179 249 180
rect 247 179 248 180
rect 246 179 247 180
rect 245 179 246 180
rect 244 179 245 180
rect 243 179 244 180
rect 242 179 243 180
rect 241 179 242 180
rect 240 179 241 180
rect 239 179 240 180
rect 238 179 239 180
rect 237 179 238 180
rect 236 179 237 180
rect 235 179 236 180
rect 234 179 235 180
rect 233 179 234 180
rect 232 179 233 180
rect 231 179 232 180
rect 230 179 231 180
rect 229 179 230 180
rect 228 179 229 180
rect 227 179 228 180
rect 226 179 227 180
rect 225 179 226 180
rect 224 179 225 180
rect 223 179 224 180
rect 203 179 204 180
rect 202 179 203 180
rect 201 179 202 180
rect 200 179 201 180
rect 199 179 200 180
rect 198 179 199 180
rect 197 179 198 180
rect 196 179 197 180
rect 195 179 196 180
rect 194 179 195 180
rect 193 179 194 180
rect 192 179 193 180
rect 191 179 192 180
rect 190 179 191 180
rect 189 179 190 180
rect 188 179 189 180
rect 187 179 188 180
rect 186 179 187 180
rect 185 179 186 180
rect 184 179 185 180
rect 183 179 184 180
rect 182 179 183 180
rect 181 179 182 180
rect 180 179 181 180
rect 179 179 180 180
rect 178 179 179 180
rect 177 179 178 180
rect 176 179 177 180
rect 175 179 176 180
rect 174 179 175 180
rect 173 179 174 180
rect 172 179 173 180
rect 171 179 172 180
rect 170 179 171 180
rect 169 179 170 180
rect 168 179 169 180
rect 167 179 168 180
rect 166 179 167 180
rect 165 179 166 180
rect 164 179 165 180
rect 163 179 164 180
rect 162 179 163 180
rect 161 179 162 180
rect 160 179 161 180
rect 159 179 160 180
rect 158 179 159 180
rect 157 179 158 180
rect 156 179 157 180
rect 155 179 156 180
rect 154 179 155 180
rect 153 179 154 180
rect 152 179 153 180
rect 151 179 152 180
rect 150 179 151 180
rect 149 179 150 180
rect 148 179 149 180
rect 147 179 148 180
rect 146 179 147 180
rect 145 179 146 180
rect 144 179 145 180
rect 143 179 144 180
rect 142 179 143 180
rect 141 179 142 180
rect 140 179 141 180
rect 139 179 140 180
rect 138 179 139 180
rect 137 179 138 180
rect 136 179 137 180
rect 135 179 136 180
rect 134 179 135 180
rect 133 179 134 180
rect 132 179 133 180
rect 131 179 132 180
rect 130 179 131 180
rect 129 179 130 180
rect 128 179 129 180
rect 127 179 128 180
rect 126 179 127 180
rect 125 179 126 180
rect 124 179 125 180
rect 123 179 124 180
rect 122 179 123 180
rect 121 179 122 180
rect 120 179 121 180
rect 119 179 120 180
rect 118 179 119 180
rect 117 179 118 180
rect 116 179 117 180
rect 52 179 53 180
rect 51 179 52 180
rect 50 179 51 180
rect 49 179 50 180
rect 48 179 49 180
rect 47 179 48 180
rect 46 179 47 180
rect 45 179 46 180
rect 44 179 45 180
rect 43 179 44 180
rect 42 179 43 180
rect 41 179 42 180
rect 40 179 41 180
rect 39 179 40 180
rect 38 179 39 180
rect 23 179 24 180
rect 22 179 23 180
rect 21 179 22 180
rect 20 179 21 180
rect 19 179 20 180
rect 18 179 19 180
rect 17 179 18 180
rect 16 179 17 180
rect 15 179 16 180
rect 14 179 15 180
rect 13 179 14 180
rect 12 179 13 180
rect 461 180 462 181
rect 460 180 461 181
rect 424 180 425 181
rect 423 180 424 181
rect 422 180 423 181
rect 421 180 422 181
rect 420 180 421 181
rect 419 180 420 181
rect 418 180 419 181
rect 417 180 418 181
rect 416 180 417 181
rect 415 180 416 181
rect 414 180 415 181
rect 413 180 414 181
rect 412 180 413 181
rect 411 180 412 181
rect 410 180 411 181
rect 317 180 318 181
rect 316 180 317 181
rect 315 180 316 181
rect 314 180 315 181
rect 313 180 314 181
rect 312 180 313 181
rect 311 180 312 181
rect 310 180 311 181
rect 309 180 310 181
rect 308 180 309 181
rect 307 180 308 181
rect 306 180 307 181
rect 305 180 306 181
rect 304 180 305 181
rect 303 180 304 181
rect 302 180 303 181
rect 301 180 302 181
rect 263 180 264 181
rect 262 180 263 181
rect 261 180 262 181
rect 260 180 261 181
rect 259 180 260 181
rect 258 180 259 181
rect 257 180 258 181
rect 256 180 257 181
rect 255 180 256 181
rect 254 180 255 181
rect 253 180 254 181
rect 252 180 253 181
rect 251 180 252 181
rect 250 180 251 181
rect 249 180 250 181
rect 248 180 249 181
rect 247 180 248 181
rect 246 180 247 181
rect 245 180 246 181
rect 244 180 245 181
rect 243 180 244 181
rect 242 180 243 181
rect 241 180 242 181
rect 240 180 241 181
rect 239 180 240 181
rect 238 180 239 181
rect 237 180 238 181
rect 236 180 237 181
rect 235 180 236 181
rect 234 180 235 181
rect 233 180 234 181
rect 232 180 233 181
rect 231 180 232 181
rect 230 180 231 181
rect 229 180 230 181
rect 228 180 229 181
rect 227 180 228 181
rect 226 180 227 181
rect 225 180 226 181
rect 224 180 225 181
rect 223 180 224 181
rect 222 180 223 181
rect 202 180 203 181
rect 201 180 202 181
rect 200 180 201 181
rect 199 180 200 181
rect 198 180 199 181
rect 197 180 198 181
rect 196 180 197 181
rect 195 180 196 181
rect 194 180 195 181
rect 193 180 194 181
rect 192 180 193 181
rect 191 180 192 181
rect 190 180 191 181
rect 189 180 190 181
rect 188 180 189 181
rect 187 180 188 181
rect 186 180 187 181
rect 185 180 186 181
rect 184 180 185 181
rect 183 180 184 181
rect 182 180 183 181
rect 181 180 182 181
rect 180 180 181 181
rect 179 180 180 181
rect 178 180 179 181
rect 177 180 178 181
rect 176 180 177 181
rect 175 180 176 181
rect 174 180 175 181
rect 173 180 174 181
rect 172 180 173 181
rect 171 180 172 181
rect 170 180 171 181
rect 169 180 170 181
rect 168 180 169 181
rect 167 180 168 181
rect 166 180 167 181
rect 165 180 166 181
rect 164 180 165 181
rect 163 180 164 181
rect 162 180 163 181
rect 161 180 162 181
rect 160 180 161 181
rect 159 180 160 181
rect 158 180 159 181
rect 157 180 158 181
rect 156 180 157 181
rect 155 180 156 181
rect 154 180 155 181
rect 153 180 154 181
rect 152 180 153 181
rect 151 180 152 181
rect 150 180 151 181
rect 149 180 150 181
rect 148 180 149 181
rect 147 180 148 181
rect 146 180 147 181
rect 145 180 146 181
rect 144 180 145 181
rect 143 180 144 181
rect 142 180 143 181
rect 141 180 142 181
rect 140 180 141 181
rect 139 180 140 181
rect 138 180 139 181
rect 137 180 138 181
rect 136 180 137 181
rect 135 180 136 181
rect 134 180 135 181
rect 133 180 134 181
rect 132 180 133 181
rect 131 180 132 181
rect 130 180 131 181
rect 129 180 130 181
rect 128 180 129 181
rect 127 180 128 181
rect 126 180 127 181
rect 125 180 126 181
rect 124 180 125 181
rect 123 180 124 181
rect 122 180 123 181
rect 121 180 122 181
rect 120 180 121 181
rect 119 180 120 181
rect 118 180 119 181
rect 117 180 118 181
rect 116 180 117 181
rect 115 180 116 181
rect 114 180 115 181
rect 113 180 114 181
rect 70 180 71 181
rect 69 180 70 181
rect 50 180 51 181
rect 49 180 50 181
rect 48 180 49 181
rect 47 180 48 181
rect 46 180 47 181
rect 45 180 46 181
rect 44 180 45 181
rect 43 180 44 181
rect 42 180 43 181
rect 41 180 42 181
rect 40 180 41 181
rect 39 180 40 181
rect 23 180 24 181
rect 22 180 23 181
rect 21 180 22 181
rect 20 180 21 181
rect 19 180 20 181
rect 18 180 19 181
rect 17 180 18 181
rect 16 180 17 181
rect 15 180 16 181
rect 14 180 15 181
rect 13 180 14 181
rect 12 180 13 181
rect 460 181 461 182
rect 425 181 426 182
rect 424 181 425 182
rect 423 181 424 182
rect 422 181 423 182
rect 421 181 422 182
rect 420 181 421 182
rect 419 181 420 182
rect 418 181 419 182
rect 417 181 418 182
rect 416 181 417 182
rect 415 181 416 182
rect 414 181 415 182
rect 413 181 414 182
rect 412 181 413 182
rect 411 181 412 182
rect 322 181 323 182
rect 321 181 322 182
rect 320 181 321 182
rect 319 181 320 182
rect 318 181 319 182
rect 317 181 318 182
rect 316 181 317 182
rect 315 181 316 182
rect 314 181 315 182
rect 313 181 314 182
rect 312 181 313 182
rect 311 181 312 182
rect 310 181 311 182
rect 309 181 310 182
rect 308 181 309 182
rect 307 181 308 182
rect 306 181 307 182
rect 305 181 306 182
rect 304 181 305 182
rect 303 181 304 182
rect 302 181 303 182
rect 301 181 302 182
rect 300 181 301 182
rect 299 181 300 182
rect 298 181 299 182
rect 297 181 298 182
rect 296 181 297 182
rect 262 181 263 182
rect 261 181 262 182
rect 260 181 261 182
rect 259 181 260 182
rect 258 181 259 182
rect 257 181 258 182
rect 256 181 257 182
rect 255 181 256 182
rect 254 181 255 182
rect 253 181 254 182
rect 252 181 253 182
rect 251 181 252 182
rect 250 181 251 182
rect 249 181 250 182
rect 248 181 249 182
rect 247 181 248 182
rect 246 181 247 182
rect 245 181 246 182
rect 244 181 245 182
rect 243 181 244 182
rect 242 181 243 182
rect 241 181 242 182
rect 240 181 241 182
rect 239 181 240 182
rect 238 181 239 182
rect 237 181 238 182
rect 236 181 237 182
rect 235 181 236 182
rect 234 181 235 182
rect 233 181 234 182
rect 232 181 233 182
rect 231 181 232 182
rect 230 181 231 182
rect 229 181 230 182
rect 228 181 229 182
rect 227 181 228 182
rect 226 181 227 182
rect 225 181 226 182
rect 224 181 225 182
rect 223 181 224 182
rect 222 181 223 182
rect 201 181 202 182
rect 200 181 201 182
rect 199 181 200 182
rect 198 181 199 182
rect 197 181 198 182
rect 196 181 197 182
rect 195 181 196 182
rect 194 181 195 182
rect 193 181 194 182
rect 192 181 193 182
rect 191 181 192 182
rect 190 181 191 182
rect 189 181 190 182
rect 188 181 189 182
rect 187 181 188 182
rect 186 181 187 182
rect 185 181 186 182
rect 184 181 185 182
rect 183 181 184 182
rect 182 181 183 182
rect 181 181 182 182
rect 180 181 181 182
rect 179 181 180 182
rect 178 181 179 182
rect 177 181 178 182
rect 176 181 177 182
rect 175 181 176 182
rect 174 181 175 182
rect 173 181 174 182
rect 172 181 173 182
rect 171 181 172 182
rect 170 181 171 182
rect 169 181 170 182
rect 168 181 169 182
rect 167 181 168 182
rect 166 181 167 182
rect 165 181 166 182
rect 164 181 165 182
rect 163 181 164 182
rect 162 181 163 182
rect 161 181 162 182
rect 160 181 161 182
rect 159 181 160 182
rect 158 181 159 182
rect 157 181 158 182
rect 156 181 157 182
rect 155 181 156 182
rect 154 181 155 182
rect 153 181 154 182
rect 152 181 153 182
rect 151 181 152 182
rect 150 181 151 182
rect 149 181 150 182
rect 148 181 149 182
rect 147 181 148 182
rect 146 181 147 182
rect 145 181 146 182
rect 144 181 145 182
rect 143 181 144 182
rect 142 181 143 182
rect 141 181 142 182
rect 140 181 141 182
rect 139 181 140 182
rect 138 181 139 182
rect 137 181 138 182
rect 136 181 137 182
rect 135 181 136 182
rect 134 181 135 182
rect 133 181 134 182
rect 132 181 133 182
rect 131 181 132 182
rect 130 181 131 182
rect 129 181 130 182
rect 128 181 129 182
rect 127 181 128 182
rect 126 181 127 182
rect 125 181 126 182
rect 124 181 125 182
rect 123 181 124 182
rect 122 181 123 182
rect 121 181 122 182
rect 120 181 121 182
rect 119 181 120 182
rect 118 181 119 182
rect 117 181 118 182
rect 116 181 117 182
rect 115 181 116 182
rect 114 181 115 182
rect 113 181 114 182
rect 112 181 113 182
rect 111 181 112 182
rect 72 181 73 182
rect 71 181 72 182
rect 70 181 71 182
rect 69 181 70 182
rect 48 181 49 182
rect 47 181 48 182
rect 46 181 47 182
rect 45 181 46 182
rect 44 181 45 182
rect 43 181 44 182
rect 42 181 43 182
rect 41 181 42 182
rect 23 181 24 182
rect 22 181 23 182
rect 21 181 22 182
rect 20 181 21 182
rect 19 181 20 182
rect 18 181 19 182
rect 17 181 18 182
rect 16 181 17 182
rect 15 181 16 182
rect 14 181 15 182
rect 13 181 14 182
rect 12 181 13 182
rect 460 182 461 183
rect 426 182 427 183
rect 425 182 426 183
rect 424 182 425 183
rect 423 182 424 183
rect 422 182 423 183
rect 421 182 422 183
rect 420 182 421 183
rect 419 182 420 183
rect 418 182 419 183
rect 417 182 418 183
rect 416 182 417 183
rect 415 182 416 183
rect 414 182 415 183
rect 413 182 414 183
rect 325 182 326 183
rect 324 182 325 183
rect 323 182 324 183
rect 322 182 323 183
rect 321 182 322 183
rect 320 182 321 183
rect 319 182 320 183
rect 318 182 319 183
rect 317 182 318 183
rect 316 182 317 183
rect 315 182 316 183
rect 314 182 315 183
rect 313 182 314 183
rect 312 182 313 183
rect 311 182 312 183
rect 310 182 311 183
rect 309 182 310 183
rect 308 182 309 183
rect 307 182 308 183
rect 306 182 307 183
rect 305 182 306 183
rect 304 182 305 183
rect 303 182 304 183
rect 302 182 303 183
rect 301 182 302 183
rect 300 182 301 183
rect 299 182 300 183
rect 298 182 299 183
rect 297 182 298 183
rect 296 182 297 183
rect 295 182 296 183
rect 294 182 295 183
rect 293 182 294 183
rect 292 182 293 183
rect 261 182 262 183
rect 260 182 261 183
rect 259 182 260 183
rect 258 182 259 183
rect 257 182 258 183
rect 256 182 257 183
rect 255 182 256 183
rect 254 182 255 183
rect 253 182 254 183
rect 252 182 253 183
rect 251 182 252 183
rect 250 182 251 183
rect 249 182 250 183
rect 248 182 249 183
rect 247 182 248 183
rect 246 182 247 183
rect 245 182 246 183
rect 244 182 245 183
rect 243 182 244 183
rect 242 182 243 183
rect 241 182 242 183
rect 240 182 241 183
rect 239 182 240 183
rect 238 182 239 183
rect 237 182 238 183
rect 236 182 237 183
rect 235 182 236 183
rect 234 182 235 183
rect 233 182 234 183
rect 232 182 233 183
rect 231 182 232 183
rect 230 182 231 183
rect 229 182 230 183
rect 228 182 229 183
rect 227 182 228 183
rect 226 182 227 183
rect 225 182 226 183
rect 224 182 225 183
rect 223 182 224 183
rect 222 182 223 183
rect 221 182 222 183
rect 201 182 202 183
rect 200 182 201 183
rect 199 182 200 183
rect 198 182 199 183
rect 197 182 198 183
rect 196 182 197 183
rect 195 182 196 183
rect 194 182 195 183
rect 193 182 194 183
rect 192 182 193 183
rect 191 182 192 183
rect 190 182 191 183
rect 189 182 190 183
rect 188 182 189 183
rect 187 182 188 183
rect 186 182 187 183
rect 185 182 186 183
rect 184 182 185 183
rect 183 182 184 183
rect 182 182 183 183
rect 181 182 182 183
rect 180 182 181 183
rect 179 182 180 183
rect 178 182 179 183
rect 177 182 178 183
rect 176 182 177 183
rect 175 182 176 183
rect 174 182 175 183
rect 173 182 174 183
rect 172 182 173 183
rect 171 182 172 183
rect 170 182 171 183
rect 169 182 170 183
rect 168 182 169 183
rect 167 182 168 183
rect 166 182 167 183
rect 165 182 166 183
rect 164 182 165 183
rect 163 182 164 183
rect 162 182 163 183
rect 161 182 162 183
rect 160 182 161 183
rect 159 182 160 183
rect 158 182 159 183
rect 157 182 158 183
rect 156 182 157 183
rect 155 182 156 183
rect 154 182 155 183
rect 153 182 154 183
rect 152 182 153 183
rect 151 182 152 183
rect 150 182 151 183
rect 149 182 150 183
rect 148 182 149 183
rect 147 182 148 183
rect 146 182 147 183
rect 145 182 146 183
rect 144 182 145 183
rect 143 182 144 183
rect 142 182 143 183
rect 141 182 142 183
rect 140 182 141 183
rect 139 182 140 183
rect 138 182 139 183
rect 137 182 138 183
rect 136 182 137 183
rect 135 182 136 183
rect 134 182 135 183
rect 133 182 134 183
rect 132 182 133 183
rect 131 182 132 183
rect 130 182 131 183
rect 129 182 130 183
rect 128 182 129 183
rect 127 182 128 183
rect 126 182 127 183
rect 125 182 126 183
rect 124 182 125 183
rect 123 182 124 183
rect 122 182 123 183
rect 121 182 122 183
rect 120 182 121 183
rect 119 182 120 183
rect 118 182 119 183
rect 117 182 118 183
rect 116 182 117 183
rect 115 182 116 183
rect 114 182 115 183
rect 113 182 114 183
rect 112 182 113 183
rect 111 182 112 183
rect 110 182 111 183
rect 109 182 110 183
rect 108 182 109 183
rect 107 182 108 183
rect 75 182 76 183
rect 74 182 75 183
rect 73 182 74 183
rect 72 182 73 183
rect 71 182 72 183
rect 70 182 71 183
rect 69 182 70 183
rect 24 182 25 183
rect 23 182 24 183
rect 22 182 23 183
rect 21 182 22 183
rect 20 182 21 183
rect 19 182 20 183
rect 18 182 19 183
rect 17 182 18 183
rect 16 182 17 183
rect 15 182 16 183
rect 14 182 15 183
rect 13 182 14 183
rect 12 182 13 183
rect 428 183 429 184
rect 427 183 428 184
rect 426 183 427 184
rect 425 183 426 184
rect 424 183 425 184
rect 423 183 424 184
rect 422 183 423 184
rect 421 183 422 184
rect 420 183 421 184
rect 419 183 420 184
rect 418 183 419 184
rect 417 183 418 184
rect 416 183 417 184
rect 415 183 416 184
rect 414 183 415 184
rect 327 183 328 184
rect 326 183 327 184
rect 325 183 326 184
rect 324 183 325 184
rect 323 183 324 184
rect 322 183 323 184
rect 321 183 322 184
rect 320 183 321 184
rect 319 183 320 184
rect 318 183 319 184
rect 317 183 318 184
rect 316 183 317 184
rect 315 183 316 184
rect 314 183 315 184
rect 313 183 314 184
rect 312 183 313 184
rect 311 183 312 184
rect 310 183 311 184
rect 309 183 310 184
rect 308 183 309 184
rect 307 183 308 184
rect 306 183 307 184
rect 305 183 306 184
rect 304 183 305 184
rect 303 183 304 184
rect 302 183 303 184
rect 301 183 302 184
rect 300 183 301 184
rect 299 183 300 184
rect 298 183 299 184
rect 297 183 298 184
rect 296 183 297 184
rect 295 183 296 184
rect 294 183 295 184
rect 293 183 294 184
rect 292 183 293 184
rect 291 183 292 184
rect 290 183 291 184
rect 289 183 290 184
rect 261 183 262 184
rect 260 183 261 184
rect 259 183 260 184
rect 258 183 259 184
rect 257 183 258 184
rect 256 183 257 184
rect 255 183 256 184
rect 254 183 255 184
rect 253 183 254 184
rect 252 183 253 184
rect 251 183 252 184
rect 250 183 251 184
rect 249 183 250 184
rect 248 183 249 184
rect 247 183 248 184
rect 246 183 247 184
rect 245 183 246 184
rect 244 183 245 184
rect 243 183 244 184
rect 242 183 243 184
rect 241 183 242 184
rect 240 183 241 184
rect 239 183 240 184
rect 238 183 239 184
rect 237 183 238 184
rect 236 183 237 184
rect 235 183 236 184
rect 234 183 235 184
rect 233 183 234 184
rect 232 183 233 184
rect 231 183 232 184
rect 230 183 231 184
rect 229 183 230 184
rect 228 183 229 184
rect 227 183 228 184
rect 226 183 227 184
rect 225 183 226 184
rect 224 183 225 184
rect 223 183 224 184
rect 222 183 223 184
rect 221 183 222 184
rect 200 183 201 184
rect 199 183 200 184
rect 198 183 199 184
rect 197 183 198 184
rect 196 183 197 184
rect 195 183 196 184
rect 194 183 195 184
rect 193 183 194 184
rect 192 183 193 184
rect 191 183 192 184
rect 190 183 191 184
rect 189 183 190 184
rect 188 183 189 184
rect 187 183 188 184
rect 186 183 187 184
rect 185 183 186 184
rect 184 183 185 184
rect 183 183 184 184
rect 182 183 183 184
rect 181 183 182 184
rect 180 183 181 184
rect 179 183 180 184
rect 178 183 179 184
rect 177 183 178 184
rect 176 183 177 184
rect 175 183 176 184
rect 174 183 175 184
rect 173 183 174 184
rect 172 183 173 184
rect 171 183 172 184
rect 170 183 171 184
rect 169 183 170 184
rect 168 183 169 184
rect 167 183 168 184
rect 166 183 167 184
rect 165 183 166 184
rect 164 183 165 184
rect 163 183 164 184
rect 162 183 163 184
rect 161 183 162 184
rect 160 183 161 184
rect 159 183 160 184
rect 158 183 159 184
rect 157 183 158 184
rect 156 183 157 184
rect 155 183 156 184
rect 154 183 155 184
rect 153 183 154 184
rect 152 183 153 184
rect 151 183 152 184
rect 150 183 151 184
rect 149 183 150 184
rect 148 183 149 184
rect 147 183 148 184
rect 146 183 147 184
rect 145 183 146 184
rect 144 183 145 184
rect 143 183 144 184
rect 142 183 143 184
rect 141 183 142 184
rect 140 183 141 184
rect 139 183 140 184
rect 138 183 139 184
rect 137 183 138 184
rect 136 183 137 184
rect 135 183 136 184
rect 134 183 135 184
rect 133 183 134 184
rect 132 183 133 184
rect 131 183 132 184
rect 130 183 131 184
rect 129 183 130 184
rect 128 183 129 184
rect 127 183 128 184
rect 126 183 127 184
rect 125 183 126 184
rect 124 183 125 184
rect 123 183 124 184
rect 122 183 123 184
rect 121 183 122 184
rect 120 183 121 184
rect 119 183 120 184
rect 118 183 119 184
rect 117 183 118 184
rect 116 183 117 184
rect 115 183 116 184
rect 114 183 115 184
rect 113 183 114 184
rect 112 183 113 184
rect 111 183 112 184
rect 110 183 111 184
rect 109 183 110 184
rect 108 183 109 184
rect 107 183 108 184
rect 106 183 107 184
rect 105 183 106 184
rect 104 183 105 184
rect 77 183 78 184
rect 76 183 77 184
rect 75 183 76 184
rect 74 183 75 184
rect 73 183 74 184
rect 72 183 73 184
rect 71 183 72 184
rect 70 183 71 184
rect 24 183 25 184
rect 23 183 24 184
rect 22 183 23 184
rect 21 183 22 184
rect 20 183 21 184
rect 19 183 20 184
rect 18 183 19 184
rect 17 183 18 184
rect 16 183 17 184
rect 15 183 16 184
rect 14 183 15 184
rect 13 183 14 184
rect 12 183 13 184
rect 429 184 430 185
rect 428 184 429 185
rect 427 184 428 185
rect 426 184 427 185
rect 425 184 426 185
rect 424 184 425 185
rect 423 184 424 185
rect 422 184 423 185
rect 421 184 422 185
rect 420 184 421 185
rect 419 184 420 185
rect 418 184 419 185
rect 417 184 418 185
rect 416 184 417 185
rect 415 184 416 185
rect 329 184 330 185
rect 328 184 329 185
rect 327 184 328 185
rect 326 184 327 185
rect 325 184 326 185
rect 324 184 325 185
rect 323 184 324 185
rect 322 184 323 185
rect 321 184 322 185
rect 320 184 321 185
rect 319 184 320 185
rect 318 184 319 185
rect 317 184 318 185
rect 316 184 317 185
rect 315 184 316 185
rect 314 184 315 185
rect 313 184 314 185
rect 312 184 313 185
rect 311 184 312 185
rect 310 184 311 185
rect 309 184 310 185
rect 308 184 309 185
rect 307 184 308 185
rect 306 184 307 185
rect 305 184 306 185
rect 304 184 305 185
rect 303 184 304 185
rect 302 184 303 185
rect 301 184 302 185
rect 300 184 301 185
rect 299 184 300 185
rect 298 184 299 185
rect 297 184 298 185
rect 296 184 297 185
rect 295 184 296 185
rect 294 184 295 185
rect 293 184 294 185
rect 292 184 293 185
rect 291 184 292 185
rect 290 184 291 185
rect 289 184 290 185
rect 288 184 289 185
rect 287 184 288 185
rect 260 184 261 185
rect 259 184 260 185
rect 258 184 259 185
rect 257 184 258 185
rect 256 184 257 185
rect 255 184 256 185
rect 254 184 255 185
rect 253 184 254 185
rect 252 184 253 185
rect 251 184 252 185
rect 250 184 251 185
rect 249 184 250 185
rect 248 184 249 185
rect 247 184 248 185
rect 246 184 247 185
rect 245 184 246 185
rect 244 184 245 185
rect 243 184 244 185
rect 242 184 243 185
rect 241 184 242 185
rect 240 184 241 185
rect 239 184 240 185
rect 238 184 239 185
rect 237 184 238 185
rect 236 184 237 185
rect 235 184 236 185
rect 234 184 235 185
rect 233 184 234 185
rect 232 184 233 185
rect 231 184 232 185
rect 230 184 231 185
rect 229 184 230 185
rect 228 184 229 185
rect 227 184 228 185
rect 226 184 227 185
rect 225 184 226 185
rect 224 184 225 185
rect 223 184 224 185
rect 222 184 223 185
rect 221 184 222 185
rect 220 184 221 185
rect 199 184 200 185
rect 198 184 199 185
rect 197 184 198 185
rect 196 184 197 185
rect 195 184 196 185
rect 194 184 195 185
rect 193 184 194 185
rect 192 184 193 185
rect 191 184 192 185
rect 190 184 191 185
rect 189 184 190 185
rect 188 184 189 185
rect 187 184 188 185
rect 186 184 187 185
rect 185 184 186 185
rect 184 184 185 185
rect 183 184 184 185
rect 182 184 183 185
rect 181 184 182 185
rect 180 184 181 185
rect 179 184 180 185
rect 178 184 179 185
rect 177 184 178 185
rect 176 184 177 185
rect 175 184 176 185
rect 174 184 175 185
rect 173 184 174 185
rect 172 184 173 185
rect 171 184 172 185
rect 170 184 171 185
rect 169 184 170 185
rect 168 184 169 185
rect 167 184 168 185
rect 166 184 167 185
rect 165 184 166 185
rect 164 184 165 185
rect 163 184 164 185
rect 162 184 163 185
rect 161 184 162 185
rect 160 184 161 185
rect 159 184 160 185
rect 158 184 159 185
rect 157 184 158 185
rect 156 184 157 185
rect 155 184 156 185
rect 154 184 155 185
rect 153 184 154 185
rect 152 184 153 185
rect 151 184 152 185
rect 150 184 151 185
rect 149 184 150 185
rect 148 184 149 185
rect 147 184 148 185
rect 146 184 147 185
rect 145 184 146 185
rect 144 184 145 185
rect 143 184 144 185
rect 142 184 143 185
rect 141 184 142 185
rect 140 184 141 185
rect 139 184 140 185
rect 138 184 139 185
rect 137 184 138 185
rect 136 184 137 185
rect 135 184 136 185
rect 134 184 135 185
rect 133 184 134 185
rect 132 184 133 185
rect 131 184 132 185
rect 130 184 131 185
rect 129 184 130 185
rect 128 184 129 185
rect 127 184 128 185
rect 126 184 127 185
rect 125 184 126 185
rect 124 184 125 185
rect 123 184 124 185
rect 122 184 123 185
rect 121 184 122 185
rect 120 184 121 185
rect 119 184 120 185
rect 118 184 119 185
rect 117 184 118 185
rect 116 184 117 185
rect 115 184 116 185
rect 114 184 115 185
rect 113 184 114 185
rect 112 184 113 185
rect 111 184 112 185
rect 110 184 111 185
rect 109 184 110 185
rect 108 184 109 185
rect 107 184 108 185
rect 106 184 107 185
rect 105 184 106 185
rect 104 184 105 185
rect 103 184 104 185
rect 102 184 103 185
rect 101 184 102 185
rect 100 184 101 185
rect 99 184 100 185
rect 81 184 82 185
rect 80 184 81 185
rect 79 184 80 185
rect 78 184 79 185
rect 77 184 78 185
rect 76 184 77 185
rect 75 184 76 185
rect 74 184 75 185
rect 73 184 74 185
rect 72 184 73 185
rect 71 184 72 185
rect 70 184 71 185
rect 24 184 25 185
rect 23 184 24 185
rect 22 184 23 185
rect 21 184 22 185
rect 20 184 21 185
rect 19 184 20 185
rect 18 184 19 185
rect 17 184 18 185
rect 16 184 17 185
rect 15 184 16 185
rect 14 184 15 185
rect 13 184 14 185
rect 12 184 13 185
rect 430 185 431 186
rect 429 185 430 186
rect 428 185 429 186
rect 427 185 428 186
rect 426 185 427 186
rect 425 185 426 186
rect 424 185 425 186
rect 423 185 424 186
rect 422 185 423 186
rect 421 185 422 186
rect 420 185 421 186
rect 419 185 420 186
rect 418 185 419 186
rect 417 185 418 186
rect 416 185 417 186
rect 331 185 332 186
rect 330 185 331 186
rect 329 185 330 186
rect 328 185 329 186
rect 327 185 328 186
rect 326 185 327 186
rect 325 185 326 186
rect 324 185 325 186
rect 323 185 324 186
rect 322 185 323 186
rect 321 185 322 186
rect 320 185 321 186
rect 319 185 320 186
rect 318 185 319 186
rect 317 185 318 186
rect 316 185 317 186
rect 315 185 316 186
rect 314 185 315 186
rect 313 185 314 186
rect 312 185 313 186
rect 311 185 312 186
rect 310 185 311 186
rect 309 185 310 186
rect 308 185 309 186
rect 307 185 308 186
rect 306 185 307 186
rect 305 185 306 186
rect 304 185 305 186
rect 303 185 304 186
rect 302 185 303 186
rect 301 185 302 186
rect 300 185 301 186
rect 299 185 300 186
rect 298 185 299 186
rect 297 185 298 186
rect 296 185 297 186
rect 295 185 296 186
rect 294 185 295 186
rect 293 185 294 186
rect 292 185 293 186
rect 291 185 292 186
rect 290 185 291 186
rect 289 185 290 186
rect 288 185 289 186
rect 287 185 288 186
rect 286 185 287 186
rect 285 185 286 186
rect 284 185 285 186
rect 259 185 260 186
rect 258 185 259 186
rect 257 185 258 186
rect 256 185 257 186
rect 255 185 256 186
rect 254 185 255 186
rect 253 185 254 186
rect 252 185 253 186
rect 251 185 252 186
rect 250 185 251 186
rect 249 185 250 186
rect 248 185 249 186
rect 247 185 248 186
rect 246 185 247 186
rect 245 185 246 186
rect 244 185 245 186
rect 243 185 244 186
rect 242 185 243 186
rect 241 185 242 186
rect 240 185 241 186
rect 239 185 240 186
rect 238 185 239 186
rect 237 185 238 186
rect 236 185 237 186
rect 235 185 236 186
rect 234 185 235 186
rect 233 185 234 186
rect 232 185 233 186
rect 231 185 232 186
rect 230 185 231 186
rect 229 185 230 186
rect 228 185 229 186
rect 227 185 228 186
rect 226 185 227 186
rect 225 185 226 186
rect 224 185 225 186
rect 223 185 224 186
rect 222 185 223 186
rect 221 185 222 186
rect 220 185 221 186
rect 219 185 220 186
rect 198 185 199 186
rect 197 185 198 186
rect 196 185 197 186
rect 195 185 196 186
rect 194 185 195 186
rect 193 185 194 186
rect 192 185 193 186
rect 191 185 192 186
rect 190 185 191 186
rect 189 185 190 186
rect 188 185 189 186
rect 187 185 188 186
rect 186 185 187 186
rect 185 185 186 186
rect 184 185 185 186
rect 183 185 184 186
rect 182 185 183 186
rect 181 185 182 186
rect 180 185 181 186
rect 179 185 180 186
rect 178 185 179 186
rect 177 185 178 186
rect 176 185 177 186
rect 175 185 176 186
rect 174 185 175 186
rect 173 185 174 186
rect 172 185 173 186
rect 171 185 172 186
rect 170 185 171 186
rect 169 185 170 186
rect 168 185 169 186
rect 167 185 168 186
rect 166 185 167 186
rect 165 185 166 186
rect 164 185 165 186
rect 163 185 164 186
rect 162 185 163 186
rect 161 185 162 186
rect 160 185 161 186
rect 159 185 160 186
rect 158 185 159 186
rect 157 185 158 186
rect 156 185 157 186
rect 155 185 156 186
rect 154 185 155 186
rect 153 185 154 186
rect 152 185 153 186
rect 151 185 152 186
rect 150 185 151 186
rect 149 185 150 186
rect 148 185 149 186
rect 147 185 148 186
rect 146 185 147 186
rect 145 185 146 186
rect 144 185 145 186
rect 143 185 144 186
rect 142 185 143 186
rect 141 185 142 186
rect 140 185 141 186
rect 139 185 140 186
rect 138 185 139 186
rect 137 185 138 186
rect 136 185 137 186
rect 135 185 136 186
rect 134 185 135 186
rect 133 185 134 186
rect 132 185 133 186
rect 131 185 132 186
rect 130 185 131 186
rect 129 185 130 186
rect 128 185 129 186
rect 127 185 128 186
rect 126 185 127 186
rect 125 185 126 186
rect 124 185 125 186
rect 123 185 124 186
rect 122 185 123 186
rect 121 185 122 186
rect 120 185 121 186
rect 119 185 120 186
rect 118 185 119 186
rect 117 185 118 186
rect 116 185 117 186
rect 115 185 116 186
rect 114 185 115 186
rect 113 185 114 186
rect 112 185 113 186
rect 111 185 112 186
rect 110 185 111 186
rect 109 185 110 186
rect 108 185 109 186
rect 107 185 108 186
rect 106 185 107 186
rect 105 185 106 186
rect 104 185 105 186
rect 103 185 104 186
rect 102 185 103 186
rect 101 185 102 186
rect 100 185 101 186
rect 99 185 100 186
rect 98 185 99 186
rect 97 185 98 186
rect 96 185 97 186
rect 95 185 96 186
rect 94 185 95 186
rect 93 185 94 186
rect 92 185 93 186
rect 91 185 92 186
rect 90 185 91 186
rect 89 185 90 186
rect 88 185 89 186
rect 87 185 88 186
rect 86 185 87 186
rect 85 185 86 186
rect 84 185 85 186
rect 83 185 84 186
rect 82 185 83 186
rect 81 185 82 186
rect 80 185 81 186
rect 79 185 80 186
rect 78 185 79 186
rect 77 185 78 186
rect 76 185 77 186
rect 75 185 76 186
rect 74 185 75 186
rect 73 185 74 186
rect 72 185 73 186
rect 71 185 72 186
rect 70 185 71 186
rect 24 185 25 186
rect 23 185 24 186
rect 22 185 23 186
rect 21 185 22 186
rect 20 185 21 186
rect 19 185 20 186
rect 18 185 19 186
rect 17 185 18 186
rect 16 185 17 186
rect 15 185 16 186
rect 14 185 15 186
rect 13 185 14 186
rect 12 185 13 186
rect 431 186 432 187
rect 430 186 431 187
rect 429 186 430 187
rect 428 186 429 187
rect 427 186 428 187
rect 426 186 427 187
rect 425 186 426 187
rect 424 186 425 187
rect 423 186 424 187
rect 422 186 423 187
rect 421 186 422 187
rect 420 186 421 187
rect 419 186 420 187
rect 418 186 419 187
rect 417 186 418 187
rect 396 186 397 187
rect 395 186 396 187
rect 333 186 334 187
rect 332 186 333 187
rect 331 186 332 187
rect 330 186 331 187
rect 329 186 330 187
rect 328 186 329 187
rect 327 186 328 187
rect 326 186 327 187
rect 325 186 326 187
rect 324 186 325 187
rect 323 186 324 187
rect 322 186 323 187
rect 321 186 322 187
rect 320 186 321 187
rect 319 186 320 187
rect 318 186 319 187
rect 317 186 318 187
rect 316 186 317 187
rect 315 186 316 187
rect 314 186 315 187
rect 313 186 314 187
rect 312 186 313 187
rect 311 186 312 187
rect 310 186 311 187
rect 309 186 310 187
rect 308 186 309 187
rect 307 186 308 187
rect 306 186 307 187
rect 305 186 306 187
rect 304 186 305 187
rect 303 186 304 187
rect 302 186 303 187
rect 301 186 302 187
rect 300 186 301 187
rect 299 186 300 187
rect 298 186 299 187
rect 297 186 298 187
rect 296 186 297 187
rect 295 186 296 187
rect 294 186 295 187
rect 293 186 294 187
rect 292 186 293 187
rect 291 186 292 187
rect 290 186 291 187
rect 289 186 290 187
rect 288 186 289 187
rect 287 186 288 187
rect 286 186 287 187
rect 285 186 286 187
rect 284 186 285 187
rect 283 186 284 187
rect 282 186 283 187
rect 259 186 260 187
rect 258 186 259 187
rect 257 186 258 187
rect 256 186 257 187
rect 255 186 256 187
rect 254 186 255 187
rect 253 186 254 187
rect 252 186 253 187
rect 251 186 252 187
rect 250 186 251 187
rect 249 186 250 187
rect 248 186 249 187
rect 247 186 248 187
rect 246 186 247 187
rect 245 186 246 187
rect 244 186 245 187
rect 243 186 244 187
rect 242 186 243 187
rect 241 186 242 187
rect 240 186 241 187
rect 239 186 240 187
rect 238 186 239 187
rect 237 186 238 187
rect 236 186 237 187
rect 235 186 236 187
rect 234 186 235 187
rect 233 186 234 187
rect 232 186 233 187
rect 231 186 232 187
rect 230 186 231 187
rect 229 186 230 187
rect 228 186 229 187
rect 227 186 228 187
rect 226 186 227 187
rect 225 186 226 187
rect 224 186 225 187
rect 223 186 224 187
rect 222 186 223 187
rect 221 186 222 187
rect 220 186 221 187
rect 219 186 220 187
rect 197 186 198 187
rect 196 186 197 187
rect 195 186 196 187
rect 194 186 195 187
rect 193 186 194 187
rect 192 186 193 187
rect 191 186 192 187
rect 190 186 191 187
rect 189 186 190 187
rect 188 186 189 187
rect 187 186 188 187
rect 186 186 187 187
rect 185 186 186 187
rect 184 186 185 187
rect 183 186 184 187
rect 182 186 183 187
rect 181 186 182 187
rect 180 186 181 187
rect 179 186 180 187
rect 178 186 179 187
rect 177 186 178 187
rect 176 186 177 187
rect 175 186 176 187
rect 174 186 175 187
rect 173 186 174 187
rect 172 186 173 187
rect 171 186 172 187
rect 170 186 171 187
rect 169 186 170 187
rect 168 186 169 187
rect 167 186 168 187
rect 166 186 167 187
rect 165 186 166 187
rect 164 186 165 187
rect 163 186 164 187
rect 162 186 163 187
rect 161 186 162 187
rect 160 186 161 187
rect 159 186 160 187
rect 158 186 159 187
rect 157 186 158 187
rect 156 186 157 187
rect 155 186 156 187
rect 154 186 155 187
rect 153 186 154 187
rect 152 186 153 187
rect 151 186 152 187
rect 150 186 151 187
rect 149 186 150 187
rect 148 186 149 187
rect 147 186 148 187
rect 146 186 147 187
rect 145 186 146 187
rect 144 186 145 187
rect 143 186 144 187
rect 142 186 143 187
rect 141 186 142 187
rect 140 186 141 187
rect 139 186 140 187
rect 138 186 139 187
rect 137 186 138 187
rect 136 186 137 187
rect 135 186 136 187
rect 134 186 135 187
rect 133 186 134 187
rect 132 186 133 187
rect 131 186 132 187
rect 130 186 131 187
rect 129 186 130 187
rect 128 186 129 187
rect 127 186 128 187
rect 126 186 127 187
rect 125 186 126 187
rect 124 186 125 187
rect 123 186 124 187
rect 122 186 123 187
rect 121 186 122 187
rect 120 186 121 187
rect 119 186 120 187
rect 118 186 119 187
rect 117 186 118 187
rect 116 186 117 187
rect 115 186 116 187
rect 114 186 115 187
rect 113 186 114 187
rect 112 186 113 187
rect 111 186 112 187
rect 110 186 111 187
rect 109 186 110 187
rect 108 186 109 187
rect 107 186 108 187
rect 106 186 107 187
rect 105 186 106 187
rect 104 186 105 187
rect 103 186 104 187
rect 102 186 103 187
rect 101 186 102 187
rect 100 186 101 187
rect 99 186 100 187
rect 98 186 99 187
rect 97 186 98 187
rect 96 186 97 187
rect 95 186 96 187
rect 94 186 95 187
rect 93 186 94 187
rect 92 186 93 187
rect 91 186 92 187
rect 90 186 91 187
rect 89 186 90 187
rect 88 186 89 187
rect 87 186 88 187
rect 86 186 87 187
rect 85 186 86 187
rect 84 186 85 187
rect 83 186 84 187
rect 82 186 83 187
rect 81 186 82 187
rect 80 186 81 187
rect 79 186 80 187
rect 78 186 79 187
rect 77 186 78 187
rect 76 186 77 187
rect 75 186 76 187
rect 74 186 75 187
rect 73 186 74 187
rect 72 186 73 187
rect 71 186 72 187
rect 70 186 71 187
rect 25 186 26 187
rect 24 186 25 187
rect 23 186 24 187
rect 22 186 23 187
rect 21 186 22 187
rect 20 186 21 187
rect 19 186 20 187
rect 18 186 19 187
rect 17 186 18 187
rect 16 186 17 187
rect 15 186 16 187
rect 14 186 15 187
rect 13 186 14 187
rect 12 186 13 187
rect 432 187 433 188
rect 431 187 432 188
rect 430 187 431 188
rect 429 187 430 188
rect 428 187 429 188
rect 427 187 428 188
rect 426 187 427 188
rect 425 187 426 188
rect 424 187 425 188
rect 423 187 424 188
rect 422 187 423 188
rect 421 187 422 188
rect 420 187 421 188
rect 419 187 420 188
rect 418 187 419 188
rect 397 187 398 188
rect 396 187 397 188
rect 395 187 396 188
rect 335 187 336 188
rect 334 187 335 188
rect 333 187 334 188
rect 332 187 333 188
rect 331 187 332 188
rect 330 187 331 188
rect 329 187 330 188
rect 328 187 329 188
rect 327 187 328 188
rect 326 187 327 188
rect 325 187 326 188
rect 324 187 325 188
rect 323 187 324 188
rect 322 187 323 188
rect 321 187 322 188
rect 320 187 321 188
rect 319 187 320 188
rect 318 187 319 188
rect 317 187 318 188
rect 316 187 317 188
rect 315 187 316 188
rect 314 187 315 188
rect 313 187 314 188
rect 312 187 313 188
rect 311 187 312 188
rect 310 187 311 188
rect 309 187 310 188
rect 308 187 309 188
rect 307 187 308 188
rect 306 187 307 188
rect 305 187 306 188
rect 304 187 305 188
rect 303 187 304 188
rect 302 187 303 188
rect 301 187 302 188
rect 300 187 301 188
rect 299 187 300 188
rect 298 187 299 188
rect 297 187 298 188
rect 296 187 297 188
rect 295 187 296 188
rect 294 187 295 188
rect 293 187 294 188
rect 292 187 293 188
rect 291 187 292 188
rect 290 187 291 188
rect 289 187 290 188
rect 288 187 289 188
rect 287 187 288 188
rect 286 187 287 188
rect 285 187 286 188
rect 284 187 285 188
rect 283 187 284 188
rect 282 187 283 188
rect 281 187 282 188
rect 280 187 281 188
rect 258 187 259 188
rect 257 187 258 188
rect 256 187 257 188
rect 255 187 256 188
rect 254 187 255 188
rect 253 187 254 188
rect 252 187 253 188
rect 251 187 252 188
rect 250 187 251 188
rect 249 187 250 188
rect 248 187 249 188
rect 247 187 248 188
rect 246 187 247 188
rect 245 187 246 188
rect 244 187 245 188
rect 243 187 244 188
rect 242 187 243 188
rect 241 187 242 188
rect 240 187 241 188
rect 239 187 240 188
rect 238 187 239 188
rect 237 187 238 188
rect 236 187 237 188
rect 235 187 236 188
rect 234 187 235 188
rect 233 187 234 188
rect 232 187 233 188
rect 231 187 232 188
rect 230 187 231 188
rect 229 187 230 188
rect 228 187 229 188
rect 227 187 228 188
rect 226 187 227 188
rect 225 187 226 188
rect 224 187 225 188
rect 223 187 224 188
rect 222 187 223 188
rect 221 187 222 188
rect 220 187 221 188
rect 219 187 220 188
rect 218 187 219 188
rect 196 187 197 188
rect 195 187 196 188
rect 194 187 195 188
rect 193 187 194 188
rect 192 187 193 188
rect 191 187 192 188
rect 190 187 191 188
rect 189 187 190 188
rect 188 187 189 188
rect 187 187 188 188
rect 186 187 187 188
rect 185 187 186 188
rect 184 187 185 188
rect 183 187 184 188
rect 182 187 183 188
rect 181 187 182 188
rect 180 187 181 188
rect 179 187 180 188
rect 178 187 179 188
rect 177 187 178 188
rect 176 187 177 188
rect 175 187 176 188
rect 174 187 175 188
rect 173 187 174 188
rect 172 187 173 188
rect 171 187 172 188
rect 170 187 171 188
rect 169 187 170 188
rect 168 187 169 188
rect 167 187 168 188
rect 166 187 167 188
rect 165 187 166 188
rect 164 187 165 188
rect 163 187 164 188
rect 162 187 163 188
rect 161 187 162 188
rect 160 187 161 188
rect 159 187 160 188
rect 158 187 159 188
rect 157 187 158 188
rect 156 187 157 188
rect 155 187 156 188
rect 154 187 155 188
rect 153 187 154 188
rect 152 187 153 188
rect 151 187 152 188
rect 150 187 151 188
rect 149 187 150 188
rect 148 187 149 188
rect 147 187 148 188
rect 146 187 147 188
rect 145 187 146 188
rect 144 187 145 188
rect 143 187 144 188
rect 142 187 143 188
rect 141 187 142 188
rect 140 187 141 188
rect 139 187 140 188
rect 138 187 139 188
rect 137 187 138 188
rect 136 187 137 188
rect 135 187 136 188
rect 134 187 135 188
rect 133 187 134 188
rect 132 187 133 188
rect 131 187 132 188
rect 130 187 131 188
rect 129 187 130 188
rect 128 187 129 188
rect 127 187 128 188
rect 126 187 127 188
rect 125 187 126 188
rect 124 187 125 188
rect 123 187 124 188
rect 122 187 123 188
rect 121 187 122 188
rect 120 187 121 188
rect 119 187 120 188
rect 118 187 119 188
rect 117 187 118 188
rect 116 187 117 188
rect 115 187 116 188
rect 114 187 115 188
rect 113 187 114 188
rect 112 187 113 188
rect 111 187 112 188
rect 110 187 111 188
rect 109 187 110 188
rect 108 187 109 188
rect 107 187 108 188
rect 106 187 107 188
rect 105 187 106 188
rect 104 187 105 188
rect 103 187 104 188
rect 102 187 103 188
rect 101 187 102 188
rect 100 187 101 188
rect 99 187 100 188
rect 98 187 99 188
rect 97 187 98 188
rect 96 187 97 188
rect 95 187 96 188
rect 94 187 95 188
rect 93 187 94 188
rect 92 187 93 188
rect 91 187 92 188
rect 90 187 91 188
rect 89 187 90 188
rect 88 187 89 188
rect 87 187 88 188
rect 86 187 87 188
rect 85 187 86 188
rect 84 187 85 188
rect 83 187 84 188
rect 82 187 83 188
rect 81 187 82 188
rect 80 187 81 188
rect 79 187 80 188
rect 78 187 79 188
rect 77 187 78 188
rect 76 187 77 188
rect 75 187 76 188
rect 74 187 75 188
rect 73 187 74 188
rect 72 187 73 188
rect 71 187 72 188
rect 70 187 71 188
rect 25 187 26 188
rect 24 187 25 188
rect 23 187 24 188
rect 22 187 23 188
rect 21 187 22 188
rect 20 187 21 188
rect 19 187 20 188
rect 18 187 19 188
rect 17 187 18 188
rect 16 187 17 188
rect 15 187 16 188
rect 14 187 15 188
rect 13 187 14 188
rect 12 187 13 188
rect 434 188 435 189
rect 433 188 434 189
rect 432 188 433 189
rect 431 188 432 189
rect 430 188 431 189
rect 429 188 430 189
rect 428 188 429 189
rect 427 188 428 189
rect 426 188 427 189
rect 425 188 426 189
rect 424 188 425 189
rect 423 188 424 189
rect 422 188 423 189
rect 421 188 422 189
rect 420 188 421 189
rect 419 188 420 189
rect 397 188 398 189
rect 396 188 397 189
rect 395 188 396 189
rect 336 188 337 189
rect 335 188 336 189
rect 334 188 335 189
rect 333 188 334 189
rect 332 188 333 189
rect 331 188 332 189
rect 330 188 331 189
rect 329 188 330 189
rect 328 188 329 189
rect 327 188 328 189
rect 326 188 327 189
rect 325 188 326 189
rect 324 188 325 189
rect 323 188 324 189
rect 322 188 323 189
rect 321 188 322 189
rect 320 188 321 189
rect 319 188 320 189
rect 318 188 319 189
rect 317 188 318 189
rect 316 188 317 189
rect 315 188 316 189
rect 314 188 315 189
rect 313 188 314 189
rect 312 188 313 189
rect 311 188 312 189
rect 310 188 311 189
rect 309 188 310 189
rect 308 188 309 189
rect 307 188 308 189
rect 306 188 307 189
rect 305 188 306 189
rect 304 188 305 189
rect 303 188 304 189
rect 302 188 303 189
rect 301 188 302 189
rect 300 188 301 189
rect 299 188 300 189
rect 298 188 299 189
rect 297 188 298 189
rect 296 188 297 189
rect 295 188 296 189
rect 294 188 295 189
rect 293 188 294 189
rect 292 188 293 189
rect 291 188 292 189
rect 290 188 291 189
rect 289 188 290 189
rect 288 188 289 189
rect 287 188 288 189
rect 286 188 287 189
rect 285 188 286 189
rect 284 188 285 189
rect 283 188 284 189
rect 282 188 283 189
rect 281 188 282 189
rect 280 188 281 189
rect 279 188 280 189
rect 278 188 279 189
rect 257 188 258 189
rect 256 188 257 189
rect 255 188 256 189
rect 254 188 255 189
rect 253 188 254 189
rect 252 188 253 189
rect 251 188 252 189
rect 250 188 251 189
rect 249 188 250 189
rect 248 188 249 189
rect 247 188 248 189
rect 246 188 247 189
rect 245 188 246 189
rect 244 188 245 189
rect 243 188 244 189
rect 242 188 243 189
rect 241 188 242 189
rect 240 188 241 189
rect 239 188 240 189
rect 238 188 239 189
rect 237 188 238 189
rect 236 188 237 189
rect 235 188 236 189
rect 234 188 235 189
rect 233 188 234 189
rect 232 188 233 189
rect 231 188 232 189
rect 230 188 231 189
rect 229 188 230 189
rect 228 188 229 189
rect 227 188 228 189
rect 226 188 227 189
rect 225 188 226 189
rect 224 188 225 189
rect 223 188 224 189
rect 222 188 223 189
rect 221 188 222 189
rect 220 188 221 189
rect 219 188 220 189
rect 218 188 219 189
rect 195 188 196 189
rect 194 188 195 189
rect 193 188 194 189
rect 192 188 193 189
rect 191 188 192 189
rect 190 188 191 189
rect 189 188 190 189
rect 188 188 189 189
rect 187 188 188 189
rect 186 188 187 189
rect 185 188 186 189
rect 184 188 185 189
rect 183 188 184 189
rect 182 188 183 189
rect 181 188 182 189
rect 180 188 181 189
rect 179 188 180 189
rect 178 188 179 189
rect 177 188 178 189
rect 176 188 177 189
rect 175 188 176 189
rect 174 188 175 189
rect 173 188 174 189
rect 172 188 173 189
rect 171 188 172 189
rect 170 188 171 189
rect 169 188 170 189
rect 168 188 169 189
rect 167 188 168 189
rect 166 188 167 189
rect 165 188 166 189
rect 164 188 165 189
rect 163 188 164 189
rect 162 188 163 189
rect 161 188 162 189
rect 160 188 161 189
rect 159 188 160 189
rect 158 188 159 189
rect 157 188 158 189
rect 156 188 157 189
rect 155 188 156 189
rect 154 188 155 189
rect 153 188 154 189
rect 152 188 153 189
rect 151 188 152 189
rect 150 188 151 189
rect 149 188 150 189
rect 148 188 149 189
rect 147 188 148 189
rect 146 188 147 189
rect 145 188 146 189
rect 144 188 145 189
rect 143 188 144 189
rect 142 188 143 189
rect 141 188 142 189
rect 140 188 141 189
rect 139 188 140 189
rect 138 188 139 189
rect 137 188 138 189
rect 136 188 137 189
rect 135 188 136 189
rect 134 188 135 189
rect 133 188 134 189
rect 132 188 133 189
rect 131 188 132 189
rect 130 188 131 189
rect 129 188 130 189
rect 128 188 129 189
rect 127 188 128 189
rect 126 188 127 189
rect 125 188 126 189
rect 124 188 125 189
rect 123 188 124 189
rect 122 188 123 189
rect 121 188 122 189
rect 120 188 121 189
rect 119 188 120 189
rect 118 188 119 189
rect 117 188 118 189
rect 116 188 117 189
rect 115 188 116 189
rect 114 188 115 189
rect 113 188 114 189
rect 112 188 113 189
rect 111 188 112 189
rect 110 188 111 189
rect 109 188 110 189
rect 108 188 109 189
rect 107 188 108 189
rect 106 188 107 189
rect 105 188 106 189
rect 104 188 105 189
rect 103 188 104 189
rect 102 188 103 189
rect 101 188 102 189
rect 100 188 101 189
rect 99 188 100 189
rect 98 188 99 189
rect 97 188 98 189
rect 96 188 97 189
rect 95 188 96 189
rect 94 188 95 189
rect 93 188 94 189
rect 92 188 93 189
rect 91 188 92 189
rect 90 188 91 189
rect 89 188 90 189
rect 88 188 89 189
rect 87 188 88 189
rect 86 188 87 189
rect 85 188 86 189
rect 84 188 85 189
rect 83 188 84 189
rect 82 188 83 189
rect 81 188 82 189
rect 80 188 81 189
rect 79 188 80 189
rect 78 188 79 189
rect 77 188 78 189
rect 76 188 77 189
rect 75 188 76 189
rect 74 188 75 189
rect 73 188 74 189
rect 72 188 73 189
rect 71 188 72 189
rect 70 188 71 189
rect 26 188 27 189
rect 25 188 26 189
rect 24 188 25 189
rect 23 188 24 189
rect 22 188 23 189
rect 21 188 22 189
rect 20 188 21 189
rect 19 188 20 189
rect 18 188 19 189
rect 17 188 18 189
rect 16 188 17 189
rect 15 188 16 189
rect 14 188 15 189
rect 13 188 14 189
rect 12 188 13 189
rect 435 189 436 190
rect 434 189 435 190
rect 433 189 434 190
rect 432 189 433 190
rect 431 189 432 190
rect 430 189 431 190
rect 429 189 430 190
rect 428 189 429 190
rect 427 189 428 190
rect 426 189 427 190
rect 425 189 426 190
rect 424 189 425 190
rect 423 189 424 190
rect 422 189 423 190
rect 421 189 422 190
rect 397 189 398 190
rect 396 189 397 190
rect 395 189 396 190
rect 338 189 339 190
rect 337 189 338 190
rect 336 189 337 190
rect 335 189 336 190
rect 334 189 335 190
rect 333 189 334 190
rect 332 189 333 190
rect 331 189 332 190
rect 330 189 331 190
rect 329 189 330 190
rect 328 189 329 190
rect 327 189 328 190
rect 326 189 327 190
rect 325 189 326 190
rect 324 189 325 190
rect 323 189 324 190
rect 322 189 323 190
rect 321 189 322 190
rect 320 189 321 190
rect 319 189 320 190
rect 318 189 319 190
rect 317 189 318 190
rect 316 189 317 190
rect 315 189 316 190
rect 314 189 315 190
rect 313 189 314 190
rect 312 189 313 190
rect 311 189 312 190
rect 310 189 311 190
rect 309 189 310 190
rect 308 189 309 190
rect 307 189 308 190
rect 306 189 307 190
rect 305 189 306 190
rect 304 189 305 190
rect 303 189 304 190
rect 302 189 303 190
rect 301 189 302 190
rect 300 189 301 190
rect 299 189 300 190
rect 298 189 299 190
rect 297 189 298 190
rect 296 189 297 190
rect 295 189 296 190
rect 294 189 295 190
rect 293 189 294 190
rect 292 189 293 190
rect 291 189 292 190
rect 290 189 291 190
rect 289 189 290 190
rect 288 189 289 190
rect 287 189 288 190
rect 286 189 287 190
rect 285 189 286 190
rect 284 189 285 190
rect 283 189 284 190
rect 282 189 283 190
rect 281 189 282 190
rect 280 189 281 190
rect 279 189 280 190
rect 278 189 279 190
rect 277 189 278 190
rect 276 189 277 190
rect 257 189 258 190
rect 256 189 257 190
rect 255 189 256 190
rect 254 189 255 190
rect 253 189 254 190
rect 252 189 253 190
rect 251 189 252 190
rect 250 189 251 190
rect 249 189 250 190
rect 248 189 249 190
rect 247 189 248 190
rect 246 189 247 190
rect 245 189 246 190
rect 244 189 245 190
rect 243 189 244 190
rect 242 189 243 190
rect 241 189 242 190
rect 240 189 241 190
rect 239 189 240 190
rect 238 189 239 190
rect 237 189 238 190
rect 236 189 237 190
rect 235 189 236 190
rect 234 189 235 190
rect 233 189 234 190
rect 232 189 233 190
rect 231 189 232 190
rect 230 189 231 190
rect 229 189 230 190
rect 228 189 229 190
rect 227 189 228 190
rect 226 189 227 190
rect 225 189 226 190
rect 224 189 225 190
rect 223 189 224 190
rect 222 189 223 190
rect 221 189 222 190
rect 220 189 221 190
rect 219 189 220 190
rect 218 189 219 190
rect 217 189 218 190
rect 194 189 195 190
rect 193 189 194 190
rect 192 189 193 190
rect 191 189 192 190
rect 190 189 191 190
rect 189 189 190 190
rect 188 189 189 190
rect 187 189 188 190
rect 186 189 187 190
rect 185 189 186 190
rect 184 189 185 190
rect 183 189 184 190
rect 182 189 183 190
rect 181 189 182 190
rect 180 189 181 190
rect 179 189 180 190
rect 178 189 179 190
rect 177 189 178 190
rect 176 189 177 190
rect 175 189 176 190
rect 174 189 175 190
rect 173 189 174 190
rect 172 189 173 190
rect 171 189 172 190
rect 170 189 171 190
rect 169 189 170 190
rect 168 189 169 190
rect 167 189 168 190
rect 166 189 167 190
rect 165 189 166 190
rect 164 189 165 190
rect 163 189 164 190
rect 162 189 163 190
rect 161 189 162 190
rect 160 189 161 190
rect 159 189 160 190
rect 158 189 159 190
rect 157 189 158 190
rect 156 189 157 190
rect 155 189 156 190
rect 154 189 155 190
rect 153 189 154 190
rect 152 189 153 190
rect 151 189 152 190
rect 150 189 151 190
rect 149 189 150 190
rect 148 189 149 190
rect 147 189 148 190
rect 146 189 147 190
rect 145 189 146 190
rect 144 189 145 190
rect 143 189 144 190
rect 142 189 143 190
rect 141 189 142 190
rect 140 189 141 190
rect 139 189 140 190
rect 138 189 139 190
rect 137 189 138 190
rect 136 189 137 190
rect 135 189 136 190
rect 134 189 135 190
rect 133 189 134 190
rect 132 189 133 190
rect 131 189 132 190
rect 130 189 131 190
rect 129 189 130 190
rect 128 189 129 190
rect 127 189 128 190
rect 126 189 127 190
rect 125 189 126 190
rect 124 189 125 190
rect 123 189 124 190
rect 122 189 123 190
rect 121 189 122 190
rect 120 189 121 190
rect 119 189 120 190
rect 118 189 119 190
rect 117 189 118 190
rect 116 189 117 190
rect 115 189 116 190
rect 114 189 115 190
rect 113 189 114 190
rect 112 189 113 190
rect 111 189 112 190
rect 110 189 111 190
rect 109 189 110 190
rect 108 189 109 190
rect 107 189 108 190
rect 106 189 107 190
rect 105 189 106 190
rect 104 189 105 190
rect 103 189 104 190
rect 102 189 103 190
rect 101 189 102 190
rect 100 189 101 190
rect 99 189 100 190
rect 98 189 99 190
rect 97 189 98 190
rect 96 189 97 190
rect 95 189 96 190
rect 94 189 95 190
rect 93 189 94 190
rect 92 189 93 190
rect 91 189 92 190
rect 90 189 91 190
rect 89 189 90 190
rect 88 189 89 190
rect 87 189 88 190
rect 86 189 87 190
rect 85 189 86 190
rect 84 189 85 190
rect 83 189 84 190
rect 82 189 83 190
rect 81 189 82 190
rect 80 189 81 190
rect 79 189 80 190
rect 78 189 79 190
rect 77 189 78 190
rect 76 189 77 190
rect 75 189 76 190
rect 74 189 75 190
rect 73 189 74 190
rect 72 189 73 190
rect 71 189 72 190
rect 70 189 71 190
rect 26 189 27 190
rect 25 189 26 190
rect 24 189 25 190
rect 23 189 24 190
rect 22 189 23 190
rect 21 189 22 190
rect 20 189 21 190
rect 19 189 20 190
rect 18 189 19 190
rect 17 189 18 190
rect 16 189 17 190
rect 15 189 16 190
rect 14 189 15 190
rect 13 189 14 190
rect 12 189 13 190
rect 480 190 481 191
rect 436 190 437 191
rect 435 190 436 191
rect 434 190 435 191
rect 433 190 434 191
rect 432 190 433 191
rect 431 190 432 191
rect 430 190 431 191
rect 429 190 430 191
rect 428 190 429 191
rect 427 190 428 191
rect 426 190 427 191
rect 425 190 426 191
rect 424 190 425 191
rect 423 190 424 191
rect 422 190 423 191
rect 397 190 398 191
rect 396 190 397 191
rect 395 190 396 191
rect 339 190 340 191
rect 338 190 339 191
rect 337 190 338 191
rect 336 190 337 191
rect 335 190 336 191
rect 334 190 335 191
rect 333 190 334 191
rect 332 190 333 191
rect 331 190 332 191
rect 330 190 331 191
rect 329 190 330 191
rect 328 190 329 191
rect 327 190 328 191
rect 326 190 327 191
rect 325 190 326 191
rect 324 190 325 191
rect 323 190 324 191
rect 322 190 323 191
rect 321 190 322 191
rect 320 190 321 191
rect 319 190 320 191
rect 318 190 319 191
rect 317 190 318 191
rect 316 190 317 191
rect 315 190 316 191
rect 314 190 315 191
rect 313 190 314 191
rect 312 190 313 191
rect 311 190 312 191
rect 310 190 311 191
rect 309 190 310 191
rect 308 190 309 191
rect 307 190 308 191
rect 306 190 307 191
rect 305 190 306 191
rect 304 190 305 191
rect 303 190 304 191
rect 302 190 303 191
rect 301 190 302 191
rect 300 190 301 191
rect 299 190 300 191
rect 298 190 299 191
rect 297 190 298 191
rect 296 190 297 191
rect 295 190 296 191
rect 294 190 295 191
rect 293 190 294 191
rect 292 190 293 191
rect 291 190 292 191
rect 290 190 291 191
rect 289 190 290 191
rect 288 190 289 191
rect 287 190 288 191
rect 286 190 287 191
rect 285 190 286 191
rect 284 190 285 191
rect 283 190 284 191
rect 282 190 283 191
rect 281 190 282 191
rect 280 190 281 191
rect 279 190 280 191
rect 278 190 279 191
rect 277 190 278 191
rect 276 190 277 191
rect 275 190 276 191
rect 256 190 257 191
rect 255 190 256 191
rect 254 190 255 191
rect 253 190 254 191
rect 252 190 253 191
rect 251 190 252 191
rect 250 190 251 191
rect 249 190 250 191
rect 248 190 249 191
rect 247 190 248 191
rect 246 190 247 191
rect 245 190 246 191
rect 244 190 245 191
rect 243 190 244 191
rect 242 190 243 191
rect 241 190 242 191
rect 240 190 241 191
rect 239 190 240 191
rect 238 190 239 191
rect 237 190 238 191
rect 236 190 237 191
rect 235 190 236 191
rect 234 190 235 191
rect 233 190 234 191
rect 232 190 233 191
rect 231 190 232 191
rect 230 190 231 191
rect 229 190 230 191
rect 228 190 229 191
rect 227 190 228 191
rect 226 190 227 191
rect 225 190 226 191
rect 224 190 225 191
rect 223 190 224 191
rect 222 190 223 191
rect 221 190 222 191
rect 220 190 221 191
rect 219 190 220 191
rect 218 190 219 191
rect 217 190 218 191
rect 216 190 217 191
rect 193 190 194 191
rect 192 190 193 191
rect 191 190 192 191
rect 190 190 191 191
rect 189 190 190 191
rect 188 190 189 191
rect 187 190 188 191
rect 186 190 187 191
rect 185 190 186 191
rect 184 190 185 191
rect 183 190 184 191
rect 182 190 183 191
rect 181 190 182 191
rect 180 190 181 191
rect 179 190 180 191
rect 178 190 179 191
rect 177 190 178 191
rect 176 190 177 191
rect 175 190 176 191
rect 174 190 175 191
rect 173 190 174 191
rect 172 190 173 191
rect 171 190 172 191
rect 170 190 171 191
rect 169 190 170 191
rect 168 190 169 191
rect 167 190 168 191
rect 166 190 167 191
rect 165 190 166 191
rect 164 190 165 191
rect 163 190 164 191
rect 162 190 163 191
rect 161 190 162 191
rect 160 190 161 191
rect 159 190 160 191
rect 158 190 159 191
rect 157 190 158 191
rect 156 190 157 191
rect 155 190 156 191
rect 154 190 155 191
rect 153 190 154 191
rect 152 190 153 191
rect 151 190 152 191
rect 150 190 151 191
rect 149 190 150 191
rect 148 190 149 191
rect 147 190 148 191
rect 146 190 147 191
rect 145 190 146 191
rect 144 190 145 191
rect 143 190 144 191
rect 142 190 143 191
rect 141 190 142 191
rect 140 190 141 191
rect 139 190 140 191
rect 138 190 139 191
rect 137 190 138 191
rect 136 190 137 191
rect 135 190 136 191
rect 134 190 135 191
rect 133 190 134 191
rect 132 190 133 191
rect 131 190 132 191
rect 130 190 131 191
rect 129 190 130 191
rect 128 190 129 191
rect 127 190 128 191
rect 126 190 127 191
rect 125 190 126 191
rect 124 190 125 191
rect 123 190 124 191
rect 122 190 123 191
rect 121 190 122 191
rect 120 190 121 191
rect 119 190 120 191
rect 118 190 119 191
rect 117 190 118 191
rect 116 190 117 191
rect 115 190 116 191
rect 114 190 115 191
rect 113 190 114 191
rect 112 190 113 191
rect 111 190 112 191
rect 110 190 111 191
rect 109 190 110 191
rect 108 190 109 191
rect 107 190 108 191
rect 106 190 107 191
rect 105 190 106 191
rect 104 190 105 191
rect 103 190 104 191
rect 102 190 103 191
rect 101 190 102 191
rect 100 190 101 191
rect 99 190 100 191
rect 98 190 99 191
rect 97 190 98 191
rect 96 190 97 191
rect 95 190 96 191
rect 94 190 95 191
rect 93 190 94 191
rect 92 190 93 191
rect 91 190 92 191
rect 90 190 91 191
rect 89 190 90 191
rect 88 190 89 191
rect 87 190 88 191
rect 86 190 87 191
rect 85 190 86 191
rect 84 190 85 191
rect 83 190 84 191
rect 82 190 83 191
rect 81 190 82 191
rect 80 190 81 191
rect 79 190 80 191
rect 78 190 79 191
rect 77 190 78 191
rect 76 190 77 191
rect 75 190 76 191
rect 74 190 75 191
rect 73 190 74 191
rect 72 190 73 191
rect 71 190 72 191
rect 70 190 71 191
rect 69 190 70 191
rect 27 190 28 191
rect 26 190 27 191
rect 25 190 26 191
rect 24 190 25 191
rect 23 190 24 191
rect 22 190 23 191
rect 21 190 22 191
rect 20 190 21 191
rect 19 190 20 191
rect 18 190 19 191
rect 17 190 18 191
rect 16 190 17 191
rect 15 190 16 191
rect 14 190 15 191
rect 13 190 14 191
rect 12 190 13 191
rect 480 191 481 192
rect 460 191 461 192
rect 437 191 438 192
rect 436 191 437 192
rect 435 191 436 192
rect 434 191 435 192
rect 433 191 434 192
rect 432 191 433 192
rect 431 191 432 192
rect 430 191 431 192
rect 429 191 430 192
rect 428 191 429 192
rect 427 191 428 192
rect 426 191 427 192
rect 425 191 426 192
rect 424 191 425 192
rect 423 191 424 192
rect 398 191 399 192
rect 397 191 398 192
rect 396 191 397 192
rect 395 191 396 192
rect 340 191 341 192
rect 339 191 340 192
rect 338 191 339 192
rect 337 191 338 192
rect 336 191 337 192
rect 335 191 336 192
rect 334 191 335 192
rect 333 191 334 192
rect 332 191 333 192
rect 331 191 332 192
rect 330 191 331 192
rect 329 191 330 192
rect 328 191 329 192
rect 327 191 328 192
rect 326 191 327 192
rect 325 191 326 192
rect 324 191 325 192
rect 323 191 324 192
rect 322 191 323 192
rect 321 191 322 192
rect 320 191 321 192
rect 319 191 320 192
rect 318 191 319 192
rect 317 191 318 192
rect 316 191 317 192
rect 315 191 316 192
rect 314 191 315 192
rect 313 191 314 192
rect 312 191 313 192
rect 311 191 312 192
rect 310 191 311 192
rect 309 191 310 192
rect 308 191 309 192
rect 307 191 308 192
rect 306 191 307 192
rect 305 191 306 192
rect 304 191 305 192
rect 303 191 304 192
rect 302 191 303 192
rect 301 191 302 192
rect 300 191 301 192
rect 299 191 300 192
rect 298 191 299 192
rect 297 191 298 192
rect 296 191 297 192
rect 295 191 296 192
rect 294 191 295 192
rect 293 191 294 192
rect 292 191 293 192
rect 291 191 292 192
rect 290 191 291 192
rect 289 191 290 192
rect 288 191 289 192
rect 287 191 288 192
rect 286 191 287 192
rect 285 191 286 192
rect 284 191 285 192
rect 283 191 284 192
rect 282 191 283 192
rect 281 191 282 192
rect 280 191 281 192
rect 279 191 280 192
rect 278 191 279 192
rect 277 191 278 192
rect 276 191 277 192
rect 275 191 276 192
rect 274 191 275 192
rect 273 191 274 192
rect 255 191 256 192
rect 254 191 255 192
rect 253 191 254 192
rect 252 191 253 192
rect 251 191 252 192
rect 250 191 251 192
rect 249 191 250 192
rect 248 191 249 192
rect 247 191 248 192
rect 246 191 247 192
rect 245 191 246 192
rect 244 191 245 192
rect 243 191 244 192
rect 242 191 243 192
rect 241 191 242 192
rect 240 191 241 192
rect 239 191 240 192
rect 238 191 239 192
rect 237 191 238 192
rect 236 191 237 192
rect 235 191 236 192
rect 234 191 235 192
rect 233 191 234 192
rect 232 191 233 192
rect 231 191 232 192
rect 230 191 231 192
rect 229 191 230 192
rect 228 191 229 192
rect 227 191 228 192
rect 226 191 227 192
rect 225 191 226 192
rect 224 191 225 192
rect 223 191 224 192
rect 222 191 223 192
rect 221 191 222 192
rect 220 191 221 192
rect 219 191 220 192
rect 218 191 219 192
rect 217 191 218 192
rect 216 191 217 192
rect 192 191 193 192
rect 191 191 192 192
rect 190 191 191 192
rect 189 191 190 192
rect 188 191 189 192
rect 187 191 188 192
rect 186 191 187 192
rect 185 191 186 192
rect 184 191 185 192
rect 183 191 184 192
rect 182 191 183 192
rect 181 191 182 192
rect 180 191 181 192
rect 179 191 180 192
rect 178 191 179 192
rect 177 191 178 192
rect 176 191 177 192
rect 175 191 176 192
rect 174 191 175 192
rect 173 191 174 192
rect 172 191 173 192
rect 171 191 172 192
rect 170 191 171 192
rect 169 191 170 192
rect 168 191 169 192
rect 167 191 168 192
rect 166 191 167 192
rect 165 191 166 192
rect 164 191 165 192
rect 163 191 164 192
rect 162 191 163 192
rect 161 191 162 192
rect 160 191 161 192
rect 159 191 160 192
rect 158 191 159 192
rect 157 191 158 192
rect 156 191 157 192
rect 155 191 156 192
rect 154 191 155 192
rect 153 191 154 192
rect 152 191 153 192
rect 151 191 152 192
rect 150 191 151 192
rect 149 191 150 192
rect 148 191 149 192
rect 147 191 148 192
rect 146 191 147 192
rect 145 191 146 192
rect 144 191 145 192
rect 143 191 144 192
rect 142 191 143 192
rect 141 191 142 192
rect 140 191 141 192
rect 139 191 140 192
rect 138 191 139 192
rect 137 191 138 192
rect 136 191 137 192
rect 135 191 136 192
rect 134 191 135 192
rect 133 191 134 192
rect 132 191 133 192
rect 131 191 132 192
rect 130 191 131 192
rect 129 191 130 192
rect 128 191 129 192
rect 127 191 128 192
rect 126 191 127 192
rect 125 191 126 192
rect 124 191 125 192
rect 123 191 124 192
rect 122 191 123 192
rect 121 191 122 192
rect 120 191 121 192
rect 119 191 120 192
rect 118 191 119 192
rect 117 191 118 192
rect 116 191 117 192
rect 115 191 116 192
rect 114 191 115 192
rect 113 191 114 192
rect 112 191 113 192
rect 111 191 112 192
rect 110 191 111 192
rect 109 191 110 192
rect 108 191 109 192
rect 107 191 108 192
rect 106 191 107 192
rect 105 191 106 192
rect 104 191 105 192
rect 103 191 104 192
rect 102 191 103 192
rect 101 191 102 192
rect 100 191 101 192
rect 99 191 100 192
rect 98 191 99 192
rect 97 191 98 192
rect 96 191 97 192
rect 95 191 96 192
rect 94 191 95 192
rect 93 191 94 192
rect 92 191 93 192
rect 91 191 92 192
rect 90 191 91 192
rect 89 191 90 192
rect 88 191 89 192
rect 87 191 88 192
rect 86 191 87 192
rect 85 191 86 192
rect 84 191 85 192
rect 83 191 84 192
rect 82 191 83 192
rect 81 191 82 192
rect 80 191 81 192
rect 79 191 80 192
rect 78 191 79 192
rect 77 191 78 192
rect 76 191 77 192
rect 75 191 76 192
rect 74 191 75 192
rect 73 191 74 192
rect 72 191 73 192
rect 71 191 72 192
rect 70 191 71 192
rect 69 191 70 192
rect 28 191 29 192
rect 27 191 28 192
rect 26 191 27 192
rect 25 191 26 192
rect 24 191 25 192
rect 23 191 24 192
rect 22 191 23 192
rect 21 191 22 192
rect 20 191 21 192
rect 19 191 20 192
rect 18 191 19 192
rect 17 191 18 192
rect 16 191 17 192
rect 15 191 16 192
rect 14 191 15 192
rect 13 191 14 192
rect 12 191 13 192
rect 480 192 481 193
rect 479 192 480 193
rect 460 192 461 193
rect 438 192 439 193
rect 437 192 438 193
rect 436 192 437 193
rect 435 192 436 193
rect 434 192 435 193
rect 433 192 434 193
rect 432 192 433 193
rect 431 192 432 193
rect 430 192 431 193
rect 429 192 430 193
rect 428 192 429 193
rect 427 192 428 193
rect 426 192 427 193
rect 425 192 426 193
rect 424 192 425 193
rect 399 192 400 193
rect 398 192 399 193
rect 397 192 398 193
rect 396 192 397 193
rect 395 192 396 193
rect 341 192 342 193
rect 340 192 341 193
rect 339 192 340 193
rect 338 192 339 193
rect 337 192 338 193
rect 336 192 337 193
rect 335 192 336 193
rect 334 192 335 193
rect 333 192 334 193
rect 332 192 333 193
rect 331 192 332 193
rect 330 192 331 193
rect 329 192 330 193
rect 328 192 329 193
rect 327 192 328 193
rect 326 192 327 193
rect 325 192 326 193
rect 324 192 325 193
rect 323 192 324 193
rect 322 192 323 193
rect 321 192 322 193
rect 320 192 321 193
rect 319 192 320 193
rect 318 192 319 193
rect 317 192 318 193
rect 316 192 317 193
rect 315 192 316 193
rect 314 192 315 193
rect 313 192 314 193
rect 312 192 313 193
rect 311 192 312 193
rect 310 192 311 193
rect 309 192 310 193
rect 308 192 309 193
rect 307 192 308 193
rect 306 192 307 193
rect 305 192 306 193
rect 304 192 305 193
rect 303 192 304 193
rect 302 192 303 193
rect 301 192 302 193
rect 300 192 301 193
rect 299 192 300 193
rect 298 192 299 193
rect 297 192 298 193
rect 296 192 297 193
rect 295 192 296 193
rect 294 192 295 193
rect 293 192 294 193
rect 292 192 293 193
rect 291 192 292 193
rect 290 192 291 193
rect 289 192 290 193
rect 288 192 289 193
rect 287 192 288 193
rect 286 192 287 193
rect 285 192 286 193
rect 284 192 285 193
rect 283 192 284 193
rect 282 192 283 193
rect 281 192 282 193
rect 280 192 281 193
rect 279 192 280 193
rect 278 192 279 193
rect 277 192 278 193
rect 276 192 277 193
rect 275 192 276 193
rect 274 192 275 193
rect 273 192 274 193
rect 272 192 273 193
rect 255 192 256 193
rect 254 192 255 193
rect 253 192 254 193
rect 252 192 253 193
rect 251 192 252 193
rect 250 192 251 193
rect 249 192 250 193
rect 248 192 249 193
rect 247 192 248 193
rect 246 192 247 193
rect 245 192 246 193
rect 244 192 245 193
rect 243 192 244 193
rect 242 192 243 193
rect 241 192 242 193
rect 240 192 241 193
rect 239 192 240 193
rect 238 192 239 193
rect 237 192 238 193
rect 236 192 237 193
rect 235 192 236 193
rect 234 192 235 193
rect 233 192 234 193
rect 232 192 233 193
rect 231 192 232 193
rect 230 192 231 193
rect 229 192 230 193
rect 228 192 229 193
rect 227 192 228 193
rect 226 192 227 193
rect 225 192 226 193
rect 224 192 225 193
rect 223 192 224 193
rect 222 192 223 193
rect 221 192 222 193
rect 220 192 221 193
rect 219 192 220 193
rect 218 192 219 193
rect 217 192 218 193
rect 216 192 217 193
rect 215 192 216 193
rect 191 192 192 193
rect 190 192 191 193
rect 189 192 190 193
rect 188 192 189 193
rect 187 192 188 193
rect 186 192 187 193
rect 185 192 186 193
rect 184 192 185 193
rect 183 192 184 193
rect 182 192 183 193
rect 181 192 182 193
rect 180 192 181 193
rect 179 192 180 193
rect 178 192 179 193
rect 177 192 178 193
rect 176 192 177 193
rect 175 192 176 193
rect 174 192 175 193
rect 173 192 174 193
rect 172 192 173 193
rect 171 192 172 193
rect 170 192 171 193
rect 169 192 170 193
rect 168 192 169 193
rect 167 192 168 193
rect 166 192 167 193
rect 165 192 166 193
rect 164 192 165 193
rect 163 192 164 193
rect 162 192 163 193
rect 161 192 162 193
rect 160 192 161 193
rect 159 192 160 193
rect 158 192 159 193
rect 157 192 158 193
rect 156 192 157 193
rect 155 192 156 193
rect 154 192 155 193
rect 153 192 154 193
rect 152 192 153 193
rect 151 192 152 193
rect 150 192 151 193
rect 149 192 150 193
rect 148 192 149 193
rect 147 192 148 193
rect 146 192 147 193
rect 145 192 146 193
rect 144 192 145 193
rect 143 192 144 193
rect 142 192 143 193
rect 141 192 142 193
rect 140 192 141 193
rect 139 192 140 193
rect 138 192 139 193
rect 137 192 138 193
rect 136 192 137 193
rect 135 192 136 193
rect 134 192 135 193
rect 133 192 134 193
rect 132 192 133 193
rect 131 192 132 193
rect 130 192 131 193
rect 129 192 130 193
rect 128 192 129 193
rect 127 192 128 193
rect 126 192 127 193
rect 125 192 126 193
rect 124 192 125 193
rect 123 192 124 193
rect 122 192 123 193
rect 121 192 122 193
rect 120 192 121 193
rect 119 192 120 193
rect 118 192 119 193
rect 117 192 118 193
rect 116 192 117 193
rect 115 192 116 193
rect 114 192 115 193
rect 113 192 114 193
rect 112 192 113 193
rect 111 192 112 193
rect 110 192 111 193
rect 109 192 110 193
rect 108 192 109 193
rect 107 192 108 193
rect 106 192 107 193
rect 105 192 106 193
rect 104 192 105 193
rect 103 192 104 193
rect 102 192 103 193
rect 101 192 102 193
rect 100 192 101 193
rect 99 192 100 193
rect 98 192 99 193
rect 97 192 98 193
rect 96 192 97 193
rect 95 192 96 193
rect 94 192 95 193
rect 93 192 94 193
rect 92 192 93 193
rect 91 192 92 193
rect 90 192 91 193
rect 89 192 90 193
rect 88 192 89 193
rect 87 192 88 193
rect 86 192 87 193
rect 85 192 86 193
rect 84 192 85 193
rect 83 192 84 193
rect 82 192 83 193
rect 81 192 82 193
rect 80 192 81 193
rect 79 192 80 193
rect 78 192 79 193
rect 77 192 78 193
rect 76 192 77 193
rect 75 192 76 193
rect 74 192 75 193
rect 73 192 74 193
rect 72 192 73 193
rect 71 192 72 193
rect 70 192 71 193
rect 69 192 70 193
rect 28 192 29 193
rect 27 192 28 193
rect 26 192 27 193
rect 25 192 26 193
rect 24 192 25 193
rect 23 192 24 193
rect 22 192 23 193
rect 21 192 22 193
rect 20 192 21 193
rect 19 192 20 193
rect 18 192 19 193
rect 17 192 18 193
rect 16 192 17 193
rect 15 192 16 193
rect 14 192 15 193
rect 13 192 14 193
rect 12 192 13 193
rect 480 193 481 194
rect 479 193 480 194
rect 478 193 479 194
rect 477 193 478 194
rect 476 193 477 194
rect 475 193 476 194
rect 474 193 475 194
rect 473 193 474 194
rect 472 193 473 194
rect 471 193 472 194
rect 470 193 471 194
rect 469 193 470 194
rect 468 193 469 194
rect 467 193 468 194
rect 466 193 467 194
rect 465 193 466 194
rect 464 193 465 194
rect 463 193 464 194
rect 462 193 463 194
rect 461 193 462 194
rect 460 193 461 194
rect 440 193 441 194
rect 439 193 440 194
rect 438 193 439 194
rect 437 193 438 194
rect 436 193 437 194
rect 435 193 436 194
rect 434 193 435 194
rect 433 193 434 194
rect 432 193 433 194
rect 431 193 432 194
rect 430 193 431 194
rect 429 193 430 194
rect 428 193 429 194
rect 427 193 428 194
rect 426 193 427 194
rect 425 193 426 194
rect 405 193 406 194
rect 404 193 405 194
rect 403 193 404 194
rect 402 193 403 194
rect 401 193 402 194
rect 400 193 401 194
rect 399 193 400 194
rect 398 193 399 194
rect 397 193 398 194
rect 396 193 397 194
rect 395 193 396 194
rect 342 193 343 194
rect 341 193 342 194
rect 340 193 341 194
rect 339 193 340 194
rect 338 193 339 194
rect 337 193 338 194
rect 336 193 337 194
rect 335 193 336 194
rect 334 193 335 194
rect 333 193 334 194
rect 332 193 333 194
rect 331 193 332 194
rect 330 193 331 194
rect 329 193 330 194
rect 328 193 329 194
rect 327 193 328 194
rect 326 193 327 194
rect 325 193 326 194
rect 324 193 325 194
rect 323 193 324 194
rect 322 193 323 194
rect 321 193 322 194
rect 320 193 321 194
rect 319 193 320 194
rect 318 193 319 194
rect 317 193 318 194
rect 316 193 317 194
rect 315 193 316 194
rect 314 193 315 194
rect 313 193 314 194
rect 312 193 313 194
rect 311 193 312 194
rect 310 193 311 194
rect 309 193 310 194
rect 308 193 309 194
rect 307 193 308 194
rect 306 193 307 194
rect 305 193 306 194
rect 304 193 305 194
rect 303 193 304 194
rect 302 193 303 194
rect 301 193 302 194
rect 300 193 301 194
rect 299 193 300 194
rect 298 193 299 194
rect 297 193 298 194
rect 296 193 297 194
rect 295 193 296 194
rect 294 193 295 194
rect 293 193 294 194
rect 292 193 293 194
rect 291 193 292 194
rect 290 193 291 194
rect 289 193 290 194
rect 288 193 289 194
rect 287 193 288 194
rect 286 193 287 194
rect 285 193 286 194
rect 284 193 285 194
rect 283 193 284 194
rect 282 193 283 194
rect 281 193 282 194
rect 280 193 281 194
rect 279 193 280 194
rect 278 193 279 194
rect 277 193 278 194
rect 276 193 277 194
rect 275 193 276 194
rect 274 193 275 194
rect 273 193 274 194
rect 272 193 273 194
rect 271 193 272 194
rect 254 193 255 194
rect 253 193 254 194
rect 252 193 253 194
rect 251 193 252 194
rect 250 193 251 194
rect 249 193 250 194
rect 248 193 249 194
rect 247 193 248 194
rect 246 193 247 194
rect 245 193 246 194
rect 244 193 245 194
rect 243 193 244 194
rect 242 193 243 194
rect 241 193 242 194
rect 240 193 241 194
rect 239 193 240 194
rect 238 193 239 194
rect 237 193 238 194
rect 236 193 237 194
rect 235 193 236 194
rect 234 193 235 194
rect 233 193 234 194
rect 232 193 233 194
rect 231 193 232 194
rect 230 193 231 194
rect 229 193 230 194
rect 228 193 229 194
rect 227 193 228 194
rect 226 193 227 194
rect 225 193 226 194
rect 224 193 225 194
rect 223 193 224 194
rect 222 193 223 194
rect 221 193 222 194
rect 220 193 221 194
rect 219 193 220 194
rect 218 193 219 194
rect 217 193 218 194
rect 216 193 217 194
rect 215 193 216 194
rect 214 193 215 194
rect 190 193 191 194
rect 189 193 190 194
rect 188 193 189 194
rect 187 193 188 194
rect 186 193 187 194
rect 185 193 186 194
rect 184 193 185 194
rect 183 193 184 194
rect 182 193 183 194
rect 181 193 182 194
rect 180 193 181 194
rect 179 193 180 194
rect 178 193 179 194
rect 177 193 178 194
rect 176 193 177 194
rect 175 193 176 194
rect 174 193 175 194
rect 173 193 174 194
rect 172 193 173 194
rect 171 193 172 194
rect 170 193 171 194
rect 169 193 170 194
rect 168 193 169 194
rect 167 193 168 194
rect 166 193 167 194
rect 165 193 166 194
rect 164 193 165 194
rect 163 193 164 194
rect 162 193 163 194
rect 161 193 162 194
rect 160 193 161 194
rect 159 193 160 194
rect 158 193 159 194
rect 157 193 158 194
rect 156 193 157 194
rect 155 193 156 194
rect 154 193 155 194
rect 153 193 154 194
rect 152 193 153 194
rect 151 193 152 194
rect 150 193 151 194
rect 149 193 150 194
rect 148 193 149 194
rect 147 193 148 194
rect 146 193 147 194
rect 145 193 146 194
rect 144 193 145 194
rect 143 193 144 194
rect 142 193 143 194
rect 141 193 142 194
rect 140 193 141 194
rect 139 193 140 194
rect 138 193 139 194
rect 137 193 138 194
rect 136 193 137 194
rect 135 193 136 194
rect 134 193 135 194
rect 133 193 134 194
rect 132 193 133 194
rect 131 193 132 194
rect 130 193 131 194
rect 129 193 130 194
rect 128 193 129 194
rect 127 193 128 194
rect 126 193 127 194
rect 125 193 126 194
rect 124 193 125 194
rect 123 193 124 194
rect 122 193 123 194
rect 121 193 122 194
rect 120 193 121 194
rect 119 193 120 194
rect 118 193 119 194
rect 117 193 118 194
rect 116 193 117 194
rect 115 193 116 194
rect 114 193 115 194
rect 113 193 114 194
rect 112 193 113 194
rect 111 193 112 194
rect 110 193 111 194
rect 109 193 110 194
rect 108 193 109 194
rect 107 193 108 194
rect 106 193 107 194
rect 105 193 106 194
rect 104 193 105 194
rect 103 193 104 194
rect 102 193 103 194
rect 101 193 102 194
rect 100 193 101 194
rect 99 193 100 194
rect 98 193 99 194
rect 97 193 98 194
rect 96 193 97 194
rect 95 193 96 194
rect 94 193 95 194
rect 93 193 94 194
rect 92 193 93 194
rect 91 193 92 194
rect 90 193 91 194
rect 89 193 90 194
rect 88 193 89 194
rect 87 193 88 194
rect 86 193 87 194
rect 85 193 86 194
rect 84 193 85 194
rect 83 193 84 194
rect 82 193 83 194
rect 81 193 82 194
rect 80 193 81 194
rect 79 193 80 194
rect 78 193 79 194
rect 77 193 78 194
rect 76 193 77 194
rect 75 193 76 194
rect 74 193 75 194
rect 73 193 74 194
rect 72 193 73 194
rect 71 193 72 194
rect 70 193 71 194
rect 50 193 51 194
rect 49 193 50 194
rect 48 193 49 194
rect 29 193 30 194
rect 28 193 29 194
rect 27 193 28 194
rect 26 193 27 194
rect 25 193 26 194
rect 24 193 25 194
rect 23 193 24 194
rect 22 193 23 194
rect 21 193 22 194
rect 20 193 21 194
rect 19 193 20 194
rect 18 193 19 194
rect 17 193 18 194
rect 16 193 17 194
rect 15 193 16 194
rect 14 193 15 194
rect 13 193 14 194
rect 12 193 13 194
rect 480 194 481 195
rect 479 194 480 195
rect 478 194 479 195
rect 477 194 478 195
rect 476 194 477 195
rect 475 194 476 195
rect 474 194 475 195
rect 473 194 474 195
rect 472 194 473 195
rect 471 194 472 195
rect 470 194 471 195
rect 469 194 470 195
rect 468 194 469 195
rect 467 194 468 195
rect 466 194 467 195
rect 465 194 466 195
rect 464 194 465 195
rect 463 194 464 195
rect 462 194 463 195
rect 461 194 462 195
rect 460 194 461 195
rect 440 194 441 195
rect 439 194 440 195
rect 438 194 439 195
rect 437 194 438 195
rect 436 194 437 195
rect 435 194 436 195
rect 434 194 435 195
rect 433 194 434 195
rect 432 194 433 195
rect 431 194 432 195
rect 430 194 431 195
rect 429 194 430 195
rect 428 194 429 195
rect 427 194 428 195
rect 426 194 427 195
rect 425 194 426 195
rect 424 194 425 195
rect 423 194 424 195
rect 422 194 423 195
rect 421 194 422 195
rect 420 194 421 195
rect 419 194 420 195
rect 418 194 419 195
rect 417 194 418 195
rect 416 194 417 195
rect 415 194 416 195
rect 414 194 415 195
rect 413 194 414 195
rect 412 194 413 195
rect 411 194 412 195
rect 410 194 411 195
rect 409 194 410 195
rect 408 194 409 195
rect 407 194 408 195
rect 406 194 407 195
rect 405 194 406 195
rect 404 194 405 195
rect 403 194 404 195
rect 402 194 403 195
rect 401 194 402 195
rect 400 194 401 195
rect 399 194 400 195
rect 398 194 399 195
rect 397 194 398 195
rect 396 194 397 195
rect 395 194 396 195
rect 343 194 344 195
rect 342 194 343 195
rect 341 194 342 195
rect 340 194 341 195
rect 339 194 340 195
rect 338 194 339 195
rect 337 194 338 195
rect 336 194 337 195
rect 335 194 336 195
rect 334 194 335 195
rect 333 194 334 195
rect 332 194 333 195
rect 331 194 332 195
rect 330 194 331 195
rect 329 194 330 195
rect 328 194 329 195
rect 327 194 328 195
rect 326 194 327 195
rect 325 194 326 195
rect 324 194 325 195
rect 323 194 324 195
rect 322 194 323 195
rect 321 194 322 195
rect 320 194 321 195
rect 319 194 320 195
rect 318 194 319 195
rect 317 194 318 195
rect 316 194 317 195
rect 315 194 316 195
rect 314 194 315 195
rect 313 194 314 195
rect 312 194 313 195
rect 311 194 312 195
rect 310 194 311 195
rect 309 194 310 195
rect 308 194 309 195
rect 307 194 308 195
rect 306 194 307 195
rect 305 194 306 195
rect 304 194 305 195
rect 303 194 304 195
rect 302 194 303 195
rect 301 194 302 195
rect 300 194 301 195
rect 299 194 300 195
rect 298 194 299 195
rect 297 194 298 195
rect 296 194 297 195
rect 295 194 296 195
rect 294 194 295 195
rect 293 194 294 195
rect 292 194 293 195
rect 291 194 292 195
rect 290 194 291 195
rect 289 194 290 195
rect 288 194 289 195
rect 287 194 288 195
rect 286 194 287 195
rect 285 194 286 195
rect 284 194 285 195
rect 283 194 284 195
rect 282 194 283 195
rect 281 194 282 195
rect 280 194 281 195
rect 279 194 280 195
rect 278 194 279 195
rect 277 194 278 195
rect 276 194 277 195
rect 275 194 276 195
rect 274 194 275 195
rect 273 194 274 195
rect 272 194 273 195
rect 271 194 272 195
rect 270 194 271 195
rect 269 194 270 195
rect 254 194 255 195
rect 253 194 254 195
rect 252 194 253 195
rect 251 194 252 195
rect 250 194 251 195
rect 249 194 250 195
rect 248 194 249 195
rect 247 194 248 195
rect 246 194 247 195
rect 245 194 246 195
rect 244 194 245 195
rect 243 194 244 195
rect 242 194 243 195
rect 241 194 242 195
rect 240 194 241 195
rect 239 194 240 195
rect 238 194 239 195
rect 237 194 238 195
rect 236 194 237 195
rect 235 194 236 195
rect 234 194 235 195
rect 233 194 234 195
rect 232 194 233 195
rect 231 194 232 195
rect 230 194 231 195
rect 229 194 230 195
rect 228 194 229 195
rect 227 194 228 195
rect 226 194 227 195
rect 225 194 226 195
rect 224 194 225 195
rect 223 194 224 195
rect 222 194 223 195
rect 221 194 222 195
rect 220 194 221 195
rect 219 194 220 195
rect 218 194 219 195
rect 217 194 218 195
rect 216 194 217 195
rect 215 194 216 195
rect 214 194 215 195
rect 189 194 190 195
rect 188 194 189 195
rect 187 194 188 195
rect 186 194 187 195
rect 185 194 186 195
rect 184 194 185 195
rect 183 194 184 195
rect 182 194 183 195
rect 181 194 182 195
rect 180 194 181 195
rect 179 194 180 195
rect 178 194 179 195
rect 177 194 178 195
rect 176 194 177 195
rect 175 194 176 195
rect 174 194 175 195
rect 173 194 174 195
rect 172 194 173 195
rect 171 194 172 195
rect 170 194 171 195
rect 169 194 170 195
rect 168 194 169 195
rect 167 194 168 195
rect 166 194 167 195
rect 165 194 166 195
rect 164 194 165 195
rect 163 194 164 195
rect 162 194 163 195
rect 161 194 162 195
rect 160 194 161 195
rect 159 194 160 195
rect 158 194 159 195
rect 157 194 158 195
rect 156 194 157 195
rect 155 194 156 195
rect 154 194 155 195
rect 153 194 154 195
rect 152 194 153 195
rect 151 194 152 195
rect 150 194 151 195
rect 149 194 150 195
rect 148 194 149 195
rect 147 194 148 195
rect 146 194 147 195
rect 145 194 146 195
rect 144 194 145 195
rect 143 194 144 195
rect 142 194 143 195
rect 141 194 142 195
rect 140 194 141 195
rect 139 194 140 195
rect 138 194 139 195
rect 137 194 138 195
rect 136 194 137 195
rect 135 194 136 195
rect 134 194 135 195
rect 133 194 134 195
rect 132 194 133 195
rect 131 194 132 195
rect 130 194 131 195
rect 129 194 130 195
rect 128 194 129 195
rect 127 194 128 195
rect 126 194 127 195
rect 125 194 126 195
rect 124 194 125 195
rect 123 194 124 195
rect 122 194 123 195
rect 121 194 122 195
rect 120 194 121 195
rect 119 194 120 195
rect 118 194 119 195
rect 117 194 118 195
rect 116 194 117 195
rect 115 194 116 195
rect 114 194 115 195
rect 113 194 114 195
rect 112 194 113 195
rect 111 194 112 195
rect 110 194 111 195
rect 109 194 110 195
rect 108 194 109 195
rect 107 194 108 195
rect 106 194 107 195
rect 105 194 106 195
rect 104 194 105 195
rect 103 194 104 195
rect 102 194 103 195
rect 101 194 102 195
rect 100 194 101 195
rect 99 194 100 195
rect 98 194 99 195
rect 97 194 98 195
rect 96 194 97 195
rect 95 194 96 195
rect 94 194 95 195
rect 93 194 94 195
rect 92 194 93 195
rect 91 194 92 195
rect 90 194 91 195
rect 89 194 90 195
rect 88 194 89 195
rect 87 194 88 195
rect 86 194 87 195
rect 85 194 86 195
rect 84 194 85 195
rect 83 194 84 195
rect 82 194 83 195
rect 81 194 82 195
rect 80 194 81 195
rect 79 194 80 195
rect 78 194 79 195
rect 77 194 78 195
rect 76 194 77 195
rect 75 194 76 195
rect 74 194 75 195
rect 73 194 74 195
rect 72 194 73 195
rect 71 194 72 195
rect 70 194 71 195
rect 51 194 52 195
rect 50 194 51 195
rect 49 194 50 195
rect 48 194 49 195
rect 47 194 48 195
rect 46 194 47 195
rect 31 194 32 195
rect 30 194 31 195
rect 29 194 30 195
rect 28 194 29 195
rect 27 194 28 195
rect 26 194 27 195
rect 25 194 26 195
rect 24 194 25 195
rect 23 194 24 195
rect 22 194 23 195
rect 21 194 22 195
rect 20 194 21 195
rect 19 194 20 195
rect 18 194 19 195
rect 17 194 18 195
rect 16 194 17 195
rect 15 194 16 195
rect 14 194 15 195
rect 13 194 14 195
rect 12 194 13 195
rect 480 195 481 196
rect 479 195 480 196
rect 478 195 479 196
rect 477 195 478 196
rect 476 195 477 196
rect 475 195 476 196
rect 474 195 475 196
rect 473 195 474 196
rect 472 195 473 196
rect 471 195 472 196
rect 470 195 471 196
rect 469 195 470 196
rect 468 195 469 196
rect 467 195 468 196
rect 466 195 467 196
rect 465 195 466 196
rect 464 195 465 196
rect 463 195 464 196
rect 462 195 463 196
rect 461 195 462 196
rect 460 195 461 196
rect 440 195 441 196
rect 439 195 440 196
rect 438 195 439 196
rect 437 195 438 196
rect 436 195 437 196
rect 435 195 436 196
rect 434 195 435 196
rect 433 195 434 196
rect 432 195 433 196
rect 431 195 432 196
rect 430 195 431 196
rect 429 195 430 196
rect 428 195 429 196
rect 427 195 428 196
rect 426 195 427 196
rect 425 195 426 196
rect 424 195 425 196
rect 423 195 424 196
rect 422 195 423 196
rect 421 195 422 196
rect 420 195 421 196
rect 419 195 420 196
rect 418 195 419 196
rect 417 195 418 196
rect 416 195 417 196
rect 415 195 416 196
rect 414 195 415 196
rect 413 195 414 196
rect 412 195 413 196
rect 411 195 412 196
rect 410 195 411 196
rect 409 195 410 196
rect 408 195 409 196
rect 407 195 408 196
rect 406 195 407 196
rect 405 195 406 196
rect 404 195 405 196
rect 403 195 404 196
rect 402 195 403 196
rect 401 195 402 196
rect 400 195 401 196
rect 399 195 400 196
rect 398 195 399 196
rect 397 195 398 196
rect 396 195 397 196
rect 395 195 396 196
rect 344 195 345 196
rect 343 195 344 196
rect 342 195 343 196
rect 341 195 342 196
rect 340 195 341 196
rect 339 195 340 196
rect 338 195 339 196
rect 337 195 338 196
rect 336 195 337 196
rect 335 195 336 196
rect 334 195 335 196
rect 333 195 334 196
rect 332 195 333 196
rect 331 195 332 196
rect 330 195 331 196
rect 329 195 330 196
rect 328 195 329 196
rect 327 195 328 196
rect 326 195 327 196
rect 325 195 326 196
rect 324 195 325 196
rect 323 195 324 196
rect 322 195 323 196
rect 321 195 322 196
rect 320 195 321 196
rect 319 195 320 196
rect 318 195 319 196
rect 317 195 318 196
rect 316 195 317 196
rect 315 195 316 196
rect 314 195 315 196
rect 313 195 314 196
rect 312 195 313 196
rect 311 195 312 196
rect 310 195 311 196
rect 309 195 310 196
rect 308 195 309 196
rect 307 195 308 196
rect 306 195 307 196
rect 305 195 306 196
rect 304 195 305 196
rect 303 195 304 196
rect 302 195 303 196
rect 301 195 302 196
rect 300 195 301 196
rect 299 195 300 196
rect 298 195 299 196
rect 297 195 298 196
rect 296 195 297 196
rect 295 195 296 196
rect 294 195 295 196
rect 293 195 294 196
rect 292 195 293 196
rect 291 195 292 196
rect 290 195 291 196
rect 289 195 290 196
rect 288 195 289 196
rect 287 195 288 196
rect 286 195 287 196
rect 285 195 286 196
rect 284 195 285 196
rect 283 195 284 196
rect 282 195 283 196
rect 281 195 282 196
rect 280 195 281 196
rect 279 195 280 196
rect 278 195 279 196
rect 277 195 278 196
rect 276 195 277 196
rect 275 195 276 196
rect 274 195 275 196
rect 273 195 274 196
rect 272 195 273 196
rect 271 195 272 196
rect 270 195 271 196
rect 269 195 270 196
rect 268 195 269 196
rect 253 195 254 196
rect 252 195 253 196
rect 251 195 252 196
rect 250 195 251 196
rect 249 195 250 196
rect 248 195 249 196
rect 247 195 248 196
rect 246 195 247 196
rect 245 195 246 196
rect 244 195 245 196
rect 243 195 244 196
rect 242 195 243 196
rect 241 195 242 196
rect 240 195 241 196
rect 239 195 240 196
rect 238 195 239 196
rect 237 195 238 196
rect 236 195 237 196
rect 235 195 236 196
rect 234 195 235 196
rect 233 195 234 196
rect 232 195 233 196
rect 231 195 232 196
rect 230 195 231 196
rect 229 195 230 196
rect 228 195 229 196
rect 227 195 228 196
rect 226 195 227 196
rect 225 195 226 196
rect 224 195 225 196
rect 223 195 224 196
rect 222 195 223 196
rect 221 195 222 196
rect 220 195 221 196
rect 219 195 220 196
rect 218 195 219 196
rect 217 195 218 196
rect 216 195 217 196
rect 215 195 216 196
rect 214 195 215 196
rect 213 195 214 196
rect 188 195 189 196
rect 187 195 188 196
rect 186 195 187 196
rect 185 195 186 196
rect 184 195 185 196
rect 183 195 184 196
rect 182 195 183 196
rect 181 195 182 196
rect 180 195 181 196
rect 179 195 180 196
rect 178 195 179 196
rect 177 195 178 196
rect 176 195 177 196
rect 175 195 176 196
rect 174 195 175 196
rect 173 195 174 196
rect 172 195 173 196
rect 171 195 172 196
rect 170 195 171 196
rect 169 195 170 196
rect 168 195 169 196
rect 167 195 168 196
rect 166 195 167 196
rect 165 195 166 196
rect 164 195 165 196
rect 163 195 164 196
rect 162 195 163 196
rect 161 195 162 196
rect 160 195 161 196
rect 159 195 160 196
rect 158 195 159 196
rect 157 195 158 196
rect 156 195 157 196
rect 155 195 156 196
rect 154 195 155 196
rect 153 195 154 196
rect 152 195 153 196
rect 151 195 152 196
rect 150 195 151 196
rect 149 195 150 196
rect 148 195 149 196
rect 147 195 148 196
rect 146 195 147 196
rect 145 195 146 196
rect 144 195 145 196
rect 143 195 144 196
rect 142 195 143 196
rect 141 195 142 196
rect 140 195 141 196
rect 139 195 140 196
rect 138 195 139 196
rect 137 195 138 196
rect 136 195 137 196
rect 135 195 136 196
rect 134 195 135 196
rect 133 195 134 196
rect 132 195 133 196
rect 131 195 132 196
rect 130 195 131 196
rect 129 195 130 196
rect 128 195 129 196
rect 127 195 128 196
rect 126 195 127 196
rect 125 195 126 196
rect 124 195 125 196
rect 123 195 124 196
rect 122 195 123 196
rect 121 195 122 196
rect 120 195 121 196
rect 119 195 120 196
rect 118 195 119 196
rect 117 195 118 196
rect 116 195 117 196
rect 115 195 116 196
rect 114 195 115 196
rect 113 195 114 196
rect 112 195 113 196
rect 111 195 112 196
rect 110 195 111 196
rect 109 195 110 196
rect 108 195 109 196
rect 107 195 108 196
rect 106 195 107 196
rect 105 195 106 196
rect 104 195 105 196
rect 103 195 104 196
rect 102 195 103 196
rect 101 195 102 196
rect 100 195 101 196
rect 99 195 100 196
rect 98 195 99 196
rect 97 195 98 196
rect 96 195 97 196
rect 95 195 96 196
rect 94 195 95 196
rect 93 195 94 196
rect 92 195 93 196
rect 91 195 92 196
rect 90 195 91 196
rect 89 195 90 196
rect 88 195 89 196
rect 87 195 88 196
rect 86 195 87 196
rect 85 195 86 196
rect 84 195 85 196
rect 83 195 84 196
rect 82 195 83 196
rect 81 195 82 196
rect 80 195 81 196
rect 79 195 80 196
rect 78 195 79 196
rect 77 195 78 196
rect 76 195 77 196
rect 75 195 76 196
rect 74 195 75 196
rect 73 195 74 196
rect 72 195 73 196
rect 71 195 72 196
rect 70 195 71 196
rect 51 195 52 196
rect 50 195 51 196
rect 49 195 50 196
rect 48 195 49 196
rect 47 195 48 196
rect 46 195 47 196
rect 45 195 46 196
rect 44 195 45 196
rect 32 195 33 196
rect 31 195 32 196
rect 30 195 31 196
rect 29 195 30 196
rect 28 195 29 196
rect 27 195 28 196
rect 26 195 27 196
rect 25 195 26 196
rect 24 195 25 196
rect 23 195 24 196
rect 22 195 23 196
rect 21 195 22 196
rect 20 195 21 196
rect 19 195 20 196
rect 18 195 19 196
rect 17 195 18 196
rect 16 195 17 196
rect 15 195 16 196
rect 14 195 15 196
rect 13 195 14 196
rect 12 195 13 196
rect 480 196 481 197
rect 479 196 480 197
rect 478 196 479 197
rect 477 196 478 197
rect 476 196 477 197
rect 475 196 476 197
rect 474 196 475 197
rect 473 196 474 197
rect 472 196 473 197
rect 471 196 472 197
rect 470 196 471 197
rect 469 196 470 197
rect 468 196 469 197
rect 467 196 468 197
rect 466 196 467 197
rect 465 196 466 197
rect 464 196 465 197
rect 463 196 464 197
rect 462 196 463 197
rect 461 196 462 197
rect 460 196 461 197
rect 440 196 441 197
rect 439 196 440 197
rect 438 196 439 197
rect 437 196 438 197
rect 436 196 437 197
rect 435 196 436 197
rect 434 196 435 197
rect 433 196 434 197
rect 432 196 433 197
rect 431 196 432 197
rect 430 196 431 197
rect 429 196 430 197
rect 428 196 429 197
rect 427 196 428 197
rect 426 196 427 197
rect 425 196 426 197
rect 424 196 425 197
rect 423 196 424 197
rect 422 196 423 197
rect 421 196 422 197
rect 420 196 421 197
rect 419 196 420 197
rect 418 196 419 197
rect 417 196 418 197
rect 416 196 417 197
rect 415 196 416 197
rect 414 196 415 197
rect 413 196 414 197
rect 412 196 413 197
rect 411 196 412 197
rect 410 196 411 197
rect 409 196 410 197
rect 408 196 409 197
rect 407 196 408 197
rect 406 196 407 197
rect 405 196 406 197
rect 404 196 405 197
rect 403 196 404 197
rect 402 196 403 197
rect 401 196 402 197
rect 400 196 401 197
rect 399 196 400 197
rect 398 196 399 197
rect 397 196 398 197
rect 396 196 397 197
rect 395 196 396 197
rect 345 196 346 197
rect 344 196 345 197
rect 343 196 344 197
rect 342 196 343 197
rect 341 196 342 197
rect 340 196 341 197
rect 339 196 340 197
rect 338 196 339 197
rect 337 196 338 197
rect 336 196 337 197
rect 335 196 336 197
rect 334 196 335 197
rect 333 196 334 197
rect 332 196 333 197
rect 331 196 332 197
rect 330 196 331 197
rect 329 196 330 197
rect 328 196 329 197
rect 327 196 328 197
rect 326 196 327 197
rect 325 196 326 197
rect 324 196 325 197
rect 323 196 324 197
rect 322 196 323 197
rect 321 196 322 197
rect 320 196 321 197
rect 319 196 320 197
rect 318 196 319 197
rect 317 196 318 197
rect 316 196 317 197
rect 315 196 316 197
rect 314 196 315 197
rect 313 196 314 197
rect 312 196 313 197
rect 311 196 312 197
rect 310 196 311 197
rect 309 196 310 197
rect 308 196 309 197
rect 307 196 308 197
rect 306 196 307 197
rect 305 196 306 197
rect 304 196 305 197
rect 303 196 304 197
rect 302 196 303 197
rect 301 196 302 197
rect 300 196 301 197
rect 299 196 300 197
rect 298 196 299 197
rect 297 196 298 197
rect 296 196 297 197
rect 295 196 296 197
rect 294 196 295 197
rect 293 196 294 197
rect 292 196 293 197
rect 291 196 292 197
rect 290 196 291 197
rect 289 196 290 197
rect 288 196 289 197
rect 287 196 288 197
rect 286 196 287 197
rect 285 196 286 197
rect 284 196 285 197
rect 283 196 284 197
rect 282 196 283 197
rect 281 196 282 197
rect 280 196 281 197
rect 279 196 280 197
rect 278 196 279 197
rect 277 196 278 197
rect 276 196 277 197
rect 275 196 276 197
rect 274 196 275 197
rect 273 196 274 197
rect 272 196 273 197
rect 271 196 272 197
rect 270 196 271 197
rect 269 196 270 197
rect 268 196 269 197
rect 267 196 268 197
rect 252 196 253 197
rect 251 196 252 197
rect 250 196 251 197
rect 249 196 250 197
rect 248 196 249 197
rect 247 196 248 197
rect 246 196 247 197
rect 245 196 246 197
rect 244 196 245 197
rect 243 196 244 197
rect 242 196 243 197
rect 241 196 242 197
rect 240 196 241 197
rect 239 196 240 197
rect 238 196 239 197
rect 237 196 238 197
rect 236 196 237 197
rect 235 196 236 197
rect 234 196 235 197
rect 233 196 234 197
rect 232 196 233 197
rect 231 196 232 197
rect 230 196 231 197
rect 229 196 230 197
rect 228 196 229 197
rect 227 196 228 197
rect 226 196 227 197
rect 225 196 226 197
rect 224 196 225 197
rect 223 196 224 197
rect 222 196 223 197
rect 221 196 222 197
rect 220 196 221 197
rect 219 196 220 197
rect 218 196 219 197
rect 217 196 218 197
rect 216 196 217 197
rect 215 196 216 197
rect 214 196 215 197
rect 213 196 214 197
rect 212 196 213 197
rect 187 196 188 197
rect 186 196 187 197
rect 185 196 186 197
rect 184 196 185 197
rect 183 196 184 197
rect 182 196 183 197
rect 181 196 182 197
rect 180 196 181 197
rect 179 196 180 197
rect 178 196 179 197
rect 177 196 178 197
rect 176 196 177 197
rect 175 196 176 197
rect 174 196 175 197
rect 173 196 174 197
rect 172 196 173 197
rect 171 196 172 197
rect 170 196 171 197
rect 169 196 170 197
rect 168 196 169 197
rect 167 196 168 197
rect 166 196 167 197
rect 165 196 166 197
rect 164 196 165 197
rect 163 196 164 197
rect 162 196 163 197
rect 161 196 162 197
rect 160 196 161 197
rect 159 196 160 197
rect 158 196 159 197
rect 157 196 158 197
rect 156 196 157 197
rect 155 196 156 197
rect 154 196 155 197
rect 153 196 154 197
rect 152 196 153 197
rect 151 196 152 197
rect 150 196 151 197
rect 149 196 150 197
rect 148 196 149 197
rect 147 196 148 197
rect 146 196 147 197
rect 145 196 146 197
rect 144 196 145 197
rect 143 196 144 197
rect 142 196 143 197
rect 141 196 142 197
rect 140 196 141 197
rect 139 196 140 197
rect 138 196 139 197
rect 137 196 138 197
rect 136 196 137 197
rect 135 196 136 197
rect 134 196 135 197
rect 133 196 134 197
rect 132 196 133 197
rect 131 196 132 197
rect 130 196 131 197
rect 129 196 130 197
rect 128 196 129 197
rect 127 196 128 197
rect 126 196 127 197
rect 125 196 126 197
rect 124 196 125 197
rect 123 196 124 197
rect 122 196 123 197
rect 121 196 122 197
rect 120 196 121 197
rect 119 196 120 197
rect 118 196 119 197
rect 117 196 118 197
rect 116 196 117 197
rect 115 196 116 197
rect 114 196 115 197
rect 113 196 114 197
rect 112 196 113 197
rect 111 196 112 197
rect 110 196 111 197
rect 109 196 110 197
rect 108 196 109 197
rect 107 196 108 197
rect 106 196 107 197
rect 105 196 106 197
rect 104 196 105 197
rect 103 196 104 197
rect 102 196 103 197
rect 101 196 102 197
rect 100 196 101 197
rect 99 196 100 197
rect 98 196 99 197
rect 97 196 98 197
rect 96 196 97 197
rect 95 196 96 197
rect 94 196 95 197
rect 93 196 94 197
rect 92 196 93 197
rect 91 196 92 197
rect 90 196 91 197
rect 89 196 90 197
rect 88 196 89 197
rect 87 196 88 197
rect 86 196 87 197
rect 85 196 86 197
rect 84 196 85 197
rect 83 196 84 197
rect 82 196 83 197
rect 81 196 82 197
rect 80 196 81 197
rect 79 196 80 197
rect 78 196 79 197
rect 77 196 78 197
rect 76 196 77 197
rect 75 196 76 197
rect 74 196 75 197
rect 73 196 74 197
rect 72 196 73 197
rect 71 196 72 197
rect 70 196 71 197
rect 52 196 53 197
rect 51 196 52 197
rect 50 196 51 197
rect 49 196 50 197
rect 48 196 49 197
rect 47 196 48 197
rect 46 196 47 197
rect 45 196 46 197
rect 44 196 45 197
rect 43 196 44 197
rect 42 196 43 197
rect 41 196 42 197
rect 40 196 41 197
rect 35 196 36 197
rect 34 196 35 197
rect 33 196 34 197
rect 32 196 33 197
rect 31 196 32 197
rect 30 196 31 197
rect 29 196 30 197
rect 28 196 29 197
rect 27 196 28 197
rect 26 196 27 197
rect 25 196 26 197
rect 24 196 25 197
rect 23 196 24 197
rect 22 196 23 197
rect 21 196 22 197
rect 20 196 21 197
rect 19 196 20 197
rect 18 196 19 197
rect 17 196 18 197
rect 16 196 17 197
rect 15 196 16 197
rect 14 196 15 197
rect 13 196 14 197
rect 12 196 13 197
rect 480 197 481 198
rect 479 197 480 198
rect 478 197 479 198
rect 477 197 478 198
rect 476 197 477 198
rect 475 197 476 198
rect 474 197 475 198
rect 473 197 474 198
rect 472 197 473 198
rect 471 197 472 198
rect 470 197 471 198
rect 469 197 470 198
rect 468 197 469 198
rect 467 197 468 198
rect 466 197 467 198
rect 465 197 466 198
rect 464 197 465 198
rect 463 197 464 198
rect 462 197 463 198
rect 461 197 462 198
rect 460 197 461 198
rect 405 197 406 198
rect 404 197 405 198
rect 403 197 404 198
rect 402 197 403 198
rect 401 197 402 198
rect 400 197 401 198
rect 399 197 400 198
rect 398 197 399 198
rect 397 197 398 198
rect 396 197 397 198
rect 395 197 396 198
rect 346 197 347 198
rect 345 197 346 198
rect 344 197 345 198
rect 343 197 344 198
rect 342 197 343 198
rect 341 197 342 198
rect 340 197 341 198
rect 339 197 340 198
rect 338 197 339 198
rect 337 197 338 198
rect 336 197 337 198
rect 335 197 336 198
rect 334 197 335 198
rect 333 197 334 198
rect 332 197 333 198
rect 331 197 332 198
rect 330 197 331 198
rect 329 197 330 198
rect 328 197 329 198
rect 327 197 328 198
rect 326 197 327 198
rect 325 197 326 198
rect 324 197 325 198
rect 323 197 324 198
rect 322 197 323 198
rect 321 197 322 198
rect 320 197 321 198
rect 319 197 320 198
rect 318 197 319 198
rect 317 197 318 198
rect 316 197 317 198
rect 315 197 316 198
rect 314 197 315 198
rect 313 197 314 198
rect 312 197 313 198
rect 311 197 312 198
rect 310 197 311 198
rect 309 197 310 198
rect 308 197 309 198
rect 307 197 308 198
rect 306 197 307 198
rect 305 197 306 198
rect 304 197 305 198
rect 303 197 304 198
rect 302 197 303 198
rect 301 197 302 198
rect 300 197 301 198
rect 299 197 300 198
rect 298 197 299 198
rect 297 197 298 198
rect 296 197 297 198
rect 295 197 296 198
rect 294 197 295 198
rect 293 197 294 198
rect 292 197 293 198
rect 291 197 292 198
rect 290 197 291 198
rect 289 197 290 198
rect 288 197 289 198
rect 287 197 288 198
rect 286 197 287 198
rect 285 197 286 198
rect 284 197 285 198
rect 283 197 284 198
rect 282 197 283 198
rect 281 197 282 198
rect 280 197 281 198
rect 279 197 280 198
rect 278 197 279 198
rect 277 197 278 198
rect 276 197 277 198
rect 275 197 276 198
rect 274 197 275 198
rect 273 197 274 198
rect 272 197 273 198
rect 271 197 272 198
rect 270 197 271 198
rect 269 197 270 198
rect 268 197 269 198
rect 267 197 268 198
rect 266 197 267 198
rect 265 197 266 198
rect 252 197 253 198
rect 251 197 252 198
rect 250 197 251 198
rect 249 197 250 198
rect 248 197 249 198
rect 247 197 248 198
rect 246 197 247 198
rect 245 197 246 198
rect 244 197 245 198
rect 243 197 244 198
rect 242 197 243 198
rect 241 197 242 198
rect 240 197 241 198
rect 239 197 240 198
rect 238 197 239 198
rect 237 197 238 198
rect 236 197 237 198
rect 235 197 236 198
rect 234 197 235 198
rect 233 197 234 198
rect 232 197 233 198
rect 231 197 232 198
rect 230 197 231 198
rect 229 197 230 198
rect 228 197 229 198
rect 227 197 228 198
rect 226 197 227 198
rect 225 197 226 198
rect 224 197 225 198
rect 223 197 224 198
rect 222 197 223 198
rect 221 197 222 198
rect 220 197 221 198
rect 219 197 220 198
rect 218 197 219 198
rect 217 197 218 198
rect 216 197 217 198
rect 215 197 216 198
rect 214 197 215 198
rect 213 197 214 198
rect 212 197 213 198
rect 211 197 212 198
rect 185 197 186 198
rect 184 197 185 198
rect 183 197 184 198
rect 182 197 183 198
rect 181 197 182 198
rect 180 197 181 198
rect 179 197 180 198
rect 178 197 179 198
rect 177 197 178 198
rect 176 197 177 198
rect 175 197 176 198
rect 174 197 175 198
rect 173 197 174 198
rect 172 197 173 198
rect 171 197 172 198
rect 170 197 171 198
rect 169 197 170 198
rect 168 197 169 198
rect 167 197 168 198
rect 166 197 167 198
rect 165 197 166 198
rect 164 197 165 198
rect 163 197 164 198
rect 162 197 163 198
rect 161 197 162 198
rect 160 197 161 198
rect 159 197 160 198
rect 158 197 159 198
rect 157 197 158 198
rect 156 197 157 198
rect 155 197 156 198
rect 154 197 155 198
rect 153 197 154 198
rect 152 197 153 198
rect 151 197 152 198
rect 150 197 151 198
rect 149 197 150 198
rect 148 197 149 198
rect 147 197 148 198
rect 146 197 147 198
rect 145 197 146 198
rect 144 197 145 198
rect 143 197 144 198
rect 142 197 143 198
rect 141 197 142 198
rect 140 197 141 198
rect 139 197 140 198
rect 138 197 139 198
rect 137 197 138 198
rect 136 197 137 198
rect 135 197 136 198
rect 134 197 135 198
rect 133 197 134 198
rect 132 197 133 198
rect 131 197 132 198
rect 130 197 131 198
rect 129 197 130 198
rect 128 197 129 198
rect 127 197 128 198
rect 126 197 127 198
rect 125 197 126 198
rect 124 197 125 198
rect 123 197 124 198
rect 122 197 123 198
rect 121 197 122 198
rect 120 197 121 198
rect 119 197 120 198
rect 118 197 119 198
rect 117 197 118 198
rect 116 197 117 198
rect 115 197 116 198
rect 114 197 115 198
rect 113 197 114 198
rect 112 197 113 198
rect 111 197 112 198
rect 110 197 111 198
rect 109 197 110 198
rect 108 197 109 198
rect 107 197 108 198
rect 106 197 107 198
rect 105 197 106 198
rect 104 197 105 198
rect 103 197 104 198
rect 102 197 103 198
rect 101 197 102 198
rect 100 197 101 198
rect 99 197 100 198
rect 98 197 99 198
rect 97 197 98 198
rect 96 197 97 198
rect 95 197 96 198
rect 94 197 95 198
rect 93 197 94 198
rect 92 197 93 198
rect 91 197 92 198
rect 90 197 91 198
rect 89 197 90 198
rect 88 197 89 198
rect 87 197 88 198
rect 86 197 87 198
rect 85 197 86 198
rect 84 197 85 198
rect 83 197 84 198
rect 82 197 83 198
rect 81 197 82 198
rect 80 197 81 198
rect 79 197 80 198
rect 78 197 79 198
rect 77 197 78 198
rect 76 197 77 198
rect 75 197 76 198
rect 74 197 75 198
rect 73 197 74 198
rect 72 197 73 198
rect 71 197 72 198
rect 70 197 71 198
rect 52 197 53 198
rect 51 197 52 198
rect 50 197 51 198
rect 49 197 50 198
rect 48 197 49 198
rect 47 197 48 198
rect 46 197 47 198
rect 45 197 46 198
rect 44 197 45 198
rect 43 197 44 198
rect 42 197 43 198
rect 41 197 42 198
rect 40 197 41 198
rect 39 197 40 198
rect 38 197 39 198
rect 37 197 38 198
rect 36 197 37 198
rect 35 197 36 198
rect 34 197 35 198
rect 33 197 34 198
rect 32 197 33 198
rect 31 197 32 198
rect 30 197 31 198
rect 29 197 30 198
rect 28 197 29 198
rect 27 197 28 198
rect 26 197 27 198
rect 25 197 26 198
rect 24 197 25 198
rect 23 197 24 198
rect 22 197 23 198
rect 21 197 22 198
rect 20 197 21 198
rect 19 197 20 198
rect 18 197 19 198
rect 17 197 18 198
rect 16 197 17 198
rect 15 197 16 198
rect 14 197 15 198
rect 13 197 14 198
rect 12 197 13 198
rect 480 198 481 199
rect 479 198 480 199
rect 470 198 471 199
rect 469 198 470 199
rect 460 198 461 199
rect 399 198 400 199
rect 398 198 399 199
rect 397 198 398 199
rect 396 198 397 199
rect 395 198 396 199
rect 347 198 348 199
rect 346 198 347 199
rect 345 198 346 199
rect 344 198 345 199
rect 343 198 344 199
rect 342 198 343 199
rect 341 198 342 199
rect 340 198 341 199
rect 339 198 340 199
rect 338 198 339 199
rect 337 198 338 199
rect 336 198 337 199
rect 335 198 336 199
rect 334 198 335 199
rect 333 198 334 199
rect 332 198 333 199
rect 331 198 332 199
rect 330 198 331 199
rect 329 198 330 199
rect 328 198 329 199
rect 327 198 328 199
rect 326 198 327 199
rect 325 198 326 199
rect 324 198 325 199
rect 323 198 324 199
rect 322 198 323 199
rect 321 198 322 199
rect 320 198 321 199
rect 319 198 320 199
rect 318 198 319 199
rect 317 198 318 199
rect 316 198 317 199
rect 315 198 316 199
rect 314 198 315 199
rect 313 198 314 199
rect 312 198 313 199
rect 311 198 312 199
rect 310 198 311 199
rect 309 198 310 199
rect 308 198 309 199
rect 307 198 308 199
rect 306 198 307 199
rect 305 198 306 199
rect 304 198 305 199
rect 303 198 304 199
rect 302 198 303 199
rect 301 198 302 199
rect 300 198 301 199
rect 299 198 300 199
rect 298 198 299 199
rect 297 198 298 199
rect 296 198 297 199
rect 295 198 296 199
rect 294 198 295 199
rect 293 198 294 199
rect 292 198 293 199
rect 291 198 292 199
rect 290 198 291 199
rect 289 198 290 199
rect 288 198 289 199
rect 287 198 288 199
rect 286 198 287 199
rect 285 198 286 199
rect 284 198 285 199
rect 283 198 284 199
rect 282 198 283 199
rect 281 198 282 199
rect 280 198 281 199
rect 279 198 280 199
rect 278 198 279 199
rect 277 198 278 199
rect 276 198 277 199
rect 275 198 276 199
rect 274 198 275 199
rect 273 198 274 199
rect 272 198 273 199
rect 271 198 272 199
rect 270 198 271 199
rect 269 198 270 199
rect 268 198 269 199
rect 267 198 268 199
rect 266 198 267 199
rect 265 198 266 199
rect 264 198 265 199
rect 251 198 252 199
rect 250 198 251 199
rect 249 198 250 199
rect 248 198 249 199
rect 247 198 248 199
rect 246 198 247 199
rect 245 198 246 199
rect 244 198 245 199
rect 243 198 244 199
rect 242 198 243 199
rect 241 198 242 199
rect 240 198 241 199
rect 239 198 240 199
rect 238 198 239 199
rect 237 198 238 199
rect 236 198 237 199
rect 235 198 236 199
rect 234 198 235 199
rect 233 198 234 199
rect 232 198 233 199
rect 231 198 232 199
rect 230 198 231 199
rect 229 198 230 199
rect 228 198 229 199
rect 227 198 228 199
rect 226 198 227 199
rect 225 198 226 199
rect 224 198 225 199
rect 223 198 224 199
rect 222 198 223 199
rect 221 198 222 199
rect 220 198 221 199
rect 219 198 220 199
rect 218 198 219 199
rect 217 198 218 199
rect 216 198 217 199
rect 215 198 216 199
rect 214 198 215 199
rect 213 198 214 199
rect 212 198 213 199
rect 211 198 212 199
rect 210 198 211 199
rect 184 198 185 199
rect 183 198 184 199
rect 182 198 183 199
rect 181 198 182 199
rect 180 198 181 199
rect 179 198 180 199
rect 178 198 179 199
rect 177 198 178 199
rect 176 198 177 199
rect 175 198 176 199
rect 174 198 175 199
rect 173 198 174 199
rect 172 198 173 199
rect 171 198 172 199
rect 170 198 171 199
rect 169 198 170 199
rect 168 198 169 199
rect 167 198 168 199
rect 166 198 167 199
rect 165 198 166 199
rect 164 198 165 199
rect 163 198 164 199
rect 162 198 163 199
rect 161 198 162 199
rect 160 198 161 199
rect 159 198 160 199
rect 158 198 159 199
rect 157 198 158 199
rect 156 198 157 199
rect 155 198 156 199
rect 154 198 155 199
rect 153 198 154 199
rect 152 198 153 199
rect 151 198 152 199
rect 150 198 151 199
rect 149 198 150 199
rect 148 198 149 199
rect 147 198 148 199
rect 146 198 147 199
rect 145 198 146 199
rect 144 198 145 199
rect 143 198 144 199
rect 142 198 143 199
rect 141 198 142 199
rect 140 198 141 199
rect 139 198 140 199
rect 138 198 139 199
rect 137 198 138 199
rect 136 198 137 199
rect 135 198 136 199
rect 134 198 135 199
rect 133 198 134 199
rect 132 198 133 199
rect 131 198 132 199
rect 130 198 131 199
rect 129 198 130 199
rect 128 198 129 199
rect 127 198 128 199
rect 126 198 127 199
rect 125 198 126 199
rect 124 198 125 199
rect 123 198 124 199
rect 122 198 123 199
rect 121 198 122 199
rect 120 198 121 199
rect 119 198 120 199
rect 118 198 119 199
rect 117 198 118 199
rect 116 198 117 199
rect 115 198 116 199
rect 114 198 115 199
rect 113 198 114 199
rect 112 198 113 199
rect 111 198 112 199
rect 110 198 111 199
rect 109 198 110 199
rect 108 198 109 199
rect 107 198 108 199
rect 106 198 107 199
rect 105 198 106 199
rect 104 198 105 199
rect 103 198 104 199
rect 102 198 103 199
rect 101 198 102 199
rect 100 198 101 199
rect 99 198 100 199
rect 98 198 99 199
rect 97 198 98 199
rect 96 198 97 199
rect 95 198 96 199
rect 94 198 95 199
rect 93 198 94 199
rect 92 198 93 199
rect 91 198 92 199
rect 90 198 91 199
rect 89 198 90 199
rect 88 198 89 199
rect 87 198 88 199
rect 86 198 87 199
rect 85 198 86 199
rect 84 198 85 199
rect 83 198 84 199
rect 82 198 83 199
rect 81 198 82 199
rect 80 198 81 199
rect 79 198 80 199
rect 78 198 79 199
rect 77 198 78 199
rect 76 198 77 199
rect 75 198 76 199
rect 74 198 75 199
rect 73 198 74 199
rect 72 198 73 199
rect 71 198 72 199
rect 53 198 54 199
rect 52 198 53 199
rect 51 198 52 199
rect 50 198 51 199
rect 49 198 50 199
rect 48 198 49 199
rect 47 198 48 199
rect 46 198 47 199
rect 45 198 46 199
rect 44 198 45 199
rect 43 198 44 199
rect 42 198 43 199
rect 41 198 42 199
rect 40 198 41 199
rect 39 198 40 199
rect 38 198 39 199
rect 37 198 38 199
rect 36 198 37 199
rect 35 198 36 199
rect 34 198 35 199
rect 33 198 34 199
rect 32 198 33 199
rect 31 198 32 199
rect 30 198 31 199
rect 29 198 30 199
rect 28 198 29 199
rect 27 198 28 199
rect 26 198 27 199
rect 25 198 26 199
rect 24 198 25 199
rect 23 198 24 199
rect 22 198 23 199
rect 21 198 22 199
rect 20 198 21 199
rect 19 198 20 199
rect 18 198 19 199
rect 17 198 18 199
rect 16 198 17 199
rect 15 198 16 199
rect 14 198 15 199
rect 13 198 14 199
rect 12 198 13 199
rect 11 198 12 199
rect 480 199 481 200
rect 470 199 471 200
rect 469 199 470 200
rect 460 199 461 200
rect 398 199 399 200
rect 397 199 398 200
rect 396 199 397 200
rect 395 199 396 200
rect 348 199 349 200
rect 347 199 348 200
rect 346 199 347 200
rect 345 199 346 200
rect 344 199 345 200
rect 343 199 344 200
rect 342 199 343 200
rect 341 199 342 200
rect 340 199 341 200
rect 339 199 340 200
rect 338 199 339 200
rect 337 199 338 200
rect 336 199 337 200
rect 335 199 336 200
rect 334 199 335 200
rect 333 199 334 200
rect 332 199 333 200
rect 331 199 332 200
rect 330 199 331 200
rect 329 199 330 200
rect 328 199 329 200
rect 327 199 328 200
rect 326 199 327 200
rect 325 199 326 200
rect 324 199 325 200
rect 323 199 324 200
rect 322 199 323 200
rect 321 199 322 200
rect 320 199 321 200
rect 319 199 320 200
rect 318 199 319 200
rect 317 199 318 200
rect 316 199 317 200
rect 315 199 316 200
rect 314 199 315 200
rect 313 199 314 200
rect 312 199 313 200
rect 311 199 312 200
rect 310 199 311 200
rect 309 199 310 200
rect 308 199 309 200
rect 307 199 308 200
rect 306 199 307 200
rect 305 199 306 200
rect 304 199 305 200
rect 303 199 304 200
rect 302 199 303 200
rect 301 199 302 200
rect 300 199 301 200
rect 299 199 300 200
rect 298 199 299 200
rect 297 199 298 200
rect 296 199 297 200
rect 295 199 296 200
rect 294 199 295 200
rect 293 199 294 200
rect 292 199 293 200
rect 291 199 292 200
rect 290 199 291 200
rect 289 199 290 200
rect 288 199 289 200
rect 287 199 288 200
rect 286 199 287 200
rect 285 199 286 200
rect 284 199 285 200
rect 283 199 284 200
rect 282 199 283 200
rect 281 199 282 200
rect 280 199 281 200
rect 279 199 280 200
rect 278 199 279 200
rect 277 199 278 200
rect 276 199 277 200
rect 275 199 276 200
rect 274 199 275 200
rect 273 199 274 200
rect 272 199 273 200
rect 271 199 272 200
rect 270 199 271 200
rect 269 199 270 200
rect 268 199 269 200
rect 267 199 268 200
rect 266 199 267 200
rect 265 199 266 200
rect 264 199 265 200
rect 263 199 264 200
rect 250 199 251 200
rect 249 199 250 200
rect 248 199 249 200
rect 247 199 248 200
rect 246 199 247 200
rect 245 199 246 200
rect 244 199 245 200
rect 243 199 244 200
rect 242 199 243 200
rect 241 199 242 200
rect 240 199 241 200
rect 239 199 240 200
rect 238 199 239 200
rect 237 199 238 200
rect 236 199 237 200
rect 235 199 236 200
rect 234 199 235 200
rect 233 199 234 200
rect 232 199 233 200
rect 231 199 232 200
rect 230 199 231 200
rect 229 199 230 200
rect 228 199 229 200
rect 227 199 228 200
rect 226 199 227 200
rect 225 199 226 200
rect 224 199 225 200
rect 223 199 224 200
rect 222 199 223 200
rect 221 199 222 200
rect 220 199 221 200
rect 219 199 220 200
rect 218 199 219 200
rect 217 199 218 200
rect 216 199 217 200
rect 215 199 216 200
rect 214 199 215 200
rect 213 199 214 200
rect 212 199 213 200
rect 211 199 212 200
rect 210 199 211 200
rect 183 199 184 200
rect 182 199 183 200
rect 181 199 182 200
rect 180 199 181 200
rect 179 199 180 200
rect 178 199 179 200
rect 177 199 178 200
rect 176 199 177 200
rect 175 199 176 200
rect 174 199 175 200
rect 173 199 174 200
rect 172 199 173 200
rect 171 199 172 200
rect 170 199 171 200
rect 169 199 170 200
rect 168 199 169 200
rect 167 199 168 200
rect 166 199 167 200
rect 165 199 166 200
rect 164 199 165 200
rect 163 199 164 200
rect 162 199 163 200
rect 161 199 162 200
rect 160 199 161 200
rect 159 199 160 200
rect 158 199 159 200
rect 157 199 158 200
rect 156 199 157 200
rect 155 199 156 200
rect 154 199 155 200
rect 153 199 154 200
rect 152 199 153 200
rect 151 199 152 200
rect 150 199 151 200
rect 149 199 150 200
rect 148 199 149 200
rect 147 199 148 200
rect 146 199 147 200
rect 145 199 146 200
rect 144 199 145 200
rect 143 199 144 200
rect 142 199 143 200
rect 141 199 142 200
rect 140 199 141 200
rect 139 199 140 200
rect 138 199 139 200
rect 137 199 138 200
rect 136 199 137 200
rect 135 199 136 200
rect 134 199 135 200
rect 133 199 134 200
rect 132 199 133 200
rect 131 199 132 200
rect 130 199 131 200
rect 129 199 130 200
rect 128 199 129 200
rect 127 199 128 200
rect 126 199 127 200
rect 125 199 126 200
rect 124 199 125 200
rect 123 199 124 200
rect 122 199 123 200
rect 121 199 122 200
rect 120 199 121 200
rect 119 199 120 200
rect 118 199 119 200
rect 117 199 118 200
rect 116 199 117 200
rect 115 199 116 200
rect 114 199 115 200
rect 113 199 114 200
rect 112 199 113 200
rect 111 199 112 200
rect 110 199 111 200
rect 109 199 110 200
rect 108 199 109 200
rect 107 199 108 200
rect 106 199 107 200
rect 105 199 106 200
rect 104 199 105 200
rect 103 199 104 200
rect 102 199 103 200
rect 101 199 102 200
rect 100 199 101 200
rect 99 199 100 200
rect 98 199 99 200
rect 97 199 98 200
rect 96 199 97 200
rect 95 199 96 200
rect 94 199 95 200
rect 93 199 94 200
rect 92 199 93 200
rect 91 199 92 200
rect 90 199 91 200
rect 89 199 90 200
rect 88 199 89 200
rect 87 199 88 200
rect 86 199 87 200
rect 85 199 86 200
rect 84 199 85 200
rect 83 199 84 200
rect 82 199 83 200
rect 81 199 82 200
rect 80 199 81 200
rect 79 199 80 200
rect 78 199 79 200
rect 77 199 78 200
rect 76 199 77 200
rect 75 199 76 200
rect 74 199 75 200
rect 73 199 74 200
rect 72 199 73 200
rect 71 199 72 200
rect 54 199 55 200
rect 53 199 54 200
rect 52 199 53 200
rect 51 199 52 200
rect 50 199 51 200
rect 49 199 50 200
rect 48 199 49 200
rect 47 199 48 200
rect 46 199 47 200
rect 45 199 46 200
rect 44 199 45 200
rect 43 199 44 200
rect 42 199 43 200
rect 41 199 42 200
rect 40 199 41 200
rect 39 199 40 200
rect 38 199 39 200
rect 37 199 38 200
rect 36 199 37 200
rect 35 199 36 200
rect 34 199 35 200
rect 33 199 34 200
rect 32 199 33 200
rect 31 199 32 200
rect 30 199 31 200
rect 29 199 30 200
rect 28 199 29 200
rect 27 199 28 200
rect 26 199 27 200
rect 25 199 26 200
rect 24 199 25 200
rect 23 199 24 200
rect 22 199 23 200
rect 21 199 22 200
rect 20 199 21 200
rect 19 199 20 200
rect 18 199 19 200
rect 17 199 18 200
rect 16 199 17 200
rect 15 199 16 200
rect 14 199 15 200
rect 13 199 14 200
rect 12 199 13 200
rect 11 199 12 200
rect 480 200 481 201
rect 470 200 471 201
rect 469 200 470 201
rect 460 200 461 201
rect 397 200 398 201
rect 396 200 397 201
rect 395 200 396 201
rect 349 200 350 201
rect 348 200 349 201
rect 347 200 348 201
rect 346 200 347 201
rect 345 200 346 201
rect 344 200 345 201
rect 343 200 344 201
rect 342 200 343 201
rect 341 200 342 201
rect 340 200 341 201
rect 339 200 340 201
rect 338 200 339 201
rect 337 200 338 201
rect 336 200 337 201
rect 335 200 336 201
rect 334 200 335 201
rect 333 200 334 201
rect 332 200 333 201
rect 331 200 332 201
rect 330 200 331 201
rect 329 200 330 201
rect 328 200 329 201
rect 327 200 328 201
rect 326 200 327 201
rect 325 200 326 201
rect 324 200 325 201
rect 323 200 324 201
rect 322 200 323 201
rect 321 200 322 201
rect 320 200 321 201
rect 319 200 320 201
rect 318 200 319 201
rect 317 200 318 201
rect 316 200 317 201
rect 315 200 316 201
rect 314 200 315 201
rect 313 200 314 201
rect 312 200 313 201
rect 311 200 312 201
rect 310 200 311 201
rect 309 200 310 201
rect 308 200 309 201
rect 307 200 308 201
rect 306 200 307 201
rect 305 200 306 201
rect 304 200 305 201
rect 303 200 304 201
rect 302 200 303 201
rect 301 200 302 201
rect 300 200 301 201
rect 299 200 300 201
rect 298 200 299 201
rect 297 200 298 201
rect 296 200 297 201
rect 295 200 296 201
rect 294 200 295 201
rect 293 200 294 201
rect 292 200 293 201
rect 291 200 292 201
rect 290 200 291 201
rect 289 200 290 201
rect 288 200 289 201
rect 287 200 288 201
rect 286 200 287 201
rect 285 200 286 201
rect 284 200 285 201
rect 283 200 284 201
rect 282 200 283 201
rect 281 200 282 201
rect 280 200 281 201
rect 279 200 280 201
rect 278 200 279 201
rect 277 200 278 201
rect 276 200 277 201
rect 275 200 276 201
rect 274 200 275 201
rect 273 200 274 201
rect 272 200 273 201
rect 271 200 272 201
rect 270 200 271 201
rect 269 200 270 201
rect 268 200 269 201
rect 267 200 268 201
rect 266 200 267 201
rect 265 200 266 201
rect 264 200 265 201
rect 263 200 264 201
rect 262 200 263 201
rect 261 200 262 201
rect 250 200 251 201
rect 249 200 250 201
rect 248 200 249 201
rect 247 200 248 201
rect 246 200 247 201
rect 245 200 246 201
rect 244 200 245 201
rect 243 200 244 201
rect 242 200 243 201
rect 241 200 242 201
rect 240 200 241 201
rect 239 200 240 201
rect 238 200 239 201
rect 237 200 238 201
rect 236 200 237 201
rect 235 200 236 201
rect 234 200 235 201
rect 233 200 234 201
rect 232 200 233 201
rect 231 200 232 201
rect 230 200 231 201
rect 229 200 230 201
rect 228 200 229 201
rect 227 200 228 201
rect 226 200 227 201
rect 225 200 226 201
rect 224 200 225 201
rect 223 200 224 201
rect 222 200 223 201
rect 221 200 222 201
rect 220 200 221 201
rect 219 200 220 201
rect 218 200 219 201
rect 217 200 218 201
rect 216 200 217 201
rect 215 200 216 201
rect 214 200 215 201
rect 213 200 214 201
rect 212 200 213 201
rect 211 200 212 201
rect 210 200 211 201
rect 209 200 210 201
rect 182 200 183 201
rect 181 200 182 201
rect 180 200 181 201
rect 179 200 180 201
rect 178 200 179 201
rect 177 200 178 201
rect 176 200 177 201
rect 175 200 176 201
rect 174 200 175 201
rect 173 200 174 201
rect 172 200 173 201
rect 171 200 172 201
rect 170 200 171 201
rect 169 200 170 201
rect 168 200 169 201
rect 167 200 168 201
rect 166 200 167 201
rect 165 200 166 201
rect 164 200 165 201
rect 163 200 164 201
rect 162 200 163 201
rect 161 200 162 201
rect 160 200 161 201
rect 159 200 160 201
rect 158 200 159 201
rect 157 200 158 201
rect 156 200 157 201
rect 155 200 156 201
rect 154 200 155 201
rect 153 200 154 201
rect 152 200 153 201
rect 151 200 152 201
rect 150 200 151 201
rect 149 200 150 201
rect 148 200 149 201
rect 147 200 148 201
rect 146 200 147 201
rect 145 200 146 201
rect 144 200 145 201
rect 143 200 144 201
rect 142 200 143 201
rect 141 200 142 201
rect 140 200 141 201
rect 139 200 140 201
rect 138 200 139 201
rect 137 200 138 201
rect 136 200 137 201
rect 135 200 136 201
rect 134 200 135 201
rect 133 200 134 201
rect 132 200 133 201
rect 131 200 132 201
rect 130 200 131 201
rect 129 200 130 201
rect 128 200 129 201
rect 127 200 128 201
rect 126 200 127 201
rect 125 200 126 201
rect 124 200 125 201
rect 123 200 124 201
rect 122 200 123 201
rect 121 200 122 201
rect 120 200 121 201
rect 119 200 120 201
rect 118 200 119 201
rect 117 200 118 201
rect 116 200 117 201
rect 115 200 116 201
rect 114 200 115 201
rect 113 200 114 201
rect 112 200 113 201
rect 111 200 112 201
rect 110 200 111 201
rect 109 200 110 201
rect 108 200 109 201
rect 107 200 108 201
rect 106 200 107 201
rect 105 200 106 201
rect 104 200 105 201
rect 103 200 104 201
rect 102 200 103 201
rect 101 200 102 201
rect 100 200 101 201
rect 99 200 100 201
rect 98 200 99 201
rect 97 200 98 201
rect 96 200 97 201
rect 95 200 96 201
rect 94 200 95 201
rect 93 200 94 201
rect 92 200 93 201
rect 91 200 92 201
rect 90 200 91 201
rect 89 200 90 201
rect 88 200 89 201
rect 87 200 88 201
rect 86 200 87 201
rect 85 200 86 201
rect 84 200 85 201
rect 83 200 84 201
rect 82 200 83 201
rect 81 200 82 201
rect 80 200 81 201
rect 79 200 80 201
rect 78 200 79 201
rect 77 200 78 201
rect 76 200 77 201
rect 75 200 76 201
rect 74 200 75 201
rect 73 200 74 201
rect 72 200 73 201
rect 71 200 72 201
rect 54 200 55 201
rect 53 200 54 201
rect 52 200 53 201
rect 51 200 52 201
rect 50 200 51 201
rect 49 200 50 201
rect 48 200 49 201
rect 47 200 48 201
rect 46 200 47 201
rect 45 200 46 201
rect 44 200 45 201
rect 43 200 44 201
rect 42 200 43 201
rect 41 200 42 201
rect 40 200 41 201
rect 39 200 40 201
rect 38 200 39 201
rect 37 200 38 201
rect 36 200 37 201
rect 35 200 36 201
rect 34 200 35 201
rect 33 200 34 201
rect 32 200 33 201
rect 31 200 32 201
rect 30 200 31 201
rect 29 200 30 201
rect 28 200 29 201
rect 27 200 28 201
rect 26 200 27 201
rect 25 200 26 201
rect 24 200 25 201
rect 23 200 24 201
rect 22 200 23 201
rect 21 200 22 201
rect 20 200 21 201
rect 19 200 20 201
rect 18 200 19 201
rect 17 200 18 201
rect 16 200 17 201
rect 15 200 16 201
rect 14 200 15 201
rect 13 200 14 201
rect 12 200 13 201
rect 11 200 12 201
rect 480 201 481 202
rect 470 201 471 202
rect 469 201 470 202
rect 460 201 461 202
rect 397 201 398 202
rect 396 201 397 202
rect 395 201 396 202
rect 350 201 351 202
rect 349 201 350 202
rect 348 201 349 202
rect 347 201 348 202
rect 346 201 347 202
rect 345 201 346 202
rect 344 201 345 202
rect 343 201 344 202
rect 342 201 343 202
rect 341 201 342 202
rect 340 201 341 202
rect 339 201 340 202
rect 338 201 339 202
rect 337 201 338 202
rect 336 201 337 202
rect 335 201 336 202
rect 334 201 335 202
rect 333 201 334 202
rect 332 201 333 202
rect 331 201 332 202
rect 330 201 331 202
rect 329 201 330 202
rect 328 201 329 202
rect 327 201 328 202
rect 326 201 327 202
rect 325 201 326 202
rect 324 201 325 202
rect 323 201 324 202
rect 322 201 323 202
rect 321 201 322 202
rect 320 201 321 202
rect 319 201 320 202
rect 318 201 319 202
rect 317 201 318 202
rect 316 201 317 202
rect 315 201 316 202
rect 314 201 315 202
rect 313 201 314 202
rect 312 201 313 202
rect 311 201 312 202
rect 310 201 311 202
rect 309 201 310 202
rect 308 201 309 202
rect 307 201 308 202
rect 306 201 307 202
rect 305 201 306 202
rect 304 201 305 202
rect 303 201 304 202
rect 302 201 303 202
rect 301 201 302 202
rect 300 201 301 202
rect 299 201 300 202
rect 298 201 299 202
rect 297 201 298 202
rect 296 201 297 202
rect 295 201 296 202
rect 294 201 295 202
rect 293 201 294 202
rect 292 201 293 202
rect 291 201 292 202
rect 290 201 291 202
rect 289 201 290 202
rect 288 201 289 202
rect 287 201 288 202
rect 286 201 287 202
rect 285 201 286 202
rect 284 201 285 202
rect 283 201 284 202
rect 282 201 283 202
rect 281 201 282 202
rect 280 201 281 202
rect 279 201 280 202
rect 278 201 279 202
rect 277 201 278 202
rect 276 201 277 202
rect 275 201 276 202
rect 274 201 275 202
rect 273 201 274 202
rect 272 201 273 202
rect 271 201 272 202
rect 270 201 271 202
rect 269 201 270 202
rect 268 201 269 202
rect 267 201 268 202
rect 266 201 267 202
rect 265 201 266 202
rect 264 201 265 202
rect 263 201 264 202
rect 262 201 263 202
rect 261 201 262 202
rect 260 201 261 202
rect 249 201 250 202
rect 248 201 249 202
rect 247 201 248 202
rect 246 201 247 202
rect 245 201 246 202
rect 244 201 245 202
rect 243 201 244 202
rect 242 201 243 202
rect 241 201 242 202
rect 240 201 241 202
rect 239 201 240 202
rect 238 201 239 202
rect 237 201 238 202
rect 236 201 237 202
rect 235 201 236 202
rect 234 201 235 202
rect 233 201 234 202
rect 232 201 233 202
rect 231 201 232 202
rect 230 201 231 202
rect 229 201 230 202
rect 228 201 229 202
rect 227 201 228 202
rect 226 201 227 202
rect 225 201 226 202
rect 224 201 225 202
rect 223 201 224 202
rect 222 201 223 202
rect 221 201 222 202
rect 220 201 221 202
rect 219 201 220 202
rect 218 201 219 202
rect 217 201 218 202
rect 216 201 217 202
rect 215 201 216 202
rect 214 201 215 202
rect 213 201 214 202
rect 212 201 213 202
rect 211 201 212 202
rect 210 201 211 202
rect 209 201 210 202
rect 208 201 209 202
rect 180 201 181 202
rect 179 201 180 202
rect 178 201 179 202
rect 177 201 178 202
rect 176 201 177 202
rect 175 201 176 202
rect 174 201 175 202
rect 173 201 174 202
rect 172 201 173 202
rect 171 201 172 202
rect 170 201 171 202
rect 169 201 170 202
rect 168 201 169 202
rect 167 201 168 202
rect 166 201 167 202
rect 165 201 166 202
rect 164 201 165 202
rect 163 201 164 202
rect 162 201 163 202
rect 161 201 162 202
rect 160 201 161 202
rect 159 201 160 202
rect 158 201 159 202
rect 157 201 158 202
rect 156 201 157 202
rect 155 201 156 202
rect 154 201 155 202
rect 153 201 154 202
rect 152 201 153 202
rect 151 201 152 202
rect 150 201 151 202
rect 149 201 150 202
rect 148 201 149 202
rect 147 201 148 202
rect 146 201 147 202
rect 145 201 146 202
rect 144 201 145 202
rect 143 201 144 202
rect 142 201 143 202
rect 141 201 142 202
rect 140 201 141 202
rect 139 201 140 202
rect 138 201 139 202
rect 137 201 138 202
rect 136 201 137 202
rect 135 201 136 202
rect 134 201 135 202
rect 133 201 134 202
rect 132 201 133 202
rect 131 201 132 202
rect 130 201 131 202
rect 129 201 130 202
rect 128 201 129 202
rect 127 201 128 202
rect 126 201 127 202
rect 125 201 126 202
rect 124 201 125 202
rect 123 201 124 202
rect 122 201 123 202
rect 121 201 122 202
rect 120 201 121 202
rect 119 201 120 202
rect 118 201 119 202
rect 117 201 118 202
rect 116 201 117 202
rect 115 201 116 202
rect 114 201 115 202
rect 113 201 114 202
rect 112 201 113 202
rect 111 201 112 202
rect 110 201 111 202
rect 109 201 110 202
rect 108 201 109 202
rect 107 201 108 202
rect 106 201 107 202
rect 105 201 106 202
rect 104 201 105 202
rect 103 201 104 202
rect 102 201 103 202
rect 101 201 102 202
rect 100 201 101 202
rect 99 201 100 202
rect 98 201 99 202
rect 97 201 98 202
rect 96 201 97 202
rect 95 201 96 202
rect 94 201 95 202
rect 93 201 94 202
rect 92 201 93 202
rect 91 201 92 202
rect 90 201 91 202
rect 89 201 90 202
rect 88 201 89 202
rect 87 201 88 202
rect 86 201 87 202
rect 85 201 86 202
rect 84 201 85 202
rect 83 201 84 202
rect 82 201 83 202
rect 81 201 82 202
rect 80 201 81 202
rect 79 201 80 202
rect 78 201 79 202
rect 77 201 78 202
rect 76 201 77 202
rect 75 201 76 202
rect 74 201 75 202
rect 73 201 74 202
rect 72 201 73 202
rect 55 201 56 202
rect 54 201 55 202
rect 53 201 54 202
rect 52 201 53 202
rect 51 201 52 202
rect 50 201 51 202
rect 49 201 50 202
rect 48 201 49 202
rect 47 201 48 202
rect 46 201 47 202
rect 45 201 46 202
rect 44 201 45 202
rect 43 201 44 202
rect 42 201 43 202
rect 41 201 42 202
rect 40 201 41 202
rect 39 201 40 202
rect 38 201 39 202
rect 37 201 38 202
rect 36 201 37 202
rect 35 201 36 202
rect 34 201 35 202
rect 33 201 34 202
rect 32 201 33 202
rect 31 201 32 202
rect 30 201 31 202
rect 29 201 30 202
rect 28 201 29 202
rect 27 201 28 202
rect 26 201 27 202
rect 25 201 26 202
rect 24 201 25 202
rect 23 201 24 202
rect 22 201 23 202
rect 21 201 22 202
rect 20 201 21 202
rect 19 201 20 202
rect 18 201 19 202
rect 17 201 18 202
rect 16 201 17 202
rect 15 201 16 202
rect 14 201 15 202
rect 13 201 14 202
rect 12 201 13 202
rect 11 201 12 202
rect 480 202 481 203
rect 470 202 471 203
rect 469 202 470 203
rect 460 202 461 203
rect 397 202 398 203
rect 396 202 397 203
rect 395 202 396 203
rect 350 202 351 203
rect 349 202 350 203
rect 348 202 349 203
rect 347 202 348 203
rect 346 202 347 203
rect 345 202 346 203
rect 344 202 345 203
rect 343 202 344 203
rect 342 202 343 203
rect 341 202 342 203
rect 340 202 341 203
rect 339 202 340 203
rect 338 202 339 203
rect 337 202 338 203
rect 336 202 337 203
rect 335 202 336 203
rect 334 202 335 203
rect 333 202 334 203
rect 332 202 333 203
rect 331 202 332 203
rect 330 202 331 203
rect 329 202 330 203
rect 328 202 329 203
rect 327 202 328 203
rect 326 202 327 203
rect 325 202 326 203
rect 324 202 325 203
rect 323 202 324 203
rect 322 202 323 203
rect 321 202 322 203
rect 320 202 321 203
rect 319 202 320 203
rect 318 202 319 203
rect 317 202 318 203
rect 316 202 317 203
rect 315 202 316 203
rect 314 202 315 203
rect 313 202 314 203
rect 312 202 313 203
rect 311 202 312 203
rect 310 202 311 203
rect 309 202 310 203
rect 308 202 309 203
rect 307 202 308 203
rect 306 202 307 203
rect 305 202 306 203
rect 304 202 305 203
rect 303 202 304 203
rect 302 202 303 203
rect 301 202 302 203
rect 300 202 301 203
rect 299 202 300 203
rect 298 202 299 203
rect 297 202 298 203
rect 296 202 297 203
rect 295 202 296 203
rect 294 202 295 203
rect 293 202 294 203
rect 292 202 293 203
rect 291 202 292 203
rect 290 202 291 203
rect 289 202 290 203
rect 288 202 289 203
rect 287 202 288 203
rect 286 202 287 203
rect 285 202 286 203
rect 284 202 285 203
rect 283 202 284 203
rect 282 202 283 203
rect 281 202 282 203
rect 280 202 281 203
rect 279 202 280 203
rect 278 202 279 203
rect 277 202 278 203
rect 276 202 277 203
rect 275 202 276 203
rect 274 202 275 203
rect 273 202 274 203
rect 272 202 273 203
rect 271 202 272 203
rect 270 202 271 203
rect 269 202 270 203
rect 268 202 269 203
rect 267 202 268 203
rect 266 202 267 203
rect 265 202 266 203
rect 264 202 265 203
rect 263 202 264 203
rect 262 202 263 203
rect 261 202 262 203
rect 260 202 261 203
rect 259 202 260 203
rect 258 202 259 203
rect 249 202 250 203
rect 248 202 249 203
rect 247 202 248 203
rect 246 202 247 203
rect 245 202 246 203
rect 244 202 245 203
rect 243 202 244 203
rect 242 202 243 203
rect 241 202 242 203
rect 240 202 241 203
rect 239 202 240 203
rect 238 202 239 203
rect 237 202 238 203
rect 236 202 237 203
rect 235 202 236 203
rect 234 202 235 203
rect 233 202 234 203
rect 232 202 233 203
rect 231 202 232 203
rect 230 202 231 203
rect 229 202 230 203
rect 228 202 229 203
rect 227 202 228 203
rect 226 202 227 203
rect 225 202 226 203
rect 224 202 225 203
rect 223 202 224 203
rect 222 202 223 203
rect 221 202 222 203
rect 220 202 221 203
rect 219 202 220 203
rect 218 202 219 203
rect 217 202 218 203
rect 216 202 217 203
rect 215 202 216 203
rect 214 202 215 203
rect 213 202 214 203
rect 212 202 213 203
rect 211 202 212 203
rect 210 202 211 203
rect 209 202 210 203
rect 208 202 209 203
rect 207 202 208 203
rect 179 202 180 203
rect 178 202 179 203
rect 177 202 178 203
rect 176 202 177 203
rect 175 202 176 203
rect 174 202 175 203
rect 173 202 174 203
rect 172 202 173 203
rect 171 202 172 203
rect 170 202 171 203
rect 169 202 170 203
rect 168 202 169 203
rect 167 202 168 203
rect 166 202 167 203
rect 165 202 166 203
rect 164 202 165 203
rect 163 202 164 203
rect 162 202 163 203
rect 161 202 162 203
rect 160 202 161 203
rect 159 202 160 203
rect 158 202 159 203
rect 157 202 158 203
rect 156 202 157 203
rect 155 202 156 203
rect 154 202 155 203
rect 153 202 154 203
rect 152 202 153 203
rect 151 202 152 203
rect 150 202 151 203
rect 149 202 150 203
rect 148 202 149 203
rect 147 202 148 203
rect 146 202 147 203
rect 145 202 146 203
rect 144 202 145 203
rect 143 202 144 203
rect 142 202 143 203
rect 141 202 142 203
rect 140 202 141 203
rect 139 202 140 203
rect 138 202 139 203
rect 137 202 138 203
rect 136 202 137 203
rect 135 202 136 203
rect 134 202 135 203
rect 133 202 134 203
rect 132 202 133 203
rect 131 202 132 203
rect 130 202 131 203
rect 129 202 130 203
rect 128 202 129 203
rect 127 202 128 203
rect 126 202 127 203
rect 125 202 126 203
rect 124 202 125 203
rect 123 202 124 203
rect 122 202 123 203
rect 121 202 122 203
rect 120 202 121 203
rect 119 202 120 203
rect 118 202 119 203
rect 117 202 118 203
rect 116 202 117 203
rect 115 202 116 203
rect 114 202 115 203
rect 113 202 114 203
rect 112 202 113 203
rect 111 202 112 203
rect 110 202 111 203
rect 109 202 110 203
rect 108 202 109 203
rect 107 202 108 203
rect 106 202 107 203
rect 105 202 106 203
rect 104 202 105 203
rect 103 202 104 203
rect 102 202 103 203
rect 101 202 102 203
rect 100 202 101 203
rect 99 202 100 203
rect 98 202 99 203
rect 97 202 98 203
rect 96 202 97 203
rect 95 202 96 203
rect 94 202 95 203
rect 93 202 94 203
rect 92 202 93 203
rect 91 202 92 203
rect 90 202 91 203
rect 89 202 90 203
rect 88 202 89 203
rect 87 202 88 203
rect 86 202 87 203
rect 85 202 86 203
rect 84 202 85 203
rect 83 202 84 203
rect 82 202 83 203
rect 81 202 82 203
rect 80 202 81 203
rect 79 202 80 203
rect 78 202 79 203
rect 77 202 78 203
rect 76 202 77 203
rect 75 202 76 203
rect 74 202 75 203
rect 73 202 74 203
rect 56 202 57 203
rect 55 202 56 203
rect 54 202 55 203
rect 53 202 54 203
rect 52 202 53 203
rect 51 202 52 203
rect 50 202 51 203
rect 49 202 50 203
rect 48 202 49 203
rect 47 202 48 203
rect 46 202 47 203
rect 45 202 46 203
rect 44 202 45 203
rect 43 202 44 203
rect 42 202 43 203
rect 41 202 42 203
rect 40 202 41 203
rect 39 202 40 203
rect 38 202 39 203
rect 37 202 38 203
rect 36 202 37 203
rect 35 202 36 203
rect 34 202 35 203
rect 33 202 34 203
rect 32 202 33 203
rect 31 202 32 203
rect 30 202 31 203
rect 29 202 30 203
rect 28 202 29 203
rect 27 202 28 203
rect 26 202 27 203
rect 25 202 26 203
rect 24 202 25 203
rect 23 202 24 203
rect 22 202 23 203
rect 21 202 22 203
rect 20 202 21 203
rect 19 202 20 203
rect 18 202 19 203
rect 17 202 18 203
rect 16 202 17 203
rect 15 202 16 203
rect 14 202 15 203
rect 13 202 14 203
rect 12 202 13 203
rect 11 202 12 203
rect 480 203 481 204
rect 472 203 473 204
rect 471 203 472 204
rect 470 203 471 204
rect 469 203 470 204
rect 468 203 469 204
rect 467 203 468 204
rect 461 203 462 204
rect 460 203 461 204
rect 396 203 397 204
rect 351 203 352 204
rect 350 203 351 204
rect 349 203 350 204
rect 348 203 349 204
rect 347 203 348 204
rect 346 203 347 204
rect 345 203 346 204
rect 344 203 345 204
rect 343 203 344 204
rect 342 203 343 204
rect 341 203 342 204
rect 340 203 341 204
rect 339 203 340 204
rect 338 203 339 204
rect 337 203 338 204
rect 336 203 337 204
rect 335 203 336 204
rect 334 203 335 204
rect 333 203 334 204
rect 332 203 333 204
rect 331 203 332 204
rect 330 203 331 204
rect 329 203 330 204
rect 328 203 329 204
rect 327 203 328 204
rect 326 203 327 204
rect 325 203 326 204
rect 324 203 325 204
rect 323 203 324 204
rect 322 203 323 204
rect 321 203 322 204
rect 320 203 321 204
rect 319 203 320 204
rect 318 203 319 204
rect 317 203 318 204
rect 316 203 317 204
rect 315 203 316 204
rect 314 203 315 204
rect 313 203 314 204
rect 312 203 313 204
rect 311 203 312 204
rect 310 203 311 204
rect 309 203 310 204
rect 308 203 309 204
rect 307 203 308 204
rect 306 203 307 204
rect 305 203 306 204
rect 304 203 305 204
rect 303 203 304 204
rect 302 203 303 204
rect 301 203 302 204
rect 300 203 301 204
rect 299 203 300 204
rect 298 203 299 204
rect 297 203 298 204
rect 296 203 297 204
rect 295 203 296 204
rect 294 203 295 204
rect 293 203 294 204
rect 292 203 293 204
rect 291 203 292 204
rect 290 203 291 204
rect 289 203 290 204
rect 288 203 289 204
rect 287 203 288 204
rect 286 203 287 204
rect 285 203 286 204
rect 284 203 285 204
rect 283 203 284 204
rect 282 203 283 204
rect 281 203 282 204
rect 280 203 281 204
rect 279 203 280 204
rect 278 203 279 204
rect 277 203 278 204
rect 276 203 277 204
rect 275 203 276 204
rect 274 203 275 204
rect 273 203 274 204
rect 272 203 273 204
rect 271 203 272 204
rect 270 203 271 204
rect 269 203 270 204
rect 268 203 269 204
rect 267 203 268 204
rect 266 203 267 204
rect 265 203 266 204
rect 264 203 265 204
rect 263 203 264 204
rect 262 203 263 204
rect 261 203 262 204
rect 260 203 261 204
rect 259 203 260 204
rect 258 203 259 204
rect 257 203 258 204
rect 248 203 249 204
rect 247 203 248 204
rect 246 203 247 204
rect 245 203 246 204
rect 244 203 245 204
rect 243 203 244 204
rect 242 203 243 204
rect 241 203 242 204
rect 240 203 241 204
rect 239 203 240 204
rect 238 203 239 204
rect 237 203 238 204
rect 236 203 237 204
rect 235 203 236 204
rect 234 203 235 204
rect 233 203 234 204
rect 232 203 233 204
rect 231 203 232 204
rect 230 203 231 204
rect 229 203 230 204
rect 228 203 229 204
rect 227 203 228 204
rect 226 203 227 204
rect 225 203 226 204
rect 224 203 225 204
rect 223 203 224 204
rect 222 203 223 204
rect 221 203 222 204
rect 220 203 221 204
rect 219 203 220 204
rect 218 203 219 204
rect 217 203 218 204
rect 216 203 217 204
rect 215 203 216 204
rect 214 203 215 204
rect 213 203 214 204
rect 212 203 213 204
rect 211 203 212 204
rect 210 203 211 204
rect 209 203 210 204
rect 208 203 209 204
rect 207 203 208 204
rect 206 203 207 204
rect 177 203 178 204
rect 176 203 177 204
rect 175 203 176 204
rect 174 203 175 204
rect 173 203 174 204
rect 172 203 173 204
rect 171 203 172 204
rect 170 203 171 204
rect 169 203 170 204
rect 168 203 169 204
rect 167 203 168 204
rect 166 203 167 204
rect 165 203 166 204
rect 164 203 165 204
rect 163 203 164 204
rect 162 203 163 204
rect 161 203 162 204
rect 160 203 161 204
rect 159 203 160 204
rect 158 203 159 204
rect 157 203 158 204
rect 156 203 157 204
rect 155 203 156 204
rect 154 203 155 204
rect 153 203 154 204
rect 152 203 153 204
rect 151 203 152 204
rect 150 203 151 204
rect 149 203 150 204
rect 148 203 149 204
rect 147 203 148 204
rect 146 203 147 204
rect 145 203 146 204
rect 144 203 145 204
rect 143 203 144 204
rect 142 203 143 204
rect 141 203 142 204
rect 140 203 141 204
rect 139 203 140 204
rect 138 203 139 204
rect 137 203 138 204
rect 136 203 137 204
rect 135 203 136 204
rect 134 203 135 204
rect 133 203 134 204
rect 132 203 133 204
rect 131 203 132 204
rect 130 203 131 204
rect 129 203 130 204
rect 128 203 129 204
rect 127 203 128 204
rect 126 203 127 204
rect 125 203 126 204
rect 124 203 125 204
rect 123 203 124 204
rect 122 203 123 204
rect 121 203 122 204
rect 120 203 121 204
rect 119 203 120 204
rect 118 203 119 204
rect 117 203 118 204
rect 116 203 117 204
rect 115 203 116 204
rect 114 203 115 204
rect 113 203 114 204
rect 112 203 113 204
rect 111 203 112 204
rect 110 203 111 204
rect 109 203 110 204
rect 108 203 109 204
rect 107 203 108 204
rect 106 203 107 204
rect 105 203 106 204
rect 104 203 105 204
rect 103 203 104 204
rect 102 203 103 204
rect 101 203 102 204
rect 100 203 101 204
rect 99 203 100 204
rect 98 203 99 204
rect 97 203 98 204
rect 96 203 97 204
rect 95 203 96 204
rect 94 203 95 204
rect 93 203 94 204
rect 92 203 93 204
rect 91 203 92 204
rect 90 203 91 204
rect 89 203 90 204
rect 88 203 89 204
rect 87 203 88 204
rect 86 203 87 204
rect 85 203 86 204
rect 84 203 85 204
rect 83 203 84 204
rect 82 203 83 204
rect 81 203 82 204
rect 80 203 81 204
rect 79 203 80 204
rect 78 203 79 204
rect 77 203 78 204
rect 76 203 77 204
rect 75 203 76 204
rect 74 203 75 204
rect 73 203 74 204
rect 56 203 57 204
rect 55 203 56 204
rect 54 203 55 204
rect 53 203 54 204
rect 52 203 53 204
rect 51 203 52 204
rect 50 203 51 204
rect 49 203 50 204
rect 48 203 49 204
rect 47 203 48 204
rect 46 203 47 204
rect 45 203 46 204
rect 44 203 45 204
rect 43 203 44 204
rect 42 203 43 204
rect 41 203 42 204
rect 40 203 41 204
rect 39 203 40 204
rect 38 203 39 204
rect 37 203 38 204
rect 36 203 37 204
rect 35 203 36 204
rect 34 203 35 204
rect 33 203 34 204
rect 32 203 33 204
rect 31 203 32 204
rect 30 203 31 204
rect 29 203 30 204
rect 28 203 29 204
rect 27 203 28 204
rect 26 203 27 204
rect 25 203 26 204
rect 24 203 25 204
rect 23 203 24 204
rect 22 203 23 204
rect 21 203 22 204
rect 20 203 21 204
rect 19 203 20 204
rect 18 203 19 204
rect 17 203 18 204
rect 16 203 17 204
rect 15 203 16 204
rect 14 203 15 204
rect 13 203 14 204
rect 12 203 13 204
rect 11 203 12 204
rect 480 204 481 205
rect 479 204 480 205
rect 473 204 474 205
rect 472 204 473 205
rect 471 204 472 205
rect 470 204 471 205
rect 469 204 470 205
rect 468 204 469 205
rect 467 204 468 205
rect 462 204 463 205
rect 461 204 462 205
rect 460 204 461 205
rect 352 204 353 205
rect 351 204 352 205
rect 350 204 351 205
rect 349 204 350 205
rect 348 204 349 205
rect 347 204 348 205
rect 346 204 347 205
rect 345 204 346 205
rect 344 204 345 205
rect 343 204 344 205
rect 342 204 343 205
rect 341 204 342 205
rect 340 204 341 205
rect 339 204 340 205
rect 338 204 339 205
rect 337 204 338 205
rect 336 204 337 205
rect 335 204 336 205
rect 334 204 335 205
rect 333 204 334 205
rect 332 204 333 205
rect 331 204 332 205
rect 330 204 331 205
rect 329 204 330 205
rect 328 204 329 205
rect 327 204 328 205
rect 326 204 327 205
rect 325 204 326 205
rect 324 204 325 205
rect 323 204 324 205
rect 322 204 323 205
rect 321 204 322 205
rect 320 204 321 205
rect 319 204 320 205
rect 318 204 319 205
rect 317 204 318 205
rect 316 204 317 205
rect 315 204 316 205
rect 314 204 315 205
rect 313 204 314 205
rect 312 204 313 205
rect 311 204 312 205
rect 310 204 311 205
rect 309 204 310 205
rect 308 204 309 205
rect 307 204 308 205
rect 306 204 307 205
rect 305 204 306 205
rect 304 204 305 205
rect 303 204 304 205
rect 302 204 303 205
rect 301 204 302 205
rect 300 204 301 205
rect 299 204 300 205
rect 298 204 299 205
rect 297 204 298 205
rect 296 204 297 205
rect 295 204 296 205
rect 294 204 295 205
rect 293 204 294 205
rect 292 204 293 205
rect 291 204 292 205
rect 290 204 291 205
rect 289 204 290 205
rect 288 204 289 205
rect 287 204 288 205
rect 286 204 287 205
rect 285 204 286 205
rect 284 204 285 205
rect 283 204 284 205
rect 282 204 283 205
rect 281 204 282 205
rect 280 204 281 205
rect 279 204 280 205
rect 278 204 279 205
rect 277 204 278 205
rect 276 204 277 205
rect 275 204 276 205
rect 274 204 275 205
rect 273 204 274 205
rect 272 204 273 205
rect 271 204 272 205
rect 270 204 271 205
rect 269 204 270 205
rect 268 204 269 205
rect 267 204 268 205
rect 266 204 267 205
rect 265 204 266 205
rect 264 204 265 205
rect 263 204 264 205
rect 262 204 263 205
rect 261 204 262 205
rect 260 204 261 205
rect 259 204 260 205
rect 258 204 259 205
rect 257 204 258 205
rect 256 204 257 205
rect 255 204 256 205
rect 247 204 248 205
rect 246 204 247 205
rect 245 204 246 205
rect 244 204 245 205
rect 243 204 244 205
rect 242 204 243 205
rect 241 204 242 205
rect 240 204 241 205
rect 239 204 240 205
rect 238 204 239 205
rect 237 204 238 205
rect 236 204 237 205
rect 235 204 236 205
rect 234 204 235 205
rect 233 204 234 205
rect 232 204 233 205
rect 231 204 232 205
rect 230 204 231 205
rect 229 204 230 205
rect 228 204 229 205
rect 227 204 228 205
rect 226 204 227 205
rect 225 204 226 205
rect 224 204 225 205
rect 223 204 224 205
rect 222 204 223 205
rect 221 204 222 205
rect 220 204 221 205
rect 219 204 220 205
rect 218 204 219 205
rect 217 204 218 205
rect 216 204 217 205
rect 215 204 216 205
rect 214 204 215 205
rect 213 204 214 205
rect 212 204 213 205
rect 211 204 212 205
rect 210 204 211 205
rect 209 204 210 205
rect 208 204 209 205
rect 207 204 208 205
rect 206 204 207 205
rect 205 204 206 205
rect 175 204 176 205
rect 174 204 175 205
rect 173 204 174 205
rect 172 204 173 205
rect 171 204 172 205
rect 170 204 171 205
rect 169 204 170 205
rect 168 204 169 205
rect 167 204 168 205
rect 166 204 167 205
rect 165 204 166 205
rect 164 204 165 205
rect 163 204 164 205
rect 162 204 163 205
rect 161 204 162 205
rect 160 204 161 205
rect 159 204 160 205
rect 158 204 159 205
rect 157 204 158 205
rect 156 204 157 205
rect 155 204 156 205
rect 154 204 155 205
rect 153 204 154 205
rect 152 204 153 205
rect 151 204 152 205
rect 150 204 151 205
rect 149 204 150 205
rect 148 204 149 205
rect 147 204 148 205
rect 146 204 147 205
rect 145 204 146 205
rect 144 204 145 205
rect 143 204 144 205
rect 142 204 143 205
rect 141 204 142 205
rect 140 204 141 205
rect 139 204 140 205
rect 138 204 139 205
rect 137 204 138 205
rect 136 204 137 205
rect 135 204 136 205
rect 134 204 135 205
rect 133 204 134 205
rect 132 204 133 205
rect 131 204 132 205
rect 130 204 131 205
rect 129 204 130 205
rect 128 204 129 205
rect 127 204 128 205
rect 126 204 127 205
rect 125 204 126 205
rect 124 204 125 205
rect 123 204 124 205
rect 122 204 123 205
rect 121 204 122 205
rect 120 204 121 205
rect 119 204 120 205
rect 118 204 119 205
rect 117 204 118 205
rect 116 204 117 205
rect 115 204 116 205
rect 114 204 115 205
rect 113 204 114 205
rect 112 204 113 205
rect 111 204 112 205
rect 110 204 111 205
rect 109 204 110 205
rect 108 204 109 205
rect 107 204 108 205
rect 106 204 107 205
rect 105 204 106 205
rect 104 204 105 205
rect 103 204 104 205
rect 102 204 103 205
rect 101 204 102 205
rect 100 204 101 205
rect 99 204 100 205
rect 98 204 99 205
rect 97 204 98 205
rect 96 204 97 205
rect 95 204 96 205
rect 94 204 95 205
rect 93 204 94 205
rect 92 204 93 205
rect 91 204 92 205
rect 90 204 91 205
rect 89 204 90 205
rect 88 204 89 205
rect 87 204 88 205
rect 86 204 87 205
rect 85 204 86 205
rect 84 204 85 205
rect 83 204 84 205
rect 82 204 83 205
rect 81 204 82 205
rect 80 204 81 205
rect 79 204 80 205
rect 78 204 79 205
rect 77 204 78 205
rect 76 204 77 205
rect 75 204 76 205
rect 74 204 75 205
rect 57 204 58 205
rect 56 204 57 205
rect 55 204 56 205
rect 54 204 55 205
rect 53 204 54 205
rect 52 204 53 205
rect 51 204 52 205
rect 50 204 51 205
rect 49 204 50 205
rect 48 204 49 205
rect 47 204 48 205
rect 46 204 47 205
rect 45 204 46 205
rect 44 204 45 205
rect 43 204 44 205
rect 42 204 43 205
rect 41 204 42 205
rect 40 204 41 205
rect 39 204 40 205
rect 38 204 39 205
rect 37 204 38 205
rect 36 204 37 205
rect 35 204 36 205
rect 34 204 35 205
rect 33 204 34 205
rect 32 204 33 205
rect 31 204 32 205
rect 30 204 31 205
rect 29 204 30 205
rect 28 204 29 205
rect 27 204 28 205
rect 26 204 27 205
rect 25 204 26 205
rect 24 204 25 205
rect 23 204 24 205
rect 22 204 23 205
rect 21 204 22 205
rect 20 204 21 205
rect 19 204 20 205
rect 18 204 19 205
rect 17 204 18 205
rect 16 204 17 205
rect 15 204 16 205
rect 14 204 15 205
rect 13 204 14 205
rect 12 204 13 205
rect 11 204 12 205
rect 10 204 11 205
rect 480 205 481 206
rect 479 205 480 206
rect 478 205 479 206
rect 464 205 465 206
rect 463 205 464 206
rect 462 205 463 206
rect 461 205 462 206
rect 460 205 461 206
rect 353 205 354 206
rect 352 205 353 206
rect 351 205 352 206
rect 350 205 351 206
rect 349 205 350 206
rect 348 205 349 206
rect 347 205 348 206
rect 346 205 347 206
rect 345 205 346 206
rect 344 205 345 206
rect 343 205 344 206
rect 342 205 343 206
rect 341 205 342 206
rect 340 205 341 206
rect 339 205 340 206
rect 338 205 339 206
rect 337 205 338 206
rect 336 205 337 206
rect 335 205 336 206
rect 334 205 335 206
rect 333 205 334 206
rect 332 205 333 206
rect 331 205 332 206
rect 330 205 331 206
rect 329 205 330 206
rect 328 205 329 206
rect 327 205 328 206
rect 326 205 327 206
rect 325 205 326 206
rect 324 205 325 206
rect 323 205 324 206
rect 322 205 323 206
rect 321 205 322 206
rect 320 205 321 206
rect 319 205 320 206
rect 318 205 319 206
rect 317 205 318 206
rect 316 205 317 206
rect 315 205 316 206
rect 314 205 315 206
rect 313 205 314 206
rect 312 205 313 206
rect 311 205 312 206
rect 310 205 311 206
rect 309 205 310 206
rect 308 205 309 206
rect 307 205 308 206
rect 306 205 307 206
rect 305 205 306 206
rect 304 205 305 206
rect 303 205 304 206
rect 302 205 303 206
rect 301 205 302 206
rect 300 205 301 206
rect 299 205 300 206
rect 298 205 299 206
rect 297 205 298 206
rect 296 205 297 206
rect 295 205 296 206
rect 294 205 295 206
rect 293 205 294 206
rect 292 205 293 206
rect 291 205 292 206
rect 290 205 291 206
rect 289 205 290 206
rect 288 205 289 206
rect 287 205 288 206
rect 286 205 287 206
rect 285 205 286 206
rect 284 205 285 206
rect 283 205 284 206
rect 282 205 283 206
rect 281 205 282 206
rect 280 205 281 206
rect 279 205 280 206
rect 278 205 279 206
rect 277 205 278 206
rect 276 205 277 206
rect 275 205 276 206
rect 274 205 275 206
rect 273 205 274 206
rect 272 205 273 206
rect 271 205 272 206
rect 270 205 271 206
rect 269 205 270 206
rect 268 205 269 206
rect 267 205 268 206
rect 266 205 267 206
rect 265 205 266 206
rect 264 205 265 206
rect 263 205 264 206
rect 262 205 263 206
rect 261 205 262 206
rect 260 205 261 206
rect 259 205 260 206
rect 258 205 259 206
rect 257 205 258 206
rect 256 205 257 206
rect 255 205 256 206
rect 254 205 255 206
rect 253 205 254 206
rect 247 205 248 206
rect 246 205 247 206
rect 245 205 246 206
rect 244 205 245 206
rect 243 205 244 206
rect 242 205 243 206
rect 241 205 242 206
rect 240 205 241 206
rect 239 205 240 206
rect 238 205 239 206
rect 237 205 238 206
rect 236 205 237 206
rect 235 205 236 206
rect 234 205 235 206
rect 233 205 234 206
rect 232 205 233 206
rect 231 205 232 206
rect 230 205 231 206
rect 229 205 230 206
rect 228 205 229 206
rect 227 205 228 206
rect 226 205 227 206
rect 225 205 226 206
rect 224 205 225 206
rect 223 205 224 206
rect 222 205 223 206
rect 221 205 222 206
rect 220 205 221 206
rect 219 205 220 206
rect 218 205 219 206
rect 217 205 218 206
rect 216 205 217 206
rect 215 205 216 206
rect 214 205 215 206
rect 213 205 214 206
rect 212 205 213 206
rect 211 205 212 206
rect 210 205 211 206
rect 209 205 210 206
rect 208 205 209 206
rect 207 205 208 206
rect 206 205 207 206
rect 205 205 206 206
rect 204 205 205 206
rect 173 205 174 206
rect 172 205 173 206
rect 171 205 172 206
rect 170 205 171 206
rect 169 205 170 206
rect 168 205 169 206
rect 167 205 168 206
rect 166 205 167 206
rect 165 205 166 206
rect 164 205 165 206
rect 163 205 164 206
rect 162 205 163 206
rect 161 205 162 206
rect 160 205 161 206
rect 159 205 160 206
rect 158 205 159 206
rect 157 205 158 206
rect 156 205 157 206
rect 155 205 156 206
rect 154 205 155 206
rect 153 205 154 206
rect 152 205 153 206
rect 151 205 152 206
rect 150 205 151 206
rect 149 205 150 206
rect 148 205 149 206
rect 147 205 148 206
rect 146 205 147 206
rect 145 205 146 206
rect 144 205 145 206
rect 143 205 144 206
rect 142 205 143 206
rect 141 205 142 206
rect 140 205 141 206
rect 139 205 140 206
rect 138 205 139 206
rect 137 205 138 206
rect 136 205 137 206
rect 135 205 136 206
rect 134 205 135 206
rect 133 205 134 206
rect 132 205 133 206
rect 131 205 132 206
rect 130 205 131 206
rect 129 205 130 206
rect 128 205 129 206
rect 127 205 128 206
rect 126 205 127 206
rect 125 205 126 206
rect 124 205 125 206
rect 123 205 124 206
rect 122 205 123 206
rect 121 205 122 206
rect 120 205 121 206
rect 119 205 120 206
rect 118 205 119 206
rect 117 205 118 206
rect 116 205 117 206
rect 115 205 116 206
rect 114 205 115 206
rect 113 205 114 206
rect 112 205 113 206
rect 111 205 112 206
rect 110 205 111 206
rect 109 205 110 206
rect 108 205 109 206
rect 107 205 108 206
rect 106 205 107 206
rect 105 205 106 206
rect 104 205 105 206
rect 103 205 104 206
rect 102 205 103 206
rect 101 205 102 206
rect 100 205 101 206
rect 99 205 100 206
rect 98 205 99 206
rect 97 205 98 206
rect 96 205 97 206
rect 95 205 96 206
rect 94 205 95 206
rect 93 205 94 206
rect 92 205 93 206
rect 91 205 92 206
rect 90 205 91 206
rect 89 205 90 206
rect 88 205 89 206
rect 87 205 88 206
rect 86 205 87 206
rect 85 205 86 206
rect 84 205 85 206
rect 83 205 84 206
rect 82 205 83 206
rect 81 205 82 206
rect 80 205 81 206
rect 79 205 80 206
rect 78 205 79 206
rect 77 205 78 206
rect 76 205 77 206
rect 75 205 76 206
rect 58 205 59 206
rect 57 205 58 206
rect 56 205 57 206
rect 55 205 56 206
rect 54 205 55 206
rect 53 205 54 206
rect 52 205 53 206
rect 51 205 52 206
rect 50 205 51 206
rect 49 205 50 206
rect 48 205 49 206
rect 47 205 48 206
rect 46 205 47 206
rect 45 205 46 206
rect 44 205 45 206
rect 43 205 44 206
rect 42 205 43 206
rect 41 205 42 206
rect 40 205 41 206
rect 39 205 40 206
rect 38 205 39 206
rect 37 205 38 206
rect 36 205 37 206
rect 35 205 36 206
rect 34 205 35 206
rect 33 205 34 206
rect 32 205 33 206
rect 31 205 32 206
rect 30 205 31 206
rect 29 205 30 206
rect 28 205 29 206
rect 27 205 28 206
rect 26 205 27 206
rect 25 205 26 206
rect 24 205 25 206
rect 23 205 24 206
rect 22 205 23 206
rect 21 205 22 206
rect 20 205 21 206
rect 19 205 20 206
rect 18 205 19 206
rect 17 205 18 206
rect 16 205 17 206
rect 15 205 16 206
rect 14 205 15 206
rect 13 205 14 206
rect 12 205 13 206
rect 11 205 12 206
rect 10 205 11 206
rect 480 206 481 207
rect 479 206 480 207
rect 478 206 479 207
rect 477 206 478 207
rect 476 206 477 207
rect 464 206 465 207
rect 463 206 464 207
rect 462 206 463 207
rect 353 206 354 207
rect 352 206 353 207
rect 351 206 352 207
rect 350 206 351 207
rect 349 206 350 207
rect 348 206 349 207
rect 347 206 348 207
rect 346 206 347 207
rect 345 206 346 207
rect 344 206 345 207
rect 343 206 344 207
rect 342 206 343 207
rect 341 206 342 207
rect 340 206 341 207
rect 339 206 340 207
rect 338 206 339 207
rect 337 206 338 207
rect 336 206 337 207
rect 335 206 336 207
rect 334 206 335 207
rect 333 206 334 207
rect 332 206 333 207
rect 331 206 332 207
rect 330 206 331 207
rect 329 206 330 207
rect 328 206 329 207
rect 327 206 328 207
rect 326 206 327 207
rect 325 206 326 207
rect 324 206 325 207
rect 323 206 324 207
rect 322 206 323 207
rect 321 206 322 207
rect 320 206 321 207
rect 319 206 320 207
rect 318 206 319 207
rect 317 206 318 207
rect 316 206 317 207
rect 315 206 316 207
rect 314 206 315 207
rect 313 206 314 207
rect 312 206 313 207
rect 311 206 312 207
rect 310 206 311 207
rect 309 206 310 207
rect 308 206 309 207
rect 307 206 308 207
rect 306 206 307 207
rect 305 206 306 207
rect 304 206 305 207
rect 303 206 304 207
rect 302 206 303 207
rect 301 206 302 207
rect 300 206 301 207
rect 299 206 300 207
rect 298 206 299 207
rect 297 206 298 207
rect 296 206 297 207
rect 295 206 296 207
rect 294 206 295 207
rect 293 206 294 207
rect 292 206 293 207
rect 291 206 292 207
rect 290 206 291 207
rect 289 206 290 207
rect 288 206 289 207
rect 287 206 288 207
rect 286 206 287 207
rect 285 206 286 207
rect 284 206 285 207
rect 283 206 284 207
rect 282 206 283 207
rect 281 206 282 207
rect 280 206 281 207
rect 279 206 280 207
rect 278 206 279 207
rect 277 206 278 207
rect 276 206 277 207
rect 275 206 276 207
rect 274 206 275 207
rect 273 206 274 207
rect 272 206 273 207
rect 271 206 272 207
rect 270 206 271 207
rect 269 206 270 207
rect 268 206 269 207
rect 267 206 268 207
rect 266 206 267 207
rect 265 206 266 207
rect 264 206 265 207
rect 263 206 264 207
rect 262 206 263 207
rect 261 206 262 207
rect 260 206 261 207
rect 259 206 260 207
rect 258 206 259 207
rect 257 206 258 207
rect 256 206 257 207
rect 255 206 256 207
rect 254 206 255 207
rect 253 206 254 207
rect 252 206 253 207
rect 251 206 252 207
rect 246 206 247 207
rect 245 206 246 207
rect 244 206 245 207
rect 243 206 244 207
rect 242 206 243 207
rect 241 206 242 207
rect 240 206 241 207
rect 239 206 240 207
rect 238 206 239 207
rect 237 206 238 207
rect 236 206 237 207
rect 235 206 236 207
rect 234 206 235 207
rect 233 206 234 207
rect 232 206 233 207
rect 231 206 232 207
rect 230 206 231 207
rect 229 206 230 207
rect 228 206 229 207
rect 227 206 228 207
rect 226 206 227 207
rect 225 206 226 207
rect 224 206 225 207
rect 223 206 224 207
rect 222 206 223 207
rect 221 206 222 207
rect 220 206 221 207
rect 219 206 220 207
rect 218 206 219 207
rect 217 206 218 207
rect 216 206 217 207
rect 215 206 216 207
rect 214 206 215 207
rect 213 206 214 207
rect 212 206 213 207
rect 211 206 212 207
rect 210 206 211 207
rect 209 206 210 207
rect 208 206 209 207
rect 207 206 208 207
rect 206 206 207 207
rect 205 206 206 207
rect 204 206 205 207
rect 203 206 204 207
rect 171 206 172 207
rect 170 206 171 207
rect 169 206 170 207
rect 168 206 169 207
rect 167 206 168 207
rect 166 206 167 207
rect 165 206 166 207
rect 164 206 165 207
rect 163 206 164 207
rect 162 206 163 207
rect 161 206 162 207
rect 160 206 161 207
rect 159 206 160 207
rect 158 206 159 207
rect 157 206 158 207
rect 156 206 157 207
rect 155 206 156 207
rect 154 206 155 207
rect 153 206 154 207
rect 152 206 153 207
rect 151 206 152 207
rect 150 206 151 207
rect 149 206 150 207
rect 148 206 149 207
rect 147 206 148 207
rect 146 206 147 207
rect 145 206 146 207
rect 144 206 145 207
rect 143 206 144 207
rect 142 206 143 207
rect 141 206 142 207
rect 140 206 141 207
rect 139 206 140 207
rect 138 206 139 207
rect 137 206 138 207
rect 136 206 137 207
rect 135 206 136 207
rect 134 206 135 207
rect 133 206 134 207
rect 132 206 133 207
rect 131 206 132 207
rect 130 206 131 207
rect 129 206 130 207
rect 128 206 129 207
rect 127 206 128 207
rect 126 206 127 207
rect 125 206 126 207
rect 124 206 125 207
rect 123 206 124 207
rect 122 206 123 207
rect 121 206 122 207
rect 120 206 121 207
rect 119 206 120 207
rect 118 206 119 207
rect 117 206 118 207
rect 116 206 117 207
rect 115 206 116 207
rect 114 206 115 207
rect 113 206 114 207
rect 112 206 113 207
rect 111 206 112 207
rect 110 206 111 207
rect 109 206 110 207
rect 108 206 109 207
rect 107 206 108 207
rect 106 206 107 207
rect 105 206 106 207
rect 104 206 105 207
rect 103 206 104 207
rect 102 206 103 207
rect 101 206 102 207
rect 100 206 101 207
rect 99 206 100 207
rect 98 206 99 207
rect 97 206 98 207
rect 96 206 97 207
rect 95 206 96 207
rect 94 206 95 207
rect 93 206 94 207
rect 92 206 93 207
rect 91 206 92 207
rect 90 206 91 207
rect 89 206 90 207
rect 88 206 89 207
rect 87 206 88 207
rect 86 206 87 207
rect 85 206 86 207
rect 84 206 85 207
rect 83 206 84 207
rect 82 206 83 207
rect 81 206 82 207
rect 80 206 81 207
rect 79 206 80 207
rect 78 206 79 207
rect 77 206 78 207
rect 76 206 77 207
rect 58 206 59 207
rect 57 206 58 207
rect 56 206 57 207
rect 55 206 56 207
rect 54 206 55 207
rect 53 206 54 207
rect 52 206 53 207
rect 51 206 52 207
rect 50 206 51 207
rect 49 206 50 207
rect 48 206 49 207
rect 47 206 48 207
rect 46 206 47 207
rect 45 206 46 207
rect 44 206 45 207
rect 43 206 44 207
rect 42 206 43 207
rect 41 206 42 207
rect 40 206 41 207
rect 39 206 40 207
rect 38 206 39 207
rect 37 206 38 207
rect 36 206 37 207
rect 35 206 36 207
rect 34 206 35 207
rect 33 206 34 207
rect 32 206 33 207
rect 31 206 32 207
rect 30 206 31 207
rect 29 206 30 207
rect 28 206 29 207
rect 27 206 28 207
rect 26 206 27 207
rect 25 206 26 207
rect 24 206 25 207
rect 23 206 24 207
rect 22 206 23 207
rect 21 206 22 207
rect 20 206 21 207
rect 19 206 20 207
rect 18 206 19 207
rect 17 206 18 207
rect 16 206 17 207
rect 15 206 16 207
rect 14 206 15 207
rect 13 206 14 207
rect 12 206 13 207
rect 11 206 12 207
rect 10 206 11 207
rect 479 207 480 208
rect 478 207 479 208
rect 477 207 478 208
rect 476 207 477 208
rect 475 207 476 208
rect 422 207 423 208
rect 421 207 422 208
rect 420 207 421 208
rect 419 207 420 208
rect 418 207 419 208
rect 417 207 418 208
rect 416 207 417 208
rect 415 207 416 208
rect 414 207 415 208
rect 413 207 414 208
rect 354 207 355 208
rect 353 207 354 208
rect 352 207 353 208
rect 351 207 352 208
rect 350 207 351 208
rect 349 207 350 208
rect 348 207 349 208
rect 347 207 348 208
rect 346 207 347 208
rect 345 207 346 208
rect 344 207 345 208
rect 343 207 344 208
rect 342 207 343 208
rect 341 207 342 208
rect 340 207 341 208
rect 339 207 340 208
rect 338 207 339 208
rect 337 207 338 208
rect 336 207 337 208
rect 335 207 336 208
rect 334 207 335 208
rect 333 207 334 208
rect 332 207 333 208
rect 331 207 332 208
rect 330 207 331 208
rect 329 207 330 208
rect 328 207 329 208
rect 327 207 328 208
rect 326 207 327 208
rect 325 207 326 208
rect 324 207 325 208
rect 323 207 324 208
rect 322 207 323 208
rect 321 207 322 208
rect 320 207 321 208
rect 319 207 320 208
rect 318 207 319 208
rect 317 207 318 208
rect 316 207 317 208
rect 315 207 316 208
rect 314 207 315 208
rect 313 207 314 208
rect 312 207 313 208
rect 311 207 312 208
rect 310 207 311 208
rect 309 207 310 208
rect 308 207 309 208
rect 307 207 308 208
rect 306 207 307 208
rect 305 207 306 208
rect 304 207 305 208
rect 303 207 304 208
rect 302 207 303 208
rect 301 207 302 208
rect 300 207 301 208
rect 299 207 300 208
rect 298 207 299 208
rect 297 207 298 208
rect 296 207 297 208
rect 295 207 296 208
rect 294 207 295 208
rect 293 207 294 208
rect 292 207 293 208
rect 291 207 292 208
rect 290 207 291 208
rect 289 207 290 208
rect 288 207 289 208
rect 287 207 288 208
rect 286 207 287 208
rect 285 207 286 208
rect 284 207 285 208
rect 283 207 284 208
rect 282 207 283 208
rect 281 207 282 208
rect 280 207 281 208
rect 279 207 280 208
rect 278 207 279 208
rect 277 207 278 208
rect 276 207 277 208
rect 275 207 276 208
rect 274 207 275 208
rect 273 207 274 208
rect 272 207 273 208
rect 271 207 272 208
rect 270 207 271 208
rect 269 207 270 208
rect 268 207 269 208
rect 267 207 268 208
rect 266 207 267 208
rect 265 207 266 208
rect 264 207 265 208
rect 263 207 264 208
rect 262 207 263 208
rect 261 207 262 208
rect 260 207 261 208
rect 259 207 260 208
rect 258 207 259 208
rect 257 207 258 208
rect 256 207 257 208
rect 255 207 256 208
rect 254 207 255 208
rect 253 207 254 208
rect 252 207 253 208
rect 251 207 252 208
rect 250 207 251 208
rect 249 207 250 208
rect 248 207 249 208
rect 247 207 248 208
rect 246 207 247 208
rect 245 207 246 208
rect 244 207 245 208
rect 243 207 244 208
rect 242 207 243 208
rect 241 207 242 208
rect 240 207 241 208
rect 239 207 240 208
rect 238 207 239 208
rect 237 207 238 208
rect 236 207 237 208
rect 235 207 236 208
rect 234 207 235 208
rect 233 207 234 208
rect 232 207 233 208
rect 231 207 232 208
rect 230 207 231 208
rect 229 207 230 208
rect 228 207 229 208
rect 227 207 228 208
rect 226 207 227 208
rect 225 207 226 208
rect 224 207 225 208
rect 223 207 224 208
rect 222 207 223 208
rect 221 207 222 208
rect 220 207 221 208
rect 219 207 220 208
rect 218 207 219 208
rect 217 207 218 208
rect 216 207 217 208
rect 215 207 216 208
rect 214 207 215 208
rect 213 207 214 208
rect 212 207 213 208
rect 211 207 212 208
rect 210 207 211 208
rect 209 207 210 208
rect 208 207 209 208
rect 207 207 208 208
rect 206 207 207 208
rect 205 207 206 208
rect 204 207 205 208
rect 203 207 204 208
rect 202 207 203 208
rect 169 207 170 208
rect 168 207 169 208
rect 167 207 168 208
rect 166 207 167 208
rect 165 207 166 208
rect 164 207 165 208
rect 163 207 164 208
rect 162 207 163 208
rect 161 207 162 208
rect 160 207 161 208
rect 159 207 160 208
rect 158 207 159 208
rect 157 207 158 208
rect 156 207 157 208
rect 155 207 156 208
rect 154 207 155 208
rect 153 207 154 208
rect 152 207 153 208
rect 151 207 152 208
rect 150 207 151 208
rect 149 207 150 208
rect 148 207 149 208
rect 147 207 148 208
rect 146 207 147 208
rect 145 207 146 208
rect 144 207 145 208
rect 143 207 144 208
rect 142 207 143 208
rect 141 207 142 208
rect 140 207 141 208
rect 139 207 140 208
rect 138 207 139 208
rect 137 207 138 208
rect 136 207 137 208
rect 135 207 136 208
rect 134 207 135 208
rect 133 207 134 208
rect 132 207 133 208
rect 131 207 132 208
rect 130 207 131 208
rect 129 207 130 208
rect 128 207 129 208
rect 127 207 128 208
rect 126 207 127 208
rect 125 207 126 208
rect 124 207 125 208
rect 123 207 124 208
rect 122 207 123 208
rect 121 207 122 208
rect 120 207 121 208
rect 119 207 120 208
rect 118 207 119 208
rect 117 207 118 208
rect 116 207 117 208
rect 115 207 116 208
rect 114 207 115 208
rect 113 207 114 208
rect 112 207 113 208
rect 111 207 112 208
rect 110 207 111 208
rect 109 207 110 208
rect 108 207 109 208
rect 107 207 108 208
rect 106 207 107 208
rect 105 207 106 208
rect 104 207 105 208
rect 103 207 104 208
rect 102 207 103 208
rect 101 207 102 208
rect 100 207 101 208
rect 99 207 100 208
rect 98 207 99 208
rect 97 207 98 208
rect 96 207 97 208
rect 95 207 96 208
rect 94 207 95 208
rect 93 207 94 208
rect 92 207 93 208
rect 91 207 92 208
rect 90 207 91 208
rect 89 207 90 208
rect 88 207 89 208
rect 87 207 88 208
rect 86 207 87 208
rect 85 207 86 208
rect 84 207 85 208
rect 83 207 84 208
rect 82 207 83 208
rect 81 207 82 208
rect 80 207 81 208
rect 79 207 80 208
rect 78 207 79 208
rect 59 207 60 208
rect 58 207 59 208
rect 57 207 58 208
rect 56 207 57 208
rect 55 207 56 208
rect 54 207 55 208
rect 53 207 54 208
rect 52 207 53 208
rect 51 207 52 208
rect 50 207 51 208
rect 49 207 50 208
rect 48 207 49 208
rect 47 207 48 208
rect 46 207 47 208
rect 45 207 46 208
rect 44 207 45 208
rect 43 207 44 208
rect 42 207 43 208
rect 41 207 42 208
rect 40 207 41 208
rect 39 207 40 208
rect 38 207 39 208
rect 37 207 38 208
rect 36 207 37 208
rect 35 207 36 208
rect 34 207 35 208
rect 33 207 34 208
rect 32 207 33 208
rect 31 207 32 208
rect 30 207 31 208
rect 29 207 30 208
rect 28 207 29 208
rect 27 207 28 208
rect 26 207 27 208
rect 25 207 26 208
rect 24 207 25 208
rect 23 207 24 208
rect 22 207 23 208
rect 21 207 22 208
rect 20 207 21 208
rect 19 207 20 208
rect 18 207 19 208
rect 17 207 18 208
rect 16 207 17 208
rect 15 207 16 208
rect 14 207 15 208
rect 13 207 14 208
rect 12 207 13 208
rect 11 207 12 208
rect 10 207 11 208
rect 426 208 427 209
rect 425 208 426 209
rect 424 208 425 209
rect 423 208 424 209
rect 422 208 423 209
rect 421 208 422 209
rect 420 208 421 209
rect 419 208 420 209
rect 418 208 419 209
rect 417 208 418 209
rect 416 208 417 209
rect 415 208 416 209
rect 414 208 415 209
rect 413 208 414 209
rect 412 208 413 209
rect 411 208 412 209
rect 410 208 411 209
rect 355 208 356 209
rect 354 208 355 209
rect 353 208 354 209
rect 352 208 353 209
rect 351 208 352 209
rect 350 208 351 209
rect 349 208 350 209
rect 348 208 349 209
rect 347 208 348 209
rect 346 208 347 209
rect 345 208 346 209
rect 344 208 345 209
rect 343 208 344 209
rect 342 208 343 209
rect 341 208 342 209
rect 340 208 341 209
rect 339 208 340 209
rect 338 208 339 209
rect 337 208 338 209
rect 336 208 337 209
rect 335 208 336 209
rect 334 208 335 209
rect 333 208 334 209
rect 332 208 333 209
rect 331 208 332 209
rect 330 208 331 209
rect 329 208 330 209
rect 328 208 329 209
rect 327 208 328 209
rect 326 208 327 209
rect 325 208 326 209
rect 324 208 325 209
rect 323 208 324 209
rect 322 208 323 209
rect 321 208 322 209
rect 320 208 321 209
rect 319 208 320 209
rect 318 208 319 209
rect 317 208 318 209
rect 316 208 317 209
rect 315 208 316 209
rect 314 208 315 209
rect 313 208 314 209
rect 312 208 313 209
rect 311 208 312 209
rect 310 208 311 209
rect 309 208 310 209
rect 308 208 309 209
rect 307 208 308 209
rect 306 208 307 209
rect 305 208 306 209
rect 304 208 305 209
rect 303 208 304 209
rect 302 208 303 209
rect 301 208 302 209
rect 300 208 301 209
rect 299 208 300 209
rect 298 208 299 209
rect 297 208 298 209
rect 296 208 297 209
rect 295 208 296 209
rect 294 208 295 209
rect 293 208 294 209
rect 292 208 293 209
rect 291 208 292 209
rect 290 208 291 209
rect 289 208 290 209
rect 288 208 289 209
rect 287 208 288 209
rect 286 208 287 209
rect 285 208 286 209
rect 284 208 285 209
rect 283 208 284 209
rect 282 208 283 209
rect 281 208 282 209
rect 280 208 281 209
rect 279 208 280 209
rect 278 208 279 209
rect 277 208 278 209
rect 276 208 277 209
rect 275 208 276 209
rect 274 208 275 209
rect 273 208 274 209
rect 272 208 273 209
rect 271 208 272 209
rect 270 208 271 209
rect 269 208 270 209
rect 268 208 269 209
rect 267 208 268 209
rect 266 208 267 209
rect 265 208 266 209
rect 264 208 265 209
rect 263 208 264 209
rect 262 208 263 209
rect 261 208 262 209
rect 260 208 261 209
rect 259 208 260 209
rect 258 208 259 209
rect 257 208 258 209
rect 256 208 257 209
rect 255 208 256 209
rect 254 208 255 209
rect 253 208 254 209
rect 252 208 253 209
rect 251 208 252 209
rect 250 208 251 209
rect 249 208 250 209
rect 248 208 249 209
rect 247 208 248 209
rect 246 208 247 209
rect 245 208 246 209
rect 244 208 245 209
rect 243 208 244 209
rect 242 208 243 209
rect 241 208 242 209
rect 240 208 241 209
rect 239 208 240 209
rect 238 208 239 209
rect 237 208 238 209
rect 236 208 237 209
rect 235 208 236 209
rect 234 208 235 209
rect 233 208 234 209
rect 232 208 233 209
rect 231 208 232 209
rect 230 208 231 209
rect 229 208 230 209
rect 228 208 229 209
rect 227 208 228 209
rect 226 208 227 209
rect 225 208 226 209
rect 224 208 225 209
rect 223 208 224 209
rect 222 208 223 209
rect 221 208 222 209
rect 220 208 221 209
rect 219 208 220 209
rect 218 208 219 209
rect 217 208 218 209
rect 216 208 217 209
rect 215 208 216 209
rect 214 208 215 209
rect 213 208 214 209
rect 212 208 213 209
rect 211 208 212 209
rect 210 208 211 209
rect 209 208 210 209
rect 208 208 209 209
rect 207 208 208 209
rect 206 208 207 209
rect 205 208 206 209
rect 204 208 205 209
rect 203 208 204 209
rect 202 208 203 209
rect 201 208 202 209
rect 200 208 201 209
rect 167 208 168 209
rect 166 208 167 209
rect 165 208 166 209
rect 164 208 165 209
rect 163 208 164 209
rect 162 208 163 209
rect 161 208 162 209
rect 160 208 161 209
rect 159 208 160 209
rect 158 208 159 209
rect 157 208 158 209
rect 156 208 157 209
rect 155 208 156 209
rect 154 208 155 209
rect 153 208 154 209
rect 152 208 153 209
rect 151 208 152 209
rect 150 208 151 209
rect 149 208 150 209
rect 148 208 149 209
rect 147 208 148 209
rect 146 208 147 209
rect 145 208 146 209
rect 144 208 145 209
rect 143 208 144 209
rect 142 208 143 209
rect 141 208 142 209
rect 140 208 141 209
rect 139 208 140 209
rect 138 208 139 209
rect 137 208 138 209
rect 136 208 137 209
rect 135 208 136 209
rect 134 208 135 209
rect 133 208 134 209
rect 132 208 133 209
rect 131 208 132 209
rect 130 208 131 209
rect 129 208 130 209
rect 128 208 129 209
rect 127 208 128 209
rect 126 208 127 209
rect 125 208 126 209
rect 124 208 125 209
rect 123 208 124 209
rect 122 208 123 209
rect 121 208 122 209
rect 120 208 121 209
rect 119 208 120 209
rect 118 208 119 209
rect 117 208 118 209
rect 116 208 117 209
rect 115 208 116 209
rect 114 208 115 209
rect 113 208 114 209
rect 112 208 113 209
rect 111 208 112 209
rect 110 208 111 209
rect 109 208 110 209
rect 108 208 109 209
rect 107 208 108 209
rect 106 208 107 209
rect 105 208 106 209
rect 104 208 105 209
rect 103 208 104 209
rect 102 208 103 209
rect 101 208 102 209
rect 100 208 101 209
rect 99 208 100 209
rect 98 208 99 209
rect 97 208 98 209
rect 96 208 97 209
rect 95 208 96 209
rect 94 208 95 209
rect 93 208 94 209
rect 92 208 93 209
rect 91 208 92 209
rect 90 208 91 209
rect 89 208 90 209
rect 88 208 89 209
rect 87 208 88 209
rect 86 208 87 209
rect 85 208 86 209
rect 84 208 85 209
rect 83 208 84 209
rect 82 208 83 209
rect 81 208 82 209
rect 80 208 81 209
rect 79 208 80 209
rect 60 208 61 209
rect 59 208 60 209
rect 58 208 59 209
rect 57 208 58 209
rect 56 208 57 209
rect 55 208 56 209
rect 54 208 55 209
rect 53 208 54 209
rect 52 208 53 209
rect 51 208 52 209
rect 50 208 51 209
rect 49 208 50 209
rect 48 208 49 209
rect 47 208 48 209
rect 46 208 47 209
rect 45 208 46 209
rect 44 208 45 209
rect 43 208 44 209
rect 42 208 43 209
rect 41 208 42 209
rect 40 208 41 209
rect 39 208 40 209
rect 38 208 39 209
rect 37 208 38 209
rect 36 208 37 209
rect 35 208 36 209
rect 34 208 35 209
rect 33 208 34 209
rect 32 208 33 209
rect 31 208 32 209
rect 30 208 31 209
rect 29 208 30 209
rect 28 208 29 209
rect 27 208 28 209
rect 26 208 27 209
rect 25 208 26 209
rect 24 208 25 209
rect 23 208 24 209
rect 22 208 23 209
rect 21 208 22 209
rect 20 208 21 209
rect 19 208 20 209
rect 18 208 19 209
rect 17 208 18 209
rect 16 208 17 209
rect 15 208 16 209
rect 14 208 15 209
rect 13 208 14 209
rect 12 208 13 209
rect 11 208 12 209
rect 10 208 11 209
rect 428 209 429 210
rect 427 209 428 210
rect 426 209 427 210
rect 425 209 426 210
rect 424 209 425 210
rect 423 209 424 210
rect 422 209 423 210
rect 421 209 422 210
rect 420 209 421 210
rect 419 209 420 210
rect 418 209 419 210
rect 417 209 418 210
rect 416 209 417 210
rect 415 209 416 210
rect 414 209 415 210
rect 413 209 414 210
rect 412 209 413 210
rect 411 209 412 210
rect 410 209 411 210
rect 409 209 410 210
rect 408 209 409 210
rect 407 209 408 210
rect 355 209 356 210
rect 354 209 355 210
rect 353 209 354 210
rect 352 209 353 210
rect 351 209 352 210
rect 350 209 351 210
rect 349 209 350 210
rect 348 209 349 210
rect 347 209 348 210
rect 346 209 347 210
rect 345 209 346 210
rect 344 209 345 210
rect 343 209 344 210
rect 342 209 343 210
rect 341 209 342 210
rect 340 209 341 210
rect 339 209 340 210
rect 338 209 339 210
rect 337 209 338 210
rect 336 209 337 210
rect 335 209 336 210
rect 334 209 335 210
rect 333 209 334 210
rect 332 209 333 210
rect 331 209 332 210
rect 330 209 331 210
rect 329 209 330 210
rect 328 209 329 210
rect 327 209 328 210
rect 326 209 327 210
rect 325 209 326 210
rect 324 209 325 210
rect 323 209 324 210
rect 322 209 323 210
rect 321 209 322 210
rect 320 209 321 210
rect 319 209 320 210
rect 318 209 319 210
rect 317 209 318 210
rect 316 209 317 210
rect 315 209 316 210
rect 314 209 315 210
rect 313 209 314 210
rect 312 209 313 210
rect 311 209 312 210
rect 310 209 311 210
rect 309 209 310 210
rect 308 209 309 210
rect 307 209 308 210
rect 306 209 307 210
rect 305 209 306 210
rect 304 209 305 210
rect 303 209 304 210
rect 302 209 303 210
rect 301 209 302 210
rect 300 209 301 210
rect 299 209 300 210
rect 298 209 299 210
rect 297 209 298 210
rect 296 209 297 210
rect 295 209 296 210
rect 294 209 295 210
rect 293 209 294 210
rect 292 209 293 210
rect 291 209 292 210
rect 290 209 291 210
rect 289 209 290 210
rect 288 209 289 210
rect 287 209 288 210
rect 286 209 287 210
rect 285 209 286 210
rect 284 209 285 210
rect 283 209 284 210
rect 282 209 283 210
rect 281 209 282 210
rect 280 209 281 210
rect 279 209 280 210
rect 278 209 279 210
rect 277 209 278 210
rect 276 209 277 210
rect 275 209 276 210
rect 274 209 275 210
rect 273 209 274 210
rect 272 209 273 210
rect 271 209 272 210
rect 270 209 271 210
rect 269 209 270 210
rect 268 209 269 210
rect 267 209 268 210
rect 266 209 267 210
rect 265 209 266 210
rect 264 209 265 210
rect 263 209 264 210
rect 262 209 263 210
rect 261 209 262 210
rect 260 209 261 210
rect 259 209 260 210
rect 258 209 259 210
rect 257 209 258 210
rect 256 209 257 210
rect 255 209 256 210
rect 254 209 255 210
rect 253 209 254 210
rect 252 209 253 210
rect 251 209 252 210
rect 250 209 251 210
rect 249 209 250 210
rect 248 209 249 210
rect 247 209 248 210
rect 246 209 247 210
rect 245 209 246 210
rect 244 209 245 210
rect 243 209 244 210
rect 242 209 243 210
rect 241 209 242 210
rect 240 209 241 210
rect 239 209 240 210
rect 238 209 239 210
rect 237 209 238 210
rect 236 209 237 210
rect 235 209 236 210
rect 234 209 235 210
rect 233 209 234 210
rect 232 209 233 210
rect 231 209 232 210
rect 230 209 231 210
rect 229 209 230 210
rect 228 209 229 210
rect 227 209 228 210
rect 226 209 227 210
rect 225 209 226 210
rect 224 209 225 210
rect 223 209 224 210
rect 222 209 223 210
rect 221 209 222 210
rect 220 209 221 210
rect 219 209 220 210
rect 218 209 219 210
rect 217 209 218 210
rect 216 209 217 210
rect 215 209 216 210
rect 214 209 215 210
rect 213 209 214 210
rect 212 209 213 210
rect 211 209 212 210
rect 210 209 211 210
rect 209 209 210 210
rect 208 209 209 210
rect 207 209 208 210
rect 206 209 207 210
rect 205 209 206 210
rect 204 209 205 210
rect 203 209 204 210
rect 202 209 203 210
rect 201 209 202 210
rect 200 209 201 210
rect 199 209 200 210
rect 165 209 166 210
rect 164 209 165 210
rect 163 209 164 210
rect 162 209 163 210
rect 161 209 162 210
rect 160 209 161 210
rect 159 209 160 210
rect 158 209 159 210
rect 157 209 158 210
rect 156 209 157 210
rect 155 209 156 210
rect 154 209 155 210
rect 153 209 154 210
rect 152 209 153 210
rect 151 209 152 210
rect 150 209 151 210
rect 149 209 150 210
rect 148 209 149 210
rect 147 209 148 210
rect 146 209 147 210
rect 145 209 146 210
rect 144 209 145 210
rect 143 209 144 210
rect 142 209 143 210
rect 141 209 142 210
rect 140 209 141 210
rect 139 209 140 210
rect 138 209 139 210
rect 137 209 138 210
rect 136 209 137 210
rect 135 209 136 210
rect 134 209 135 210
rect 133 209 134 210
rect 132 209 133 210
rect 131 209 132 210
rect 130 209 131 210
rect 129 209 130 210
rect 128 209 129 210
rect 127 209 128 210
rect 126 209 127 210
rect 125 209 126 210
rect 124 209 125 210
rect 123 209 124 210
rect 122 209 123 210
rect 121 209 122 210
rect 120 209 121 210
rect 119 209 120 210
rect 118 209 119 210
rect 117 209 118 210
rect 116 209 117 210
rect 115 209 116 210
rect 114 209 115 210
rect 113 209 114 210
rect 112 209 113 210
rect 111 209 112 210
rect 110 209 111 210
rect 109 209 110 210
rect 108 209 109 210
rect 107 209 108 210
rect 106 209 107 210
rect 105 209 106 210
rect 104 209 105 210
rect 103 209 104 210
rect 102 209 103 210
rect 101 209 102 210
rect 100 209 101 210
rect 99 209 100 210
rect 98 209 99 210
rect 97 209 98 210
rect 96 209 97 210
rect 95 209 96 210
rect 94 209 95 210
rect 93 209 94 210
rect 92 209 93 210
rect 91 209 92 210
rect 90 209 91 210
rect 89 209 90 210
rect 88 209 89 210
rect 87 209 88 210
rect 86 209 87 210
rect 85 209 86 210
rect 84 209 85 210
rect 83 209 84 210
rect 82 209 83 210
rect 81 209 82 210
rect 61 209 62 210
rect 60 209 61 210
rect 59 209 60 210
rect 58 209 59 210
rect 57 209 58 210
rect 56 209 57 210
rect 55 209 56 210
rect 54 209 55 210
rect 53 209 54 210
rect 52 209 53 210
rect 51 209 52 210
rect 50 209 51 210
rect 49 209 50 210
rect 48 209 49 210
rect 47 209 48 210
rect 46 209 47 210
rect 45 209 46 210
rect 44 209 45 210
rect 43 209 44 210
rect 42 209 43 210
rect 41 209 42 210
rect 40 209 41 210
rect 39 209 40 210
rect 38 209 39 210
rect 37 209 38 210
rect 36 209 37 210
rect 35 209 36 210
rect 34 209 35 210
rect 33 209 34 210
rect 32 209 33 210
rect 31 209 32 210
rect 30 209 31 210
rect 29 209 30 210
rect 28 209 29 210
rect 27 209 28 210
rect 26 209 27 210
rect 25 209 26 210
rect 24 209 25 210
rect 23 209 24 210
rect 22 209 23 210
rect 21 209 22 210
rect 20 209 21 210
rect 19 209 20 210
rect 18 209 19 210
rect 17 209 18 210
rect 16 209 17 210
rect 15 209 16 210
rect 14 209 15 210
rect 13 209 14 210
rect 12 209 13 210
rect 11 209 12 210
rect 10 209 11 210
rect 9 209 10 210
rect 430 210 431 211
rect 429 210 430 211
rect 428 210 429 211
rect 427 210 428 211
rect 426 210 427 211
rect 425 210 426 211
rect 424 210 425 211
rect 423 210 424 211
rect 422 210 423 211
rect 421 210 422 211
rect 420 210 421 211
rect 419 210 420 211
rect 418 210 419 211
rect 417 210 418 211
rect 416 210 417 211
rect 415 210 416 211
rect 414 210 415 211
rect 413 210 414 211
rect 412 210 413 211
rect 411 210 412 211
rect 410 210 411 211
rect 409 210 410 211
rect 408 210 409 211
rect 407 210 408 211
rect 406 210 407 211
rect 405 210 406 211
rect 356 210 357 211
rect 355 210 356 211
rect 354 210 355 211
rect 353 210 354 211
rect 352 210 353 211
rect 351 210 352 211
rect 350 210 351 211
rect 349 210 350 211
rect 348 210 349 211
rect 347 210 348 211
rect 346 210 347 211
rect 345 210 346 211
rect 344 210 345 211
rect 343 210 344 211
rect 342 210 343 211
rect 341 210 342 211
rect 340 210 341 211
rect 339 210 340 211
rect 338 210 339 211
rect 337 210 338 211
rect 336 210 337 211
rect 335 210 336 211
rect 334 210 335 211
rect 333 210 334 211
rect 332 210 333 211
rect 331 210 332 211
rect 330 210 331 211
rect 329 210 330 211
rect 328 210 329 211
rect 327 210 328 211
rect 326 210 327 211
rect 325 210 326 211
rect 324 210 325 211
rect 323 210 324 211
rect 322 210 323 211
rect 321 210 322 211
rect 320 210 321 211
rect 319 210 320 211
rect 318 210 319 211
rect 317 210 318 211
rect 316 210 317 211
rect 315 210 316 211
rect 314 210 315 211
rect 313 210 314 211
rect 312 210 313 211
rect 311 210 312 211
rect 310 210 311 211
rect 309 210 310 211
rect 308 210 309 211
rect 307 210 308 211
rect 306 210 307 211
rect 305 210 306 211
rect 304 210 305 211
rect 303 210 304 211
rect 302 210 303 211
rect 301 210 302 211
rect 300 210 301 211
rect 299 210 300 211
rect 298 210 299 211
rect 297 210 298 211
rect 296 210 297 211
rect 295 210 296 211
rect 294 210 295 211
rect 293 210 294 211
rect 292 210 293 211
rect 291 210 292 211
rect 290 210 291 211
rect 289 210 290 211
rect 288 210 289 211
rect 287 210 288 211
rect 286 210 287 211
rect 285 210 286 211
rect 284 210 285 211
rect 283 210 284 211
rect 282 210 283 211
rect 281 210 282 211
rect 280 210 281 211
rect 279 210 280 211
rect 278 210 279 211
rect 277 210 278 211
rect 276 210 277 211
rect 275 210 276 211
rect 274 210 275 211
rect 273 210 274 211
rect 272 210 273 211
rect 271 210 272 211
rect 270 210 271 211
rect 269 210 270 211
rect 268 210 269 211
rect 267 210 268 211
rect 266 210 267 211
rect 265 210 266 211
rect 264 210 265 211
rect 263 210 264 211
rect 262 210 263 211
rect 261 210 262 211
rect 260 210 261 211
rect 259 210 260 211
rect 258 210 259 211
rect 257 210 258 211
rect 256 210 257 211
rect 255 210 256 211
rect 254 210 255 211
rect 253 210 254 211
rect 252 210 253 211
rect 251 210 252 211
rect 250 210 251 211
rect 249 210 250 211
rect 248 210 249 211
rect 247 210 248 211
rect 246 210 247 211
rect 245 210 246 211
rect 244 210 245 211
rect 243 210 244 211
rect 242 210 243 211
rect 241 210 242 211
rect 240 210 241 211
rect 239 210 240 211
rect 238 210 239 211
rect 237 210 238 211
rect 236 210 237 211
rect 235 210 236 211
rect 234 210 235 211
rect 233 210 234 211
rect 232 210 233 211
rect 231 210 232 211
rect 230 210 231 211
rect 229 210 230 211
rect 228 210 229 211
rect 227 210 228 211
rect 226 210 227 211
rect 225 210 226 211
rect 224 210 225 211
rect 223 210 224 211
rect 222 210 223 211
rect 221 210 222 211
rect 220 210 221 211
rect 219 210 220 211
rect 218 210 219 211
rect 217 210 218 211
rect 216 210 217 211
rect 215 210 216 211
rect 214 210 215 211
rect 213 210 214 211
rect 212 210 213 211
rect 211 210 212 211
rect 210 210 211 211
rect 209 210 210 211
rect 208 210 209 211
rect 207 210 208 211
rect 206 210 207 211
rect 205 210 206 211
rect 204 210 205 211
rect 203 210 204 211
rect 202 210 203 211
rect 201 210 202 211
rect 200 210 201 211
rect 199 210 200 211
rect 198 210 199 211
rect 162 210 163 211
rect 161 210 162 211
rect 160 210 161 211
rect 159 210 160 211
rect 158 210 159 211
rect 157 210 158 211
rect 156 210 157 211
rect 155 210 156 211
rect 154 210 155 211
rect 153 210 154 211
rect 152 210 153 211
rect 151 210 152 211
rect 150 210 151 211
rect 149 210 150 211
rect 148 210 149 211
rect 147 210 148 211
rect 146 210 147 211
rect 145 210 146 211
rect 144 210 145 211
rect 143 210 144 211
rect 142 210 143 211
rect 141 210 142 211
rect 140 210 141 211
rect 139 210 140 211
rect 138 210 139 211
rect 137 210 138 211
rect 136 210 137 211
rect 135 210 136 211
rect 134 210 135 211
rect 133 210 134 211
rect 132 210 133 211
rect 131 210 132 211
rect 130 210 131 211
rect 129 210 130 211
rect 128 210 129 211
rect 127 210 128 211
rect 126 210 127 211
rect 125 210 126 211
rect 124 210 125 211
rect 123 210 124 211
rect 122 210 123 211
rect 121 210 122 211
rect 120 210 121 211
rect 119 210 120 211
rect 118 210 119 211
rect 117 210 118 211
rect 116 210 117 211
rect 115 210 116 211
rect 114 210 115 211
rect 113 210 114 211
rect 112 210 113 211
rect 111 210 112 211
rect 110 210 111 211
rect 109 210 110 211
rect 108 210 109 211
rect 107 210 108 211
rect 106 210 107 211
rect 105 210 106 211
rect 104 210 105 211
rect 103 210 104 211
rect 102 210 103 211
rect 101 210 102 211
rect 100 210 101 211
rect 99 210 100 211
rect 98 210 99 211
rect 97 210 98 211
rect 96 210 97 211
rect 95 210 96 211
rect 94 210 95 211
rect 93 210 94 211
rect 92 210 93 211
rect 91 210 92 211
rect 90 210 91 211
rect 89 210 90 211
rect 88 210 89 211
rect 87 210 88 211
rect 86 210 87 211
rect 85 210 86 211
rect 84 210 85 211
rect 83 210 84 211
rect 82 210 83 211
rect 61 210 62 211
rect 60 210 61 211
rect 59 210 60 211
rect 58 210 59 211
rect 57 210 58 211
rect 56 210 57 211
rect 55 210 56 211
rect 54 210 55 211
rect 53 210 54 211
rect 52 210 53 211
rect 51 210 52 211
rect 50 210 51 211
rect 49 210 50 211
rect 48 210 49 211
rect 47 210 48 211
rect 46 210 47 211
rect 45 210 46 211
rect 44 210 45 211
rect 43 210 44 211
rect 42 210 43 211
rect 41 210 42 211
rect 40 210 41 211
rect 39 210 40 211
rect 38 210 39 211
rect 37 210 38 211
rect 36 210 37 211
rect 35 210 36 211
rect 34 210 35 211
rect 33 210 34 211
rect 32 210 33 211
rect 31 210 32 211
rect 30 210 31 211
rect 29 210 30 211
rect 28 210 29 211
rect 27 210 28 211
rect 26 210 27 211
rect 25 210 26 211
rect 24 210 25 211
rect 23 210 24 211
rect 22 210 23 211
rect 21 210 22 211
rect 20 210 21 211
rect 19 210 20 211
rect 18 210 19 211
rect 17 210 18 211
rect 16 210 17 211
rect 15 210 16 211
rect 14 210 15 211
rect 13 210 14 211
rect 12 210 13 211
rect 11 210 12 211
rect 10 210 11 211
rect 9 210 10 211
rect 431 211 432 212
rect 430 211 431 212
rect 429 211 430 212
rect 428 211 429 212
rect 427 211 428 212
rect 426 211 427 212
rect 425 211 426 212
rect 424 211 425 212
rect 423 211 424 212
rect 422 211 423 212
rect 421 211 422 212
rect 420 211 421 212
rect 419 211 420 212
rect 418 211 419 212
rect 417 211 418 212
rect 416 211 417 212
rect 415 211 416 212
rect 414 211 415 212
rect 413 211 414 212
rect 412 211 413 212
rect 411 211 412 212
rect 410 211 411 212
rect 409 211 410 212
rect 408 211 409 212
rect 407 211 408 212
rect 406 211 407 212
rect 405 211 406 212
rect 404 211 405 212
rect 356 211 357 212
rect 355 211 356 212
rect 354 211 355 212
rect 353 211 354 212
rect 352 211 353 212
rect 351 211 352 212
rect 350 211 351 212
rect 349 211 350 212
rect 348 211 349 212
rect 347 211 348 212
rect 346 211 347 212
rect 345 211 346 212
rect 344 211 345 212
rect 343 211 344 212
rect 342 211 343 212
rect 341 211 342 212
rect 340 211 341 212
rect 339 211 340 212
rect 338 211 339 212
rect 337 211 338 212
rect 336 211 337 212
rect 335 211 336 212
rect 334 211 335 212
rect 333 211 334 212
rect 332 211 333 212
rect 331 211 332 212
rect 330 211 331 212
rect 329 211 330 212
rect 328 211 329 212
rect 327 211 328 212
rect 326 211 327 212
rect 325 211 326 212
rect 324 211 325 212
rect 323 211 324 212
rect 322 211 323 212
rect 321 211 322 212
rect 320 211 321 212
rect 319 211 320 212
rect 318 211 319 212
rect 317 211 318 212
rect 316 211 317 212
rect 315 211 316 212
rect 314 211 315 212
rect 313 211 314 212
rect 312 211 313 212
rect 311 211 312 212
rect 310 211 311 212
rect 309 211 310 212
rect 308 211 309 212
rect 307 211 308 212
rect 306 211 307 212
rect 305 211 306 212
rect 304 211 305 212
rect 303 211 304 212
rect 302 211 303 212
rect 301 211 302 212
rect 300 211 301 212
rect 299 211 300 212
rect 298 211 299 212
rect 297 211 298 212
rect 296 211 297 212
rect 295 211 296 212
rect 294 211 295 212
rect 293 211 294 212
rect 292 211 293 212
rect 291 211 292 212
rect 290 211 291 212
rect 289 211 290 212
rect 288 211 289 212
rect 287 211 288 212
rect 286 211 287 212
rect 285 211 286 212
rect 284 211 285 212
rect 283 211 284 212
rect 282 211 283 212
rect 281 211 282 212
rect 280 211 281 212
rect 279 211 280 212
rect 278 211 279 212
rect 277 211 278 212
rect 276 211 277 212
rect 275 211 276 212
rect 274 211 275 212
rect 273 211 274 212
rect 272 211 273 212
rect 271 211 272 212
rect 270 211 271 212
rect 269 211 270 212
rect 268 211 269 212
rect 267 211 268 212
rect 266 211 267 212
rect 265 211 266 212
rect 264 211 265 212
rect 263 211 264 212
rect 262 211 263 212
rect 261 211 262 212
rect 260 211 261 212
rect 259 211 260 212
rect 258 211 259 212
rect 257 211 258 212
rect 256 211 257 212
rect 255 211 256 212
rect 254 211 255 212
rect 253 211 254 212
rect 252 211 253 212
rect 251 211 252 212
rect 250 211 251 212
rect 249 211 250 212
rect 248 211 249 212
rect 247 211 248 212
rect 246 211 247 212
rect 245 211 246 212
rect 244 211 245 212
rect 243 211 244 212
rect 242 211 243 212
rect 241 211 242 212
rect 240 211 241 212
rect 239 211 240 212
rect 238 211 239 212
rect 237 211 238 212
rect 236 211 237 212
rect 235 211 236 212
rect 234 211 235 212
rect 233 211 234 212
rect 232 211 233 212
rect 231 211 232 212
rect 230 211 231 212
rect 229 211 230 212
rect 228 211 229 212
rect 227 211 228 212
rect 226 211 227 212
rect 225 211 226 212
rect 224 211 225 212
rect 223 211 224 212
rect 222 211 223 212
rect 221 211 222 212
rect 220 211 221 212
rect 219 211 220 212
rect 218 211 219 212
rect 217 211 218 212
rect 216 211 217 212
rect 215 211 216 212
rect 214 211 215 212
rect 213 211 214 212
rect 212 211 213 212
rect 211 211 212 212
rect 210 211 211 212
rect 209 211 210 212
rect 208 211 209 212
rect 207 211 208 212
rect 206 211 207 212
rect 205 211 206 212
rect 204 211 205 212
rect 203 211 204 212
rect 202 211 203 212
rect 201 211 202 212
rect 200 211 201 212
rect 199 211 200 212
rect 198 211 199 212
rect 197 211 198 212
rect 196 211 197 212
rect 159 211 160 212
rect 158 211 159 212
rect 157 211 158 212
rect 156 211 157 212
rect 155 211 156 212
rect 154 211 155 212
rect 153 211 154 212
rect 152 211 153 212
rect 151 211 152 212
rect 150 211 151 212
rect 149 211 150 212
rect 148 211 149 212
rect 147 211 148 212
rect 146 211 147 212
rect 145 211 146 212
rect 144 211 145 212
rect 143 211 144 212
rect 142 211 143 212
rect 141 211 142 212
rect 140 211 141 212
rect 139 211 140 212
rect 138 211 139 212
rect 137 211 138 212
rect 136 211 137 212
rect 135 211 136 212
rect 134 211 135 212
rect 133 211 134 212
rect 132 211 133 212
rect 131 211 132 212
rect 130 211 131 212
rect 129 211 130 212
rect 128 211 129 212
rect 127 211 128 212
rect 126 211 127 212
rect 125 211 126 212
rect 124 211 125 212
rect 123 211 124 212
rect 122 211 123 212
rect 121 211 122 212
rect 120 211 121 212
rect 119 211 120 212
rect 118 211 119 212
rect 117 211 118 212
rect 116 211 117 212
rect 115 211 116 212
rect 114 211 115 212
rect 113 211 114 212
rect 112 211 113 212
rect 111 211 112 212
rect 110 211 111 212
rect 109 211 110 212
rect 108 211 109 212
rect 107 211 108 212
rect 106 211 107 212
rect 105 211 106 212
rect 104 211 105 212
rect 103 211 104 212
rect 102 211 103 212
rect 101 211 102 212
rect 100 211 101 212
rect 99 211 100 212
rect 98 211 99 212
rect 97 211 98 212
rect 96 211 97 212
rect 95 211 96 212
rect 94 211 95 212
rect 93 211 94 212
rect 92 211 93 212
rect 91 211 92 212
rect 90 211 91 212
rect 89 211 90 212
rect 88 211 89 212
rect 87 211 88 212
rect 86 211 87 212
rect 85 211 86 212
rect 84 211 85 212
rect 62 211 63 212
rect 61 211 62 212
rect 60 211 61 212
rect 59 211 60 212
rect 58 211 59 212
rect 57 211 58 212
rect 56 211 57 212
rect 55 211 56 212
rect 54 211 55 212
rect 53 211 54 212
rect 52 211 53 212
rect 51 211 52 212
rect 50 211 51 212
rect 49 211 50 212
rect 48 211 49 212
rect 47 211 48 212
rect 46 211 47 212
rect 45 211 46 212
rect 44 211 45 212
rect 43 211 44 212
rect 42 211 43 212
rect 41 211 42 212
rect 40 211 41 212
rect 39 211 40 212
rect 38 211 39 212
rect 37 211 38 212
rect 36 211 37 212
rect 35 211 36 212
rect 34 211 35 212
rect 33 211 34 212
rect 32 211 33 212
rect 31 211 32 212
rect 30 211 31 212
rect 29 211 30 212
rect 28 211 29 212
rect 27 211 28 212
rect 26 211 27 212
rect 25 211 26 212
rect 24 211 25 212
rect 23 211 24 212
rect 22 211 23 212
rect 21 211 22 212
rect 20 211 21 212
rect 19 211 20 212
rect 18 211 19 212
rect 17 211 18 212
rect 16 211 17 212
rect 15 211 16 212
rect 14 211 15 212
rect 13 211 14 212
rect 12 211 13 212
rect 11 211 12 212
rect 10 211 11 212
rect 9 211 10 212
rect 432 212 433 213
rect 431 212 432 213
rect 430 212 431 213
rect 429 212 430 213
rect 428 212 429 213
rect 427 212 428 213
rect 426 212 427 213
rect 425 212 426 213
rect 424 212 425 213
rect 423 212 424 213
rect 422 212 423 213
rect 421 212 422 213
rect 420 212 421 213
rect 419 212 420 213
rect 418 212 419 213
rect 417 212 418 213
rect 416 212 417 213
rect 415 212 416 213
rect 414 212 415 213
rect 413 212 414 213
rect 412 212 413 213
rect 411 212 412 213
rect 410 212 411 213
rect 409 212 410 213
rect 408 212 409 213
rect 407 212 408 213
rect 406 212 407 213
rect 405 212 406 213
rect 404 212 405 213
rect 403 212 404 213
rect 357 212 358 213
rect 356 212 357 213
rect 355 212 356 213
rect 354 212 355 213
rect 353 212 354 213
rect 352 212 353 213
rect 351 212 352 213
rect 350 212 351 213
rect 349 212 350 213
rect 348 212 349 213
rect 347 212 348 213
rect 346 212 347 213
rect 345 212 346 213
rect 344 212 345 213
rect 343 212 344 213
rect 342 212 343 213
rect 341 212 342 213
rect 340 212 341 213
rect 339 212 340 213
rect 338 212 339 213
rect 337 212 338 213
rect 336 212 337 213
rect 335 212 336 213
rect 334 212 335 213
rect 333 212 334 213
rect 332 212 333 213
rect 331 212 332 213
rect 330 212 331 213
rect 329 212 330 213
rect 328 212 329 213
rect 327 212 328 213
rect 326 212 327 213
rect 325 212 326 213
rect 324 212 325 213
rect 323 212 324 213
rect 322 212 323 213
rect 321 212 322 213
rect 320 212 321 213
rect 319 212 320 213
rect 318 212 319 213
rect 317 212 318 213
rect 316 212 317 213
rect 315 212 316 213
rect 314 212 315 213
rect 313 212 314 213
rect 312 212 313 213
rect 311 212 312 213
rect 310 212 311 213
rect 309 212 310 213
rect 308 212 309 213
rect 307 212 308 213
rect 306 212 307 213
rect 305 212 306 213
rect 304 212 305 213
rect 303 212 304 213
rect 302 212 303 213
rect 301 212 302 213
rect 300 212 301 213
rect 299 212 300 213
rect 298 212 299 213
rect 297 212 298 213
rect 296 212 297 213
rect 295 212 296 213
rect 294 212 295 213
rect 293 212 294 213
rect 292 212 293 213
rect 291 212 292 213
rect 290 212 291 213
rect 289 212 290 213
rect 288 212 289 213
rect 287 212 288 213
rect 286 212 287 213
rect 285 212 286 213
rect 284 212 285 213
rect 283 212 284 213
rect 282 212 283 213
rect 281 212 282 213
rect 280 212 281 213
rect 279 212 280 213
rect 278 212 279 213
rect 277 212 278 213
rect 276 212 277 213
rect 275 212 276 213
rect 274 212 275 213
rect 273 212 274 213
rect 272 212 273 213
rect 271 212 272 213
rect 270 212 271 213
rect 269 212 270 213
rect 268 212 269 213
rect 267 212 268 213
rect 266 212 267 213
rect 265 212 266 213
rect 264 212 265 213
rect 263 212 264 213
rect 262 212 263 213
rect 261 212 262 213
rect 260 212 261 213
rect 259 212 260 213
rect 258 212 259 213
rect 257 212 258 213
rect 256 212 257 213
rect 255 212 256 213
rect 254 212 255 213
rect 253 212 254 213
rect 252 212 253 213
rect 251 212 252 213
rect 250 212 251 213
rect 249 212 250 213
rect 248 212 249 213
rect 247 212 248 213
rect 246 212 247 213
rect 245 212 246 213
rect 244 212 245 213
rect 243 212 244 213
rect 242 212 243 213
rect 241 212 242 213
rect 240 212 241 213
rect 239 212 240 213
rect 238 212 239 213
rect 237 212 238 213
rect 236 212 237 213
rect 235 212 236 213
rect 234 212 235 213
rect 233 212 234 213
rect 232 212 233 213
rect 231 212 232 213
rect 230 212 231 213
rect 229 212 230 213
rect 228 212 229 213
rect 227 212 228 213
rect 226 212 227 213
rect 225 212 226 213
rect 224 212 225 213
rect 223 212 224 213
rect 222 212 223 213
rect 221 212 222 213
rect 220 212 221 213
rect 219 212 220 213
rect 218 212 219 213
rect 217 212 218 213
rect 216 212 217 213
rect 215 212 216 213
rect 214 212 215 213
rect 213 212 214 213
rect 212 212 213 213
rect 211 212 212 213
rect 210 212 211 213
rect 209 212 210 213
rect 208 212 209 213
rect 207 212 208 213
rect 206 212 207 213
rect 205 212 206 213
rect 204 212 205 213
rect 203 212 204 213
rect 202 212 203 213
rect 201 212 202 213
rect 200 212 201 213
rect 199 212 200 213
rect 198 212 199 213
rect 197 212 198 213
rect 196 212 197 213
rect 195 212 196 213
rect 156 212 157 213
rect 155 212 156 213
rect 154 212 155 213
rect 153 212 154 213
rect 152 212 153 213
rect 151 212 152 213
rect 150 212 151 213
rect 149 212 150 213
rect 148 212 149 213
rect 147 212 148 213
rect 146 212 147 213
rect 145 212 146 213
rect 144 212 145 213
rect 143 212 144 213
rect 142 212 143 213
rect 141 212 142 213
rect 140 212 141 213
rect 139 212 140 213
rect 138 212 139 213
rect 137 212 138 213
rect 136 212 137 213
rect 135 212 136 213
rect 134 212 135 213
rect 133 212 134 213
rect 132 212 133 213
rect 131 212 132 213
rect 130 212 131 213
rect 129 212 130 213
rect 128 212 129 213
rect 127 212 128 213
rect 126 212 127 213
rect 125 212 126 213
rect 124 212 125 213
rect 123 212 124 213
rect 122 212 123 213
rect 121 212 122 213
rect 120 212 121 213
rect 119 212 120 213
rect 118 212 119 213
rect 117 212 118 213
rect 116 212 117 213
rect 115 212 116 213
rect 114 212 115 213
rect 113 212 114 213
rect 112 212 113 213
rect 111 212 112 213
rect 110 212 111 213
rect 109 212 110 213
rect 108 212 109 213
rect 107 212 108 213
rect 106 212 107 213
rect 105 212 106 213
rect 104 212 105 213
rect 103 212 104 213
rect 102 212 103 213
rect 101 212 102 213
rect 100 212 101 213
rect 99 212 100 213
rect 98 212 99 213
rect 97 212 98 213
rect 96 212 97 213
rect 95 212 96 213
rect 94 212 95 213
rect 93 212 94 213
rect 92 212 93 213
rect 91 212 92 213
rect 90 212 91 213
rect 89 212 90 213
rect 88 212 89 213
rect 87 212 88 213
rect 86 212 87 213
rect 63 212 64 213
rect 62 212 63 213
rect 61 212 62 213
rect 60 212 61 213
rect 59 212 60 213
rect 58 212 59 213
rect 57 212 58 213
rect 56 212 57 213
rect 55 212 56 213
rect 54 212 55 213
rect 53 212 54 213
rect 52 212 53 213
rect 51 212 52 213
rect 50 212 51 213
rect 49 212 50 213
rect 48 212 49 213
rect 47 212 48 213
rect 46 212 47 213
rect 45 212 46 213
rect 44 212 45 213
rect 43 212 44 213
rect 42 212 43 213
rect 41 212 42 213
rect 40 212 41 213
rect 39 212 40 213
rect 38 212 39 213
rect 37 212 38 213
rect 36 212 37 213
rect 35 212 36 213
rect 34 212 35 213
rect 33 212 34 213
rect 32 212 33 213
rect 31 212 32 213
rect 30 212 31 213
rect 29 212 30 213
rect 28 212 29 213
rect 27 212 28 213
rect 26 212 27 213
rect 25 212 26 213
rect 24 212 25 213
rect 23 212 24 213
rect 22 212 23 213
rect 21 212 22 213
rect 20 212 21 213
rect 19 212 20 213
rect 18 212 19 213
rect 17 212 18 213
rect 16 212 17 213
rect 15 212 16 213
rect 14 212 15 213
rect 13 212 14 213
rect 12 212 13 213
rect 11 212 12 213
rect 10 212 11 213
rect 9 212 10 213
rect 433 213 434 214
rect 432 213 433 214
rect 431 213 432 214
rect 430 213 431 214
rect 429 213 430 214
rect 428 213 429 214
rect 427 213 428 214
rect 426 213 427 214
rect 425 213 426 214
rect 424 213 425 214
rect 423 213 424 214
rect 422 213 423 214
rect 421 213 422 214
rect 420 213 421 214
rect 419 213 420 214
rect 418 213 419 214
rect 417 213 418 214
rect 416 213 417 214
rect 415 213 416 214
rect 414 213 415 214
rect 413 213 414 214
rect 412 213 413 214
rect 411 213 412 214
rect 410 213 411 214
rect 409 213 410 214
rect 408 213 409 214
rect 407 213 408 214
rect 406 213 407 214
rect 405 213 406 214
rect 404 213 405 214
rect 403 213 404 214
rect 402 213 403 214
rect 358 213 359 214
rect 357 213 358 214
rect 356 213 357 214
rect 355 213 356 214
rect 354 213 355 214
rect 353 213 354 214
rect 352 213 353 214
rect 351 213 352 214
rect 350 213 351 214
rect 349 213 350 214
rect 348 213 349 214
rect 347 213 348 214
rect 346 213 347 214
rect 345 213 346 214
rect 344 213 345 214
rect 343 213 344 214
rect 342 213 343 214
rect 341 213 342 214
rect 340 213 341 214
rect 339 213 340 214
rect 338 213 339 214
rect 337 213 338 214
rect 336 213 337 214
rect 335 213 336 214
rect 334 213 335 214
rect 333 213 334 214
rect 332 213 333 214
rect 331 213 332 214
rect 330 213 331 214
rect 329 213 330 214
rect 328 213 329 214
rect 327 213 328 214
rect 326 213 327 214
rect 325 213 326 214
rect 324 213 325 214
rect 323 213 324 214
rect 322 213 323 214
rect 321 213 322 214
rect 320 213 321 214
rect 319 213 320 214
rect 318 213 319 214
rect 317 213 318 214
rect 316 213 317 214
rect 315 213 316 214
rect 314 213 315 214
rect 313 213 314 214
rect 312 213 313 214
rect 311 213 312 214
rect 310 213 311 214
rect 309 213 310 214
rect 308 213 309 214
rect 307 213 308 214
rect 306 213 307 214
rect 305 213 306 214
rect 304 213 305 214
rect 303 213 304 214
rect 302 213 303 214
rect 301 213 302 214
rect 300 213 301 214
rect 299 213 300 214
rect 298 213 299 214
rect 297 213 298 214
rect 296 213 297 214
rect 295 213 296 214
rect 294 213 295 214
rect 293 213 294 214
rect 292 213 293 214
rect 291 213 292 214
rect 290 213 291 214
rect 289 213 290 214
rect 288 213 289 214
rect 287 213 288 214
rect 286 213 287 214
rect 285 213 286 214
rect 284 213 285 214
rect 283 213 284 214
rect 282 213 283 214
rect 281 213 282 214
rect 280 213 281 214
rect 279 213 280 214
rect 278 213 279 214
rect 277 213 278 214
rect 276 213 277 214
rect 275 213 276 214
rect 274 213 275 214
rect 273 213 274 214
rect 272 213 273 214
rect 271 213 272 214
rect 270 213 271 214
rect 269 213 270 214
rect 268 213 269 214
rect 267 213 268 214
rect 266 213 267 214
rect 265 213 266 214
rect 264 213 265 214
rect 263 213 264 214
rect 262 213 263 214
rect 261 213 262 214
rect 260 213 261 214
rect 259 213 260 214
rect 258 213 259 214
rect 257 213 258 214
rect 256 213 257 214
rect 255 213 256 214
rect 254 213 255 214
rect 253 213 254 214
rect 252 213 253 214
rect 251 213 252 214
rect 250 213 251 214
rect 249 213 250 214
rect 248 213 249 214
rect 247 213 248 214
rect 246 213 247 214
rect 245 213 246 214
rect 244 213 245 214
rect 243 213 244 214
rect 242 213 243 214
rect 241 213 242 214
rect 240 213 241 214
rect 239 213 240 214
rect 238 213 239 214
rect 237 213 238 214
rect 236 213 237 214
rect 235 213 236 214
rect 234 213 235 214
rect 233 213 234 214
rect 232 213 233 214
rect 231 213 232 214
rect 230 213 231 214
rect 229 213 230 214
rect 228 213 229 214
rect 227 213 228 214
rect 226 213 227 214
rect 225 213 226 214
rect 224 213 225 214
rect 223 213 224 214
rect 222 213 223 214
rect 221 213 222 214
rect 220 213 221 214
rect 219 213 220 214
rect 218 213 219 214
rect 217 213 218 214
rect 216 213 217 214
rect 215 213 216 214
rect 214 213 215 214
rect 213 213 214 214
rect 212 213 213 214
rect 211 213 212 214
rect 210 213 211 214
rect 209 213 210 214
rect 208 213 209 214
rect 207 213 208 214
rect 206 213 207 214
rect 205 213 206 214
rect 204 213 205 214
rect 203 213 204 214
rect 202 213 203 214
rect 201 213 202 214
rect 200 213 201 214
rect 199 213 200 214
rect 198 213 199 214
rect 197 213 198 214
rect 196 213 197 214
rect 195 213 196 214
rect 194 213 195 214
rect 193 213 194 214
rect 153 213 154 214
rect 152 213 153 214
rect 151 213 152 214
rect 150 213 151 214
rect 149 213 150 214
rect 148 213 149 214
rect 147 213 148 214
rect 146 213 147 214
rect 145 213 146 214
rect 144 213 145 214
rect 143 213 144 214
rect 142 213 143 214
rect 141 213 142 214
rect 140 213 141 214
rect 139 213 140 214
rect 138 213 139 214
rect 137 213 138 214
rect 136 213 137 214
rect 135 213 136 214
rect 134 213 135 214
rect 133 213 134 214
rect 132 213 133 214
rect 131 213 132 214
rect 130 213 131 214
rect 129 213 130 214
rect 128 213 129 214
rect 127 213 128 214
rect 126 213 127 214
rect 125 213 126 214
rect 124 213 125 214
rect 123 213 124 214
rect 122 213 123 214
rect 121 213 122 214
rect 120 213 121 214
rect 119 213 120 214
rect 118 213 119 214
rect 117 213 118 214
rect 116 213 117 214
rect 115 213 116 214
rect 114 213 115 214
rect 113 213 114 214
rect 112 213 113 214
rect 111 213 112 214
rect 110 213 111 214
rect 109 213 110 214
rect 108 213 109 214
rect 107 213 108 214
rect 106 213 107 214
rect 105 213 106 214
rect 104 213 105 214
rect 103 213 104 214
rect 102 213 103 214
rect 101 213 102 214
rect 100 213 101 214
rect 99 213 100 214
rect 98 213 99 214
rect 97 213 98 214
rect 96 213 97 214
rect 95 213 96 214
rect 94 213 95 214
rect 93 213 94 214
rect 92 213 93 214
rect 91 213 92 214
rect 90 213 91 214
rect 89 213 90 214
rect 88 213 89 214
rect 64 213 65 214
rect 63 213 64 214
rect 62 213 63 214
rect 61 213 62 214
rect 60 213 61 214
rect 59 213 60 214
rect 58 213 59 214
rect 57 213 58 214
rect 56 213 57 214
rect 55 213 56 214
rect 54 213 55 214
rect 53 213 54 214
rect 52 213 53 214
rect 51 213 52 214
rect 50 213 51 214
rect 49 213 50 214
rect 48 213 49 214
rect 47 213 48 214
rect 46 213 47 214
rect 45 213 46 214
rect 44 213 45 214
rect 43 213 44 214
rect 42 213 43 214
rect 41 213 42 214
rect 40 213 41 214
rect 39 213 40 214
rect 38 213 39 214
rect 37 213 38 214
rect 36 213 37 214
rect 35 213 36 214
rect 34 213 35 214
rect 33 213 34 214
rect 32 213 33 214
rect 31 213 32 214
rect 30 213 31 214
rect 29 213 30 214
rect 28 213 29 214
rect 27 213 28 214
rect 26 213 27 214
rect 25 213 26 214
rect 24 213 25 214
rect 23 213 24 214
rect 22 213 23 214
rect 21 213 22 214
rect 20 213 21 214
rect 19 213 20 214
rect 18 213 19 214
rect 17 213 18 214
rect 16 213 17 214
rect 15 213 16 214
rect 14 213 15 214
rect 13 213 14 214
rect 12 213 13 214
rect 11 213 12 214
rect 10 213 11 214
rect 9 213 10 214
rect 8 213 9 214
rect 434 214 435 215
rect 433 214 434 215
rect 432 214 433 215
rect 431 214 432 215
rect 430 214 431 215
rect 429 214 430 215
rect 428 214 429 215
rect 427 214 428 215
rect 426 214 427 215
rect 425 214 426 215
rect 424 214 425 215
rect 423 214 424 215
rect 422 214 423 215
rect 421 214 422 215
rect 420 214 421 215
rect 419 214 420 215
rect 418 214 419 215
rect 417 214 418 215
rect 416 214 417 215
rect 415 214 416 215
rect 414 214 415 215
rect 413 214 414 215
rect 412 214 413 215
rect 411 214 412 215
rect 410 214 411 215
rect 409 214 410 215
rect 408 214 409 215
rect 407 214 408 215
rect 406 214 407 215
rect 405 214 406 215
rect 404 214 405 215
rect 403 214 404 215
rect 402 214 403 215
rect 401 214 402 215
rect 358 214 359 215
rect 357 214 358 215
rect 356 214 357 215
rect 355 214 356 215
rect 354 214 355 215
rect 353 214 354 215
rect 352 214 353 215
rect 351 214 352 215
rect 350 214 351 215
rect 349 214 350 215
rect 348 214 349 215
rect 347 214 348 215
rect 346 214 347 215
rect 345 214 346 215
rect 344 214 345 215
rect 343 214 344 215
rect 342 214 343 215
rect 341 214 342 215
rect 340 214 341 215
rect 339 214 340 215
rect 338 214 339 215
rect 337 214 338 215
rect 336 214 337 215
rect 335 214 336 215
rect 334 214 335 215
rect 333 214 334 215
rect 332 214 333 215
rect 331 214 332 215
rect 330 214 331 215
rect 329 214 330 215
rect 328 214 329 215
rect 327 214 328 215
rect 326 214 327 215
rect 325 214 326 215
rect 324 214 325 215
rect 323 214 324 215
rect 322 214 323 215
rect 321 214 322 215
rect 320 214 321 215
rect 319 214 320 215
rect 318 214 319 215
rect 317 214 318 215
rect 316 214 317 215
rect 315 214 316 215
rect 314 214 315 215
rect 313 214 314 215
rect 312 214 313 215
rect 311 214 312 215
rect 310 214 311 215
rect 309 214 310 215
rect 308 214 309 215
rect 307 214 308 215
rect 306 214 307 215
rect 305 214 306 215
rect 304 214 305 215
rect 303 214 304 215
rect 302 214 303 215
rect 301 214 302 215
rect 300 214 301 215
rect 299 214 300 215
rect 298 214 299 215
rect 297 214 298 215
rect 296 214 297 215
rect 295 214 296 215
rect 294 214 295 215
rect 293 214 294 215
rect 292 214 293 215
rect 291 214 292 215
rect 290 214 291 215
rect 289 214 290 215
rect 288 214 289 215
rect 287 214 288 215
rect 286 214 287 215
rect 285 214 286 215
rect 284 214 285 215
rect 283 214 284 215
rect 282 214 283 215
rect 281 214 282 215
rect 280 214 281 215
rect 279 214 280 215
rect 278 214 279 215
rect 277 214 278 215
rect 276 214 277 215
rect 275 214 276 215
rect 274 214 275 215
rect 273 214 274 215
rect 272 214 273 215
rect 271 214 272 215
rect 270 214 271 215
rect 269 214 270 215
rect 268 214 269 215
rect 267 214 268 215
rect 266 214 267 215
rect 265 214 266 215
rect 264 214 265 215
rect 263 214 264 215
rect 262 214 263 215
rect 261 214 262 215
rect 260 214 261 215
rect 259 214 260 215
rect 258 214 259 215
rect 257 214 258 215
rect 256 214 257 215
rect 255 214 256 215
rect 254 214 255 215
rect 253 214 254 215
rect 252 214 253 215
rect 251 214 252 215
rect 250 214 251 215
rect 249 214 250 215
rect 248 214 249 215
rect 247 214 248 215
rect 246 214 247 215
rect 245 214 246 215
rect 244 214 245 215
rect 243 214 244 215
rect 242 214 243 215
rect 241 214 242 215
rect 240 214 241 215
rect 239 214 240 215
rect 238 214 239 215
rect 237 214 238 215
rect 236 214 237 215
rect 235 214 236 215
rect 234 214 235 215
rect 233 214 234 215
rect 232 214 233 215
rect 231 214 232 215
rect 230 214 231 215
rect 229 214 230 215
rect 228 214 229 215
rect 227 214 228 215
rect 226 214 227 215
rect 225 214 226 215
rect 224 214 225 215
rect 223 214 224 215
rect 222 214 223 215
rect 221 214 222 215
rect 220 214 221 215
rect 219 214 220 215
rect 218 214 219 215
rect 217 214 218 215
rect 216 214 217 215
rect 215 214 216 215
rect 214 214 215 215
rect 213 214 214 215
rect 212 214 213 215
rect 211 214 212 215
rect 210 214 211 215
rect 209 214 210 215
rect 208 214 209 215
rect 207 214 208 215
rect 206 214 207 215
rect 205 214 206 215
rect 204 214 205 215
rect 203 214 204 215
rect 202 214 203 215
rect 201 214 202 215
rect 200 214 201 215
rect 199 214 200 215
rect 198 214 199 215
rect 197 214 198 215
rect 196 214 197 215
rect 195 214 196 215
rect 194 214 195 215
rect 193 214 194 215
rect 192 214 193 215
rect 151 214 152 215
rect 150 214 151 215
rect 149 214 150 215
rect 148 214 149 215
rect 147 214 148 215
rect 146 214 147 215
rect 145 214 146 215
rect 144 214 145 215
rect 143 214 144 215
rect 142 214 143 215
rect 141 214 142 215
rect 140 214 141 215
rect 139 214 140 215
rect 138 214 139 215
rect 137 214 138 215
rect 136 214 137 215
rect 135 214 136 215
rect 134 214 135 215
rect 133 214 134 215
rect 132 214 133 215
rect 131 214 132 215
rect 130 214 131 215
rect 129 214 130 215
rect 128 214 129 215
rect 127 214 128 215
rect 126 214 127 215
rect 125 214 126 215
rect 124 214 125 215
rect 123 214 124 215
rect 122 214 123 215
rect 121 214 122 215
rect 120 214 121 215
rect 119 214 120 215
rect 118 214 119 215
rect 117 214 118 215
rect 116 214 117 215
rect 115 214 116 215
rect 114 214 115 215
rect 113 214 114 215
rect 112 214 113 215
rect 111 214 112 215
rect 110 214 111 215
rect 109 214 110 215
rect 108 214 109 215
rect 107 214 108 215
rect 106 214 107 215
rect 105 214 106 215
rect 104 214 105 215
rect 103 214 104 215
rect 102 214 103 215
rect 101 214 102 215
rect 100 214 101 215
rect 99 214 100 215
rect 98 214 99 215
rect 97 214 98 215
rect 96 214 97 215
rect 95 214 96 215
rect 94 214 95 215
rect 93 214 94 215
rect 92 214 93 215
rect 91 214 92 215
rect 90 214 91 215
rect 65 214 66 215
rect 64 214 65 215
rect 63 214 64 215
rect 62 214 63 215
rect 61 214 62 215
rect 60 214 61 215
rect 59 214 60 215
rect 58 214 59 215
rect 57 214 58 215
rect 56 214 57 215
rect 55 214 56 215
rect 54 214 55 215
rect 53 214 54 215
rect 52 214 53 215
rect 51 214 52 215
rect 50 214 51 215
rect 49 214 50 215
rect 48 214 49 215
rect 47 214 48 215
rect 46 214 47 215
rect 45 214 46 215
rect 44 214 45 215
rect 43 214 44 215
rect 42 214 43 215
rect 41 214 42 215
rect 40 214 41 215
rect 39 214 40 215
rect 38 214 39 215
rect 37 214 38 215
rect 36 214 37 215
rect 35 214 36 215
rect 34 214 35 215
rect 33 214 34 215
rect 32 214 33 215
rect 31 214 32 215
rect 30 214 31 215
rect 29 214 30 215
rect 28 214 29 215
rect 27 214 28 215
rect 26 214 27 215
rect 25 214 26 215
rect 24 214 25 215
rect 23 214 24 215
rect 22 214 23 215
rect 21 214 22 215
rect 20 214 21 215
rect 19 214 20 215
rect 18 214 19 215
rect 17 214 18 215
rect 16 214 17 215
rect 15 214 16 215
rect 14 214 15 215
rect 13 214 14 215
rect 12 214 13 215
rect 11 214 12 215
rect 10 214 11 215
rect 9 214 10 215
rect 8 214 9 215
rect 435 215 436 216
rect 434 215 435 216
rect 433 215 434 216
rect 432 215 433 216
rect 431 215 432 216
rect 430 215 431 216
rect 429 215 430 216
rect 428 215 429 216
rect 427 215 428 216
rect 426 215 427 216
rect 425 215 426 216
rect 424 215 425 216
rect 423 215 424 216
rect 422 215 423 216
rect 421 215 422 216
rect 420 215 421 216
rect 419 215 420 216
rect 418 215 419 216
rect 417 215 418 216
rect 416 215 417 216
rect 415 215 416 216
rect 414 215 415 216
rect 413 215 414 216
rect 412 215 413 216
rect 411 215 412 216
rect 410 215 411 216
rect 409 215 410 216
rect 408 215 409 216
rect 407 215 408 216
rect 406 215 407 216
rect 405 215 406 216
rect 404 215 405 216
rect 403 215 404 216
rect 402 215 403 216
rect 401 215 402 216
rect 400 215 401 216
rect 359 215 360 216
rect 358 215 359 216
rect 357 215 358 216
rect 356 215 357 216
rect 355 215 356 216
rect 354 215 355 216
rect 353 215 354 216
rect 352 215 353 216
rect 351 215 352 216
rect 350 215 351 216
rect 349 215 350 216
rect 348 215 349 216
rect 347 215 348 216
rect 346 215 347 216
rect 345 215 346 216
rect 344 215 345 216
rect 343 215 344 216
rect 342 215 343 216
rect 341 215 342 216
rect 340 215 341 216
rect 339 215 340 216
rect 338 215 339 216
rect 337 215 338 216
rect 336 215 337 216
rect 335 215 336 216
rect 334 215 335 216
rect 333 215 334 216
rect 332 215 333 216
rect 331 215 332 216
rect 311 215 312 216
rect 310 215 311 216
rect 309 215 310 216
rect 308 215 309 216
rect 307 215 308 216
rect 306 215 307 216
rect 305 215 306 216
rect 304 215 305 216
rect 303 215 304 216
rect 302 215 303 216
rect 301 215 302 216
rect 300 215 301 216
rect 299 215 300 216
rect 298 215 299 216
rect 297 215 298 216
rect 296 215 297 216
rect 295 215 296 216
rect 294 215 295 216
rect 293 215 294 216
rect 292 215 293 216
rect 291 215 292 216
rect 290 215 291 216
rect 289 215 290 216
rect 288 215 289 216
rect 287 215 288 216
rect 286 215 287 216
rect 285 215 286 216
rect 284 215 285 216
rect 283 215 284 216
rect 282 215 283 216
rect 281 215 282 216
rect 280 215 281 216
rect 279 215 280 216
rect 278 215 279 216
rect 277 215 278 216
rect 276 215 277 216
rect 275 215 276 216
rect 274 215 275 216
rect 273 215 274 216
rect 272 215 273 216
rect 271 215 272 216
rect 270 215 271 216
rect 269 215 270 216
rect 268 215 269 216
rect 267 215 268 216
rect 266 215 267 216
rect 265 215 266 216
rect 264 215 265 216
rect 263 215 264 216
rect 262 215 263 216
rect 261 215 262 216
rect 260 215 261 216
rect 259 215 260 216
rect 258 215 259 216
rect 257 215 258 216
rect 256 215 257 216
rect 255 215 256 216
rect 254 215 255 216
rect 253 215 254 216
rect 252 215 253 216
rect 251 215 252 216
rect 250 215 251 216
rect 249 215 250 216
rect 248 215 249 216
rect 247 215 248 216
rect 246 215 247 216
rect 245 215 246 216
rect 244 215 245 216
rect 243 215 244 216
rect 242 215 243 216
rect 241 215 242 216
rect 240 215 241 216
rect 239 215 240 216
rect 238 215 239 216
rect 237 215 238 216
rect 236 215 237 216
rect 235 215 236 216
rect 234 215 235 216
rect 233 215 234 216
rect 232 215 233 216
rect 231 215 232 216
rect 230 215 231 216
rect 229 215 230 216
rect 228 215 229 216
rect 227 215 228 216
rect 226 215 227 216
rect 225 215 226 216
rect 224 215 225 216
rect 223 215 224 216
rect 222 215 223 216
rect 221 215 222 216
rect 220 215 221 216
rect 219 215 220 216
rect 218 215 219 216
rect 217 215 218 216
rect 216 215 217 216
rect 215 215 216 216
rect 214 215 215 216
rect 213 215 214 216
rect 212 215 213 216
rect 211 215 212 216
rect 210 215 211 216
rect 209 215 210 216
rect 208 215 209 216
rect 207 215 208 216
rect 206 215 207 216
rect 205 215 206 216
rect 204 215 205 216
rect 203 215 204 216
rect 202 215 203 216
rect 201 215 202 216
rect 200 215 201 216
rect 199 215 200 216
rect 198 215 199 216
rect 197 215 198 216
rect 196 215 197 216
rect 195 215 196 216
rect 194 215 195 216
rect 193 215 194 216
rect 192 215 193 216
rect 191 215 192 216
rect 190 215 191 216
rect 149 215 150 216
rect 148 215 149 216
rect 147 215 148 216
rect 146 215 147 216
rect 145 215 146 216
rect 144 215 145 216
rect 143 215 144 216
rect 142 215 143 216
rect 141 215 142 216
rect 140 215 141 216
rect 139 215 140 216
rect 138 215 139 216
rect 137 215 138 216
rect 136 215 137 216
rect 135 215 136 216
rect 134 215 135 216
rect 133 215 134 216
rect 132 215 133 216
rect 131 215 132 216
rect 130 215 131 216
rect 129 215 130 216
rect 128 215 129 216
rect 127 215 128 216
rect 126 215 127 216
rect 125 215 126 216
rect 124 215 125 216
rect 123 215 124 216
rect 122 215 123 216
rect 121 215 122 216
rect 120 215 121 216
rect 119 215 120 216
rect 118 215 119 216
rect 117 215 118 216
rect 116 215 117 216
rect 115 215 116 216
rect 114 215 115 216
rect 113 215 114 216
rect 112 215 113 216
rect 111 215 112 216
rect 110 215 111 216
rect 109 215 110 216
rect 108 215 109 216
rect 107 215 108 216
rect 106 215 107 216
rect 105 215 106 216
rect 104 215 105 216
rect 103 215 104 216
rect 102 215 103 216
rect 101 215 102 216
rect 100 215 101 216
rect 99 215 100 216
rect 98 215 99 216
rect 97 215 98 216
rect 96 215 97 216
rect 95 215 96 216
rect 94 215 95 216
rect 93 215 94 216
rect 66 215 67 216
rect 65 215 66 216
rect 64 215 65 216
rect 63 215 64 216
rect 62 215 63 216
rect 61 215 62 216
rect 60 215 61 216
rect 59 215 60 216
rect 58 215 59 216
rect 57 215 58 216
rect 56 215 57 216
rect 55 215 56 216
rect 54 215 55 216
rect 53 215 54 216
rect 52 215 53 216
rect 51 215 52 216
rect 50 215 51 216
rect 49 215 50 216
rect 48 215 49 216
rect 47 215 48 216
rect 46 215 47 216
rect 45 215 46 216
rect 44 215 45 216
rect 43 215 44 216
rect 42 215 43 216
rect 41 215 42 216
rect 40 215 41 216
rect 39 215 40 216
rect 38 215 39 216
rect 37 215 38 216
rect 36 215 37 216
rect 35 215 36 216
rect 34 215 35 216
rect 33 215 34 216
rect 32 215 33 216
rect 31 215 32 216
rect 30 215 31 216
rect 29 215 30 216
rect 28 215 29 216
rect 27 215 28 216
rect 26 215 27 216
rect 25 215 26 216
rect 24 215 25 216
rect 23 215 24 216
rect 22 215 23 216
rect 21 215 22 216
rect 20 215 21 216
rect 19 215 20 216
rect 18 215 19 216
rect 17 215 18 216
rect 16 215 17 216
rect 15 215 16 216
rect 14 215 15 216
rect 13 215 14 216
rect 12 215 13 216
rect 11 215 12 216
rect 10 215 11 216
rect 9 215 10 216
rect 8 215 9 216
rect 480 216 481 217
rect 460 216 461 217
rect 436 216 437 217
rect 435 216 436 217
rect 434 216 435 217
rect 433 216 434 217
rect 432 216 433 217
rect 431 216 432 217
rect 430 216 431 217
rect 429 216 430 217
rect 428 216 429 217
rect 427 216 428 217
rect 426 216 427 217
rect 425 216 426 217
rect 424 216 425 217
rect 423 216 424 217
rect 422 216 423 217
rect 421 216 422 217
rect 420 216 421 217
rect 419 216 420 217
rect 418 216 419 217
rect 417 216 418 217
rect 416 216 417 217
rect 415 216 416 217
rect 414 216 415 217
rect 413 216 414 217
rect 412 216 413 217
rect 411 216 412 217
rect 410 216 411 217
rect 409 216 410 217
rect 408 216 409 217
rect 407 216 408 217
rect 406 216 407 217
rect 405 216 406 217
rect 404 216 405 217
rect 403 216 404 217
rect 402 216 403 217
rect 401 216 402 217
rect 400 216 401 217
rect 399 216 400 217
rect 359 216 360 217
rect 358 216 359 217
rect 357 216 358 217
rect 356 216 357 217
rect 355 216 356 217
rect 354 216 355 217
rect 353 216 354 217
rect 352 216 353 217
rect 351 216 352 217
rect 350 216 351 217
rect 349 216 350 217
rect 348 216 349 217
rect 347 216 348 217
rect 346 216 347 217
rect 345 216 346 217
rect 344 216 345 217
rect 343 216 344 217
rect 342 216 343 217
rect 341 216 342 217
rect 340 216 341 217
rect 339 216 340 217
rect 338 216 339 217
rect 337 216 338 217
rect 305 216 306 217
rect 304 216 305 217
rect 303 216 304 217
rect 302 216 303 217
rect 301 216 302 217
rect 300 216 301 217
rect 299 216 300 217
rect 298 216 299 217
rect 297 216 298 217
rect 296 216 297 217
rect 295 216 296 217
rect 294 216 295 217
rect 293 216 294 217
rect 292 216 293 217
rect 291 216 292 217
rect 290 216 291 217
rect 289 216 290 217
rect 288 216 289 217
rect 287 216 288 217
rect 286 216 287 217
rect 285 216 286 217
rect 284 216 285 217
rect 283 216 284 217
rect 282 216 283 217
rect 281 216 282 217
rect 280 216 281 217
rect 279 216 280 217
rect 278 216 279 217
rect 277 216 278 217
rect 276 216 277 217
rect 275 216 276 217
rect 274 216 275 217
rect 273 216 274 217
rect 272 216 273 217
rect 271 216 272 217
rect 270 216 271 217
rect 269 216 270 217
rect 268 216 269 217
rect 267 216 268 217
rect 266 216 267 217
rect 265 216 266 217
rect 264 216 265 217
rect 263 216 264 217
rect 262 216 263 217
rect 261 216 262 217
rect 260 216 261 217
rect 259 216 260 217
rect 258 216 259 217
rect 257 216 258 217
rect 256 216 257 217
rect 255 216 256 217
rect 254 216 255 217
rect 253 216 254 217
rect 252 216 253 217
rect 251 216 252 217
rect 250 216 251 217
rect 249 216 250 217
rect 248 216 249 217
rect 247 216 248 217
rect 246 216 247 217
rect 245 216 246 217
rect 244 216 245 217
rect 243 216 244 217
rect 242 216 243 217
rect 241 216 242 217
rect 240 216 241 217
rect 239 216 240 217
rect 238 216 239 217
rect 237 216 238 217
rect 236 216 237 217
rect 235 216 236 217
rect 234 216 235 217
rect 233 216 234 217
rect 232 216 233 217
rect 231 216 232 217
rect 230 216 231 217
rect 229 216 230 217
rect 228 216 229 217
rect 227 216 228 217
rect 226 216 227 217
rect 225 216 226 217
rect 224 216 225 217
rect 223 216 224 217
rect 222 216 223 217
rect 221 216 222 217
rect 220 216 221 217
rect 219 216 220 217
rect 218 216 219 217
rect 217 216 218 217
rect 216 216 217 217
rect 215 216 216 217
rect 214 216 215 217
rect 213 216 214 217
rect 212 216 213 217
rect 211 216 212 217
rect 210 216 211 217
rect 209 216 210 217
rect 208 216 209 217
rect 207 216 208 217
rect 206 216 207 217
rect 205 216 206 217
rect 204 216 205 217
rect 203 216 204 217
rect 202 216 203 217
rect 201 216 202 217
rect 200 216 201 217
rect 199 216 200 217
rect 198 216 199 217
rect 197 216 198 217
rect 196 216 197 217
rect 195 216 196 217
rect 194 216 195 217
rect 193 216 194 217
rect 192 216 193 217
rect 191 216 192 217
rect 190 216 191 217
rect 189 216 190 217
rect 188 216 189 217
rect 148 216 149 217
rect 147 216 148 217
rect 146 216 147 217
rect 145 216 146 217
rect 144 216 145 217
rect 143 216 144 217
rect 142 216 143 217
rect 141 216 142 217
rect 140 216 141 217
rect 139 216 140 217
rect 138 216 139 217
rect 137 216 138 217
rect 136 216 137 217
rect 135 216 136 217
rect 134 216 135 217
rect 133 216 134 217
rect 132 216 133 217
rect 131 216 132 217
rect 130 216 131 217
rect 129 216 130 217
rect 128 216 129 217
rect 127 216 128 217
rect 126 216 127 217
rect 125 216 126 217
rect 124 216 125 217
rect 123 216 124 217
rect 122 216 123 217
rect 121 216 122 217
rect 120 216 121 217
rect 119 216 120 217
rect 118 216 119 217
rect 117 216 118 217
rect 116 216 117 217
rect 115 216 116 217
rect 114 216 115 217
rect 113 216 114 217
rect 112 216 113 217
rect 111 216 112 217
rect 110 216 111 217
rect 109 216 110 217
rect 108 216 109 217
rect 107 216 108 217
rect 106 216 107 217
rect 105 216 106 217
rect 104 216 105 217
rect 103 216 104 217
rect 102 216 103 217
rect 101 216 102 217
rect 100 216 101 217
rect 99 216 100 217
rect 98 216 99 217
rect 97 216 98 217
rect 96 216 97 217
rect 95 216 96 217
rect 67 216 68 217
rect 66 216 67 217
rect 65 216 66 217
rect 64 216 65 217
rect 63 216 64 217
rect 62 216 63 217
rect 61 216 62 217
rect 60 216 61 217
rect 59 216 60 217
rect 58 216 59 217
rect 57 216 58 217
rect 56 216 57 217
rect 55 216 56 217
rect 54 216 55 217
rect 53 216 54 217
rect 52 216 53 217
rect 51 216 52 217
rect 50 216 51 217
rect 49 216 50 217
rect 48 216 49 217
rect 47 216 48 217
rect 46 216 47 217
rect 45 216 46 217
rect 44 216 45 217
rect 43 216 44 217
rect 42 216 43 217
rect 41 216 42 217
rect 40 216 41 217
rect 39 216 40 217
rect 38 216 39 217
rect 37 216 38 217
rect 36 216 37 217
rect 35 216 36 217
rect 34 216 35 217
rect 33 216 34 217
rect 32 216 33 217
rect 31 216 32 217
rect 30 216 31 217
rect 29 216 30 217
rect 28 216 29 217
rect 27 216 28 217
rect 26 216 27 217
rect 25 216 26 217
rect 24 216 25 217
rect 23 216 24 217
rect 22 216 23 217
rect 21 216 22 217
rect 20 216 21 217
rect 19 216 20 217
rect 18 216 19 217
rect 17 216 18 217
rect 16 216 17 217
rect 15 216 16 217
rect 14 216 15 217
rect 13 216 14 217
rect 12 216 13 217
rect 11 216 12 217
rect 10 216 11 217
rect 9 216 10 217
rect 8 216 9 217
rect 480 217 481 218
rect 460 217 461 218
rect 436 217 437 218
rect 435 217 436 218
rect 434 217 435 218
rect 433 217 434 218
rect 432 217 433 218
rect 431 217 432 218
rect 430 217 431 218
rect 429 217 430 218
rect 428 217 429 218
rect 427 217 428 218
rect 426 217 427 218
rect 425 217 426 218
rect 424 217 425 218
rect 423 217 424 218
rect 422 217 423 218
rect 421 217 422 218
rect 420 217 421 218
rect 419 217 420 218
rect 418 217 419 218
rect 417 217 418 218
rect 416 217 417 218
rect 415 217 416 218
rect 414 217 415 218
rect 413 217 414 218
rect 412 217 413 218
rect 411 217 412 218
rect 410 217 411 218
rect 409 217 410 218
rect 408 217 409 218
rect 407 217 408 218
rect 406 217 407 218
rect 405 217 406 218
rect 404 217 405 218
rect 403 217 404 218
rect 402 217 403 218
rect 401 217 402 218
rect 400 217 401 218
rect 399 217 400 218
rect 360 217 361 218
rect 359 217 360 218
rect 358 217 359 218
rect 357 217 358 218
rect 356 217 357 218
rect 355 217 356 218
rect 354 217 355 218
rect 353 217 354 218
rect 352 217 353 218
rect 351 217 352 218
rect 350 217 351 218
rect 349 217 350 218
rect 348 217 349 218
rect 347 217 348 218
rect 346 217 347 218
rect 345 217 346 218
rect 344 217 345 218
rect 343 217 344 218
rect 342 217 343 218
rect 301 217 302 218
rect 300 217 301 218
rect 299 217 300 218
rect 298 217 299 218
rect 297 217 298 218
rect 296 217 297 218
rect 295 217 296 218
rect 294 217 295 218
rect 293 217 294 218
rect 292 217 293 218
rect 291 217 292 218
rect 290 217 291 218
rect 289 217 290 218
rect 288 217 289 218
rect 287 217 288 218
rect 286 217 287 218
rect 285 217 286 218
rect 284 217 285 218
rect 283 217 284 218
rect 282 217 283 218
rect 281 217 282 218
rect 280 217 281 218
rect 279 217 280 218
rect 278 217 279 218
rect 277 217 278 218
rect 276 217 277 218
rect 275 217 276 218
rect 274 217 275 218
rect 273 217 274 218
rect 272 217 273 218
rect 271 217 272 218
rect 270 217 271 218
rect 269 217 270 218
rect 268 217 269 218
rect 267 217 268 218
rect 266 217 267 218
rect 265 217 266 218
rect 264 217 265 218
rect 263 217 264 218
rect 262 217 263 218
rect 261 217 262 218
rect 260 217 261 218
rect 259 217 260 218
rect 258 217 259 218
rect 257 217 258 218
rect 256 217 257 218
rect 255 217 256 218
rect 254 217 255 218
rect 253 217 254 218
rect 252 217 253 218
rect 251 217 252 218
rect 250 217 251 218
rect 249 217 250 218
rect 248 217 249 218
rect 247 217 248 218
rect 246 217 247 218
rect 245 217 246 218
rect 244 217 245 218
rect 243 217 244 218
rect 242 217 243 218
rect 241 217 242 218
rect 240 217 241 218
rect 239 217 240 218
rect 238 217 239 218
rect 237 217 238 218
rect 236 217 237 218
rect 235 217 236 218
rect 234 217 235 218
rect 233 217 234 218
rect 232 217 233 218
rect 231 217 232 218
rect 230 217 231 218
rect 229 217 230 218
rect 228 217 229 218
rect 227 217 228 218
rect 226 217 227 218
rect 225 217 226 218
rect 224 217 225 218
rect 223 217 224 218
rect 222 217 223 218
rect 221 217 222 218
rect 220 217 221 218
rect 219 217 220 218
rect 218 217 219 218
rect 217 217 218 218
rect 216 217 217 218
rect 215 217 216 218
rect 214 217 215 218
rect 213 217 214 218
rect 212 217 213 218
rect 211 217 212 218
rect 210 217 211 218
rect 209 217 210 218
rect 208 217 209 218
rect 207 217 208 218
rect 206 217 207 218
rect 205 217 206 218
rect 204 217 205 218
rect 203 217 204 218
rect 202 217 203 218
rect 201 217 202 218
rect 200 217 201 218
rect 199 217 200 218
rect 198 217 199 218
rect 197 217 198 218
rect 196 217 197 218
rect 195 217 196 218
rect 194 217 195 218
rect 193 217 194 218
rect 192 217 193 218
rect 191 217 192 218
rect 190 217 191 218
rect 189 217 190 218
rect 188 217 189 218
rect 187 217 188 218
rect 186 217 187 218
rect 147 217 148 218
rect 146 217 147 218
rect 145 217 146 218
rect 144 217 145 218
rect 143 217 144 218
rect 142 217 143 218
rect 141 217 142 218
rect 140 217 141 218
rect 139 217 140 218
rect 138 217 139 218
rect 137 217 138 218
rect 136 217 137 218
rect 135 217 136 218
rect 134 217 135 218
rect 133 217 134 218
rect 132 217 133 218
rect 131 217 132 218
rect 130 217 131 218
rect 129 217 130 218
rect 128 217 129 218
rect 127 217 128 218
rect 126 217 127 218
rect 125 217 126 218
rect 124 217 125 218
rect 123 217 124 218
rect 122 217 123 218
rect 121 217 122 218
rect 120 217 121 218
rect 119 217 120 218
rect 118 217 119 218
rect 117 217 118 218
rect 116 217 117 218
rect 115 217 116 218
rect 114 217 115 218
rect 113 217 114 218
rect 112 217 113 218
rect 111 217 112 218
rect 110 217 111 218
rect 109 217 110 218
rect 108 217 109 218
rect 107 217 108 218
rect 106 217 107 218
rect 105 217 106 218
rect 104 217 105 218
rect 103 217 104 218
rect 102 217 103 218
rect 101 217 102 218
rect 100 217 101 218
rect 99 217 100 218
rect 98 217 99 218
rect 97 217 98 218
rect 68 217 69 218
rect 67 217 68 218
rect 66 217 67 218
rect 65 217 66 218
rect 64 217 65 218
rect 63 217 64 218
rect 62 217 63 218
rect 61 217 62 218
rect 60 217 61 218
rect 59 217 60 218
rect 58 217 59 218
rect 57 217 58 218
rect 56 217 57 218
rect 55 217 56 218
rect 54 217 55 218
rect 53 217 54 218
rect 52 217 53 218
rect 51 217 52 218
rect 50 217 51 218
rect 49 217 50 218
rect 48 217 49 218
rect 47 217 48 218
rect 46 217 47 218
rect 45 217 46 218
rect 44 217 45 218
rect 43 217 44 218
rect 42 217 43 218
rect 41 217 42 218
rect 40 217 41 218
rect 39 217 40 218
rect 38 217 39 218
rect 37 217 38 218
rect 36 217 37 218
rect 35 217 36 218
rect 34 217 35 218
rect 33 217 34 218
rect 32 217 33 218
rect 31 217 32 218
rect 30 217 31 218
rect 29 217 30 218
rect 28 217 29 218
rect 27 217 28 218
rect 26 217 27 218
rect 25 217 26 218
rect 24 217 25 218
rect 23 217 24 218
rect 22 217 23 218
rect 21 217 22 218
rect 20 217 21 218
rect 19 217 20 218
rect 18 217 19 218
rect 17 217 18 218
rect 16 217 17 218
rect 15 217 16 218
rect 14 217 15 218
rect 13 217 14 218
rect 12 217 13 218
rect 11 217 12 218
rect 10 217 11 218
rect 9 217 10 218
rect 8 217 9 218
rect 7 217 8 218
rect 480 218 481 219
rect 479 218 480 219
rect 478 218 479 219
rect 462 218 463 219
rect 461 218 462 219
rect 460 218 461 219
rect 437 218 438 219
rect 436 218 437 219
rect 435 218 436 219
rect 434 218 435 219
rect 433 218 434 219
rect 432 218 433 219
rect 431 218 432 219
rect 430 218 431 219
rect 429 218 430 219
rect 428 218 429 219
rect 427 218 428 219
rect 426 218 427 219
rect 425 218 426 219
rect 424 218 425 219
rect 423 218 424 219
rect 410 218 411 219
rect 409 218 410 219
rect 408 218 409 219
rect 407 218 408 219
rect 406 218 407 219
rect 405 218 406 219
rect 404 218 405 219
rect 403 218 404 219
rect 402 218 403 219
rect 401 218 402 219
rect 400 218 401 219
rect 399 218 400 219
rect 398 218 399 219
rect 360 218 361 219
rect 359 218 360 219
rect 358 218 359 219
rect 357 218 358 219
rect 356 218 357 219
rect 355 218 356 219
rect 354 218 355 219
rect 353 218 354 219
rect 352 218 353 219
rect 351 218 352 219
rect 350 218 351 219
rect 349 218 350 219
rect 348 218 349 219
rect 347 218 348 219
rect 346 218 347 219
rect 298 218 299 219
rect 297 218 298 219
rect 296 218 297 219
rect 295 218 296 219
rect 294 218 295 219
rect 293 218 294 219
rect 292 218 293 219
rect 291 218 292 219
rect 290 218 291 219
rect 289 218 290 219
rect 288 218 289 219
rect 287 218 288 219
rect 286 218 287 219
rect 285 218 286 219
rect 284 218 285 219
rect 283 218 284 219
rect 282 218 283 219
rect 281 218 282 219
rect 280 218 281 219
rect 279 218 280 219
rect 278 218 279 219
rect 277 218 278 219
rect 276 218 277 219
rect 275 218 276 219
rect 274 218 275 219
rect 273 218 274 219
rect 272 218 273 219
rect 271 218 272 219
rect 270 218 271 219
rect 269 218 270 219
rect 268 218 269 219
rect 267 218 268 219
rect 266 218 267 219
rect 265 218 266 219
rect 264 218 265 219
rect 263 218 264 219
rect 262 218 263 219
rect 261 218 262 219
rect 260 218 261 219
rect 259 218 260 219
rect 258 218 259 219
rect 257 218 258 219
rect 256 218 257 219
rect 255 218 256 219
rect 254 218 255 219
rect 253 218 254 219
rect 252 218 253 219
rect 251 218 252 219
rect 250 218 251 219
rect 249 218 250 219
rect 248 218 249 219
rect 247 218 248 219
rect 246 218 247 219
rect 245 218 246 219
rect 244 218 245 219
rect 243 218 244 219
rect 242 218 243 219
rect 241 218 242 219
rect 240 218 241 219
rect 239 218 240 219
rect 238 218 239 219
rect 237 218 238 219
rect 236 218 237 219
rect 235 218 236 219
rect 234 218 235 219
rect 233 218 234 219
rect 232 218 233 219
rect 231 218 232 219
rect 230 218 231 219
rect 229 218 230 219
rect 228 218 229 219
rect 227 218 228 219
rect 226 218 227 219
rect 225 218 226 219
rect 224 218 225 219
rect 223 218 224 219
rect 222 218 223 219
rect 221 218 222 219
rect 220 218 221 219
rect 219 218 220 219
rect 218 218 219 219
rect 217 218 218 219
rect 216 218 217 219
rect 215 218 216 219
rect 214 218 215 219
rect 213 218 214 219
rect 212 218 213 219
rect 211 218 212 219
rect 210 218 211 219
rect 209 218 210 219
rect 208 218 209 219
rect 207 218 208 219
rect 206 218 207 219
rect 205 218 206 219
rect 204 218 205 219
rect 203 218 204 219
rect 202 218 203 219
rect 201 218 202 219
rect 200 218 201 219
rect 199 218 200 219
rect 198 218 199 219
rect 197 218 198 219
rect 196 218 197 219
rect 195 218 196 219
rect 194 218 195 219
rect 193 218 194 219
rect 192 218 193 219
rect 191 218 192 219
rect 190 218 191 219
rect 189 218 190 219
rect 188 218 189 219
rect 187 218 188 219
rect 186 218 187 219
rect 185 218 186 219
rect 184 218 185 219
rect 183 218 184 219
rect 146 218 147 219
rect 145 218 146 219
rect 144 218 145 219
rect 143 218 144 219
rect 142 218 143 219
rect 141 218 142 219
rect 140 218 141 219
rect 139 218 140 219
rect 138 218 139 219
rect 137 218 138 219
rect 136 218 137 219
rect 135 218 136 219
rect 134 218 135 219
rect 133 218 134 219
rect 132 218 133 219
rect 131 218 132 219
rect 130 218 131 219
rect 129 218 130 219
rect 128 218 129 219
rect 127 218 128 219
rect 126 218 127 219
rect 125 218 126 219
rect 124 218 125 219
rect 123 218 124 219
rect 122 218 123 219
rect 121 218 122 219
rect 120 218 121 219
rect 119 218 120 219
rect 118 218 119 219
rect 117 218 118 219
rect 116 218 117 219
rect 115 218 116 219
rect 114 218 115 219
rect 113 218 114 219
rect 112 218 113 219
rect 111 218 112 219
rect 110 218 111 219
rect 109 218 110 219
rect 108 218 109 219
rect 107 218 108 219
rect 106 218 107 219
rect 105 218 106 219
rect 104 218 105 219
rect 103 218 104 219
rect 102 218 103 219
rect 101 218 102 219
rect 100 218 101 219
rect 99 218 100 219
rect 69 218 70 219
rect 68 218 69 219
rect 67 218 68 219
rect 66 218 67 219
rect 65 218 66 219
rect 64 218 65 219
rect 63 218 64 219
rect 62 218 63 219
rect 61 218 62 219
rect 60 218 61 219
rect 59 218 60 219
rect 58 218 59 219
rect 57 218 58 219
rect 56 218 57 219
rect 55 218 56 219
rect 54 218 55 219
rect 53 218 54 219
rect 52 218 53 219
rect 51 218 52 219
rect 50 218 51 219
rect 49 218 50 219
rect 48 218 49 219
rect 47 218 48 219
rect 46 218 47 219
rect 45 218 46 219
rect 44 218 45 219
rect 43 218 44 219
rect 42 218 43 219
rect 41 218 42 219
rect 40 218 41 219
rect 39 218 40 219
rect 38 218 39 219
rect 37 218 38 219
rect 36 218 37 219
rect 35 218 36 219
rect 34 218 35 219
rect 33 218 34 219
rect 32 218 33 219
rect 31 218 32 219
rect 30 218 31 219
rect 29 218 30 219
rect 28 218 29 219
rect 27 218 28 219
rect 26 218 27 219
rect 25 218 26 219
rect 24 218 25 219
rect 23 218 24 219
rect 22 218 23 219
rect 21 218 22 219
rect 20 218 21 219
rect 19 218 20 219
rect 18 218 19 219
rect 17 218 18 219
rect 16 218 17 219
rect 15 218 16 219
rect 14 218 15 219
rect 13 218 14 219
rect 12 218 13 219
rect 11 218 12 219
rect 10 218 11 219
rect 9 218 10 219
rect 8 218 9 219
rect 7 218 8 219
rect 480 219 481 220
rect 479 219 480 220
rect 478 219 479 220
rect 477 219 478 220
rect 476 219 477 220
rect 475 219 476 220
rect 474 219 475 220
rect 473 219 474 220
rect 472 219 473 220
rect 471 219 472 220
rect 470 219 471 220
rect 469 219 470 220
rect 468 219 469 220
rect 467 219 468 220
rect 466 219 467 220
rect 465 219 466 220
rect 464 219 465 220
rect 463 219 464 220
rect 462 219 463 220
rect 461 219 462 220
rect 460 219 461 220
rect 437 219 438 220
rect 436 219 437 220
rect 435 219 436 220
rect 434 219 435 220
rect 433 219 434 220
rect 432 219 433 220
rect 431 219 432 220
rect 430 219 431 220
rect 429 219 430 220
rect 428 219 429 220
rect 427 219 428 220
rect 406 219 407 220
rect 405 219 406 220
rect 404 219 405 220
rect 403 219 404 220
rect 402 219 403 220
rect 401 219 402 220
rect 400 219 401 220
rect 399 219 400 220
rect 398 219 399 220
rect 397 219 398 220
rect 361 219 362 220
rect 360 219 361 220
rect 359 219 360 220
rect 358 219 359 220
rect 357 219 358 220
rect 356 219 357 220
rect 355 219 356 220
rect 354 219 355 220
rect 353 219 354 220
rect 352 219 353 220
rect 351 219 352 220
rect 350 219 351 220
rect 349 219 350 220
rect 295 219 296 220
rect 294 219 295 220
rect 293 219 294 220
rect 292 219 293 220
rect 291 219 292 220
rect 290 219 291 220
rect 289 219 290 220
rect 288 219 289 220
rect 287 219 288 220
rect 286 219 287 220
rect 285 219 286 220
rect 284 219 285 220
rect 283 219 284 220
rect 282 219 283 220
rect 281 219 282 220
rect 280 219 281 220
rect 279 219 280 220
rect 278 219 279 220
rect 277 219 278 220
rect 276 219 277 220
rect 275 219 276 220
rect 274 219 275 220
rect 273 219 274 220
rect 272 219 273 220
rect 271 219 272 220
rect 270 219 271 220
rect 269 219 270 220
rect 268 219 269 220
rect 267 219 268 220
rect 266 219 267 220
rect 265 219 266 220
rect 264 219 265 220
rect 263 219 264 220
rect 262 219 263 220
rect 261 219 262 220
rect 260 219 261 220
rect 259 219 260 220
rect 258 219 259 220
rect 257 219 258 220
rect 256 219 257 220
rect 255 219 256 220
rect 254 219 255 220
rect 253 219 254 220
rect 252 219 253 220
rect 251 219 252 220
rect 250 219 251 220
rect 249 219 250 220
rect 248 219 249 220
rect 247 219 248 220
rect 246 219 247 220
rect 245 219 246 220
rect 244 219 245 220
rect 243 219 244 220
rect 242 219 243 220
rect 241 219 242 220
rect 240 219 241 220
rect 239 219 240 220
rect 238 219 239 220
rect 237 219 238 220
rect 236 219 237 220
rect 235 219 236 220
rect 234 219 235 220
rect 233 219 234 220
rect 232 219 233 220
rect 231 219 232 220
rect 230 219 231 220
rect 229 219 230 220
rect 228 219 229 220
rect 227 219 228 220
rect 226 219 227 220
rect 225 219 226 220
rect 224 219 225 220
rect 223 219 224 220
rect 222 219 223 220
rect 221 219 222 220
rect 220 219 221 220
rect 219 219 220 220
rect 218 219 219 220
rect 217 219 218 220
rect 216 219 217 220
rect 215 219 216 220
rect 214 219 215 220
rect 213 219 214 220
rect 212 219 213 220
rect 211 219 212 220
rect 210 219 211 220
rect 209 219 210 220
rect 208 219 209 220
rect 207 219 208 220
rect 206 219 207 220
rect 205 219 206 220
rect 204 219 205 220
rect 203 219 204 220
rect 202 219 203 220
rect 201 219 202 220
rect 200 219 201 220
rect 199 219 200 220
rect 198 219 199 220
rect 197 219 198 220
rect 196 219 197 220
rect 195 219 196 220
rect 194 219 195 220
rect 193 219 194 220
rect 192 219 193 220
rect 191 219 192 220
rect 190 219 191 220
rect 189 219 190 220
rect 188 219 189 220
rect 187 219 188 220
rect 186 219 187 220
rect 185 219 186 220
rect 184 219 185 220
rect 183 219 184 220
rect 182 219 183 220
rect 181 219 182 220
rect 145 219 146 220
rect 144 219 145 220
rect 143 219 144 220
rect 142 219 143 220
rect 141 219 142 220
rect 140 219 141 220
rect 139 219 140 220
rect 138 219 139 220
rect 137 219 138 220
rect 136 219 137 220
rect 135 219 136 220
rect 134 219 135 220
rect 133 219 134 220
rect 132 219 133 220
rect 131 219 132 220
rect 130 219 131 220
rect 129 219 130 220
rect 128 219 129 220
rect 127 219 128 220
rect 126 219 127 220
rect 125 219 126 220
rect 124 219 125 220
rect 123 219 124 220
rect 122 219 123 220
rect 121 219 122 220
rect 120 219 121 220
rect 119 219 120 220
rect 118 219 119 220
rect 117 219 118 220
rect 116 219 117 220
rect 115 219 116 220
rect 114 219 115 220
rect 113 219 114 220
rect 112 219 113 220
rect 111 219 112 220
rect 110 219 111 220
rect 109 219 110 220
rect 108 219 109 220
rect 107 219 108 220
rect 106 219 107 220
rect 105 219 106 220
rect 104 219 105 220
rect 103 219 104 220
rect 102 219 103 220
rect 101 219 102 220
rect 70 219 71 220
rect 69 219 70 220
rect 68 219 69 220
rect 67 219 68 220
rect 66 219 67 220
rect 65 219 66 220
rect 64 219 65 220
rect 63 219 64 220
rect 62 219 63 220
rect 61 219 62 220
rect 60 219 61 220
rect 59 219 60 220
rect 58 219 59 220
rect 57 219 58 220
rect 56 219 57 220
rect 55 219 56 220
rect 54 219 55 220
rect 53 219 54 220
rect 52 219 53 220
rect 51 219 52 220
rect 50 219 51 220
rect 49 219 50 220
rect 48 219 49 220
rect 47 219 48 220
rect 46 219 47 220
rect 45 219 46 220
rect 44 219 45 220
rect 43 219 44 220
rect 42 219 43 220
rect 41 219 42 220
rect 40 219 41 220
rect 39 219 40 220
rect 38 219 39 220
rect 37 219 38 220
rect 36 219 37 220
rect 35 219 36 220
rect 34 219 35 220
rect 33 219 34 220
rect 32 219 33 220
rect 31 219 32 220
rect 30 219 31 220
rect 29 219 30 220
rect 28 219 29 220
rect 27 219 28 220
rect 26 219 27 220
rect 25 219 26 220
rect 24 219 25 220
rect 23 219 24 220
rect 22 219 23 220
rect 21 219 22 220
rect 20 219 21 220
rect 19 219 20 220
rect 18 219 19 220
rect 17 219 18 220
rect 16 219 17 220
rect 15 219 16 220
rect 14 219 15 220
rect 13 219 14 220
rect 12 219 13 220
rect 11 219 12 220
rect 10 219 11 220
rect 9 219 10 220
rect 8 219 9 220
rect 7 219 8 220
rect 480 220 481 221
rect 479 220 480 221
rect 478 220 479 221
rect 477 220 478 221
rect 476 220 477 221
rect 475 220 476 221
rect 474 220 475 221
rect 473 220 474 221
rect 472 220 473 221
rect 471 220 472 221
rect 470 220 471 221
rect 469 220 470 221
rect 468 220 469 221
rect 467 220 468 221
rect 466 220 467 221
rect 465 220 466 221
rect 464 220 465 221
rect 463 220 464 221
rect 462 220 463 221
rect 461 220 462 221
rect 460 220 461 221
rect 438 220 439 221
rect 437 220 438 221
rect 436 220 437 221
rect 435 220 436 221
rect 434 220 435 221
rect 433 220 434 221
rect 432 220 433 221
rect 431 220 432 221
rect 430 220 431 221
rect 429 220 430 221
rect 404 220 405 221
rect 403 220 404 221
rect 402 220 403 221
rect 401 220 402 221
rect 400 220 401 221
rect 399 220 400 221
rect 398 220 399 221
rect 397 220 398 221
rect 361 220 362 221
rect 360 220 361 221
rect 359 220 360 221
rect 358 220 359 221
rect 357 220 358 221
rect 356 220 357 221
rect 355 220 356 221
rect 354 220 355 221
rect 353 220 354 221
rect 352 220 353 221
rect 293 220 294 221
rect 292 220 293 221
rect 291 220 292 221
rect 290 220 291 221
rect 289 220 290 221
rect 288 220 289 221
rect 287 220 288 221
rect 286 220 287 221
rect 285 220 286 221
rect 284 220 285 221
rect 283 220 284 221
rect 282 220 283 221
rect 281 220 282 221
rect 280 220 281 221
rect 279 220 280 221
rect 278 220 279 221
rect 277 220 278 221
rect 276 220 277 221
rect 275 220 276 221
rect 274 220 275 221
rect 273 220 274 221
rect 272 220 273 221
rect 271 220 272 221
rect 270 220 271 221
rect 269 220 270 221
rect 268 220 269 221
rect 267 220 268 221
rect 266 220 267 221
rect 265 220 266 221
rect 264 220 265 221
rect 263 220 264 221
rect 262 220 263 221
rect 261 220 262 221
rect 260 220 261 221
rect 259 220 260 221
rect 258 220 259 221
rect 257 220 258 221
rect 256 220 257 221
rect 255 220 256 221
rect 254 220 255 221
rect 253 220 254 221
rect 252 220 253 221
rect 251 220 252 221
rect 250 220 251 221
rect 249 220 250 221
rect 248 220 249 221
rect 247 220 248 221
rect 246 220 247 221
rect 245 220 246 221
rect 244 220 245 221
rect 243 220 244 221
rect 242 220 243 221
rect 241 220 242 221
rect 240 220 241 221
rect 239 220 240 221
rect 238 220 239 221
rect 237 220 238 221
rect 236 220 237 221
rect 235 220 236 221
rect 234 220 235 221
rect 233 220 234 221
rect 232 220 233 221
rect 231 220 232 221
rect 230 220 231 221
rect 229 220 230 221
rect 228 220 229 221
rect 227 220 228 221
rect 226 220 227 221
rect 225 220 226 221
rect 224 220 225 221
rect 223 220 224 221
rect 222 220 223 221
rect 221 220 222 221
rect 220 220 221 221
rect 219 220 220 221
rect 218 220 219 221
rect 217 220 218 221
rect 216 220 217 221
rect 215 220 216 221
rect 214 220 215 221
rect 213 220 214 221
rect 212 220 213 221
rect 211 220 212 221
rect 210 220 211 221
rect 209 220 210 221
rect 208 220 209 221
rect 207 220 208 221
rect 206 220 207 221
rect 205 220 206 221
rect 204 220 205 221
rect 203 220 204 221
rect 202 220 203 221
rect 201 220 202 221
rect 200 220 201 221
rect 199 220 200 221
rect 198 220 199 221
rect 197 220 198 221
rect 196 220 197 221
rect 195 220 196 221
rect 194 220 195 221
rect 193 220 194 221
rect 192 220 193 221
rect 191 220 192 221
rect 190 220 191 221
rect 189 220 190 221
rect 188 220 189 221
rect 187 220 188 221
rect 186 220 187 221
rect 185 220 186 221
rect 184 220 185 221
rect 183 220 184 221
rect 182 220 183 221
rect 181 220 182 221
rect 180 220 181 221
rect 179 220 180 221
rect 145 220 146 221
rect 144 220 145 221
rect 143 220 144 221
rect 142 220 143 221
rect 141 220 142 221
rect 140 220 141 221
rect 139 220 140 221
rect 138 220 139 221
rect 137 220 138 221
rect 136 220 137 221
rect 135 220 136 221
rect 134 220 135 221
rect 133 220 134 221
rect 132 220 133 221
rect 131 220 132 221
rect 130 220 131 221
rect 129 220 130 221
rect 128 220 129 221
rect 127 220 128 221
rect 126 220 127 221
rect 125 220 126 221
rect 124 220 125 221
rect 123 220 124 221
rect 122 220 123 221
rect 121 220 122 221
rect 120 220 121 221
rect 119 220 120 221
rect 118 220 119 221
rect 117 220 118 221
rect 116 220 117 221
rect 115 220 116 221
rect 114 220 115 221
rect 113 220 114 221
rect 112 220 113 221
rect 111 220 112 221
rect 110 220 111 221
rect 109 220 110 221
rect 108 220 109 221
rect 107 220 108 221
rect 106 220 107 221
rect 105 220 106 221
rect 104 220 105 221
rect 103 220 104 221
rect 71 220 72 221
rect 70 220 71 221
rect 69 220 70 221
rect 68 220 69 221
rect 67 220 68 221
rect 66 220 67 221
rect 65 220 66 221
rect 64 220 65 221
rect 63 220 64 221
rect 62 220 63 221
rect 61 220 62 221
rect 60 220 61 221
rect 59 220 60 221
rect 58 220 59 221
rect 57 220 58 221
rect 56 220 57 221
rect 55 220 56 221
rect 54 220 55 221
rect 53 220 54 221
rect 52 220 53 221
rect 51 220 52 221
rect 50 220 51 221
rect 49 220 50 221
rect 48 220 49 221
rect 47 220 48 221
rect 46 220 47 221
rect 45 220 46 221
rect 44 220 45 221
rect 43 220 44 221
rect 42 220 43 221
rect 41 220 42 221
rect 40 220 41 221
rect 39 220 40 221
rect 38 220 39 221
rect 37 220 38 221
rect 36 220 37 221
rect 35 220 36 221
rect 34 220 35 221
rect 33 220 34 221
rect 32 220 33 221
rect 31 220 32 221
rect 30 220 31 221
rect 29 220 30 221
rect 28 220 29 221
rect 27 220 28 221
rect 26 220 27 221
rect 25 220 26 221
rect 24 220 25 221
rect 23 220 24 221
rect 22 220 23 221
rect 21 220 22 221
rect 20 220 21 221
rect 19 220 20 221
rect 18 220 19 221
rect 17 220 18 221
rect 16 220 17 221
rect 15 220 16 221
rect 14 220 15 221
rect 13 220 14 221
rect 12 220 13 221
rect 11 220 12 221
rect 10 220 11 221
rect 9 220 10 221
rect 8 220 9 221
rect 7 220 8 221
rect 480 221 481 222
rect 479 221 480 222
rect 478 221 479 222
rect 477 221 478 222
rect 476 221 477 222
rect 475 221 476 222
rect 474 221 475 222
rect 473 221 474 222
rect 472 221 473 222
rect 471 221 472 222
rect 470 221 471 222
rect 469 221 470 222
rect 468 221 469 222
rect 467 221 468 222
rect 466 221 467 222
rect 465 221 466 222
rect 464 221 465 222
rect 463 221 464 222
rect 462 221 463 222
rect 461 221 462 222
rect 460 221 461 222
rect 438 221 439 222
rect 437 221 438 222
rect 436 221 437 222
rect 435 221 436 222
rect 434 221 435 222
rect 433 221 434 222
rect 432 221 433 222
rect 431 221 432 222
rect 403 221 404 222
rect 402 221 403 222
rect 401 221 402 222
rect 400 221 401 222
rect 399 221 400 222
rect 398 221 399 222
rect 397 221 398 222
rect 396 221 397 222
rect 361 221 362 222
rect 360 221 361 222
rect 359 221 360 222
rect 358 221 359 222
rect 357 221 358 222
rect 356 221 357 222
rect 355 221 356 222
rect 290 221 291 222
rect 289 221 290 222
rect 288 221 289 222
rect 287 221 288 222
rect 286 221 287 222
rect 285 221 286 222
rect 284 221 285 222
rect 283 221 284 222
rect 282 221 283 222
rect 281 221 282 222
rect 280 221 281 222
rect 279 221 280 222
rect 278 221 279 222
rect 277 221 278 222
rect 276 221 277 222
rect 275 221 276 222
rect 274 221 275 222
rect 273 221 274 222
rect 272 221 273 222
rect 271 221 272 222
rect 270 221 271 222
rect 269 221 270 222
rect 268 221 269 222
rect 267 221 268 222
rect 266 221 267 222
rect 265 221 266 222
rect 264 221 265 222
rect 263 221 264 222
rect 262 221 263 222
rect 261 221 262 222
rect 260 221 261 222
rect 259 221 260 222
rect 258 221 259 222
rect 257 221 258 222
rect 256 221 257 222
rect 255 221 256 222
rect 254 221 255 222
rect 253 221 254 222
rect 252 221 253 222
rect 251 221 252 222
rect 250 221 251 222
rect 249 221 250 222
rect 248 221 249 222
rect 247 221 248 222
rect 246 221 247 222
rect 245 221 246 222
rect 244 221 245 222
rect 243 221 244 222
rect 242 221 243 222
rect 241 221 242 222
rect 240 221 241 222
rect 239 221 240 222
rect 238 221 239 222
rect 237 221 238 222
rect 236 221 237 222
rect 235 221 236 222
rect 234 221 235 222
rect 233 221 234 222
rect 232 221 233 222
rect 231 221 232 222
rect 230 221 231 222
rect 229 221 230 222
rect 228 221 229 222
rect 227 221 228 222
rect 226 221 227 222
rect 225 221 226 222
rect 224 221 225 222
rect 223 221 224 222
rect 222 221 223 222
rect 221 221 222 222
rect 220 221 221 222
rect 219 221 220 222
rect 218 221 219 222
rect 217 221 218 222
rect 216 221 217 222
rect 215 221 216 222
rect 214 221 215 222
rect 213 221 214 222
rect 212 221 213 222
rect 211 221 212 222
rect 210 221 211 222
rect 209 221 210 222
rect 208 221 209 222
rect 207 221 208 222
rect 206 221 207 222
rect 205 221 206 222
rect 204 221 205 222
rect 203 221 204 222
rect 202 221 203 222
rect 201 221 202 222
rect 200 221 201 222
rect 199 221 200 222
rect 198 221 199 222
rect 197 221 198 222
rect 196 221 197 222
rect 195 221 196 222
rect 194 221 195 222
rect 193 221 194 222
rect 192 221 193 222
rect 191 221 192 222
rect 190 221 191 222
rect 189 221 190 222
rect 188 221 189 222
rect 187 221 188 222
rect 186 221 187 222
rect 185 221 186 222
rect 184 221 185 222
rect 183 221 184 222
rect 182 221 183 222
rect 181 221 182 222
rect 180 221 181 222
rect 179 221 180 222
rect 178 221 179 222
rect 177 221 178 222
rect 144 221 145 222
rect 143 221 144 222
rect 142 221 143 222
rect 141 221 142 222
rect 140 221 141 222
rect 139 221 140 222
rect 138 221 139 222
rect 137 221 138 222
rect 136 221 137 222
rect 135 221 136 222
rect 134 221 135 222
rect 133 221 134 222
rect 132 221 133 222
rect 131 221 132 222
rect 130 221 131 222
rect 129 221 130 222
rect 128 221 129 222
rect 127 221 128 222
rect 126 221 127 222
rect 125 221 126 222
rect 124 221 125 222
rect 123 221 124 222
rect 122 221 123 222
rect 121 221 122 222
rect 120 221 121 222
rect 119 221 120 222
rect 118 221 119 222
rect 117 221 118 222
rect 116 221 117 222
rect 115 221 116 222
rect 114 221 115 222
rect 113 221 114 222
rect 112 221 113 222
rect 111 221 112 222
rect 110 221 111 222
rect 109 221 110 222
rect 108 221 109 222
rect 107 221 108 222
rect 106 221 107 222
rect 105 221 106 222
rect 104 221 105 222
rect 72 221 73 222
rect 71 221 72 222
rect 70 221 71 222
rect 69 221 70 222
rect 68 221 69 222
rect 67 221 68 222
rect 66 221 67 222
rect 65 221 66 222
rect 64 221 65 222
rect 63 221 64 222
rect 62 221 63 222
rect 61 221 62 222
rect 60 221 61 222
rect 59 221 60 222
rect 58 221 59 222
rect 57 221 58 222
rect 56 221 57 222
rect 55 221 56 222
rect 54 221 55 222
rect 53 221 54 222
rect 52 221 53 222
rect 51 221 52 222
rect 50 221 51 222
rect 49 221 50 222
rect 48 221 49 222
rect 47 221 48 222
rect 46 221 47 222
rect 45 221 46 222
rect 44 221 45 222
rect 43 221 44 222
rect 42 221 43 222
rect 41 221 42 222
rect 40 221 41 222
rect 39 221 40 222
rect 38 221 39 222
rect 37 221 38 222
rect 36 221 37 222
rect 35 221 36 222
rect 34 221 35 222
rect 33 221 34 222
rect 32 221 33 222
rect 31 221 32 222
rect 30 221 31 222
rect 29 221 30 222
rect 28 221 29 222
rect 27 221 28 222
rect 26 221 27 222
rect 25 221 26 222
rect 24 221 25 222
rect 23 221 24 222
rect 22 221 23 222
rect 21 221 22 222
rect 20 221 21 222
rect 19 221 20 222
rect 18 221 19 222
rect 17 221 18 222
rect 16 221 17 222
rect 15 221 16 222
rect 14 221 15 222
rect 13 221 14 222
rect 12 221 13 222
rect 11 221 12 222
rect 10 221 11 222
rect 9 221 10 222
rect 8 221 9 222
rect 7 221 8 222
rect 480 222 481 223
rect 479 222 480 223
rect 478 222 479 223
rect 477 222 478 223
rect 476 222 477 223
rect 475 222 476 223
rect 474 222 475 223
rect 473 222 474 223
rect 472 222 473 223
rect 471 222 472 223
rect 470 222 471 223
rect 469 222 470 223
rect 468 222 469 223
rect 467 222 468 223
rect 466 222 467 223
rect 465 222 466 223
rect 464 222 465 223
rect 463 222 464 223
rect 462 222 463 223
rect 461 222 462 223
rect 460 222 461 223
rect 439 222 440 223
rect 438 222 439 223
rect 437 222 438 223
rect 436 222 437 223
rect 435 222 436 223
rect 434 222 435 223
rect 433 222 434 223
rect 432 222 433 223
rect 401 222 402 223
rect 400 222 401 223
rect 399 222 400 223
rect 398 222 399 223
rect 397 222 398 223
rect 396 222 397 223
rect 362 222 363 223
rect 361 222 362 223
rect 360 222 361 223
rect 359 222 360 223
rect 358 222 359 223
rect 289 222 290 223
rect 288 222 289 223
rect 287 222 288 223
rect 286 222 287 223
rect 285 222 286 223
rect 284 222 285 223
rect 283 222 284 223
rect 282 222 283 223
rect 281 222 282 223
rect 280 222 281 223
rect 279 222 280 223
rect 278 222 279 223
rect 277 222 278 223
rect 276 222 277 223
rect 275 222 276 223
rect 274 222 275 223
rect 273 222 274 223
rect 272 222 273 223
rect 271 222 272 223
rect 270 222 271 223
rect 269 222 270 223
rect 268 222 269 223
rect 267 222 268 223
rect 266 222 267 223
rect 265 222 266 223
rect 264 222 265 223
rect 263 222 264 223
rect 262 222 263 223
rect 261 222 262 223
rect 260 222 261 223
rect 259 222 260 223
rect 258 222 259 223
rect 257 222 258 223
rect 256 222 257 223
rect 255 222 256 223
rect 254 222 255 223
rect 253 222 254 223
rect 252 222 253 223
rect 251 222 252 223
rect 250 222 251 223
rect 249 222 250 223
rect 248 222 249 223
rect 247 222 248 223
rect 246 222 247 223
rect 245 222 246 223
rect 244 222 245 223
rect 243 222 244 223
rect 242 222 243 223
rect 241 222 242 223
rect 240 222 241 223
rect 239 222 240 223
rect 238 222 239 223
rect 237 222 238 223
rect 236 222 237 223
rect 235 222 236 223
rect 234 222 235 223
rect 233 222 234 223
rect 232 222 233 223
rect 231 222 232 223
rect 230 222 231 223
rect 229 222 230 223
rect 228 222 229 223
rect 227 222 228 223
rect 226 222 227 223
rect 225 222 226 223
rect 224 222 225 223
rect 223 222 224 223
rect 222 222 223 223
rect 221 222 222 223
rect 220 222 221 223
rect 219 222 220 223
rect 218 222 219 223
rect 217 222 218 223
rect 216 222 217 223
rect 215 222 216 223
rect 214 222 215 223
rect 213 222 214 223
rect 212 222 213 223
rect 211 222 212 223
rect 210 222 211 223
rect 209 222 210 223
rect 208 222 209 223
rect 207 222 208 223
rect 206 222 207 223
rect 205 222 206 223
rect 204 222 205 223
rect 203 222 204 223
rect 202 222 203 223
rect 201 222 202 223
rect 200 222 201 223
rect 199 222 200 223
rect 198 222 199 223
rect 197 222 198 223
rect 196 222 197 223
rect 195 222 196 223
rect 194 222 195 223
rect 193 222 194 223
rect 192 222 193 223
rect 191 222 192 223
rect 190 222 191 223
rect 189 222 190 223
rect 188 222 189 223
rect 187 222 188 223
rect 186 222 187 223
rect 185 222 186 223
rect 184 222 185 223
rect 183 222 184 223
rect 182 222 183 223
rect 181 222 182 223
rect 180 222 181 223
rect 179 222 180 223
rect 178 222 179 223
rect 177 222 178 223
rect 176 222 177 223
rect 175 222 176 223
rect 144 222 145 223
rect 143 222 144 223
rect 142 222 143 223
rect 141 222 142 223
rect 140 222 141 223
rect 139 222 140 223
rect 138 222 139 223
rect 137 222 138 223
rect 136 222 137 223
rect 135 222 136 223
rect 134 222 135 223
rect 133 222 134 223
rect 132 222 133 223
rect 131 222 132 223
rect 130 222 131 223
rect 129 222 130 223
rect 128 222 129 223
rect 127 222 128 223
rect 126 222 127 223
rect 125 222 126 223
rect 124 222 125 223
rect 123 222 124 223
rect 122 222 123 223
rect 121 222 122 223
rect 120 222 121 223
rect 119 222 120 223
rect 118 222 119 223
rect 117 222 118 223
rect 116 222 117 223
rect 115 222 116 223
rect 114 222 115 223
rect 113 222 114 223
rect 112 222 113 223
rect 111 222 112 223
rect 110 222 111 223
rect 109 222 110 223
rect 108 222 109 223
rect 107 222 108 223
rect 106 222 107 223
rect 73 222 74 223
rect 72 222 73 223
rect 71 222 72 223
rect 70 222 71 223
rect 69 222 70 223
rect 68 222 69 223
rect 67 222 68 223
rect 66 222 67 223
rect 65 222 66 223
rect 64 222 65 223
rect 63 222 64 223
rect 62 222 63 223
rect 61 222 62 223
rect 60 222 61 223
rect 59 222 60 223
rect 58 222 59 223
rect 57 222 58 223
rect 56 222 57 223
rect 55 222 56 223
rect 54 222 55 223
rect 53 222 54 223
rect 52 222 53 223
rect 51 222 52 223
rect 50 222 51 223
rect 49 222 50 223
rect 48 222 49 223
rect 47 222 48 223
rect 46 222 47 223
rect 45 222 46 223
rect 44 222 45 223
rect 43 222 44 223
rect 42 222 43 223
rect 41 222 42 223
rect 40 222 41 223
rect 39 222 40 223
rect 38 222 39 223
rect 37 222 38 223
rect 36 222 37 223
rect 35 222 36 223
rect 34 222 35 223
rect 33 222 34 223
rect 32 222 33 223
rect 31 222 32 223
rect 30 222 31 223
rect 29 222 30 223
rect 28 222 29 223
rect 27 222 28 223
rect 26 222 27 223
rect 25 222 26 223
rect 24 222 25 223
rect 23 222 24 223
rect 22 222 23 223
rect 21 222 22 223
rect 20 222 21 223
rect 19 222 20 223
rect 18 222 19 223
rect 17 222 18 223
rect 16 222 17 223
rect 15 222 16 223
rect 14 222 15 223
rect 13 222 14 223
rect 12 222 13 223
rect 11 222 12 223
rect 10 222 11 223
rect 9 222 10 223
rect 8 222 9 223
rect 7 222 8 223
rect 6 222 7 223
rect 480 223 481 224
rect 479 223 480 224
rect 471 223 472 224
rect 470 223 471 224
rect 461 223 462 224
rect 460 223 461 224
rect 439 223 440 224
rect 438 223 439 224
rect 437 223 438 224
rect 436 223 437 224
rect 435 223 436 224
rect 434 223 435 224
rect 400 223 401 224
rect 399 223 400 224
rect 398 223 399 224
rect 397 223 398 224
rect 396 223 397 224
rect 362 223 363 224
rect 361 223 362 224
rect 360 223 361 224
rect 287 223 288 224
rect 286 223 287 224
rect 285 223 286 224
rect 284 223 285 224
rect 283 223 284 224
rect 282 223 283 224
rect 281 223 282 224
rect 280 223 281 224
rect 279 223 280 224
rect 278 223 279 224
rect 277 223 278 224
rect 276 223 277 224
rect 275 223 276 224
rect 274 223 275 224
rect 273 223 274 224
rect 272 223 273 224
rect 271 223 272 224
rect 270 223 271 224
rect 269 223 270 224
rect 268 223 269 224
rect 267 223 268 224
rect 266 223 267 224
rect 265 223 266 224
rect 264 223 265 224
rect 263 223 264 224
rect 262 223 263 224
rect 261 223 262 224
rect 260 223 261 224
rect 259 223 260 224
rect 258 223 259 224
rect 257 223 258 224
rect 256 223 257 224
rect 255 223 256 224
rect 254 223 255 224
rect 253 223 254 224
rect 252 223 253 224
rect 251 223 252 224
rect 250 223 251 224
rect 249 223 250 224
rect 248 223 249 224
rect 247 223 248 224
rect 246 223 247 224
rect 245 223 246 224
rect 244 223 245 224
rect 243 223 244 224
rect 242 223 243 224
rect 241 223 242 224
rect 240 223 241 224
rect 239 223 240 224
rect 238 223 239 224
rect 237 223 238 224
rect 236 223 237 224
rect 235 223 236 224
rect 234 223 235 224
rect 233 223 234 224
rect 232 223 233 224
rect 231 223 232 224
rect 230 223 231 224
rect 229 223 230 224
rect 228 223 229 224
rect 227 223 228 224
rect 226 223 227 224
rect 225 223 226 224
rect 224 223 225 224
rect 223 223 224 224
rect 222 223 223 224
rect 221 223 222 224
rect 220 223 221 224
rect 219 223 220 224
rect 218 223 219 224
rect 217 223 218 224
rect 216 223 217 224
rect 215 223 216 224
rect 214 223 215 224
rect 213 223 214 224
rect 212 223 213 224
rect 211 223 212 224
rect 210 223 211 224
rect 209 223 210 224
rect 208 223 209 224
rect 207 223 208 224
rect 206 223 207 224
rect 205 223 206 224
rect 204 223 205 224
rect 203 223 204 224
rect 202 223 203 224
rect 201 223 202 224
rect 200 223 201 224
rect 199 223 200 224
rect 198 223 199 224
rect 197 223 198 224
rect 196 223 197 224
rect 195 223 196 224
rect 194 223 195 224
rect 193 223 194 224
rect 192 223 193 224
rect 191 223 192 224
rect 190 223 191 224
rect 189 223 190 224
rect 188 223 189 224
rect 187 223 188 224
rect 186 223 187 224
rect 185 223 186 224
rect 184 223 185 224
rect 183 223 184 224
rect 182 223 183 224
rect 181 223 182 224
rect 180 223 181 224
rect 179 223 180 224
rect 178 223 179 224
rect 177 223 178 224
rect 176 223 177 224
rect 175 223 176 224
rect 174 223 175 224
rect 173 223 174 224
rect 144 223 145 224
rect 143 223 144 224
rect 142 223 143 224
rect 141 223 142 224
rect 140 223 141 224
rect 139 223 140 224
rect 138 223 139 224
rect 137 223 138 224
rect 136 223 137 224
rect 135 223 136 224
rect 134 223 135 224
rect 133 223 134 224
rect 132 223 133 224
rect 131 223 132 224
rect 130 223 131 224
rect 129 223 130 224
rect 128 223 129 224
rect 127 223 128 224
rect 126 223 127 224
rect 125 223 126 224
rect 124 223 125 224
rect 123 223 124 224
rect 122 223 123 224
rect 121 223 122 224
rect 120 223 121 224
rect 119 223 120 224
rect 118 223 119 224
rect 117 223 118 224
rect 116 223 117 224
rect 115 223 116 224
rect 114 223 115 224
rect 113 223 114 224
rect 112 223 113 224
rect 111 223 112 224
rect 110 223 111 224
rect 109 223 110 224
rect 108 223 109 224
rect 107 223 108 224
rect 75 223 76 224
rect 74 223 75 224
rect 73 223 74 224
rect 72 223 73 224
rect 71 223 72 224
rect 70 223 71 224
rect 69 223 70 224
rect 68 223 69 224
rect 67 223 68 224
rect 66 223 67 224
rect 65 223 66 224
rect 64 223 65 224
rect 63 223 64 224
rect 62 223 63 224
rect 61 223 62 224
rect 60 223 61 224
rect 59 223 60 224
rect 58 223 59 224
rect 57 223 58 224
rect 56 223 57 224
rect 55 223 56 224
rect 54 223 55 224
rect 53 223 54 224
rect 52 223 53 224
rect 51 223 52 224
rect 50 223 51 224
rect 49 223 50 224
rect 48 223 49 224
rect 47 223 48 224
rect 46 223 47 224
rect 45 223 46 224
rect 44 223 45 224
rect 43 223 44 224
rect 42 223 43 224
rect 41 223 42 224
rect 40 223 41 224
rect 39 223 40 224
rect 38 223 39 224
rect 37 223 38 224
rect 36 223 37 224
rect 35 223 36 224
rect 34 223 35 224
rect 33 223 34 224
rect 32 223 33 224
rect 31 223 32 224
rect 30 223 31 224
rect 29 223 30 224
rect 28 223 29 224
rect 27 223 28 224
rect 26 223 27 224
rect 25 223 26 224
rect 24 223 25 224
rect 23 223 24 224
rect 22 223 23 224
rect 21 223 22 224
rect 20 223 21 224
rect 19 223 20 224
rect 18 223 19 224
rect 17 223 18 224
rect 16 223 17 224
rect 15 223 16 224
rect 14 223 15 224
rect 13 223 14 224
rect 12 223 13 224
rect 11 223 12 224
rect 10 223 11 224
rect 9 223 10 224
rect 8 223 9 224
rect 7 223 8 224
rect 6 223 7 224
rect 480 224 481 225
rect 471 224 472 225
rect 460 224 461 225
rect 439 224 440 225
rect 438 224 439 225
rect 437 224 438 225
rect 436 224 437 225
rect 435 224 436 225
rect 399 224 400 225
rect 398 224 399 225
rect 397 224 398 225
rect 396 224 397 225
rect 395 224 396 225
rect 362 224 363 225
rect 285 224 286 225
rect 284 224 285 225
rect 283 224 284 225
rect 282 224 283 225
rect 281 224 282 225
rect 280 224 281 225
rect 279 224 280 225
rect 278 224 279 225
rect 277 224 278 225
rect 276 224 277 225
rect 275 224 276 225
rect 274 224 275 225
rect 273 224 274 225
rect 272 224 273 225
rect 271 224 272 225
rect 270 224 271 225
rect 269 224 270 225
rect 268 224 269 225
rect 267 224 268 225
rect 266 224 267 225
rect 265 224 266 225
rect 264 224 265 225
rect 263 224 264 225
rect 262 224 263 225
rect 261 224 262 225
rect 260 224 261 225
rect 259 224 260 225
rect 258 224 259 225
rect 257 224 258 225
rect 256 224 257 225
rect 255 224 256 225
rect 254 224 255 225
rect 253 224 254 225
rect 252 224 253 225
rect 251 224 252 225
rect 250 224 251 225
rect 249 224 250 225
rect 248 224 249 225
rect 247 224 248 225
rect 246 224 247 225
rect 245 224 246 225
rect 244 224 245 225
rect 243 224 244 225
rect 242 224 243 225
rect 241 224 242 225
rect 240 224 241 225
rect 239 224 240 225
rect 238 224 239 225
rect 237 224 238 225
rect 236 224 237 225
rect 235 224 236 225
rect 234 224 235 225
rect 233 224 234 225
rect 232 224 233 225
rect 231 224 232 225
rect 230 224 231 225
rect 229 224 230 225
rect 228 224 229 225
rect 227 224 228 225
rect 226 224 227 225
rect 225 224 226 225
rect 224 224 225 225
rect 223 224 224 225
rect 222 224 223 225
rect 221 224 222 225
rect 220 224 221 225
rect 219 224 220 225
rect 218 224 219 225
rect 217 224 218 225
rect 216 224 217 225
rect 215 224 216 225
rect 214 224 215 225
rect 213 224 214 225
rect 212 224 213 225
rect 211 224 212 225
rect 210 224 211 225
rect 209 224 210 225
rect 208 224 209 225
rect 207 224 208 225
rect 206 224 207 225
rect 205 224 206 225
rect 204 224 205 225
rect 203 224 204 225
rect 202 224 203 225
rect 201 224 202 225
rect 200 224 201 225
rect 199 224 200 225
rect 198 224 199 225
rect 197 224 198 225
rect 196 224 197 225
rect 195 224 196 225
rect 194 224 195 225
rect 193 224 194 225
rect 192 224 193 225
rect 191 224 192 225
rect 190 224 191 225
rect 189 224 190 225
rect 188 224 189 225
rect 187 224 188 225
rect 186 224 187 225
rect 185 224 186 225
rect 184 224 185 225
rect 183 224 184 225
rect 182 224 183 225
rect 181 224 182 225
rect 180 224 181 225
rect 179 224 180 225
rect 178 224 179 225
rect 177 224 178 225
rect 176 224 177 225
rect 175 224 176 225
rect 174 224 175 225
rect 173 224 174 225
rect 172 224 173 225
rect 171 224 172 225
rect 144 224 145 225
rect 143 224 144 225
rect 142 224 143 225
rect 141 224 142 225
rect 140 224 141 225
rect 139 224 140 225
rect 138 224 139 225
rect 137 224 138 225
rect 136 224 137 225
rect 135 224 136 225
rect 134 224 135 225
rect 133 224 134 225
rect 132 224 133 225
rect 131 224 132 225
rect 130 224 131 225
rect 129 224 130 225
rect 128 224 129 225
rect 127 224 128 225
rect 126 224 127 225
rect 125 224 126 225
rect 124 224 125 225
rect 123 224 124 225
rect 122 224 123 225
rect 121 224 122 225
rect 120 224 121 225
rect 119 224 120 225
rect 118 224 119 225
rect 117 224 118 225
rect 116 224 117 225
rect 115 224 116 225
rect 114 224 115 225
rect 113 224 114 225
rect 112 224 113 225
rect 111 224 112 225
rect 110 224 111 225
rect 109 224 110 225
rect 76 224 77 225
rect 75 224 76 225
rect 74 224 75 225
rect 73 224 74 225
rect 72 224 73 225
rect 71 224 72 225
rect 70 224 71 225
rect 69 224 70 225
rect 68 224 69 225
rect 67 224 68 225
rect 66 224 67 225
rect 65 224 66 225
rect 64 224 65 225
rect 63 224 64 225
rect 62 224 63 225
rect 61 224 62 225
rect 60 224 61 225
rect 59 224 60 225
rect 58 224 59 225
rect 57 224 58 225
rect 56 224 57 225
rect 55 224 56 225
rect 54 224 55 225
rect 53 224 54 225
rect 52 224 53 225
rect 51 224 52 225
rect 50 224 51 225
rect 49 224 50 225
rect 48 224 49 225
rect 47 224 48 225
rect 46 224 47 225
rect 45 224 46 225
rect 44 224 45 225
rect 43 224 44 225
rect 42 224 43 225
rect 41 224 42 225
rect 40 224 41 225
rect 39 224 40 225
rect 38 224 39 225
rect 37 224 38 225
rect 36 224 37 225
rect 35 224 36 225
rect 34 224 35 225
rect 33 224 34 225
rect 32 224 33 225
rect 31 224 32 225
rect 30 224 31 225
rect 29 224 30 225
rect 28 224 29 225
rect 27 224 28 225
rect 26 224 27 225
rect 25 224 26 225
rect 24 224 25 225
rect 23 224 24 225
rect 22 224 23 225
rect 21 224 22 225
rect 20 224 21 225
rect 19 224 20 225
rect 18 224 19 225
rect 17 224 18 225
rect 16 224 17 225
rect 15 224 16 225
rect 14 224 15 225
rect 13 224 14 225
rect 12 224 13 225
rect 11 224 12 225
rect 10 224 11 225
rect 9 224 10 225
rect 8 224 9 225
rect 7 224 8 225
rect 6 224 7 225
rect 480 225 481 226
rect 472 225 473 226
rect 471 225 472 226
rect 470 225 471 226
rect 460 225 461 226
rect 439 225 440 226
rect 438 225 439 226
rect 437 225 438 226
rect 436 225 437 226
rect 435 225 436 226
rect 399 225 400 226
rect 398 225 399 226
rect 397 225 398 226
rect 396 225 397 226
rect 395 225 396 226
rect 284 225 285 226
rect 283 225 284 226
rect 282 225 283 226
rect 281 225 282 226
rect 280 225 281 226
rect 279 225 280 226
rect 278 225 279 226
rect 277 225 278 226
rect 276 225 277 226
rect 275 225 276 226
rect 274 225 275 226
rect 273 225 274 226
rect 272 225 273 226
rect 271 225 272 226
rect 270 225 271 226
rect 269 225 270 226
rect 268 225 269 226
rect 267 225 268 226
rect 266 225 267 226
rect 265 225 266 226
rect 264 225 265 226
rect 263 225 264 226
rect 262 225 263 226
rect 261 225 262 226
rect 260 225 261 226
rect 259 225 260 226
rect 258 225 259 226
rect 257 225 258 226
rect 256 225 257 226
rect 255 225 256 226
rect 254 225 255 226
rect 253 225 254 226
rect 252 225 253 226
rect 251 225 252 226
rect 250 225 251 226
rect 249 225 250 226
rect 248 225 249 226
rect 247 225 248 226
rect 246 225 247 226
rect 245 225 246 226
rect 244 225 245 226
rect 243 225 244 226
rect 242 225 243 226
rect 241 225 242 226
rect 240 225 241 226
rect 239 225 240 226
rect 238 225 239 226
rect 237 225 238 226
rect 236 225 237 226
rect 235 225 236 226
rect 234 225 235 226
rect 233 225 234 226
rect 232 225 233 226
rect 231 225 232 226
rect 230 225 231 226
rect 229 225 230 226
rect 228 225 229 226
rect 227 225 228 226
rect 226 225 227 226
rect 225 225 226 226
rect 224 225 225 226
rect 223 225 224 226
rect 222 225 223 226
rect 221 225 222 226
rect 220 225 221 226
rect 219 225 220 226
rect 218 225 219 226
rect 217 225 218 226
rect 216 225 217 226
rect 215 225 216 226
rect 214 225 215 226
rect 213 225 214 226
rect 212 225 213 226
rect 211 225 212 226
rect 210 225 211 226
rect 209 225 210 226
rect 208 225 209 226
rect 207 225 208 226
rect 206 225 207 226
rect 205 225 206 226
rect 204 225 205 226
rect 203 225 204 226
rect 202 225 203 226
rect 201 225 202 226
rect 200 225 201 226
rect 199 225 200 226
rect 198 225 199 226
rect 197 225 198 226
rect 196 225 197 226
rect 195 225 196 226
rect 194 225 195 226
rect 193 225 194 226
rect 192 225 193 226
rect 191 225 192 226
rect 190 225 191 226
rect 189 225 190 226
rect 188 225 189 226
rect 187 225 188 226
rect 186 225 187 226
rect 185 225 186 226
rect 184 225 185 226
rect 183 225 184 226
rect 182 225 183 226
rect 181 225 182 226
rect 180 225 181 226
rect 179 225 180 226
rect 178 225 179 226
rect 177 225 178 226
rect 176 225 177 226
rect 175 225 176 226
rect 174 225 175 226
rect 173 225 174 226
rect 172 225 173 226
rect 171 225 172 226
rect 170 225 171 226
rect 169 225 170 226
rect 144 225 145 226
rect 143 225 144 226
rect 142 225 143 226
rect 141 225 142 226
rect 140 225 141 226
rect 139 225 140 226
rect 138 225 139 226
rect 137 225 138 226
rect 136 225 137 226
rect 135 225 136 226
rect 134 225 135 226
rect 133 225 134 226
rect 132 225 133 226
rect 131 225 132 226
rect 130 225 131 226
rect 129 225 130 226
rect 128 225 129 226
rect 127 225 128 226
rect 126 225 127 226
rect 125 225 126 226
rect 124 225 125 226
rect 123 225 124 226
rect 122 225 123 226
rect 121 225 122 226
rect 120 225 121 226
rect 119 225 120 226
rect 118 225 119 226
rect 117 225 118 226
rect 116 225 117 226
rect 115 225 116 226
rect 114 225 115 226
rect 113 225 114 226
rect 112 225 113 226
rect 111 225 112 226
rect 110 225 111 226
rect 77 225 78 226
rect 76 225 77 226
rect 75 225 76 226
rect 74 225 75 226
rect 73 225 74 226
rect 72 225 73 226
rect 71 225 72 226
rect 70 225 71 226
rect 69 225 70 226
rect 68 225 69 226
rect 67 225 68 226
rect 66 225 67 226
rect 65 225 66 226
rect 64 225 65 226
rect 63 225 64 226
rect 62 225 63 226
rect 61 225 62 226
rect 60 225 61 226
rect 59 225 60 226
rect 58 225 59 226
rect 57 225 58 226
rect 56 225 57 226
rect 55 225 56 226
rect 54 225 55 226
rect 53 225 54 226
rect 52 225 53 226
rect 51 225 52 226
rect 50 225 51 226
rect 49 225 50 226
rect 48 225 49 226
rect 47 225 48 226
rect 46 225 47 226
rect 45 225 46 226
rect 44 225 45 226
rect 43 225 44 226
rect 42 225 43 226
rect 41 225 42 226
rect 40 225 41 226
rect 39 225 40 226
rect 38 225 39 226
rect 37 225 38 226
rect 36 225 37 226
rect 35 225 36 226
rect 34 225 35 226
rect 33 225 34 226
rect 32 225 33 226
rect 31 225 32 226
rect 30 225 31 226
rect 29 225 30 226
rect 28 225 29 226
rect 27 225 28 226
rect 26 225 27 226
rect 25 225 26 226
rect 24 225 25 226
rect 23 225 24 226
rect 22 225 23 226
rect 21 225 22 226
rect 20 225 21 226
rect 19 225 20 226
rect 18 225 19 226
rect 17 225 18 226
rect 16 225 17 226
rect 15 225 16 226
rect 14 225 15 226
rect 13 225 14 226
rect 12 225 13 226
rect 11 225 12 226
rect 10 225 11 226
rect 9 225 10 226
rect 8 225 9 226
rect 7 225 8 226
rect 6 225 7 226
rect 474 226 475 227
rect 473 226 474 227
rect 472 226 473 227
rect 471 226 472 227
rect 470 226 471 227
rect 461 226 462 227
rect 460 226 461 227
rect 440 226 441 227
rect 439 226 440 227
rect 438 226 439 227
rect 437 226 438 227
rect 436 226 437 227
rect 398 226 399 227
rect 397 226 398 227
rect 396 226 397 227
rect 395 226 396 227
rect 282 226 283 227
rect 281 226 282 227
rect 280 226 281 227
rect 279 226 280 227
rect 278 226 279 227
rect 277 226 278 227
rect 276 226 277 227
rect 275 226 276 227
rect 274 226 275 227
rect 273 226 274 227
rect 272 226 273 227
rect 271 226 272 227
rect 270 226 271 227
rect 269 226 270 227
rect 268 226 269 227
rect 267 226 268 227
rect 266 226 267 227
rect 265 226 266 227
rect 264 226 265 227
rect 263 226 264 227
rect 262 226 263 227
rect 261 226 262 227
rect 260 226 261 227
rect 259 226 260 227
rect 258 226 259 227
rect 257 226 258 227
rect 256 226 257 227
rect 255 226 256 227
rect 254 226 255 227
rect 253 226 254 227
rect 252 226 253 227
rect 251 226 252 227
rect 250 226 251 227
rect 249 226 250 227
rect 248 226 249 227
rect 247 226 248 227
rect 246 226 247 227
rect 245 226 246 227
rect 244 226 245 227
rect 243 226 244 227
rect 242 226 243 227
rect 241 226 242 227
rect 240 226 241 227
rect 239 226 240 227
rect 238 226 239 227
rect 237 226 238 227
rect 236 226 237 227
rect 235 226 236 227
rect 234 226 235 227
rect 233 226 234 227
rect 232 226 233 227
rect 231 226 232 227
rect 230 226 231 227
rect 229 226 230 227
rect 228 226 229 227
rect 227 226 228 227
rect 226 226 227 227
rect 225 226 226 227
rect 224 226 225 227
rect 223 226 224 227
rect 222 226 223 227
rect 221 226 222 227
rect 220 226 221 227
rect 219 226 220 227
rect 218 226 219 227
rect 217 226 218 227
rect 216 226 217 227
rect 215 226 216 227
rect 214 226 215 227
rect 213 226 214 227
rect 212 226 213 227
rect 211 226 212 227
rect 210 226 211 227
rect 209 226 210 227
rect 208 226 209 227
rect 207 226 208 227
rect 206 226 207 227
rect 205 226 206 227
rect 204 226 205 227
rect 203 226 204 227
rect 202 226 203 227
rect 201 226 202 227
rect 200 226 201 227
rect 199 226 200 227
rect 198 226 199 227
rect 197 226 198 227
rect 196 226 197 227
rect 195 226 196 227
rect 194 226 195 227
rect 193 226 194 227
rect 192 226 193 227
rect 191 226 192 227
rect 190 226 191 227
rect 189 226 190 227
rect 188 226 189 227
rect 187 226 188 227
rect 186 226 187 227
rect 185 226 186 227
rect 184 226 185 227
rect 183 226 184 227
rect 182 226 183 227
rect 181 226 182 227
rect 180 226 181 227
rect 179 226 180 227
rect 178 226 179 227
rect 177 226 178 227
rect 176 226 177 227
rect 175 226 176 227
rect 174 226 175 227
rect 173 226 174 227
rect 172 226 173 227
rect 171 226 172 227
rect 170 226 171 227
rect 169 226 170 227
rect 168 226 169 227
rect 167 226 168 227
rect 144 226 145 227
rect 143 226 144 227
rect 142 226 143 227
rect 141 226 142 227
rect 140 226 141 227
rect 139 226 140 227
rect 138 226 139 227
rect 137 226 138 227
rect 136 226 137 227
rect 135 226 136 227
rect 134 226 135 227
rect 133 226 134 227
rect 132 226 133 227
rect 131 226 132 227
rect 130 226 131 227
rect 129 226 130 227
rect 128 226 129 227
rect 127 226 128 227
rect 126 226 127 227
rect 125 226 126 227
rect 124 226 125 227
rect 123 226 124 227
rect 122 226 123 227
rect 121 226 122 227
rect 120 226 121 227
rect 119 226 120 227
rect 118 226 119 227
rect 117 226 118 227
rect 116 226 117 227
rect 115 226 116 227
rect 114 226 115 227
rect 113 226 114 227
rect 112 226 113 227
rect 111 226 112 227
rect 79 226 80 227
rect 78 226 79 227
rect 77 226 78 227
rect 76 226 77 227
rect 75 226 76 227
rect 74 226 75 227
rect 73 226 74 227
rect 72 226 73 227
rect 71 226 72 227
rect 70 226 71 227
rect 69 226 70 227
rect 68 226 69 227
rect 67 226 68 227
rect 66 226 67 227
rect 65 226 66 227
rect 64 226 65 227
rect 63 226 64 227
rect 62 226 63 227
rect 61 226 62 227
rect 60 226 61 227
rect 59 226 60 227
rect 58 226 59 227
rect 57 226 58 227
rect 56 226 57 227
rect 55 226 56 227
rect 54 226 55 227
rect 53 226 54 227
rect 52 226 53 227
rect 51 226 52 227
rect 50 226 51 227
rect 49 226 50 227
rect 48 226 49 227
rect 47 226 48 227
rect 46 226 47 227
rect 45 226 46 227
rect 44 226 45 227
rect 43 226 44 227
rect 42 226 43 227
rect 41 226 42 227
rect 40 226 41 227
rect 39 226 40 227
rect 38 226 39 227
rect 37 226 38 227
rect 36 226 37 227
rect 35 226 36 227
rect 34 226 35 227
rect 33 226 34 227
rect 32 226 33 227
rect 31 226 32 227
rect 30 226 31 227
rect 29 226 30 227
rect 28 226 29 227
rect 27 226 28 227
rect 26 226 27 227
rect 25 226 26 227
rect 24 226 25 227
rect 23 226 24 227
rect 22 226 23 227
rect 21 226 22 227
rect 20 226 21 227
rect 19 226 20 227
rect 18 226 19 227
rect 17 226 18 227
rect 16 226 17 227
rect 15 226 16 227
rect 14 226 15 227
rect 13 226 14 227
rect 12 226 13 227
rect 11 226 12 227
rect 10 226 11 227
rect 9 226 10 227
rect 8 226 9 227
rect 7 226 8 227
rect 6 226 7 227
rect 5 226 6 227
rect 476 227 477 228
rect 475 227 476 228
rect 474 227 475 228
rect 473 227 474 228
rect 472 227 473 228
rect 471 227 472 228
rect 470 227 471 228
rect 469 227 470 228
rect 461 227 462 228
rect 460 227 461 228
rect 440 227 441 228
rect 439 227 440 228
rect 438 227 439 228
rect 437 227 438 228
rect 397 227 398 228
rect 396 227 397 228
rect 395 227 396 228
rect 281 227 282 228
rect 280 227 281 228
rect 279 227 280 228
rect 278 227 279 228
rect 277 227 278 228
rect 276 227 277 228
rect 275 227 276 228
rect 274 227 275 228
rect 273 227 274 228
rect 272 227 273 228
rect 271 227 272 228
rect 270 227 271 228
rect 269 227 270 228
rect 268 227 269 228
rect 267 227 268 228
rect 266 227 267 228
rect 265 227 266 228
rect 264 227 265 228
rect 263 227 264 228
rect 262 227 263 228
rect 261 227 262 228
rect 260 227 261 228
rect 259 227 260 228
rect 258 227 259 228
rect 257 227 258 228
rect 256 227 257 228
rect 255 227 256 228
rect 254 227 255 228
rect 253 227 254 228
rect 252 227 253 228
rect 251 227 252 228
rect 250 227 251 228
rect 249 227 250 228
rect 248 227 249 228
rect 247 227 248 228
rect 246 227 247 228
rect 245 227 246 228
rect 244 227 245 228
rect 243 227 244 228
rect 242 227 243 228
rect 241 227 242 228
rect 240 227 241 228
rect 239 227 240 228
rect 238 227 239 228
rect 237 227 238 228
rect 236 227 237 228
rect 235 227 236 228
rect 234 227 235 228
rect 233 227 234 228
rect 232 227 233 228
rect 231 227 232 228
rect 230 227 231 228
rect 229 227 230 228
rect 228 227 229 228
rect 227 227 228 228
rect 226 227 227 228
rect 225 227 226 228
rect 224 227 225 228
rect 223 227 224 228
rect 222 227 223 228
rect 221 227 222 228
rect 220 227 221 228
rect 219 227 220 228
rect 218 227 219 228
rect 217 227 218 228
rect 216 227 217 228
rect 215 227 216 228
rect 214 227 215 228
rect 213 227 214 228
rect 212 227 213 228
rect 211 227 212 228
rect 210 227 211 228
rect 209 227 210 228
rect 208 227 209 228
rect 207 227 208 228
rect 206 227 207 228
rect 205 227 206 228
rect 204 227 205 228
rect 203 227 204 228
rect 202 227 203 228
rect 201 227 202 228
rect 200 227 201 228
rect 199 227 200 228
rect 198 227 199 228
rect 197 227 198 228
rect 196 227 197 228
rect 195 227 196 228
rect 194 227 195 228
rect 193 227 194 228
rect 192 227 193 228
rect 191 227 192 228
rect 190 227 191 228
rect 189 227 190 228
rect 188 227 189 228
rect 187 227 188 228
rect 186 227 187 228
rect 185 227 186 228
rect 184 227 185 228
rect 183 227 184 228
rect 182 227 183 228
rect 181 227 182 228
rect 180 227 181 228
rect 179 227 180 228
rect 178 227 179 228
rect 177 227 178 228
rect 176 227 177 228
rect 175 227 176 228
rect 174 227 175 228
rect 173 227 174 228
rect 172 227 173 228
rect 171 227 172 228
rect 170 227 171 228
rect 169 227 170 228
rect 168 227 169 228
rect 167 227 168 228
rect 166 227 167 228
rect 165 227 166 228
rect 164 227 165 228
rect 144 227 145 228
rect 143 227 144 228
rect 142 227 143 228
rect 141 227 142 228
rect 140 227 141 228
rect 139 227 140 228
rect 138 227 139 228
rect 137 227 138 228
rect 136 227 137 228
rect 135 227 136 228
rect 134 227 135 228
rect 133 227 134 228
rect 132 227 133 228
rect 131 227 132 228
rect 130 227 131 228
rect 129 227 130 228
rect 128 227 129 228
rect 127 227 128 228
rect 126 227 127 228
rect 125 227 126 228
rect 124 227 125 228
rect 123 227 124 228
rect 122 227 123 228
rect 121 227 122 228
rect 120 227 121 228
rect 119 227 120 228
rect 118 227 119 228
rect 117 227 118 228
rect 116 227 117 228
rect 115 227 116 228
rect 114 227 115 228
rect 113 227 114 228
rect 112 227 113 228
rect 80 227 81 228
rect 79 227 80 228
rect 78 227 79 228
rect 77 227 78 228
rect 76 227 77 228
rect 75 227 76 228
rect 74 227 75 228
rect 73 227 74 228
rect 72 227 73 228
rect 71 227 72 228
rect 70 227 71 228
rect 69 227 70 228
rect 68 227 69 228
rect 67 227 68 228
rect 66 227 67 228
rect 65 227 66 228
rect 64 227 65 228
rect 63 227 64 228
rect 62 227 63 228
rect 61 227 62 228
rect 60 227 61 228
rect 59 227 60 228
rect 58 227 59 228
rect 57 227 58 228
rect 56 227 57 228
rect 55 227 56 228
rect 54 227 55 228
rect 53 227 54 228
rect 52 227 53 228
rect 51 227 52 228
rect 50 227 51 228
rect 49 227 50 228
rect 48 227 49 228
rect 47 227 48 228
rect 46 227 47 228
rect 45 227 46 228
rect 44 227 45 228
rect 43 227 44 228
rect 42 227 43 228
rect 41 227 42 228
rect 40 227 41 228
rect 39 227 40 228
rect 38 227 39 228
rect 37 227 38 228
rect 36 227 37 228
rect 35 227 36 228
rect 34 227 35 228
rect 33 227 34 228
rect 32 227 33 228
rect 31 227 32 228
rect 30 227 31 228
rect 29 227 30 228
rect 28 227 29 228
rect 27 227 28 228
rect 26 227 27 228
rect 25 227 26 228
rect 24 227 25 228
rect 23 227 24 228
rect 22 227 23 228
rect 21 227 22 228
rect 20 227 21 228
rect 19 227 20 228
rect 18 227 19 228
rect 17 227 18 228
rect 16 227 17 228
rect 15 227 16 228
rect 14 227 15 228
rect 13 227 14 228
rect 12 227 13 228
rect 11 227 12 228
rect 10 227 11 228
rect 9 227 10 228
rect 8 227 9 228
rect 7 227 8 228
rect 6 227 7 228
rect 5 227 6 228
rect 478 228 479 229
rect 477 228 478 229
rect 476 228 477 229
rect 475 228 476 229
rect 474 228 475 229
rect 473 228 474 229
rect 472 228 473 229
rect 471 228 472 229
rect 470 228 471 229
rect 469 228 470 229
rect 468 228 469 229
rect 467 228 468 229
rect 464 228 465 229
rect 463 228 464 229
rect 462 228 463 229
rect 461 228 462 229
rect 460 228 461 229
rect 440 228 441 229
rect 439 228 440 229
rect 438 228 439 229
rect 437 228 438 229
rect 397 228 398 229
rect 396 228 397 229
rect 395 228 396 229
rect 394 228 395 229
rect 280 228 281 229
rect 279 228 280 229
rect 278 228 279 229
rect 277 228 278 229
rect 276 228 277 229
rect 275 228 276 229
rect 274 228 275 229
rect 273 228 274 229
rect 272 228 273 229
rect 271 228 272 229
rect 270 228 271 229
rect 269 228 270 229
rect 268 228 269 229
rect 267 228 268 229
rect 266 228 267 229
rect 265 228 266 229
rect 264 228 265 229
rect 263 228 264 229
rect 262 228 263 229
rect 261 228 262 229
rect 260 228 261 229
rect 259 228 260 229
rect 258 228 259 229
rect 257 228 258 229
rect 256 228 257 229
rect 255 228 256 229
rect 254 228 255 229
rect 253 228 254 229
rect 252 228 253 229
rect 251 228 252 229
rect 250 228 251 229
rect 249 228 250 229
rect 248 228 249 229
rect 247 228 248 229
rect 246 228 247 229
rect 245 228 246 229
rect 244 228 245 229
rect 243 228 244 229
rect 242 228 243 229
rect 241 228 242 229
rect 240 228 241 229
rect 239 228 240 229
rect 238 228 239 229
rect 237 228 238 229
rect 236 228 237 229
rect 235 228 236 229
rect 234 228 235 229
rect 233 228 234 229
rect 232 228 233 229
rect 231 228 232 229
rect 230 228 231 229
rect 229 228 230 229
rect 228 228 229 229
rect 227 228 228 229
rect 226 228 227 229
rect 225 228 226 229
rect 224 228 225 229
rect 223 228 224 229
rect 222 228 223 229
rect 221 228 222 229
rect 220 228 221 229
rect 219 228 220 229
rect 218 228 219 229
rect 217 228 218 229
rect 216 228 217 229
rect 215 228 216 229
rect 214 228 215 229
rect 213 228 214 229
rect 212 228 213 229
rect 211 228 212 229
rect 210 228 211 229
rect 209 228 210 229
rect 208 228 209 229
rect 207 228 208 229
rect 206 228 207 229
rect 205 228 206 229
rect 204 228 205 229
rect 203 228 204 229
rect 202 228 203 229
rect 201 228 202 229
rect 200 228 201 229
rect 199 228 200 229
rect 198 228 199 229
rect 197 228 198 229
rect 196 228 197 229
rect 195 228 196 229
rect 194 228 195 229
rect 193 228 194 229
rect 192 228 193 229
rect 191 228 192 229
rect 190 228 191 229
rect 189 228 190 229
rect 188 228 189 229
rect 187 228 188 229
rect 186 228 187 229
rect 185 228 186 229
rect 184 228 185 229
rect 183 228 184 229
rect 182 228 183 229
rect 181 228 182 229
rect 180 228 181 229
rect 179 228 180 229
rect 178 228 179 229
rect 177 228 178 229
rect 176 228 177 229
rect 175 228 176 229
rect 174 228 175 229
rect 173 228 174 229
rect 172 228 173 229
rect 171 228 172 229
rect 170 228 171 229
rect 169 228 170 229
rect 168 228 169 229
rect 167 228 168 229
rect 166 228 167 229
rect 165 228 166 229
rect 164 228 165 229
rect 163 228 164 229
rect 162 228 163 229
rect 144 228 145 229
rect 143 228 144 229
rect 142 228 143 229
rect 141 228 142 229
rect 140 228 141 229
rect 139 228 140 229
rect 138 228 139 229
rect 137 228 138 229
rect 136 228 137 229
rect 135 228 136 229
rect 134 228 135 229
rect 133 228 134 229
rect 132 228 133 229
rect 131 228 132 229
rect 130 228 131 229
rect 129 228 130 229
rect 128 228 129 229
rect 127 228 128 229
rect 126 228 127 229
rect 125 228 126 229
rect 124 228 125 229
rect 123 228 124 229
rect 122 228 123 229
rect 121 228 122 229
rect 120 228 121 229
rect 119 228 120 229
rect 118 228 119 229
rect 117 228 118 229
rect 116 228 117 229
rect 115 228 116 229
rect 114 228 115 229
rect 113 228 114 229
rect 112 228 113 229
rect 82 228 83 229
rect 81 228 82 229
rect 80 228 81 229
rect 79 228 80 229
rect 78 228 79 229
rect 77 228 78 229
rect 76 228 77 229
rect 75 228 76 229
rect 74 228 75 229
rect 73 228 74 229
rect 72 228 73 229
rect 71 228 72 229
rect 70 228 71 229
rect 69 228 70 229
rect 68 228 69 229
rect 67 228 68 229
rect 66 228 67 229
rect 65 228 66 229
rect 64 228 65 229
rect 63 228 64 229
rect 62 228 63 229
rect 61 228 62 229
rect 60 228 61 229
rect 59 228 60 229
rect 58 228 59 229
rect 57 228 58 229
rect 56 228 57 229
rect 55 228 56 229
rect 54 228 55 229
rect 53 228 54 229
rect 52 228 53 229
rect 51 228 52 229
rect 50 228 51 229
rect 49 228 50 229
rect 48 228 49 229
rect 47 228 48 229
rect 46 228 47 229
rect 45 228 46 229
rect 44 228 45 229
rect 43 228 44 229
rect 42 228 43 229
rect 41 228 42 229
rect 40 228 41 229
rect 39 228 40 229
rect 38 228 39 229
rect 37 228 38 229
rect 36 228 37 229
rect 35 228 36 229
rect 34 228 35 229
rect 33 228 34 229
rect 32 228 33 229
rect 31 228 32 229
rect 30 228 31 229
rect 29 228 30 229
rect 28 228 29 229
rect 27 228 28 229
rect 26 228 27 229
rect 25 228 26 229
rect 24 228 25 229
rect 23 228 24 229
rect 22 228 23 229
rect 21 228 22 229
rect 20 228 21 229
rect 19 228 20 229
rect 18 228 19 229
rect 17 228 18 229
rect 16 228 17 229
rect 15 228 16 229
rect 14 228 15 229
rect 13 228 14 229
rect 12 228 13 229
rect 11 228 12 229
rect 10 228 11 229
rect 9 228 10 229
rect 8 228 9 229
rect 7 228 8 229
rect 6 228 7 229
rect 5 228 6 229
rect 479 229 480 230
rect 478 229 479 230
rect 477 229 478 230
rect 476 229 477 230
rect 475 229 476 230
rect 474 229 475 230
rect 473 229 474 230
rect 472 229 473 230
rect 471 229 472 230
rect 470 229 471 230
rect 469 229 470 230
rect 468 229 469 230
rect 467 229 468 230
rect 466 229 467 230
rect 465 229 466 230
rect 464 229 465 230
rect 463 229 464 230
rect 462 229 463 230
rect 461 229 462 230
rect 460 229 461 230
rect 440 229 441 230
rect 439 229 440 230
rect 438 229 439 230
rect 437 229 438 230
rect 397 229 398 230
rect 396 229 397 230
rect 395 229 396 230
rect 394 229 395 230
rect 278 229 279 230
rect 277 229 278 230
rect 276 229 277 230
rect 275 229 276 230
rect 274 229 275 230
rect 273 229 274 230
rect 272 229 273 230
rect 271 229 272 230
rect 270 229 271 230
rect 269 229 270 230
rect 268 229 269 230
rect 267 229 268 230
rect 266 229 267 230
rect 265 229 266 230
rect 264 229 265 230
rect 263 229 264 230
rect 262 229 263 230
rect 261 229 262 230
rect 260 229 261 230
rect 259 229 260 230
rect 258 229 259 230
rect 257 229 258 230
rect 256 229 257 230
rect 255 229 256 230
rect 254 229 255 230
rect 253 229 254 230
rect 252 229 253 230
rect 251 229 252 230
rect 250 229 251 230
rect 249 229 250 230
rect 248 229 249 230
rect 247 229 248 230
rect 246 229 247 230
rect 245 229 246 230
rect 244 229 245 230
rect 243 229 244 230
rect 242 229 243 230
rect 241 229 242 230
rect 240 229 241 230
rect 239 229 240 230
rect 238 229 239 230
rect 237 229 238 230
rect 236 229 237 230
rect 235 229 236 230
rect 234 229 235 230
rect 233 229 234 230
rect 232 229 233 230
rect 231 229 232 230
rect 230 229 231 230
rect 229 229 230 230
rect 228 229 229 230
rect 227 229 228 230
rect 226 229 227 230
rect 225 229 226 230
rect 224 229 225 230
rect 223 229 224 230
rect 222 229 223 230
rect 221 229 222 230
rect 220 229 221 230
rect 219 229 220 230
rect 218 229 219 230
rect 217 229 218 230
rect 216 229 217 230
rect 215 229 216 230
rect 214 229 215 230
rect 213 229 214 230
rect 212 229 213 230
rect 211 229 212 230
rect 210 229 211 230
rect 209 229 210 230
rect 208 229 209 230
rect 207 229 208 230
rect 206 229 207 230
rect 205 229 206 230
rect 204 229 205 230
rect 203 229 204 230
rect 202 229 203 230
rect 201 229 202 230
rect 200 229 201 230
rect 199 229 200 230
rect 198 229 199 230
rect 197 229 198 230
rect 196 229 197 230
rect 195 229 196 230
rect 194 229 195 230
rect 193 229 194 230
rect 192 229 193 230
rect 191 229 192 230
rect 190 229 191 230
rect 189 229 190 230
rect 188 229 189 230
rect 187 229 188 230
rect 186 229 187 230
rect 185 229 186 230
rect 184 229 185 230
rect 183 229 184 230
rect 182 229 183 230
rect 181 229 182 230
rect 180 229 181 230
rect 179 229 180 230
rect 178 229 179 230
rect 177 229 178 230
rect 176 229 177 230
rect 175 229 176 230
rect 174 229 175 230
rect 173 229 174 230
rect 172 229 173 230
rect 171 229 172 230
rect 170 229 171 230
rect 169 229 170 230
rect 168 229 169 230
rect 167 229 168 230
rect 166 229 167 230
rect 165 229 166 230
rect 164 229 165 230
rect 163 229 164 230
rect 162 229 163 230
rect 144 229 145 230
rect 143 229 144 230
rect 142 229 143 230
rect 141 229 142 230
rect 140 229 141 230
rect 139 229 140 230
rect 138 229 139 230
rect 137 229 138 230
rect 136 229 137 230
rect 135 229 136 230
rect 134 229 135 230
rect 133 229 134 230
rect 132 229 133 230
rect 131 229 132 230
rect 130 229 131 230
rect 129 229 130 230
rect 128 229 129 230
rect 127 229 128 230
rect 126 229 127 230
rect 125 229 126 230
rect 124 229 125 230
rect 123 229 124 230
rect 122 229 123 230
rect 121 229 122 230
rect 120 229 121 230
rect 119 229 120 230
rect 118 229 119 230
rect 117 229 118 230
rect 116 229 117 230
rect 115 229 116 230
rect 114 229 115 230
rect 113 229 114 230
rect 83 229 84 230
rect 82 229 83 230
rect 81 229 82 230
rect 80 229 81 230
rect 79 229 80 230
rect 78 229 79 230
rect 77 229 78 230
rect 76 229 77 230
rect 75 229 76 230
rect 74 229 75 230
rect 73 229 74 230
rect 72 229 73 230
rect 71 229 72 230
rect 70 229 71 230
rect 69 229 70 230
rect 68 229 69 230
rect 67 229 68 230
rect 66 229 67 230
rect 65 229 66 230
rect 64 229 65 230
rect 63 229 64 230
rect 62 229 63 230
rect 61 229 62 230
rect 60 229 61 230
rect 59 229 60 230
rect 58 229 59 230
rect 57 229 58 230
rect 56 229 57 230
rect 55 229 56 230
rect 54 229 55 230
rect 53 229 54 230
rect 52 229 53 230
rect 51 229 52 230
rect 50 229 51 230
rect 49 229 50 230
rect 48 229 49 230
rect 47 229 48 230
rect 46 229 47 230
rect 45 229 46 230
rect 44 229 45 230
rect 43 229 44 230
rect 42 229 43 230
rect 41 229 42 230
rect 40 229 41 230
rect 39 229 40 230
rect 38 229 39 230
rect 37 229 38 230
rect 36 229 37 230
rect 35 229 36 230
rect 34 229 35 230
rect 33 229 34 230
rect 32 229 33 230
rect 31 229 32 230
rect 30 229 31 230
rect 29 229 30 230
rect 28 229 29 230
rect 27 229 28 230
rect 26 229 27 230
rect 25 229 26 230
rect 24 229 25 230
rect 23 229 24 230
rect 22 229 23 230
rect 21 229 22 230
rect 20 229 21 230
rect 19 229 20 230
rect 18 229 19 230
rect 17 229 18 230
rect 16 229 17 230
rect 15 229 16 230
rect 14 229 15 230
rect 13 229 14 230
rect 12 229 13 230
rect 11 229 12 230
rect 10 229 11 230
rect 9 229 10 230
rect 8 229 9 230
rect 7 229 8 230
rect 6 229 7 230
rect 5 229 6 230
rect 480 230 481 231
rect 479 230 480 231
rect 478 230 479 231
rect 477 230 478 231
rect 476 230 477 231
rect 475 230 476 231
rect 474 230 475 231
rect 473 230 474 231
rect 469 230 470 231
rect 468 230 469 231
rect 467 230 468 231
rect 466 230 467 231
rect 465 230 466 231
rect 464 230 465 231
rect 463 230 464 231
rect 462 230 463 231
rect 461 230 462 231
rect 460 230 461 231
rect 440 230 441 231
rect 439 230 440 231
rect 438 230 439 231
rect 396 230 397 231
rect 395 230 396 231
rect 394 230 395 231
rect 277 230 278 231
rect 276 230 277 231
rect 275 230 276 231
rect 274 230 275 231
rect 273 230 274 231
rect 272 230 273 231
rect 271 230 272 231
rect 270 230 271 231
rect 269 230 270 231
rect 268 230 269 231
rect 267 230 268 231
rect 266 230 267 231
rect 265 230 266 231
rect 264 230 265 231
rect 263 230 264 231
rect 262 230 263 231
rect 261 230 262 231
rect 260 230 261 231
rect 259 230 260 231
rect 258 230 259 231
rect 257 230 258 231
rect 256 230 257 231
rect 255 230 256 231
rect 254 230 255 231
rect 253 230 254 231
rect 252 230 253 231
rect 251 230 252 231
rect 250 230 251 231
rect 249 230 250 231
rect 248 230 249 231
rect 247 230 248 231
rect 246 230 247 231
rect 245 230 246 231
rect 244 230 245 231
rect 243 230 244 231
rect 242 230 243 231
rect 241 230 242 231
rect 240 230 241 231
rect 239 230 240 231
rect 238 230 239 231
rect 237 230 238 231
rect 236 230 237 231
rect 235 230 236 231
rect 234 230 235 231
rect 233 230 234 231
rect 232 230 233 231
rect 231 230 232 231
rect 230 230 231 231
rect 229 230 230 231
rect 228 230 229 231
rect 227 230 228 231
rect 226 230 227 231
rect 225 230 226 231
rect 224 230 225 231
rect 223 230 224 231
rect 222 230 223 231
rect 221 230 222 231
rect 220 230 221 231
rect 219 230 220 231
rect 218 230 219 231
rect 217 230 218 231
rect 216 230 217 231
rect 215 230 216 231
rect 214 230 215 231
rect 213 230 214 231
rect 212 230 213 231
rect 211 230 212 231
rect 210 230 211 231
rect 209 230 210 231
rect 208 230 209 231
rect 207 230 208 231
rect 206 230 207 231
rect 205 230 206 231
rect 204 230 205 231
rect 203 230 204 231
rect 202 230 203 231
rect 201 230 202 231
rect 200 230 201 231
rect 199 230 200 231
rect 198 230 199 231
rect 197 230 198 231
rect 196 230 197 231
rect 195 230 196 231
rect 194 230 195 231
rect 193 230 194 231
rect 192 230 193 231
rect 191 230 192 231
rect 190 230 191 231
rect 189 230 190 231
rect 188 230 189 231
rect 187 230 188 231
rect 186 230 187 231
rect 185 230 186 231
rect 184 230 185 231
rect 183 230 184 231
rect 182 230 183 231
rect 181 230 182 231
rect 180 230 181 231
rect 179 230 180 231
rect 178 230 179 231
rect 177 230 178 231
rect 176 230 177 231
rect 175 230 176 231
rect 174 230 175 231
rect 173 230 174 231
rect 172 230 173 231
rect 171 230 172 231
rect 170 230 171 231
rect 169 230 170 231
rect 168 230 169 231
rect 167 230 168 231
rect 166 230 167 231
rect 165 230 166 231
rect 164 230 165 231
rect 163 230 164 231
rect 145 230 146 231
rect 144 230 145 231
rect 143 230 144 231
rect 142 230 143 231
rect 141 230 142 231
rect 140 230 141 231
rect 139 230 140 231
rect 138 230 139 231
rect 137 230 138 231
rect 136 230 137 231
rect 135 230 136 231
rect 134 230 135 231
rect 133 230 134 231
rect 132 230 133 231
rect 131 230 132 231
rect 130 230 131 231
rect 129 230 130 231
rect 128 230 129 231
rect 127 230 128 231
rect 126 230 127 231
rect 125 230 126 231
rect 124 230 125 231
rect 123 230 124 231
rect 122 230 123 231
rect 121 230 122 231
rect 120 230 121 231
rect 119 230 120 231
rect 118 230 119 231
rect 117 230 118 231
rect 116 230 117 231
rect 115 230 116 231
rect 114 230 115 231
rect 85 230 86 231
rect 84 230 85 231
rect 83 230 84 231
rect 82 230 83 231
rect 81 230 82 231
rect 80 230 81 231
rect 79 230 80 231
rect 78 230 79 231
rect 77 230 78 231
rect 76 230 77 231
rect 75 230 76 231
rect 74 230 75 231
rect 73 230 74 231
rect 72 230 73 231
rect 71 230 72 231
rect 70 230 71 231
rect 69 230 70 231
rect 68 230 69 231
rect 67 230 68 231
rect 66 230 67 231
rect 65 230 66 231
rect 64 230 65 231
rect 63 230 64 231
rect 62 230 63 231
rect 61 230 62 231
rect 60 230 61 231
rect 59 230 60 231
rect 58 230 59 231
rect 57 230 58 231
rect 56 230 57 231
rect 55 230 56 231
rect 54 230 55 231
rect 53 230 54 231
rect 52 230 53 231
rect 51 230 52 231
rect 50 230 51 231
rect 49 230 50 231
rect 48 230 49 231
rect 47 230 48 231
rect 46 230 47 231
rect 45 230 46 231
rect 44 230 45 231
rect 43 230 44 231
rect 42 230 43 231
rect 41 230 42 231
rect 40 230 41 231
rect 39 230 40 231
rect 38 230 39 231
rect 37 230 38 231
rect 36 230 37 231
rect 35 230 36 231
rect 34 230 35 231
rect 33 230 34 231
rect 32 230 33 231
rect 31 230 32 231
rect 30 230 31 231
rect 29 230 30 231
rect 28 230 29 231
rect 27 230 28 231
rect 26 230 27 231
rect 25 230 26 231
rect 24 230 25 231
rect 23 230 24 231
rect 22 230 23 231
rect 21 230 22 231
rect 20 230 21 231
rect 19 230 20 231
rect 18 230 19 231
rect 17 230 18 231
rect 16 230 17 231
rect 15 230 16 231
rect 14 230 15 231
rect 13 230 14 231
rect 12 230 13 231
rect 11 230 12 231
rect 10 230 11 231
rect 9 230 10 231
rect 8 230 9 231
rect 7 230 8 231
rect 6 230 7 231
rect 5 230 6 231
rect 480 231 481 232
rect 479 231 480 232
rect 478 231 479 232
rect 477 231 478 232
rect 476 231 477 232
rect 475 231 476 232
rect 474 231 475 232
rect 469 231 470 232
rect 468 231 469 232
rect 467 231 468 232
rect 466 231 467 232
rect 465 231 466 232
rect 464 231 465 232
rect 463 231 464 232
rect 462 231 463 232
rect 461 231 462 232
rect 440 231 441 232
rect 439 231 440 232
rect 438 231 439 232
rect 396 231 397 232
rect 395 231 396 232
rect 394 231 395 232
rect 276 231 277 232
rect 275 231 276 232
rect 274 231 275 232
rect 273 231 274 232
rect 272 231 273 232
rect 271 231 272 232
rect 270 231 271 232
rect 269 231 270 232
rect 268 231 269 232
rect 267 231 268 232
rect 266 231 267 232
rect 265 231 266 232
rect 264 231 265 232
rect 263 231 264 232
rect 262 231 263 232
rect 261 231 262 232
rect 260 231 261 232
rect 259 231 260 232
rect 258 231 259 232
rect 257 231 258 232
rect 256 231 257 232
rect 255 231 256 232
rect 254 231 255 232
rect 253 231 254 232
rect 252 231 253 232
rect 251 231 252 232
rect 250 231 251 232
rect 249 231 250 232
rect 248 231 249 232
rect 247 231 248 232
rect 246 231 247 232
rect 245 231 246 232
rect 244 231 245 232
rect 243 231 244 232
rect 242 231 243 232
rect 241 231 242 232
rect 240 231 241 232
rect 239 231 240 232
rect 238 231 239 232
rect 237 231 238 232
rect 236 231 237 232
rect 235 231 236 232
rect 234 231 235 232
rect 233 231 234 232
rect 232 231 233 232
rect 231 231 232 232
rect 230 231 231 232
rect 229 231 230 232
rect 228 231 229 232
rect 227 231 228 232
rect 226 231 227 232
rect 225 231 226 232
rect 224 231 225 232
rect 223 231 224 232
rect 222 231 223 232
rect 221 231 222 232
rect 220 231 221 232
rect 219 231 220 232
rect 218 231 219 232
rect 217 231 218 232
rect 216 231 217 232
rect 215 231 216 232
rect 214 231 215 232
rect 213 231 214 232
rect 212 231 213 232
rect 211 231 212 232
rect 210 231 211 232
rect 209 231 210 232
rect 208 231 209 232
rect 207 231 208 232
rect 206 231 207 232
rect 205 231 206 232
rect 204 231 205 232
rect 203 231 204 232
rect 202 231 203 232
rect 201 231 202 232
rect 200 231 201 232
rect 199 231 200 232
rect 198 231 199 232
rect 197 231 198 232
rect 196 231 197 232
rect 195 231 196 232
rect 194 231 195 232
rect 193 231 194 232
rect 192 231 193 232
rect 191 231 192 232
rect 190 231 191 232
rect 189 231 190 232
rect 188 231 189 232
rect 187 231 188 232
rect 186 231 187 232
rect 185 231 186 232
rect 184 231 185 232
rect 183 231 184 232
rect 182 231 183 232
rect 181 231 182 232
rect 180 231 181 232
rect 179 231 180 232
rect 178 231 179 232
rect 177 231 178 232
rect 176 231 177 232
rect 175 231 176 232
rect 174 231 175 232
rect 173 231 174 232
rect 172 231 173 232
rect 171 231 172 232
rect 170 231 171 232
rect 169 231 170 232
rect 168 231 169 232
rect 167 231 168 232
rect 166 231 167 232
rect 165 231 166 232
rect 164 231 165 232
rect 145 231 146 232
rect 144 231 145 232
rect 143 231 144 232
rect 142 231 143 232
rect 141 231 142 232
rect 140 231 141 232
rect 139 231 140 232
rect 138 231 139 232
rect 137 231 138 232
rect 136 231 137 232
rect 135 231 136 232
rect 134 231 135 232
rect 133 231 134 232
rect 132 231 133 232
rect 131 231 132 232
rect 130 231 131 232
rect 129 231 130 232
rect 128 231 129 232
rect 127 231 128 232
rect 126 231 127 232
rect 125 231 126 232
rect 124 231 125 232
rect 123 231 124 232
rect 122 231 123 232
rect 121 231 122 232
rect 120 231 121 232
rect 119 231 120 232
rect 118 231 119 232
rect 117 231 118 232
rect 116 231 117 232
rect 115 231 116 232
rect 114 231 115 232
rect 87 231 88 232
rect 86 231 87 232
rect 85 231 86 232
rect 84 231 85 232
rect 83 231 84 232
rect 82 231 83 232
rect 81 231 82 232
rect 80 231 81 232
rect 79 231 80 232
rect 78 231 79 232
rect 77 231 78 232
rect 76 231 77 232
rect 75 231 76 232
rect 74 231 75 232
rect 73 231 74 232
rect 72 231 73 232
rect 71 231 72 232
rect 70 231 71 232
rect 69 231 70 232
rect 68 231 69 232
rect 67 231 68 232
rect 66 231 67 232
rect 65 231 66 232
rect 64 231 65 232
rect 63 231 64 232
rect 62 231 63 232
rect 61 231 62 232
rect 60 231 61 232
rect 59 231 60 232
rect 58 231 59 232
rect 57 231 58 232
rect 56 231 57 232
rect 55 231 56 232
rect 54 231 55 232
rect 53 231 54 232
rect 52 231 53 232
rect 51 231 52 232
rect 50 231 51 232
rect 49 231 50 232
rect 48 231 49 232
rect 47 231 48 232
rect 46 231 47 232
rect 45 231 46 232
rect 44 231 45 232
rect 43 231 44 232
rect 42 231 43 232
rect 41 231 42 232
rect 40 231 41 232
rect 39 231 40 232
rect 38 231 39 232
rect 37 231 38 232
rect 36 231 37 232
rect 35 231 36 232
rect 34 231 35 232
rect 33 231 34 232
rect 32 231 33 232
rect 31 231 32 232
rect 30 231 31 232
rect 29 231 30 232
rect 28 231 29 232
rect 27 231 28 232
rect 26 231 27 232
rect 25 231 26 232
rect 24 231 25 232
rect 23 231 24 232
rect 22 231 23 232
rect 21 231 22 232
rect 20 231 21 232
rect 19 231 20 232
rect 18 231 19 232
rect 17 231 18 232
rect 16 231 17 232
rect 15 231 16 232
rect 14 231 15 232
rect 13 231 14 232
rect 12 231 13 232
rect 11 231 12 232
rect 10 231 11 232
rect 9 231 10 232
rect 8 231 9 232
rect 7 231 8 232
rect 6 231 7 232
rect 5 231 6 232
rect 480 232 481 233
rect 479 232 480 233
rect 478 232 479 233
rect 477 232 478 233
rect 476 232 477 233
rect 468 232 469 233
rect 467 232 468 233
rect 466 232 467 233
rect 465 232 466 233
rect 464 232 465 233
rect 463 232 464 233
rect 462 232 463 233
rect 440 232 441 233
rect 439 232 440 233
rect 438 232 439 233
rect 420 232 421 233
rect 419 232 420 233
rect 418 232 419 233
rect 396 232 397 233
rect 395 232 396 233
rect 394 232 395 233
rect 275 232 276 233
rect 274 232 275 233
rect 273 232 274 233
rect 272 232 273 233
rect 271 232 272 233
rect 270 232 271 233
rect 269 232 270 233
rect 268 232 269 233
rect 267 232 268 233
rect 266 232 267 233
rect 265 232 266 233
rect 264 232 265 233
rect 263 232 264 233
rect 262 232 263 233
rect 261 232 262 233
rect 260 232 261 233
rect 259 232 260 233
rect 258 232 259 233
rect 257 232 258 233
rect 256 232 257 233
rect 255 232 256 233
rect 254 232 255 233
rect 253 232 254 233
rect 252 232 253 233
rect 251 232 252 233
rect 250 232 251 233
rect 249 232 250 233
rect 248 232 249 233
rect 247 232 248 233
rect 246 232 247 233
rect 245 232 246 233
rect 244 232 245 233
rect 243 232 244 233
rect 242 232 243 233
rect 241 232 242 233
rect 240 232 241 233
rect 239 232 240 233
rect 238 232 239 233
rect 237 232 238 233
rect 236 232 237 233
rect 235 232 236 233
rect 234 232 235 233
rect 233 232 234 233
rect 232 232 233 233
rect 231 232 232 233
rect 230 232 231 233
rect 229 232 230 233
rect 228 232 229 233
rect 227 232 228 233
rect 226 232 227 233
rect 225 232 226 233
rect 224 232 225 233
rect 223 232 224 233
rect 222 232 223 233
rect 221 232 222 233
rect 220 232 221 233
rect 219 232 220 233
rect 218 232 219 233
rect 217 232 218 233
rect 216 232 217 233
rect 215 232 216 233
rect 214 232 215 233
rect 213 232 214 233
rect 212 232 213 233
rect 211 232 212 233
rect 210 232 211 233
rect 209 232 210 233
rect 208 232 209 233
rect 207 232 208 233
rect 206 232 207 233
rect 205 232 206 233
rect 204 232 205 233
rect 203 232 204 233
rect 202 232 203 233
rect 201 232 202 233
rect 200 232 201 233
rect 199 232 200 233
rect 198 232 199 233
rect 197 232 198 233
rect 196 232 197 233
rect 195 232 196 233
rect 194 232 195 233
rect 193 232 194 233
rect 192 232 193 233
rect 191 232 192 233
rect 190 232 191 233
rect 189 232 190 233
rect 188 232 189 233
rect 187 232 188 233
rect 186 232 187 233
rect 185 232 186 233
rect 184 232 185 233
rect 183 232 184 233
rect 182 232 183 233
rect 181 232 182 233
rect 180 232 181 233
rect 179 232 180 233
rect 178 232 179 233
rect 177 232 178 233
rect 176 232 177 233
rect 175 232 176 233
rect 174 232 175 233
rect 173 232 174 233
rect 172 232 173 233
rect 171 232 172 233
rect 170 232 171 233
rect 169 232 170 233
rect 168 232 169 233
rect 167 232 168 233
rect 166 232 167 233
rect 165 232 166 233
rect 145 232 146 233
rect 144 232 145 233
rect 143 232 144 233
rect 142 232 143 233
rect 141 232 142 233
rect 140 232 141 233
rect 139 232 140 233
rect 138 232 139 233
rect 137 232 138 233
rect 136 232 137 233
rect 135 232 136 233
rect 134 232 135 233
rect 133 232 134 233
rect 132 232 133 233
rect 131 232 132 233
rect 130 232 131 233
rect 129 232 130 233
rect 128 232 129 233
rect 127 232 128 233
rect 126 232 127 233
rect 125 232 126 233
rect 124 232 125 233
rect 123 232 124 233
rect 122 232 123 233
rect 121 232 122 233
rect 120 232 121 233
rect 119 232 120 233
rect 118 232 119 233
rect 117 232 118 233
rect 116 232 117 233
rect 115 232 116 233
rect 89 232 90 233
rect 88 232 89 233
rect 87 232 88 233
rect 86 232 87 233
rect 85 232 86 233
rect 84 232 85 233
rect 83 232 84 233
rect 82 232 83 233
rect 81 232 82 233
rect 80 232 81 233
rect 79 232 80 233
rect 78 232 79 233
rect 77 232 78 233
rect 76 232 77 233
rect 75 232 76 233
rect 74 232 75 233
rect 73 232 74 233
rect 72 232 73 233
rect 71 232 72 233
rect 70 232 71 233
rect 69 232 70 233
rect 68 232 69 233
rect 67 232 68 233
rect 66 232 67 233
rect 65 232 66 233
rect 64 232 65 233
rect 63 232 64 233
rect 62 232 63 233
rect 61 232 62 233
rect 60 232 61 233
rect 59 232 60 233
rect 58 232 59 233
rect 57 232 58 233
rect 56 232 57 233
rect 55 232 56 233
rect 54 232 55 233
rect 53 232 54 233
rect 52 232 53 233
rect 51 232 52 233
rect 50 232 51 233
rect 49 232 50 233
rect 48 232 49 233
rect 47 232 48 233
rect 46 232 47 233
rect 45 232 46 233
rect 44 232 45 233
rect 43 232 44 233
rect 42 232 43 233
rect 41 232 42 233
rect 40 232 41 233
rect 39 232 40 233
rect 38 232 39 233
rect 37 232 38 233
rect 36 232 37 233
rect 35 232 36 233
rect 34 232 35 233
rect 33 232 34 233
rect 32 232 33 233
rect 31 232 32 233
rect 30 232 31 233
rect 29 232 30 233
rect 28 232 29 233
rect 27 232 28 233
rect 26 232 27 233
rect 23 232 24 233
rect 22 232 23 233
rect 21 232 22 233
rect 20 232 21 233
rect 19 232 20 233
rect 18 232 19 233
rect 17 232 18 233
rect 16 232 17 233
rect 15 232 16 233
rect 14 232 15 233
rect 13 232 14 233
rect 12 232 13 233
rect 11 232 12 233
rect 10 232 11 233
rect 9 232 10 233
rect 8 232 9 233
rect 7 232 8 233
rect 6 232 7 233
rect 5 232 6 233
rect 4 232 5 233
rect 481 233 482 234
rect 480 233 481 234
rect 479 233 480 234
rect 478 233 479 234
rect 440 233 441 234
rect 439 233 440 234
rect 438 233 439 234
rect 420 233 421 234
rect 419 233 420 234
rect 418 233 419 234
rect 396 233 397 234
rect 395 233 396 234
rect 394 233 395 234
rect 274 233 275 234
rect 273 233 274 234
rect 272 233 273 234
rect 271 233 272 234
rect 270 233 271 234
rect 269 233 270 234
rect 268 233 269 234
rect 267 233 268 234
rect 266 233 267 234
rect 265 233 266 234
rect 264 233 265 234
rect 263 233 264 234
rect 262 233 263 234
rect 261 233 262 234
rect 260 233 261 234
rect 259 233 260 234
rect 258 233 259 234
rect 257 233 258 234
rect 256 233 257 234
rect 255 233 256 234
rect 254 233 255 234
rect 253 233 254 234
rect 252 233 253 234
rect 251 233 252 234
rect 250 233 251 234
rect 249 233 250 234
rect 248 233 249 234
rect 247 233 248 234
rect 246 233 247 234
rect 245 233 246 234
rect 244 233 245 234
rect 243 233 244 234
rect 242 233 243 234
rect 241 233 242 234
rect 240 233 241 234
rect 239 233 240 234
rect 238 233 239 234
rect 237 233 238 234
rect 236 233 237 234
rect 235 233 236 234
rect 234 233 235 234
rect 233 233 234 234
rect 232 233 233 234
rect 231 233 232 234
rect 230 233 231 234
rect 229 233 230 234
rect 228 233 229 234
rect 227 233 228 234
rect 226 233 227 234
rect 225 233 226 234
rect 224 233 225 234
rect 223 233 224 234
rect 222 233 223 234
rect 221 233 222 234
rect 220 233 221 234
rect 219 233 220 234
rect 218 233 219 234
rect 217 233 218 234
rect 216 233 217 234
rect 215 233 216 234
rect 214 233 215 234
rect 213 233 214 234
rect 212 233 213 234
rect 211 233 212 234
rect 210 233 211 234
rect 209 233 210 234
rect 208 233 209 234
rect 207 233 208 234
rect 206 233 207 234
rect 205 233 206 234
rect 204 233 205 234
rect 203 233 204 234
rect 202 233 203 234
rect 201 233 202 234
rect 200 233 201 234
rect 199 233 200 234
rect 198 233 199 234
rect 197 233 198 234
rect 196 233 197 234
rect 195 233 196 234
rect 194 233 195 234
rect 193 233 194 234
rect 192 233 193 234
rect 191 233 192 234
rect 190 233 191 234
rect 189 233 190 234
rect 188 233 189 234
rect 187 233 188 234
rect 186 233 187 234
rect 185 233 186 234
rect 184 233 185 234
rect 183 233 184 234
rect 182 233 183 234
rect 181 233 182 234
rect 180 233 181 234
rect 179 233 180 234
rect 178 233 179 234
rect 177 233 178 234
rect 176 233 177 234
rect 175 233 176 234
rect 174 233 175 234
rect 173 233 174 234
rect 172 233 173 234
rect 171 233 172 234
rect 170 233 171 234
rect 169 233 170 234
rect 168 233 169 234
rect 167 233 168 234
rect 145 233 146 234
rect 144 233 145 234
rect 143 233 144 234
rect 142 233 143 234
rect 141 233 142 234
rect 140 233 141 234
rect 139 233 140 234
rect 138 233 139 234
rect 137 233 138 234
rect 136 233 137 234
rect 135 233 136 234
rect 134 233 135 234
rect 133 233 134 234
rect 132 233 133 234
rect 131 233 132 234
rect 130 233 131 234
rect 129 233 130 234
rect 128 233 129 234
rect 127 233 128 234
rect 126 233 127 234
rect 125 233 126 234
rect 124 233 125 234
rect 123 233 124 234
rect 122 233 123 234
rect 121 233 122 234
rect 120 233 121 234
rect 119 233 120 234
rect 118 233 119 234
rect 117 233 118 234
rect 116 233 117 234
rect 92 233 93 234
rect 91 233 92 234
rect 90 233 91 234
rect 89 233 90 234
rect 88 233 89 234
rect 87 233 88 234
rect 86 233 87 234
rect 85 233 86 234
rect 84 233 85 234
rect 83 233 84 234
rect 82 233 83 234
rect 81 233 82 234
rect 80 233 81 234
rect 79 233 80 234
rect 78 233 79 234
rect 77 233 78 234
rect 76 233 77 234
rect 75 233 76 234
rect 74 233 75 234
rect 73 233 74 234
rect 72 233 73 234
rect 71 233 72 234
rect 70 233 71 234
rect 69 233 70 234
rect 68 233 69 234
rect 67 233 68 234
rect 66 233 67 234
rect 65 233 66 234
rect 64 233 65 234
rect 63 233 64 234
rect 62 233 63 234
rect 61 233 62 234
rect 60 233 61 234
rect 59 233 60 234
rect 58 233 59 234
rect 57 233 58 234
rect 56 233 57 234
rect 55 233 56 234
rect 54 233 55 234
rect 53 233 54 234
rect 52 233 53 234
rect 51 233 52 234
rect 50 233 51 234
rect 49 233 50 234
rect 48 233 49 234
rect 47 233 48 234
rect 46 233 47 234
rect 45 233 46 234
rect 44 233 45 234
rect 43 233 44 234
rect 42 233 43 234
rect 41 233 42 234
rect 40 233 41 234
rect 39 233 40 234
rect 38 233 39 234
rect 37 233 38 234
rect 36 233 37 234
rect 35 233 36 234
rect 34 233 35 234
rect 33 233 34 234
rect 32 233 33 234
rect 31 233 32 234
rect 30 233 31 234
rect 29 233 30 234
rect 28 233 29 234
rect 27 233 28 234
rect 26 233 27 234
rect 22 233 23 234
rect 21 233 22 234
rect 20 233 21 234
rect 19 233 20 234
rect 18 233 19 234
rect 17 233 18 234
rect 16 233 17 234
rect 15 233 16 234
rect 14 233 15 234
rect 13 233 14 234
rect 12 233 13 234
rect 11 233 12 234
rect 10 233 11 234
rect 9 233 10 234
rect 8 233 9 234
rect 7 233 8 234
rect 6 233 7 234
rect 5 233 6 234
rect 4 233 5 234
rect 481 234 482 235
rect 480 234 481 235
rect 479 234 480 235
rect 440 234 441 235
rect 439 234 440 235
rect 438 234 439 235
rect 420 234 421 235
rect 419 234 420 235
rect 418 234 419 235
rect 396 234 397 235
rect 395 234 396 235
rect 394 234 395 235
rect 273 234 274 235
rect 272 234 273 235
rect 271 234 272 235
rect 270 234 271 235
rect 269 234 270 235
rect 268 234 269 235
rect 267 234 268 235
rect 266 234 267 235
rect 265 234 266 235
rect 264 234 265 235
rect 263 234 264 235
rect 262 234 263 235
rect 261 234 262 235
rect 260 234 261 235
rect 259 234 260 235
rect 258 234 259 235
rect 257 234 258 235
rect 256 234 257 235
rect 255 234 256 235
rect 254 234 255 235
rect 253 234 254 235
rect 252 234 253 235
rect 251 234 252 235
rect 250 234 251 235
rect 249 234 250 235
rect 248 234 249 235
rect 247 234 248 235
rect 246 234 247 235
rect 245 234 246 235
rect 244 234 245 235
rect 243 234 244 235
rect 242 234 243 235
rect 241 234 242 235
rect 240 234 241 235
rect 239 234 240 235
rect 238 234 239 235
rect 237 234 238 235
rect 236 234 237 235
rect 235 234 236 235
rect 234 234 235 235
rect 233 234 234 235
rect 232 234 233 235
rect 231 234 232 235
rect 230 234 231 235
rect 229 234 230 235
rect 228 234 229 235
rect 227 234 228 235
rect 226 234 227 235
rect 225 234 226 235
rect 224 234 225 235
rect 223 234 224 235
rect 222 234 223 235
rect 221 234 222 235
rect 220 234 221 235
rect 219 234 220 235
rect 218 234 219 235
rect 217 234 218 235
rect 216 234 217 235
rect 215 234 216 235
rect 214 234 215 235
rect 213 234 214 235
rect 212 234 213 235
rect 211 234 212 235
rect 210 234 211 235
rect 209 234 210 235
rect 208 234 209 235
rect 207 234 208 235
rect 206 234 207 235
rect 205 234 206 235
rect 204 234 205 235
rect 203 234 204 235
rect 202 234 203 235
rect 201 234 202 235
rect 200 234 201 235
rect 199 234 200 235
rect 198 234 199 235
rect 197 234 198 235
rect 196 234 197 235
rect 195 234 196 235
rect 194 234 195 235
rect 193 234 194 235
rect 192 234 193 235
rect 191 234 192 235
rect 190 234 191 235
rect 189 234 190 235
rect 188 234 189 235
rect 187 234 188 235
rect 186 234 187 235
rect 185 234 186 235
rect 184 234 185 235
rect 183 234 184 235
rect 182 234 183 235
rect 181 234 182 235
rect 180 234 181 235
rect 179 234 180 235
rect 178 234 179 235
rect 177 234 178 235
rect 176 234 177 235
rect 175 234 176 235
rect 174 234 175 235
rect 173 234 174 235
rect 172 234 173 235
rect 171 234 172 235
rect 170 234 171 235
rect 169 234 170 235
rect 168 234 169 235
rect 146 234 147 235
rect 145 234 146 235
rect 144 234 145 235
rect 143 234 144 235
rect 142 234 143 235
rect 141 234 142 235
rect 140 234 141 235
rect 139 234 140 235
rect 138 234 139 235
rect 137 234 138 235
rect 136 234 137 235
rect 135 234 136 235
rect 134 234 135 235
rect 133 234 134 235
rect 132 234 133 235
rect 131 234 132 235
rect 130 234 131 235
rect 129 234 130 235
rect 128 234 129 235
rect 127 234 128 235
rect 126 234 127 235
rect 125 234 126 235
rect 124 234 125 235
rect 123 234 124 235
rect 122 234 123 235
rect 121 234 122 235
rect 120 234 121 235
rect 119 234 120 235
rect 118 234 119 235
rect 117 234 118 235
rect 116 234 117 235
rect 94 234 95 235
rect 93 234 94 235
rect 92 234 93 235
rect 91 234 92 235
rect 90 234 91 235
rect 89 234 90 235
rect 88 234 89 235
rect 87 234 88 235
rect 86 234 87 235
rect 85 234 86 235
rect 84 234 85 235
rect 83 234 84 235
rect 82 234 83 235
rect 81 234 82 235
rect 80 234 81 235
rect 79 234 80 235
rect 78 234 79 235
rect 77 234 78 235
rect 76 234 77 235
rect 75 234 76 235
rect 74 234 75 235
rect 73 234 74 235
rect 72 234 73 235
rect 71 234 72 235
rect 70 234 71 235
rect 69 234 70 235
rect 68 234 69 235
rect 67 234 68 235
rect 66 234 67 235
rect 65 234 66 235
rect 64 234 65 235
rect 63 234 64 235
rect 62 234 63 235
rect 61 234 62 235
rect 60 234 61 235
rect 59 234 60 235
rect 58 234 59 235
rect 57 234 58 235
rect 56 234 57 235
rect 55 234 56 235
rect 54 234 55 235
rect 53 234 54 235
rect 52 234 53 235
rect 51 234 52 235
rect 50 234 51 235
rect 49 234 50 235
rect 48 234 49 235
rect 47 234 48 235
rect 46 234 47 235
rect 45 234 46 235
rect 44 234 45 235
rect 43 234 44 235
rect 42 234 43 235
rect 41 234 42 235
rect 40 234 41 235
rect 39 234 40 235
rect 38 234 39 235
rect 37 234 38 235
rect 36 234 37 235
rect 35 234 36 235
rect 34 234 35 235
rect 33 234 34 235
rect 32 234 33 235
rect 31 234 32 235
rect 30 234 31 235
rect 29 234 30 235
rect 28 234 29 235
rect 27 234 28 235
rect 22 234 23 235
rect 21 234 22 235
rect 20 234 21 235
rect 19 234 20 235
rect 18 234 19 235
rect 17 234 18 235
rect 16 234 17 235
rect 15 234 16 235
rect 14 234 15 235
rect 13 234 14 235
rect 12 234 13 235
rect 11 234 12 235
rect 10 234 11 235
rect 9 234 10 235
rect 8 234 9 235
rect 7 234 8 235
rect 6 234 7 235
rect 5 234 6 235
rect 4 234 5 235
rect 481 235 482 236
rect 480 235 481 236
rect 440 235 441 236
rect 439 235 440 236
rect 438 235 439 236
rect 421 235 422 236
rect 420 235 421 236
rect 419 235 420 236
rect 418 235 419 236
rect 396 235 397 236
rect 395 235 396 236
rect 394 235 395 236
rect 272 235 273 236
rect 271 235 272 236
rect 270 235 271 236
rect 269 235 270 236
rect 268 235 269 236
rect 267 235 268 236
rect 266 235 267 236
rect 265 235 266 236
rect 264 235 265 236
rect 263 235 264 236
rect 262 235 263 236
rect 261 235 262 236
rect 260 235 261 236
rect 259 235 260 236
rect 258 235 259 236
rect 257 235 258 236
rect 256 235 257 236
rect 255 235 256 236
rect 254 235 255 236
rect 253 235 254 236
rect 252 235 253 236
rect 251 235 252 236
rect 250 235 251 236
rect 249 235 250 236
rect 248 235 249 236
rect 247 235 248 236
rect 246 235 247 236
rect 245 235 246 236
rect 244 235 245 236
rect 243 235 244 236
rect 242 235 243 236
rect 241 235 242 236
rect 240 235 241 236
rect 239 235 240 236
rect 238 235 239 236
rect 237 235 238 236
rect 236 235 237 236
rect 235 235 236 236
rect 234 235 235 236
rect 233 235 234 236
rect 232 235 233 236
rect 231 235 232 236
rect 230 235 231 236
rect 229 235 230 236
rect 228 235 229 236
rect 227 235 228 236
rect 226 235 227 236
rect 225 235 226 236
rect 224 235 225 236
rect 223 235 224 236
rect 222 235 223 236
rect 221 235 222 236
rect 220 235 221 236
rect 219 235 220 236
rect 218 235 219 236
rect 217 235 218 236
rect 216 235 217 236
rect 215 235 216 236
rect 214 235 215 236
rect 213 235 214 236
rect 212 235 213 236
rect 211 235 212 236
rect 210 235 211 236
rect 209 235 210 236
rect 208 235 209 236
rect 207 235 208 236
rect 206 235 207 236
rect 205 235 206 236
rect 204 235 205 236
rect 203 235 204 236
rect 202 235 203 236
rect 201 235 202 236
rect 200 235 201 236
rect 199 235 200 236
rect 198 235 199 236
rect 197 235 198 236
rect 196 235 197 236
rect 195 235 196 236
rect 194 235 195 236
rect 193 235 194 236
rect 192 235 193 236
rect 191 235 192 236
rect 190 235 191 236
rect 189 235 190 236
rect 188 235 189 236
rect 187 235 188 236
rect 186 235 187 236
rect 185 235 186 236
rect 184 235 185 236
rect 183 235 184 236
rect 182 235 183 236
rect 181 235 182 236
rect 180 235 181 236
rect 179 235 180 236
rect 178 235 179 236
rect 177 235 178 236
rect 176 235 177 236
rect 175 235 176 236
rect 174 235 175 236
rect 173 235 174 236
rect 172 235 173 236
rect 171 235 172 236
rect 170 235 171 236
rect 146 235 147 236
rect 145 235 146 236
rect 144 235 145 236
rect 143 235 144 236
rect 142 235 143 236
rect 141 235 142 236
rect 140 235 141 236
rect 139 235 140 236
rect 138 235 139 236
rect 137 235 138 236
rect 136 235 137 236
rect 135 235 136 236
rect 134 235 135 236
rect 133 235 134 236
rect 132 235 133 236
rect 131 235 132 236
rect 130 235 131 236
rect 129 235 130 236
rect 128 235 129 236
rect 127 235 128 236
rect 126 235 127 236
rect 125 235 126 236
rect 124 235 125 236
rect 123 235 124 236
rect 122 235 123 236
rect 121 235 122 236
rect 120 235 121 236
rect 119 235 120 236
rect 118 235 119 236
rect 117 235 118 236
rect 96 235 97 236
rect 95 235 96 236
rect 94 235 95 236
rect 93 235 94 236
rect 92 235 93 236
rect 91 235 92 236
rect 90 235 91 236
rect 89 235 90 236
rect 88 235 89 236
rect 87 235 88 236
rect 86 235 87 236
rect 85 235 86 236
rect 84 235 85 236
rect 83 235 84 236
rect 82 235 83 236
rect 81 235 82 236
rect 80 235 81 236
rect 79 235 80 236
rect 78 235 79 236
rect 77 235 78 236
rect 76 235 77 236
rect 75 235 76 236
rect 74 235 75 236
rect 73 235 74 236
rect 72 235 73 236
rect 71 235 72 236
rect 70 235 71 236
rect 69 235 70 236
rect 68 235 69 236
rect 67 235 68 236
rect 66 235 67 236
rect 65 235 66 236
rect 64 235 65 236
rect 63 235 64 236
rect 62 235 63 236
rect 61 235 62 236
rect 60 235 61 236
rect 59 235 60 236
rect 58 235 59 236
rect 57 235 58 236
rect 56 235 57 236
rect 55 235 56 236
rect 54 235 55 236
rect 53 235 54 236
rect 52 235 53 236
rect 51 235 52 236
rect 50 235 51 236
rect 49 235 50 236
rect 48 235 49 236
rect 47 235 48 236
rect 46 235 47 236
rect 45 235 46 236
rect 44 235 45 236
rect 43 235 44 236
rect 42 235 43 236
rect 41 235 42 236
rect 40 235 41 236
rect 39 235 40 236
rect 38 235 39 236
rect 37 235 38 236
rect 36 235 37 236
rect 35 235 36 236
rect 34 235 35 236
rect 33 235 34 236
rect 32 235 33 236
rect 31 235 32 236
rect 30 235 31 236
rect 29 235 30 236
rect 28 235 29 236
rect 27 235 28 236
rect 22 235 23 236
rect 21 235 22 236
rect 20 235 21 236
rect 19 235 20 236
rect 18 235 19 236
rect 17 235 18 236
rect 16 235 17 236
rect 15 235 16 236
rect 14 235 15 236
rect 13 235 14 236
rect 12 235 13 236
rect 11 235 12 236
rect 10 235 11 236
rect 9 235 10 236
rect 8 235 9 236
rect 7 235 8 236
rect 6 235 7 236
rect 5 235 6 236
rect 4 235 5 236
rect 440 236 441 237
rect 439 236 440 237
rect 438 236 439 237
rect 421 236 422 237
rect 420 236 421 237
rect 419 236 420 237
rect 418 236 419 237
rect 396 236 397 237
rect 395 236 396 237
rect 394 236 395 237
rect 271 236 272 237
rect 270 236 271 237
rect 269 236 270 237
rect 268 236 269 237
rect 267 236 268 237
rect 266 236 267 237
rect 265 236 266 237
rect 264 236 265 237
rect 263 236 264 237
rect 262 236 263 237
rect 261 236 262 237
rect 260 236 261 237
rect 259 236 260 237
rect 258 236 259 237
rect 257 236 258 237
rect 256 236 257 237
rect 255 236 256 237
rect 254 236 255 237
rect 253 236 254 237
rect 252 236 253 237
rect 251 236 252 237
rect 250 236 251 237
rect 249 236 250 237
rect 248 236 249 237
rect 247 236 248 237
rect 246 236 247 237
rect 245 236 246 237
rect 244 236 245 237
rect 243 236 244 237
rect 242 236 243 237
rect 241 236 242 237
rect 240 236 241 237
rect 239 236 240 237
rect 238 236 239 237
rect 237 236 238 237
rect 236 236 237 237
rect 235 236 236 237
rect 234 236 235 237
rect 233 236 234 237
rect 232 236 233 237
rect 231 236 232 237
rect 230 236 231 237
rect 229 236 230 237
rect 228 236 229 237
rect 227 236 228 237
rect 226 236 227 237
rect 225 236 226 237
rect 224 236 225 237
rect 223 236 224 237
rect 222 236 223 237
rect 221 236 222 237
rect 220 236 221 237
rect 219 236 220 237
rect 218 236 219 237
rect 217 236 218 237
rect 216 236 217 237
rect 215 236 216 237
rect 214 236 215 237
rect 213 236 214 237
rect 212 236 213 237
rect 211 236 212 237
rect 210 236 211 237
rect 209 236 210 237
rect 208 236 209 237
rect 207 236 208 237
rect 206 236 207 237
rect 205 236 206 237
rect 204 236 205 237
rect 203 236 204 237
rect 202 236 203 237
rect 201 236 202 237
rect 200 236 201 237
rect 199 236 200 237
rect 198 236 199 237
rect 197 236 198 237
rect 196 236 197 237
rect 195 236 196 237
rect 194 236 195 237
rect 193 236 194 237
rect 192 236 193 237
rect 191 236 192 237
rect 190 236 191 237
rect 189 236 190 237
rect 188 236 189 237
rect 187 236 188 237
rect 186 236 187 237
rect 185 236 186 237
rect 184 236 185 237
rect 183 236 184 237
rect 182 236 183 237
rect 181 236 182 237
rect 180 236 181 237
rect 179 236 180 237
rect 178 236 179 237
rect 177 236 178 237
rect 176 236 177 237
rect 175 236 176 237
rect 174 236 175 237
rect 173 236 174 237
rect 172 236 173 237
rect 171 236 172 237
rect 147 236 148 237
rect 146 236 147 237
rect 145 236 146 237
rect 144 236 145 237
rect 143 236 144 237
rect 142 236 143 237
rect 141 236 142 237
rect 140 236 141 237
rect 139 236 140 237
rect 138 236 139 237
rect 137 236 138 237
rect 136 236 137 237
rect 135 236 136 237
rect 134 236 135 237
rect 133 236 134 237
rect 132 236 133 237
rect 131 236 132 237
rect 130 236 131 237
rect 129 236 130 237
rect 128 236 129 237
rect 127 236 128 237
rect 126 236 127 237
rect 125 236 126 237
rect 124 236 125 237
rect 123 236 124 237
rect 122 236 123 237
rect 121 236 122 237
rect 120 236 121 237
rect 119 236 120 237
rect 118 236 119 237
rect 117 236 118 237
rect 97 236 98 237
rect 96 236 97 237
rect 95 236 96 237
rect 94 236 95 237
rect 93 236 94 237
rect 92 236 93 237
rect 91 236 92 237
rect 90 236 91 237
rect 89 236 90 237
rect 88 236 89 237
rect 87 236 88 237
rect 86 236 87 237
rect 85 236 86 237
rect 84 236 85 237
rect 83 236 84 237
rect 82 236 83 237
rect 81 236 82 237
rect 80 236 81 237
rect 79 236 80 237
rect 78 236 79 237
rect 77 236 78 237
rect 76 236 77 237
rect 75 236 76 237
rect 74 236 75 237
rect 73 236 74 237
rect 72 236 73 237
rect 71 236 72 237
rect 70 236 71 237
rect 69 236 70 237
rect 68 236 69 237
rect 67 236 68 237
rect 66 236 67 237
rect 65 236 66 237
rect 64 236 65 237
rect 63 236 64 237
rect 62 236 63 237
rect 61 236 62 237
rect 60 236 61 237
rect 59 236 60 237
rect 58 236 59 237
rect 57 236 58 237
rect 56 236 57 237
rect 55 236 56 237
rect 54 236 55 237
rect 53 236 54 237
rect 52 236 53 237
rect 51 236 52 237
rect 50 236 51 237
rect 49 236 50 237
rect 48 236 49 237
rect 47 236 48 237
rect 46 236 47 237
rect 45 236 46 237
rect 44 236 45 237
rect 43 236 44 237
rect 42 236 43 237
rect 41 236 42 237
rect 40 236 41 237
rect 39 236 40 237
rect 38 236 39 237
rect 37 236 38 237
rect 36 236 37 237
rect 35 236 36 237
rect 34 236 35 237
rect 33 236 34 237
rect 32 236 33 237
rect 31 236 32 237
rect 30 236 31 237
rect 29 236 30 237
rect 28 236 29 237
rect 27 236 28 237
rect 21 236 22 237
rect 20 236 21 237
rect 19 236 20 237
rect 18 236 19 237
rect 17 236 18 237
rect 16 236 17 237
rect 15 236 16 237
rect 14 236 15 237
rect 13 236 14 237
rect 12 236 13 237
rect 11 236 12 237
rect 10 236 11 237
rect 9 236 10 237
rect 8 236 9 237
rect 7 236 8 237
rect 6 236 7 237
rect 5 236 6 237
rect 4 236 5 237
rect 440 237 441 238
rect 439 237 440 238
rect 438 237 439 238
rect 421 237 422 238
rect 420 237 421 238
rect 419 237 420 238
rect 418 237 419 238
rect 397 237 398 238
rect 396 237 397 238
rect 395 237 396 238
rect 394 237 395 238
rect 271 237 272 238
rect 270 237 271 238
rect 269 237 270 238
rect 268 237 269 238
rect 267 237 268 238
rect 266 237 267 238
rect 265 237 266 238
rect 264 237 265 238
rect 263 237 264 238
rect 262 237 263 238
rect 261 237 262 238
rect 260 237 261 238
rect 259 237 260 238
rect 258 237 259 238
rect 257 237 258 238
rect 256 237 257 238
rect 255 237 256 238
rect 254 237 255 238
rect 253 237 254 238
rect 252 237 253 238
rect 251 237 252 238
rect 250 237 251 238
rect 249 237 250 238
rect 248 237 249 238
rect 247 237 248 238
rect 246 237 247 238
rect 245 237 246 238
rect 244 237 245 238
rect 243 237 244 238
rect 242 237 243 238
rect 241 237 242 238
rect 240 237 241 238
rect 239 237 240 238
rect 238 237 239 238
rect 237 237 238 238
rect 236 237 237 238
rect 235 237 236 238
rect 234 237 235 238
rect 233 237 234 238
rect 232 237 233 238
rect 231 237 232 238
rect 230 237 231 238
rect 229 237 230 238
rect 228 237 229 238
rect 227 237 228 238
rect 226 237 227 238
rect 225 237 226 238
rect 224 237 225 238
rect 223 237 224 238
rect 222 237 223 238
rect 221 237 222 238
rect 220 237 221 238
rect 219 237 220 238
rect 218 237 219 238
rect 217 237 218 238
rect 216 237 217 238
rect 215 237 216 238
rect 214 237 215 238
rect 213 237 214 238
rect 212 237 213 238
rect 211 237 212 238
rect 210 237 211 238
rect 209 237 210 238
rect 208 237 209 238
rect 207 237 208 238
rect 206 237 207 238
rect 205 237 206 238
rect 204 237 205 238
rect 203 237 204 238
rect 202 237 203 238
rect 201 237 202 238
rect 200 237 201 238
rect 199 237 200 238
rect 198 237 199 238
rect 197 237 198 238
rect 196 237 197 238
rect 195 237 196 238
rect 194 237 195 238
rect 193 237 194 238
rect 192 237 193 238
rect 191 237 192 238
rect 190 237 191 238
rect 189 237 190 238
rect 188 237 189 238
rect 187 237 188 238
rect 186 237 187 238
rect 185 237 186 238
rect 184 237 185 238
rect 183 237 184 238
rect 182 237 183 238
rect 181 237 182 238
rect 180 237 181 238
rect 179 237 180 238
rect 178 237 179 238
rect 177 237 178 238
rect 176 237 177 238
rect 175 237 176 238
rect 174 237 175 238
rect 173 237 174 238
rect 147 237 148 238
rect 146 237 147 238
rect 145 237 146 238
rect 144 237 145 238
rect 143 237 144 238
rect 142 237 143 238
rect 141 237 142 238
rect 140 237 141 238
rect 139 237 140 238
rect 138 237 139 238
rect 137 237 138 238
rect 136 237 137 238
rect 135 237 136 238
rect 134 237 135 238
rect 133 237 134 238
rect 132 237 133 238
rect 131 237 132 238
rect 130 237 131 238
rect 129 237 130 238
rect 128 237 129 238
rect 127 237 128 238
rect 126 237 127 238
rect 125 237 126 238
rect 124 237 125 238
rect 123 237 124 238
rect 122 237 123 238
rect 121 237 122 238
rect 120 237 121 238
rect 119 237 120 238
rect 118 237 119 238
rect 117 237 118 238
rect 99 237 100 238
rect 98 237 99 238
rect 97 237 98 238
rect 96 237 97 238
rect 95 237 96 238
rect 94 237 95 238
rect 93 237 94 238
rect 92 237 93 238
rect 91 237 92 238
rect 90 237 91 238
rect 89 237 90 238
rect 88 237 89 238
rect 87 237 88 238
rect 86 237 87 238
rect 85 237 86 238
rect 84 237 85 238
rect 83 237 84 238
rect 82 237 83 238
rect 81 237 82 238
rect 80 237 81 238
rect 79 237 80 238
rect 78 237 79 238
rect 77 237 78 238
rect 76 237 77 238
rect 75 237 76 238
rect 74 237 75 238
rect 73 237 74 238
rect 72 237 73 238
rect 71 237 72 238
rect 70 237 71 238
rect 69 237 70 238
rect 68 237 69 238
rect 67 237 68 238
rect 66 237 67 238
rect 65 237 66 238
rect 64 237 65 238
rect 63 237 64 238
rect 62 237 63 238
rect 61 237 62 238
rect 60 237 61 238
rect 59 237 60 238
rect 58 237 59 238
rect 57 237 58 238
rect 56 237 57 238
rect 55 237 56 238
rect 54 237 55 238
rect 53 237 54 238
rect 52 237 53 238
rect 51 237 52 238
rect 50 237 51 238
rect 49 237 50 238
rect 48 237 49 238
rect 47 237 48 238
rect 46 237 47 238
rect 45 237 46 238
rect 44 237 45 238
rect 43 237 44 238
rect 42 237 43 238
rect 41 237 42 238
rect 40 237 41 238
rect 39 237 40 238
rect 38 237 39 238
rect 37 237 38 238
rect 36 237 37 238
rect 35 237 36 238
rect 34 237 35 238
rect 33 237 34 238
rect 32 237 33 238
rect 31 237 32 238
rect 30 237 31 238
rect 29 237 30 238
rect 28 237 29 238
rect 27 237 28 238
rect 21 237 22 238
rect 20 237 21 238
rect 19 237 20 238
rect 18 237 19 238
rect 17 237 18 238
rect 16 237 17 238
rect 15 237 16 238
rect 14 237 15 238
rect 13 237 14 238
rect 12 237 13 238
rect 11 237 12 238
rect 10 237 11 238
rect 9 237 10 238
rect 8 237 9 238
rect 7 237 8 238
rect 6 237 7 238
rect 5 237 6 238
rect 4 237 5 238
rect 440 238 441 239
rect 439 238 440 239
rect 438 238 439 239
rect 437 238 438 239
rect 422 238 423 239
rect 421 238 422 239
rect 420 238 421 239
rect 419 238 420 239
rect 418 238 419 239
rect 397 238 398 239
rect 396 238 397 239
rect 395 238 396 239
rect 394 238 395 239
rect 270 238 271 239
rect 269 238 270 239
rect 268 238 269 239
rect 267 238 268 239
rect 266 238 267 239
rect 265 238 266 239
rect 264 238 265 239
rect 263 238 264 239
rect 262 238 263 239
rect 261 238 262 239
rect 260 238 261 239
rect 259 238 260 239
rect 258 238 259 239
rect 257 238 258 239
rect 256 238 257 239
rect 255 238 256 239
rect 254 238 255 239
rect 253 238 254 239
rect 252 238 253 239
rect 251 238 252 239
rect 250 238 251 239
rect 249 238 250 239
rect 248 238 249 239
rect 247 238 248 239
rect 246 238 247 239
rect 245 238 246 239
rect 244 238 245 239
rect 243 238 244 239
rect 242 238 243 239
rect 241 238 242 239
rect 240 238 241 239
rect 239 238 240 239
rect 238 238 239 239
rect 237 238 238 239
rect 236 238 237 239
rect 235 238 236 239
rect 234 238 235 239
rect 233 238 234 239
rect 232 238 233 239
rect 231 238 232 239
rect 230 238 231 239
rect 229 238 230 239
rect 228 238 229 239
rect 227 238 228 239
rect 226 238 227 239
rect 225 238 226 239
rect 224 238 225 239
rect 223 238 224 239
rect 222 238 223 239
rect 221 238 222 239
rect 220 238 221 239
rect 219 238 220 239
rect 218 238 219 239
rect 217 238 218 239
rect 216 238 217 239
rect 215 238 216 239
rect 214 238 215 239
rect 213 238 214 239
rect 212 238 213 239
rect 211 238 212 239
rect 210 238 211 239
rect 209 238 210 239
rect 208 238 209 239
rect 207 238 208 239
rect 206 238 207 239
rect 205 238 206 239
rect 204 238 205 239
rect 203 238 204 239
rect 202 238 203 239
rect 201 238 202 239
rect 200 238 201 239
rect 199 238 200 239
rect 198 238 199 239
rect 197 238 198 239
rect 196 238 197 239
rect 195 238 196 239
rect 194 238 195 239
rect 193 238 194 239
rect 192 238 193 239
rect 191 238 192 239
rect 190 238 191 239
rect 189 238 190 239
rect 188 238 189 239
rect 187 238 188 239
rect 186 238 187 239
rect 185 238 186 239
rect 184 238 185 239
rect 183 238 184 239
rect 182 238 183 239
rect 181 238 182 239
rect 180 238 181 239
rect 179 238 180 239
rect 178 238 179 239
rect 177 238 178 239
rect 176 238 177 239
rect 175 238 176 239
rect 148 238 149 239
rect 147 238 148 239
rect 146 238 147 239
rect 145 238 146 239
rect 144 238 145 239
rect 143 238 144 239
rect 142 238 143 239
rect 141 238 142 239
rect 140 238 141 239
rect 139 238 140 239
rect 138 238 139 239
rect 137 238 138 239
rect 136 238 137 239
rect 135 238 136 239
rect 134 238 135 239
rect 133 238 134 239
rect 132 238 133 239
rect 131 238 132 239
rect 130 238 131 239
rect 129 238 130 239
rect 128 238 129 239
rect 127 238 128 239
rect 126 238 127 239
rect 125 238 126 239
rect 124 238 125 239
rect 123 238 124 239
rect 122 238 123 239
rect 121 238 122 239
rect 120 238 121 239
rect 119 238 120 239
rect 118 238 119 239
rect 100 238 101 239
rect 99 238 100 239
rect 98 238 99 239
rect 97 238 98 239
rect 96 238 97 239
rect 95 238 96 239
rect 94 238 95 239
rect 93 238 94 239
rect 92 238 93 239
rect 91 238 92 239
rect 90 238 91 239
rect 89 238 90 239
rect 88 238 89 239
rect 87 238 88 239
rect 86 238 87 239
rect 85 238 86 239
rect 84 238 85 239
rect 83 238 84 239
rect 82 238 83 239
rect 81 238 82 239
rect 80 238 81 239
rect 79 238 80 239
rect 78 238 79 239
rect 77 238 78 239
rect 76 238 77 239
rect 75 238 76 239
rect 74 238 75 239
rect 73 238 74 239
rect 72 238 73 239
rect 71 238 72 239
rect 70 238 71 239
rect 69 238 70 239
rect 68 238 69 239
rect 67 238 68 239
rect 66 238 67 239
rect 65 238 66 239
rect 64 238 65 239
rect 63 238 64 239
rect 62 238 63 239
rect 61 238 62 239
rect 60 238 61 239
rect 59 238 60 239
rect 58 238 59 239
rect 57 238 58 239
rect 56 238 57 239
rect 55 238 56 239
rect 54 238 55 239
rect 53 238 54 239
rect 52 238 53 239
rect 51 238 52 239
rect 50 238 51 239
rect 49 238 50 239
rect 48 238 49 239
rect 47 238 48 239
rect 46 238 47 239
rect 45 238 46 239
rect 44 238 45 239
rect 43 238 44 239
rect 42 238 43 239
rect 41 238 42 239
rect 40 238 41 239
rect 39 238 40 239
rect 38 238 39 239
rect 37 238 38 239
rect 36 238 37 239
rect 35 238 36 239
rect 34 238 35 239
rect 33 238 34 239
rect 32 238 33 239
rect 31 238 32 239
rect 30 238 31 239
rect 29 238 30 239
rect 28 238 29 239
rect 27 238 28 239
rect 21 238 22 239
rect 20 238 21 239
rect 19 238 20 239
rect 18 238 19 239
rect 17 238 18 239
rect 16 238 17 239
rect 15 238 16 239
rect 14 238 15 239
rect 13 238 14 239
rect 12 238 13 239
rect 11 238 12 239
rect 10 238 11 239
rect 9 238 10 239
rect 8 238 9 239
rect 7 238 8 239
rect 6 238 7 239
rect 5 238 6 239
rect 4 238 5 239
rect 440 239 441 240
rect 439 239 440 240
rect 438 239 439 240
rect 437 239 438 240
rect 436 239 437 240
rect 435 239 436 240
rect 434 239 435 240
rect 424 239 425 240
rect 423 239 424 240
rect 422 239 423 240
rect 421 239 422 240
rect 420 239 421 240
rect 419 239 420 240
rect 418 239 419 240
rect 397 239 398 240
rect 396 239 397 240
rect 395 239 396 240
rect 394 239 395 240
rect 308 239 309 240
rect 307 239 308 240
rect 306 239 307 240
rect 305 239 306 240
rect 304 239 305 240
rect 303 239 304 240
rect 302 239 303 240
rect 301 239 302 240
rect 300 239 301 240
rect 299 239 300 240
rect 298 239 299 240
rect 297 239 298 240
rect 296 239 297 240
rect 295 239 296 240
rect 294 239 295 240
rect 293 239 294 240
rect 292 239 293 240
rect 269 239 270 240
rect 268 239 269 240
rect 267 239 268 240
rect 266 239 267 240
rect 265 239 266 240
rect 264 239 265 240
rect 263 239 264 240
rect 262 239 263 240
rect 261 239 262 240
rect 260 239 261 240
rect 259 239 260 240
rect 258 239 259 240
rect 257 239 258 240
rect 256 239 257 240
rect 255 239 256 240
rect 254 239 255 240
rect 253 239 254 240
rect 252 239 253 240
rect 251 239 252 240
rect 250 239 251 240
rect 249 239 250 240
rect 248 239 249 240
rect 247 239 248 240
rect 246 239 247 240
rect 245 239 246 240
rect 244 239 245 240
rect 243 239 244 240
rect 242 239 243 240
rect 241 239 242 240
rect 240 239 241 240
rect 239 239 240 240
rect 238 239 239 240
rect 237 239 238 240
rect 236 239 237 240
rect 235 239 236 240
rect 234 239 235 240
rect 233 239 234 240
rect 232 239 233 240
rect 231 239 232 240
rect 230 239 231 240
rect 229 239 230 240
rect 228 239 229 240
rect 227 239 228 240
rect 226 239 227 240
rect 225 239 226 240
rect 224 239 225 240
rect 223 239 224 240
rect 222 239 223 240
rect 221 239 222 240
rect 220 239 221 240
rect 219 239 220 240
rect 218 239 219 240
rect 217 239 218 240
rect 216 239 217 240
rect 215 239 216 240
rect 214 239 215 240
rect 213 239 214 240
rect 212 239 213 240
rect 211 239 212 240
rect 210 239 211 240
rect 209 239 210 240
rect 208 239 209 240
rect 207 239 208 240
rect 206 239 207 240
rect 205 239 206 240
rect 204 239 205 240
rect 203 239 204 240
rect 202 239 203 240
rect 201 239 202 240
rect 200 239 201 240
rect 199 239 200 240
rect 198 239 199 240
rect 197 239 198 240
rect 196 239 197 240
rect 195 239 196 240
rect 194 239 195 240
rect 193 239 194 240
rect 192 239 193 240
rect 191 239 192 240
rect 190 239 191 240
rect 189 239 190 240
rect 188 239 189 240
rect 187 239 188 240
rect 186 239 187 240
rect 185 239 186 240
rect 184 239 185 240
rect 183 239 184 240
rect 182 239 183 240
rect 181 239 182 240
rect 180 239 181 240
rect 179 239 180 240
rect 178 239 179 240
rect 177 239 178 240
rect 176 239 177 240
rect 148 239 149 240
rect 147 239 148 240
rect 146 239 147 240
rect 145 239 146 240
rect 144 239 145 240
rect 143 239 144 240
rect 142 239 143 240
rect 141 239 142 240
rect 140 239 141 240
rect 139 239 140 240
rect 138 239 139 240
rect 137 239 138 240
rect 136 239 137 240
rect 135 239 136 240
rect 134 239 135 240
rect 133 239 134 240
rect 132 239 133 240
rect 131 239 132 240
rect 130 239 131 240
rect 129 239 130 240
rect 128 239 129 240
rect 127 239 128 240
rect 126 239 127 240
rect 125 239 126 240
rect 124 239 125 240
rect 123 239 124 240
rect 122 239 123 240
rect 121 239 122 240
rect 120 239 121 240
rect 119 239 120 240
rect 118 239 119 240
rect 101 239 102 240
rect 100 239 101 240
rect 99 239 100 240
rect 98 239 99 240
rect 97 239 98 240
rect 96 239 97 240
rect 95 239 96 240
rect 94 239 95 240
rect 93 239 94 240
rect 92 239 93 240
rect 91 239 92 240
rect 90 239 91 240
rect 89 239 90 240
rect 88 239 89 240
rect 87 239 88 240
rect 86 239 87 240
rect 85 239 86 240
rect 84 239 85 240
rect 83 239 84 240
rect 82 239 83 240
rect 81 239 82 240
rect 80 239 81 240
rect 79 239 80 240
rect 78 239 79 240
rect 77 239 78 240
rect 76 239 77 240
rect 75 239 76 240
rect 74 239 75 240
rect 73 239 74 240
rect 72 239 73 240
rect 71 239 72 240
rect 70 239 71 240
rect 69 239 70 240
rect 68 239 69 240
rect 67 239 68 240
rect 66 239 67 240
rect 65 239 66 240
rect 64 239 65 240
rect 63 239 64 240
rect 62 239 63 240
rect 61 239 62 240
rect 60 239 61 240
rect 59 239 60 240
rect 58 239 59 240
rect 57 239 58 240
rect 56 239 57 240
rect 55 239 56 240
rect 54 239 55 240
rect 53 239 54 240
rect 52 239 53 240
rect 51 239 52 240
rect 50 239 51 240
rect 49 239 50 240
rect 48 239 49 240
rect 47 239 48 240
rect 46 239 47 240
rect 45 239 46 240
rect 44 239 45 240
rect 43 239 44 240
rect 42 239 43 240
rect 41 239 42 240
rect 40 239 41 240
rect 39 239 40 240
rect 38 239 39 240
rect 37 239 38 240
rect 36 239 37 240
rect 35 239 36 240
rect 34 239 35 240
rect 33 239 34 240
rect 32 239 33 240
rect 31 239 32 240
rect 30 239 31 240
rect 29 239 30 240
rect 28 239 29 240
rect 21 239 22 240
rect 20 239 21 240
rect 19 239 20 240
rect 18 239 19 240
rect 17 239 18 240
rect 16 239 17 240
rect 15 239 16 240
rect 14 239 15 240
rect 13 239 14 240
rect 12 239 13 240
rect 11 239 12 240
rect 10 239 11 240
rect 9 239 10 240
rect 8 239 9 240
rect 7 239 8 240
rect 6 239 7 240
rect 5 239 6 240
rect 4 239 5 240
rect 440 240 441 241
rect 439 240 440 241
rect 438 240 439 241
rect 437 240 438 241
rect 436 240 437 241
rect 435 240 436 241
rect 434 240 435 241
rect 433 240 434 241
rect 432 240 433 241
rect 431 240 432 241
rect 430 240 431 241
rect 429 240 430 241
rect 428 240 429 241
rect 427 240 428 241
rect 426 240 427 241
rect 425 240 426 241
rect 424 240 425 241
rect 423 240 424 241
rect 422 240 423 241
rect 421 240 422 241
rect 420 240 421 241
rect 419 240 420 241
rect 418 240 419 241
rect 398 240 399 241
rect 397 240 398 241
rect 396 240 397 241
rect 395 240 396 241
rect 394 240 395 241
rect 316 240 317 241
rect 315 240 316 241
rect 314 240 315 241
rect 313 240 314 241
rect 312 240 313 241
rect 311 240 312 241
rect 310 240 311 241
rect 309 240 310 241
rect 308 240 309 241
rect 307 240 308 241
rect 306 240 307 241
rect 305 240 306 241
rect 304 240 305 241
rect 303 240 304 241
rect 302 240 303 241
rect 301 240 302 241
rect 300 240 301 241
rect 299 240 300 241
rect 298 240 299 241
rect 297 240 298 241
rect 296 240 297 241
rect 295 240 296 241
rect 294 240 295 241
rect 293 240 294 241
rect 292 240 293 241
rect 291 240 292 241
rect 290 240 291 241
rect 289 240 290 241
rect 288 240 289 241
rect 287 240 288 241
rect 286 240 287 241
rect 285 240 286 241
rect 268 240 269 241
rect 267 240 268 241
rect 266 240 267 241
rect 265 240 266 241
rect 264 240 265 241
rect 263 240 264 241
rect 262 240 263 241
rect 261 240 262 241
rect 260 240 261 241
rect 259 240 260 241
rect 258 240 259 241
rect 257 240 258 241
rect 256 240 257 241
rect 255 240 256 241
rect 254 240 255 241
rect 253 240 254 241
rect 252 240 253 241
rect 251 240 252 241
rect 250 240 251 241
rect 249 240 250 241
rect 248 240 249 241
rect 247 240 248 241
rect 246 240 247 241
rect 245 240 246 241
rect 244 240 245 241
rect 243 240 244 241
rect 242 240 243 241
rect 241 240 242 241
rect 240 240 241 241
rect 239 240 240 241
rect 238 240 239 241
rect 237 240 238 241
rect 236 240 237 241
rect 235 240 236 241
rect 234 240 235 241
rect 233 240 234 241
rect 232 240 233 241
rect 231 240 232 241
rect 230 240 231 241
rect 229 240 230 241
rect 228 240 229 241
rect 227 240 228 241
rect 226 240 227 241
rect 225 240 226 241
rect 224 240 225 241
rect 223 240 224 241
rect 222 240 223 241
rect 221 240 222 241
rect 220 240 221 241
rect 219 240 220 241
rect 218 240 219 241
rect 217 240 218 241
rect 216 240 217 241
rect 215 240 216 241
rect 214 240 215 241
rect 213 240 214 241
rect 212 240 213 241
rect 211 240 212 241
rect 210 240 211 241
rect 209 240 210 241
rect 208 240 209 241
rect 207 240 208 241
rect 206 240 207 241
rect 205 240 206 241
rect 204 240 205 241
rect 203 240 204 241
rect 202 240 203 241
rect 201 240 202 241
rect 200 240 201 241
rect 199 240 200 241
rect 198 240 199 241
rect 197 240 198 241
rect 196 240 197 241
rect 195 240 196 241
rect 194 240 195 241
rect 193 240 194 241
rect 192 240 193 241
rect 191 240 192 241
rect 190 240 191 241
rect 189 240 190 241
rect 188 240 189 241
rect 187 240 188 241
rect 186 240 187 241
rect 185 240 186 241
rect 184 240 185 241
rect 183 240 184 241
rect 182 240 183 241
rect 181 240 182 241
rect 180 240 181 241
rect 179 240 180 241
rect 149 240 150 241
rect 148 240 149 241
rect 147 240 148 241
rect 146 240 147 241
rect 145 240 146 241
rect 144 240 145 241
rect 143 240 144 241
rect 142 240 143 241
rect 141 240 142 241
rect 140 240 141 241
rect 139 240 140 241
rect 138 240 139 241
rect 137 240 138 241
rect 136 240 137 241
rect 135 240 136 241
rect 134 240 135 241
rect 133 240 134 241
rect 132 240 133 241
rect 131 240 132 241
rect 130 240 131 241
rect 129 240 130 241
rect 128 240 129 241
rect 127 240 128 241
rect 126 240 127 241
rect 125 240 126 241
rect 124 240 125 241
rect 123 240 124 241
rect 122 240 123 241
rect 121 240 122 241
rect 120 240 121 241
rect 119 240 120 241
rect 118 240 119 241
rect 102 240 103 241
rect 101 240 102 241
rect 100 240 101 241
rect 99 240 100 241
rect 98 240 99 241
rect 97 240 98 241
rect 96 240 97 241
rect 95 240 96 241
rect 94 240 95 241
rect 93 240 94 241
rect 92 240 93 241
rect 91 240 92 241
rect 90 240 91 241
rect 89 240 90 241
rect 88 240 89 241
rect 87 240 88 241
rect 86 240 87 241
rect 85 240 86 241
rect 84 240 85 241
rect 83 240 84 241
rect 82 240 83 241
rect 81 240 82 241
rect 80 240 81 241
rect 79 240 80 241
rect 78 240 79 241
rect 77 240 78 241
rect 76 240 77 241
rect 75 240 76 241
rect 74 240 75 241
rect 73 240 74 241
rect 72 240 73 241
rect 71 240 72 241
rect 70 240 71 241
rect 69 240 70 241
rect 68 240 69 241
rect 67 240 68 241
rect 66 240 67 241
rect 65 240 66 241
rect 64 240 65 241
rect 63 240 64 241
rect 62 240 63 241
rect 61 240 62 241
rect 60 240 61 241
rect 59 240 60 241
rect 58 240 59 241
rect 57 240 58 241
rect 56 240 57 241
rect 55 240 56 241
rect 54 240 55 241
rect 53 240 54 241
rect 52 240 53 241
rect 51 240 52 241
rect 50 240 51 241
rect 49 240 50 241
rect 48 240 49 241
rect 47 240 48 241
rect 46 240 47 241
rect 45 240 46 241
rect 44 240 45 241
rect 43 240 44 241
rect 42 240 43 241
rect 41 240 42 241
rect 40 240 41 241
rect 39 240 40 241
rect 38 240 39 241
rect 37 240 38 241
rect 36 240 37 241
rect 35 240 36 241
rect 34 240 35 241
rect 33 240 34 241
rect 32 240 33 241
rect 31 240 32 241
rect 30 240 31 241
rect 29 240 30 241
rect 28 240 29 241
rect 21 240 22 241
rect 20 240 21 241
rect 19 240 20 241
rect 18 240 19 241
rect 17 240 18 241
rect 16 240 17 241
rect 15 240 16 241
rect 14 240 15 241
rect 13 240 14 241
rect 12 240 13 241
rect 11 240 12 241
rect 10 240 11 241
rect 9 240 10 241
rect 8 240 9 241
rect 7 240 8 241
rect 6 240 7 241
rect 5 240 6 241
rect 4 240 5 241
rect 3 240 4 241
rect 439 241 440 242
rect 438 241 439 242
rect 437 241 438 242
rect 436 241 437 242
rect 435 241 436 242
rect 434 241 435 242
rect 433 241 434 242
rect 432 241 433 242
rect 431 241 432 242
rect 430 241 431 242
rect 429 241 430 242
rect 428 241 429 242
rect 427 241 428 242
rect 426 241 427 242
rect 425 241 426 242
rect 424 241 425 242
rect 423 241 424 242
rect 422 241 423 242
rect 421 241 422 242
rect 420 241 421 242
rect 419 241 420 242
rect 418 241 419 242
rect 399 241 400 242
rect 398 241 399 242
rect 397 241 398 242
rect 396 241 397 242
rect 395 241 396 242
rect 320 241 321 242
rect 319 241 320 242
rect 318 241 319 242
rect 317 241 318 242
rect 316 241 317 242
rect 315 241 316 242
rect 314 241 315 242
rect 313 241 314 242
rect 312 241 313 242
rect 311 241 312 242
rect 310 241 311 242
rect 309 241 310 242
rect 308 241 309 242
rect 307 241 308 242
rect 306 241 307 242
rect 305 241 306 242
rect 304 241 305 242
rect 303 241 304 242
rect 302 241 303 242
rect 301 241 302 242
rect 300 241 301 242
rect 299 241 300 242
rect 298 241 299 242
rect 297 241 298 242
rect 296 241 297 242
rect 295 241 296 242
rect 294 241 295 242
rect 293 241 294 242
rect 292 241 293 242
rect 291 241 292 242
rect 290 241 291 242
rect 289 241 290 242
rect 288 241 289 242
rect 287 241 288 242
rect 286 241 287 242
rect 285 241 286 242
rect 284 241 285 242
rect 283 241 284 242
rect 282 241 283 242
rect 281 241 282 242
rect 280 241 281 242
rect 267 241 268 242
rect 266 241 267 242
rect 265 241 266 242
rect 264 241 265 242
rect 263 241 264 242
rect 262 241 263 242
rect 261 241 262 242
rect 260 241 261 242
rect 259 241 260 242
rect 258 241 259 242
rect 257 241 258 242
rect 256 241 257 242
rect 255 241 256 242
rect 254 241 255 242
rect 253 241 254 242
rect 252 241 253 242
rect 251 241 252 242
rect 250 241 251 242
rect 249 241 250 242
rect 248 241 249 242
rect 247 241 248 242
rect 246 241 247 242
rect 245 241 246 242
rect 244 241 245 242
rect 243 241 244 242
rect 242 241 243 242
rect 241 241 242 242
rect 240 241 241 242
rect 239 241 240 242
rect 238 241 239 242
rect 237 241 238 242
rect 236 241 237 242
rect 235 241 236 242
rect 234 241 235 242
rect 233 241 234 242
rect 232 241 233 242
rect 231 241 232 242
rect 230 241 231 242
rect 229 241 230 242
rect 228 241 229 242
rect 227 241 228 242
rect 226 241 227 242
rect 225 241 226 242
rect 224 241 225 242
rect 223 241 224 242
rect 222 241 223 242
rect 221 241 222 242
rect 220 241 221 242
rect 219 241 220 242
rect 218 241 219 242
rect 217 241 218 242
rect 216 241 217 242
rect 215 241 216 242
rect 214 241 215 242
rect 213 241 214 242
rect 212 241 213 242
rect 211 241 212 242
rect 210 241 211 242
rect 209 241 210 242
rect 208 241 209 242
rect 207 241 208 242
rect 206 241 207 242
rect 205 241 206 242
rect 204 241 205 242
rect 203 241 204 242
rect 202 241 203 242
rect 201 241 202 242
rect 200 241 201 242
rect 199 241 200 242
rect 198 241 199 242
rect 197 241 198 242
rect 196 241 197 242
rect 195 241 196 242
rect 194 241 195 242
rect 193 241 194 242
rect 192 241 193 242
rect 191 241 192 242
rect 190 241 191 242
rect 189 241 190 242
rect 188 241 189 242
rect 187 241 188 242
rect 186 241 187 242
rect 185 241 186 242
rect 184 241 185 242
rect 183 241 184 242
rect 182 241 183 242
rect 181 241 182 242
rect 150 241 151 242
rect 149 241 150 242
rect 148 241 149 242
rect 147 241 148 242
rect 146 241 147 242
rect 145 241 146 242
rect 144 241 145 242
rect 143 241 144 242
rect 142 241 143 242
rect 141 241 142 242
rect 140 241 141 242
rect 139 241 140 242
rect 138 241 139 242
rect 137 241 138 242
rect 136 241 137 242
rect 135 241 136 242
rect 134 241 135 242
rect 133 241 134 242
rect 132 241 133 242
rect 131 241 132 242
rect 130 241 131 242
rect 129 241 130 242
rect 128 241 129 242
rect 127 241 128 242
rect 126 241 127 242
rect 125 241 126 242
rect 124 241 125 242
rect 123 241 124 242
rect 122 241 123 242
rect 121 241 122 242
rect 120 241 121 242
rect 119 241 120 242
rect 103 241 104 242
rect 102 241 103 242
rect 101 241 102 242
rect 100 241 101 242
rect 99 241 100 242
rect 98 241 99 242
rect 97 241 98 242
rect 96 241 97 242
rect 95 241 96 242
rect 94 241 95 242
rect 93 241 94 242
rect 92 241 93 242
rect 91 241 92 242
rect 90 241 91 242
rect 89 241 90 242
rect 88 241 89 242
rect 87 241 88 242
rect 86 241 87 242
rect 85 241 86 242
rect 84 241 85 242
rect 83 241 84 242
rect 82 241 83 242
rect 81 241 82 242
rect 80 241 81 242
rect 79 241 80 242
rect 78 241 79 242
rect 77 241 78 242
rect 76 241 77 242
rect 75 241 76 242
rect 74 241 75 242
rect 73 241 74 242
rect 72 241 73 242
rect 71 241 72 242
rect 70 241 71 242
rect 69 241 70 242
rect 68 241 69 242
rect 67 241 68 242
rect 66 241 67 242
rect 65 241 66 242
rect 64 241 65 242
rect 63 241 64 242
rect 62 241 63 242
rect 61 241 62 242
rect 60 241 61 242
rect 59 241 60 242
rect 58 241 59 242
rect 57 241 58 242
rect 56 241 57 242
rect 55 241 56 242
rect 54 241 55 242
rect 53 241 54 242
rect 52 241 53 242
rect 51 241 52 242
rect 50 241 51 242
rect 49 241 50 242
rect 48 241 49 242
rect 47 241 48 242
rect 46 241 47 242
rect 45 241 46 242
rect 44 241 45 242
rect 43 241 44 242
rect 42 241 43 242
rect 41 241 42 242
rect 40 241 41 242
rect 39 241 40 242
rect 38 241 39 242
rect 37 241 38 242
rect 36 241 37 242
rect 35 241 36 242
rect 34 241 35 242
rect 33 241 34 242
rect 32 241 33 242
rect 31 241 32 242
rect 30 241 31 242
rect 29 241 30 242
rect 28 241 29 242
rect 21 241 22 242
rect 20 241 21 242
rect 19 241 20 242
rect 18 241 19 242
rect 17 241 18 242
rect 16 241 17 242
rect 15 241 16 242
rect 14 241 15 242
rect 13 241 14 242
rect 12 241 13 242
rect 11 241 12 242
rect 10 241 11 242
rect 9 241 10 242
rect 8 241 9 242
rect 7 241 8 242
rect 6 241 7 242
rect 5 241 6 242
rect 4 241 5 242
rect 3 241 4 242
rect 439 242 440 243
rect 438 242 439 243
rect 437 242 438 243
rect 436 242 437 243
rect 435 242 436 243
rect 434 242 435 243
rect 433 242 434 243
rect 432 242 433 243
rect 431 242 432 243
rect 430 242 431 243
rect 429 242 430 243
rect 428 242 429 243
rect 427 242 428 243
rect 426 242 427 243
rect 425 242 426 243
rect 424 242 425 243
rect 423 242 424 243
rect 422 242 423 243
rect 421 242 422 243
rect 420 242 421 243
rect 419 242 420 243
rect 418 242 419 243
rect 400 242 401 243
rect 399 242 400 243
rect 398 242 399 243
rect 397 242 398 243
rect 396 242 397 243
rect 395 242 396 243
rect 324 242 325 243
rect 323 242 324 243
rect 322 242 323 243
rect 321 242 322 243
rect 320 242 321 243
rect 319 242 320 243
rect 318 242 319 243
rect 317 242 318 243
rect 316 242 317 243
rect 315 242 316 243
rect 314 242 315 243
rect 313 242 314 243
rect 312 242 313 243
rect 311 242 312 243
rect 310 242 311 243
rect 309 242 310 243
rect 308 242 309 243
rect 307 242 308 243
rect 306 242 307 243
rect 305 242 306 243
rect 304 242 305 243
rect 303 242 304 243
rect 302 242 303 243
rect 301 242 302 243
rect 300 242 301 243
rect 299 242 300 243
rect 298 242 299 243
rect 297 242 298 243
rect 296 242 297 243
rect 295 242 296 243
rect 294 242 295 243
rect 293 242 294 243
rect 292 242 293 243
rect 291 242 292 243
rect 290 242 291 243
rect 289 242 290 243
rect 288 242 289 243
rect 287 242 288 243
rect 286 242 287 243
rect 285 242 286 243
rect 284 242 285 243
rect 283 242 284 243
rect 282 242 283 243
rect 281 242 282 243
rect 280 242 281 243
rect 279 242 280 243
rect 278 242 279 243
rect 277 242 278 243
rect 276 242 277 243
rect 267 242 268 243
rect 266 242 267 243
rect 265 242 266 243
rect 264 242 265 243
rect 263 242 264 243
rect 262 242 263 243
rect 261 242 262 243
rect 260 242 261 243
rect 259 242 260 243
rect 258 242 259 243
rect 257 242 258 243
rect 256 242 257 243
rect 255 242 256 243
rect 254 242 255 243
rect 253 242 254 243
rect 252 242 253 243
rect 251 242 252 243
rect 250 242 251 243
rect 249 242 250 243
rect 248 242 249 243
rect 247 242 248 243
rect 246 242 247 243
rect 245 242 246 243
rect 244 242 245 243
rect 243 242 244 243
rect 242 242 243 243
rect 241 242 242 243
rect 240 242 241 243
rect 239 242 240 243
rect 238 242 239 243
rect 237 242 238 243
rect 236 242 237 243
rect 235 242 236 243
rect 234 242 235 243
rect 233 242 234 243
rect 232 242 233 243
rect 228 242 229 243
rect 227 242 228 243
rect 226 242 227 243
rect 225 242 226 243
rect 224 242 225 243
rect 223 242 224 243
rect 222 242 223 243
rect 221 242 222 243
rect 220 242 221 243
rect 219 242 220 243
rect 218 242 219 243
rect 217 242 218 243
rect 216 242 217 243
rect 215 242 216 243
rect 214 242 215 243
rect 213 242 214 243
rect 212 242 213 243
rect 211 242 212 243
rect 210 242 211 243
rect 209 242 210 243
rect 208 242 209 243
rect 207 242 208 243
rect 206 242 207 243
rect 205 242 206 243
rect 204 242 205 243
rect 203 242 204 243
rect 202 242 203 243
rect 201 242 202 243
rect 200 242 201 243
rect 199 242 200 243
rect 198 242 199 243
rect 197 242 198 243
rect 196 242 197 243
rect 195 242 196 243
rect 194 242 195 243
rect 193 242 194 243
rect 192 242 193 243
rect 191 242 192 243
rect 190 242 191 243
rect 189 242 190 243
rect 188 242 189 243
rect 187 242 188 243
rect 186 242 187 243
rect 185 242 186 243
rect 184 242 185 243
rect 150 242 151 243
rect 149 242 150 243
rect 148 242 149 243
rect 147 242 148 243
rect 146 242 147 243
rect 145 242 146 243
rect 144 242 145 243
rect 143 242 144 243
rect 142 242 143 243
rect 141 242 142 243
rect 140 242 141 243
rect 139 242 140 243
rect 138 242 139 243
rect 137 242 138 243
rect 136 242 137 243
rect 135 242 136 243
rect 134 242 135 243
rect 133 242 134 243
rect 132 242 133 243
rect 131 242 132 243
rect 130 242 131 243
rect 129 242 130 243
rect 128 242 129 243
rect 127 242 128 243
rect 126 242 127 243
rect 125 242 126 243
rect 124 242 125 243
rect 123 242 124 243
rect 122 242 123 243
rect 121 242 122 243
rect 120 242 121 243
rect 119 242 120 243
rect 104 242 105 243
rect 103 242 104 243
rect 102 242 103 243
rect 101 242 102 243
rect 100 242 101 243
rect 99 242 100 243
rect 98 242 99 243
rect 97 242 98 243
rect 96 242 97 243
rect 95 242 96 243
rect 94 242 95 243
rect 93 242 94 243
rect 92 242 93 243
rect 91 242 92 243
rect 90 242 91 243
rect 89 242 90 243
rect 88 242 89 243
rect 87 242 88 243
rect 86 242 87 243
rect 85 242 86 243
rect 84 242 85 243
rect 83 242 84 243
rect 82 242 83 243
rect 81 242 82 243
rect 80 242 81 243
rect 79 242 80 243
rect 78 242 79 243
rect 77 242 78 243
rect 76 242 77 243
rect 75 242 76 243
rect 74 242 75 243
rect 73 242 74 243
rect 72 242 73 243
rect 71 242 72 243
rect 70 242 71 243
rect 69 242 70 243
rect 68 242 69 243
rect 67 242 68 243
rect 66 242 67 243
rect 65 242 66 243
rect 64 242 65 243
rect 63 242 64 243
rect 62 242 63 243
rect 61 242 62 243
rect 60 242 61 243
rect 59 242 60 243
rect 58 242 59 243
rect 57 242 58 243
rect 56 242 57 243
rect 55 242 56 243
rect 54 242 55 243
rect 53 242 54 243
rect 52 242 53 243
rect 51 242 52 243
rect 50 242 51 243
rect 49 242 50 243
rect 48 242 49 243
rect 47 242 48 243
rect 46 242 47 243
rect 45 242 46 243
rect 44 242 45 243
rect 43 242 44 243
rect 42 242 43 243
rect 41 242 42 243
rect 40 242 41 243
rect 39 242 40 243
rect 38 242 39 243
rect 37 242 38 243
rect 36 242 37 243
rect 35 242 36 243
rect 34 242 35 243
rect 33 242 34 243
rect 32 242 33 243
rect 31 242 32 243
rect 30 242 31 243
rect 29 242 30 243
rect 21 242 22 243
rect 20 242 21 243
rect 19 242 20 243
rect 18 242 19 243
rect 17 242 18 243
rect 16 242 17 243
rect 15 242 16 243
rect 14 242 15 243
rect 13 242 14 243
rect 12 242 13 243
rect 11 242 12 243
rect 10 242 11 243
rect 9 242 10 243
rect 8 242 9 243
rect 7 242 8 243
rect 6 242 7 243
rect 5 242 6 243
rect 4 242 5 243
rect 3 242 4 243
rect 439 243 440 244
rect 438 243 439 244
rect 437 243 438 244
rect 436 243 437 244
rect 435 243 436 244
rect 434 243 435 244
rect 433 243 434 244
rect 432 243 433 244
rect 431 243 432 244
rect 430 243 431 244
rect 429 243 430 244
rect 428 243 429 244
rect 427 243 428 244
rect 426 243 427 244
rect 425 243 426 244
rect 424 243 425 244
rect 423 243 424 244
rect 422 243 423 244
rect 421 243 422 244
rect 420 243 421 244
rect 419 243 420 244
rect 418 243 419 244
rect 401 243 402 244
rect 400 243 401 244
rect 399 243 400 244
rect 398 243 399 244
rect 397 243 398 244
rect 396 243 397 244
rect 395 243 396 244
rect 327 243 328 244
rect 326 243 327 244
rect 325 243 326 244
rect 324 243 325 244
rect 323 243 324 244
rect 322 243 323 244
rect 321 243 322 244
rect 320 243 321 244
rect 319 243 320 244
rect 318 243 319 244
rect 317 243 318 244
rect 316 243 317 244
rect 315 243 316 244
rect 314 243 315 244
rect 313 243 314 244
rect 312 243 313 244
rect 311 243 312 244
rect 310 243 311 244
rect 309 243 310 244
rect 308 243 309 244
rect 307 243 308 244
rect 306 243 307 244
rect 305 243 306 244
rect 304 243 305 244
rect 303 243 304 244
rect 302 243 303 244
rect 301 243 302 244
rect 300 243 301 244
rect 299 243 300 244
rect 298 243 299 244
rect 297 243 298 244
rect 296 243 297 244
rect 295 243 296 244
rect 294 243 295 244
rect 293 243 294 244
rect 292 243 293 244
rect 291 243 292 244
rect 290 243 291 244
rect 289 243 290 244
rect 288 243 289 244
rect 287 243 288 244
rect 286 243 287 244
rect 285 243 286 244
rect 284 243 285 244
rect 283 243 284 244
rect 282 243 283 244
rect 281 243 282 244
rect 280 243 281 244
rect 279 243 280 244
rect 278 243 279 244
rect 277 243 278 244
rect 276 243 277 244
rect 275 243 276 244
rect 274 243 275 244
rect 273 243 274 244
rect 266 243 267 244
rect 265 243 266 244
rect 264 243 265 244
rect 263 243 264 244
rect 262 243 263 244
rect 261 243 262 244
rect 260 243 261 244
rect 259 243 260 244
rect 258 243 259 244
rect 257 243 258 244
rect 256 243 257 244
rect 255 243 256 244
rect 254 243 255 244
rect 253 243 254 244
rect 252 243 253 244
rect 251 243 252 244
rect 250 243 251 244
rect 249 243 250 244
rect 248 243 249 244
rect 247 243 248 244
rect 246 243 247 244
rect 245 243 246 244
rect 244 243 245 244
rect 243 243 244 244
rect 242 243 243 244
rect 241 243 242 244
rect 240 243 241 244
rect 239 243 240 244
rect 238 243 239 244
rect 237 243 238 244
rect 236 243 237 244
rect 235 243 236 244
rect 234 243 235 244
rect 233 243 234 244
rect 232 243 233 244
rect 224 243 225 244
rect 223 243 224 244
rect 222 243 223 244
rect 221 243 222 244
rect 220 243 221 244
rect 219 243 220 244
rect 218 243 219 244
rect 217 243 218 244
rect 216 243 217 244
rect 215 243 216 244
rect 214 243 215 244
rect 213 243 214 244
rect 212 243 213 244
rect 211 243 212 244
rect 210 243 211 244
rect 209 243 210 244
rect 208 243 209 244
rect 207 243 208 244
rect 206 243 207 244
rect 205 243 206 244
rect 204 243 205 244
rect 203 243 204 244
rect 202 243 203 244
rect 201 243 202 244
rect 200 243 201 244
rect 199 243 200 244
rect 198 243 199 244
rect 197 243 198 244
rect 196 243 197 244
rect 195 243 196 244
rect 194 243 195 244
rect 193 243 194 244
rect 192 243 193 244
rect 191 243 192 244
rect 190 243 191 244
rect 189 243 190 244
rect 188 243 189 244
rect 187 243 188 244
rect 151 243 152 244
rect 150 243 151 244
rect 149 243 150 244
rect 148 243 149 244
rect 147 243 148 244
rect 146 243 147 244
rect 145 243 146 244
rect 144 243 145 244
rect 143 243 144 244
rect 142 243 143 244
rect 141 243 142 244
rect 140 243 141 244
rect 139 243 140 244
rect 138 243 139 244
rect 137 243 138 244
rect 136 243 137 244
rect 135 243 136 244
rect 134 243 135 244
rect 133 243 134 244
rect 132 243 133 244
rect 131 243 132 244
rect 130 243 131 244
rect 129 243 130 244
rect 128 243 129 244
rect 127 243 128 244
rect 126 243 127 244
rect 125 243 126 244
rect 124 243 125 244
rect 123 243 124 244
rect 122 243 123 244
rect 121 243 122 244
rect 120 243 121 244
rect 119 243 120 244
rect 104 243 105 244
rect 103 243 104 244
rect 102 243 103 244
rect 101 243 102 244
rect 100 243 101 244
rect 99 243 100 244
rect 98 243 99 244
rect 97 243 98 244
rect 96 243 97 244
rect 95 243 96 244
rect 94 243 95 244
rect 93 243 94 244
rect 92 243 93 244
rect 91 243 92 244
rect 90 243 91 244
rect 89 243 90 244
rect 88 243 89 244
rect 87 243 88 244
rect 86 243 87 244
rect 85 243 86 244
rect 84 243 85 244
rect 83 243 84 244
rect 82 243 83 244
rect 81 243 82 244
rect 80 243 81 244
rect 79 243 80 244
rect 78 243 79 244
rect 77 243 78 244
rect 76 243 77 244
rect 75 243 76 244
rect 74 243 75 244
rect 73 243 74 244
rect 72 243 73 244
rect 71 243 72 244
rect 70 243 71 244
rect 69 243 70 244
rect 68 243 69 244
rect 67 243 68 244
rect 66 243 67 244
rect 65 243 66 244
rect 64 243 65 244
rect 63 243 64 244
rect 62 243 63 244
rect 61 243 62 244
rect 60 243 61 244
rect 59 243 60 244
rect 58 243 59 244
rect 57 243 58 244
rect 56 243 57 244
rect 55 243 56 244
rect 54 243 55 244
rect 53 243 54 244
rect 52 243 53 244
rect 51 243 52 244
rect 50 243 51 244
rect 49 243 50 244
rect 48 243 49 244
rect 47 243 48 244
rect 46 243 47 244
rect 45 243 46 244
rect 44 243 45 244
rect 43 243 44 244
rect 42 243 43 244
rect 41 243 42 244
rect 40 243 41 244
rect 39 243 40 244
rect 38 243 39 244
rect 37 243 38 244
rect 36 243 37 244
rect 35 243 36 244
rect 34 243 35 244
rect 33 243 34 244
rect 32 243 33 244
rect 31 243 32 244
rect 30 243 31 244
rect 29 243 30 244
rect 21 243 22 244
rect 20 243 21 244
rect 19 243 20 244
rect 18 243 19 244
rect 17 243 18 244
rect 16 243 17 244
rect 15 243 16 244
rect 14 243 15 244
rect 13 243 14 244
rect 12 243 13 244
rect 11 243 12 244
rect 10 243 11 244
rect 9 243 10 244
rect 8 243 9 244
rect 7 243 8 244
rect 6 243 7 244
rect 5 243 6 244
rect 4 243 5 244
rect 3 243 4 244
rect 479 244 480 245
rect 478 244 479 245
rect 477 244 478 245
rect 476 244 477 245
rect 475 244 476 245
rect 466 244 467 245
rect 465 244 466 245
rect 464 244 465 245
rect 439 244 440 245
rect 438 244 439 245
rect 437 244 438 245
rect 436 244 437 245
rect 435 244 436 245
rect 434 244 435 245
rect 433 244 434 245
rect 432 244 433 245
rect 431 244 432 245
rect 430 244 431 245
rect 429 244 430 245
rect 428 244 429 245
rect 427 244 428 245
rect 426 244 427 245
rect 425 244 426 245
rect 424 244 425 245
rect 423 244 424 245
rect 422 244 423 245
rect 421 244 422 245
rect 420 244 421 245
rect 419 244 420 245
rect 418 244 419 245
rect 402 244 403 245
rect 401 244 402 245
rect 400 244 401 245
rect 399 244 400 245
rect 398 244 399 245
rect 397 244 398 245
rect 396 244 397 245
rect 395 244 396 245
rect 327 244 328 245
rect 326 244 327 245
rect 325 244 326 245
rect 324 244 325 245
rect 323 244 324 245
rect 322 244 323 245
rect 321 244 322 245
rect 320 244 321 245
rect 319 244 320 245
rect 318 244 319 245
rect 317 244 318 245
rect 316 244 317 245
rect 315 244 316 245
rect 314 244 315 245
rect 313 244 314 245
rect 312 244 313 245
rect 311 244 312 245
rect 310 244 311 245
rect 309 244 310 245
rect 308 244 309 245
rect 307 244 308 245
rect 306 244 307 245
rect 305 244 306 245
rect 304 244 305 245
rect 303 244 304 245
rect 302 244 303 245
rect 301 244 302 245
rect 300 244 301 245
rect 299 244 300 245
rect 298 244 299 245
rect 297 244 298 245
rect 296 244 297 245
rect 295 244 296 245
rect 294 244 295 245
rect 293 244 294 245
rect 292 244 293 245
rect 291 244 292 245
rect 290 244 291 245
rect 289 244 290 245
rect 288 244 289 245
rect 287 244 288 245
rect 286 244 287 245
rect 285 244 286 245
rect 284 244 285 245
rect 283 244 284 245
rect 282 244 283 245
rect 281 244 282 245
rect 280 244 281 245
rect 279 244 280 245
rect 278 244 279 245
rect 277 244 278 245
rect 276 244 277 245
rect 275 244 276 245
rect 274 244 275 245
rect 273 244 274 245
rect 272 244 273 245
rect 271 244 272 245
rect 265 244 266 245
rect 264 244 265 245
rect 263 244 264 245
rect 262 244 263 245
rect 261 244 262 245
rect 260 244 261 245
rect 259 244 260 245
rect 258 244 259 245
rect 257 244 258 245
rect 256 244 257 245
rect 255 244 256 245
rect 254 244 255 245
rect 253 244 254 245
rect 252 244 253 245
rect 251 244 252 245
rect 250 244 251 245
rect 249 244 250 245
rect 248 244 249 245
rect 247 244 248 245
rect 246 244 247 245
rect 245 244 246 245
rect 244 244 245 245
rect 243 244 244 245
rect 242 244 243 245
rect 241 244 242 245
rect 240 244 241 245
rect 239 244 240 245
rect 238 244 239 245
rect 237 244 238 245
rect 236 244 237 245
rect 235 244 236 245
rect 234 244 235 245
rect 233 244 234 245
rect 232 244 233 245
rect 220 244 221 245
rect 219 244 220 245
rect 218 244 219 245
rect 217 244 218 245
rect 216 244 217 245
rect 215 244 216 245
rect 214 244 215 245
rect 213 244 214 245
rect 212 244 213 245
rect 211 244 212 245
rect 210 244 211 245
rect 209 244 210 245
rect 208 244 209 245
rect 207 244 208 245
rect 206 244 207 245
rect 205 244 206 245
rect 204 244 205 245
rect 203 244 204 245
rect 202 244 203 245
rect 201 244 202 245
rect 200 244 201 245
rect 199 244 200 245
rect 198 244 199 245
rect 197 244 198 245
rect 196 244 197 245
rect 195 244 196 245
rect 194 244 195 245
rect 193 244 194 245
rect 192 244 193 245
rect 191 244 192 245
rect 152 244 153 245
rect 151 244 152 245
rect 150 244 151 245
rect 149 244 150 245
rect 148 244 149 245
rect 147 244 148 245
rect 146 244 147 245
rect 145 244 146 245
rect 144 244 145 245
rect 143 244 144 245
rect 142 244 143 245
rect 141 244 142 245
rect 140 244 141 245
rect 139 244 140 245
rect 138 244 139 245
rect 137 244 138 245
rect 136 244 137 245
rect 135 244 136 245
rect 134 244 135 245
rect 133 244 134 245
rect 132 244 133 245
rect 131 244 132 245
rect 130 244 131 245
rect 129 244 130 245
rect 128 244 129 245
rect 127 244 128 245
rect 126 244 127 245
rect 125 244 126 245
rect 124 244 125 245
rect 123 244 124 245
rect 122 244 123 245
rect 121 244 122 245
rect 120 244 121 245
rect 119 244 120 245
rect 105 244 106 245
rect 104 244 105 245
rect 103 244 104 245
rect 102 244 103 245
rect 101 244 102 245
rect 100 244 101 245
rect 99 244 100 245
rect 98 244 99 245
rect 97 244 98 245
rect 96 244 97 245
rect 95 244 96 245
rect 94 244 95 245
rect 93 244 94 245
rect 92 244 93 245
rect 91 244 92 245
rect 90 244 91 245
rect 89 244 90 245
rect 88 244 89 245
rect 87 244 88 245
rect 86 244 87 245
rect 85 244 86 245
rect 84 244 85 245
rect 83 244 84 245
rect 82 244 83 245
rect 81 244 82 245
rect 80 244 81 245
rect 79 244 80 245
rect 78 244 79 245
rect 77 244 78 245
rect 76 244 77 245
rect 75 244 76 245
rect 74 244 75 245
rect 73 244 74 245
rect 72 244 73 245
rect 71 244 72 245
rect 70 244 71 245
rect 69 244 70 245
rect 68 244 69 245
rect 67 244 68 245
rect 66 244 67 245
rect 65 244 66 245
rect 64 244 65 245
rect 63 244 64 245
rect 62 244 63 245
rect 61 244 62 245
rect 60 244 61 245
rect 59 244 60 245
rect 58 244 59 245
rect 57 244 58 245
rect 56 244 57 245
rect 55 244 56 245
rect 54 244 55 245
rect 53 244 54 245
rect 52 244 53 245
rect 51 244 52 245
rect 50 244 51 245
rect 49 244 50 245
rect 48 244 49 245
rect 47 244 48 245
rect 46 244 47 245
rect 45 244 46 245
rect 44 244 45 245
rect 43 244 44 245
rect 42 244 43 245
rect 41 244 42 245
rect 40 244 41 245
rect 39 244 40 245
rect 38 244 39 245
rect 37 244 38 245
rect 36 244 37 245
rect 35 244 36 245
rect 34 244 35 245
rect 33 244 34 245
rect 32 244 33 245
rect 31 244 32 245
rect 30 244 31 245
rect 29 244 30 245
rect 21 244 22 245
rect 20 244 21 245
rect 19 244 20 245
rect 18 244 19 245
rect 17 244 18 245
rect 16 244 17 245
rect 15 244 16 245
rect 14 244 15 245
rect 13 244 14 245
rect 12 244 13 245
rect 11 244 12 245
rect 10 244 11 245
rect 9 244 10 245
rect 8 244 9 245
rect 7 244 8 245
rect 6 244 7 245
rect 5 244 6 245
rect 4 244 5 245
rect 3 244 4 245
rect 480 245 481 246
rect 479 245 480 246
rect 478 245 479 246
rect 477 245 478 246
rect 476 245 477 246
rect 468 245 469 246
rect 467 245 468 246
rect 466 245 467 246
rect 465 245 466 246
rect 464 245 465 246
rect 463 245 464 246
rect 462 245 463 246
rect 439 245 440 246
rect 438 245 439 246
rect 437 245 438 246
rect 436 245 437 246
rect 435 245 436 246
rect 434 245 435 246
rect 433 245 434 246
rect 432 245 433 246
rect 431 245 432 246
rect 430 245 431 246
rect 429 245 430 246
rect 428 245 429 246
rect 427 245 428 246
rect 426 245 427 246
rect 425 245 426 246
rect 424 245 425 246
rect 423 245 424 246
rect 422 245 423 246
rect 421 245 422 246
rect 420 245 421 246
rect 419 245 420 246
rect 418 245 419 246
rect 404 245 405 246
rect 403 245 404 246
rect 402 245 403 246
rect 401 245 402 246
rect 400 245 401 246
rect 399 245 400 246
rect 398 245 399 246
rect 397 245 398 246
rect 396 245 397 246
rect 395 245 396 246
rect 325 245 326 246
rect 324 245 325 246
rect 323 245 324 246
rect 322 245 323 246
rect 321 245 322 246
rect 320 245 321 246
rect 319 245 320 246
rect 318 245 319 246
rect 317 245 318 246
rect 316 245 317 246
rect 315 245 316 246
rect 314 245 315 246
rect 313 245 314 246
rect 312 245 313 246
rect 311 245 312 246
rect 310 245 311 246
rect 309 245 310 246
rect 308 245 309 246
rect 307 245 308 246
rect 306 245 307 246
rect 305 245 306 246
rect 304 245 305 246
rect 303 245 304 246
rect 302 245 303 246
rect 301 245 302 246
rect 300 245 301 246
rect 299 245 300 246
rect 298 245 299 246
rect 297 245 298 246
rect 296 245 297 246
rect 295 245 296 246
rect 294 245 295 246
rect 293 245 294 246
rect 292 245 293 246
rect 291 245 292 246
rect 290 245 291 246
rect 289 245 290 246
rect 288 245 289 246
rect 287 245 288 246
rect 286 245 287 246
rect 285 245 286 246
rect 284 245 285 246
rect 283 245 284 246
rect 282 245 283 246
rect 281 245 282 246
rect 280 245 281 246
rect 279 245 280 246
rect 278 245 279 246
rect 277 245 278 246
rect 276 245 277 246
rect 275 245 276 246
rect 274 245 275 246
rect 273 245 274 246
rect 272 245 273 246
rect 271 245 272 246
rect 270 245 271 246
rect 269 245 270 246
rect 265 245 266 246
rect 264 245 265 246
rect 263 245 264 246
rect 262 245 263 246
rect 261 245 262 246
rect 260 245 261 246
rect 259 245 260 246
rect 258 245 259 246
rect 257 245 258 246
rect 256 245 257 246
rect 255 245 256 246
rect 254 245 255 246
rect 253 245 254 246
rect 252 245 253 246
rect 251 245 252 246
rect 250 245 251 246
rect 249 245 250 246
rect 248 245 249 246
rect 247 245 248 246
rect 246 245 247 246
rect 245 245 246 246
rect 244 245 245 246
rect 243 245 244 246
rect 242 245 243 246
rect 241 245 242 246
rect 240 245 241 246
rect 239 245 240 246
rect 238 245 239 246
rect 237 245 238 246
rect 236 245 237 246
rect 235 245 236 246
rect 234 245 235 246
rect 233 245 234 246
rect 232 245 233 246
rect 214 245 215 246
rect 213 245 214 246
rect 212 245 213 246
rect 211 245 212 246
rect 210 245 211 246
rect 209 245 210 246
rect 208 245 209 246
rect 207 245 208 246
rect 206 245 207 246
rect 205 245 206 246
rect 204 245 205 246
rect 203 245 204 246
rect 202 245 203 246
rect 201 245 202 246
rect 200 245 201 246
rect 199 245 200 246
rect 198 245 199 246
rect 197 245 198 246
rect 196 245 197 246
rect 153 245 154 246
rect 152 245 153 246
rect 151 245 152 246
rect 150 245 151 246
rect 149 245 150 246
rect 148 245 149 246
rect 147 245 148 246
rect 146 245 147 246
rect 145 245 146 246
rect 144 245 145 246
rect 143 245 144 246
rect 142 245 143 246
rect 141 245 142 246
rect 140 245 141 246
rect 139 245 140 246
rect 138 245 139 246
rect 137 245 138 246
rect 136 245 137 246
rect 135 245 136 246
rect 134 245 135 246
rect 133 245 134 246
rect 132 245 133 246
rect 131 245 132 246
rect 130 245 131 246
rect 129 245 130 246
rect 128 245 129 246
rect 127 245 128 246
rect 126 245 127 246
rect 125 245 126 246
rect 124 245 125 246
rect 123 245 124 246
rect 122 245 123 246
rect 121 245 122 246
rect 120 245 121 246
rect 105 245 106 246
rect 104 245 105 246
rect 103 245 104 246
rect 102 245 103 246
rect 101 245 102 246
rect 100 245 101 246
rect 99 245 100 246
rect 98 245 99 246
rect 97 245 98 246
rect 96 245 97 246
rect 95 245 96 246
rect 94 245 95 246
rect 93 245 94 246
rect 92 245 93 246
rect 91 245 92 246
rect 90 245 91 246
rect 89 245 90 246
rect 88 245 89 246
rect 87 245 88 246
rect 86 245 87 246
rect 85 245 86 246
rect 84 245 85 246
rect 83 245 84 246
rect 82 245 83 246
rect 81 245 82 246
rect 80 245 81 246
rect 79 245 80 246
rect 78 245 79 246
rect 77 245 78 246
rect 76 245 77 246
rect 75 245 76 246
rect 74 245 75 246
rect 73 245 74 246
rect 72 245 73 246
rect 71 245 72 246
rect 70 245 71 246
rect 69 245 70 246
rect 68 245 69 246
rect 67 245 68 246
rect 66 245 67 246
rect 65 245 66 246
rect 64 245 65 246
rect 63 245 64 246
rect 62 245 63 246
rect 61 245 62 246
rect 60 245 61 246
rect 59 245 60 246
rect 58 245 59 246
rect 57 245 58 246
rect 56 245 57 246
rect 55 245 56 246
rect 54 245 55 246
rect 53 245 54 246
rect 52 245 53 246
rect 51 245 52 246
rect 50 245 51 246
rect 49 245 50 246
rect 48 245 49 246
rect 47 245 48 246
rect 46 245 47 246
rect 45 245 46 246
rect 44 245 45 246
rect 43 245 44 246
rect 42 245 43 246
rect 41 245 42 246
rect 40 245 41 246
rect 39 245 40 246
rect 38 245 39 246
rect 37 245 38 246
rect 36 245 37 246
rect 35 245 36 246
rect 34 245 35 246
rect 33 245 34 246
rect 32 245 33 246
rect 31 245 32 246
rect 30 245 31 246
rect 29 245 30 246
rect 21 245 22 246
rect 20 245 21 246
rect 19 245 20 246
rect 18 245 19 246
rect 17 245 18 246
rect 16 245 17 246
rect 15 245 16 246
rect 14 245 15 246
rect 13 245 14 246
rect 12 245 13 246
rect 11 245 12 246
rect 10 245 11 246
rect 9 245 10 246
rect 8 245 9 246
rect 7 245 8 246
rect 6 245 7 246
rect 5 245 6 246
rect 4 245 5 246
rect 3 245 4 246
rect 480 246 481 247
rect 479 246 480 247
rect 478 246 479 247
rect 477 246 478 247
rect 469 246 470 247
rect 468 246 469 247
rect 467 246 468 247
rect 466 246 467 247
rect 465 246 466 247
rect 464 246 465 247
rect 463 246 464 247
rect 462 246 463 247
rect 461 246 462 247
rect 438 246 439 247
rect 437 246 438 247
rect 436 246 437 247
rect 435 246 436 247
rect 434 246 435 247
rect 433 246 434 247
rect 432 246 433 247
rect 431 246 432 247
rect 430 246 431 247
rect 429 246 430 247
rect 428 246 429 247
rect 427 246 428 247
rect 426 246 427 247
rect 425 246 426 247
rect 424 246 425 247
rect 423 246 424 247
rect 422 246 423 247
rect 421 246 422 247
rect 420 246 421 247
rect 419 246 420 247
rect 418 246 419 247
rect 407 246 408 247
rect 406 246 407 247
rect 405 246 406 247
rect 404 246 405 247
rect 403 246 404 247
rect 402 246 403 247
rect 401 246 402 247
rect 400 246 401 247
rect 399 246 400 247
rect 398 246 399 247
rect 397 246 398 247
rect 396 246 397 247
rect 323 246 324 247
rect 322 246 323 247
rect 321 246 322 247
rect 320 246 321 247
rect 319 246 320 247
rect 318 246 319 247
rect 317 246 318 247
rect 316 246 317 247
rect 315 246 316 247
rect 314 246 315 247
rect 313 246 314 247
rect 312 246 313 247
rect 311 246 312 247
rect 310 246 311 247
rect 309 246 310 247
rect 308 246 309 247
rect 307 246 308 247
rect 306 246 307 247
rect 305 246 306 247
rect 304 246 305 247
rect 303 246 304 247
rect 302 246 303 247
rect 301 246 302 247
rect 300 246 301 247
rect 299 246 300 247
rect 298 246 299 247
rect 297 246 298 247
rect 296 246 297 247
rect 295 246 296 247
rect 294 246 295 247
rect 293 246 294 247
rect 292 246 293 247
rect 291 246 292 247
rect 290 246 291 247
rect 289 246 290 247
rect 288 246 289 247
rect 287 246 288 247
rect 286 246 287 247
rect 285 246 286 247
rect 284 246 285 247
rect 283 246 284 247
rect 282 246 283 247
rect 281 246 282 247
rect 280 246 281 247
rect 279 246 280 247
rect 278 246 279 247
rect 277 246 278 247
rect 276 246 277 247
rect 275 246 276 247
rect 274 246 275 247
rect 273 246 274 247
rect 272 246 273 247
rect 271 246 272 247
rect 270 246 271 247
rect 269 246 270 247
rect 268 246 269 247
rect 267 246 268 247
rect 264 246 265 247
rect 263 246 264 247
rect 262 246 263 247
rect 261 246 262 247
rect 260 246 261 247
rect 259 246 260 247
rect 258 246 259 247
rect 257 246 258 247
rect 256 246 257 247
rect 255 246 256 247
rect 254 246 255 247
rect 253 246 254 247
rect 252 246 253 247
rect 251 246 252 247
rect 250 246 251 247
rect 249 246 250 247
rect 248 246 249 247
rect 247 246 248 247
rect 246 246 247 247
rect 245 246 246 247
rect 244 246 245 247
rect 243 246 244 247
rect 242 246 243 247
rect 241 246 242 247
rect 240 246 241 247
rect 239 246 240 247
rect 238 246 239 247
rect 237 246 238 247
rect 236 246 237 247
rect 235 246 236 247
rect 234 246 235 247
rect 233 246 234 247
rect 232 246 233 247
rect 154 246 155 247
rect 153 246 154 247
rect 152 246 153 247
rect 151 246 152 247
rect 150 246 151 247
rect 149 246 150 247
rect 148 246 149 247
rect 147 246 148 247
rect 146 246 147 247
rect 145 246 146 247
rect 144 246 145 247
rect 143 246 144 247
rect 142 246 143 247
rect 141 246 142 247
rect 140 246 141 247
rect 139 246 140 247
rect 138 246 139 247
rect 137 246 138 247
rect 136 246 137 247
rect 135 246 136 247
rect 134 246 135 247
rect 133 246 134 247
rect 132 246 133 247
rect 131 246 132 247
rect 130 246 131 247
rect 129 246 130 247
rect 128 246 129 247
rect 127 246 128 247
rect 126 246 127 247
rect 125 246 126 247
rect 124 246 125 247
rect 123 246 124 247
rect 122 246 123 247
rect 121 246 122 247
rect 120 246 121 247
rect 106 246 107 247
rect 105 246 106 247
rect 104 246 105 247
rect 103 246 104 247
rect 102 246 103 247
rect 101 246 102 247
rect 100 246 101 247
rect 99 246 100 247
rect 98 246 99 247
rect 97 246 98 247
rect 96 246 97 247
rect 95 246 96 247
rect 94 246 95 247
rect 93 246 94 247
rect 92 246 93 247
rect 91 246 92 247
rect 90 246 91 247
rect 89 246 90 247
rect 88 246 89 247
rect 87 246 88 247
rect 86 246 87 247
rect 85 246 86 247
rect 84 246 85 247
rect 83 246 84 247
rect 82 246 83 247
rect 81 246 82 247
rect 80 246 81 247
rect 79 246 80 247
rect 78 246 79 247
rect 77 246 78 247
rect 76 246 77 247
rect 75 246 76 247
rect 74 246 75 247
rect 73 246 74 247
rect 72 246 73 247
rect 71 246 72 247
rect 70 246 71 247
rect 69 246 70 247
rect 68 246 69 247
rect 67 246 68 247
rect 66 246 67 247
rect 65 246 66 247
rect 64 246 65 247
rect 63 246 64 247
rect 62 246 63 247
rect 61 246 62 247
rect 60 246 61 247
rect 59 246 60 247
rect 58 246 59 247
rect 57 246 58 247
rect 56 246 57 247
rect 55 246 56 247
rect 54 246 55 247
rect 53 246 54 247
rect 52 246 53 247
rect 51 246 52 247
rect 50 246 51 247
rect 49 246 50 247
rect 48 246 49 247
rect 47 246 48 247
rect 46 246 47 247
rect 45 246 46 247
rect 44 246 45 247
rect 43 246 44 247
rect 42 246 43 247
rect 41 246 42 247
rect 40 246 41 247
rect 39 246 40 247
rect 38 246 39 247
rect 37 246 38 247
rect 36 246 37 247
rect 35 246 36 247
rect 34 246 35 247
rect 33 246 34 247
rect 32 246 33 247
rect 31 246 32 247
rect 30 246 31 247
rect 21 246 22 247
rect 20 246 21 247
rect 19 246 20 247
rect 18 246 19 247
rect 17 246 18 247
rect 16 246 17 247
rect 15 246 16 247
rect 14 246 15 247
rect 13 246 14 247
rect 12 246 13 247
rect 11 246 12 247
rect 10 246 11 247
rect 9 246 10 247
rect 8 246 9 247
rect 7 246 8 247
rect 6 246 7 247
rect 5 246 6 247
rect 4 246 5 247
rect 3 246 4 247
rect 481 247 482 248
rect 480 247 481 248
rect 479 247 480 248
rect 470 247 471 248
rect 469 247 470 248
rect 468 247 469 248
rect 467 247 468 248
rect 466 247 467 248
rect 465 247 466 248
rect 464 247 465 248
rect 463 247 464 248
rect 462 247 463 248
rect 461 247 462 248
rect 460 247 461 248
rect 438 247 439 248
rect 437 247 438 248
rect 436 247 437 248
rect 435 247 436 248
rect 434 247 435 248
rect 433 247 434 248
rect 432 247 433 248
rect 431 247 432 248
rect 430 247 431 248
rect 429 247 430 248
rect 428 247 429 248
rect 427 247 428 248
rect 426 247 427 248
rect 425 247 426 248
rect 424 247 425 248
rect 423 247 424 248
rect 422 247 423 248
rect 421 247 422 248
rect 420 247 421 248
rect 419 247 420 248
rect 418 247 419 248
rect 407 247 408 248
rect 406 247 407 248
rect 405 247 406 248
rect 404 247 405 248
rect 403 247 404 248
rect 402 247 403 248
rect 401 247 402 248
rect 400 247 401 248
rect 399 247 400 248
rect 398 247 399 248
rect 397 247 398 248
rect 396 247 397 248
rect 321 247 322 248
rect 320 247 321 248
rect 319 247 320 248
rect 318 247 319 248
rect 317 247 318 248
rect 316 247 317 248
rect 315 247 316 248
rect 314 247 315 248
rect 313 247 314 248
rect 312 247 313 248
rect 311 247 312 248
rect 310 247 311 248
rect 309 247 310 248
rect 308 247 309 248
rect 307 247 308 248
rect 306 247 307 248
rect 305 247 306 248
rect 304 247 305 248
rect 303 247 304 248
rect 302 247 303 248
rect 301 247 302 248
rect 300 247 301 248
rect 299 247 300 248
rect 298 247 299 248
rect 297 247 298 248
rect 296 247 297 248
rect 295 247 296 248
rect 294 247 295 248
rect 293 247 294 248
rect 292 247 293 248
rect 291 247 292 248
rect 290 247 291 248
rect 289 247 290 248
rect 288 247 289 248
rect 287 247 288 248
rect 286 247 287 248
rect 285 247 286 248
rect 284 247 285 248
rect 283 247 284 248
rect 282 247 283 248
rect 281 247 282 248
rect 280 247 281 248
rect 279 247 280 248
rect 278 247 279 248
rect 277 247 278 248
rect 276 247 277 248
rect 275 247 276 248
rect 274 247 275 248
rect 273 247 274 248
rect 272 247 273 248
rect 271 247 272 248
rect 270 247 271 248
rect 269 247 270 248
rect 268 247 269 248
rect 267 247 268 248
rect 266 247 267 248
rect 265 247 266 248
rect 263 247 264 248
rect 262 247 263 248
rect 261 247 262 248
rect 260 247 261 248
rect 259 247 260 248
rect 258 247 259 248
rect 257 247 258 248
rect 256 247 257 248
rect 255 247 256 248
rect 254 247 255 248
rect 253 247 254 248
rect 252 247 253 248
rect 251 247 252 248
rect 250 247 251 248
rect 249 247 250 248
rect 248 247 249 248
rect 247 247 248 248
rect 246 247 247 248
rect 245 247 246 248
rect 244 247 245 248
rect 243 247 244 248
rect 242 247 243 248
rect 241 247 242 248
rect 240 247 241 248
rect 239 247 240 248
rect 238 247 239 248
rect 237 247 238 248
rect 236 247 237 248
rect 235 247 236 248
rect 234 247 235 248
rect 233 247 234 248
rect 232 247 233 248
rect 155 247 156 248
rect 154 247 155 248
rect 153 247 154 248
rect 152 247 153 248
rect 151 247 152 248
rect 150 247 151 248
rect 149 247 150 248
rect 148 247 149 248
rect 147 247 148 248
rect 146 247 147 248
rect 145 247 146 248
rect 144 247 145 248
rect 143 247 144 248
rect 142 247 143 248
rect 141 247 142 248
rect 140 247 141 248
rect 139 247 140 248
rect 138 247 139 248
rect 137 247 138 248
rect 136 247 137 248
rect 135 247 136 248
rect 134 247 135 248
rect 133 247 134 248
rect 132 247 133 248
rect 131 247 132 248
rect 130 247 131 248
rect 129 247 130 248
rect 128 247 129 248
rect 127 247 128 248
rect 126 247 127 248
rect 125 247 126 248
rect 124 247 125 248
rect 123 247 124 248
rect 122 247 123 248
rect 121 247 122 248
rect 120 247 121 248
rect 106 247 107 248
rect 105 247 106 248
rect 104 247 105 248
rect 103 247 104 248
rect 102 247 103 248
rect 101 247 102 248
rect 100 247 101 248
rect 99 247 100 248
rect 98 247 99 248
rect 97 247 98 248
rect 96 247 97 248
rect 95 247 96 248
rect 94 247 95 248
rect 93 247 94 248
rect 92 247 93 248
rect 91 247 92 248
rect 90 247 91 248
rect 89 247 90 248
rect 88 247 89 248
rect 87 247 88 248
rect 86 247 87 248
rect 85 247 86 248
rect 84 247 85 248
rect 83 247 84 248
rect 82 247 83 248
rect 81 247 82 248
rect 80 247 81 248
rect 79 247 80 248
rect 78 247 79 248
rect 77 247 78 248
rect 76 247 77 248
rect 75 247 76 248
rect 74 247 75 248
rect 73 247 74 248
rect 72 247 73 248
rect 71 247 72 248
rect 70 247 71 248
rect 69 247 70 248
rect 68 247 69 248
rect 67 247 68 248
rect 66 247 67 248
rect 65 247 66 248
rect 64 247 65 248
rect 63 247 64 248
rect 62 247 63 248
rect 61 247 62 248
rect 60 247 61 248
rect 59 247 60 248
rect 58 247 59 248
rect 57 247 58 248
rect 56 247 57 248
rect 55 247 56 248
rect 54 247 55 248
rect 53 247 54 248
rect 52 247 53 248
rect 51 247 52 248
rect 50 247 51 248
rect 49 247 50 248
rect 48 247 49 248
rect 47 247 48 248
rect 46 247 47 248
rect 45 247 46 248
rect 44 247 45 248
rect 43 247 44 248
rect 42 247 43 248
rect 41 247 42 248
rect 40 247 41 248
rect 39 247 40 248
rect 38 247 39 248
rect 37 247 38 248
rect 36 247 37 248
rect 35 247 36 248
rect 34 247 35 248
rect 33 247 34 248
rect 32 247 33 248
rect 31 247 32 248
rect 30 247 31 248
rect 21 247 22 248
rect 20 247 21 248
rect 19 247 20 248
rect 18 247 19 248
rect 17 247 18 248
rect 16 247 17 248
rect 15 247 16 248
rect 14 247 15 248
rect 13 247 14 248
rect 12 247 13 248
rect 11 247 12 248
rect 10 247 11 248
rect 9 247 10 248
rect 8 247 9 248
rect 7 247 8 248
rect 6 247 7 248
rect 5 247 6 248
rect 4 247 5 248
rect 3 247 4 248
rect 481 248 482 249
rect 480 248 481 249
rect 471 248 472 249
rect 470 248 471 249
rect 469 248 470 249
rect 468 248 469 249
rect 467 248 468 249
rect 466 248 467 249
rect 465 248 466 249
rect 462 248 463 249
rect 461 248 462 249
rect 460 248 461 249
rect 438 248 439 249
rect 437 248 438 249
rect 436 248 437 249
rect 435 248 436 249
rect 434 248 435 249
rect 433 248 434 249
rect 432 248 433 249
rect 431 248 432 249
rect 430 248 431 249
rect 429 248 430 249
rect 428 248 429 249
rect 427 248 428 249
rect 426 248 427 249
rect 425 248 426 249
rect 424 248 425 249
rect 423 248 424 249
rect 422 248 423 249
rect 421 248 422 249
rect 420 248 421 249
rect 419 248 420 249
rect 418 248 419 249
rect 407 248 408 249
rect 406 248 407 249
rect 405 248 406 249
rect 404 248 405 249
rect 403 248 404 249
rect 402 248 403 249
rect 401 248 402 249
rect 400 248 401 249
rect 399 248 400 249
rect 319 248 320 249
rect 318 248 319 249
rect 317 248 318 249
rect 316 248 317 249
rect 315 248 316 249
rect 314 248 315 249
rect 313 248 314 249
rect 312 248 313 249
rect 311 248 312 249
rect 310 248 311 249
rect 309 248 310 249
rect 308 248 309 249
rect 307 248 308 249
rect 306 248 307 249
rect 305 248 306 249
rect 304 248 305 249
rect 303 248 304 249
rect 302 248 303 249
rect 301 248 302 249
rect 300 248 301 249
rect 299 248 300 249
rect 298 248 299 249
rect 297 248 298 249
rect 296 248 297 249
rect 295 248 296 249
rect 294 248 295 249
rect 293 248 294 249
rect 292 248 293 249
rect 291 248 292 249
rect 290 248 291 249
rect 289 248 290 249
rect 288 248 289 249
rect 287 248 288 249
rect 286 248 287 249
rect 285 248 286 249
rect 284 248 285 249
rect 283 248 284 249
rect 282 248 283 249
rect 281 248 282 249
rect 280 248 281 249
rect 279 248 280 249
rect 278 248 279 249
rect 277 248 278 249
rect 276 248 277 249
rect 275 248 276 249
rect 274 248 275 249
rect 273 248 274 249
rect 272 248 273 249
rect 271 248 272 249
rect 270 248 271 249
rect 269 248 270 249
rect 268 248 269 249
rect 267 248 268 249
rect 266 248 267 249
rect 265 248 266 249
rect 264 248 265 249
rect 263 248 264 249
rect 262 248 263 249
rect 261 248 262 249
rect 260 248 261 249
rect 259 248 260 249
rect 258 248 259 249
rect 257 248 258 249
rect 256 248 257 249
rect 255 248 256 249
rect 254 248 255 249
rect 253 248 254 249
rect 252 248 253 249
rect 251 248 252 249
rect 250 248 251 249
rect 249 248 250 249
rect 248 248 249 249
rect 247 248 248 249
rect 246 248 247 249
rect 245 248 246 249
rect 244 248 245 249
rect 243 248 244 249
rect 242 248 243 249
rect 241 248 242 249
rect 240 248 241 249
rect 239 248 240 249
rect 238 248 239 249
rect 237 248 238 249
rect 236 248 237 249
rect 235 248 236 249
rect 234 248 235 249
rect 233 248 234 249
rect 232 248 233 249
rect 156 248 157 249
rect 155 248 156 249
rect 154 248 155 249
rect 153 248 154 249
rect 152 248 153 249
rect 151 248 152 249
rect 150 248 151 249
rect 149 248 150 249
rect 148 248 149 249
rect 147 248 148 249
rect 146 248 147 249
rect 145 248 146 249
rect 144 248 145 249
rect 143 248 144 249
rect 142 248 143 249
rect 141 248 142 249
rect 140 248 141 249
rect 139 248 140 249
rect 138 248 139 249
rect 137 248 138 249
rect 136 248 137 249
rect 135 248 136 249
rect 134 248 135 249
rect 133 248 134 249
rect 132 248 133 249
rect 131 248 132 249
rect 130 248 131 249
rect 129 248 130 249
rect 128 248 129 249
rect 127 248 128 249
rect 126 248 127 249
rect 125 248 126 249
rect 124 248 125 249
rect 123 248 124 249
rect 122 248 123 249
rect 121 248 122 249
rect 120 248 121 249
rect 107 248 108 249
rect 106 248 107 249
rect 105 248 106 249
rect 104 248 105 249
rect 103 248 104 249
rect 102 248 103 249
rect 101 248 102 249
rect 100 248 101 249
rect 99 248 100 249
rect 98 248 99 249
rect 97 248 98 249
rect 96 248 97 249
rect 95 248 96 249
rect 94 248 95 249
rect 93 248 94 249
rect 92 248 93 249
rect 91 248 92 249
rect 90 248 91 249
rect 89 248 90 249
rect 88 248 89 249
rect 87 248 88 249
rect 86 248 87 249
rect 85 248 86 249
rect 84 248 85 249
rect 83 248 84 249
rect 82 248 83 249
rect 81 248 82 249
rect 80 248 81 249
rect 79 248 80 249
rect 78 248 79 249
rect 77 248 78 249
rect 76 248 77 249
rect 75 248 76 249
rect 74 248 75 249
rect 73 248 74 249
rect 72 248 73 249
rect 71 248 72 249
rect 70 248 71 249
rect 69 248 70 249
rect 68 248 69 249
rect 67 248 68 249
rect 66 248 67 249
rect 65 248 66 249
rect 64 248 65 249
rect 63 248 64 249
rect 62 248 63 249
rect 61 248 62 249
rect 60 248 61 249
rect 59 248 60 249
rect 58 248 59 249
rect 57 248 58 249
rect 56 248 57 249
rect 55 248 56 249
rect 54 248 55 249
rect 53 248 54 249
rect 52 248 53 249
rect 51 248 52 249
rect 50 248 51 249
rect 49 248 50 249
rect 48 248 49 249
rect 47 248 48 249
rect 46 248 47 249
rect 45 248 46 249
rect 44 248 45 249
rect 43 248 44 249
rect 42 248 43 249
rect 41 248 42 249
rect 40 248 41 249
rect 39 248 40 249
rect 38 248 39 249
rect 37 248 38 249
rect 36 248 37 249
rect 35 248 36 249
rect 34 248 35 249
rect 33 248 34 249
rect 32 248 33 249
rect 31 248 32 249
rect 30 248 31 249
rect 21 248 22 249
rect 20 248 21 249
rect 19 248 20 249
rect 18 248 19 249
rect 17 248 18 249
rect 16 248 17 249
rect 15 248 16 249
rect 14 248 15 249
rect 13 248 14 249
rect 12 248 13 249
rect 11 248 12 249
rect 10 248 11 249
rect 9 248 10 249
rect 8 248 9 249
rect 7 248 8 249
rect 6 248 7 249
rect 5 248 6 249
rect 4 248 5 249
rect 3 248 4 249
rect 481 249 482 250
rect 480 249 481 250
rect 471 249 472 250
rect 470 249 471 250
rect 469 249 470 250
rect 468 249 469 250
rect 467 249 468 250
rect 466 249 467 250
rect 460 249 461 250
rect 459 249 460 250
rect 422 249 423 250
rect 421 249 422 250
rect 420 249 421 250
rect 419 249 420 250
rect 418 249 419 250
rect 318 249 319 250
rect 317 249 318 250
rect 316 249 317 250
rect 315 249 316 250
rect 314 249 315 250
rect 313 249 314 250
rect 312 249 313 250
rect 311 249 312 250
rect 310 249 311 250
rect 309 249 310 250
rect 308 249 309 250
rect 307 249 308 250
rect 306 249 307 250
rect 305 249 306 250
rect 304 249 305 250
rect 303 249 304 250
rect 302 249 303 250
rect 301 249 302 250
rect 300 249 301 250
rect 299 249 300 250
rect 298 249 299 250
rect 297 249 298 250
rect 296 249 297 250
rect 295 249 296 250
rect 294 249 295 250
rect 293 249 294 250
rect 292 249 293 250
rect 291 249 292 250
rect 290 249 291 250
rect 289 249 290 250
rect 288 249 289 250
rect 287 249 288 250
rect 286 249 287 250
rect 285 249 286 250
rect 284 249 285 250
rect 283 249 284 250
rect 282 249 283 250
rect 281 249 282 250
rect 280 249 281 250
rect 279 249 280 250
rect 278 249 279 250
rect 277 249 278 250
rect 276 249 277 250
rect 275 249 276 250
rect 274 249 275 250
rect 273 249 274 250
rect 272 249 273 250
rect 271 249 272 250
rect 270 249 271 250
rect 269 249 270 250
rect 268 249 269 250
rect 267 249 268 250
rect 266 249 267 250
rect 265 249 266 250
rect 264 249 265 250
rect 263 249 264 250
rect 262 249 263 250
rect 261 249 262 250
rect 260 249 261 250
rect 259 249 260 250
rect 258 249 259 250
rect 257 249 258 250
rect 256 249 257 250
rect 255 249 256 250
rect 254 249 255 250
rect 253 249 254 250
rect 252 249 253 250
rect 251 249 252 250
rect 250 249 251 250
rect 249 249 250 250
rect 248 249 249 250
rect 247 249 248 250
rect 246 249 247 250
rect 245 249 246 250
rect 244 249 245 250
rect 243 249 244 250
rect 242 249 243 250
rect 241 249 242 250
rect 240 249 241 250
rect 239 249 240 250
rect 238 249 239 250
rect 237 249 238 250
rect 236 249 237 250
rect 235 249 236 250
rect 234 249 235 250
rect 233 249 234 250
rect 232 249 233 250
rect 231 249 232 250
rect 157 249 158 250
rect 156 249 157 250
rect 155 249 156 250
rect 154 249 155 250
rect 153 249 154 250
rect 152 249 153 250
rect 151 249 152 250
rect 150 249 151 250
rect 149 249 150 250
rect 148 249 149 250
rect 147 249 148 250
rect 146 249 147 250
rect 145 249 146 250
rect 144 249 145 250
rect 143 249 144 250
rect 142 249 143 250
rect 141 249 142 250
rect 140 249 141 250
rect 139 249 140 250
rect 138 249 139 250
rect 137 249 138 250
rect 136 249 137 250
rect 135 249 136 250
rect 134 249 135 250
rect 133 249 134 250
rect 132 249 133 250
rect 131 249 132 250
rect 130 249 131 250
rect 129 249 130 250
rect 128 249 129 250
rect 127 249 128 250
rect 126 249 127 250
rect 125 249 126 250
rect 124 249 125 250
rect 123 249 124 250
rect 122 249 123 250
rect 121 249 122 250
rect 120 249 121 250
rect 107 249 108 250
rect 106 249 107 250
rect 105 249 106 250
rect 104 249 105 250
rect 103 249 104 250
rect 102 249 103 250
rect 101 249 102 250
rect 100 249 101 250
rect 99 249 100 250
rect 98 249 99 250
rect 97 249 98 250
rect 96 249 97 250
rect 95 249 96 250
rect 94 249 95 250
rect 93 249 94 250
rect 92 249 93 250
rect 91 249 92 250
rect 90 249 91 250
rect 89 249 90 250
rect 88 249 89 250
rect 87 249 88 250
rect 86 249 87 250
rect 85 249 86 250
rect 84 249 85 250
rect 83 249 84 250
rect 82 249 83 250
rect 81 249 82 250
rect 80 249 81 250
rect 79 249 80 250
rect 78 249 79 250
rect 77 249 78 250
rect 76 249 77 250
rect 75 249 76 250
rect 74 249 75 250
rect 73 249 74 250
rect 72 249 73 250
rect 71 249 72 250
rect 70 249 71 250
rect 69 249 70 250
rect 68 249 69 250
rect 67 249 68 250
rect 66 249 67 250
rect 65 249 66 250
rect 64 249 65 250
rect 63 249 64 250
rect 62 249 63 250
rect 61 249 62 250
rect 60 249 61 250
rect 59 249 60 250
rect 58 249 59 250
rect 57 249 58 250
rect 56 249 57 250
rect 55 249 56 250
rect 54 249 55 250
rect 53 249 54 250
rect 52 249 53 250
rect 51 249 52 250
rect 50 249 51 250
rect 49 249 50 250
rect 48 249 49 250
rect 47 249 48 250
rect 46 249 47 250
rect 45 249 46 250
rect 44 249 45 250
rect 43 249 44 250
rect 42 249 43 250
rect 41 249 42 250
rect 40 249 41 250
rect 39 249 40 250
rect 38 249 39 250
rect 37 249 38 250
rect 36 249 37 250
rect 35 249 36 250
rect 34 249 35 250
rect 33 249 34 250
rect 32 249 33 250
rect 31 249 32 250
rect 21 249 22 250
rect 20 249 21 250
rect 19 249 20 250
rect 18 249 19 250
rect 17 249 18 250
rect 16 249 17 250
rect 15 249 16 250
rect 14 249 15 250
rect 13 249 14 250
rect 12 249 13 250
rect 11 249 12 250
rect 10 249 11 250
rect 9 249 10 250
rect 8 249 9 250
rect 7 249 8 250
rect 6 249 7 250
rect 5 249 6 250
rect 4 249 5 250
rect 3 249 4 250
rect 481 250 482 251
rect 480 250 481 251
rect 472 250 473 251
rect 471 250 472 251
rect 470 250 471 251
rect 469 250 470 251
rect 468 250 469 251
rect 467 250 468 251
rect 460 250 461 251
rect 459 250 460 251
rect 421 250 422 251
rect 420 250 421 251
rect 419 250 420 251
rect 418 250 419 251
rect 316 250 317 251
rect 315 250 316 251
rect 314 250 315 251
rect 313 250 314 251
rect 312 250 313 251
rect 311 250 312 251
rect 310 250 311 251
rect 309 250 310 251
rect 308 250 309 251
rect 307 250 308 251
rect 306 250 307 251
rect 305 250 306 251
rect 304 250 305 251
rect 303 250 304 251
rect 302 250 303 251
rect 301 250 302 251
rect 300 250 301 251
rect 299 250 300 251
rect 298 250 299 251
rect 297 250 298 251
rect 296 250 297 251
rect 295 250 296 251
rect 294 250 295 251
rect 293 250 294 251
rect 292 250 293 251
rect 291 250 292 251
rect 290 250 291 251
rect 289 250 290 251
rect 288 250 289 251
rect 287 250 288 251
rect 286 250 287 251
rect 285 250 286 251
rect 284 250 285 251
rect 283 250 284 251
rect 282 250 283 251
rect 281 250 282 251
rect 280 250 281 251
rect 279 250 280 251
rect 278 250 279 251
rect 277 250 278 251
rect 276 250 277 251
rect 275 250 276 251
rect 274 250 275 251
rect 273 250 274 251
rect 272 250 273 251
rect 271 250 272 251
rect 270 250 271 251
rect 269 250 270 251
rect 268 250 269 251
rect 267 250 268 251
rect 266 250 267 251
rect 265 250 266 251
rect 264 250 265 251
rect 263 250 264 251
rect 262 250 263 251
rect 261 250 262 251
rect 260 250 261 251
rect 259 250 260 251
rect 258 250 259 251
rect 257 250 258 251
rect 256 250 257 251
rect 255 250 256 251
rect 254 250 255 251
rect 253 250 254 251
rect 252 250 253 251
rect 251 250 252 251
rect 250 250 251 251
rect 249 250 250 251
rect 248 250 249 251
rect 247 250 248 251
rect 246 250 247 251
rect 245 250 246 251
rect 244 250 245 251
rect 243 250 244 251
rect 242 250 243 251
rect 241 250 242 251
rect 240 250 241 251
rect 239 250 240 251
rect 238 250 239 251
rect 237 250 238 251
rect 236 250 237 251
rect 235 250 236 251
rect 234 250 235 251
rect 233 250 234 251
rect 232 250 233 251
rect 231 250 232 251
rect 158 250 159 251
rect 157 250 158 251
rect 156 250 157 251
rect 155 250 156 251
rect 154 250 155 251
rect 153 250 154 251
rect 152 250 153 251
rect 151 250 152 251
rect 150 250 151 251
rect 149 250 150 251
rect 148 250 149 251
rect 147 250 148 251
rect 146 250 147 251
rect 145 250 146 251
rect 144 250 145 251
rect 143 250 144 251
rect 142 250 143 251
rect 141 250 142 251
rect 140 250 141 251
rect 139 250 140 251
rect 138 250 139 251
rect 137 250 138 251
rect 136 250 137 251
rect 135 250 136 251
rect 134 250 135 251
rect 133 250 134 251
rect 132 250 133 251
rect 131 250 132 251
rect 130 250 131 251
rect 129 250 130 251
rect 128 250 129 251
rect 127 250 128 251
rect 126 250 127 251
rect 125 250 126 251
rect 124 250 125 251
rect 123 250 124 251
rect 122 250 123 251
rect 121 250 122 251
rect 108 250 109 251
rect 107 250 108 251
rect 106 250 107 251
rect 105 250 106 251
rect 104 250 105 251
rect 103 250 104 251
rect 102 250 103 251
rect 101 250 102 251
rect 100 250 101 251
rect 99 250 100 251
rect 98 250 99 251
rect 97 250 98 251
rect 96 250 97 251
rect 95 250 96 251
rect 94 250 95 251
rect 93 250 94 251
rect 92 250 93 251
rect 91 250 92 251
rect 90 250 91 251
rect 89 250 90 251
rect 88 250 89 251
rect 87 250 88 251
rect 86 250 87 251
rect 85 250 86 251
rect 84 250 85 251
rect 83 250 84 251
rect 82 250 83 251
rect 81 250 82 251
rect 80 250 81 251
rect 79 250 80 251
rect 78 250 79 251
rect 77 250 78 251
rect 76 250 77 251
rect 75 250 76 251
rect 74 250 75 251
rect 73 250 74 251
rect 72 250 73 251
rect 71 250 72 251
rect 70 250 71 251
rect 69 250 70 251
rect 68 250 69 251
rect 67 250 68 251
rect 66 250 67 251
rect 65 250 66 251
rect 64 250 65 251
rect 63 250 64 251
rect 62 250 63 251
rect 61 250 62 251
rect 60 250 61 251
rect 59 250 60 251
rect 58 250 59 251
rect 57 250 58 251
rect 56 250 57 251
rect 55 250 56 251
rect 54 250 55 251
rect 53 250 54 251
rect 52 250 53 251
rect 51 250 52 251
rect 50 250 51 251
rect 49 250 50 251
rect 48 250 49 251
rect 47 250 48 251
rect 46 250 47 251
rect 45 250 46 251
rect 44 250 45 251
rect 43 250 44 251
rect 42 250 43 251
rect 41 250 42 251
rect 40 250 41 251
rect 39 250 40 251
rect 38 250 39 251
rect 37 250 38 251
rect 36 250 37 251
rect 35 250 36 251
rect 34 250 35 251
rect 33 250 34 251
rect 32 250 33 251
rect 31 250 32 251
rect 21 250 22 251
rect 20 250 21 251
rect 19 250 20 251
rect 18 250 19 251
rect 17 250 18 251
rect 16 250 17 251
rect 15 250 16 251
rect 14 250 15 251
rect 13 250 14 251
rect 12 250 13 251
rect 11 250 12 251
rect 10 250 11 251
rect 9 250 10 251
rect 8 250 9 251
rect 7 250 8 251
rect 6 250 7 251
rect 5 250 6 251
rect 4 250 5 251
rect 3 250 4 251
rect 481 251 482 252
rect 480 251 481 252
rect 472 251 473 252
rect 471 251 472 252
rect 470 251 471 252
rect 469 251 470 252
rect 468 251 469 252
rect 460 251 461 252
rect 459 251 460 252
rect 420 251 421 252
rect 419 251 420 252
rect 418 251 419 252
rect 315 251 316 252
rect 314 251 315 252
rect 313 251 314 252
rect 312 251 313 252
rect 311 251 312 252
rect 310 251 311 252
rect 309 251 310 252
rect 308 251 309 252
rect 307 251 308 252
rect 306 251 307 252
rect 305 251 306 252
rect 304 251 305 252
rect 303 251 304 252
rect 302 251 303 252
rect 301 251 302 252
rect 300 251 301 252
rect 299 251 300 252
rect 298 251 299 252
rect 297 251 298 252
rect 296 251 297 252
rect 295 251 296 252
rect 294 251 295 252
rect 293 251 294 252
rect 292 251 293 252
rect 291 251 292 252
rect 290 251 291 252
rect 289 251 290 252
rect 288 251 289 252
rect 287 251 288 252
rect 286 251 287 252
rect 285 251 286 252
rect 284 251 285 252
rect 283 251 284 252
rect 282 251 283 252
rect 281 251 282 252
rect 280 251 281 252
rect 279 251 280 252
rect 278 251 279 252
rect 277 251 278 252
rect 276 251 277 252
rect 275 251 276 252
rect 274 251 275 252
rect 273 251 274 252
rect 272 251 273 252
rect 271 251 272 252
rect 270 251 271 252
rect 269 251 270 252
rect 268 251 269 252
rect 267 251 268 252
rect 266 251 267 252
rect 265 251 266 252
rect 264 251 265 252
rect 263 251 264 252
rect 262 251 263 252
rect 261 251 262 252
rect 260 251 261 252
rect 259 251 260 252
rect 258 251 259 252
rect 257 251 258 252
rect 256 251 257 252
rect 255 251 256 252
rect 254 251 255 252
rect 253 251 254 252
rect 252 251 253 252
rect 251 251 252 252
rect 250 251 251 252
rect 249 251 250 252
rect 248 251 249 252
rect 247 251 248 252
rect 246 251 247 252
rect 245 251 246 252
rect 244 251 245 252
rect 243 251 244 252
rect 242 251 243 252
rect 241 251 242 252
rect 240 251 241 252
rect 239 251 240 252
rect 238 251 239 252
rect 237 251 238 252
rect 236 251 237 252
rect 235 251 236 252
rect 234 251 235 252
rect 233 251 234 252
rect 232 251 233 252
rect 231 251 232 252
rect 159 251 160 252
rect 158 251 159 252
rect 157 251 158 252
rect 156 251 157 252
rect 155 251 156 252
rect 154 251 155 252
rect 153 251 154 252
rect 152 251 153 252
rect 151 251 152 252
rect 150 251 151 252
rect 149 251 150 252
rect 148 251 149 252
rect 147 251 148 252
rect 146 251 147 252
rect 145 251 146 252
rect 144 251 145 252
rect 143 251 144 252
rect 142 251 143 252
rect 141 251 142 252
rect 140 251 141 252
rect 139 251 140 252
rect 138 251 139 252
rect 137 251 138 252
rect 136 251 137 252
rect 135 251 136 252
rect 134 251 135 252
rect 133 251 134 252
rect 132 251 133 252
rect 131 251 132 252
rect 130 251 131 252
rect 129 251 130 252
rect 128 251 129 252
rect 127 251 128 252
rect 126 251 127 252
rect 125 251 126 252
rect 124 251 125 252
rect 123 251 124 252
rect 122 251 123 252
rect 121 251 122 252
rect 108 251 109 252
rect 107 251 108 252
rect 106 251 107 252
rect 105 251 106 252
rect 104 251 105 252
rect 103 251 104 252
rect 102 251 103 252
rect 101 251 102 252
rect 100 251 101 252
rect 99 251 100 252
rect 98 251 99 252
rect 97 251 98 252
rect 96 251 97 252
rect 95 251 96 252
rect 94 251 95 252
rect 93 251 94 252
rect 92 251 93 252
rect 91 251 92 252
rect 90 251 91 252
rect 89 251 90 252
rect 88 251 89 252
rect 87 251 88 252
rect 86 251 87 252
rect 85 251 86 252
rect 84 251 85 252
rect 83 251 84 252
rect 82 251 83 252
rect 81 251 82 252
rect 80 251 81 252
rect 79 251 80 252
rect 78 251 79 252
rect 77 251 78 252
rect 76 251 77 252
rect 75 251 76 252
rect 74 251 75 252
rect 73 251 74 252
rect 72 251 73 252
rect 71 251 72 252
rect 70 251 71 252
rect 69 251 70 252
rect 68 251 69 252
rect 67 251 68 252
rect 66 251 67 252
rect 65 251 66 252
rect 64 251 65 252
rect 63 251 64 252
rect 62 251 63 252
rect 61 251 62 252
rect 60 251 61 252
rect 59 251 60 252
rect 58 251 59 252
rect 57 251 58 252
rect 56 251 57 252
rect 55 251 56 252
rect 54 251 55 252
rect 53 251 54 252
rect 52 251 53 252
rect 51 251 52 252
rect 50 251 51 252
rect 49 251 50 252
rect 48 251 49 252
rect 47 251 48 252
rect 46 251 47 252
rect 45 251 46 252
rect 44 251 45 252
rect 43 251 44 252
rect 42 251 43 252
rect 41 251 42 252
rect 40 251 41 252
rect 39 251 40 252
rect 38 251 39 252
rect 37 251 38 252
rect 36 251 37 252
rect 35 251 36 252
rect 34 251 35 252
rect 33 251 34 252
rect 32 251 33 252
rect 31 251 32 252
rect 21 251 22 252
rect 20 251 21 252
rect 19 251 20 252
rect 18 251 19 252
rect 17 251 18 252
rect 16 251 17 252
rect 15 251 16 252
rect 14 251 15 252
rect 13 251 14 252
rect 12 251 13 252
rect 11 251 12 252
rect 10 251 11 252
rect 9 251 10 252
rect 8 251 9 252
rect 7 251 8 252
rect 6 251 7 252
rect 5 251 6 252
rect 4 251 5 252
rect 3 251 4 252
rect 481 252 482 253
rect 480 252 481 253
rect 473 252 474 253
rect 472 252 473 253
rect 471 252 472 253
rect 470 252 471 253
rect 469 252 470 253
rect 468 252 469 253
rect 460 252 461 253
rect 459 252 460 253
rect 420 252 421 253
rect 419 252 420 253
rect 313 252 314 253
rect 312 252 313 253
rect 311 252 312 253
rect 310 252 311 253
rect 309 252 310 253
rect 308 252 309 253
rect 307 252 308 253
rect 306 252 307 253
rect 305 252 306 253
rect 304 252 305 253
rect 303 252 304 253
rect 302 252 303 253
rect 301 252 302 253
rect 300 252 301 253
rect 299 252 300 253
rect 298 252 299 253
rect 297 252 298 253
rect 296 252 297 253
rect 295 252 296 253
rect 294 252 295 253
rect 293 252 294 253
rect 292 252 293 253
rect 291 252 292 253
rect 290 252 291 253
rect 289 252 290 253
rect 288 252 289 253
rect 287 252 288 253
rect 286 252 287 253
rect 285 252 286 253
rect 284 252 285 253
rect 283 252 284 253
rect 282 252 283 253
rect 281 252 282 253
rect 280 252 281 253
rect 279 252 280 253
rect 278 252 279 253
rect 277 252 278 253
rect 276 252 277 253
rect 275 252 276 253
rect 274 252 275 253
rect 273 252 274 253
rect 272 252 273 253
rect 271 252 272 253
rect 270 252 271 253
rect 269 252 270 253
rect 268 252 269 253
rect 267 252 268 253
rect 266 252 267 253
rect 265 252 266 253
rect 264 252 265 253
rect 263 252 264 253
rect 262 252 263 253
rect 261 252 262 253
rect 260 252 261 253
rect 259 252 260 253
rect 258 252 259 253
rect 257 252 258 253
rect 256 252 257 253
rect 255 252 256 253
rect 254 252 255 253
rect 253 252 254 253
rect 252 252 253 253
rect 251 252 252 253
rect 250 252 251 253
rect 249 252 250 253
rect 248 252 249 253
rect 247 252 248 253
rect 246 252 247 253
rect 245 252 246 253
rect 244 252 245 253
rect 243 252 244 253
rect 242 252 243 253
rect 241 252 242 253
rect 240 252 241 253
rect 239 252 240 253
rect 238 252 239 253
rect 237 252 238 253
rect 236 252 237 253
rect 235 252 236 253
rect 234 252 235 253
rect 233 252 234 253
rect 232 252 233 253
rect 231 252 232 253
rect 160 252 161 253
rect 159 252 160 253
rect 158 252 159 253
rect 157 252 158 253
rect 156 252 157 253
rect 155 252 156 253
rect 154 252 155 253
rect 153 252 154 253
rect 152 252 153 253
rect 151 252 152 253
rect 150 252 151 253
rect 149 252 150 253
rect 148 252 149 253
rect 147 252 148 253
rect 146 252 147 253
rect 145 252 146 253
rect 144 252 145 253
rect 143 252 144 253
rect 142 252 143 253
rect 141 252 142 253
rect 140 252 141 253
rect 139 252 140 253
rect 138 252 139 253
rect 137 252 138 253
rect 136 252 137 253
rect 135 252 136 253
rect 134 252 135 253
rect 133 252 134 253
rect 132 252 133 253
rect 131 252 132 253
rect 130 252 131 253
rect 129 252 130 253
rect 128 252 129 253
rect 127 252 128 253
rect 126 252 127 253
rect 125 252 126 253
rect 124 252 125 253
rect 123 252 124 253
rect 122 252 123 253
rect 121 252 122 253
rect 108 252 109 253
rect 107 252 108 253
rect 106 252 107 253
rect 105 252 106 253
rect 104 252 105 253
rect 103 252 104 253
rect 102 252 103 253
rect 101 252 102 253
rect 100 252 101 253
rect 99 252 100 253
rect 98 252 99 253
rect 97 252 98 253
rect 96 252 97 253
rect 95 252 96 253
rect 94 252 95 253
rect 93 252 94 253
rect 92 252 93 253
rect 91 252 92 253
rect 90 252 91 253
rect 89 252 90 253
rect 88 252 89 253
rect 87 252 88 253
rect 86 252 87 253
rect 85 252 86 253
rect 84 252 85 253
rect 83 252 84 253
rect 82 252 83 253
rect 81 252 82 253
rect 80 252 81 253
rect 79 252 80 253
rect 78 252 79 253
rect 77 252 78 253
rect 76 252 77 253
rect 75 252 76 253
rect 74 252 75 253
rect 73 252 74 253
rect 72 252 73 253
rect 71 252 72 253
rect 70 252 71 253
rect 69 252 70 253
rect 68 252 69 253
rect 67 252 68 253
rect 66 252 67 253
rect 65 252 66 253
rect 64 252 65 253
rect 63 252 64 253
rect 62 252 63 253
rect 61 252 62 253
rect 60 252 61 253
rect 59 252 60 253
rect 58 252 59 253
rect 57 252 58 253
rect 56 252 57 253
rect 55 252 56 253
rect 54 252 55 253
rect 53 252 54 253
rect 52 252 53 253
rect 51 252 52 253
rect 50 252 51 253
rect 49 252 50 253
rect 48 252 49 253
rect 47 252 48 253
rect 46 252 47 253
rect 45 252 46 253
rect 44 252 45 253
rect 43 252 44 253
rect 42 252 43 253
rect 41 252 42 253
rect 40 252 41 253
rect 39 252 40 253
rect 38 252 39 253
rect 37 252 38 253
rect 36 252 37 253
rect 35 252 36 253
rect 34 252 35 253
rect 33 252 34 253
rect 32 252 33 253
rect 21 252 22 253
rect 20 252 21 253
rect 19 252 20 253
rect 18 252 19 253
rect 17 252 18 253
rect 16 252 17 253
rect 15 252 16 253
rect 14 252 15 253
rect 13 252 14 253
rect 12 252 13 253
rect 11 252 12 253
rect 10 252 11 253
rect 9 252 10 253
rect 8 252 9 253
rect 7 252 8 253
rect 6 252 7 253
rect 5 252 6 253
rect 4 252 5 253
rect 3 252 4 253
rect 480 253 481 254
rect 479 253 480 254
rect 474 253 475 254
rect 473 253 474 254
rect 472 253 473 254
rect 471 253 472 254
rect 470 253 471 254
rect 469 253 470 254
rect 460 253 461 254
rect 459 253 460 254
rect 312 253 313 254
rect 311 253 312 254
rect 310 253 311 254
rect 309 253 310 254
rect 308 253 309 254
rect 307 253 308 254
rect 306 253 307 254
rect 305 253 306 254
rect 304 253 305 254
rect 303 253 304 254
rect 302 253 303 254
rect 301 253 302 254
rect 300 253 301 254
rect 299 253 300 254
rect 298 253 299 254
rect 297 253 298 254
rect 296 253 297 254
rect 295 253 296 254
rect 294 253 295 254
rect 293 253 294 254
rect 292 253 293 254
rect 291 253 292 254
rect 290 253 291 254
rect 289 253 290 254
rect 288 253 289 254
rect 287 253 288 254
rect 286 253 287 254
rect 285 253 286 254
rect 284 253 285 254
rect 283 253 284 254
rect 282 253 283 254
rect 281 253 282 254
rect 280 253 281 254
rect 279 253 280 254
rect 278 253 279 254
rect 277 253 278 254
rect 276 253 277 254
rect 275 253 276 254
rect 274 253 275 254
rect 273 253 274 254
rect 272 253 273 254
rect 271 253 272 254
rect 270 253 271 254
rect 269 253 270 254
rect 268 253 269 254
rect 267 253 268 254
rect 266 253 267 254
rect 265 253 266 254
rect 264 253 265 254
rect 263 253 264 254
rect 262 253 263 254
rect 261 253 262 254
rect 260 253 261 254
rect 259 253 260 254
rect 258 253 259 254
rect 257 253 258 254
rect 256 253 257 254
rect 255 253 256 254
rect 254 253 255 254
rect 253 253 254 254
rect 252 253 253 254
rect 251 253 252 254
rect 250 253 251 254
rect 249 253 250 254
rect 248 253 249 254
rect 247 253 248 254
rect 246 253 247 254
rect 245 253 246 254
rect 244 253 245 254
rect 243 253 244 254
rect 242 253 243 254
rect 241 253 242 254
rect 240 253 241 254
rect 239 253 240 254
rect 238 253 239 254
rect 237 253 238 254
rect 236 253 237 254
rect 235 253 236 254
rect 234 253 235 254
rect 233 253 234 254
rect 232 253 233 254
rect 231 253 232 254
rect 230 253 231 254
rect 162 253 163 254
rect 161 253 162 254
rect 160 253 161 254
rect 159 253 160 254
rect 158 253 159 254
rect 157 253 158 254
rect 156 253 157 254
rect 155 253 156 254
rect 154 253 155 254
rect 153 253 154 254
rect 152 253 153 254
rect 151 253 152 254
rect 150 253 151 254
rect 149 253 150 254
rect 148 253 149 254
rect 147 253 148 254
rect 146 253 147 254
rect 145 253 146 254
rect 144 253 145 254
rect 143 253 144 254
rect 142 253 143 254
rect 141 253 142 254
rect 140 253 141 254
rect 139 253 140 254
rect 138 253 139 254
rect 137 253 138 254
rect 136 253 137 254
rect 135 253 136 254
rect 134 253 135 254
rect 133 253 134 254
rect 132 253 133 254
rect 131 253 132 254
rect 130 253 131 254
rect 129 253 130 254
rect 128 253 129 254
rect 127 253 128 254
rect 126 253 127 254
rect 125 253 126 254
rect 124 253 125 254
rect 123 253 124 254
rect 122 253 123 254
rect 121 253 122 254
rect 108 253 109 254
rect 107 253 108 254
rect 106 253 107 254
rect 105 253 106 254
rect 104 253 105 254
rect 103 253 104 254
rect 102 253 103 254
rect 101 253 102 254
rect 100 253 101 254
rect 99 253 100 254
rect 98 253 99 254
rect 97 253 98 254
rect 96 253 97 254
rect 95 253 96 254
rect 94 253 95 254
rect 93 253 94 254
rect 92 253 93 254
rect 91 253 92 254
rect 90 253 91 254
rect 89 253 90 254
rect 88 253 89 254
rect 87 253 88 254
rect 86 253 87 254
rect 85 253 86 254
rect 84 253 85 254
rect 83 253 84 254
rect 82 253 83 254
rect 81 253 82 254
rect 80 253 81 254
rect 79 253 80 254
rect 78 253 79 254
rect 77 253 78 254
rect 76 253 77 254
rect 75 253 76 254
rect 74 253 75 254
rect 73 253 74 254
rect 72 253 73 254
rect 71 253 72 254
rect 70 253 71 254
rect 69 253 70 254
rect 68 253 69 254
rect 67 253 68 254
rect 66 253 67 254
rect 65 253 66 254
rect 64 253 65 254
rect 63 253 64 254
rect 62 253 63 254
rect 61 253 62 254
rect 60 253 61 254
rect 59 253 60 254
rect 58 253 59 254
rect 57 253 58 254
rect 56 253 57 254
rect 55 253 56 254
rect 54 253 55 254
rect 53 253 54 254
rect 52 253 53 254
rect 51 253 52 254
rect 50 253 51 254
rect 49 253 50 254
rect 48 253 49 254
rect 47 253 48 254
rect 46 253 47 254
rect 45 253 46 254
rect 44 253 45 254
rect 43 253 44 254
rect 42 253 43 254
rect 41 253 42 254
rect 40 253 41 254
rect 39 253 40 254
rect 38 253 39 254
rect 37 253 38 254
rect 36 253 37 254
rect 35 253 36 254
rect 34 253 35 254
rect 33 253 34 254
rect 32 253 33 254
rect 21 253 22 254
rect 20 253 21 254
rect 19 253 20 254
rect 18 253 19 254
rect 17 253 18 254
rect 16 253 17 254
rect 15 253 16 254
rect 14 253 15 254
rect 13 253 14 254
rect 12 253 13 254
rect 11 253 12 254
rect 10 253 11 254
rect 9 253 10 254
rect 8 253 9 254
rect 7 253 8 254
rect 6 253 7 254
rect 5 253 6 254
rect 4 253 5 254
rect 3 253 4 254
rect 480 254 481 255
rect 479 254 480 255
rect 478 254 479 255
rect 477 254 478 255
rect 476 254 477 255
rect 475 254 476 255
rect 474 254 475 255
rect 473 254 474 255
rect 472 254 473 255
rect 471 254 472 255
rect 470 254 471 255
rect 469 254 470 255
rect 461 254 462 255
rect 460 254 461 255
rect 459 254 460 255
rect 311 254 312 255
rect 310 254 311 255
rect 309 254 310 255
rect 308 254 309 255
rect 307 254 308 255
rect 306 254 307 255
rect 305 254 306 255
rect 304 254 305 255
rect 303 254 304 255
rect 302 254 303 255
rect 301 254 302 255
rect 300 254 301 255
rect 299 254 300 255
rect 298 254 299 255
rect 297 254 298 255
rect 296 254 297 255
rect 295 254 296 255
rect 294 254 295 255
rect 293 254 294 255
rect 292 254 293 255
rect 291 254 292 255
rect 290 254 291 255
rect 289 254 290 255
rect 288 254 289 255
rect 287 254 288 255
rect 286 254 287 255
rect 285 254 286 255
rect 284 254 285 255
rect 283 254 284 255
rect 282 254 283 255
rect 281 254 282 255
rect 280 254 281 255
rect 279 254 280 255
rect 278 254 279 255
rect 277 254 278 255
rect 276 254 277 255
rect 275 254 276 255
rect 274 254 275 255
rect 273 254 274 255
rect 272 254 273 255
rect 271 254 272 255
rect 270 254 271 255
rect 269 254 270 255
rect 268 254 269 255
rect 267 254 268 255
rect 266 254 267 255
rect 265 254 266 255
rect 264 254 265 255
rect 263 254 264 255
rect 262 254 263 255
rect 261 254 262 255
rect 260 254 261 255
rect 259 254 260 255
rect 258 254 259 255
rect 257 254 258 255
rect 256 254 257 255
rect 255 254 256 255
rect 254 254 255 255
rect 253 254 254 255
rect 252 254 253 255
rect 251 254 252 255
rect 250 254 251 255
rect 249 254 250 255
rect 248 254 249 255
rect 247 254 248 255
rect 246 254 247 255
rect 245 254 246 255
rect 244 254 245 255
rect 243 254 244 255
rect 242 254 243 255
rect 241 254 242 255
rect 240 254 241 255
rect 239 254 240 255
rect 238 254 239 255
rect 237 254 238 255
rect 236 254 237 255
rect 235 254 236 255
rect 234 254 235 255
rect 233 254 234 255
rect 232 254 233 255
rect 231 254 232 255
rect 230 254 231 255
rect 164 254 165 255
rect 163 254 164 255
rect 162 254 163 255
rect 161 254 162 255
rect 160 254 161 255
rect 159 254 160 255
rect 158 254 159 255
rect 157 254 158 255
rect 156 254 157 255
rect 155 254 156 255
rect 154 254 155 255
rect 153 254 154 255
rect 152 254 153 255
rect 151 254 152 255
rect 150 254 151 255
rect 149 254 150 255
rect 148 254 149 255
rect 147 254 148 255
rect 146 254 147 255
rect 145 254 146 255
rect 144 254 145 255
rect 143 254 144 255
rect 142 254 143 255
rect 141 254 142 255
rect 140 254 141 255
rect 139 254 140 255
rect 138 254 139 255
rect 137 254 138 255
rect 136 254 137 255
rect 135 254 136 255
rect 134 254 135 255
rect 133 254 134 255
rect 132 254 133 255
rect 131 254 132 255
rect 130 254 131 255
rect 129 254 130 255
rect 128 254 129 255
rect 127 254 128 255
rect 126 254 127 255
rect 125 254 126 255
rect 124 254 125 255
rect 123 254 124 255
rect 122 254 123 255
rect 121 254 122 255
rect 109 254 110 255
rect 108 254 109 255
rect 107 254 108 255
rect 106 254 107 255
rect 105 254 106 255
rect 104 254 105 255
rect 103 254 104 255
rect 102 254 103 255
rect 101 254 102 255
rect 100 254 101 255
rect 99 254 100 255
rect 98 254 99 255
rect 97 254 98 255
rect 96 254 97 255
rect 95 254 96 255
rect 94 254 95 255
rect 93 254 94 255
rect 92 254 93 255
rect 91 254 92 255
rect 90 254 91 255
rect 89 254 90 255
rect 88 254 89 255
rect 87 254 88 255
rect 86 254 87 255
rect 85 254 86 255
rect 84 254 85 255
rect 83 254 84 255
rect 82 254 83 255
rect 81 254 82 255
rect 80 254 81 255
rect 79 254 80 255
rect 78 254 79 255
rect 77 254 78 255
rect 76 254 77 255
rect 75 254 76 255
rect 74 254 75 255
rect 73 254 74 255
rect 72 254 73 255
rect 71 254 72 255
rect 70 254 71 255
rect 69 254 70 255
rect 68 254 69 255
rect 67 254 68 255
rect 66 254 67 255
rect 65 254 66 255
rect 64 254 65 255
rect 63 254 64 255
rect 62 254 63 255
rect 61 254 62 255
rect 60 254 61 255
rect 59 254 60 255
rect 58 254 59 255
rect 54 254 55 255
rect 53 254 54 255
rect 52 254 53 255
rect 51 254 52 255
rect 50 254 51 255
rect 49 254 50 255
rect 48 254 49 255
rect 47 254 48 255
rect 46 254 47 255
rect 45 254 46 255
rect 44 254 45 255
rect 43 254 44 255
rect 42 254 43 255
rect 41 254 42 255
rect 40 254 41 255
rect 39 254 40 255
rect 38 254 39 255
rect 37 254 38 255
rect 36 254 37 255
rect 35 254 36 255
rect 34 254 35 255
rect 33 254 34 255
rect 32 254 33 255
rect 22 254 23 255
rect 21 254 22 255
rect 20 254 21 255
rect 19 254 20 255
rect 18 254 19 255
rect 17 254 18 255
rect 16 254 17 255
rect 15 254 16 255
rect 14 254 15 255
rect 13 254 14 255
rect 12 254 13 255
rect 11 254 12 255
rect 10 254 11 255
rect 9 254 10 255
rect 8 254 9 255
rect 7 254 8 255
rect 6 254 7 255
rect 5 254 6 255
rect 4 254 5 255
rect 3 254 4 255
rect 479 255 480 256
rect 478 255 479 256
rect 477 255 478 256
rect 476 255 477 256
rect 475 255 476 256
rect 474 255 475 256
rect 473 255 474 256
rect 472 255 473 256
rect 471 255 472 256
rect 470 255 471 256
rect 463 255 464 256
rect 462 255 463 256
rect 461 255 462 256
rect 460 255 461 256
rect 309 255 310 256
rect 308 255 309 256
rect 307 255 308 256
rect 306 255 307 256
rect 305 255 306 256
rect 304 255 305 256
rect 303 255 304 256
rect 302 255 303 256
rect 301 255 302 256
rect 300 255 301 256
rect 299 255 300 256
rect 298 255 299 256
rect 297 255 298 256
rect 296 255 297 256
rect 295 255 296 256
rect 294 255 295 256
rect 293 255 294 256
rect 292 255 293 256
rect 291 255 292 256
rect 290 255 291 256
rect 289 255 290 256
rect 288 255 289 256
rect 287 255 288 256
rect 286 255 287 256
rect 285 255 286 256
rect 284 255 285 256
rect 283 255 284 256
rect 282 255 283 256
rect 281 255 282 256
rect 280 255 281 256
rect 279 255 280 256
rect 278 255 279 256
rect 277 255 278 256
rect 276 255 277 256
rect 275 255 276 256
rect 274 255 275 256
rect 273 255 274 256
rect 272 255 273 256
rect 271 255 272 256
rect 270 255 271 256
rect 269 255 270 256
rect 268 255 269 256
rect 267 255 268 256
rect 266 255 267 256
rect 265 255 266 256
rect 264 255 265 256
rect 263 255 264 256
rect 262 255 263 256
rect 261 255 262 256
rect 260 255 261 256
rect 259 255 260 256
rect 258 255 259 256
rect 257 255 258 256
rect 256 255 257 256
rect 255 255 256 256
rect 254 255 255 256
rect 253 255 254 256
rect 252 255 253 256
rect 251 255 252 256
rect 250 255 251 256
rect 249 255 250 256
rect 248 255 249 256
rect 247 255 248 256
rect 246 255 247 256
rect 245 255 246 256
rect 244 255 245 256
rect 243 255 244 256
rect 242 255 243 256
rect 241 255 242 256
rect 240 255 241 256
rect 239 255 240 256
rect 238 255 239 256
rect 237 255 238 256
rect 236 255 237 256
rect 235 255 236 256
rect 234 255 235 256
rect 233 255 234 256
rect 232 255 233 256
rect 231 255 232 256
rect 230 255 231 256
rect 166 255 167 256
rect 165 255 166 256
rect 164 255 165 256
rect 163 255 164 256
rect 162 255 163 256
rect 161 255 162 256
rect 160 255 161 256
rect 159 255 160 256
rect 158 255 159 256
rect 157 255 158 256
rect 156 255 157 256
rect 155 255 156 256
rect 154 255 155 256
rect 153 255 154 256
rect 152 255 153 256
rect 151 255 152 256
rect 150 255 151 256
rect 149 255 150 256
rect 148 255 149 256
rect 147 255 148 256
rect 146 255 147 256
rect 145 255 146 256
rect 144 255 145 256
rect 143 255 144 256
rect 142 255 143 256
rect 141 255 142 256
rect 140 255 141 256
rect 139 255 140 256
rect 138 255 139 256
rect 137 255 138 256
rect 136 255 137 256
rect 135 255 136 256
rect 134 255 135 256
rect 133 255 134 256
rect 132 255 133 256
rect 131 255 132 256
rect 130 255 131 256
rect 129 255 130 256
rect 128 255 129 256
rect 127 255 128 256
rect 126 255 127 256
rect 125 255 126 256
rect 124 255 125 256
rect 123 255 124 256
rect 122 255 123 256
rect 109 255 110 256
rect 108 255 109 256
rect 107 255 108 256
rect 106 255 107 256
rect 105 255 106 256
rect 104 255 105 256
rect 103 255 104 256
rect 102 255 103 256
rect 101 255 102 256
rect 100 255 101 256
rect 99 255 100 256
rect 98 255 99 256
rect 97 255 98 256
rect 96 255 97 256
rect 95 255 96 256
rect 94 255 95 256
rect 93 255 94 256
rect 92 255 93 256
rect 91 255 92 256
rect 90 255 91 256
rect 89 255 90 256
rect 88 255 89 256
rect 87 255 88 256
rect 86 255 87 256
rect 85 255 86 256
rect 84 255 85 256
rect 83 255 84 256
rect 82 255 83 256
rect 81 255 82 256
rect 80 255 81 256
rect 79 255 80 256
rect 78 255 79 256
rect 77 255 78 256
rect 76 255 77 256
rect 75 255 76 256
rect 74 255 75 256
rect 73 255 74 256
rect 72 255 73 256
rect 71 255 72 256
rect 70 255 71 256
rect 69 255 70 256
rect 68 255 69 256
rect 67 255 68 256
rect 66 255 67 256
rect 65 255 66 256
rect 64 255 65 256
rect 63 255 64 256
rect 54 255 55 256
rect 53 255 54 256
rect 52 255 53 256
rect 51 255 52 256
rect 50 255 51 256
rect 49 255 50 256
rect 48 255 49 256
rect 47 255 48 256
rect 46 255 47 256
rect 45 255 46 256
rect 44 255 45 256
rect 43 255 44 256
rect 42 255 43 256
rect 41 255 42 256
rect 40 255 41 256
rect 39 255 40 256
rect 38 255 39 256
rect 37 255 38 256
rect 36 255 37 256
rect 35 255 36 256
rect 34 255 35 256
rect 33 255 34 256
rect 22 255 23 256
rect 21 255 22 256
rect 20 255 21 256
rect 19 255 20 256
rect 18 255 19 256
rect 17 255 18 256
rect 16 255 17 256
rect 15 255 16 256
rect 14 255 15 256
rect 13 255 14 256
rect 12 255 13 256
rect 11 255 12 256
rect 10 255 11 256
rect 9 255 10 256
rect 8 255 9 256
rect 7 255 8 256
rect 6 255 7 256
rect 5 255 6 256
rect 4 255 5 256
rect 3 255 4 256
rect 478 256 479 257
rect 477 256 478 257
rect 476 256 477 257
rect 475 256 476 257
rect 474 256 475 257
rect 473 256 474 257
rect 472 256 473 257
rect 471 256 472 257
rect 464 256 465 257
rect 463 256 464 257
rect 462 256 463 257
rect 461 256 462 257
rect 460 256 461 257
rect 308 256 309 257
rect 307 256 308 257
rect 306 256 307 257
rect 305 256 306 257
rect 304 256 305 257
rect 303 256 304 257
rect 302 256 303 257
rect 301 256 302 257
rect 300 256 301 257
rect 299 256 300 257
rect 298 256 299 257
rect 297 256 298 257
rect 296 256 297 257
rect 295 256 296 257
rect 294 256 295 257
rect 293 256 294 257
rect 292 256 293 257
rect 291 256 292 257
rect 290 256 291 257
rect 289 256 290 257
rect 288 256 289 257
rect 287 256 288 257
rect 286 256 287 257
rect 285 256 286 257
rect 284 256 285 257
rect 283 256 284 257
rect 282 256 283 257
rect 281 256 282 257
rect 280 256 281 257
rect 279 256 280 257
rect 278 256 279 257
rect 277 256 278 257
rect 276 256 277 257
rect 275 256 276 257
rect 274 256 275 257
rect 273 256 274 257
rect 272 256 273 257
rect 271 256 272 257
rect 270 256 271 257
rect 269 256 270 257
rect 268 256 269 257
rect 267 256 268 257
rect 266 256 267 257
rect 265 256 266 257
rect 264 256 265 257
rect 263 256 264 257
rect 262 256 263 257
rect 261 256 262 257
rect 260 256 261 257
rect 259 256 260 257
rect 258 256 259 257
rect 257 256 258 257
rect 256 256 257 257
rect 255 256 256 257
rect 254 256 255 257
rect 253 256 254 257
rect 252 256 253 257
rect 251 256 252 257
rect 250 256 251 257
rect 249 256 250 257
rect 248 256 249 257
rect 247 256 248 257
rect 246 256 247 257
rect 245 256 246 257
rect 244 256 245 257
rect 243 256 244 257
rect 242 256 243 257
rect 241 256 242 257
rect 240 256 241 257
rect 239 256 240 257
rect 238 256 239 257
rect 237 256 238 257
rect 236 256 237 257
rect 235 256 236 257
rect 234 256 235 257
rect 233 256 234 257
rect 232 256 233 257
rect 231 256 232 257
rect 230 256 231 257
rect 168 256 169 257
rect 167 256 168 257
rect 166 256 167 257
rect 165 256 166 257
rect 164 256 165 257
rect 163 256 164 257
rect 162 256 163 257
rect 161 256 162 257
rect 160 256 161 257
rect 159 256 160 257
rect 158 256 159 257
rect 157 256 158 257
rect 156 256 157 257
rect 155 256 156 257
rect 154 256 155 257
rect 153 256 154 257
rect 152 256 153 257
rect 151 256 152 257
rect 150 256 151 257
rect 149 256 150 257
rect 148 256 149 257
rect 147 256 148 257
rect 146 256 147 257
rect 145 256 146 257
rect 144 256 145 257
rect 143 256 144 257
rect 142 256 143 257
rect 141 256 142 257
rect 140 256 141 257
rect 139 256 140 257
rect 138 256 139 257
rect 137 256 138 257
rect 136 256 137 257
rect 135 256 136 257
rect 134 256 135 257
rect 133 256 134 257
rect 132 256 133 257
rect 131 256 132 257
rect 130 256 131 257
rect 129 256 130 257
rect 128 256 129 257
rect 127 256 128 257
rect 126 256 127 257
rect 125 256 126 257
rect 124 256 125 257
rect 123 256 124 257
rect 122 256 123 257
rect 109 256 110 257
rect 108 256 109 257
rect 107 256 108 257
rect 106 256 107 257
rect 105 256 106 257
rect 104 256 105 257
rect 103 256 104 257
rect 102 256 103 257
rect 101 256 102 257
rect 100 256 101 257
rect 99 256 100 257
rect 98 256 99 257
rect 97 256 98 257
rect 96 256 97 257
rect 95 256 96 257
rect 94 256 95 257
rect 93 256 94 257
rect 92 256 93 257
rect 91 256 92 257
rect 90 256 91 257
rect 89 256 90 257
rect 88 256 89 257
rect 87 256 88 257
rect 86 256 87 257
rect 85 256 86 257
rect 84 256 85 257
rect 83 256 84 257
rect 82 256 83 257
rect 81 256 82 257
rect 80 256 81 257
rect 79 256 80 257
rect 78 256 79 257
rect 77 256 78 257
rect 76 256 77 257
rect 75 256 76 257
rect 74 256 75 257
rect 73 256 74 257
rect 72 256 73 257
rect 71 256 72 257
rect 70 256 71 257
rect 69 256 70 257
rect 68 256 69 257
rect 67 256 68 257
rect 66 256 67 257
rect 65 256 66 257
rect 54 256 55 257
rect 53 256 54 257
rect 52 256 53 257
rect 51 256 52 257
rect 50 256 51 257
rect 49 256 50 257
rect 48 256 49 257
rect 47 256 48 257
rect 46 256 47 257
rect 45 256 46 257
rect 44 256 45 257
rect 43 256 44 257
rect 42 256 43 257
rect 41 256 42 257
rect 40 256 41 257
rect 39 256 40 257
rect 38 256 39 257
rect 37 256 38 257
rect 36 256 37 257
rect 35 256 36 257
rect 34 256 35 257
rect 33 256 34 257
rect 22 256 23 257
rect 21 256 22 257
rect 20 256 21 257
rect 19 256 20 257
rect 18 256 19 257
rect 17 256 18 257
rect 16 256 17 257
rect 15 256 16 257
rect 14 256 15 257
rect 13 256 14 257
rect 12 256 13 257
rect 11 256 12 257
rect 10 256 11 257
rect 9 256 10 257
rect 8 256 9 257
rect 7 256 8 257
rect 6 256 7 257
rect 5 256 6 257
rect 4 256 5 257
rect 3 256 4 257
rect 477 257 478 258
rect 476 257 477 258
rect 475 257 476 258
rect 474 257 475 258
rect 473 257 474 258
rect 472 257 473 258
rect 307 257 308 258
rect 306 257 307 258
rect 305 257 306 258
rect 304 257 305 258
rect 303 257 304 258
rect 302 257 303 258
rect 301 257 302 258
rect 300 257 301 258
rect 299 257 300 258
rect 298 257 299 258
rect 297 257 298 258
rect 296 257 297 258
rect 295 257 296 258
rect 294 257 295 258
rect 293 257 294 258
rect 292 257 293 258
rect 291 257 292 258
rect 290 257 291 258
rect 289 257 290 258
rect 288 257 289 258
rect 287 257 288 258
rect 286 257 287 258
rect 285 257 286 258
rect 284 257 285 258
rect 283 257 284 258
rect 282 257 283 258
rect 281 257 282 258
rect 280 257 281 258
rect 279 257 280 258
rect 278 257 279 258
rect 277 257 278 258
rect 276 257 277 258
rect 275 257 276 258
rect 274 257 275 258
rect 273 257 274 258
rect 272 257 273 258
rect 271 257 272 258
rect 270 257 271 258
rect 269 257 270 258
rect 268 257 269 258
rect 267 257 268 258
rect 266 257 267 258
rect 265 257 266 258
rect 264 257 265 258
rect 263 257 264 258
rect 262 257 263 258
rect 261 257 262 258
rect 260 257 261 258
rect 259 257 260 258
rect 258 257 259 258
rect 257 257 258 258
rect 256 257 257 258
rect 255 257 256 258
rect 254 257 255 258
rect 253 257 254 258
rect 252 257 253 258
rect 251 257 252 258
rect 250 257 251 258
rect 249 257 250 258
rect 248 257 249 258
rect 247 257 248 258
rect 246 257 247 258
rect 245 257 246 258
rect 244 257 245 258
rect 243 257 244 258
rect 242 257 243 258
rect 241 257 242 258
rect 240 257 241 258
rect 239 257 240 258
rect 238 257 239 258
rect 237 257 238 258
rect 236 257 237 258
rect 235 257 236 258
rect 234 257 235 258
rect 233 257 234 258
rect 232 257 233 258
rect 231 257 232 258
rect 230 257 231 258
rect 229 257 230 258
rect 170 257 171 258
rect 169 257 170 258
rect 168 257 169 258
rect 167 257 168 258
rect 166 257 167 258
rect 165 257 166 258
rect 164 257 165 258
rect 163 257 164 258
rect 162 257 163 258
rect 161 257 162 258
rect 160 257 161 258
rect 159 257 160 258
rect 158 257 159 258
rect 157 257 158 258
rect 156 257 157 258
rect 155 257 156 258
rect 154 257 155 258
rect 153 257 154 258
rect 152 257 153 258
rect 151 257 152 258
rect 150 257 151 258
rect 149 257 150 258
rect 148 257 149 258
rect 147 257 148 258
rect 146 257 147 258
rect 145 257 146 258
rect 144 257 145 258
rect 143 257 144 258
rect 142 257 143 258
rect 141 257 142 258
rect 140 257 141 258
rect 139 257 140 258
rect 138 257 139 258
rect 137 257 138 258
rect 136 257 137 258
rect 135 257 136 258
rect 134 257 135 258
rect 133 257 134 258
rect 132 257 133 258
rect 131 257 132 258
rect 130 257 131 258
rect 129 257 130 258
rect 128 257 129 258
rect 127 257 128 258
rect 126 257 127 258
rect 125 257 126 258
rect 124 257 125 258
rect 123 257 124 258
rect 122 257 123 258
rect 109 257 110 258
rect 108 257 109 258
rect 107 257 108 258
rect 106 257 107 258
rect 105 257 106 258
rect 104 257 105 258
rect 103 257 104 258
rect 102 257 103 258
rect 101 257 102 258
rect 100 257 101 258
rect 99 257 100 258
rect 98 257 99 258
rect 97 257 98 258
rect 96 257 97 258
rect 95 257 96 258
rect 94 257 95 258
rect 93 257 94 258
rect 92 257 93 258
rect 91 257 92 258
rect 90 257 91 258
rect 89 257 90 258
rect 88 257 89 258
rect 87 257 88 258
rect 86 257 87 258
rect 85 257 86 258
rect 84 257 85 258
rect 83 257 84 258
rect 82 257 83 258
rect 81 257 82 258
rect 80 257 81 258
rect 79 257 80 258
rect 78 257 79 258
rect 77 257 78 258
rect 76 257 77 258
rect 75 257 76 258
rect 74 257 75 258
rect 73 257 74 258
rect 72 257 73 258
rect 71 257 72 258
rect 70 257 71 258
rect 69 257 70 258
rect 68 257 69 258
rect 67 257 68 258
rect 55 257 56 258
rect 54 257 55 258
rect 53 257 54 258
rect 52 257 53 258
rect 51 257 52 258
rect 50 257 51 258
rect 49 257 50 258
rect 48 257 49 258
rect 47 257 48 258
rect 46 257 47 258
rect 45 257 46 258
rect 44 257 45 258
rect 43 257 44 258
rect 42 257 43 258
rect 41 257 42 258
rect 40 257 41 258
rect 39 257 40 258
rect 38 257 39 258
rect 37 257 38 258
rect 36 257 37 258
rect 35 257 36 258
rect 34 257 35 258
rect 33 257 34 258
rect 22 257 23 258
rect 21 257 22 258
rect 20 257 21 258
rect 19 257 20 258
rect 18 257 19 258
rect 17 257 18 258
rect 16 257 17 258
rect 15 257 16 258
rect 14 257 15 258
rect 13 257 14 258
rect 12 257 13 258
rect 11 257 12 258
rect 10 257 11 258
rect 9 257 10 258
rect 8 257 9 258
rect 7 257 8 258
rect 6 257 7 258
rect 5 257 6 258
rect 4 257 5 258
rect 3 257 4 258
rect 306 258 307 259
rect 305 258 306 259
rect 304 258 305 259
rect 303 258 304 259
rect 302 258 303 259
rect 301 258 302 259
rect 300 258 301 259
rect 299 258 300 259
rect 298 258 299 259
rect 297 258 298 259
rect 296 258 297 259
rect 295 258 296 259
rect 294 258 295 259
rect 293 258 294 259
rect 292 258 293 259
rect 291 258 292 259
rect 290 258 291 259
rect 289 258 290 259
rect 288 258 289 259
rect 287 258 288 259
rect 286 258 287 259
rect 285 258 286 259
rect 284 258 285 259
rect 283 258 284 259
rect 282 258 283 259
rect 281 258 282 259
rect 280 258 281 259
rect 279 258 280 259
rect 278 258 279 259
rect 277 258 278 259
rect 276 258 277 259
rect 275 258 276 259
rect 274 258 275 259
rect 273 258 274 259
rect 272 258 273 259
rect 271 258 272 259
rect 270 258 271 259
rect 269 258 270 259
rect 268 258 269 259
rect 267 258 268 259
rect 266 258 267 259
rect 265 258 266 259
rect 264 258 265 259
rect 263 258 264 259
rect 262 258 263 259
rect 261 258 262 259
rect 260 258 261 259
rect 259 258 260 259
rect 258 258 259 259
rect 257 258 258 259
rect 256 258 257 259
rect 255 258 256 259
rect 254 258 255 259
rect 253 258 254 259
rect 252 258 253 259
rect 251 258 252 259
rect 250 258 251 259
rect 249 258 250 259
rect 248 258 249 259
rect 247 258 248 259
rect 246 258 247 259
rect 245 258 246 259
rect 244 258 245 259
rect 243 258 244 259
rect 242 258 243 259
rect 241 258 242 259
rect 240 258 241 259
rect 239 258 240 259
rect 238 258 239 259
rect 237 258 238 259
rect 236 258 237 259
rect 235 258 236 259
rect 234 258 235 259
rect 233 258 234 259
rect 232 258 233 259
rect 231 258 232 259
rect 230 258 231 259
rect 229 258 230 259
rect 173 258 174 259
rect 172 258 173 259
rect 171 258 172 259
rect 170 258 171 259
rect 169 258 170 259
rect 168 258 169 259
rect 167 258 168 259
rect 166 258 167 259
rect 165 258 166 259
rect 164 258 165 259
rect 163 258 164 259
rect 162 258 163 259
rect 161 258 162 259
rect 160 258 161 259
rect 159 258 160 259
rect 158 258 159 259
rect 157 258 158 259
rect 156 258 157 259
rect 155 258 156 259
rect 154 258 155 259
rect 153 258 154 259
rect 152 258 153 259
rect 151 258 152 259
rect 150 258 151 259
rect 149 258 150 259
rect 148 258 149 259
rect 147 258 148 259
rect 146 258 147 259
rect 145 258 146 259
rect 144 258 145 259
rect 143 258 144 259
rect 142 258 143 259
rect 141 258 142 259
rect 140 258 141 259
rect 139 258 140 259
rect 138 258 139 259
rect 137 258 138 259
rect 136 258 137 259
rect 135 258 136 259
rect 134 258 135 259
rect 133 258 134 259
rect 132 258 133 259
rect 131 258 132 259
rect 130 258 131 259
rect 129 258 130 259
rect 128 258 129 259
rect 127 258 128 259
rect 126 258 127 259
rect 125 258 126 259
rect 124 258 125 259
rect 123 258 124 259
rect 122 258 123 259
rect 109 258 110 259
rect 108 258 109 259
rect 107 258 108 259
rect 106 258 107 259
rect 105 258 106 259
rect 104 258 105 259
rect 103 258 104 259
rect 102 258 103 259
rect 101 258 102 259
rect 100 258 101 259
rect 99 258 100 259
rect 98 258 99 259
rect 97 258 98 259
rect 96 258 97 259
rect 95 258 96 259
rect 94 258 95 259
rect 93 258 94 259
rect 92 258 93 259
rect 91 258 92 259
rect 90 258 91 259
rect 89 258 90 259
rect 88 258 89 259
rect 87 258 88 259
rect 86 258 87 259
rect 85 258 86 259
rect 84 258 85 259
rect 83 258 84 259
rect 82 258 83 259
rect 81 258 82 259
rect 80 258 81 259
rect 79 258 80 259
rect 78 258 79 259
rect 77 258 78 259
rect 76 258 77 259
rect 75 258 76 259
rect 74 258 75 259
rect 73 258 74 259
rect 72 258 73 259
rect 71 258 72 259
rect 70 258 71 259
rect 69 258 70 259
rect 68 258 69 259
rect 55 258 56 259
rect 54 258 55 259
rect 53 258 54 259
rect 52 258 53 259
rect 51 258 52 259
rect 50 258 51 259
rect 49 258 50 259
rect 48 258 49 259
rect 47 258 48 259
rect 46 258 47 259
rect 45 258 46 259
rect 44 258 45 259
rect 43 258 44 259
rect 42 258 43 259
rect 41 258 42 259
rect 40 258 41 259
rect 39 258 40 259
rect 38 258 39 259
rect 37 258 38 259
rect 36 258 37 259
rect 35 258 36 259
rect 34 258 35 259
rect 22 258 23 259
rect 21 258 22 259
rect 20 258 21 259
rect 19 258 20 259
rect 18 258 19 259
rect 17 258 18 259
rect 16 258 17 259
rect 15 258 16 259
rect 14 258 15 259
rect 13 258 14 259
rect 12 258 13 259
rect 11 258 12 259
rect 10 258 11 259
rect 9 258 10 259
rect 8 258 9 259
rect 7 258 8 259
rect 6 258 7 259
rect 5 258 6 259
rect 4 258 5 259
rect 3 258 4 259
rect 305 259 306 260
rect 304 259 305 260
rect 303 259 304 260
rect 302 259 303 260
rect 301 259 302 260
rect 300 259 301 260
rect 299 259 300 260
rect 298 259 299 260
rect 297 259 298 260
rect 296 259 297 260
rect 295 259 296 260
rect 294 259 295 260
rect 293 259 294 260
rect 292 259 293 260
rect 291 259 292 260
rect 290 259 291 260
rect 289 259 290 260
rect 288 259 289 260
rect 287 259 288 260
rect 286 259 287 260
rect 285 259 286 260
rect 284 259 285 260
rect 283 259 284 260
rect 282 259 283 260
rect 281 259 282 260
rect 280 259 281 260
rect 279 259 280 260
rect 278 259 279 260
rect 277 259 278 260
rect 276 259 277 260
rect 275 259 276 260
rect 274 259 275 260
rect 273 259 274 260
rect 272 259 273 260
rect 271 259 272 260
rect 270 259 271 260
rect 269 259 270 260
rect 268 259 269 260
rect 267 259 268 260
rect 266 259 267 260
rect 265 259 266 260
rect 264 259 265 260
rect 263 259 264 260
rect 262 259 263 260
rect 261 259 262 260
rect 260 259 261 260
rect 259 259 260 260
rect 258 259 259 260
rect 257 259 258 260
rect 256 259 257 260
rect 255 259 256 260
rect 254 259 255 260
rect 253 259 254 260
rect 252 259 253 260
rect 251 259 252 260
rect 250 259 251 260
rect 249 259 250 260
rect 248 259 249 260
rect 247 259 248 260
rect 246 259 247 260
rect 245 259 246 260
rect 244 259 245 260
rect 243 259 244 260
rect 242 259 243 260
rect 241 259 242 260
rect 240 259 241 260
rect 239 259 240 260
rect 238 259 239 260
rect 237 259 238 260
rect 236 259 237 260
rect 235 259 236 260
rect 234 259 235 260
rect 233 259 234 260
rect 232 259 233 260
rect 231 259 232 260
rect 230 259 231 260
rect 229 259 230 260
rect 177 259 178 260
rect 176 259 177 260
rect 175 259 176 260
rect 174 259 175 260
rect 173 259 174 260
rect 172 259 173 260
rect 171 259 172 260
rect 170 259 171 260
rect 169 259 170 260
rect 168 259 169 260
rect 167 259 168 260
rect 166 259 167 260
rect 165 259 166 260
rect 164 259 165 260
rect 163 259 164 260
rect 162 259 163 260
rect 161 259 162 260
rect 160 259 161 260
rect 159 259 160 260
rect 158 259 159 260
rect 157 259 158 260
rect 156 259 157 260
rect 155 259 156 260
rect 154 259 155 260
rect 153 259 154 260
rect 152 259 153 260
rect 151 259 152 260
rect 150 259 151 260
rect 149 259 150 260
rect 148 259 149 260
rect 147 259 148 260
rect 146 259 147 260
rect 145 259 146 260
rect 144 259 145 260
rect 143 259 144 260
rect 142 259 143 260
rect 141 259 142 260
rect 140 259 141 260
rect 139 259 140 260
rect 138 259 139 260
rect 137 259 138 260
rect 136 259 137 260
rect 135 259 136 260
rect 134 259 135 260
rect 133 259 134 260
rect 132 259 133 260
rect 131 259 132 260
rect 130 259 131 260
rect 129 259 130 260
rect 128 259 129 260
rect 127 259 128 260
rect 126 259 127 260
rect 125 259 126 260
rect 124 259 125 260
rect 123 259 124 260
rect 122 259 123 260
rect 110 259 111 260
rect 109 259 110 260
rect 108 259 109 260
rect 107 259 108 260
rect 106 259 107 260
rect 105 259 106 260
rect 104 259 105 260
rect 103 259 104 260
rect 102 259 103 260
rect 101 259 102 260
rect 100 259 101 260
rect 99 259 100 260
rect 98 259 99 260
rect 97 259 98 260
rect 96 259 97 260
rect 95 259 96 260
rect 94 259 95 260
rect 93 259 94 260
rect 92 259 93 260
rect 91 259 92 260
rect 90 259 91 260
rect 89 259 90 260
rect 88 259 89 260
rect 87 259 88 260
rect 86 259 87 260
rect 85 259 86 260
rect 84 259 85 260
rect 83 259 84 260
rect 82 259 83 260
rect 81 259 82 260
rect 80 259 81 260
rect 79 259 80 260
rect 78 259 79 260
rect 77 259 78 260
rect 76 259 77 260
rect 75 259 76 260
rect 74 259 75 260
rect 73 259 74 260
rect 72 259 73 260
rect 71 259 72 260
rect 70 259 71 260
rect 69 259 70 260
rect 55 259 56 260
rect 54 259 55 260
rect 53 259 54 260
rect 52 259 53 260
rect 51 259 52 260
rect 50 259 51 260
rect 49 259 50 260
rect 48 259 49 260
rect 47 259 48 260
rect 46 259 47 260
rect 45 259 46 260
rect 44 259 45 260
rect 43 259 44 260
rect 42 259 43 260
rect 41 259 42 260
rect 40 259 41 260
rect 39 259 40 260
rect 38 259 39 260
rect 37 259 38 260
rect 36 259 37 260
rect 35 259 36 260
rect 34 259 35 260
rect 23 259 24 260
rect 22 259 23 260
rect 21 259 22 260
rect 20 259 21 260
rect 19 259 20 260
rect 18 259 19 260
rect 17 259 18 260
rect 16 259 17 260
rect 15 259 16 260
rect 14 259 15 260
rect 13 259 14 260
rect 12 259 13 260
rect 11 259 12 260
rect 10 259 11 260
rect 9 259 10 260
rect 8 259 9 260
rect 7 259 8 260
rect 6 259 7 260
rect 5 259 6 260
rect 4 259 5 260
rect 3 259 4 260
rect 304 260 305 261
rect 303 260 304 261
rect 302 260 303 261
rect 301 260 302 261
rect 300 260 301 261
rect 299 260 300 261
rect 298 260 299 261
rect 297 260 298 261
rect 296 260 297 261
rect 295 260 296 261
rect 294 260 295 261
rect 293 260 294 261
rect 292 260 293 261
rect 291 260 292 261
rect 290 260 291 261
rect 289 260 290 261
rect 288 260 289 261
rect 287 260 288 261
rect 286 260 287 261
rect 285 260 286 261
rect 284 260 285 261
rect 283 260 284 261
rect 282 260 283 261
rect 281 260 282 261
rect 280 260 281 261
rect 279 260 280 261
rect 278 260 279 261
rect 277 260 278 261
rect 276 260 277 261
rect 275 260 276 261
rect 274 260 275 261
rect 273 260 274 261
rect 272 260 273 261
rect 271 260 272 261
rect 270 260 271 261
rect 269 260 270 261
rect 268 260 269 261
rect 267 260 268 261
rect 266 260 267 261
rect 265 260 266 261
rect 264 260 265 261
rect 263 260 264 261
rect 262 260 263 261
rect 261 260 262 261
rect 260 260 261 261
rect 259 260 260 261
rect 258 260 259 261
rect 257 260 258 261
rect 256 260 257 261
rect 255 260 256 261
rect 254 260 255 261
rect 253 260 254 261
rect 252 260 253 261
rect 251 260 252 261
rect 250 260 251 261
rect 249 260 250 261
rect 248 260 249 261
rect 247 260 248 261
rect 246 260 247 261
rect 245 260 246 261
rect 244 260 245 261
rect 243 260 244 261
rect 242 260 243 261
rect 241 260 242 261
rect 240 260 241 261
rect 239 260 240 261
rect 238 260 239 261
rect 237 260 238 261
rect 236 260 237 261
rect 235 260 236 261
rect 234 260 235 261
rect 233 260 234 261
rect 232 260 233 261
rect 231 260 232 261
rect 230 260 231 261
rect 229 260 230 261
rect 228 260 229 261
rect 181 260 182 261
rect 180 260 181 261
rect 179 260 180 261
rect 178 260 179 261
rect 177 260 178 261
rect 176 260 177 261
rect 175 260 176 261
rect 174 260 175 261
rect 173 260 174 261
rect 172 260 173 261
rect 171 260 172 261
rect 170 260 171 261
rect 169 260 170 261
rect 168 260 169 261
rect 167 260 168 261
rect 166 260 167 261
rect 165 260 166 261
rect 164 260 165 261
rect 163 260 164 261
rect 162 260 163 261
rect 161 260 162 261
rect 160 260 161 261
rect 159 260 160 261
rect 158 260 159 261
rect 157 260 158 261
rect 156 260 157 261
rect 155 260 156 261
rect 154 260 155 261
rect 153 260 154 261
rect 152 260 153 261
rect 151 260 152 261
rect 150 260 151 261
rect 149 260 150 261
rect 148 260 149 261
rect 147 260 148 261
rect 146 260 147 261
rect 145 260 146 261
rect 144 260 145 261
rect 143 260 144 261
rect 142 260 143 261
rect 141 260 142 261
rect 140 260 141 261
rect 139 260 140 261
rect 138 260 139 261
rect 137 260 138 261
rect 136 260 137 261
rect 135 260 136 261
rect 134 260 135 261
rect 133 260 134 261
rect 132 260 133 261
rect 131 260 132 261
rect 130 260 131 261
rect 129 260 130 261
rect 128 260 129 261
rect 127 260 128 261
rect 126 260 127 261
rect 125 260 126 261
rect 124 260 125 261
rect 123 260 124 261
rect 122 260 123 261
rect 110 260 111 261
rect 109 260 110 261
rect 108 260 109 261
rect 107 260 108 261
rect 106 260 107 261
rect 105 260 106 261
rect 104 260 105 261
rect 103 260 104 261
rect 102 260 103 261
rect 101 260 102 261
rect 100 260 101 261
rect 99 260 100 261
rect 98 260 99 261
rect 97 260 98 261
rect 96 260 97 261
rect 95 260 96 261
rect 94 260 95 261
rect 93 260 94 261
rect 92 260 93 261
rect 91 260 92 261
rect 90 260 91 261
rect 89 260 90 261
rect 88 260 89 261
rect 87 260 88 261
rect 86 260 87 261
rect 85 260 86 261
rect 84 260 85 261
rect 83 260 84 261
rect 82 260 83 261
rect 81 260 82 261
rect 80 260 81 261
rect 79 260 80 261
rect 78 260 79 261
rect 77 260 78 261
rect 76 260 77 261
rect 75 260 76 261
rect 74 260 75 261
rect 73 260 74 261
rect 72 260 73 261
rect 71 260 72 261
rect 70 260 71 261
rect 55 260 56 261
rect 54 260 55 261
rect 53 260 54 261
rect 52 260 53 261
rect 51 260 52 261
rect 50 260 51 261
rect 49 260 50 261
rect 48 260 49 261
rect 47 260 48 261
rect 46 260 47 261
rect 45 260 46 261
rect 44 260 45 261
rect 43 260 44 261
rect 42 260 43 261
rect 41 260 42 261
rect 40 260 41 261
rect 39 260 40 261
rect 38 260 39 261
rect 37 260 38 261
rect 36 260 37 261
rect 35 260 36 261
rect 34 260 35 261
rect 23 260 24 261
rect 22 260 23 261
rect 21 260 22 261
rect 20 260 21 261
rect 19 260 20 261
rect 18 260 19 261
rect 17 260 18 261
rect 16 260 17 261
rect 15 260 16 261
rect 14 260 15 261
rect 13 260 14 261
rect 12 260 13 261
rect 11 260 12 261
rect 10 260 11 261
rect 9 260 10 261
rect 8 260 9 261
rect 7 260 8 261
rect 6 260 7 261
rect 5 260 6 261
rect 4 260 5 261
rect 3 260 4 261
rect 303 261 304 262
rect 302 261 303 262
rect 301 261 302 262
rect 300 261 301 262
rect 299 261 300 262
rect 298 261 299 262
rect 297 261 298 262
rect 296 261 297 262
rect 295 261 296 262
rect 294 261 295 262
rect 293 261 294 262
rect 292 261 293 262
rect 291 261 292 262
rect 290 261 291 262
rect 289 261 290 262
rect 288 261 289 262
rect 287 261 288 262
rect 286 261 287 262
rect 285 261 286 262
rect 284 261 285 262
rect 283 261 284 262
rect 282 261 283 262
rect 281 261 282 262
rect 280 261 281 262
rect 279 261 280 262
rect 278 261 279 262
rect 277 261 278 262
rect 276 261 277 262
rect 275 261 276 262
rect 274 261 275 262
rect 273 261 274 262
rect 272 261 273 262
rect 271 261 272 262
rect 270 261 271 262
rect 269 261 270 262
rect 268 261 269 262
rect 267 261 268 262
rect 266 261 267 262
rect 265 261 266 262
rect 264 261 265 262
rect 263 261 264 262
rect 262 261 263 262
rect 261 261 262 262
rect 260 261 261 262
rect 259 261 260 262
rect 258 261 259 262
rect 257 261 258 262
rect 256 261 257 262
rect 255 261 256 262
rect 254 261 255 262
rect 253 261 254 262
rect 252 261 253 262
rect 251 261 252 262
rect 250 261 251 262
rect 249 261 250 262
rect 248 261 249 262
rect 247 261 248 262
rect 246 261 247 262
rect 245 261 246 262
rect 244 261 245 262
rect 243 261 244 262
rect 242 261 243 262
rect 241 261 242 262
rect 240 261 241 262
rect 239 261 240 262
rect 238 261 239 262
rect 237 261 238 262
rect 236 261 237 262
rect 235 261 236 262
rect 234 261 235 262
rect 233 261 234 262
rect 232 261 233 262
rect 231 261 232 262
rect 230 261 231 262
rect 229 261 230 262
rect 228 261 229 262
rect 185 261 186 262
rect 184 261 185 262
rect 183 261 184 262
rect 182 261 183 262
rect 181 261 182 262
rect 180 261 181 262
rect 179 261 180 262
rect 178 261 179 262
rect 177 261 178 262
rect 176 261 177 262
rect 175 261 176 262
rect 174 261 175 262
rect 173 261 174 262
rect 172 261 173 262
rect 171 261 172 262
rect 170 261 171 262
rect 169 261 170 262
rect 168 261 169 262
rect 167 261 168 262
rect 166 261 167 262
rect 165 261 166 262
rect 164 261 165 262
rect 163 261 164 262
rect 162 261 163 262
rect 161 261 162 262
rect 160 261 161 262
rect 159 261 160 262
rect 158 261 159 262
rect 157 261 158 262
rect 156 261 157 262
rect 155 261 156 262
rect 154 261 155 262
rect 153 261 154 262
rect 152 261 153 262
rect 151 261 152 262
rect 150 261 151 262
rect 149 261 150 262
rect 148 261 149 262
rect 147 261 148 262
rect 146 261 147 262
rect 145 261 146 262
rect 144 261 145 262
rect 143 261 144 262
rect 142 261 143 262
rect 141 261 142 262
rect 140 261 141 262
rect 139 261 140 262
rect 138 261 139 262
rect 137 261 138 262
rect 136 261 137 262
rect 135 261 136 262
rect 134 261 135 262
rect 133 261 134 262
rect 132 261 133 262
rect 131 261 132 262
rect 130 261 131 262
rect 129 261 130 262
rect 128 261 129 262
rect 127 261 128 262
rect 126 261 127 262
rect 125 261 126 262
rect 124 261 125 262
rect 123 261 124 262
rect 110 261 111 262
rect 109 261 110 262
rect 108 261 109 262
rect 107 261 108 262
rect 106 261 107 262
rect 105 261 106 262
rect 104 261 105 262
rect 103 261 104 262
rect 102 261 103 262
rect 101 261 102 262
rect 100 261 101 262
rect 99 261 100 262
rect 98 261 99 262
rect 97 261 98 262
rect 96 261 97 262
rect 95 261 96 262
rect 94 261 95 262
rect 93 261 94 262
rect 92 261 93 262
rect 91 261 92 262
rect 90 261 91 262
rect 89 261 90 262
rect 88 261 89 262
rect 87 261 88 262
rect 86 261 87 262
rect 85 261 86 262
rect 84 261 85 262
rect 83 261 84 262
rect 82 261 83 262
rect 81 261 82 262
rect 80 261 81 262
rect 79 261 80 262
rect 78 261 79 262
rect 77 261 78 262
rect 76 261 77 262
rect 75 261 76 262
rect 74 261 75 262
rect 73 261 74 262
rect 72 261 73 262
rect 71 261 72 262
rect 56 261 57 262
rect 55 261 56 262
rect 54 261 55 262
rect 53 261 54 262
rect 52 261 53 262
rect 51 261 52 262
rect 50 261 51 262
rect 49 261 50 262
rect 48 261 49 262
rect 47 261 48 262
rect 46 261 47 262
rect 45 261 46 262
rect 44 261 45 262
rect 43 261 44 262
rect 42 261 43 262
rect 41 261 42 262
rect 40 261 41 262
rect 39 261 40 262
rect 38 261 39 262
rect 37 261 38 262
rect 36 261 37 262
rect 35 261 36 262
rect 23 261 24 262
rect 22 261 23 262
rect 21 261 22 262
rect 20 261 21 262
rect 19 261 20 262
rect 18 261 19 262
rect 17 261 18 262
rect 16 261 17 262
rect 15 261 16 262
rect 14 261 15 262
rect 13 261 14 262
rect 12 261 13 262
rect 11 261 12 262
rect 10 261 11 262
rect 9 261 10 262
rect 8 261 9 262
rect 7 261 8 262
rect 6 261 7 262
rect 5 261 6 262
rect 4 261 5 262
rect 3 261 4 262
rect 302 262 303 263
rect 301 262 302 263
rect 300 262 301 263
rect 299 262 300 263
rect 298 262 299 263
rect 297 262 298 263
rect 296 262 297 263
rect 295 262 296 263
rect 294 262 295 263
rect 293 262 294 263
rect 292 262 293 263
rect 291 262 292 263
rect 290 262 291 263
rect 289 262 290 263
rect 288 262 289 263
rect 287 262 288 263
rect 286 262 287 263
rect 285 262 286 263
rect 284 262 285 263
rect 283 262 284 263
rect 282 262 283 263
rect 281 262 282 263
rect 280 262 281 263
rect 279 262 280 263
rect 278 262 279 263
rect 277 262 278 263
rect 276 262 277 263
rect 275 262 276 263
rect 274 262 275 263
rect 273 262 274 263
rect 272 262 273 263
rect 271 262 272 263
rect 270 262 271 263
rect 269 262 270 263
rect 268 262 269 263
rect 267 262 268 263
rect 266 262 267 263
rect 265 262 266 263
rect 264 262 265 263
rect 263 262 264 263
rect 262 262 263 263
rect 261 262 262 263
rect 260 262 261 263
rect 259 262 260 263
rect 258 262 259 263
rect 257 262 258 263
rect 256 262 257 263
rect 255 262 256 263
rect 254 262 255 263
rect 253 262 254 263
rect 252 262 253 263
rect 251 262 252 263
rect 250 262 251 263
rect 249 262 250 263
rect 248 262 249 263
rect 247 262 248 263
rect 246 262 247 263
rect 245 262 246 263
rect 244 262 245 263
rect 243 262 244 263
rect 242 262 243 263
rect 241 262 242 263
rect 240 262 241 263
rect 239 262 240 263
rect 238 262 239 263
rect 237 262 238 263
rect 236 262 237 263
rect 235 262 236 263
rect 234 262 235 263
rect 233 262 234 263
rect 232 262 233 263
rect 231 262 232 263
rect 230 262 231 263
rect 229 262 230 263
rect 228 262 229 263
rect 207 262 208 263
rect 206 262 207 263
rect 205 262 206 263
rect 204 262 205 263
rect 203 262 204 263
rect 202 262 203 263
rect 192 262 193 263
rect 191 262 192 263
rect 190 262 191 263
rect 189 262 190 263
rect 188 262 189 263
rect 187 262 188 263
rect 186 262 187 263
rect 185 262 186 263
rect 184 262 185 263
rect 183 262 184 263
rect 182 262 183 263
rect 181 262 182 263
rect 180 262 181 263
rect 179 262 180 263
rect 178 262 179 263
rect 177 262 178 263
rect 176 262 177 263
rect 175 262 176 263
rect 174 262 175 263
rect 173 262 174 263
rect 172 262 173 263
rect 171 262 172 263
rect 170 262 171 263
rect 169 262 170 263
rect 168 262 169 263
rect 167 262 168 263
rect 166 262 167 263
rect 165 262 166 263
rect 164 262 165 263
rect 163 262 164 263
rect 162 262 163 263
rect 161 262 162 263
rect 160 262 161 263
rect 159 262 160 263
rect 158 262 159 263
rect 157 262 158 263
rect 156 262 157 263
rect 155 262 156 263
rect 154 262 155 263
rect 153 262 154 263
rect 152 262 153 263
rect 151 262 152 263
rect 150 262 151 263
rect 149 262 150 263
rect 148 262 149 263
rect 147 262 148 263
rect 146 262 147 263
rect 145 262 146 263
rect 144 262 145 263
rect 143 262 144 263
rect 142 262 143 263
rect 141 262 142 263
rect 140 262 141 263
rect 139 262 140 263
rect 138 262 139 263
rect 137 262 138 263
rect 136 262 137 263
rect 135 262 136 263
rect 134 262 135 263
rect 133 262 134 263
rect 132 262 133 263
rect 131 262 132 263
rect 130 262 131 263
rect 129 262 130 263
rect 128 262 129 263
rect 127 262 128 263
rect 126 262 127 263
rect 125 262 126 263
rect 124 262 125 263
rect 123 262 124 263
rect 110 262 111 263
rect 109 262 110 263
rect 108 262 109 263
rect 107 262 108 263
rect 106 262 107 263
rect 105 262 106 263
rect 104 262 105 263
rect 103 262 104 263
rect 102 262 103 263
rect 101 262 102 263
rect 100 262 101 263
rect 99 262 100 263
rect 98 262 99 263
rect 97 262 98 263
rect 96 262 97 263
rect 95 262 96 263
rect 94 262 95 263
rect 93 262 94 263
rect 92 262 93 263
rect 91 262 92 263
rect 90 262 91 263
rect 89 262 90 263
rect 88 262 89 263
rect 87 262 88 263
rect 86 262 87 263
rect 85 262 86 263
rect 84 262 85 263
rect 83 262 84 263
rect 82 262 83 263
rect 81 262 82 263
rect 80 262 81 263
rect 79 262 80 263
rect 78 262 79 263
rect 77 262 78 263
rect 76 262 77 263
rect 75 262 76 263
rect 74 262 75 263
rect 73 262 74 263
rect 72 262 73 263
rect 56 262 57 263
rect 55 262 56 263
rect 54 262 55 263
rect 53 262 54 263
rect 52 262 53 263
rect 51 262 52 263
rect 50 262 51 263
rect 49 262 50 263
rect 48 262 49 263
rect 47 262 48 263
rect 46 262 47 263
rect 45 262 46 263
rect 44 262 45 263
rect 43 262 44 263
rect 42 262 43 263
rect 41 262 42 263
rect 40 262 41 263
rect 39 262 40 263
rect 38 262 39 263
rect 37 262 38 263
rect 36 262 37 263
rect 35 262 36 263
rect 24 262 25 263
rect 23 262 24 263
rect 22 262 23 263
rect 21 262 22 263
rect 20 262 21 263
rect 19 262 20 263
rect 18 262 19 263
rect 17 262 18 263
rect 16 262 17 263
rect 15 262 16 263
rect 14 262 15 263
rect 13 262 14 263
rect 12 262 13 263
rect 11 262 12 263
rect 10 262 11 263
rect 9 262 10 263
rect 8 262 9 263
rect 7 262 8 263
rect 6 262 7 263
rect 5 262 6 263
rect 4 262 5 263
rect 3 262 4 263
rect 302 263 303 264
rect 301 263 302 264
rect 300 263 301 264
rect 299 263 300 264
rect 298 263 299 264
rect 297 263 298 264
rect 296 263 297 264
rect 295 263 296 264
rect 294 263 295 264
rect 293 263 294 264
rect 292 263 293 264
rect 291 263 292 264
rect 290 263 291 264
rect 289 263 290 264
rect 288 263 289 264
rect 287 263 288 264
rect 286 263 287 264
rect 285 263 286 264
rect 284 263 285 264
rect 283 263 284 264
rect 282 263 283 264
rect 281 263 282 264
rect 280 263 281 264
rect 279 263 280 264
rect 278 263 279 264
rect 277 263 278 264
rect 276 263 277 264
rect 275 263 276 264
rect 274 263 275 264
rect 273 263 274 264
rect 272 263 273 264
rect 271 263 272 264
rect 270 263 271 264
rect 269 263 270 264
rect 268 263 269 264
rect 267 263 268 264
rect 266 263 267 264
rect 265 263 266 264
rect 264 263 265 264
rect 263 263 264 264
rect 262 263 263 264
rect 261 263 262 264
rect 260 263 261 264
rect 259 263 260 264
rect 258 263 259 264
rect 257 263 258 264
rect 256 263 257 264
rect 255 263 256 264
rect 254 263 255 264
rect 253 263 254 264
rect 252 263 253 264
rect 251 263 252 264
rect 250 263 251 264
rect 249 263 250 264
rect 248 263 249 264
rect 247 263 248 264
rect 246 263 247 264
rect 245 263 246 264
rect 244 263 245 264
rect 243 263 244 264
rect 242 263 243 264
rect 241 263 242 264
rect 240 263 241 264
rect 239 263 240 264
rect 238 263 239 264
rect 237 263 238 264
rect 236 263 237 264
rect 235 263 236 264
rect 234 263 235 264
rect 233 263 234 264
rect 232 263 233 264
rect 231 263 232 264
rect 230 263 231 264
rect 229 263 230 264
rect 228 263 229 264
rect 227 263 228 264
rect 206 263 207 264
rect 205 263 206 264
rect 204 263 205 264
rect 203 263 204 264
rect 202 263 203 264
rect 201 263 202 264
rect 200 263 201 264
rect 199 263 200 264
rect 198 263 199 264
rect 197 263 198 264
rect 196 263 197 264
rect 195 263 196 264
rect 194 263 195 264
rect 193 263 194 264
rect 192 263 193 264
rect 191 263 192 264
rect 190 263 191 264
rect 189 263 190 264
rect 188 263 189 264
rect 187 263 188 264
rect 186 263 187 264
rect 185 263 186 264
rect 184 263 185 264
rect 183 263 184 264
rect 182 263 183 264
rect 181 263 182 264
rect 180 263 181 264
rect 179 263 180 264
rect 178 263 179 264
rect 177 263 178 264
rect 176 263 177 264
rect 175 263 176 264
rect 174 263 175 264
rect 173 263 174 264
rect 172 263 173 264
rect 171 263 172 264
rect 170 263 171 264
rect 169 263 170 264
rect 168 263 169 264
rect 167 263 168 264
rect 166 263 167 264
rect 165 263 166 264
rect 164 263 165 264
rect 163 263 164 264
rect 162 263 163 264
rect 161 263 162 264
rect 160 263 161 264
rect 159 263 160 264
rect 158 263 159 264
rect 157 263 158 264
rect 156 263 157 264
rect 155 263 156 264
rect 154 263 155 264
rect 153 263 154 264
rect 152 263 153 264
rect 151 263 152 264
rect 150 263 151 264
rect 149 263 150 264
rect 148 263 149 264
rect 147 263 148 264
rect 146 263 147 264
rect 145 263 146 264
rect 144 263 145 264
rect 143 263 144 264
rect 142 263 143 264
rect 141 263 142 264
rect 140 263 141 264
rect 139 263 140 264
rect 138 263 139 264
rect 137 263 138 264
rect 136 263 137 264
rect 135 263 136 264
rect 134 263 135 264
rect 133 263 134 264
rect 132 263 133 264
rect 131 263 132 264
rect 130 263 131 264
rect 129 263 130 264
rect 128 263 129 264
rect 127 263 128 264
rect 126 263 127 264
rect 125 263 126 264
rect 124 263 125 264
rect 123 263 124 264
rect 110 263 111 264
rect 109 263 110 264
rect 108 263 109 264
rect 107 263 108 264
rect 106 263 107 264
rect 105 263 106 264
rect 104 263 105 264
rect 103 263 104 264
rect 102 263 103 264
rect 101 263 102 264
rect 100 263 101 264
rect 99 263 100 264
rect 98 263 99 264
rect 97 263 98 264
rect 96 263 97 264
rect 95 263 96 264
rect 94 263 95 264
rect 93 263 94 264
rect 92 263 93 264
rect 91 263 92 264
rect 90 263 91 264
rect 89 263 90 264
rect 88 263 89 264
rect 87 263 88 264
rect 86 263 87 264
rect 85 263 86 264
rect 84 263 85 264
rect 83 263 84 264
rect 82 263 83 264
rect 81 263 82 264
rect 80 263 81 264
rect 79 263 80 264
rect 78 263 79 264
rect 77 263 78 264
rect 76 263 77 264
rect 75 263 76 264
rect 74 263 75 264
rect 73 263 74 264
rect 72 263 73 264
rect 57 263 58 264
rect 56 263 57 264
rect 55 263 56 264
rect 54 263 55 264
rect 53 263 54 264
rect 52 263 53 264
rect 51 263 52 264
rect 50 263 51 264
rect 49 263 50 264
rect 48 263 49 264
rect 47 263 48 264
rect 46 263 47 264
rect 45 263 46 264
rect 44 263 45 264
rect 43 263 44 264
rect 42 263 43 264
rect 41 263 42 264
rect 40 263 41 264
rect 39 263 40 264
rect 38 263 39 264
rect 37 263 38 264
rect 36 263 37 264
rect 35 263 36 264
rect 24 263 25 264
rect 23 263 24 264
rect 22 263 23 264
rect 21 263 22 264
rect 20 263 21 264
rect 19 263 20 264
rect 18 263 19 264
rect 17 263 18 264
rect 16 263 17 264
rect 15 263 16 264
rect 14 263 15 264
rect 13 263 14 264
rect 12 263 13 264
rect 11 263 12 264
rect 10 263 11 264
rect 9 263 10 264
rect 8 263 9 264
rect 7 263 8 264
rect 6 263 7 264
rect 5 263 6 264
rect 4 263 5 264
rect 3 263 4 264
rect 301 264 302 265
rect 300 264 301 265
rect 299 264 300 265
rect 298 264 299 265
rect 297 264 298 265
rect 296 264 297 265
rect 295 264 296 265
rect 294 264 295 265
rect 293 264 294 265
rect 292 264 293 265
rect 291 264 292 265
rect 290 264 291 265
rect 289 264 290 265
rect 288 264 289 265
rect 287 264 288 265
rect 286 264 287 265
rect 285 264 286 265
rect 284 264 285 265
rect 283 264 284 265
rect 282 264 283 265
rect 281 264 282 265
rect 280 264 281 265
rect 279 264 280 265
rect 278 264 279 265
rect 277 264 278 265
rect 276 264 277 265
rect 275 264 276 265
rect 274 264 275 265
rect 273 264 274 265
rect 272 264 273 265
rect 271 264 272 265
rect 270 264 271 265
rect 269 264 270 265
rect 268 264 269 265
rect 267 264 268 265
rect 266 264 267 265
rect 265 264 266 265
rect 264 264 265 265
rect 263 264 264 265
rect 262 264 263 265
rect 261 264 262 265
rect 260 264 261 265
rect 259 264 260 265
rect 258 264 259 265
rect 257 264 258 265
rect 256 264 257 265
rect 255 264 256 265
rect 254 264 255 265
rect 253 264 254 265
rect 252 264 253 265
rect 251 264 252 265
rect 250 264 251 265
rect 249 264 250 265
rect 248 264 249 265
rect 247 264 248 265
rect 246 264 247 265
rect 245 264 246 265
rect 244 264 245 265
rect 243 264 244 265
rect 242 264 243 265
rect 241 264 242 265
rect 240 264 241 265
rect 239 264 240 265
rect 238 264 239 265
rect 237 264 238 265
rect 236 264 237 265
rect 235 264 236 265
rect 234 264 235 265
rect 233 264 234 265
rect 232 264 233 265
rect 231 264 232 265
rect 230 264 231 265
rect 229 264 230 265
rect 228 264 229 265
rect 227 264 228 265
rect 206 264 207 265
rect 205 264 206 265
rect 204 264 205 265
rect 203 264 204 265
rect 202 264 203 265
rect 201 264 202 265
rect 200 264 201 265
rect 199 264 200 265
rect 198 264 199 265
rect 197 264 198 265
rect 196 264 197 265
rect 195 264 196 265
rect 194 264 195 265
rect 193 264 194 265
rect 192 264 193 265
rect 191 264 192 265
rect 190 264 191 265
rect 189 264 190 265
rect 188 264 189 265
rect 187 264 188 265
rect 186 264 187 265
rect 185 264 186 265
rect 184 264 185 265
rect 183 264 184 265
rect 182 264 183 265
rect 181 264 182 265
rect 180 264 181 265
rect 179 264 180 265
rect 178 264 179 265
rect 177 264 178 265
rect 176 264 177 265
rect 175 264 176 265
rect 174 264 175 265
rect 173 264 174 265
rect 172 264 173 265
rect 171 264 172 265
rect 170 264 171 265
rect 169 264 170 265
rect 168 264 169 265
rect 167 264 168 265
rect 166 264 167 265
rect 165 264 166 265
rect 164 264 165 265
rect 163 264 164 265
rect 162 264 163 265
rect 161 264 162 265
rect 160 264 161 265
rect 159 264 160 265
rect 158 264 159 265
rect 157 264 158 265
rect 156 264 157 265
rect 155 264 156 265
rect 154 264 155 265
rect 153 264 154 265
rect 152 264 153 265
rect 151 264 152 265
rect 150 264 151 265
rect 149 264 150 265
rect 148 264 149 265
rect 147 264 148 265
rect 146 264 147 265
rect 145 264 146 265
rect 144 264 145 265
rect 143 264 144 265
rect 142 264 143 265
rect 141 264 142 265
rect 140 264 141 265
rect 139 264 140 265
rect 138 264 139 265
rect 137 264 138 265
rect 136 264 137 265
rect 135 264 136 265
rect 134 264 135 265
rect 133 264 134 265
rect 132 264 133 265
rect 131 264 132 265
rect 130 264 131 265
rect 129 264 130 265
rect 128 264 129 265
rect 127 264 128 265
rect 126 264 127 265
rect 125 264 126 265
rect 124 264 125 265
rect 123 264 124 265
rect 110 264 111 265
rect 109 264 110 265
rect 108 264 109 265
rect 107 264 108 265
rect 106 264 107 265
rect 105 264 106 265
rect 104 264 105 265
rect 103 264 104 265
rect 102 264 103 265
rect 101 264 102 265
rect 100 264 101 265
rect 99 264 100 265
rect 98 264 99 265
rect 97 264 98 265
rect 96 264 97 265
rect 95 264 96 265
rect 94 264 95 265
rect 93 264 94 265
rect 92 264 93 265
rect 91 264 92 265
rect 90 264 91 265
rect 89 264 90 265
rect 88 264 89 265
rect 87 264 88 265
rect 86 264 87 265
rect 85 264 86 265
rect 84 264 85 265
rect 83 264 84 265
rect 82 264 83 265
rect 81 264 82 265
rect 80 264 81 265
rect 79 264 80 265
rect 78 264 79 265
rect 77 264 78 265
rect 76 264 77 265
rect 75 264 76 265
rect 74 264 75 265
rect 73 264 74 265
rect 57 264 58 265
rect 56 264 57 265
rect 55 264 56 265
rect 54 264 55 265
rect 53 264 54 265
rect 52 264 53 265
rect 51 264 52 265
rect 50 264 51 265
rect 49 264 50 265
rect 48 264 49 265
rect 47 264 48 265
rect 46 264 47 265
rect 45 264 46 265
rect 44 264 45 265
rect 43 264 44 265
rect 42 264 43 265
rect 41 264 42 265
rect 40 264 41 265
rect 39 264 40 265
rect 38 264 39 265
rect 37 264 38 265
rect 36 264 37 265
rect 35 264 36 265
rect 24 264 25 265
rect 23 264 24 265
rect 22 264 23 265
rect 21 264 22 265
rect 20 264 21 265
rect 19 264 20 265
rect 18 264 19 265
rect 17 264 18 265
rect 16 264 17 265
rect 15 264 16 265
rect 14 264 15 265
rect 13 264 14 265
rect 12 264 13 265
rect 11 264 12 265
rect 10 264 11 265
rect 9 264 10 265
rect 8 264 9 265
rect 7 264 8 265
rect 6 264 7 265
rect 5 264 6 265
rect 4 264 5 265
rect 3 264 4 265
rect 300 265 301 266
rect 299 265 300 266
rect 298 265 299 266
rect 297 265 298 266
rect 296 265 297 266
rect 295 265 296 266
rect 294 265 295 266
rect 293 265 294 266
rect 292 265 293 266
rect 291 265 292 266
rect 290 265 291 266
rect 289 265 290 266
rect 288 265 289 266
rect 287 265 288 266
rect 286 265 287 266
rect 285 265 286 266
rect 284 265 285 266
rect 283 265 284 266
rect 282 265 283 266
rect 281 265 282 266
rect 280 265 281 266
rect 279 265 280 266
rect 278 265 279 266
rect 277 265 278 266
rect 276 265 277 266
rect 275 265 276 266
rect 274 265 275 266
rect 273 265 274 266
rect 272 265 273 266
rect 271 265 272 266
rect 270 265 271 266
rect 269 265 270 266
rect 268 265 269 266
rect 267 265 268 266
rect 266 265 267 266
rect 265 265 266 266
rect 264 265 265 266
rect 263 265 264 266
rect 262 265 263 266
rect 261 265 262 266
rect 260 265 261 266
rect 259 265 260 266
rect 258 265 259 266
rect 257 265 258 266
rect 256 265 257 266
rect 255 265 256 266
rect 254 265 255 266
rect 253 265 254 266
rect 252 265 253 266
rect 251 265 252 266
rect 250 265 251 266
rect 249 265 250 266
rect 248 265 249 266
rect 247 265 248 266
rect 246 265 247 266
rect 245 265 246 266
rect 244 265 245 266
rect 243 265 244 266
rect 242 265 243 266
rect 241 265 242 266
rect 240 265 241 266
rect 239 265 240 266
rect 238 265 239 266
rect 237 265 238 266
rect 236 265 237 266
rect 235 265 236 266
rect 234 265 235 266
rect 233 265 234 266
rect 232 265 233 266
rect 231 265 232 266
rect 230 265 231 266
rect 229 265 230 266
rect 228 265 229 266
rect 227 265 228 266
rect 206 265 207 266
rect 205 265 206 266
rect 204 265 205 266
rect 203 265 204 266
rect 202 265 203 266
rect 201 265 202 266
rect 200 265 201 266
rect 199 265 200 266
rect 198 265 199 266
rect 197 265 198 266
rect 196 265 197 266
rect 195 265 196 266
rect 194 265 195 266
rect 193 265 194 266
rect 192 265 193 266
rect 191 265 192 266
rect 190 265 191 266
rect 189 265 190 266
rect 188 265 189 266
rect 187 265 188 266
rect 186 265 187 266
rect 185 265 186 266
rect 184 265 185 266
rect 183 265 184 266
rect 182 265 183 266
rect 181 265 182 266
rect 180 265 181 266
rect 179 265 180 266
rect 178 265 179 266
rect 177 265 178 266
rect 176 265 177 266
rect 175 265 176 266
rect 174 265 175 266
rect 173 265 174 266
rect 172 265 173 266
rect 171 265 172 266
rect 170 265 171 266
rect 169 265 170 266
rect 168 265 169 266
rect 167 265 168 266
rect 166 265 167 266
rect 165 265 166 266
rect 164 265 165 266
rect 163 265 164 266
rect 162 265 163 266
rect 161 265 162 266
rect 160 265 161 266
rect 159 265 160 266
rect 158 265 159 266
rect 157 265 158 266
rect 156 265 157 266
rect 155 265 156 266
rect 154 265 155 266
rect 153 265 154 266
rect 152 265 153 266
rect 151 265 152 266
rect 150 265 151 266
rect 149 265 150 266
rect 148 265 149 266
rect 147 265 148 266
rect 146 265 147 266
rect 145 265 146 266
rect 144 265 145 266
rect 143 265 144 266
rect 142 265 143 266
rect 141 265 142 266
rect 140 265 141 266
rect 139 265 140 266
rect 138 265 139 266
rect 137 265 138 266
rect 136 265 137 266
rect 135 265 136 266
rect 134 265 135 266
rect 133 265 134 266
rect 132 265 133 266
rect 131 265 132 266
rect 130 265 131 266
rect 129 265 130 266
rect 128 265 129 266
rect 127 265 128 266
rect 126 265 127 266
rect 125 265 126 266
rect 124 265 125 266
rect 111 265 112 266
rect 110 265 111 266
rect 109 265 110 266
rect 108 265 109 266
rect 107 265 108 266
rect 106 265 107 266
rect 105 265 106 266
rect 104 265 105 266
rect 103 265 104 266
rect 102 265 103 266
rect 101 265 102 266
rect 100 265 101 266
rect 99 265 100 266
rect 98 265 99 266
rect 97 265 98 266
rect 96 265 97 266
rect 95 265 96 266
rect 94 265 95 266
rect 93 265 94 266
rect 92 265 93 266
rect 91 265 92 266
rect 90 265 91 266
rect 89 265 90 266
rect 88 265 89 266
rect 87 265 88 266
rect 86 265 87 266
rect 85 265 86 266
rect 84 265 85 266
rect 83 265 84 266
rect 82 265 83 266
rect 81 265 82 266
rect 80 265 81 266
rect 79 265 80 266
rect 78 265 79 266
rect 77 265 78 266
rect 76 265 77 266
rect 75 265 76 266
rect 74 265 75 266
rect 57 265 58 266
rect 56 265 57 266
rect 55 265 56 266
rect 54 265 55 266
rect 53 265 54 266
rect 52 265 53 266
rect 51 265 52 266
rect 50 265 51 266
rect 49 265 50 266
rect 48 265 49 266
rect 47 265 48 266
rect 46 265 47 266
rect 45 265 46 266
rect 44 265 45 266
rect 43 265 44 266
rect 42 265 43 266
rect 41 265 42 266
rect 40 265 41 266
rect 39 265 40 266
rect 38 265 39 266
rect 37 265 38 266
rect 36 265 37 266
rect 24 265 25 266
rect 23 265 24 266
rect 22 265 23 266
rect 21 265 22 266
rect 20 265 21 266
rect 19 265 20 266
rect 18 265 19 266
rect 17 265 18 266
rect 16 265 17 266
rect 15 265 16 266
rect 14 265 15 266
rect 13 265 14 266
rect 12 265 13 266
rect 11 265 12 266
rect 10 265 11 266
rect 9 265 10 266
rect 8 265 9 266
rect 7 265 8 266
rect 6 265 7 266
rect 5 265 6 266
rect 4 265 5 266
rect 3 265 4 266
rect 480 266 481 267
rect 460 266 461 267
rect 299 266 300 267
rect 298 266 299 267
rect 297 266 298 267
rect 296 266 297 267
rect 295 266 296 267
rect 294 266 295 267
rect 293 266 294 267
rect 292 266 293 267
rect 291 266 292 267
rect 290 266 291 267
rect 289 266 290 267
rect 288 266 289 267
rect 287 266 288 267
rect 286 266 287 267
rect 285 266 286 267
rect 284 266 285 267
rect 283 266 284 267
rect 282 266 283 267
rect 281 266 282 267
rect 280 266 281 267
rect 279 266 280 267
rect 278 266 279 267
rect 277 266 278 267
rect 276 266 277 267
rect 275 266 276 267
rect 274 266 275 267
rect 273 266 274 267
rect 272 266 273 267
rect 271 266 272 267
rect 270 266 271 267
rect 269 266 270 267
rect 268 266 269 267
rect 267 266 268 267
rect 266 266 267 267
rect 265 266 266 267
rect 264 266 265 267
rect 263 266 264 267
rect 262 266 263 267
rect 261 266 262 267
rect 260 266 261 267
rect 259 266 260 267
rect 258 266 259 267
rect 257 266 258 267
rect 256 266 257 267
rect 255 266 256 267
rect 254 266 255 267
rect 253 266 254 267
rect 252 266 253 267
rect 251 266 252 267
rect 250 266 251 267
rect 249 266 250 267
rect 248 266 249 267
rect 247 266 248 267
rect 246 266 247 267
rect 245 266 246 267
rect 244 266 245 267
rect 243 266 244 267
rect 242 266 243 267
rect 241 266 242 267
rect 240 266 241 267
rect 239 266 240 267
rect 238 266 239 267
rect 237 266 238 267
rect 236 266 237 267
rect 235 266 236 267
rect 234 266 235 267
rect 233 266 234 267
rect 232 266 233 267
rect 231 266 232 267
rect 230 266 231 267
rect 229 266 230 267
rect 228 266 229 267
rect 227 266 228 267
rect 226 266 227 267
rect 205 266 206 267
rect 204 266 205 267
rect 203 266 204 267
rect 202 266 203 267
rect 201 266 202 267
rect 200 266 201 267
rect 199 266 200 267
rect 198 266 199 267
rect 197 266 198 267
rect 196 266 197 267
rect 195 266 196 267
rect 194 266 195 267
rect 193 266 194 267
rect 192 266 193 267
rect 191 266 192 267
rect 190 266 191 267
rect 189 266 190 267
rect 188 266 189 267
rect 187 266 188 267
rect 186 266 187 267
rect 185 266 186 267
rect 184 266 185 267
rect 183 266 184 267
rect 182 266 183 267
rect 181 266 182 267
rect 180 266 181 267
rect 179 266 180 267
rect 178 266 179 267
rect 177 266 178 267
rect 176 266 177 267
rect 175 266 176 267
rect 174 266 175 267
rect 173 266 174 267
rect 172 266 173 267
rect 171 266 172 267
rect 170 266 171 267
rect 169 266 170 267
rect 168 266 169 267
rect 167 266 168 267
rect 166 266 167 267
rect 165 266 166 267
rect 164 266 165 267
rect 163 266 164 267
rect 162 266 163 267
rect 161 266 162 267
rect 160 266 161 267
rect 159 266 160 267
rect 158 266 159 267
rect 157 266 158 267
rect 156 266 157 267
rect 155 266 156 267
rect 154 266 155 267
rect 153 266 154 267
rect 152 266 153 267
rect 151 266 152 267
rect 150 266 151 267
rect 149 266 150 267
rect 148 266 149 267
rect 147 266 148 267
rect 146 266 147 267
rect 145 266 146 267
rect 144 266 145 267
rect 143 266 144 267
rect 142 266 143 267
rect 141 266 142 267
rect 140 266 141 267
rect 139 266 140 267
rect 138 266 139 267
rect 137 266 138 267
rect 136 266 137 267
rect 135 266 136 267
rect 134 266 135 267
rect 133 266 134 267
rect 132 266 133 267
rect 131 266 132 267
rect 130 266 131 267
rect 129 266 130 267
rect 128 266 129 267
rect 127 266 128 267
rect 126 266 127 267
rect 125 266 126 267
rect 124 266 125 267
rect 111 266 112 267
rect 110 266 111 267
rect 109 266 110 267
rect 108 266 109 267
rect 107 266 108 267
rect 106 266 107 267
rect 105 266 106 267
rect 104 266 105 267
rect 103 266 104 267
rect 102 266 103 267
rect 101 266 102 267
rect 100 266 101 267
rect 99 266 100 267
rect 98 266 99 267
rect 97 266 98 267
rect 96 266 97 267
rect 95 266 96 267
rect 94 266 95 267
rect 93 266 94 267
rect 92 266 93 267
rect 91 266 92 267
rect 90 266 91 267
rect 89 266 90 267
rect 88 266 89 267
rect 87 266 88 267
rect 86 266 87 267
rect 85 266 86 267
rect 84 266 85 267
rect 83 266 84 267
rect 82 266 83 267
rect 81 266 82 267
rect 80 266 81 267
rect 79 266 80 267
rect 78 266 79 267
rect 77 266 78 267
rect 76 266 77 267
rect 75 266 76 267
rect 74 266 75 267
rect 58 266 59 267
rect 57 266 58 267
rect 56 266 57 267
rect 55 266 56 267
rect 54 266 55 267
rect 53 266 54 267
rect 52 266 53 267
rect 51 266 52 267
rect 50 266 51 267
rect 49 266 50 267
rect 48 266 49 267
rect 47 266 48 267
rect 46 266 47 267
rect 45 266 46 267
rect 44 266 45 267
rect 43 266 44 267
rect 42 266 43 267
rect 41 266 42 267
rect 40 266 41 267
rect 39 266 40 267
rect 38 266 39 267
rect 37 266 38 267
rect 36 266 37 267
rect 25 266 26 267
rect 24 266 25 267
rect 23 266 24 267
rect 22 266 23 267
rect 21 266 22 267
rect 20 266 21 267
rect 19 266 20 267
rect 18 266 19 267
rect 17 266 18 267
rect 16 266 17 267
rect 15 266 16 267
rect 14 266 15 267
rect 13 266 14 267
rect 12 266 13 267
rect 11 266 12 267
rect 10 266 11 267
rect 9 266 10 267
rect 8 266 9 267
rect 7 266 8 267
rect 6 266 7 267
rect 5 266 6 267
rect 4 266 5 267
rect 3 266 4 267
rect 480 267 481 268
rect 460 267 461 268
rect 299 267 300 268
rect 298 267 299 268
rect 297 267 298 268
rect 296 267 297 268
rect 295 267 296 268
rect 294 267 295 268
rect 293 267 294 268
rect 292 267 293 268
rect 291 267 292 268
rect 290 267 291 268
rect 289 267 290 268
rect 288 267 289 268
rect 287 267 288 268
rect 286 267 287 268
rect 285 267 286 268
rect 284 267 285 268
rect 283 267 284 268
rect 282 267 283 268
rect 281 267 282 268
rect 280 267 281 268
rect 279 267 280 268
rect 278 267 279 268
rect 277 267 278 268
rect 276 267 277 268
rect 275 267 276 268
rect 274 267 275 268
rect 273 267 274 268
rect 272 267 273 268
rect 271 267 272 268
rect 270 267 271 268
rect 269 267 270 268
rect 268 267 269 268
rect 267 267 268 268
rect 266 267 267 268
rect 265 267 266 268
rect 264 267 265 268
rect 263 267 264 268
rect 262 267 263 268
rect 261 267 262 268
rect 260 267 261 268
rect 259 267 260 268
rect 258 267 259 268
rect 257 267 258 268
rect 256 267 257 268
rect 255 267 256 268
rect 254 267 255 268
rect 253 267 254 268
rect 252 267 253 268
rect 251 267 252 268
rect 250 267 251 268
rect 249 267 250 268
rect 248 267 249 268
rect 247 267 248 268
rect 246 267 247 268
rect 245 267 246 268
rect 244 267 245 268
rect 243 267 244 268
rect 242 267 243 268
rect 241 267 242 268
rect 240 267 241 268
rect 239 267 240 268
rect 238 267 239 268
rect 237 267 238 268
rect 236 267 237 268
rect 235 267 236 268
rect 234 267 235 268
rect 233 267 234 268
rect 232 267 233 268
rect 231 267 232 268
rect 230 267 231 268
rect 229 267 230 268
rect 228 267 229 268
rect 227 267 228 268
rect 226 267 227 268
rect 205 267 206 268
rect 204 267 205 268
rect 203 267 204 268
rect 202 267 203 268
rect 201 267 202 268
rect 200 267 201 268
rect 199 267 200 268
rect 198 267 199 268
rect 197 267 198 268
rect 196 267 197 268
rect 195 267 196 268
rect 194 267 195 268
rect 193 267 194 268
rect 192 267 193 268
rect 191 267 192 268
rect 190 267 191 268
rect 189 267 190 268
rect 188 267 189 268
rect 187 267 188 268
rect 186 267 187 268
rect 185 267 186 268
rect 184 267 185 268
rect 183 267 184 268
rect 182 267 183 268
rect 181 267 182 268
rect 180 267 181 268
rect 179 267 180 268
rect 178 267 179 268
rect 177 267 178 268
rect 176 267 177 268
rect 175 267 176 268
rect 174 267 175 268
rect 173 267 174 268
rect 172 267 173 268
rect 171 267 172 268
rect 170 267 171 268
rect 169 267 170 268
rect 168 267 169 268
rect 167 267 168 268
rect 166 267 167 268
rect 165 267 166 268
rect 164 267 165 268
rect 163 267 164 268
rect 162 267 163 268
rect 161 267 162 268
rect 160 267 161 268
rect 159 267 160 268
rect 158 267 159 268
rect 157 267 158 268
rect 156 267 157 268
rect 155 267 156 268
rect 154 267 155 268
rect 153 267 154 268
rect 152 267 153 268
rect 151 267 152 268
rect 150 267 151 268
rect 149 267 150 268
rect 148 267 149 268
rect 147 267 148 268
rect 146 267 147 268
rect 145 267 146 268
rect 144 267 145 268
rect 143 267 144 268
rect 142 267 143 268
rect 141 267 142 268
rect 140 267 141 268
rect 139 267 140 268
rect 138 267 139 268
rect 137 267 138 268
rect 136 267 137 268
rect 135 267 136 268
rect 134 267 135 268
rect 133 267 134 268
rect 132 267 133 268
rect 131 267 132 268
rect 130 267 131 268
rect 129 267 130 268
rect 128 267 129 268
rect 127 267 128 268
rect 126 267 127 268
rect 125 267 126 268
rect 124 267 125 268
rect 111 267 112 268
rect 110 267 111 268
rect 109 267 110 268
rect 108 267 109 268
rect 107 267 108 268
rect 106 267 107 268
rect 105 267 106 268
rect 104 267 105 268
rect 103 267 104 268
rect 102 267 103 268
rect 101 267 102 268
rect 100 267 101 268
rect 99 267 100 268
rect 98 267 99 268
rect 97 267 98 268
rect 96 267 97 268
rect 95 267 96 268
rect 94 267 95 268
rect 93 267 94 268
rect 92 267 93 268
rect 91 267 92 268
rect 90 267 91 268
rect 89 267 90 268
rect 88 267 89 268
rect 87 267 88 268
rect 86 267 87 268
rect 85 267 86 268
rect 84 267 85 268
rect 83 267 84 268
rect 82 267 83 268
rect 81 267 82 268
rect 80 267 81 268
rect 79 267 80 268
rect 78 267 79 268
rect 77 267 78 268
rect 76 267 77 268
rect 75 267 76 268
rect 58 267 59 268
rect 57 267 58 268
rect 56 267 57 268
rect 55 267 56 268
rect 54 267 55 268
rect 53 267 54 268
rect 52 267 53 268
rect 51 267 52 268
rect 50 267 51 268
rect 49 267 50 268
rect 48 267 49 268
rect 47 267 48 268
rect 46 267 47 268
rect 45 267 46 268
rect 44 267 45 268
rect 43 267 44 268
rect 42 267 43 268
rect 41 267 42 268
rect 40 267 41 268
rect 39 267 40 268
rect 38 267 39 268
rect 37 267 38 268
rect 36 267 37 268
rect 25 267 26 268
rect 24 267 25 268
rect 23 267 24 268
rect 22 267 23 268
rect 21 267 22 268
rect 20 267 21 268
rect 19 267 20 268
rect 18 267 19 268
rect 17 267 18 268
rect 16 267 17 268
rect 15 267 16 268
rect 14 267 15 268
rect 13 267 14 268
rect 12 267 13 268
rect 11 267 12 268
rect 10 267 11 268
rect 9 267 10 268
rect 8 267 9 268
rect 7 267 8 268
rect 6 267 7 268
rect 5 267 6 268
rect 4 267 5 268
rect 3 267 4 268
rect 480 268 481 269
rect 479 268 480 269
rect 461 268 462 269
rect 460 268 461 269
rect 298 268 299 269
rect 297 268 298 269
rect 296 268 297 269
rect 295 268 296 269
rect 294 268 295 269
rect 293 268 294 269
rect 292 268 293 269
rect 291 268 292 269
rect 290 268 291 269
rect 289 268 290 269
rect 288 268 289 269
rect 287 268 288 269
rect 286 268 287 269
rect 285 268 286 269
rect 284 268 285 269
rect 283 268 284 269
rect 282 268 283 269
rect 281 268 282 269
rect 280 268 281 269
rect 279 268 280 269
rect 278 268 279 269
rect 277 268 278 269
rect 276 268 277 269
rect 275 268 276 269
rect 274 268 275 269
rect 273 268 274 269
rect 272 268 273 269
rect 271 268 272 269
rect 270 268 271 269
rect 269 268 270 269
rect 268 268 269 269
rect 267 268 268 269
rect 266 268 267 269
rect 265 268 266 269
rect 264 268 265 269
rect 263 268 264 269
rect 262 268 263 269
rect 261 268 262 269
rect 260 268 261 269
rect 259 268 260 269
rect 258 268 259 269
rect 257 268 258 269
rect 256 268 257 269
rect 255 268 256 269
rect 254 268 255 269
rect 253 268 254 269
rect 252 268 253 269
rect 251 268 252 269
rect 250 268 251 269
rect 249 268 250 269
rect 248 268 249 269
rect 247 268 248 269
rect 246 268 247 269
rect 245 268 246 269
rect 244 268 245 269
rect 243 268 244 269
rect 242 268 243 269
rect 241 268 242 269
rect 240 268 241 269
rect 239 268 240 269
rect 238 268 239 269
rect 237 268 238 269
rect 236 268 237 269
rect 235 268 236 269
rect 234 268 235 269
rect 233 268 234 269
rect 232 268 233 269
rect 231 268 232 269
rect 230 268 231 269
rect 229 268 230 269
rect 228 268 229 269
rect 227 268 228 269
rect 226 268 227 269
rect 225 268 226 269
rect 204 268 205 269
rect 203 268 204 269
rect 202 268 203 269
rect 201 268 202 269
rect 200 268 201 269
rect 199 268 200 269
rect 198 268 199 269
rect 197 268 198 269
rect 196 268 197 269
rect 195 268 196 269
rect 194 268 195 269
rect 193 268 194 269
rect 192 268 193 269
rect 191 268 192 269
rect 190 268 191 269
rect 189 268 190 269
rect 188 268 189 269
rect 187 268 188 269
rect 186 268 187 269
rect 185 268 186 269
rect 184 268 185 269
rect 183 268 184 269
rect 182 268 183 269
rect 181 268 182 269
rect 180 268 181 269
rect 179 268 180 269
rect 178 268 179 269
rect 177 268 178 269
rect 176 268 177 269
rect 175 268 176 269
rect 174 268 175 269
rect 173 268 174 269
rect 172 268 173 269
rect 171 268 172 269
rect 170 268 171 269
rect 169 268 170 269
rect 168 268 169 269
rect 167 268 168 269
rect 166 268 167 269
rect 165 268 166 269
rect 164 268 165 269
rect 163 268 164 269
rect 162 268 163 269
rect 161 268 162 269
rect 160 268 161 269
rect 159 268 160 269
rect 158 268 159 269
rect 157 268 158 269
rect 156 268 157 269
rect 155 268 156 269
rect 154 268 155 269
rect 153 268 154 269
rect 152 268 153 269
rect 151 268 152 269
rect 150 268 151 269
rect 149 268 150 269
rect 148 268 149 269
rect 147 268 148 269
rect 146 268 147 269
rect 145 268 146 269
rect 144 268 145 269
rect 143 268 144 269
rect 142 268 143 269
rect 141 268 142 269
rect 140 268 141 269
rect 139 268 140 269
rect 138 268 139 269
rect 137 268 138 269
rect 136 268 137 269
rect 135 268 136 269
rect 134 268 135 269
rect 133 268 134 269
rect 132 268 133 269
rect 131 268 132 269
rect 130 268 131 269
rect 129 268 130 269
rect 128 268 129 269
rect 127 268 128 269
rect 126 268 127 269
rect 125 268 126 269
rect 124 268 125 269
rect 111 268 112 269
rect 110 268 111 269
rect 109 268 110 269
rect 108 268 109 269
rect 107 268 108 269
rect 106 268 107 269
rect 105 268 106 269
rect 104 268 105 269
rect 103 268 104 269
rect 102 268 103 269
rect 101 268 102 269
rect 100 268 101 269
rect 99 268 100 269
rect 98 268 99 269
rect 97 268 98 269
rect 96 268 97 269
rect 95 268 96 269
rect 94 268 95 269
rect 93 268 94 269
rect 92 268 93 269
rect 91 268 92 269
rect 90 268 91 269
rect 89 268 90 269
rect 88 268 89 269
rect 87 268 88 269
rect 86 268 87 269
rect 85 268 86 269
rect 84 268 85 269
rect 83 268 84 269
rect 82 268 83 269
rect 81 268 82 269
rect 80 268 81 269
rect 79 268 80 269
rect 78 268 79 269
rect 77 268 78 269
rect 76 268 77 269
rect 75 268 76 269
rect 59 268 60 269
rect 58 268 59 269
rect 57 268 58 269
rect 56 268 57 269
rect 55 268 56 269
rect 54 268 55 269
rect 53 268 54 269
rect 52 268 53 269
rect 51 268 52 269
rect 50 268 51 269
rect 49 268 50 269
rect 48 268 49 269
rect 47 268 48 269
rect 46 268 47 269
rect 45 268 46 269
rect 44 268 45 269
rect 43 268 44 269
rect 42 268 43 269
rect 41 268 42 269
rect 40 268 41 269
rect 39 268 40 269
rect 38 268 39 269
rect 37 268 38 269
rect 36 268 37 269
rect 25 268 26 269
rect 24 268 25 269
rect 23 268 24 269
rect 22 268 23 269
rect 21 268 22 269
rect 20 268 21 269
rect 19 268 20 269
rect 18 268 19 269
rect 17 268 18 269
rect 16 268 17 269
rect 15 268 16 269
rect 14 268 15 269
rect 13 268 14 269
rect 12 268 13 269
rect 11 268 12 269
rect 10 268 11 269
rect 9 268 10 269
rect 8 268 9 269
rect 7 268 8 269
rect 6 268 7 269
rect 5 268 6 269
rect 4 268 5 269
rect 3 268 4 269
rect 480 269 481 270
rect 479 269 480 270
rect 478 269 479 270
rect 477 269 478 270
rect 476 269 477 270
rect 475 269 476 270
rect 474 269 475 270
rect 473 269 474 270
rect 472 269 473 270
rect 471 269 472 270
rect 470 269 471 270
rect 469 269 470 270
rect 468 269 469 270
rect 467 269 468 270
rect 466 269 467 270
rect 465 269 466 270
rect 464 269 465 270
rect 463 269 464 270
rect 462 269 463 270
rect 461 269 462 270
rect 460 269 461 270
rect 297 269 298 270
rect 296 269 297 270
rect 295 269 296 270
rect 294 269 295 270
rect 293 269 294 270
rect 292 269 293 270
rect 291 269 292 270
rect 290 269 291 270
rect 289 269 290 270
rect 288 269 289 270
rect 287 269 288 270
rect 286 269 287 270
rect 285 269 286 270
rect 284 269 285 270
rect 283 269 284 270
rect 282 269 283 270
rect 281 269 282 270
rect 280 269 281 270
rect 279 269 280 270
rect 278 269 279 270
rect 277 269 278 270
rect 276 269 277 270
rect 275 269 276 270
rect 274 269 275 270
rect 273 269 274 270
rect 272 269 273 270
rect 271 269 272 270
rect 270 269 271 270
rect 269 269 270 270
rect 268 269 269 270
rect 267 269 268 270
rect 266 269 267 270
rect 265 269 266 270
rect 264 269 265 270
rect 263 269 264 270
rect 262 269 263 270
rect 261 269 262 270
rect 260 269 261 270
rect 259 269 260 270
rect 258 269 259 270
rect 257 269 258 270
rect 256 269 257 270
rect 255 269 256 270
rect 254 269 255 270
rect 253 269 254 270
rect 252 269 253 270
rect 251 269 252 270
rect 250 269 251 270
rect 249 269 250 270
rect 248 269 249 270
rect 247 269 248 270
rect 246 269 247 270
rect 245 269 246 270
rect 244 269 245 270
rect 243 269 244 270
rect 242 269 243 270
rect 241 269 242 270
rect 240 269 241 270
rect 239 269 240 270
rect 238 269 239 270
rect 237 269 238 270
rect 236 269 237 270
rect 235 269 236 270
rect 234 269 235 270
rect 233 269 234 270
rect 232 269 233 270
rect 231 269 232 270
rect 230 269 231 270
rect 229 269 230 270
rect 228 269 229 270
rect 227 269 228 270
rect 226 269 227 270
rect 225 269 226 270
rect 204 269 205 270
rect 203 269 204 270
rect 202 269 203 270
rect 201 269 202 270
rect 200 269 201 270
rect 199 269 200 270
rect 198 269 199 270
rect 197 269 198 270
rect 196 269 197 270
rect 195 269 196 270
rect 194 269 195 270
rect 193 269 194 270
rect 192 269 193 270
rect 191 269 192 270
rect 190 269 191 270
rect 189 269 190 270
rect 188 269 189 270
rect 187 269 188 270
rect 186 269 187 270
rect 185 269 186 270
rect 184 269 185 270
rect 183 269 184 270
rect 182 269 183 270
rect 181 269 182 270
rect 180 269 181 270
rect 179 269 180 270
rect 178 269 179 270
rect 177 269 178 270
rect 176 269 177 270
rect 175 269 176 270
rect 174 269 175 270
rect 173 269 174 270
rect 172 269 173 270
rect 171 269 172 270
rect 170 269 171 270
rect 169 269 170 270
rect 168 269 169 270
rect 167 269 168 270
rect 166 269 167 270
rect 165 269 166 270
rect 164 269 165 270
rect 163 269 164 270
rect 162 269 163 270
rect 161 269 162 270
rect 160 269 161 270
rect 159 269 160 270
rect 158 269 159 270
rect 157 269 158 270
rect 156 269 157 270
rect 155 269 156 270
rect 154 269 155 270
rect 153 269 154 270
rect 152 269 153 270
rect 151 269 152 270
rect 150 269 151 270
rect 149 269 150 270
rect 148 269 149 270
rect 147 269 148 270
rect 146 269 147 270
rect 145 269 146 270
rect 144 269 145 270
rect 143 269 144 270
rect 142 269 143 270
rect 141 269 142 270
rect 140 269 141 270
rect 139 269 140 270
rect 138 269 139 270
rect 137 269 138 270
rect 136 269 137 270
rect 135 269 136 270
rect 134 269 135 270
rect 133 269 134 270
rect 132 269 133 270
rect 131 269 132 270
rect 130 269 131 270
rect 129 269 130 270
rect 128 269 129 270
rect 127 269 128 270
rect 126 269 127 270
rect 125 269 126 270
rect 111 269 112 270
rect 110 269 111 270
rect 109 269 110 270
rect 108 269 109 270
rect 107 269 108 270
rect 106 269 107 270
rect 105 269 106 270
rect 104 269 105 270
rect 103 269 104 270
rect 102 269 103 270
rect 101 269 102 270
rect 100 269 101 270
rect 99 269 100 270
rect 98 269 99 270
rect 97 269 98 270
rect 96 269 97 270
rect 95 269 96 270
rect 94 269 95 270
rect 93 269 94 270
rect 92 269 93 270
rect 91 269 92 270
rect 90 269 91 270
rect 89 269 90 270
rect 88 269 89 270
rect 87 269 88 270
rect 86 269 87 270
rect 85 269 86 270
rect 84 269 85 270
rect 83 269 84 270
rect 82 269 83 270
rect 81 269 82 270
rect 80 269 81 270
rect 79 269 80 270
rect 78 269 79 270
rect 77 269 78 270
rect 76 269 77 270
rect 59 269 60 270
rect 58 269 59 270
rect 57 269 58 270
rect 56 269 57 270
rect 55 269 56 270
rect 54 269 55 270
rect 53 269 54 270
rect 52 269 53 270
rect 51 269 52 270
rect 50 269 51 270
rect 49 269 50 270
rect 48 269 49 270
rect 47 269 48 270
rect 46 269 47 270
rect 45 269 46 270
rect 44 269 45 270
rect 43 269 44 270
rect 42 269 43 270
rect 41 269 42 270
rect 40 269 41 270
rect 39 269 40 270
rect 38 269 39 270
rect 37 269 38 270
rect 25 269 26 270
rect 24 269 25 270
rect 23 269 24 270
rect 22 269 23 270
rect 21 269 22 270
rect 20 269 21 270
rect 19 269 20 270
rect 18 269 19 270
rect 17 269 18 270
rect 16 269 17 270
rect 15 269 16 270
rect 14 269 15 270
rect 13 269 14 270
rect 12 269 13 270
rect 11 269 12 270
rect 10 269 11 270
rect 9 269 10 270
rect 8 269 9 270
rect 7 269 8 270
rect 6 269 7 270
rect 5 269 6 270
rect 4 269 5 270
rect 3 269 4 270
rect 480 270 481 271
rect 479 270 480 271
rect 478 270 479 271
rect 477 270 478 271
rect 476 270 477 271
rect 475 270 476 271
rect 474 270 475 271
rect 473 270 474 271
rect 472 270 473 271
rect 471 270 472 271
rect 470 270 471 271
rect 469 270 470 271
rect 468 270 469 271
rect 467 270 468 271
rect 466 270 467 271
rect 465 270 466 271
rect 464 270 465 271
rect 463 270 464 271
rect 462 270 463 271
rect 461 270 462 271
rect 460 270 461 271
rect 297 270 298 271
rect 296 270 297 271
rect 295 270 296 271
rect 294 270 295 271
rect 293 270 294 271
rect 292 270 293 271
rect 291 270 292 271
rect 290 270 291 271
rect 289 270 290 271
rect 288 270 289 271
rect 287 270 288 271
rect 286 270 287 271
rect 285 270 286 271
rect 284 270 285 271
rect 283 270 284 271
rect 282 270 283 271
rect 281 270 282 271
rect 280 270 281 271
rect 279 270 280 271
rect 278 270 279 271
rect 277 270 278 271
rect 276 270 277 271
rect 275 270 276 271
rect 274 270 275 271
rect 273 270 274 271
rect 272 270 273 271
rect 271 270 272 271
rect 270 270 271 271
rect 269 270 270 271
rect 268 270 269 271
rect 267 270 268 271
rect 266 270 267 271
rect 265 270 266 271
rect 264 270 265 271
rect 263 270 264 271
rect 262 270 263 271
rect 261 270 262 271
rect 260 270 261 271
rect 259 270 260 271
rect 258 270 259 271
rect 257 270 258 271
rect 256 270 257 271
rect 255 270 256 271
rect 254 270 255 271
rect 253 270 254 271
rect 252 270 253 271
rect 251 270 252 271
rect 250 270 251 271
rect 249 270 250 271
rect 248 270 249 271
rect 247 270 248 271
rect 246 270 247 271
rect 245 270 246 271
rect 244 270 245 271
rect 243 270 244 271
rect 242 270 243 271
rect 241 270 242 271
rect 240 270 241 271
rect 239 270 240 271
rect 238 270 239 271
rect 237 270 238 271
rect 236 270 237 271
rect 235 270 236 271
rect 234 270 235 271
rect 233 270 234 271
rect 232 270 233 271
rect 231 270 232 271
rect 230 270 231 271
rect 229 270 230 271
rect 228 270 229 271
rect 227 270 228 271
rect 226 270 227 271
rect 225 270 226 271
rect 204 270 205 271
rect 203 270 204 271
rect 202 270 203 271
rect 201 270 202 271
rect 200 270 201 271
rect 199 270 200 271
rect 198 270 199 271
rect 197 270 198 271
rect 196 270 197 271
rect 195 270 196 271
rect 194 270 195 271
rect 193 270 194 271
rect 192 270 193 271
rect 191 270 192 271
rect 190 270 191 271
rect 189 270 190 271
rect 188 270 189 271
rect 187 270 188 271
rect 186 270 187 271
rect 185 270 186 271
rect 184 270 185 271
rect 183 270 184 271
rect 182 270 183 271
rect 181 270 182 271
rect 180 270 181 271
rect 179 270 180 271
rect 178 270 179 271
rect 177 270 178 271
rect 176 270 177 271
rect 175 270 176 271
rect 174 270 175 271
rect 173 270 174 271
rect 172 270 173 271
rect 171 270 172 271
rect 170 270 171 271
rect 169 270 170 271
rect 168 270 169 271
rect 167 270 168 271
rect 166 270 167 271
rect 165 270 166 271
rect 164 270 165 271
rect 163 270 164 271
rect 162 270 163 271
rect 161 270 162 271
rect 160 270 161 271
rect 159 270 160 271
rect 158 270 159 271
rect 157 270 158 271
rect 156 270 157 271
rect 155 270 156 271
rect 154 270 155 271
rect 153 270 154 271
rect 152 270 153 271
rect 151 270 152 271
rect 150 270 151 271
rect 149 270 150 271
rect 148 270 149 271
rect 147 270 148 271
rect 146 270 147 271
rect 145 270 146 271
rect 144 270 145 271
rect 143 270 144 271
rect 142 270 143 271
rect 141 270 142 271
rect 140 270 141 271
rect 139 270 140 271
rect 138 270 139 271
rect 137 270 138 271
rect 136 270 137 271
rect 135 270 136 271
rect 134 270 135 271
rect 133 270 134 271
rect 132 270 133 271
rect 131 270 132 271
rect 130 270 131 271
rect 129 270 130 271
rect 128 270 129 271
rect 127 270 128 271
rect 126 270 127 271
rect 125 270 126 271
rect 111 270 112 271
rect 110 270 111 271
rect 109 270 110 271
rect 108 270 109 271
rect 107 270 108 271
rect 106 270 107 271
rect 105 270 106 271
rect 104 270 105 271
rect 103 270 104 271
rect 102 270 103 271
rect 101 270 102 271
rect 100 270 101 271
rect 99 270 100 271
rect 98 270 99 271
rect 97 270 98 271
rect 96 270 97 271
rect 95 270 96 271
rect 94 270 95 271
rect 93 270 94 271
rect 92 270 93 271
rect 91 270 92 271
rect 90 270 91 271
rect 89 270 90 271
rect 88 270 89 271
rect 87 270 88 271
rect 86 270 87 271
rect 85 270 86 271
rect 84 270 85 271
rect 83 270 84 271
rect 82 270 83 271
rect 81 270 82 271
rect 80 270 81 271
rect 79 270 80 271
rect 78 270 79 271
rect 77 270 78 271
rect 76 270 77 271
rect 59 270 60 271
rect 58 270 59 271
rect 57 270 58 271
rect 56 270 57 271
rect 55 270 56 271
rect 54 270 55 271
rect 53 270 54 271
rect 52 270 53 271
rect 51 270 52 271
rect 50 270 51 271
rect 49 270 50 271
rect 48 270 49 271
rect 47 270 48 271
rect 46 270 47 271
rect 45 270 46 271
rect 44 270 45 271
rect 43 270 44 271
rect 42 270 43 271
rect 41 270 42 271
rect 40 270 41 271
rect 39 270 40 271
rect 38 270 39 271
rect 37 270 38 271
rect 25 270 26 271
rect 24 270 25 271
rect 23 270 24 271
rect 22 270 23 271
rect 21 270 22 271
rect 20 270 21 271
rect 19 270 20 271
rect 18 270 19 271
rect 17 270 18 271
rect 16 270 17 271
rect 15 270 16 271
rect 14 270 15 271
rect 13 270 14 271
rect 12 270 13 271
rect 11 270 12 271
rect 10 270 11 271
rect 9 270 10 271
rect 8 270 9 271
rect 7 270 8 271
rect 6 270 7 271
rect 5 270 6 271
rect 4 270 5 271
rect 3 270 4 271
rect 480 271 481 272
rect 479 271 480 272
rect 478 271 479 272
rect 477 271 478 272
rect 476 271 477 272
rect 475 271 476 272
rect 474 271 475 272
rect 473 271 474 272
rect 472 271 473 272
rect 471 271 472 272
rect 470 271 471 272
rect 469 271 470 272
rect 468 271 469 272
rect 467 271 468 272
rect 466 271 467 272
rect 465 271 466 272
rect 464 271 465 272
rect 463 271 464 272
rect 462 271 463 272
rect 461 271 462 272
rect 460 271 461 272
rect 296 271 297 272
rect 295 271 296 272
rect 294 271 295 272
rect 293 271 294 272
rect 292 271 293 272
rect 291 271 292 272
rect 290 271 291 272
rect 289 271 290 272
rect 288 271 289 272
rect 287 271 288 272
rect 286 271 287 272
rect 285 271 286 272
rect 284 271 285 272
rect 283 271 284 272
rect 282 271 283 272
rect 281 271 282 272
rect 280 271 281 272
rect 279 271 280 272
rect 278 271 279 272
rect 277 271 278 272
rect 276 271 277 272
rect 275 271 276 272
rect 274 271 275 272
rect 273 271 274 272
rect 272 271 273 272
rect 271 271 272 272
rect 270 271 271 272
rect 269 271 270 272
rect 268 271 269 272
rect 267 271 268 272
rect 266 271 267 272
rect 265 271 266 272
rect 264 271 265 272
rect 263 271 264 272
rect 262 271 263 272
rect 261 271 262 272
rect 260 271 261 272
rect 259 271 260 272
rect 258 271 259 272
rect 257 271 258 272
rect 256 271 257 272
rect 255 271 256 272
rect 254 271 255 272
rect 253 271 254 272
rect 252 271 253 272
rect 251 271 252 272
rect 250 271 251 272
rect 249 271 250 272
rect 248 271 249 272
rect 247 271 248 272
rect 246 271 247 272
rect 245 271 246 272
rect 244 271 245 272
rect 243 271 244 272
rect 242 271 243 272
rect 241 271 242 272
rect 240 271 241 272
rect 239 271 240 272
rect 238 271 239 272
rect 237 271 238 272
rect 236 271 237 272
rect 235 271 236 272
rect 234 271 235 272
rect 233 271 234 272
rect 232 271 233 272
rect 231 271 232 272
rect 230 271 231 272
rect 229 271 230 272
rect 228 271 229 272
rect 227 271 228 272
rect 226 271 227 272
rect 225 271 226 272
rect 224 271 225 272
rect 203 271 204 272
rect 202 271 203 272
rect 201 271 202 272
rect 200 271 201 272
rect 199 271 200 272
rect 198 271 199 272
rect 197 271 198 272
rect 196 271 197 272
rect 195 271 196 272
rect 194 271 195 272
rect 193 271 194 272
rect 192 271 193 272
rect 191 271 192 272
rect 190 271 191 272
rect 189 271 190 272
rect 188 271 189 272
rect 187 271 188 272
rect 186 271 187 272
rect 185 271 186 272
rect 184 271 185 272
rect 183 271 184 272
rect 182 271 183 272
rect 181 271 182 272
rect 180 271 181 272
rect 179 271 180 272
rect 178 271 179 272
rect 177 271 178 272
rect 176 271 177 272
rect 175 271 176 272
rect 174 271 175 272
rect 173 271 174 272
rect 172 271 173 272
rect 171 271 172 272
rect 170 271 171 272
rect 169 271 170 272
rect 168 271 169 272
rect 167 271 168 272
rect 166 271 167 272
rect 165 271 166 272
rect 164 271 165 272
rect 163 271 164 272
rect 162 271 163 272
rect 161 271 162 272
rect 160 271 161 272
rect 159 271 160 272
rect 158 271 159 272
rect 157 271 158 272
rect 156 271 157 272
rect 155 271 156 272
rect 154 271 155 272
rect 153 271 154 272
rect 152 271 153 272
rect 151 271 152 272
rect 150 271 151 272
rect 149 271 150 272
rect 148 271 149 272
rect 147 271 148 272
rect 146 271 147 272
rect 145 271 146 272
rect 144 271 145 272
rect 143 271 144 272
rect 142 271 143 272
rect 141 271 142 272
rect 140 271 141 272
rect 139 271 140 272
rect 138 271 139 272
rect 137 271 138 272
rect 136 271 137 272
rect 135 271 136 272
rect 134 271 135 272
rect 133 271 134 272
rect 132 271 133 272
rect 131 271 132 272
rect 130 271 131 272
rect 129 271 130 272
rect 128 271 129 272
rect 127 271 128 272
rect 126 271 127 272
rect 112 271 113 272
rect 111 271 112 272
rect 110 271 111 272
rect 109 271 110 272
rect 108 271 109 272
rect 107 271 108 272
rect 106 271 107 272
rect 105 271 106 272
rect 104 271 105 272
rect 103 271 104 272
rect 102 271 103 272
rect 101 271 102 272
rect 100 271 101 272
rect 99 271 100 272
rect 98 271 99 272
rect 97 271 98 272
rect 96 271 97 272
rect 95 271 96 272
rect 94 271 95 272
rect 93 271 94 272
rect 92 271 93 272
rect 91 271 92 272
rect 90 271 91 272
rect 89 271 90 272
rect 88 271 89 272
rect 87 271 88 272
rect 86 271 87 272
rect 85 271 86 272
rect 84 271 85 272
rect 83 271 84 272
rect 82 271 83 272
rect 81 271 82 272
rect 80 271 81 272
rect 79 271 80 272
rect 78 271 79 272
rect 77 271 78 272
rect 60 271 61 272
rect 59 271 60 272
rect 58 271 59 272
rect 57 271 58 272
rect 56 271 57 272
rect 55 271 56 272
rect 54 271 55 272
rect 53 271 54 272
rect 52 271 53 272
rect 51 271 52 272
rect 50 271 51 272
rect 49 271 50 272
rect 48 271 49 272
rect 47 271 48 272
rect 46 271 47 272
rect 45 271 46 272
rect 44 271 45 272
rect 43 271 44 272
rect 42 271 43 272
rect 41 271 42 272
rect 40 271 41 272
rect 39 271 40 272
rect 38 271 39 272
rect 37 271 38 272
rect 26 271 27 272
rect 25 271 26 272
rect 24 271 25 272
rect 23 271 24 272
rect 22 271 23 272
rect 21 271 22 272
rect 20 271 21 272
rect 19 271 20 272
rect 18 271 19 272
rect 17 271 18 272
rect 16 271 17 272
rect 15 271 16 272
rect 14 271 15 272
rect 13 271 14 272
rect 12 271 13 272
rect 11 271 12 272
rect 10 271 11 272
rect 9 271 10 272
rect 8 271 9 272
rect 7 271 8 272
rect 6 271 7 272
rect 5 271 6 272
rect 4 271 5 272
rect 3 271 4 272
rect 480 272 481 273
rect 479 272 480 273
rect 478 272 479 273
rect 477 272 478 273
rect 476 272 477 273
rect 475 272 476 273
rect 474 272 475 273
rect 473 272 474 273
rect 472 272 473 273
rect 471 272 472 273
rect 470 272 471 273
rect 469 272 470 273
rect 468 272 469 273
rect 467 272 468 273
rect 466 272 467 273
rect 465 272 466 273
rect 464 272 465 273
rect 463 272 464 273
rect 462 272 463 273
rect 461 272 462 273
rect 460 272 461 273
rect 295 272 296 273
rect 294 272 295 273
rect 293 272 294 273
rect 292 272 293 273
rect 291 272 292 273
rect 290 272 291 273
rect 289 272 290 273
rect 288 272 289 273
rect 287 272 288 273
rect 286 272 287 273
rect 285 272 286 273
rect 284 272 285 273
rect 283 272 284 273
rect 282 272 283 273
rect 281 272 282 273
rect 280 272 281 273
rect 279 272 280 273
rect 278 272 279 273
rect 277 272 278 273
rect 276 272 277 273
rect 275 272 276 273
rect 274 272 275 273
rect 273 272 274 273
rect 272 272 273 273
rect 271 272 272 273
rect 270 272 271 273
rect 269 272 270 273
rect 268 272 269 273
rect 267 272 268 273
rect 266 272 267 273
rect 265 272 266 273
rect 264 272 265 273
rect 263 272 264 273
rect 262 272 263 273
rect 261 272 262 273
rect 260 272 261 273
rect 259 272 260 273
rect 258 272 259 273
rect 257 272 258 273
rect 256 272 257 273
rect 255 272 256 273
rect 254 272 255 273
rect 253 272 254 273
rect 252 272 253 273
rect 251 272 252 273
rect 250 272 251 273
rect 249 272 250 273
rect 248 272 249 273
rect 247 272 248 273
rect 246 272 247 273
rect 245 272 246 273
rect 244 272 245 273
rect 243 272 244 273
rect 242 272 243 273
rect 241 272 242 273
rect 240 272 241 273
rect 239 272 240 273
rect 238 272 239 273
rect 237 272 238 273
rect 236 272 237 273
rect 235 272 236 273
rect 234 272 235 273
rect 233 272 234 273
rect 232 272 233 273
rect 231 272 232 273
rect 230 272 231 273
rect 229 272 230 273
rect 228 272 229 273
rect 227 272 228 273
rect 226 272 227 273
rect 225 272 226 273
rect 224 272 225 273
rect 203 272 204 273
rect 202 272 203 273
rect 201 272 202 273
rect 200 272 201 273
rect 199 272 200 273
rect 198 272 199 273
rect 197 272 198 273
rect 196 272 197 273
rect 195 272 196 273
rect 194 272 195 273
rect 193 272 194 273
rect 192 272 193 273
rect 191 272 192 273
rect 190 272 191 273
rect 189 272 190 273
rect 188 272 189 273
rect 187 272 188 273
rect 186 272 187 273
rect 185 272 186 273
rect 184 272 185 273
rect 183 272 184 273
rect 182 272 183 273
rect 181 272 182 273
rect 180 272 181 273
rect 179 272 180 273
rect 178 272 179 273
rect 177 272 178 273
rect 176 272 177 273
rect 175 272 176 273
rect 174 272 175 273
rect 173 272 174 273
rect 172 272 173 273
rect 171 272 172 273
rect 170 272 171 273
rect 169 272 170 273
rect 168 272 169 273
rect 167 272 168 273
rect 166 272 167 273
rect 165 272 166 273
rect 164 272 165 273
rect 163 272 164 273
rect 162 272 163 273
rect 161 272 162 273
rect 160 272 161 273
rect 159 272 160 273
rect 158 272 159 273
rect 157 272 158 273
rect 156 272 157 273
rect 155 272 156 273
rect 154 272 155 273
rect 153 272 154 273
rect 152 272 153 273
rect 151 272 152 273
rect 150 272 151 273
rect 149 272 150 273
rect 148 272 149 273
rect 147 272 148 273
rect 146 272 147 273
rect 145 272 146 273
rect 144 272 145 273
rect 143 272 144 273
rect 142 272 143 273
rect 141 272 142 273
rect 140 272 141 273
rect 139 272 140 273
rect 138 272 139 273
rect 137 272 138 273
rect 136 272 137 273
rect 135 272 136 273
rect 134 272 135 273
rect 133 272 134 273
rect 132 272 133 273
rect 131 272 132 273
rect 130 272 131 273
rect 129 272 130 273
rect 128 272 129 273
rect 127 272 128 273
rect 126 272 127 273
rect 112 272 113 273
rect 111 272 112 273
rect 110 272 111 273
rect 109 272 110 273
rect 108 272 109 273
rect 107 272 108 273
rect 106 272 107 273
rect 105 272 106 273
rect 104 272 105 273
rect 103 272 104 273
rect 102 272 103 273
rect 101 272 102 273
rect 100 272 101 273
rect 99 272 100 273
rect 98 272 99 273
rect 97 272 98 273
rect 96 272 97 273
rect 95 272 96 273
rect 94 272 95 273
rect 93 272 94 273
rect 92 272 93 273
rect 91 272 92 273
rect 90 272 91 273
rect 89 272 90 273
rect 88 272 89 273
rect 87 272 88 273
rect 86 272 87 273
rect 85 272 86 273
rect 84 272 85 273
rect 83 272 84 273
rect 82 272 83 273
rect 81 272 82 273
rect 80 272 81 273
rect 79 272 80 273
rect 78 272 79 273
rect 77 272 78 273
rect 60 272 61 273
rect 59 272 60 273
rect 58 272 59 273
rect 57 272 58 273
rect 56 272 57 273
rect 55 272 56 273
rect 54 272 55 273
rect 53 272 54 273
rect 52 272 53 273
rect 51 272 52 273
rect 50 272 51 273
rect 49 272 50 273
rect 48 272 49 273
rect 47 272 48 273
rect 46 272 47 273
rect 45 272 46 273
rect 44 272 45 273
rect 43 272 44 273
rect 42 272 43 273
rect 41 272 42 273
rect 40 272 41 273
rect 39 272 40 273
rect 38 272 39 273
rect 37 272 38 273
rect 26 272 27 273
rect 25 272 26 273
rect 24 272 25 273
rect 23 272 24 273
rect 22 272 23 273
rect 21 272 22 273
rect 20 272 21 273
rect 19 272 20 273
rect 18 272 19 273
rect 17 272 18 273
rect 16 272 17 273
rect 15 272 16 273
rect 14 272 15 273
rect 13 272 14 273
rect 12 272 13 273
rect 11 272 12 273
rect 10 272 11 273
rect 9 272 10 273
rect 8 272 9 273
rect 7 272 8 273
rect 6 272 7 273
rect 5 272 6 273
rect 4 272 5 273
rect 3 272 4 273
rect 480 273 481 274
rect 479 273 480 274
rect 478 273 479 274
rect 477 273 478 274
rect 476 273 477 274
rect 475 273 476 274
rect 474 273 475 274
rect 473 273 474 274
rect 472 273 473 274
rect 471 273 472 274
rect 470 273 471 274
rect 469 273 470 274
rect 468 273 469 274
rect 467 273 468 274
rect 466 273 467 274
rect 465 273 466 274
rect 464 273 465 274
rect 463 273 464 274
rect 462 273 463 274
rect 461 273 462 274
rect 460 273 461 274
rect 294 273 295 274
rect 293 273 294 274
rect 292 273 293 274
rect 291 273 292 274
rect 290 273 291 274
rect 289 273 290 274
rect 288 273 289 274
rect 287 273 288 274
rect 286 273 287 274
rect 285 273 286 274
rect 284 273 285 274
rect 283 273 284 274
rect 282 273 283 274
rect 281 273 282 274
rect 280 273 281 274
rect 279 273 280 274
rect 278 273 279 274
rect 277 273 278 274
rect 276 273 277 274
rect 275 273 276 274
rect 274 273 275 274
rect 273 273 274 274
rect 272 273 273 274
rect 271 273 272 274
rect 270 273 271 274
rect 269 273 270 274
rect 268 273 269 274
rect 267 273 268 274
rect 266 273 267 274
rect 265 273 266 274
rect 264 273 265 274
rect 263 273 264 274
rect 262 273 263 274
rect 261 273 262 274
rect 260 273 261 274
rect 259 273 260 274
rect 258 273 259 274
rect 257 273 258 274
rect 256 273 257 274
rect 255 273 256 274
rect 254 273 255 274
rect 253 273 254 274
rect 252 273 253 274
rect 251 273 252 274
rect 250 273 251 274
rect 249 273 250 274
rect 248 273 249 274
rect 247 273 248 274
rect 246 273 247 274
rect 245 273 246 274
rect 244 273 245 274
rect 243 273 244 274
rect 242 273 243 274
rect 241 273 242 274
rect 240 273 241 274
rect 239 273 240 274
rect 238 273 239 274
rect 237 273 238 274
rect 236 273 237 274
rect 235 273 236 274
rect 234 273 235 274
rect 233 273 234 274
rect 232 273 233 274
rect 231 273 232 274
rect 230 273 231 274
rect 229 273 230 274
rect 228 273 229 274
rect 227 273 228 274
rect 226 273 227 274
rect 225 273 226 274
rect 224 273 225 274
rect 223 273 224 274
rect 202 273 203 274
rect 201 273 202 274
rect 200 273 201 274
rect 199 273 200 274
rect 198 273 199 274
rect 197 273 198 274
rect 196 273 197 274
rect 195 273 196 274
rect 194 273 195 274
rect 193 273 194 274
rect 192 273 193 274
rect 191 273 192 274
rect 190 273 191 274
rect 189 273 190 274
rect 188 273 189 274
rect 187 273 188 274
rect 186 273 187 274
rect 185 273 186 274
rect 184 273 185 274
rect 183 273 184 274
rect 182 273 183 274
rect 181 273 182 274
rect 180 273 181 274
rect 179 273 180 274
rect 178 273 179 274
rect 177 273 178 274
rect 176 273 177 274
rect 175 273 176 274
rect 174 273 175 274
rect 173 273 174 274
rect 172 273 173 274
rect 171 273 172 274
rect 170 273 171 274
rect 169 273 170 274
rect 168 273 169 274
rect 167 273 168 274
rect 166 273 167 274
rect 165 273 166 274
rect 164 273 165 274
rect 163 273 164 274
rect 162 273 163 274
rect 161 273 162 274
rect 160 273 161 274
rect 159 273 160 274
rect 158 273 159 274
rect 157 273 158 274
rect 156 273 157 274
rect 155 273 156 274
rect 154 273 155 274
rect 153 273 154 274
rect 152 273 153 274
rect 151 273 152 274
rect 150 273 151 274
rect 149 273 150 274
rect 148 273 149 274
rect 147 273 148 274
rect 146 273 147 274
rect 145 273 146 274
rect 144 273 145 274
rect 143 273 144 274
rect 142 273 143 274
rect 141 273 142 274
rect 140 273 141 274
rect 139 273 140 274
rect 138 273 139 274
rect 137 273 138 274
rect 136 273 137 274
rect 135 273 136 274
rect 134 273 135 274
rect 133 273 134 274
rect 132 273 133 274
rect 131 273 132 274
rect 130 273 131 274
rect 129 273 130 274
rect 128 273 129 274
rect 127 273 128 274
rect 126 273 127 274
rect 112 273 113 274
rect 111 273 112 274
rect 110 273 111 274
rect 109 273 110 274
rect 108 273 109 274
rect 107 273 108 274
rect 106 273 107 274
rect 105 273 106 274
rect 104 273 105 274
rect 103 273 104 274
rect 102 273 103 274
rect 101 273 102 274
rect 100 273 101 274
rect 99 273 100 274
rect 98 273 99 274
rect 97 273 98 274
rect 96 273 97 274
rect 95 273 96 274
rect 94 273 95 274
rect 93 273 94 274
rect 92 273 93 274
rect 91 273 92 274
rect 90 273 91 274
rect 89 273 90 274
rect 88 273 89 274
rect 87 273 88 274
rect 86 273 87 274
rect 85 273 86 274
rect 84 273 85 274
rect 83 273 84 274
rect 82 273 83 274
rect 81 273 82 274
rect 80 273 81 274
rect 79 273 80 274
rect 78 273 79 274
rect 61 273 62 274
rect 60 273 61 274
rect 59 273 60 274
rect 58 273 59 274
rect 57 273 58 274
rect 56 273 57 274
rect 55 273 56 274
rect 54 273 55 274
rect 53 273 54 274
rect 52 273 53 274
rect 51 273 52 274
rect 50 273 51 274
rect 49 273 50 274
rect 48 273 49 274
rect 47 273 48 274
rect 46 273 47 274
rect 45 273 46 274
rect 44 273 45 274
rect 43 273 44 274
rect 42 273 43 274
rect 41 273 42 274
rect 40 273 41 274
rect 39 273 40 274
rect 38 273 39 274
rect 37 273 38 274
rect 26 273 27 274
rect 25 273 26 274
rect 24 273 25 274
rect 23 273 24 274
rect 22 273 23 274
rect 21 273 22 274
rect 20 273 21 274
rect 19 273 20 274
rect 18 273 19 274
rect 17 273 18 274
rect 16 273 17 274
rect 15 273 16 274
rect 14 273 15 274
rect 13 273 14 274
rect 12 273 13 274
rect 11 273 12 274
rect 10 273 11 274
rect 9 273 10 274
rect 8 273 9 274
rect 7 273 8 274
rect 6 273 7 274
rect 5 273 6 274
rect 4 273 5 274
rect 3 273 4 274
rect 480 274 481 275
rect 460 274 461 275
rect 439 274 440 275
rect 438 274 439 275
rect 397 274 398 275
rect 396 274 397 275
rect 395 274 396 275
rect 294 274 295 275
rect 293 274 294 275
rect 292 274 293 275
rect 291 274 292 275
rect 290 274 291 275
rect 289 274 290 275
rect 288 274 289 275
rect 287 274 288 275
rect 286 274 287 275
rect 285 274 286 275
rect 284 274 285 275
rect 283 274 284 275
rect 282 274 283 275
rect 281 274 282 275
rect 280 274 281 275
rect 279 274 280 275
rect 278 274 279 275
rect 277 274 278 275
rect 276 274 277 275
rect 275 274 276 275
rect 274 274 275 275
rect 273 274 274 275
rect 272 274 273 275
rect 271 274 272 275
rect 270 274 271 275
rect 269 274 270 275
rect 268 274 269 275
rect 267 274 268 275
rect 266 274 267 275
rect 265 274 266 275
rect 264 274 265 275
rect 263 274 264 275
rect 262 274 263 275
rect 261 274 262 275
rect 260 274 261 275
rect 259 274 260 275
rect 258 274 259 275
rect 257 274 258 275
rect 256 274 257 275
rect 255 274 256 275
rect 254 274 255 275
rect 253 274 254 275
rect 252 274 253 275
rect 251 274 252 275
rect 250 274 251 275
rect 249 274 250 275
rect 248 274 249 275
rect 247 274 248 275
rect 246 274 247 275
rect 245 274 246 275
rect 244 274 245 275
rect 243 274 244 275
rect 242 274 243 275
rect 241 274 242 275
rect 240 274 241 275
rect 239 274 240 275
rect 238 274 239 275
rect 237 274 238 275
rect 236 274 237 275
rect 235 274 236 275
rect 234 274 235 275
rect 233 274 234 275
rect 232 274 233 275
rect 231 274 232 275
rect 230 274 231 275
rect 229 274 230 275
rect 228 274 229 275
rect 227 274 228 275
rect 226 274 227 275
rect 225 274 226 275
rect 224 274 225 275
rect 223 274 224 275
rect 202 274 203 275
rect 201 274 202 275
rect 200 274 201 275
rect 199 274 200 275
rect 198 274 199 275
rect 197 274 198 275
rect 196 274 197 275
rect 195 274 196 275
rect 194 274 195 275
rect 193 274 194 275
rect 192 274 193 275
rect 191 274 192 275
rect 190 274 191 275
rect 189 274 190 275
rect 188 274 189 275
rect 187 274 188 275
rect 186 274 187 275
rect 185 274 186 275
rect 184 274 185 275
rect 183 274 184 275
rect 182 274 183 275
rect 181 274 182 275
rect 180 274 181 275
rect 179 274 180 275
rect 178 274 179 275
rect 177 274 178 275
rect 176 274 177 275
rect 175 274 176 275
rect 174 274 175 275
rect 173 274 174 275
rect 172 274 173 275
rect 171 274 172 275
rect 170 274 171 275
rect 169 274 170 275
rect 168 274 169 275
rect 167 274 168 275
rect 166 274 167 275
rect 165 274 166 275
rect 164 274 165 275
rect 163 274 164 275
rect 162 274 163 275
rect 161 274 162 275
rect 160 274 161 275
rect 159 274 160 275
rect 158 274 159 275
rect 157 274 158 275
rect 156 274 157 275
rect 155 274 156 275
rect 154 274 155 275
rect 153 274 154 275
rect 152 274 153 275
rect 151 274 152 275
rect 150 274 151 275
rect 149 274 150 275
rect 148 274 149 275
rect 147 274 148 275
rect 146 274 147 275
rect 145 274 146 275
rect 144 274 145 275
rect 143 274 144 275
rect 142 274 143 275
rect 141 274 142 275
rect 140 274 141 275
rect 139 274 140 275
rect 138 274 139 275
rect 137 274 138 275
rect 136 274 137 275
rect 135 274 136 275
rect 134 274 135 275
rect 133 274 134 275
rect 132 274 133 275
rect 131 274 132 275
rect 130 274 131 275
rect 129 274 130 275
rect 128 274 129 275
rect 127 274 128 275
rect 112 274 113 275
rect 111 274 112 275
rect 110 274 111 275
rect 109 274 110 275
rect 108 274 109 275
rect 107 274 108 275
rect 106 274 107 275
rect 105 274 106 275
rect 104 274 105 275
rect 103 274 104 275
rect 102 274 103 275
rect 101 274 102 275
rect 100 274 101 275
rect 99 274 100 275
rect 98 274 99 275
rect 97 274 98 275
rect 96 274 97 275
rect 95 274 96 275
rect 94 274 95 275
rect 93 274 94 275
rect 92 274 93 275
rect 91 274 92 275
rect 90 274 91 275
rect 89 274 90 275
rect 88 274 89 275
rect 87 274 88 275
rect 86 274 87 275
rect 85 274 86 275
rect 84 274 85 275
rect 83 274 84 275
rect 82 274 83 275
rect 81 274 82 275
rect 80 274 81 275
rect 79 274 80 275
rect 78 274 79 275
rect 61 274 62 275
rect 60 274 61 275
rect 59 274 60 275
rect 58 274 59 275
rect 57 274 58 275
rect 56 274 57 275
rect 55 274 56 275
rect 54 274 55 275
rect 53 274 54 275
rect 52 274 53 275
rect 51 274 52 275
rect 50 274 51 275
rect 49 274 50 275
rect 48 274 49 275
rect 47 274 48 275
rect 46 274 47 275
rect 45 274 46 275
rect 44 274 45 275
rect 43 274 44 275
rect 42 274 43 275
rect 41 274 42 275
rect 40 274 41 275
rect 39 274 40 275
rect 38 274 39 275
rect 37 274 38 275
rect 26 274 27 275
rect 25 274 26 275
rect 24 274 25 275
rect 23 274 24 275
rect 22 274 23 275
rect 21 274 22 275
rect 20 274 21 275
rect 19 274 20 275
rect 18 274 19 275
rect 17 274 18 275
rect 16 274 17 275
rect 15 274 16 275
rect 14 274 15 275
rect 13 274 14 275
rect 12 274 13 275
rect 11 274 12 275
rect 10 274 11 275
rect 9 274 10 275
rect 8 274 9 275
rect 7 274 8 275
rect 6 274 7 275
rect 5 274 6 275
rect 4 274 5 275
rect 3 274 4 275
rect 480 275 481 276
rect 460 275 461 276
rect 439 275 440 276
rect 438 275 439 276
rect 437 275 438 276
rect 397 275 398 276
rect 396 275 397 276
rect 395 275 396 276
rect 293 275 294 276
rect 292 275 293 276
rect 291 275 292 276
rect 290 275 291 276
rect 289 275 290 276
rect 288 275 289 276
rect 287 275 288 276
rect 286 275 287 276
rect 285 275 286 276
rect 284 275 285 276
rect 283 275 284 276
rect 282 275 283 276
rect 281 275 282 276
rect 280 275 281 276
rect 279 275 280 276
rect 278 275 279 276
rect 277 275 278 276
rect 276 275 277 276
rect 275 275 276 276
rect 274 275 275 276
rect 273 275 274 276
rect 272 275 273 276
rect 271 275 272 276
rect 270 275 271 276
rect 269 275 270 276
rect 268 275 269 276
rect 267 275 268 276
rect 266 275 267 276
rect 265 275 266 276
rect 264 275 265 276
rect 263 275 264 276
rect 262 275 263 276
rect 261 275 262 276
rect 260 275 261 276
rect 259 275 260 276
rect 258 275 259 276
rect 257 275 258 276
rect 256 275 257 276
rect 255 275 256 276
rect 254 275 255 276
rect 253 275 254 276
rect 252 275 253 276
rect 251 275 252 276
rect 250 275 251 276
rect 249 275 250 276
rect 248 275 249 276
rect 247 275 248 276
rect 246 275 247 276
rect 245 275 246 276
rect 244 275 245 276
rect 243 275 244 276
rect 242 275 243 276
rect 241 275 242 276
rect 240 275 241 276
rect 239 275 240 276
rect 238 275 239 276
rect 237 275 238 276
rect 236 275 237 276
rect 235 275 236 276
rect 234 275 235 276
rect 233 275 234 276
rect 232 275 233 276
rect 231 275 232 276
rect 230 275 231 276
rect 229 275 230 276
rect 228 275 229 276
rect 227 275 228 276
rect 226 275 227 276
rect 225 275 226 276
rect 224 275 225 276
rect 223 275 224 276
rect 222 275 223 276
rect 201 275 202 276
rect 200 275 201 276
rect 199 275 200 276
rect 198 275 199 276
rect 197 275 198 276
rect 196 275 197 276
rect 195 275 196 276
rect 194 275 195 276
rect 193 275 194 276
rect 192 275 193 276
rect 191 275 192 276
rect 190 275 191 276
rect 189 275 190 276
rect 188 275 189 276
rect 187 275 188 276
rect 186 275 187 276
rect 185 275 186 276
rect 184 275 185 276
rect 183 275 184 276
rect 182 275 183 276
rect 181 275 182 276
rect 180 275 181 276
rect 179 275 180 276
rect 178 275 179 276
rect 177 275 178 276
rect 176 275 177 276
rect 175 275 176 276
rect 174 275 175 276
rect 173 275 174 276
rect 172 275 173 276
rect 171 275 172 276
rect 170 275 171 276
rect 169 275 170 276
rect 168 275 169 276
rect 167 275 168 276
rect 166 275 167 276
rect 165 275 166 276
rect 164 275 165 276
rect 163 275 164 276
rect 162 275 163 276
rect 161 275 162 276
rect 160 275 161 276
rect 159 275 160 276
rect 158 275 159 276
rect 157 275 158 276
rect 156 275 157 276
rect 155 275 156 276
rect 154 275 155 276
rect 153 275 154 276
rect 152 275 153 276
rect 151 275 152 276
rect 150 275 151 276
rect 149 275 150 276
rect 148 275 149 276
rect 147 275 148 276
rect 146 275 147 276
rect 145 275 146 276
rect 144 275 145 276
rect 143 275 144 276
rect 142 275 143 276
rect 141 275 142 276
rect 140 275 141 276
rect 139 275 140 276
rect 138 275 139 276
rect 137 275 138 276
rect 136 275 137 276
rect 135 275 136 276
rect 134 275 135 276
rect 133 275 134 276
rect 132 275 133 276
rect 131 275 132 276
rect 130 275 131 276
rect 129 275 130 276
rect 128 275 129 276
rect 127 275 128 276
rect 112 275 113 276
rect 111 275 112 276
rect 110 275 111 276
rect 109 275 110 276
rect 108 275 109 276
rect 107 275 108 276
rect 106 275 107 276
rect 105 275 106 276
rect 104 275 105 276
rect 103 275 104 276
rect 102 275 103 276
rect 101 275 102 276
rect 100 275 101 276
rect 99 275 100 276
rect 98 275 99 276
rect 97 275 98 276
rect 96 275 97 276
rect 95 275 96 276
rect 94 275 95 276
rect 93 275 94 276
rect 92 275 93 276
rect 91 275 92 276
rect 90 275 91 276
rect 89 275 90 276
rect 88 275 89 276
rect 87 275 88 276
rect 86 275 87 276
rect 85 275 86 276
rect 84 275 85 276
rect 83 275 84 276
rect 82 275 83 276
rect 81 275 82 276
rect 80 275 81 276
rect 79 275 80 276
rect 62 275 63 276
rect 61 275 62 276
rect 60 275 61 276
rect 59 275 60 276
rect 58 275 59 276
rect 57 275 58 276
rect 56 275 57 276
rect 55 275 56 276
rect 54 275 55 276
rect 53 275 54 276
rect 52 275 53 276
rect 51 275 52 276
rect 50 275 51 276
rect 49 275 50 276
rect 48 275 49 276
rect 47 275 48 276
rect 46 275 47 276
rect 45 275 46 276
rect 44 275 45 276
rect 43 275 44 276
rect 42 275 43 276
rect 41 275 42 276
rect 40 275 41 276
rect 39 275 40 276
rect 38 275 39 276
rect 27 275 28 276
rect 26 275 27 276
rect 25 275 26 276
rect 24 275 25 276
rect 23 275 24 276
rect 22 275 23 276
rect 21 275 22 276
rect 20 275 21 276
rect 19 275 20 276
rect 18 275 19 276
rect 17 275 18 276
rect 16 275 17 276
rect 15 275 16 276
rect 14 275 15 276
rect 13 275 14 276
rect 12 275 13 276
rect 11 275 12 276
rect 10 275 11 276
rect 9 275 10 276
rect 8 275 9 276
rect 7 275 8 276
rect 6 275 7 276
rect 5 275 6 276
rect 4 275 5 276
rect 3 275 4 276
rect 439 276 440 277
rect 438 276 439 277
rect 437 276 438 277
rect 397 276 398 277
rect 396 276 397 277
rect 395 276 396 277
rect 292 276 293 277
rect 291 276 292 277
rect 290 276 291 277
rect 289 276 290 277
rect 288 276 289 277
rect 287 276 288 277
rect 286 276 287 277
rect 285 276 286 277
rect 284 276 285 277
rect 283 276 284 277
rect 282 276 283 277
rect 281 276 282 277
rect 280 276 281 277
rect 279 276 280 277
rect 278 276 279 277
rect 277 276 278 277
rect 276 276 277 277
rect 275 276 276 277
rect 274 276 275 277
rect 273 276 274 277
rect 272 276 273 277
rect 271 276 272 277
rect 270 276 271 277
rect 269 276 270 277
rect 268 276 269 277
rect 267 276 268 277
rect 266 276 267 277
rect 265 276 266 277
rect 264 276 265 277
rect 263 276 264 277
rect 262 276 263 277
rect 261 276 262 277
rect 260 276 261 277
rect 259 276 260 277
rect 258 276 259 277
rect 257 276 258 277
rect 256 276 257 277
rect 255 276 256 277
rect 254 276 255 277
rect 253 276 254 277
rect 252 276 253 277
rect 251 276 252 277
rect 250 276 251 277
rect 249 276 250 277
rect 248 276 249 277
rect 247 276 248 277
rect 246 276 247 277
rect 245 276 246 277
rect 244 276 245 277
rect 243 276 244 277
rect 242 276 243 277
rect 241 276 242 277
rect 240 276 241 277
rect 239 276 240 277
rect 238 276 239 277
rect 237 276 238 277
rect 236 276 237 277
rect 235 276 236 277
rect 234 276 235 277
rect 233 276 234 277
rect 232 276 233 277
rect 231 276 232 277
rect 230 276 231 277
rect 229 276 230 277
rect 228 276 229 277
rect 227 276 228 277
rect 226 276 227 277
rect 225 276 226 277
rect 224 276 225 277
rect 223 276 224 277
rect 222 276 223 277
rect 201 276 202 277
rect 200 276 201 277
rect 199 276 200 277
rect 198 276 199 277
rect 197 276 198 277
rect 196 276 197 277
rect 195 276 196 277
rect 194 276 195 277
rect 193 276 194 277
rect 192 276 193 277
rect 191 276 192 277
rect 190 276 191 277
rect 189 276 190 277
rect 188 276 189 277
rect 187 276 188 277
rect 186 276 187 277
rect 185 276 186 277
rect 184 276 185 277
rect 183 276 184 277
rect 182 276 183 277
rect 181 276 182 277
rect 180 276 181 277
rect 179 276 180 277
rect 178 276 179 277
rect 177 276 178 277
rect 176 276 177 277
rect 175 276 176 277
rect 174 276 175 277
rect 173 276 174 277
rect 172 276 173 277
rect 171 276 172 277
rect 170 276 171 277
rect 169 276 170 277
rect 168 276 169 277
rect 167 276 168 277
rect 166 276 167 277
rect 165 276 166 277
rect 164 276 165 277
rect 163 276 164 277
rect 162 276 163 277
rect 161 276 162 277
rect 160 276 161 277
rect 159 276 160 277
rect 158 276 159 277
rect 157 276 158 277
rect 156 276 157 277
rect 155 276 156 277
rect 154 276 155 277
rect 153 276 154 277
rect 152 276 153 277
rect 151 276 152 277
rect 150 276 151 277
rect 149 276 150 277
rect 148 276 149 277
rect 147 276 148 277
rect 146 276 147 277
rect 145 276 146 277
rect 144 276 145 277
rect 143 276 144 277
rect 142 276 143 277
rect 141 276 142 277
rect 140 276 141 277
rect 139 276 140 277
rect 138 276 139 277
rect 137 276 138 277
rect 136 276 137 277
rect 135 276 136 277
rect 134 276 135 277
rect 133 276 134 277
rect 132 276 133 277
rect 131 276 132 277
rect 130 276 131 277
rect 129 276 130 277
rect 128 276 129 277
rect 127 276 128 277
rect 113 276 114 277
rect 112 276 113 277
rect 111 276 112 277
rect 110 276 111 277
rect 109 276 110 277
rect 108 276 109 277
rect 107 276 108 277
rect 106 276 107 277
rect 105 276 106 277
rect 104 276 105 277
rect 103 276 104 277
rect 102 276 103 277
rect 101 276 102 277
rect 100 276 101 277
rect 99 276 100 277
rect 98 276 99 277
rect 97 276 98 277
rect 96 276 97 277
rect 95 276 96 277
rect 94 276 95 277
rect 93 276 94 277
rect 92 276 93 277
rect 91 276 92 277
rect 90 276 91 277
rect 89 276 90 277
rect 88 276 89 277
rect 87 276 88 277
rect 86 276 87 277
rect 85 276 86 277
rect 84 276 85 277
rect 83 276 84 277
rect 82 276 83 277
rect 81 276 82 277
rect 80 276 81 277
rect 79 276 80 277
rect 62 276 63 277
rect 61 276 62 277
rect 60 276 61 277
rect 59 276 60 277
rect 58 276 59 277
rect 57 276 58 277
rect 56 276 57 277
rect 55 276 56 277
rect 54 276 55 277
rect 53 276 54 277
rect 52 276 53 277
rect 51 276 52 277
rect 50 276 51 277
rect 49 276 50 277
rect 48 276 49 277
rect 47 276 48 277
rect 46 276 47 277
rect 45 276 46 277
rect 44 276 45 277
rect 43 276 44 277
rect 42 276 43 277
rect 41 276 42 277
rect 40 276 41 277
rect 39 276 40 277
rect 38 276 39 277
rect 27 276 28 277
rect 26 276 27 277
rect 25 276 26 277
rect 24 276 25 277
rect 23 276 24 277
rect 22 276 23 277
rect 21 276 22 277
rect 20 276 21 277
rect 19 276 20 277
rect 18 276 19 277
rect 17 276 18 277
rect 16 276 17 277
rect 15 276 16 277
rect 14 276 15 277
rect 13 276 14 277
rect 12 276 13 277
rect 11 276 12 277
rect 10 276 11 277
rect 9 276 10 277
rect 8 276 9 277
rect 7 276 8 277
rect 6 276 7 277
rect 5 276 6 277
rect 4 276 5 277
rect 3 276 4 277
rect 439 277 440 278
rect 438 277 439 278
rect 437 277 438 278
rect 397 277 398 278
rect 396 277 397 278
rect 395 277 396 278
rect 291 277 292 278
rect 290 277 291 278
rect 289 277 290 278
rect 288 277 289 278
rect 287 277 288 278
rect 286 277 287 278
rect 285 277 286 278
rect 284 277 285 278
rect 283 277 284 278
rect 282 277 283 278
rect 281 277 282 278
rect 280 277 281 278
rect 279 277 280 278
rect 278 277 279 278
rect 277 277 278 278
rect 276 277 277 278
rect 275 277 276 278
rect 274 277 275 278
rect 273 277 274 278
rect 272 277 273 278
rect 271 277 272 278
rect 270 277 271 278
rect 269 277 270 278
rect 268 277 269 278
rect 267 277 268 278
rect 266 277 267 278
rect 265 277 266 278
rect 264 277 265 278
rect 263 277 264 278
rect 262 277 263 278
rect 261 277 262 278
rect 260 277 261 278
rect 259 277 260 278
rect 258 277 259 278
rect 257 277 258 278
rect 256 277 257 278
rect 255 277 256 278
rect 254 277 255 278
rect 253 277 254 278
rect 252 277 253 278
rect 251 277 252 278
rect 250 277 251 278
rect 249 277 250 278
rect 248 277 249 278
rect 247 277 248 278
rect 246 277 247 278
rect 245 277 246 278
rect 244 277 245 278
rect 243 277 244 278
rect 242 277 243 278
rect 241 277 242 278
rect 240 277 241 278
rect 239 277 240 278
rect 238 277 239 278
rect 237 277 238 278
rect 236 277 237 278
rect 235 277 236 278
rect 234 277 235 278
rect 233 277 234 278
rect 232 277 233 278
rect 231 277 232 278
rect 230 277 231 278
rect 229 277 230 278
rect 228 277 229 278
rect 227 277 228 278
rect 226 277 227 278
rect 225 277 226 278
rect 224 277 225 278
rect 223 277 224 278
rect 222 277 223 278
rect 200 277 201 278
rect 199 277 200 278
rect 198 277 199 278
rect 197 277 198 278
rect 196 277 197 278
rect 195 277 196 278
rect 194 277 195 278
rect 193 277 194 278
rect 192 277 193 278
rect 191 277 192 278
rect 190 277 191 278
rect 189 277 190 278
rect 188 277 189 278
rect 187 277 188 278
rect 186 277 187 278
rect 185 277 186 278
rect 184 277 185 278
rect 183 277 184 278
rect 182 277 183 278
rect 181 277 182 278
rect 180 277 181 278
rect 179 277 180 278
rect 178 277 179 278
rect 177 277 178 278
rect 176 277 177 278
rect 175 277 176 278
rect 174 277 175 278
rect 173 277 174 278
rect 172 277 173 278
rect 171 277 172 278
rect 170 277 171 278
rect 169 277 170 278
rect 168 277 169 278
rect 167 277 168 278
rect 166 277 167 278
rect 165 277 166 278
rect 164 277 165 278
rect 163 277 164 278
rect 162 277 163 278
rect 161 277 162 278
rect 160 277 161 278
rect 159 277 160 278
rect 158 277 159 278
rect 157 277 158 278
rect 156 277 157 278
rect 155 277 156 278
rect 154 277 155 278
rect 153 277 154 278
rect 152 277 153 278
rect 151 277 152 278
rect 150 277 151 278
rect 149 277 150 278
rect 148 277 149 278
rect 147 277 148 278
rect 146 277 147 278
rect 145 277 146 278
rect 144 277 145 278
rect 143 277 144 278
rect 142 277 143 278
rect 141 277 142 278
rect 140 277 141 278
rect 139 277 140 278
rect 138 277 139 278
rect 137 277 138 278
rect 136 277 137 278
rect 135 277 136 278
rect 134 277 135 278
rect 133 277 134 278
rect 132 277 133 278
rect 131 277 132 278
rect 130 277 131 278
rect 129 277 130 278
rect 128 277 129 278
rect 113 277 114 278
rect 112 277 113 278
rect 111 277 112 278
rect 110 277 111 278
rect 109 277 110 278
rect 108 277 109 278
rect 107 277 108 278
rect 106 277 107 278
rect 105 277 106 278
rect 104 277 105 278
rect 103 277 104 278
rect 102 277 103 278
rect 101 277 102 278
rect 100 277 101 278
rect 99 277 100 278
rect 98 277 99 278
rect 97 277 98 278
rect 96 277 97 278
rect 95 277 96 278
rect 94 277 95 278
rect 93 277 94 278
rect 92 277 93 278
rect 91 277 92 278
rect 90 277 91 278
rect 89 277 90 278
rect 88 277 89 278
rect 87 277 88 278
rect 86 277 87 278
rect 85 277 86 278
rect 84 277 85 278
rect 83 277 84 278
rect 82 277 83 278
rect 81 277 82 278
rect 80 277 81 278
rect 79 277 80 278
rect 62 277 63 278
rect 61 277 62 278
rect 60 277 61 278
rect 59 277 60 278
rect 58 277 59 278
rect 57 277 58 278
rect 56 277 57 278
rect 55 277 56 278
rect 54 277 55 278
rect 53 277 54 278
rect 52 277 53 278
rect 51 277 52 278
rect 50 277 51 278
rect 49 277 50 278
rect 48 277 49 278
rect 47 277 48 278
rect 46 277 47 278
rect 45 277 46 278
rect 44 277 45 278
rect 43 277 44 278
rect 42 277 43 278
rect 41 277 42 278
rect 40 277 41 278
rect 39 277 40 278
rect 38 277 39 278
rect 27 277 28 278
rect 26 277 27 278
rect 25 277 26 278
rect 24 277 25 278
rect 23 277 24 278
rect 22 277 23 278
rect 21 277 22 278
rect 20 277 21 278
rect 19 277 20 278
rect 18 277 19 278
rect 17 277 18 278
rect 16 277 17 278
rect 15 277 16 278
rect 14 277 15 278
rect 13 277 14 278
rect 12 277 13 278
rect 11 277 12 278
rect 10 277 11 278
rect 9 277 10 278
rect 8 277 9 278
rect 7 277 8 278
rect 6 277 7 278
rect 5 277 6 278
rect 4 277 5 278
rect 3 277 4 278
rect 439 278 440 279
rect 438 278 439 279
rect 437 278 438 279
rect 398 278 399 279
rect 397 278 398 279
rect 396 278 397 279
rect 395 278 396 279
rect 290 278 291 279
rect 289 278 290 279
rect 288 278 289 279
rect 287 278 288 279
rect 286 278 287 279
rect 285 278 286 279
rect 284 278 285 279
rect 283 278 284 279
rect 282 278 283 279
rect 281 278 282 279
rect 280 278 281 279
rect 279 278 280 279
rect 278 278 279 279
rect 277 278 278 279
rect 276 278 277 279
rect 275 278 276 279
rect 274 278 275 279
rect 273 278 274 279
rect 272 278 273 279
rect 271 278 272 279
rect 270 278 271 279
rect 269 278 270 279
rect 268 278 269 279
rect 267 278 268 279
rect 266 278 267 279
rect 265 278 266 279
rect 264 278 265 279
rect 263 278 264 279
rect 262 278 263 279
rect 261 278 262 279
rect 260 278 261 279
rect 259 278 260 279
rect 258 278 259 279
rect 257 278 258 279
rect 256 278 257 279
rect 255 278 256 279
rect 254 278 255 279
rect 253 278 254 279
rect 252 278 253 279
rect 251 278 252 279
rect 250 278 251 279
rect 249 278 250 279
rect 248 278 249 279
rect 247 278 248 279
rect 246 278 247 279
rect 245 278 246 279
rect 244 278 245 279
rect 243 278 244 279
rect 242 278 243 279
rect 241 278 242 279
rect 240 278 241 279
rect 239 278 240 279
rect 238 278 239 279
rect 237 278 238 279
rect 236 278 237 279
rect 235 278 236 279
rect 234 278 235 279
rect 233 278 234 279
rect 232 278 233 279
rect 231 278 232 279
rect 230 278 231 279
rect 229 278 230 279
rect 228 278 229 279
rect 227 278 228 279
rect 226 278 227 279
rect 225 278 226 279
rect 224 278 225 279
rect 223 278 224 279
rect 222 278 223 279
rect 221 278 222 279
rect 199 278 200 279
rect 198 278 199 279
rect 197 278 198 279
rect 196 278 197 279
rect 195 278 196 279
rect 194 278 195 279
rect 193 278 194 279
rect 192 278 193 279
rect 191 278 192 279
rect 190 278 191 279
rect 189 278 190 279
rect 188 278 189 279
rect 187 278 188 279
rect 186 278 187 279
rect 185 278 186 279
rect 184 278 185 279
rect 183 278 184 279
rect 182 278 183 279
rect 181 278 182 279
rect 180 278 181 279
rect 179 278 180 279
rect 178 278 179 279
rect 177 278 178 279
rect 176 278 177 279
rect 175 278 176 279
rect 174 278 175 279
rect 173 278 174 279
rect 172 278 173 279
rect 171 278 172 279
rect 170 278 171 279
rect 169 278 170 279
rect 168 278 169 279
rect 167 278 168 279
rect 166 278 167 279
rect 165 278 166 279
rect 164 278 165 279
rect 163 278 164 279
rect 162 278 163 279
rect 161 278 162 279
rect 160 278 161 279
rect 159 278 160 279
rect 158 278 159 279
rect 157 278 158 279
rect 156 278 157 279
rect 155 278 156 279
rect 154 278 155 279
rect 153 278 154 279
rect 152 278 153 279
rect 151 278 152 279
rect 150 278 151 279
rect 149 278 150 279
rect 148 278 149 279
rect 147 278 148 279
rect 146 278 147 279
rect 145 278 146 279
rect 144 278 145 279
rect 143 278 144 279
rect 142 278 143 279
rect 141 278 142 279
rect 140 278 141 279
rect 139 278 140 279
rect 138 278 139 279
rect 137 278 138 279
rect 136 278 137 279
rect 135 278 136 279
rect 134 278 135 279
rect 133 278 134 279
rect 132 278 133 279
rect 131 278 132 279
rect 130 278 131 279
rect 129 278 130 279
rect 128 278 129 279
rect 113 278 114 279
rect 112 278 113 279
rect 111 278 112 279
rect 110 278 111 279
rect 109 278 110 279
rect 108 278 109 279
rect 107 278 108 279
rect 106 278 107 279
rect 105 278 106 279
rect 104 278 105 279
rect 103 278 104 279
rect 102 278 103 279
rect 101 278 102 279
rect 100 278 101 279
rect 99 278 100 279
rect 98 278 99 279
rect 97 278 98 279
rect 96 278 97 279
rect 95 278 96 279
rect 94 278 95 279
rect 93 278 94 279
rect 92 278 93 279
rect 91 278 92 279
rect 90 278 91 279
rect 89 278 90 279
rect 88 278 89 279
rect 87 278 88 279
rect 86 278 87 279
rect 85 278 86 279
rect 84 278 85 279
rect 83 278 84 279
rect 82 278 83 279
rect 81 278 82 279
rect 80 278 81 279
rect 63 278 64 279
rect 62 278 63 279
rect 61 278 62 279
rect 60 278 61 279
rect 59 278 60 279
rect 58 278 59 279
rect 57 278 58 279
rect 56 278 57 279
rect 55 278 56 279
rect 54 278 55 279
rect 53 278 54 279
rect 52 278 53 279
rect 51 278 52 279
rect 50 278 51 279
rect 49 278 50 279
rect 48 278 49 279
rect 47 278 48 279
rect 46 278 47 279
rect 45 278 46 279
rect 44 278 45 279
rect 43 278 44 279
rect 42 278 43 279
rect 41 278 42 279
rect 40 278 41 279
rect 39 278 40 279
rect 38 278 39 279
rect 27 278 28 279
rect 26 278 27 279
rect 25 278 26 279
rect 24 278 25 279
rect 23 278 24 279
rect 22 278 23 279
rect 21 278 22 279
rect 20 278 21 279
rect 19 278 20 279
rect 18 278 19 279
rect 17 278 18 279
rect 16 278 17 279
rect 15 278 16 279
rect 14 278 15 279
rect 13 278 14 279
rect 12 278 13 279
rect 11 278 12 279
rect 10 278 11 279
rect 9 278 10 279
rect 8 278 9 279
rect 7 278 8 279
rect 6 278 7 279
rect 5 278 6 279
rect 4 278 5 279
rect 3 278 4 279
rect 439 279 440 280
rect 438 279 439 280
rect 437 279 438 280
rect 436 279 437 280
rect 435 279 436 280
rect 399 279 400 280
rect 398 279 399 280
rect 397 279 398 280
rect 396 279 397 280
rect 395 279 396 280
rect 290 279 291 280
rect 289 279 290 280
rect 288 279 289 280
rect 287 279 288 280
rect 286 279 287 280
rect 285 279 286 280
rect 284 279 285 280
rect 283 279 284 280
rect 282 279 283 280
rect 281 279 282 280
rect 280 279 281 280
rect 279 279 280 280
rect 278 279 279 280
rect 277 279 278 280
rect 276 279 277 280
rect 275 279 276 280
rect 274 279 275 280
rect 273 279 274 280
rect 272 279 273 280
rect 271 279 272 280
rect 270 279 271 280
rect 269 279 270 280
rect 268 279 269 280
rect 267 279 268 280
rect 266 279 267 280
rect 265 279 266 280
rect 264 279 265 280
rect 263 279 264 280
rect 262 279 263 280
rect 261 279 262 280
rect 260 279 261 280
rect 259 279 260 280
rect 258 279 259 280
rect 257 279 258 280
rect 256 279 257 280
rect 255 279 256 280
rect 254 279 255 280
rect 253 279 254 280
rect 252 279 253 280
rect 251 279 252 280
rect 250 279 251 280
rect 249 279 250 280
rect 248 279 249 280
rect 247 279 248 280
rect 246 279 247 280
rect 245 279 246 280
rect 244 279 245 280
rect 243 279 244 280
rect 242 279 243 280
rect 241 279 242 280
rect 240 279 241 280
rect 239 279 240 280
rect 238 279 239 280
rect 237 279 238 280
rect 236 279 237 280
rect 235 279 236 280
rect 234 279 235 280
rect 233 279 234 280
rect 232 279 233 280
rect 231 279 232 280
rect 230 279 231 280
rect 229 279 230 280
rect 228 279 229 280
rect 227 279 228 280
rect 226 279 227 280
rect 225 279 226 280
rect 224 279 225 280
rect 223 279 224 280
rect 222 279 223 280
rect 221 279 222 280
rect 199 279 200 280
rect 198 279 199 280
rect 197 279 198 280
rect 196 279 197 280
rect 195 279 196 280
rect 194 279 195 280
rect 193 279 194 280
rect 192 279 193 280
rect 191 279 192 280
rect 190 279 191 280
rect 189 279 190 280
rect 188 279 189 280
rect 187 279 188 280
rect 186 279 187 280
rect 185 279 186 280
rect 184 279 185 280
rect 183 279 184 280
rect 182 279 183 280
rect 181 279 182 280
rect 180 279 181 280
rect 179 279 180 280
rect 178 279 179 280
rect 177 279 178 280
rect 176 279 177 280
rect 175 279 176 280
rect 174 279 175 280
rect 173 279 174 280
rect 172 279 173 280
rect 171 279 172 280
rect 170 279 171 280
rect 169 279 170 280
rect 168 279 169 280
rect 167 279 168 280
rect 166 279 167 280
rect 165 279 166 280
rect 164 279 165 280
rect 163 279 164 280
rect 162 279 163 280
rect 161 279 162 280
rect 160 279 161 280
rect 159 279 160 280
rect 158 279 159 280
rect 157 279 158 280
rect 156 279 157 280
rect 155 279 156 280
rect 154 279 155 280
rect 153 279 154 280
rect 152 279 153 280
rect 151 279 152 280
rect 150 279 151 280
rect 149 279 150 280
rect 148 279 149 280
rect 147 279 148 280
rect 146 279 147 280
rect 145 279 146 280
rect 144 279 145 280
rect 143 279 144 280
rect 142 279 143 280
rect 141 279 142 280
rect 140 279 141 280
rect 139 279 140 280
rect 138 279 139 280
rect 137 279 138 280
rect 136 279 137 280
rect 135 279 136 280
rect 134 279 135 280
rect 133 279 134 280
rect 132 279 133 280
rect 131 279 132 280
rect 130 279 131 280
rect 129 279 130 280
rect 114 279 115 280
rect 113 279 114 280
rect 112 279 113 280
rect 111 279 112 280
rect 110 279 111 280
rect 109 279 110 280
rect 108 279 109 280
rect 107 279 108 280
rect 106 279 107 280
rect 105 279 106 280
rect 104 279 105 280
rect 103 279 104 280
rect 102 279 103 280
rect 101 279 102 280
rect 100 279 101 280
rect 99 279 100 280
rect 98 279 99 280
rect 97 279 98 280
rect 96 279 97 280
rect 95 279 96 280
rect 94 279 95 280
rect 93 279 94 280
rect 92 279 93 280
rect 91 279 92 280
rect 90 279 91 280
rect 89 279 90 280
rect 88 279 89 280
rect 87 279 88 280
rect 86 279 87 280
rect 85 279 86 280
rect 84 279 85 280
rect 83 279 84 280
rect 82 279 83 280
rect 81 279 82 280
rect 80 279 81 280
rect 63 279 64 280
rect 62 279 63 280
rect 61 279 62 280
rect 60 279 61 280
rect 59 279 60 280
rect 58 279 59 280
rect 57 279 58 280
rect 56 279 57 280
rect 55 279 56 280
rect 54 279 55 280
rect 53 279 54 280
rect 52 279 53 280
rect 51 279 52 280
rect 50 279 51 280
rect 49 279 50 280
rect 48 279 49 280
rect 47 279 48 280
rect 46 279 47 280
rect 45 279 46 280
rect 44 279 45 280
rect 43 279 44 280
rect 42 279 43 280
rect 41 279 42 280
rect 40 279 41 280
rect 39 279 40 280
rect 38 279 39 280
rect 27 279 28 280
rect 26 279 27 280
rect 25 279 26 280
rect 24 279 25 280
rect 23 279 24 280
rect 22 279 23 280
rect 21 279 22 280
rect 20 279 21 280
rect 19 279 20 280
rect 18 279 19 280
rect 17 279 18 280
rect 16 279 17 280
rect 15 279 16 280
rect 14 279 15 280
rect 13 279 14 280
rect 12 279 13 280
rect 11 279 12 280
rect 10 279 11 280
rect 9 279 10 280
rect 8 279 9 280
rect 7 279 8 280
rect 6 279 7 280
rect 5 279 6 280
rect 4 279 5 280
rect 3 279 4 280
rect 439 280 440 281
rect 438 280 439 281
rect 437 280 438 281
rect 436 280 437 281
rect 435 280 436 281
rect 434 280 435 281
rect 433 280 434 281
rect 432 280 433 281
rect 431 280 432 281
rect 430 280 431 281
rect 429 280 430 281
rect 428 280 429 281
rect 427 280 428 281
rect 426 280 427 281
rect 425 280 426 281
rect 424 280 425 281
rect 423 280 424 281
rect 422 280 423 281
rect 421 280 422 281
rect 420 280 421 281
rect 419 280 420 281
rect 418 280 419 281
rect 417 280 418 281
rect 416 280 417 281
rect 415 280 416 281
rect 414 280 415 281
rect 413 280 414 281
rect 412 280 413 281
rect 411 280 412 281
rect 410 280 411 281
rect 409 280 410 281
rect 408 280 409 281
rect 407 280 408 281
rect 406 280 407 281
rect 405 280 406 281
rect 404 280 405 281
rect 403 280 404 281
rect 402 280 403 281
rect 401 280 402 281
rect 400 280 401 281
rect 399 280 400 281
rect 398 280 399 281
rect 397 280 398 281
rect 396 280 397 281
rect 395 280 396 281
rect 289 280 290 281
rect 288 280 289 281
rect 287 280 288 281
rect 286 280 287 281
rect 285 280 286 281
rect 284 280 285 281
rect 283 280 284 281
rect 282 280 283 281
rect 281 280 282 281
rect 280 280 281 281
rect 279 280 280 281
rect 278 280 279 281
rect 277 280 278 281
rect 276 280 277 281
rect 275 280 276 281
rect 274 280 275 281
rect 273 280 274 281
rect 272 280 273 281
rect 271 280 272 281
rect 270 280 271 281
rect 269 280 270 281
rect 268 280 269 281
rect 267 280 268 281
rect 266 280 267 281
rect 265 280 266 281
rect 264 280 265 281
rect 263 280 264 281
rect 262 280 263 281
rect 261 280 262 281
rect 260 280 261 281
rect 259 280 260 281
rect 258 280 259 281
rect 257 280 258 281
rect 256 280 257 281
rect 255 280 256 281
rect 254 280 255 281
rect 253 280 254 281
rect 252 280 253 281
rect 251 280 252 281
rect 250 280 251 281
rect 249 280 250 281
rect 248 280 249 281
rect 247 280 248 281
rect 246 280 247 281
rect 245 280 246 281
rect 244 280 245 281
rect 243 280 244 281
rect 242 280 243 281
rect 241 280 242 281
rect 240 280 241 281
rect 239 280 240 281
rect 238 280 239 281
rect 237 280 238 281
rect 236 280 237 281
rect 235 280 236 281
rect 234 280 235 281
rect 233 280 234 281
rect 232 280 233 281
rect 231 280 232 281
rect 230 280 231 281
rect 229 280 230 281
rect 228 280 229 281
rect 227 280 228 281
rect 226 280 227 281
rect 225 280 226 281
rect 224 280 225 281
rect 223 280 224 281
rect 222 280 223 281
rect 221 280 222 281
rect 220 280 221 281
rect 198 280 199 281
rect 197 280 198 281
rect 196 280 197 281
rect 195 280 196 281
rect 194 280 195 281
rect 193 280 194 281
rect 192 280 193 281
rect 191 280 192 281
rect 190 280 191 281
rect 189 280 190 281
rect 188 280 189 281
rect 187 280 188 281
rect 186 280 187 281
rect 185 280 186 281
rect 184 280 185 281
rect 183 280 184 281
rect 182 280 183 281
rect 181 280 182 281
rect 180 280 181 281
rect 179 280 180 281
rect 178 280 179 281
rect 177 280 178 281
rect 176 280 177 281
rect 175 280 176 281
rect 174 280 175 281
rect 173 280 174 281
rect 172 280 173 281
rect 171 280 172 281
rect 170 280 171 281
rect 169 280 170 281
rect 168 280 169 281
rect 167 280 168 281
rect 166 280 167 281
rect 165 280 166 281
rect 164 280 165 281
rect 163 280 164 281
rect 162 280 163 281
rect 161 280 162 281
rect 160 280 161 281
rect 159 280 160 281
rect 158 280 159 281
rect 157 280 158 281
rect 156 280 157 281
rect 155 280 156 281
rect 154 280 155 281
rect 153 280 154 281
rect 152 280 153 281
rect 151 280 152 281
rect 150 280 151 281
rect 149 280 150 281
rect 148 280 149 281
rect 147 280 148 281
rect 146 280 147 281
rect 145 280 146 281
rect 144 280 145 281
rect 143 280 144 281
rect 142 280 143 281
rect 141 280 142 281
rect 140 280 141 281
rect 139 280 140 281
rect 138 280 139 281
rect 137 280 138 281
rect 136 280 137 281
rect 135 280 136 281
rect 134 280 135 281
rect 133 280 134 281
rect 132 280 133 281
rect 131 280 132 281
rect 130 280 131 281
rect 129 280 130 281
rect 114 280 115 281
rect 113 280 114 281
rect 112 280 113 281
rect 111 280 112 281
rect 110 280 111 281
rect 109 280 110 281
rect 108 280 109 281
rect 107 280 108 281
rect 106 280 107 281
rect 105 280 106 281
rect 104 280 105 281
rect 103 280 104 281
rect 102 280 103 281
rect 101 280 102 281
rect 100 280 101 281
rect 99 280 100 281
rect 98 280 99 281
rect 97 280 98 281
rect 96 280 97 281
rect 95 280 96 281
rect 94 280 95 281
rect 93 280 94 281
rect 92 280 93 281
rect 91 280 92 281
rect 90 280 91 281
rect 89 280 90 281
rect 88 280 89 281
rect 87 280 88 281
rect 86 280 87 281
rect 85 280 86 281
rect 84 280 85 281
rect 83 280 84 281
rect 82 280 83 281
rect 81 280 82 281
rect 80 280 81 281
rect 64 280 65 281
rect 63 280 64 281
rect 62 280 63 281
rect 61 280 62 281
rect 60 280 61 281
rect 59 280 60 281
rect 58 280 59 281
rect 57 280 58 281
rect 56 280 57 281
rect 55 280 56 281
rect 54 280 55 281
rect 53 280 54 281
rect 52 280 53 281
rect 51 280 52 281
rect 50 280 51 281
rect 49 280 50 281
rect 48 280 49 281
rect 47 280 48 281
rect 46 280 47 281
rect 45 280 46 281
rect 44 280 45 281
rect 43 280 44 281
rect 42 280 43 281
rect 41 280 42 281
rect 40 280 41 281
rect 39 280 40 281
rect 38 280 39 281
rect 28 280 29 281
rect 27 280 28 281
rect 26 280 27 281
rect 25 280 26 281
rect 24 280 25 281
rect 23 280 24 281
rect 22 280 23 281
rect 21 280 22 281
rect 20 280 21 281
rect 19 280 20 281
rect 18 280 19 281
rect 17 280 18 281
rect 16 280 17 281
rect 15 280 16 281
rect 14 280 15 281
rect 13 280 14 281
rect 12 280 13 281
rect 11 280 12 281
rect 10 280 11 281
rect 9 280 10 281
rect 8 280 9 281
rect 7 280 8 281
rect 6 280 7 281
rect 5 280 6 281
rect 4 280 5 281
rect 3 280 4 281
rect 439 281 440 282
rect 438 281 439 282
rect 437 281 438 282
rect 436 281 437 282
rect 435 281 436 282
rect 434 281 435 282
rect 433 281 434 282
rect 432 281 433 282
rect 431 281 432 282
rect 430 281 431 282
rect 429 281 430 282
rect 428 281 429 282
rect 427 281 428 282
rect 426 281 427 282
rect 425 281 426 282
rect 424 281 425 282
rect 423 281 424 282
rect 422 281 423 282
rect 421 281 422 282
rect 420 281 421 282
rect 419 281 420 282
rect 418 281 419 282
rect 417 281 418 282
rect 416 281 417 282
rect 415 281 416 282
rect 414 281 415 282
rect 413 281 414 282
rect 412 281 413 282
rect 411 281 412 282
rect 410 281 411 282
rect 409 281 410 282
rect 408 281 409 282
rect 407 281 408 282
rect 406 281 407 282
rect 405 281 406 282
rect 404 281 405 282
rect 403 281 404 282
rect 402 281 403 282
rect 401 281 402 282
rect 400 281 401 282
rect 399 281 400 282
rect 398 281 399 282
rect 397 281 398 282
rect 396 281 397 282
rect 395 281 396 282
rect 288 281 289 282
rect 287 281 288 282
rect 286 281 287 282
rect 285 281 286 282
rect 284 281 285 282
rect 283 281 284 282
rect 282 281 283 282
rect 281 281 282 282
rect 280 281 281 282
rect 279 281 280 282
rect 278 281 279 282
rect 277 281 278 282
rect 276 281 277 282
rect 275 281 276 282
rect 274 281 275 282
rect 273 281 274 282
rect 272 281 273 282
rect 271 281 272 282
rect 270 281 271 282
rect 269 281 270 282
rect 268 281 269 282
rect 267 281 268 282
rect 266 281 267 282
rect 265 281 266 282
rect 264 281 265 282
rect 263 281 264 282
rect 262 281 263 282
rect 261 281 262 282
rect 260 281 261 282
rect 259 281 260 282
rect 258 281 259 282
rect 257 281 258 282
rect 256 281 257 282
rect 255 281 256 282
rect 254 281 255 282
rect 253 281 254 282
rect 252 281 253 282
rect 251 281 252 282
rect 250 281 251 282
rect 249 281 250 282
rect 248 281 249 282
rect 247 281 248 282
rect 246 281 247 282
rect 245 281 246 282
rect 244 281 245 282
rect 243 281 244 282
rect 242 281 243 282
rect 241 281 242 282
rect 240 281 241 282
rect 239 281 240 282
rect 238 281 239 282
rect 237 281 238 282
rect 236 281 237 282
rect 235 281 236 282
rect 234 281 235 282
rect 233 281 234 282
rect 232 281 233 282
rect 231 281 232 282
rect 230 281 231 282
rect 229 281 230 282
rect 228 281 229 282
rect 227 281 228 282
rect 226 281 227 282
rect 225 281 226 282
rect 224 281 225 282
rect 223 281 224 282
rect 222 281 223 282
rect 221 281 222 282
rect 220 281 221 282
rect 198 281 199 282
rect 197 281 198 282
rect 196 281 197 282
rect 195 281 196 282
rect 194 281 195 282
rect 193 281 194 282
rect 192 281 193 282
rect 191 281 192 282
rect 190 281 191 282
rect 189 281 190 282
rect 188 281 189 282
rect 187 281 188 282
rect 186 281 187 282
rect 185 281 186 282
rect 184 281 185 282
rect 183 281 184 282
rect 182 281 183 282
rect 181 281 182 282
rect 180 281 181 282
rect 179 281 180 282
rect 178 281 179 282
rect 177 281 178 282
rect 176 281 177 282
rect 175 281 176 282
rect 174 281 175 282
rect 173 281 174 282
rect 172 281 173 282
rect 171 281 172 282
rect 170 281 171 282
rect 169 281 170 282
rect 168 281 169 282
rect 167 281 168 282
rect 166 281 167 282
rect 165 281 166 282
rect 164 281 165 282
rect 163 281 164 282
rect 162 281 163 282
rect 161 281 162 282
rect 160 281 161 282
rect 159 281 160 282
rect 158 281 159 282
rect 157 281 158 282
rect 156 281 157 282
rect 155 281 156 282
rect 154 281 155 282
rect 153 281 154 282
rect 152 281 153 282
rect 151 281 152 282
rect 150 281 151 282
rect 149 281 150 282
rect 148 281 149 282
rect 147 281 148 282
rect 146 281 147 282
rect 145 281 146 282
rect 144 281 145 282
rect 143 281 144 282
rect 142 281 143 282
rect 141 281 142 282
rect 140 281 141 282
rect 139 281 140 282
rect 138 281 139 282
rect 137 281 138 282
rect 136 281 137 282
rect 135 281 136 282
rect 134 281 135 282
rect 133 281 134 282
rect 132 281 133 282
rect 131 281 132 282
rect 130 281 131 282
rect 114 281 115 282
rect 113 281 114 282
rect 112 281 113 282
rect 111 281 112 282
rect 110 281 111 282
rect 109 281 110 282
rect 108 281 109 282
rect 107 281 108 282
rect 106 281 107 282
rect 105 281 106 282
rect 104 281 105 282
rect 103 281 104 282
rect 102 281 103 282
rect 101 281 102 282
rect 100 281 101 282
rect 99 281 100 282
rect 98 281 99 282
rect 97 281 98 282
rect 96 281 97 282
rect 95 281 96 282
rect 94 281 95 282
rect 93 281 94 282
rect 92 281 93 282
rect 91 281 92 282
rect 90 281 91 282
rect 89 281 90 282
rect 88 281 89 282
rect 87 281 88 282
rect 86 281 87 282
rect 85 281 86 282
rect 84 281 85 282
rect 83 281 84 282
rect 82 281 83 282
rect 81 281 82 282
rect 80 281 81 282
rect 64 281 65 282
rect 63 281 64 282
rect 62 281 63 282
rect 61 281 62 282
rect 60 281 61 282
rect 59 281 60 282
rect 58 281 59 282
rect 57 281 58 282
rect 56 281 57 282
rect 55 281 56 282
rect 54 281 55 282
rect 53 281 54 282
rect 52 281 53 282
rect 51 281 52 282
rect 50 281 51 282
rect 49 281 50 282
rect 48 281 49 282
rect 47 281 48 282
rect 46 281 47 282
rect 45 281 46 282
rect 44 281 45 282
rect 43 281 44 282
rect 42 281 43 282
rect 41 281 42 282
rect 40 281 41 282
rect 39 281 40 282
rect 38 281 39 282
rect 28 281 29 282
rect 27 281 28 282
rect 26 281 27 282
rect 25 281 26 282
rect 24 281 25 282
rect 23 281 24 282
rect 22 281 23 282
rect 21 281 22 282
rect 20 281 21 282
rect 19 281 20 282
rect 18 281 19 282
rect 17 281 18 282
rect 16 281 17 282
rect 15 281 16 282
rect 14 281 15 282
rect 13 281 14 282
rect 12 281 13 282
rect 11 281 12 282
rect 10 281 11 282
rect 9 281 10 282
rect 8 281 9 282
rect 7 281 8 282
rect 6 281 7 282
rect 5 281 6 282
rect 4 281 5 282
rect 3 281 4 282
rect 439 282 440 283
rect 438 282 439 283
rect 437 282 438 283
rect 436 282 437 283
rect 435 282 436 283
rect 434 282 435 283
rect 433 282 434 283
rect 432 282 433 283
rect 431 282 432 283
rect 430 282 431 283
rect 429 282 430 283
rect 428 282 429 283
rect 427 282 428 283
rect 426 282 427 283
rect 425 282 426 283
rect 424 282 425 283
rect 423 282 424 283
rect 422 282 423 283
rect 421 282 422 283
rect 420 282 421 283
rect 419 282 420 283
rect 418 282 419 283
rect 417 282 418 283
rect 416 282 417 283
rect 415 282 416 283
rect 414 282 415 283
rect 413 282 414 283
rect 412 282 413 283
rect 411 282 412 283
rect 410 282 411 283
rect 409 282 410 283
rect 408 282 409 283
rect 407 282 408 283
rect 406 282 407 283
rect 405 282 406 283
rect 404 282 405 283
rect 403 282 404 283
rect 402 282 403 283
rect 401 282 402 283
rect 400 282 401 283
rect 399 282 400 283
rect 398 282 399 283
rect 397 282 398 283
rect 396 282 397 283
rect 395 282 396 283
rect 287 282 288 283
rect 286 282 287 283
rect 285 282 286 283
rect 284 282 285 283
rect 283 282 284 283
rect 282 282 283 283
rect 281 282 282 283
rect 280 282 281 283
rect 279 282 280 283
rect 278 282 279 283
rect 277 282 278 283
rect 276 282 277 283
rect 275 282 276 283
rect 274 282 275 283
rect 273 282 274 283
rect 272 282 273 283
rect 271 282 272 283
rect 270 282 271 283
rect 269 282 270 283
rect 268 282 269 283
rect 267 282 268 283
rect 266 282 267 283
rect 265 282 266 283
rect 264 282 265 283
rect 263 282 264 283
rect 262 282 263 283
rect 261 282 262 283
rect 260 282 261 283
rect 259 282 260 283
rect 258 282 259 283
rect 257 282 258 283
rect 256 282 257 283
rect 255 282 256 283
rect 254 282 255 283
rect 253 282 254 283
rect 252 282 253 283
rect 251 282 252 283
rect 250 282 251 283
rect 249 282 250 283
rect 248 282 249 283
rect 247 282 248 283
rect 246 282 247 283
rect 245 282 246 283
rect 244 282 245 283
rect 243 282 244 283
rect 242 282 243 283
rect 241 282 242 283
rect 240 282 241 283
rect 239 282 240 283
rect 238 282 239 283
rect 237 282 238 283
rect 236 282 237 283
rect 235 282 236 283
rect 234 282 235 283
rect 233 282 234 283
rect 232 282 233 283
rect 231 282 232 283
rect 230 282 231 283
rect 229 282 230 283
rect 228 282 229 283
rect 227 282 228 283
rect 226 282 227 283
rect 225 282 226 283
rect 224 282 225 283
rect 223 282 224 283
rect 222 282 223 283
rect 221 282 222 283
rect 220 282 221 283
rect 219 282 220 283
rect 197 282 198 283
rect 196 282 197 283
rect 195 282 196 283
rect 194 282 195 283
rect 193 282 194 283
rect 192 282 193 283
rect 191 282 192 283
rect 190 282 191 283
rect 189 282 190 283
rect 188 282 189 283
rect 187 282 188 283
rect 186 282 187 283
rect 185 282 186 283
rect 184 282 185 283
rect 183 282 184 283
rect 182 282 183 283
rect 181 282 182 283
rect 180 282 181 283
rect 179 282 180 283
rect 178 282 179 283
rect 177 282 178 283
rect 176 282 177 283
rect 175 282 176 283
rect 174 282 175 283
rect 173 282 174 283
rect 172 282 173 283
rect 171 282 172 283
rect 170 282 171 283
rect 169 282 170 283
rect 168 282 169 283
rect 167 282 168 283
rect 166 282 167 283
rect 165 282 166 283
rect 164 282 165 283
rect 163 282 164 283
rect 162 282 163 283
rect 161 282 162 283
rect 160 282 161 283
rect 159 282 160 283
rect 158 282 159 283
rect 157 282 158 283
rect 156 282 157 283
rect 155 282 156 283
rect 154 282 155 283
rect 153 282 154 283
rect 152 282 153 283
rect 151 282 152 283
rect 150 282 151 283
rect 149 282 150 283
rect 148 282 149 283
rect 147 282 148 283
rect 146 282 147 283
rect 145 282 146 283
rect 144 282 145 283
rect 143 282 144 283
rect 142 282 143 283
rect 141 282 142 283
rect 140 282 141 283
rect 139 282 140 283
rect 138 282 139 283
rect 137 282 138 283
rect 136 282 137 283
rect 135 282 136 283
rect 134 282 135 283
rect 133 282 134 283
rect 132 282 133 283
rect 131 282 132 283
rect 130 282 131 283
rect 115 282 116 283
rect 114 282 115 283
rect 113 282 114 283
rect 112 282 113 283
rect 111 282 112 283
rect 110 282 111 283
rect 109 282 110 283
rect 108 282 109 283
rect 107 282 108 283
rect 106 282 107 283
rect 105 282 106 283
rect 104 282 105 283
rect 103 282 104 283
rect 102 282 103 283
rect 101 282 102 283
rect 100 282 101 283
rect 99 282 100 283
rect 98 282 99 283
rect 97 282 98 283
rect 96 282 97 283
rect 95 282 96 283
rect 94 282 95 283
rect 93 282 94 283
rect 92 282 93 283
rect 91 282 92 283
rect 90 282 91 283
rect 89 282 90 283
rect 88 282 89 283
rect 87 282 88 283
rect 86 282 87 283
rect 85 282 86 283
rect 84 282 85 283
rect 83 282 84 283
rect 82 282 83 283
rect 81 282 82 283
rect 64 282 65 283
rect 63 282 64 283
rect 62 282 63 283
rect 61 282 62 283
rect 60 282 61 283
rect 59 282 60 283
rect 58 282 59 283
rect 57 282 58 283
rect 56 282 57 283
rect 55 282 56 283
rect 54 282 55 283
rect 53 282 54 283
rect 52 282 53 283
rect 51 282 52 283
rect 50 282 51 283
rect 49 282 50 283
rect 48 282 49 283
rect 47 282 48 283
rect 46 282 47 283
rect 45 282 46 283
rect 44 282 45 283
rect 43 282 44 283
rect 42 282 43 283
rect 41 282 42 283
rect 40 282 41 283
rect 39 282 40 283
rect 38 282 39 283
rect 28 282 29 283
rect 27 282 28 283
rect 26 282 27 283
rect 25 282 26 283
rect 24 282 25 283
rect 23 282 24 283
rect 22 282 23 283
rect 21 282 22 283
rect 20 282 21 283
rect 19 282 20 283
rect 18 282 19 283
rect 17 282 18 283
rect 16 282 17 283
rect 15 282 16 283
rect 14 282 15 283
rect 13 282 14 283
rect 12 282 13 283
rect 11 282 12 283
rect 10 282 11 283
rect 9 282 10 283
rect 8 282 9 283
rect 7 282 8 283
rect 6 282 7 283
rect 5 282 6 283
rect 4 282 5 283
rect 3 282 4 283
rect 439 283 440 284
rect 438 283 439 284
rect 437 283 438 284
rect 436 283 437 284
rect 435 283 436 284
rect 434 283 435 284
rect 433 283 434 284
rect 432 283 433 284
rect 431 283 432 284
rect 430 283 431 284
rect 429 283 430 284
rect 428 283 429 284
rect 427 283 428 284
rect 426 283 427 284
rect 425 283 426 284
rect 424 283 425 284
rect 423 283 424 284
rect 422 283 423 284
rect 421 283 422 284
rect 420 283 421 284
rect 419 283 420 284
rect 418 283 419 284
rect 417 283 418 284
rect 416 283 417 284
rect 415 283 416 284
rect 414 283 415 284
rect 413 283 414 284
rect 412 283 413 284
rect 411 283 412 284
rect 410 283 411 284
rect 409 283 410 284
rect 408 283 409 284
rect 407 283 408 284
rect 406 283 407 284
rect 405 283 406 284
rect 404 283 405 284
rect 403 283 404 284
rect 402 283 403 284
rect 401 283 402 284
rect 400 283 401 284
rect 399 283 400 284
rect 398 283 399 284
rect 397 283 398 284
rect 396 283 397 284
rect 395 283 396 284
rect 286 283 287 284
rect 285 283 286 284
rect 284 283 285 284
rect 283 283 284 284
rect 282 283 283 284
rect 281 283 282 284
rect 280 283 281 284
rect 279 283 280 284
rect 278 283 279 284
rect 277 283 278 284
rect 276 283 277 284
rect 275 283 276 284
rect 274 283 275 284
rect 273 283 274 284
rect 272 283 273 284
rect 271 283 272 284
rect 270 283 271 284
rect 269 283 270 284
rect 268 283 269 284
rect 267 283 268 284
rect 266 283 267 284
rect 265 283 266 284
rect 264 283 265 284
rect 263 283 264 284
rect 262 283 263 284
rect 261 283 262 284
rect 260 283 261 284
rect 259 283 260 284
rect 258 283 259 284
rect 257 283 258 284
rect 256 283 257 284
rect 255 283 256 284
rect 254 283 255 284
rect 253 283 254 284
rect 252 283 253 284
rect 251 283 252 284
rect 250 283 251 284
rect 249 283 250 284
rect 248 283 249 284
rect 247 283 248 284
rect 246 283 247 284
rect 245 283 246 284
rect 244 283 245 284
rect 243 283 244 284
rect 242 283 243 284
rect 241 283 242 284
rect 240 283 241 284
rect 239 283 240 284
rect 238 283 239 284
rect 237 283 238 284
rect 236 283 237 284
rect 235 283 236 284
rect 234 283 235 284
rect 233 283 234 284
rect 232 283 233 284
rect 231 283 232 284
rect 230 283 231 284
rect 229 283 230 284
rect 228 283 229 284
rect 227 283 228 284
rect 226 283 227 284
rect 225 283 226 284
rect 224 283 225 284
rect 223 283 224 284
rect 222 283 223 284
rect 221 283 222 284
rect 220 283 221 284
rect 219 283 220 284
rect 196 283 197 284
rect 195 283 196 284
rect 194 283 195 284
rect 193 283 194 284
rect 192 283 193 284
rect 191 283 192 284
rect 190 283 191 284
rect 189 283 190 284
rect 188 283 189 284
rect 187 283 188 284
rect 186 283 187 284
rect 185 283 186 284
rect 184 283 185 284
rect 183 283 184 284
rect 182 283 183 284
rect 181 283 182 284
rect 180 283 181 284
rect 179 283 180 284
rect 178 283 179 284
rect 177 283 178 284
rect 176 283 177 284
rect 175 283 176 284
rect 174 283 175 284
rect 173 283 174 284
rect 172 283 173 284
rect 171 283 172 284
rect 170 283 171 284
rect 169 283 170 284
rect 168 283 169 284
rect 167 283 168 284
rect 166 283 167 284
rect 165 283 166 284
rect 164 283 165 284
rect 163 283 164 284
rect 162 283 163 284
rect 161 283 162 284
rect 160 283 161 284
rect 159 283 160 284
rect 158 283 159 284
rect 157 283 158 284
rect 156 283 157 284
rect 155 283 156 284
rect 154 283 155 284
rect 153 283 154 284
rect 152 283 153 284
rect 151 283 152 284
rect 150 283 151 284
rect 149 283 150 284
rect 148 283 149 284
rect 147 283 148 284
rect 146 283 147 284
rect 145 283 146 284
rect 144 283 145 284
rect 143 283 144 284
rect 142 283 143 284
rect 141 283 142 284
rect 140 283 141 284
rect 139 283 140 284
rect 138 283 139 284
rect 137 283 138 284
rect 136 283 137 284
rect 135 283 136 284
rect 134 283 135 284
rect 133 283 134 284
rect 132 283 133 284
rect 131 283 132 284
rect 115 283 116 284
rect 114 283 115 284
rect 113 283 114 284
rect 112 283 113 284
rect 111 283 112 284
rect 110 283 111 284
rect 109 283 110 284
rect 108 283 109 284
rect 107 283 108 284
rect 106 283 107 284
rect 105 283 106 284
rect 104 283 105 284
rect 103 283 104 284
rect 102 283 103 284
rect 101 283 102 284
rect 100 283 101 284
rect 99 283 100 284
rect 98 283 99 284
rect 97 283 98 284
rect 96 283 97 284
rect 95 283 96 284
rect 94 283 95 284
rect 93 283 94 284
rect 92 283 93 284
rect 91 283 92 284
rect 90 283 91 284
rect 89 283 90 284
rect 88 283 89 284
rect 87 283 88 284
rect 86 283 87 284
rect 85 283 86 284
rect 84 283 85 284
rect 83 283 84 284
rect 82 283 83 284
rect 81 283 82 284
rect 65 283 66 284
rect 64 283 65 284
rect 63 283 64 284
rect 62 283 63 284
rect 61 283 62 284
rect 60 283 61 284
rect 59 283 60 284
rect 58 283 59 284
rect 57 283 58 284
rect 56 283 57 284
rect 55 283 56 284
rect 54 283 55 284
rect 53 283 54 284
rect 52 283 53 284
rect 51 283 52 284
rect 50 283 51 284
rect 49 283 50 284
rect 48 283 49 284
rect 47 283 48 284
rect 46 283 47 284
rect 45 283 46 284
rect 44 283 45 284
rect 43 283 44 284
rect 42 283 43 284
rect 41 283 42 284
rect 40 283 41 284
rect 39 283 40 284
rect 38 283 39 284
rect 28 283 29 284
rect 27 283 28 284
rect 26 283 27 284
rect 25 283 26 284
rect 24 283 25 284
rect 23 283 24 284
rect 22 283 23 284
rect 21 283 22 284
rect 20 283 21 284
rect 19 283 20 284
rect 18 283 19 284
rect 17 283 18 284
rect 16 283 17 284
rect 15 283 16 284
rect 14 283 15 284
rect 13 283 14 284
rect 12 283 13 284
rect 11 283 12 284
rect 10 283 11 284
rect 9 283 10 284
rect 8 283 9 284
rect 7 283 8 284
rect 6 283 7 284
rect 5 283 6 284
rect 4 283 5 284
rect 3 283 4 284
rect 464 284 465 285
rect 439 284 440 285
rect 438 284 439 285
rect 437 284 438 285
rect 436 284 437 285
rect 435 284 436 285
rect 434 284 435 285
rect 433 284 434 285
rect 432 284 433 285
rect 431 284 432 285
rect 430 284 431 285
rect 429 284 430 285
rect 428 284 429 285
rect 427 284 428 285
rect 426 284 427 285
rect 425 284 426 285
rect 424 284 425 285
rect 423 284 424 285
rect 422 284 423 285
rect 421 284 422 285
rect 420 284 421 285
rect 419 284 420 285
rect 418 284 419 285
rect 417 284 418 285
rect 416 284 417 285
rect 415 284 416 285
rect 414 284 415 285
rect 413 284 414 285
rect 412 284 413 285
rect 411 284 412 285
rect 410 284 411 285
rect 409 284 410 285
rect 408 284 409 285
rect 407 284 408 285
rect 406 284 407 285
rect 405 284 406 285
rect 404 284 405 285
rect 403 284 404 285
rect 402 284 403 285
rect 401 284 402 285
rect 400 284 401 285
rect 399 284 400 285
rect 398 284 399 285
rect 397 284 398 285
rect 396 284 397 285
rect 395 284 396 285
rect 285 284 286 285
rect 284 284 285 285
rect 283 284 284 285
rect 282 284 283 285
rect 281 284 282 285
rect 280 284 281 285
rect 279 284 280 285
rect 278 284 279 285
rect 277 284 278 285
rect 276 284 277 285
rect 275 284 276 285
rect 274 284 275 285
rect 273 284 274 285
rect 272 284 273 285
rect 271 284 272 285
rect 270 284 271 285
rect 269 284 270 285
rect 268 284 269 285
rect 267 284 268 285
rect 266 284 267 285
rect 265 284 266 285
rect 264 284 265 285
rect 263 284 264 285
rect 262 284 263 285
rect 261 284 262 285
rect 260 284 261 285
rect 259 284 260 285
rect 258 284 259 285
rect 257 284 258 285
rect 256 284 257 285
rect 255 284 256 285
rect 254 284 255 285
rect 253 284 254 285
rect 252 284 253 285
rect 251 284 252 285
rect 250 284 251 285
rect 249 284 250 285
rect 248 284 249 285
rect 247 284 248 285
rect 246 284 247 285
rect 245 284 246 285
rect 244 284 245 285
rect 243 284 244 285
rect 242 284 243 285
rect 241 284 242 285
rect 240 284 241 285
rect 239 284 240 285
rect 238 284 239 285
rect 237 284 238 285
rect 236 284 237 285
rect 235 284 236 285
rect 234 284 235 285
rect 233 284 234 285
rect 232 284 233 285
rect 231 284 232 285
rect 230 284 231 285
rect 229 284 230 285
rect 228 284 229 285
rect 227 284 228 285
rect 226 284 227 285
rect 225 284 226 285
rect 224 284 225 285
rect 223 284 224 285
rect 222 284 223 285
rect 221 284 222 285
rect 220 284 221 285
rect 219 284 220 285
rect 218 284 219 285
rect 196 284 197 285
rect 195 284 196 285
rect 194 284 195 285
rect 193 284 194 285
rect 192 284 193 285
rect 191 284 192 285
rect 190 284 191 285
rect 189 284 190 285
rect 188 284 189 285
rect 187 284 188 285
rect 186 284 187 285
rect 185 284 186 285
rect 184 284 185 285
rect 183 284 184 285
rect 182 284 183 285
rect 181 284 182 285
rect 180 284 181 285
rect 179 284 180 285
rect 178 284 179 285
rect 177 284 178 285
rect 176 284 177 285
rect 175 284 176 285
rect 174 284 175 285
rect 173 284 174 285
rect 172 284 173 285
rect 171 284 172 285
rect 170 284 171 285
rect 169 284 170 285
rect 168 284 169 285
rect 167 284 168 285
rect 166 284 167 285
rect 165 284 166 285
rect 164 284 165 285
rect 163 284 164 285
rect 162 284 163 285
rect 161 284 162 285
rect 160 284 161 285
rect 159 284 160 285
rect 158 284 159 285
rect 157 284 158 285
rect 156 284 157 285
rect 155 284 156 285
rect 154 284 155 285
rect 153 284 154 285
rect 152 284 153 285
rect 151 284 152 285
rect 150 284 151 285
rect 149 284 150 285
rect 148 284 149 285
rect 147 284 148 285
rect 146 284 147 285
rect 145 284 146 285
rect 144 284 145 285
rect 143 284 144 285
rect 142 284 143 285
rect 141 284 142 285
rect 140 284 141 285
rect 139 284 140 285
rect 138 284 139 285
rect 137 284 138 285
rect 136 284 137 285
rect 135 284 136 285
rect 134 284 135 285
rect 133 284 134 285
rect 132 284 133 285
rect 131 284 132 285
rect 115 284 116 285
rect 114 284 115 285
rect 113 284 114 285
rect 112 284 113 285
rect 111 284 112 285
rect 110 284 111 285
rect 109 284 110 285
rect 108 284 109 285
rect 107 284 108 285
rect 106 284 107 285
rect 105 284 106 285
rect 104 284 105 285
rect 103 284 104 285
rect 102 284 103 285
rect 101 284 102 285
rect 100 284 101 285
rect 99 284 100 285
rect 98 284 99 285
rect 97 284 98 285
rect 96 284 97 285
rect 95 284 96 285
rect 94 284 95 285
rect 93 284 94 285
rect 92 284 93 285
rect 91 284 92 285
rect 90 284 91 285
rect 89 284 90 285
rect 88 284 89 285
rect 87 284 88 285
rect 86 284 87 285
rect 85 284 86 285
rect 84 284 85 285
rect 83 284 84 285
rect 82 284 83 285
rect 81 284 82 285
rect 65 284 66 285
rect 64 284 65 285
rect 63 284 64 285
rect 62 284 63 285
rect 61 284 62 285
rect 60 284 61 285
rect 59 284 60 285
rect 58 284 59 285
rect 57 284 58 285
rect 56 284 57 285
rect 55 284 56 285
rect 54 284 55 285
rect 53 284 54 285
rect 52 284 53 285
rect 51 284 52 285
rect 50 284 51 285
rect 49 284 50 285
rect 48 284 49 285
rect 47 284 48 285
rect 46 284 47 285
rect 45 284 46 285
rect 44 284 45 285
rect 43 284 44 285
rect 42 284 43 285
rect 41 284 42 285
rect 40 284 41 285
rect 39 284 40 285
rect 38 284 39 285
rect 28 284 29 285
rect 27 284 28 285
rect 26 284 27 285
rect 25 284 26 285
rect 24 284 25 285
rect 23 284 24 285
rect 22 284 23 285
rect 21 284 22 285
rect 20 284 21 285
rect 19 284 20 285
rect 18 284 19 285
rect 17 284 18 285
rect 16 284 17 285
rect 15 284 16 285
rect 14 284 15 285
rect 13 284 14 285
rect 12 284 13 285
rect 11 284 12 285
rect 10 284 11 285
rect 9 284 10 285
rect 8 284 9 285
rect 7 284 8 285
rect 6 284 7 285
rect 5 284 6 285
rect 4 284 5 285
rect 3 284 4 285
rect 465 285 466 286
rect 464 285 465 286
rect 463 285 464 286
rect 462 285 463 286
rect 461 285 462 286
rect 460 285 461 286
rect 459 285 460 286
rect 439 285 440 286
rect 438 285 439 286
rect 437 285 438 286
rect 436 285 437 286
rect 435 285 436 286
rect 434 285 435 286
rect 433 285 434 286
rect 432 285 433 286
rect 431 285 432 286
rect 430 285 431 286
rect 429 285 430 286
rect 428 285 429 286
rect 427 285 428 286
rect 426 285 427 286
rect 425 285 426 286
rect 424 285 425 286
rect 423 285 424 286
rect 422 285 423 286
rect 421 285 422 286
rect 420 285 421 286
rect 419 285 420 286
rect 418 285 419 286
rect 417 285 418 286
rect 416 285 417 286
rect 415 285 416 286
rect 414 285 415 286
rect 413 285 414 286
rect 412 285 413 286
rect 411 285 412 286
rect 410 285 411 286
rect 409 285 410 286
rect 408 285 409 286
rect 407 285 408 286
rect 406 285 407 286
rect 405 285 406 286
rect 404 285 405 286
rect 403 285 404 286
rect 402 285 403 286
rect 401 285 402 286
rect 400 285 401 286
rect 399 285 400 286
rect 398 285 399 286
rect 397 285 398 286
rect 396 285 397 286
rect 395 285 396 286
rect 284 285 285 286
rect 283 285 284 286
rect 282 285 283 286
rect 281 285 282 286
rect 280 285 281 286
rect 279 285 280 286
rect 278 285 279 286
rect 277 285 278 286
rect 276 285 277 286
rect 275 285 276 286
rect 274 285 275 286
rect 273 285 274 286
rect 272 285 273 286
rect 271 285 272 286
rect 270 285 271 286
rect 269 285 270 286
rect 268 285 269 286
rect 267 285 268 286
rect 266 285 267 286
rect 265 285 266 286
rect 264 285 265 286
rect 263 285 264 286
rect 262 285 263 286
rect 261 285 262 286
rect 260 285 261 286
rect 259 285 260 286
rect 258 285 259 286
rect 257 285 258 286
rect 256 285 257 286
rect 255 285 256 286
rect 254 285 255 286
rect 253 285 254 286
rect 252 285 253 286
rect 251 285 252 286
rect 250 285 251 286
rect 249 285 250 286
rect 248 285 249 286
rect 247 285 248 286
rect 246 285 247 286
rect 245 285 246 286
rect 244 285 245 286
rect 243 285 244 286
rect 242 285 243 286
rect 241 285 242 286
rect 240 285 241 286
rect 239 285 240 286
rect 238 285 239 286
rect 237 285 238 286
rect 236 285 237 286
rect 235 285 236 286
rect 234 285 235 286
rect 233 285 234 286
rect 232 285 233 286
rect 231 285 232 286
rect 230 285 231 286
rect 229 285 230 286
rect 228 285 229 286
rect 227 285 228 286
rect 226 285 227 286
rect 225 285 226 286
rect 224 285 225 286
rect 223 285 224 286
rect 222 285 223 286
rect 221 285 222 286
rect 220 285 221 286
rect 219 285 220 286
rect 218 285 219 286
rect 217 285 218 286
rect 195 285 196 286
rect 194 285 195 286
rect 193 285 194 286
rect 192 285 193 286
rect 191 285 192 286
rect 190 285 191 286
rect 189 285 190 286
rect 188 285 189 286
rect 187 285 188 286
rect 186 285 187 286
rect 185 285 186 286
rect 184 285 185 286
rect 183 285 184 286
rect 182 285 183 286
rect 181 285 182 286
rect 180 285 181 286
rect 179 285 180 286
rect 178 285 179 286
rect 177 285 178 286
rect 176 285 177 286
rect 175 285 176 286
rect 174 285 175 286
rect 173 285 174 286
rect 172 285 173 286
rect 171 285 172 286
rect 170 285 171 286
rect 169 285 170 286
rect 168 285 169 286
rect 167 285 168 286
rect 166 285 167 286
rect 165 285 166 286
rect 164 285 165 286
rect 163 285 164 286
rect 162 285 163 286
rect 161 285 162 286
rect 160 285 161 286
rect 159 285 160 286
rect 158 285 159 286
rect 157 285 158 286
rect 156 285 157 286
rect 155 285 156 286
rect 154 285 155 286
rect 153 285 154 286
rect 152 285 153 286
rect 151 285 152 286
rect 150 285 151 286
rect 149 285 150 286
rect 148 285 149 286
rect 147 285 148 286
rect 146 285 147 286
rect 145 285 146 286
rect 144 285 145 286
rect 143 285 144 286
rect 142 285 143 286
rect 141 285 142 286
rect 140 285 141 286
rect 139 285 140 286
rect 138 285 139 286
rect 137 285 138 286
rect 136 285 137 286
rect 135 285 136 286
rect 134 285 135 286
rect 133 285 134 286
rect 132 285 133 286
rect 116 285 117 286
rect 115 285 116 286
rect 114 285 115 286
rect 113 285 114 286
rect 112 285 113 286
rect 111 285 112 286
rect 110 285 111 286
rect 109 285 110 286
rect 108 285 109 286
rect 107 285 108 286
rect 106 285 107 286
rect 105 285 106 286
rect 104 285 105 286
rect 103 285 104 286
rect 102 285 103 286
rect 101 285 102 286
rect 100 285 101 286
rect 99 285 100 286
rect 98 285 99 286
rect 97 285 98 286
rect 96 285 97 286
rect 95 285 96 286
rect 94 285 95 286
rect 93 285 94 286
rect 92 285 93 286
rect 91 285 92 286
rect 90 285 91 286
rect 89 285 90 286
rect 88 285 89 286
rect 87 285 88 286
rect 86 285 87 286
rect 85 285 86 286
rect 84 285 85 286
rect 83 285 84 286
rect 82 285 83 286
rect 66 285 67 286
rect 65 285 66 286
rect 64 285 65 286
rect 63 285 64 286
rect 62 285 63 286
rect 61 285 62 286
rect 60 285 61 286
rect 59 285 60 286
rect 58 285 59 286
rect 57 285 58 286
rect 56 285 57 286
rect 55 285 56 286
rect 54 285 55 286
rect 53 285 54 286
rect 52 285 53 286
rect 51 285 52 286
rect 50 285 51 286
rect 49 285 50 286
rect 48 285 49 286
rect 47 285 48 286
rect 46 285 47 286
rect 45 285 46 286
rect 44 285 45 286
rect 43 285 44 286
rect 42 285 43 286
rect 41 285 42 286
rect 40 285 41 286
rect 39 285 40 286
rect 38 285 39 286
rect 28 285 29 286
rect 27 285 28 286
rect 26 285 27 286
rect 25 285 26 286
rect 24 285 25 286
rect 23 285 24 286
rect 22 285 23 286
rect 21 285 22 286
rect 20 285 21 286
rect 19 285 20 286
rect 18 285 19 286
rect 17 285 18 286
rect 16 285 17 286
rect 15 285 16 286
rect 14 285 15 286
rect 13 285 14 286
rect 12 285 13 286
rect 11 285 12 286
rect 10 285 11 286
rect 9 285 10 286
rect 8 285 9 286
rect 7 285 8 286
rect 6 285 7 286
rect 5 285 6 286
rect 4 285 5 286
rect 3 285 4 286
rect 462 286 463 287
rect 461 286 462 287
rect 460 286 461 287
rect 459 286 460 287
rect 439 286 440 287
rect 438 286 439 287
rect 437 286 438 287
rect 436 286 437 287
rect 435 286 436 287
rect 434 286 435 287
rect 433 286 434 287
rect 432 286 433 287
rect 431 286 432 287
rect 430 286 431 287
rect 429 286 430 287
rect 428 286 429 287
rect 427 286 428 287
rect 426 286 427 287
rect 425 286 426 287
rect 424 286 425 287
rect 423 286 424 287
rect 422 286 423 287
rect 421 286 422 287
rect 420 286 421 287
rect 419 286 420 287
rect 418 286 419 287
rect 417 286 418 287
rect 416 286 417 287
rect 415 286 416 287
rect 414 286 415 287
rect 413 286 414 287
rect 412 286 413 287
rect 411 286 412 287
rect 410 286 411 287
rect 409 286 410 287
rect 408 286 409 287
rect 407 286 408 287
rect 406 286 407 287
rect 405 286 406 287
rect 404 286 405 287
rect 403 286 404 287
rect 402 286 403 287
rect 401 286 402 287
rect 400 286 401 287
rect 399 286 400 287
rect 398 286 399 287
rect 397 286 398 287
rect 396 286 397 287
rect 395 286 396 287
rect 284 286 285 287
rect 283 286 284 287
rect 282 286 283 287
rect 281 286 282 287
rect 280 286 281 287
rect 279 286 280 287
rect 278 286 279 287
rect 277 286 278 287
rect 276 286 277 287
rect 275 286 276 287
rect 274 286 275 287
rect 273 286 274 287
rect 272 286 273 287
rect 271 286 272 287
rect 270 286 271 287
rect 269 286 270 287
rect 268 286 269 287
rect 267 286 268 287
rect 266 286 267 287
rect 265 286 266 287
rect 264 286 265 287
rect 263 286 264 287
rect 262 286 263 287
rect 261 286 262 287
rect 260 286 261 287
rect 259 286 260 287
rect 258 286 259 287
rect 257 286 258 287
rect 256 286 257 287
rect 255 286 256 287
rect 254 286 255 287
rect 253 286 254 287
rect 252 286 253 287
rect 251 286 252 287
rect 250 286 251 287
rect 249 286 250 287
rect 248 286 249 287
rect 247 286 248 287
rect 246 286 247 287
rect 245 286 246 287
rect 244 286 245 287
rect 243 286 244 287
rect 242 286 243 287
rect 241 286 242 287
rect 240 286 241 287
rect 239 286 240 287
rect 238 286 239 287
rect 237 286 238 287
rect 236 286 237 287
rect 235 286 236 287
rect 234 286 235 287
rect 233 286 234 287
rect 232 286 233 287
rect 231 286 232 287
rect 230 286 231 287
rect 229 286 230 287
rect 228 286 229 287
rect 227 286 228 287
rect 226 286 227 287
rect 225 286 226 287
rect 224 286 225 287
rect 223 286 224 287
rect 222 286 223 287
rect 221 286 222 287
rect 220 286 221 287
rect 219 286 220 287
rect 218 286 219 287
rect 217 286 218 287
rect 194 286 195 287
rect 193 286 194 287
rect 192 286 193 287
rect 191 286 192 287
rect 190 286 191 287
rect 189 286 190 287
rect 188 286 189 287
rect 187 286 188 287
rect 186 286 187 287
rect 185 286 186 287
rect 184 286 185 287
rect 183 286 184 287
rect 182 286 183 287
rect 181 286 182 287
rect 180 286 181 287
rect 179 286 180 287
rect 178 286 179 287
rect 177 286 178 287
rect 176 286 177 287
rect 175 286 176 287
rect 174 286 175 287
rect 173 286 174 287
rect 172 286 173 287
rect 171 286 172 287
rect 170 286 171 287
rect 169 286 170 287
rect 168 286 169 287
rect 167 286 168 287
rect 166 286 167 287
rect 165 286 166 287
rect 164 286 165 287
rect 163 286 164 287
rect 162 286 163 287
rect 161 286 162 287
rect 160 286 161 287
rect 159 286 160 287
rect 158 286 159 287
rect 157 286 158 287
rect 156 286 157 287
rect 155 286 156 287
rect 154 286 155 287
rect 153 286 154 287
rect 152 286 153 287
rect 151 286 152 287
rect 150 286 151 287
rect 149 286 150 287
rect 148 286 149 287
rect 147 286 148 287
rect 146 286 147 287
rect 145 286 146 287
rect 144 286 145 287
rect 143 286 144 287
rect 142 286 143 287
rect 141 286 142 287
rect 140 286 141 287
rect 139 286 140 287
rect 138 286 139 287
rect 137 286 138 287
rect 136 286 137 287
rect 135 286 136 287
rect 134 286 135 287
rect 133 286 134 287
rect 132 286 133 287
rect 116 286 117 287
rect 115 286 116 287
rect 114 286 115 287
rect 113 286 114 287
rect 112 286 113 287
rect 111 286 112 287
rect 110 286 111 287
rect 109 286 110 287
rect 108 286 109 287
rect 107 286 108 287
rect 106 286 107 287
rect 105 286 106 287
rect 104 286 105 287
rect 103 286 104 287
rect 102 286 103 287
rect 101 286 102 287
rect 100 286 101 287
rect 99 286 100 287
rect 98 286 99 287
rect 97 286 98 287
rect 96 286 97 287
rect 95 286 96 287
rect 94 286 95 287
rect 93 286 94 287
rect 92 286 93 287
rect 91 286 92 287
rect 90 286 91 287
rect 89 286 90 287
rect 88 286 89 287
rect 87 286 88 287
rect 86 286 87 287
rect 85 286 86 287
rect 84 286 85 287
rect 83 286 84 287
rect 82 286 83 287
rect 66 286 67 287
rect 65 286 66 287
rect 64 286 65 287
rect 63 286 64 287
rect 62 286 63 287
rect 61 286 62 287
rect 60 286 61 287
rect 59 286 60 287
rect 58 286 59 287
rect 57 286 58 287
rect 56 286 57 287
rect 55 286 56 287
rect 54 286 55 287
rect 53 286 54 287
rect 52 286 53 287
rect 51 286 52 287
rect 50 286 51 287
rect 49 286 50 287
rect 48 286 49 287
rect 47 286 48 287
rect 46 286 47 287
rect 45 286 46 287
rect 44 286 45 287
rect 43 286 44 287
rect 42 286 43 287
rect 41 286 42 287
rect 40 286 41 287
rect 39 286 40 287
rect 38 286 39 287
rect 28 286 29 287
rect 27 286 28 287
rect 26 286 27 287
rect 25 286 26 287
rect 24 286 25 287
rect 23 286 24 287
rect 22 286 23 287
rect 21 286 22 287
rect 20 286 21 287
rect 19 286 20 287
rect 18 286 19 287
rect 17 286 18 287
rect 16 286 17 287
rect 15 286 16 287
rect 14 286 15 287
rect 13 286 14 287
rect 12 286 13 287
rect 11 286 12 287
rect 10 286 11 287
rect 9 286 10 287
rect 8 286 9 287
rect 7 286 8 287
rect 6 286 7 287
rect 5 286 6 287
rect 4 286 5 287
rect 3 286 4 287
rect 461 287 462 288
rect 460 287 461 288
rect 439 287 440 288
rect 438 287 439 288
rect 437 287 438 288
rect 436 287 437 288
rect 435 287 436 288
rect 434 287 435 288
rect 433 287 434 288
rect 432 287 433 288
rect 431 287 432 288
rect 430 287 431 288
rect 429 287 430 288
rect 428 287 429 288
rect 427 287 428 288
rect 426 287 427 288
rect 425 287 426 288
rect 424 287 425 288
rect 423 287 424 288
rect 422 287 423 288
rect 421 287 422 288
rect 420 287 421 288
rect 419 287 420 288
rect 418 287 419 288
rect 417 287 418 288
rect 416 287 417 288
rect 415 287 416 288
rect 414 287 415 288
rect 413 287 414 288
rect 412 287 413 288
rect 411 287 412 288
rect 410 287 411 288
rect 409 287 410 288
rect 408 287 409 288
rect 407 287 408 288
rect 406 287 407 288
rect 405 287 406 288
rect 404 287 405 288
rect 403 287 404 288
rect 402 287 403 288
rect 401 287 402 288
rect 400 287 401 288
rect 399 287 400 288
rect 398 287 399 288
rect 397 287 398 288
rect 396 287 397 288
rect 395 287 396 288
rect 283 287 284 288
rect 282 287 283 288
rect 281 287 282 288
rect 280 287 281 288
rect 279 287 280 288
rect 278 287 279 288
rect 277 287 278 288
rect 276 287 277 288
rect 275 287 276 288
rect 274 287 275 288
rect 273 287 274 288
rect 272 287 273 288
rect 271 287 272 288
rect 270 287 271 288
rect 269 287 270 288
rect 268 287 269 288
rect 267 287 268 288
rect 266 287 267 288
rect 265 287 266 288
rect 264 287 265 288
rect 263 287 264 288
rect 262 287 263 288
rect 261 287 262 288
rect 260 287 261 288
rect 259 287 260 288
rect 258 287 259 288
rect 257 287 258 288
rect 256 287 257 288
rect 255 287 256 288
rect 254 287 255 288
rect 253 287 254 288
rect 252 287 253 288
rect 251 287 252 288
rect 250 287 251 288
rect 249 287 250 288
rect 248 287 249 288
rect 247 287 248 288
rect 246 287 247 288
rect 245 287 246 288
rect 244 287 245 288
rect 243 287 244 288
rect 242 287 243 288
rect 241 287 242 288
rect 240 287 241 288
rect 239 287 240 288
rect 238 287 239 288
rect 237 287 238 288
rect 236 287 237 288
rect 235 287 236 288
rect 234 287 235 288
rect 233 287 234 288
rect 232 287 233 288
rect 231 287 232 288
rect 230 287 231 288
rect 229 287 230 288
rect 228 287 229 288
rect 227 287 228 288
rect 226 287 227 288
rect 225 287 226 288
rect 224 287 225 288
rect 223 287 224 288
rect 222 287 223 288
rect 221 287 222 288
rect 220 287 221 288
rect 219 287 220 288
rect 218 287 219 288
rect 217 287 218 288
rect 216 287 217 288
rect 194 287 195 288
rect 193 287 194 288
rect 192 287 193 288
rect 191 287 192 288
rect 190 287 191 288
rect 189 287 190 288
rect 188 287 189 288
rect 187 287 188 288
rect 186 287 187 288
rect 185 287 186 288
rect 184 287 185 288
rect 183 287 184 288
rect 182 287 183 288
rect 181 287 182 288
rect 180 287 181 288
rect 179 287 180 288
rect 178 287 179 288
rect 177 287 178 288
rect 176 287 177 288
rect 175 287 176 288
rect 174 287 175 288
rect 173 287 174 288
rect 172 287 173 288
rect 171 287 172 288
rect 170 287 171 288
rect 169 287 170 288
rect 168 287 169 288
rect 167 287 168 288
rect 166 287 167 288
rect 165 287 166 288
rect 164 287 165 288
rect 163 287 164 288
rect 162 287 163 288
rect 161 287 162 288
rect 160 287 161 288
rect 159 287 160 288
rect 158 287 159 288
rect 157 287 158 288
rect 156 287 157 288
rect 155 287 156 288
rect 154 287 155 288
rect 153 287 154 288
rect 152 287 153 288
rect 151 287 152 288
rect 150 287 151 288
rect 149 287 150 288
rect 148 287 149 288
rect 147 287 148 288
rect 146 287 147 288
rect 145 287 146 288
rect 144 287 145 288
rect 143 287 144 288
rect 142 287 143 288
rect 141 287 142 288
rect 140 287 141 288
rect 139 287 140 288
rect 138 287 139 288
rect 137 287 138 288
rect 136 287 137 288
rect 135 287 136 288
rect 134 287 135 288
rect 133 287 134 288
rect 116 287 117 288
rect 115 287 116 288
rect 114 287 115 288
rect 113 287 114 288
rect 112 287 113 288
rect 111 287 112 288
rect 110 287 111 288
rect 109 287 110 288
rect 108 287 109 288
rect 107 287 108 288
rect 106 287 107 288
rect 105 287 106 288
rect 104 287 105 288
rect 103 287 104 288
rect 102 287 103 288
rect 101 287 102 288
rect 100 287 101 288
rect 99 287 100 288
rect 98 287 99 288
rect 97 287 98 288
rect 96 287 97 288
rect 95 287 96 288
rect 94 287 95 288
rect 93 287 94 288
rect 92 287 93 288
rect 91 287 92 288
rect 90 287 91 288
rect 89 287 90 288
rect 88 287 89 288
rect 87 287 88 288
rect 86 287 87 288
rect 85 287 86 288
rect 84 287 85 288
rect 83 287 84 288
rect 82 287 83 288
rect 66 287 67 288
rect 65 287 66 288
rect 64 287 65 288
rect 63 287 64 288
rect 62 287 63 288
rect 61 287 62 288
rect 60 287 61 288
rect 59 287 60 288
rect 58 287 59 288
rect 57 287 58 288
rect 56 287 57 288
rect 55 287 56 288
rect 54 287 55 288
rect 53 287 54 288
rect 52 287 53 288
rect 51 287 52 288
rect 50 287 51 288
rect 49 287 50 288
rect 48 287 49 288
rect 47 287 48 288
rect 46 287 47 288
rect 45 287 46 288
rect 44 287 45 288
rect 43 287 44 288
rect 42 287 43 288
rect 41 287 42 288
rect 40 287 41 288
rect 39 287 40 288
rect 38 287 39 288
rect 29 287 30 288
rect 28 287 29 288
rect 27 287 28 288
rect 26 287 27 288
rect 25 287 26 288
rect 24 287 25 288
rect 23 287 24 288
rect 22 287 23 288
rect 21 287 22 288
rect 20 287 21 288
rect 19 287 20 288
rect 18 287 19 288
rect 17 287 18 288
rect 16 287 17 288
rect 15 287 16 288
rect 14 287 15 288
rect 13 287 14 288
rect 12 287 13 288
rect 11 287 12 288
rect 10 287 11 288
rect 9 287 10 288
rect 8 287 9 288
rect 7 287 8 288
rect 6 287 7 288
rect 5 287 6 288
rect 4 287 5 288
rect 3 287 4 288
rect 460 288 461 289
rect 439 288 440 289
rect 438 288 439 289
rect 437 288 438 289
rect 436 288 437 289
rect 435 288 436 289
rect 434 288 435 289
rect 433 288 434 289
rect 432 288 433 289
rect 431 288 432 289
rect 430 288 431 289
rect 429 288 430 289
rect 428 288 429 289
rect 427 288 428 289
rect 426 288 427 289
rect 425 288 426 289
rect 424 288 425 289
rect 423 288 424 289
rect 422 288 423 289
rect 421 288 422 289
rect 420 288 421 289
rect 419 288 420 289
rect 418 288 419 289
rect 417 288 418 289
rect 416 288 417 289
rect 415 288 416 289
rect 414 288 415 289
rect 413 288 414 289
rect 412 288 413 289
rect 411 288 412 289
rect 410 288 411 289
rect 409 288 410 289
rect 408 288 409 289
rect 407 288 408 289
rect 406 288 407 289
rect 405 288 406 289
rect 404 288 405 289
rect 403 288 404 289
rect 402 288 403 289
rect 401 288 402 289
rect 400 288 401 289
rect 399 288 400 289
rect 398 288 399 289
rect 397 288 398 289
rect 396 288 397 289
rect 395 288 396 289
rect 282 288 283 289
rect 281 288 282 289
rect 280 288 281 289
rect 279 288 280 289
rect 278 288 279 289
rect 277 288 278 289
rect 276 288 277 289
rect 275 288 276 289
rect 274 288 275 289
rect 273 288 274 289
rect 272 288 273 289
rect 271 288 272 289
rect 270 288 271 289
rect 269 288 270 289
rect 268 288 269 289
rect 267 288 268 289
rect 266 288 267 289
rect 265 288 266 289
rect 264 288 265 289
rect 263 288 264 289
rect 262 288 263 289
rect 261 288 262 289
rect 260 288 261 289
rect 259 288 260 289
rect 258 288 259 289
rect 257 288 258 289
rect 256 288 257 289
rect 255 288 256 289
rect 254 288 255 289
rect 253 288 254 289
rect 252 288 253 289
rect 251 288 252 289
rect 250 288 251 289
rect 249 288 250 289
rect 248 288 249 289
rect 247 288 248 289
rect 246 288 247 289
rect 245 288 246 289
rect 244 288 245 289
rect 243 288 244 289
rect 242 288 243 289
rect 241 288 242 289
rect 240 288 241 289
rect 239 288 240 289
rect 238 288 239 289
rect 237 288 238 289
rect 236 288 237 289
rect 235 288 236 289
rect 234 288 235 289
rect 233 288 234 289
rect 232 288 233 289
rect 231 288 232 289
rect 230 288 231 289
rect 229 288 230 289
rect 228 288 229 289
rect 227 288 228 289
rect 226 288 227 289
rect 225 288 226 289
rect 224 288 225 289
rect 223 288 224 289
rect 222 288 223 289
rect 221 288 222 289
rect 220 288 221 289
rect 219 288 220 289
rect 218 288 219 289
rect 217 288 218 289
rect 216 288 217 289
rect 193 288 194 289
rect 192 288 193 289
rect 191 288 192 289
rect 190 288 191 289
rect 189 288 190 289
rect 188 288 189 289
rect 187 288 188 289
rect 186 288 187 289
rect 185 288 186 289
rect 184 288 185 289
rect 183 288 184 289
rect 182 288 183 289
rect 181 288 182 289
rect 180 288 181 289
rect 179 288 180 289
rect 178 288 179 289
rect 177 288 178 289
rect 176 288 177 289
rect 175 288 176 289
rect 174 288 175 289
rect 173 288 174 289
rect 172 288 173 289
rect 171 288 172 289
rect 170 288 171 289
rect 169 288 170 289
rect 168 288 169 289
rect 167 288 168 289
rect 166 288 167 289
rect 165 288 166 289
rect 164 288 165 289
rect 163 288 164 289
rect 162 288 163 289
rect 161 288 162 289
rect 160 288 161 289
rect 159 288 160 289
rect 158 288 159 289
rect 157 288 158 289
rect 156 288 157 289
rect 155 288 156 289
rect 154 288 155 289
rect 153 288 154 289
rect 152 288 153 289
rect 151 288 152 289
rect 150 288 151 289
rect 149 288 150 289
rect 148 288 149 289
rect 147 288 148 289
rect 146 288 147 289
rect 145 288 146 289
rect 144 288 145 289
rect 143 288 144 289
rect 142 288 143 289
rect 141 288 142 289
rect 140 288 141 289
rect 139 288 140 289
rect 138 288 139 289
rect 137 288 138 289
rect 136 288 137 289
rect 135 288 136 289
rect 134 288 135 289
rect 133 288 134 289
rect 117 288 118 289
rect 116 288 117 289
rect 115 288 116 289
rect 114 288 115 289
rect 113 288 114 289
rect 112 288 113 289
rect 111 288 112 289
rect 110 288 111 289
rect 109 288 110 289
rect 108 288 109 289
rect 107 288 108 289
rect 106 288 107 289
rect 105 288 106 289
rect 104 288 105 289
rect 103 288 104 289
rect 102 288 103 289
rect 101 288 102 289
rect 100 288 101 289
rect 99 288 100 289
rect 98 288 99 289
rect 97 288 98 289
rect 96 288 97 289
rect 95 288 96 289
rect 94 288 95 289
rect 93 288 94 289
rect 92 288 93 289
rect 91 288 92 289
rect 90 288 91 289
rect 89 288 90 289
rect 88 288 89 289
rect 87 288 88 289
rect 86 288 87 289
rect 85 288 86 289
rect 84 288 85 289
rect 83 288 84 289
rect 82 288 83 289
rect 66 288 67 289
rect 65 288 66 289
rect 64 288 65 289
rect 63 288 64 289
rect 62 288 63 289
rect 61 288 62 289
rect 60 288 61 289
rect 59 288 60 289
rect 58 288 59 289
rect 57 288 58 289
rect 56 288 57 289
rect 55 288 56 289
rect 54 288 55 289
rect 53 288 54 289
rect 52 288 53 289
rect 51 288 52 289
rect 50 288 51 289
rect 49 288 50 289
rect 48 288 49 289
rect 47 288 48 289
rect 46 288 47 289
rect 45 288 46 289
rect 44 288 45 289
rect 43 288 44 289
rect 42 288 43 289
rect 41 288 42 289
rect 40 288 41 289
rect 39 288 40 289
rect 38 288 39 289
rect 29 288 30 289
rect 28 288 29 289
rect 27 288 28 289
rect 26 288 27 289
rect 25 288 26 289
rect 24 288 25 289
rect 23 288 24 289
rect 22 288 23 289
rect 21 288 22 289
rect 20 288 21 289
rect 19 288 20 289
rect 18 288 19 289
rect 17 288 18 289
rect 16 288 17 289
rect 15 288 16 289
rect 14 288 15 289
rect 13 288 14 289
rect 12 288 13 289
rect 11 288 12 289
rect 10 288 11 289
rect 9 288 10 289
rect 8 288 9 289
rect 7 288 8 289
rect 6 288 7 289
rect 5 288 6 289
rect 4 288 5 289
rect 3 288 4 289
rect 480 289 481 290
rect 460 289 461 290
rect 439 289 440 290
rect 438 289 439 290
rect 437 289 438 290
rect 436 289 437 290
rect 435 289 436 290
rect 434 289 435 290
rect 418 289 419 290
rect 417 289 418 290
rect 416 289 417 290
rect 415 289 416 290
rect 414 289 415 290
rect 401 289 402 290
rect 400 289 401 290
rect 399 289 400 290
rect 398 289 399 290
rect 397 289 398 290
rect 396 289 397 290
rect 395 289 396 290
rect 281 289 282 290
rect 280 289 281 290
rect 279 289 280 290
rect 278 289 279 290
rect 277 289 278 290
rect 276 289 277 290
rect 275 289 276 290
rect 274 289 275 290
rect 273 289 274 290
rect 272 289 273 290
rect 271 289 272 290
rect 270 289 271 290
rect 269 289 270 290
rect 268 289 269 290
rect 267 289 268 290
rect 266 289 267 290
rect 265 289 266 290
rect 264 289 265 290
rect 263 289 264 290
rect 262 289 263 290
rect 261 289 262 290
rect 260 289 261 290
rect 259 289 260 290
rect 258 289 259 290
rect 257 289 258 290
rect 256 289 257 290
rect 255 289 256 290
rect 254 289 255 290
rect 253 289 254 290
rect 252 289 253 290
rect 251 289 252 290
rect 250 289 251 290
rect 249 289 250 290
rect 248 289 249 290
rect 247 289 248 290
rect 246 289 247 290
rect 245 289 246 290
rect 244 289 245 290
rect 243 289 244 290
rect 242 289 243 290
rect 241 289 242 290
rect 240 289 241 290
rect 239 289 240 290
rect 238 289 239 290
rect 237 289 238 290
rect 236 289 237 290
rect 235 289 236 290
rect 234 289 235 290
rect 233 289 234 290
rect 232 289 233 290
rect 231 289 232 290
rect 230 289 231 290
rect 229 289 230 290
rect 228 289 229 290
rect 227 289 228 290
rect 226 289 227 290
rect 225 289 226 290
rect 224 289 225 290
rect 223 289 224 290
rect 222 289 223 290
rect 221 289 222 290
rect 220 289 221 290
rect 219 289 220 290
rect 218 289 219 290
rect 217 289 218 290
rect 216 289 217 290
rect 215 289 216 290
rect 192 289 193 290
rect 191 289 192 290
rect 190 289 191 290
rect 189 289 190 290
rect 188 289 189 290
rect 187 289 188 290
rect 186 289 187 290
rect 185 289 186 290
rect 184 289 185 290
rect 183 289 184 290
rect 182 289 183 290
rect 181 289 182 290
rect 180 289 181 290
rect 179 289 180 290
rect 178 289 179 290
rect 177 289 178 290
rect 176 289 177 290
rect 175 289 176 290
rect 174 289 175 290
rect 173 289 174 290
rect 172 289 173 290
rect 171 289 172 290
rect 170 289 171 290
rect 169 289 170 290
rect 168 289 169 290
rect 167 289 168 290
rect 166 289 167 290
rect 165 289 166 290
rect 164 289 165 290
rect 163 289 164 290
rect 162 289 163 290
rect 161 289 162 290
rect 160 289 161 290
rect 159 289 160 290
rect 158 289 159 290
rect 157 289 158 290
rect 156 289 157 290
rect 155 289 156 290
rect 154 289 155 290
rect 153 289 154 290
rect 152 289 153 290
rect 151 289 152 290
rect 150 289 151 290
rect 149 289 150 290
rect 148 289 149 290
rect 147 289 148 290
rect 146 289 147 290
rect 145 289 146 290
rect 144 289 145 290
rect 143 289 144 290
rect 142 289 143 290
rect 141 289 142 290
rect 140 289 141 290
rect 139 289 140 290
rect 138 289 139 290
rect 137 289 138 290
rect 136 289 137 290
rect 135 289 136 290
rect 134 289 135 290
rect 117 289 118 290
rect 116 289 117 290
rect 115 289 116 290
rect 114 289 115 290
rect 113 289 114 290
rect 112 289 113 290
rect 111 289 112 290
rect 110 289 111 290
rect 109 289 110 290
rect 108 289 109 290
rect 107 289 108 290
rect 106 289 107 290
rect 105 289 106 290
rect 104 289 105 290
rect 103 289 104 290
rect 102 289 103 290
rect 101 289 102 290
rect 100 289 101 290
rect 99 289 100 290
rect 98 289 99 290
rect 97 289 98 290
rect 96 289 97 290
rect 95 289 96 290
rect 94 289 95 290
rect 93 289 94 290
rect 92 289 93 290
rect 91 289 92 290
rect 90 289 91 290
rect 89 289 90 290
rect 88 289 89 290
rect 87 289 88 290
rect 86 289 87 290
rect 85 289 86 290
rect 84 289 85 290
rect 83 289 84 290
rect 67 289 68 290
rect 66 289 67 290
rect 65 289 66 290
rect 64 289 65 290
rect 63 289 64 290
rect 62 289 63 290
rect 61 289 62 290
rect 60 289 61 290
rect 59 289 60 290
rect 58 289 59 290
rect 57 289 58 290
rect 56 289 57 290
rect 55 289 56 290
rect 54 289 55 290
rect 53 289 54 290
rect 52 289 53 290
rect 51 289 52 290
rect 50 289 51 290
rect 49 289 50 290
rect 48 289 49 290
rect 47 289 48 290
rect 46 289 47 290
rect 45 289 46 290
rect 44 289 45 290
rect 43 289 44 290
rect 42 289 43 290
rect 41 289 42 290
rect 40 289 41 290
rect 39 289 40 290
rect 38 289 39 290
rect 29 289 30 290
rect 28 289 29 290
rect 27 289 28 290
rect 26 289 27 290
rect 25 289 26 290
rect 24 289 25 290
rect 23 289 24 290
rect 22 289 23 290
rect 21 289 22 290
rect 20 289 21 290
rect 19 289 20 290
rect 18 289 19 290
rect 17 289 18 290
rect 16 289 17 290
rect 15 289 16 290
rect 14 289 15 290
rect 13 289 14 290
rect 12 289 13 290
rect 11 289 12 290
rect 10 289 11 290
rect 9 289 10 290
rect 8 289 9 290
rect 7 289 8 290
rect 6 289 7 290
rect 5 289 6 290
rect 4 289 5 290
rect 3 289 4 290
rect 480 290 481 291
rect 460 290 461 291
rect 439 290 440 291
rect 438 290 439 291
rect 437 290 438 291
rect 436 290 437 291
rect 417 290 418 291
rect 416 290 417 291
rect 415 290 416 291
rect 414 290 415 291
rect 398 290 399 291
rect 397 290 398 291
rect 396 290 397 291
rect 395 290 396 291
rect 280 290 281 291
rect 279 290 280 291
rect 278 290 279 291
rect 277 290 278 291
rect 276 290 277 291
rect 275 290 276 291
rect 274 290 275 291
rect 273 290 274 291
rect 272 290 273 291
rect 271 290 272 291
rect 270 290 271 291
rect 269 290 270 291
rect 268 290 269 291
rect 267 290 268 291
rect 266 290 267 291
rect 265 290 266 291
rect 264 290 265 291
rect 263 290 264 291
rect 262 290 263 291
rect 261 290 262 291
rect 260 290 261 291
rect 259 290 260 291
rect 258 290 259 291
rect 257 290 258 291
rect 256 290 257 291
rect 255 290 256 291
rect 254 290 255 291
rect 253 290 254 291
rect 252 290 253 291
rect 251 290 252 291
rect 250 290 251 291
rect 249 290 250 291
rect 248 290 249 291
rect 247 290 248 291
rect 246 290 247 291
rect 245 290 246 291
rect 244 290 245 291
rect 243 290 244 291
rect 242 290 243 291
rect 241 290 242 291
rect 240 290 241 291
rect 239 290 240 291
rect 238 290 239 291
rect 237 290 238 291
rect 236 290 237 291
rect 235 290 236 291
rect 234 290 235 291
rect 233 290 234 291
rect 232 290 233 291
rect 231 290 232 291
rect 230 290 231 291
rect 229 290 230 291
rect 228 290 229 291
rect 227 290 228 291
rect 226 290 227 291
rect 225 290 226 291
rect 224 290 225 291
rect 223 290 224 291
rect 222 290 223 291
rect 221 290 222 291
rect 220 290 221 291
rect 219 290 220 291
rect 218 290 219 291
rect 217 290 218 291
rect 216 290 217 291
rect 215 290 216 291
rect 191 290 192 291
rect 190 290 191 291
rect 189 290 190 291
rect 188 290 189 291
rect 187 290 188 291
rect 186 290 187 291
rect 185 290 186 291
rect 184 290 185 291
rect 183 290 184 291
rect 182 290 183 291
rect 181 290 182 291
rect 180 290 181 291
rect 179 290 180 291
rect 178 290 179 291
rect 177 290 178 291
rect 176 290 177 291
rect 175 290 176 291
rect 174 290 175 291
rect 173 290 174 291
rect 172 290 173 291
rect 171 290 172 291
rect 170 290 171 291
rect 169 290 170 291
rect 168 290 169 291
rect 167 290 168 291
rect 166 290 167 291
rect 165 290 166 291
rect 164 290 165 291
rect 163 290 164 291
rect 162 290 163 291
rect 161 290 162 291
rect 160 290 161 291
rect 159 290 160 291
rect 158 290 159 291
rect 157 290 158 291
rect 156 290 157 291
rect 155 290 156 291
rect 154 290 155 291
rect 153 290 154 291
rect 152 290 153 291
rect 151 290 152 291
rect 150 290 151 291
rect 149 290 150 291
rect 148 290 149 291
rect 147 290 148 291
rect 146 290 147 291
rect 145 290 146 291
rect 144 290 145 291
rect 143 290 144 291
rect 142 290 143 291
rect 141 290 142 291
rect 140 290 141 291
rect 139 290 140 291
rect 138 290 139 291
rect 137 290 138 291
rect 136 290 137 291
rect 135 290 136 291
rect 118 290 119 291
rect 117 290 118 291
rect 116 290 117 291
rect 115 290 116 291
rect 114 290 115 291
rect 113 290 114 291
rect 112 290 113 291
rect 111 290 112 291
rect 110 290 111 291
rect 109 290 110 291
rect 108 290 109 291
rect 107 290 108 291
rect 106 290 107 291
rect 105 290 106 291
rect 104 290 105 291
rect 103 290 104 291
rect 102 290 103 291
rect 101 290 102 291
rect 100 290 101 291
rect 99 290 100 291
rect 98 290 99 291
rect 97 290 98 291
rect 96 290 97 291
rect 95 290 96 291
rect 94 290 95 291
rect 93 290 94 291
rect 92 290 93 291
rect 91 290 92 291
rect 90 290 91 291
rect 89 290 90 291
rect 88 290 89 291
rect 87 290 88 291
rect 86 290 87 291
rect 85 290 86 291
rect 84 290 85 291
rect 83 290 84 291
rect 67 290 68 291
rect 66 290 67 291
rect 65 290 66 291
rect 64 290 65 291
rect 63 290 64 291
rect 62 290 63 291
rect 61 290 62 291
rect 60 290 61 291
rect 59 290 60 291
rect 58 290 59 291
rect 57 290 58 291
rect 56 290 57 291
rect 55 290 56 291
rect 54 290 55 291
rect 53 290 54 291
rect 52 290 53 291
rect 51 290 52 291
rect 50 290 51 291
rect 49 290 50 291
rect 48 290 49 291
rect 47 290 48 291
rect 46 290 47 291
rect 45 290 46 291
rect 44 290 45 291
rect 43 290 44 291
rect 42 290 43 291
rect 41 290 42 291
rect 40 290 41 291
rect 39 290 40 291
rect 38 290 39 291
rect 29 290 30 291
rect 28 290 29 291
rect 27 290 28 291
rect 26 290 27 291
rect 25 290 26 291
rect 24 290 25 291
rect 23 290 24 291
rect 22 290 23 291
rect 21 290 22 291
rect 20 290 21 291
rect 19 290 20 291
rect 18 290 19 291
rect 17 290 18 291
rect 16 290 17 291
rect 15 290 16 291
rect 14 290 15 291
rect 13 290 14 291
rect 12 290 13 291
rect 11 290 12 291
rect 10 290 11 291
rect 9 290 10 291
rect 8 290 9 291
rect 7 290 8 291
rect 6 290 7 291
rect 5 290 6 291
rect 4 290 5 291
rect 3 290 4 291
rect 480 291 481 292
rect 479 291 480 292
rect 460 291 461 292
rect 439 291 440 292
rect 438 291 439 292
rect 437 291 438 292
rect 417 291 418 292
rect 416 291 417 292
rect 415 291 416 292
rect 414 291 415 292
rect 397 291 398 292
rect 396 291 397 292
rect 395 291 396 292
rect 279 291 280 292
rect 278 291 279 292
rect 277 291 278 292
rect 276 291 277 292
rect 275 291 276 292
rect 274 291 275 292
rect 273 291 274 292
rect 272 291 273 292
rect 271 291 272 292
rect 270 291 271 292
rect 269 291 270 292
rect 268 291 269 292
rect 267 291 268 292
rect 266 291 267 292
rect 265 291 266 292
rect 264 291 265 292
rect 263 291 264 292
rect 262 291 263 292
rect 261 291 262 292
rect 260 291 261 292
rect 259 291 260 292
rect 258 291 259 292
rect 257 291 258 292
rect 256 291 257 292
rect 255 291 256 292
rect 254 291 255 292
rect 253 291 254 292
rect 252 291 253 292
rect 251 291 252 292
rect 250 291 251 292
rect 249 291 250 292
rect 248 291 249 292
rect 247 291 248 292
rect 246 291 247 292
rect 245 291 246 292
rect 244 291 245 292
rect 243 291 244 292
rect 242 291 243 292
rect 241 291 242 292
rect 240 291 241 292
rect 239 291 240 292
rect 238 291 239 292
rect 237 291 238 292
rect 236 291 237 292
rect 235 291 236 292
rect 234 291 235 292
rect 233 291 234 292
rect 232 291 233 292
rect 231 291 232 292
rect 230 291 231 292
rect 229 291 230 292
rect 228 291 229 292
rect 227 291 228 292
rect 226 291 227 292
rect 225 291 226 292
rect 224 291 225 292
rect 223 291 224 292
rect 222 291 223 292
rect 221 291 222 292
rect 220 291 221 292
rect 219 291 220 292
rect 218 291 219 292
rect 217 291 218 292
rect 216 291 217 292
rect 215 291 216 292
rect 214 291 215 292
rect 191 291 192 292
rect 190 291 191 292
rect 189 291 190 292
rect 188 291 189 292
rect 187 291 188 292
rect 186 291 187 292
rect 185 291 186 292
rect 184 291 185 292
rect 183 291 184 292
rect 182 291 183 292
rect 181 291 182 292
rect 180 291 181 292
rect 179 291 180 292
rect 178 291 179 292
rect 177 291 178 292
rect 176 291 177 292
rect 175 291 176 292
rect 174 291 175 292
rect 173 291 174 292
rect 172 291 173 292
rect 171 291 172 292
rect 170 291 171 292
rect 169 291 170 292
rect 168 291 169 292
rect 167 291 168 292
rect 166 291 167 292
rect 165 291 166 292
rect 164 291 165 292
rect 163 291 164 292
rect 162 291 163 292
rect 161 291 162 292
rect 160 291 161 292
rect 159 291 160 292
rect 158 291 159 292
rect 157 291 158 292
rect 156 291 157 292
rect 155 291 156 292
rect 154 291 155 292
rect 153 291 154 292
rect 152 291 153 292
rect 151 291 152 292
rect 150 291 151 292
rect 149 291 150 292
rect 148 291 149 292
rect 147 291 148 292
rect 146 291 147 292
rect 145 291 146 292
rect 144 291 145 292
rect 143 291 144 292
rect 142 291 143 292
rect 141 291 142 292
rect 140 291 141 292
rect 139 291 140 292
rect 138 291 139 292
rect 137 291 138 292
rect 136 291 137 292
rect 135 291 136 292
rect 118 291 119 292
rect 117 291 118 292
rect 116 291 117 292
rect 115 291 116 292
rect 114 291 115 292
rect 113 291 114 292
rect 112 291 113 292
rect 111 291 112 292
rect 110 291 111 292
rect 109 291 110 292
rect 108 291 109 292
rect 107 291 108 292
rect 106 291 107 292
rect 105 291 106 292
rect 104 291 105 292
rect 103 291 104 292
rect 102 291 103 292
rect 101 291 102 292
rect 100 291 101 292
rect 99 291 100 292
rect 98 291 99 292
rect 97 291 98 292
rect 96 291 97 292
rect 95 291 96 292
rect 94 291 95 292
rect 93 291 94 292
rect 92 291 93 292
rect 91 291 92 292
rect 90 291 91 292
rect 89 291 90 292
rect 88 291 89 292
rect 87 291 88 292
rect 86 291 87 292
rect 85 291 86 292
rect 84 291 85 292
rect 83 291 84 292
rect 67 291 68 292
rect 66 291 67 292
rect 65 291 66 292
rect 64 291 65 292
rect 63 291 64 292
rect 62 291 63 292
rect 61 291 62 292
rect 60 291 61 292
rect 59 291 60 292
rect 58 291 59 292
rect 57 291 58 292
rect 56 291 57 292
rect 55 291 56 292
rect 54 291 55 292
rect 53 291 54 292
rect 52 291 53 292
rect 51 291 52 292
rect 50 291 51 292
rect 49 291 50 292
rect 48 291 49 292
rect 47 291 48 292
rect 46 291 47 292
rect 45 291 46 292
rect 44 291 45 292
rect 43 291 44 292
rect 42 291 43 292
rect 41 291 42 292
rect 40 291 41 292
rect 39 291 40 292
rect 38 291 39 292
rect 29 291 30 292
rect 28 291 29 292
rect 27 291 28 292
rect 26 291 27 292
rect 25 291 26 292
rect 24 291 25 292
rect 23 291 24 292
rect 22 291 23 292
rect 21 291 22 292
rect 20 291 21 292
rect 19 291 20 292
rect 18 291 19 292
rect 17 291 18 292
rect 16 291 17 292
rect 15 291 16 292
rect 14 291 15 292
rect 13 291 14 292
rect 12 291 13 292
rect 11 291 12 292
rect 10 291 11 292
rect 9 291 10 292
rect 8 291 9 292
rect 7 291 8 292
rect 6 291 7 292
rect 5 291 6 292
rect 4 291 5 292
rect 3 291 4 292
rect 480 292 481 293
rect 479 292 480 293
rect 478 292 479 293
rect 477 292 478 293
rect 476 292 477 293
rect 475 292 476 293
rect 474 292 475 293
rect 473 292 474 293
rect 472 292 473 293
rect 471 292 472 293
rect 470 292 471 293
rect 469 292 470 293
rect 468 292 469 293
rect 467 292 468 293
rect 466 292 467 293
rect 465 292 466 293
rect 464 292 465 293
rect 463 292 464 293
rect 462 292 463 293
rect 461 292 462 293
rect 460 292 461 293
rect 439 292 440 293
rect 438 292 439 293
rect 437 292 438 293
rect 417 292 418 293
rect 416 292 417 293
rect 415 292 416 293
rect 414 292 415 293
rect 397 292 398 293
rect 396 292 397 293
rect 395 292 396 293
rect 278 292 279 293
rect 277 292 278 293
rect 276 292 277 293
rect 275 292 276 293
rect 274 292 275 293
rect 273 292 274 293
rect 272 292 273 293
rect 271 292 272 293
rect 270 292 271 293
rect 269 292 270 293
rect 268 292 269 293
rect 267 292 268 293
rect 266 292 267 293
rect 265 292 266 293
rect 264 292 265 293
rect 263 292 264 293
rect 262 292 263 293
rect 261 292 262 293
rect 260 292 261 293
rect 259 292 260 293
rect 258 292 259 293
rect 257 292 258 293
rect 256 292 257 293
rect 255 292 256 293
rect 254 292 255 293
rect 253 292 254 293
rect 252 292 253 293
rect 251 292 252 293
rect 250 292 251 293
rect 249 292 250 293
rect 248 292 249 293
rect 247 292 248 293
rect 246 292 247 293
rect 245 292 246 293
rect 244 292 245 293
rect 243 292 244 293
rect 242 292 243 293
rect 241 292 242 293
rect 240 292 241 293
rect 239 292 240 293
rect 238 292 239 293
rect 237 292 238 293
rect 236 292 237 293
rect 235 292 236 293
rect 234 292 235 293
rect 233 292 234 293
rect 232 292 233 293
rect 231 292 232 293
rect 230 292 231 293
rect 229 292 230 293
rect 228 292 229 293
rect 227 292 228 293
rect 226 292 227 293
rect 225 292 226 293
rect 224 292 225 293
rect 223 292 224 293
rect 222 292 223 293
rect 221 292 222 293
rect 220 292 221 293
rect 219 292 220 293
rect 218 292 219 293
rect 217 292 218 293
rect 216 292 217 293
rect 215 292 216 293
rect 214 292 215 293
rect 213 292 214 293
rect 190 292 191 293
rect 189 292 190 293
rect 188 292 189 293
rect 187 292 188 293
rect 186 292 187 293
rect 185 292 186 293
rect 184 292 185 293
rect 183 292 184 293
rect 182 292 183 293
rect 181 292 182 293
rect 180 292 181 293
rect 179 292 180 293
rect 178 292 179 293
rect 177 292 178 293
rect 176 292 177 293
rect 175 292 176 293
rect 174 292 175 293
rect 173 292 174 293
rect 172 292 173 293
rect 171 292 172 293
rect 170 292 171 293
rect 169 292 170 293
rect 168 292 169 293
rect 167 292 168 293
rect 166 292 167 293
rect 165 292 166 293
rect 164 292 165 293
rect 163 292 164 293
rect 162 292 163 293
rect 161 292 162 293
rect 160 292 161 293
rect 159 292 160 293
rect 158 292 159 293
rect 157 292 158 293
rect 156 292 157 293
rect 155 292 156 293
rect 154 292 155 293
rect 153 292 154 293
rect 152 292 153 293
rect 151 292 152 293
rect 150 292 151 293
rect 149 292 150 293
rect 148 292 149 293
rect 147 292 148 293
rect 146 292 147 293
rect 145 292 146 293
rect 144 292 145 293
rect 143 292 144 293
rect 142 292 143 293
rect 141 292 142 293
rect 140 292 141 293
rect 139 292 140 293
rect 138 292 139 293
rect 137 292 138 293
rect 136 292 137 293
rect 118 292 119 293
rect 117 292 118 293
rect 116 292 117 293
rect 115 292 116 293
rect 114 292 115 293
rect 113 292 114 293
rect 112 292 113 293
rect 111 292 112 293
rect 110 292 111 293
rect 109 292 110 293
rect 108 292 109 293
rect 107 292 108 293
rect 106 292 107 293
rect 105 292 106 293
rect 104 292 105 293
rect 103 292 104 293
rect 102 292 103 293
rect 101 292 102 293
rect 100 292 101 293
rect 99 292 100 293
rect 98 292 99 293
rect 97 292 98 293
rect 96 292 97 293
rect 95 292 96 293
rect 94 292 95 293
rect 93 292 94 293
rect 92 292 93 293
rect 91 292 92 293
rect 90 292 91 293
rect 89 292 90 293
rect 88 292 89 293
rect 87 292 88 293
rect 86 292 87 293
rect 85 292 86 293
rect 84 292 85 293
rect 83 292 84 293
rect 67 292 68 293
rect 66 292 67 293
rect 65 292 66 293
rect 64 292 65 293
rect 63 292 64 293
rect 62 292 63 293
rect 61 292 62 293
rect 60 292 61 293
rect 59 292 60 293
rect 58 292 59 293
rect 57 292 58 293
rect 56 292 57 293
rect 55 292 56 293
rect 54 292 55 293
rect 53 292 54 293
rect 52 292 53 293
rect 51 292 52 293
rect 50 292 51 293
rect 49 292 50 293
rect 48 292 49 293
rect 47 292 48 293
rect 46 292 47 293
rect 45 292 46 293
rect 44 292 45 293
rect 43 292 44 293
rect 42 292 43 293
rect 41 292 42 293
rect 40 292 41 293
rect 39 292 40 293
rect 29 292 30 293
rect 28 292 29 293
rect 27 292 28 293
rect 26 292 27 293
rect 25 292 26 293
rect 24 292 25 293
rect 23 292 24 293
rect 22 292 23 293
rect 21 292 22 293
rect 20 292 21 293
rect 19 292 20 293
rect 18 292 19 293
rect 17 292 18 293
rect 16 292 17 293
rect 15 292 16 293
rect 14 292 15 293
rect 13 292 14 293
rect 12 292 13 293
rect 11 292 12 293
rect 10 292 11 293
rect 9 292 10 293
rect 8 292 9 293
rect 7 292 8 293
rect 6 292 7 293
rect 5 292 6 293
rect 4 292 5 293
rect 3 292 4 293
rect 480 293 481 294
rect 479 293 480 294
rect 478 293 479 294
rect 477 293 478 294
rect 476 293 477 294
rect 475 293 476 294
rect 474 293 475 294
rect 473 293 474 294
rect 472 293 473 294
rect 471 293 472 294
rect 470 293 471 294
rect 469 293 470 294
rect 468 293 469 294
rect 467 293 468 294
rect 466 293 467 294
rect 465 293 466 294
rect 464 293 465 294
rect 463 293 464 294
rect 462 293 463 294
rect 461 293 462 294
rect 460 293 461 294
rect 439 293 440 294
rect 438 293 439 294
rect 437 293 438 294
rect 417 293 418 294
rect 416 293 417 294
rect 415 293 416 294
rect 414 293 415 294
rect 397 293 398 294
rect 396 293 397 294
rect 395 293 396 294
rect 277 293 278 294
rect 276 293 277 294
rect 275 293 276 294
rect 274 293 275 294
rect 273 293 274 294
rect 272 293 273 294
rect 271 293 272 294
rect 270 293 271 294
rect 269 293 270 294
rect 268 293 269 294
rect 267 293 268 294
rect 266 293 267 294
rect 265 293 266 294
rect 264 293 265 294
rect 263 293 264 294
rect 262 293 263 294
rect 261 293 262 294
rect 260 293 261 294
rect 259 293 260 294
rect 258 293 259 294
rect 257 293 258 294
rect 256 293 257 294
rect 255 293 256 294
rect 254 293 255 294
rect 253 293 254 294
rect 252 293 253 294
rect 251 293 252 294
rect 250 293 251 294
rect 249 293 250 294
rect 248 293 249 294
rect 247 293 248 294
rect 246 293 247 294
rect 245 293 246 294
rect 244 293 245 294
rect 243 293 244 294
rect 242 293 243 294
rect 241 293 242 294
rect 240 293 241 294
rect 239 293 240 294
rect 238 293 239 294
rect 237 293 238 294
rect 236 293 237 294
rect 235 293 236 294
rect 234 293 235 294
rect 233 293 234 294
rect 232 293 233 294
rect 231 293 232 294
rect 230 293 231 294
rect 229 293 230 294
rect 228 293 229 294
rect 227 293 228 294
rect 226 293 227 294
rect 225 293 226 294
rect 224 293 225 294
rect 223 293 224 294
rect 222 293 223 294
rect 221 293 222 294
rect 220 293 221 294
rect 219 293 220 294
rect 218 293 219 294
rect 217 293 218 294
rect 216 293 217 294
rect 215 293 216 294
rect 214 293 215 294
rect 213 293 214 294
rect 189 293 190 294
rect 188 293 189 294
rect 187 293 188 294
rect 186 293 187 294
rect 185 293 186 294
rect 184 293 185 294
rect 183 293 184 294
rect 182 293 183 294
rect 181 293 182 294
rect 180 293 181 294
rect 179 293 180 294
rect 178 293 179 294
rect 177 293 178 294
rect 176 293 177 294
rect 175 293 176 294
rect 174 293 175 294
rect 173 293 174 294
rect 172 293 173 294
rect 171 293 172 294
rect 170 293 171 294
rect 169 293 170 294
rect 168 293 169 294
rect 167 293 168 294
rect 166 293 167 294
rect 165 293 166 294
rect 164 293 165 294
rect 163 293 164 294
rect 162 293 163 294
rect 161 293 162 294
rect 160 293 161 294
rect 159 293 160 294
rect 158 293 159 294
rect 157 293 158 294
rect 156 293 157 294
rect 155 293 156 294
rect 154 293 155 294
rect 153 293 154 294
rect 152 293 153 294
rect 151 293 152 294
rect 150 293 151 294
rect 149 293 150 294
rect 148 293 149 294
rect 147 293 148 294
rect 146 293 147 294
rect 145 293 146 294
rect 144 293 145 294
rect 143 293 144 294
rect 142 293 143 294
rect 141 293 142 294
rect 140 293 141 294
rect 139 293 140 294
rect 138 293 139 294
rect 137 293 138 294
rect 119 293 120 294
rect 118 293 119 294
rect 117 293 118 294
rect 116 293 117 294
rect 115 293 116 294
rect 114 293 115 294
rect 113 293 114 294
rect 112 293 113 294
rect 111 293 112 294
rect 110 293 111 294
rect 109 293 110 294
rect 108 293 109 294
rect 107 293 108 294
rect 106 293 107 294
rect 105 293 106 294
rect 104 293 105 294
rect 103 293 104 294
rect 102 293 103 294
rect 101 293 102 294
rect 100 293 101 294
rect 99 293 100 294
rect 98 293 99 294
rect 97 293 98 294
rect 96 293 97 294
rect 95 293 96 294
rect 94 293 95 294
rect 93 293 94 294
rect 92 293 93 294
rect 91 293 92 294
rect 90 293 91 294
rect 89 293 90 294
rect 88 293 89 294
rect 87 293 88 294
rect 86 293 87 294
rect 85 293 86 294
rect 84 293 85 294
rect 68 293 69 294
rect 67 293 68 294
rect 66 293 67 294
rect 65 293 66 294
rect 64 293 65 294
rect 63 293 64 294
rect 62 293 63 294
rect 61 293 62 294
rect 60 293 61 294
rect 59 293 60 294
rect 58 293 59 294
rect 57 293 58 294
rect 56 293 57 294
rect 55 293 56 294
rect 54 293 55 294
rect 53 293 54 294
rect 52 293 53 294
rect 51 293 52 294
rect 50 293 51 294
rect 49 293 50 294
rect 48 293 49 294
rect 47 293 48 294
rect 46 293 47 294
rect 45 293 46 294
rect 44 293 45 294
rect 43 293 44 294
rect 42 293 43 294
rect 41 293 42 294
rect 40 293 41 294
rect 39 293 40 294
rect 29 293 30 294
rect 28 293 29 294
rect 27 293 28 294
rect 26 293 27 294
rect 25 293 26 294
rect 24 293 25 294
rect 23 293 24 294
rect 22 293 23 294
rect 21 293 22 294
rect 20 293 21 294
rect 19 293 20 294
rect 18 293 19 294
rect 17 293 18 294
rect 16 293 17 294
rect 15 293 16 294
rect 14 293 15 294
rect 13 293 14 294
rect 12 293 13 294
rect 11 293 12 294
rect 10 293 11 294
rect 9 293 10 294
rect 8 293 9 294
rect 7 293 8 294
rect 6 293 7 294
rect 5 293 6 294
rect 4 293 5 294
rect 3 293 4 294
rect 480 294 481 295
rect 479 294 480 295
rect 478 294 479 295
rect 477 294 478 295
rect 476 294 477 295
rect 475 294 476 295
rect 474 294 475 295
rect 473 294 474 295
rect 472 294 473 295
rect 471 294 472 295
rect 470 294 471 295
rect 469 294 470 295
rect 468 294 469 295
rect 467 294 468 295
rect 466 294 467 295
rect 465 294 466 295
rect 464 294 465 295
rect 463 294 464 295
rect 462 294 463 295
rect 461 294 462 295
rect 460 294 461 295
rect 439 294 440 295
rect 438 294 439 295
rect 417 294 418 295
rect 416 294 417 295
rect 415 294 416 295
rect 414 294 415 295
rect 397 294 398 295
rect 396 294 397 295
rect 395 294 396 295
rect 276 294 277 295
rect 275 294 276 295
rect 274 294 275 295
rect 273 294 274 295
rect 272 294 273 295
rect 271 294 272 295
rect 270 294 271 295
rect 269 294 270 295
rect 268 294 269 295
rect 267 294 268 295
rect 266 294 267 295
rect 265 294 266 295
rect 264 294 265 295
rect 263 294 264 295
rect 262 294 263 295
rect 261 294 262 295
rect 260 294 261 295
rect 259 294 260 295
rect 258 294 259 295
rect 257 294 258 295
rect 256 294 257 295
rect 255 294 256 295
rect 254 294 255 295
rect 253 294 254 295
rect 252 294 253 295
rect 251 294 252 295
rect 250 294 251 295
rect 249 294 250 295
rect 248 294 249 295
rect 247 294 248 295
rect 246 294 247 295
rect 245 294 246 295
rect 244 294 245 295
rect 243 294 244 295
rect 242 294 243 295
rect 241 294 242 295
rect 240 294 241 295
rect 239 294 240 295
rect 238 294 239 295
rect 237 294 238 295
rect 236 294 237 295
rect 235 294 236 295
rect 234 294 235 295
rect 233 294 234 295
rect 232 294 233 295
rect 231 294 232 295
rect 230 294 231 295
rect 229 294 230 295
rect 228 294 229 295
rect 227 294 228 295
rect 226 294 227 295
rect 225 294 226 295
rect 224 294 225 295
rect 223 294 224 295
rect 222 294 223 295
rect 221 294 222 295
rect 220 294 221 295
rect 219 294 220 295
rect 218 294 219 295
rect 217 294 218 295
rect 216 294 217 295
rect 215 294 216 295
rect 214 294 215 295
rect 213 294 214 295
rect 212 294 213 295
rect 188 294 189 295
rect 187 294 188 295
rect 186 294 187 295
rect 185 294 186 295
rect 184 294 185 295
rect 183 294 184 295
rect 182 294 183 295
rect 181 294 182 295
rect 180 294 181 295
rect 179 294 180 295
rect 178 294 179 295
rect 177 294 178 295
rect 176 294 177 295
rect 175 294 176 295
rect 174 294 175 295
rect 173 294 174 295
rect 172 294 173 295
rect 171 294 172 295
rect 170 294 171 295
rect 169 294 170 295
rect 168 294 169 295
rect 167 294 168 295
rect 166 294 167 295
rect 165 294 166 295
rect 164 294 165 295
rect 163 294 164 295
rect 162 294 163 295
rect 161 294 162 295
rect 160 294 161 295
rect 159 294 160 295
rect 158 294 159 295
rect 157 294 158 295
rect 156 294 157 295
rect 155 294 156 295
rect 154 294 155 295
rect 153 294 154 295
rect 152 294 153 295
rect 151 294 152 295
rect 150 294 151 295
rect 149 294 150 295
rect 148 294 149 295
rect 147 294 148 295
rect 146 294 147 295
rect 145 294 146 295
rect 144 294 145 295
rect 143 294 144 295
rect 142 294 143 295
rect 141 294 142 295
rect 140 294 141 295
rect 139 294 140 295
rect 138 294 139 295
rect 119 294 120 295
rect 118 294 119 295
rect 117 294 118 295
rect 116 294 117 295
rect 115 294 116 295
rect 114 294 115 295
rect 113 294 114 295
rect 112 294 113 295
rect 111 294 112 295
rect 110 294 111 295
rect 109 294 110 295
rect 108 294 109 295
rect 107 294 108 295
rect 106 294 107 295
rect 105 294 106 295
rect 104 294 105 295
rect 103 294 104 295
rect 102 294 103 295
rect 101 294 102 295
rect 100 294 101 295
rect 99 294 100 295
rect 98 294 99 295
rect 97 294 98 295
rect 96 294 97 295
rect 95 294 96 295
rect 94 294 95 295
rect 93 294 94 295
rect 92 294 93 295
rect 91 294 92 295
rect 90 294 91 295
rect 89 294 90 295
rect 88 294 89 295
rect 87 294 88 295
rect 86 294 87 295
rect 85 294 86 295
rect 84 294 85 295
rect 68 294 69 295
rect 67 294 68 295
rect 66 294 67 295
rect 65 294 66 295
rect 64 294 65 295
rect 63 294 64 295
rect 62 294 63 295
rect 61 294 62 295
rect 60 294 61 295
rect 59 294 60 295
rect 58 294 59 295
rect 57 294 58 295
rect 56 294 57 295
rect 55 294 56 295
rect 54 294 55 295
rect 53 294 54 295
rect 52 294 53 295
rect 51 294 52 295
rect 50 294 51 295
rect 49 294 50 295
rect 48 294 49 295
rect 47 294 48 295
rect 46 294 47 295
rect 45 294 46 295
rect 44 294 45 295
rect 43 294 44 295
rect 42 294 43 295
rect 41 294 42 295
rect 40 294 41 295
rect 39 294 40 295
rect 29 294 30 295
rect 28 294 29 295
rect 27 294 28 295
rect 26 294 27 295
rect 25 294 26 295
rect 24 294 25 295
rect 23 294 24 295
rect 22 294 23 295
rect 21 294 22 295
rect 20 294 21 295
rect 19 294 20 295
rect 18 294 19 295
rect 17 294 18 295
rect 16 294 17 295
rect 15 294 16 295
rect 14 294 15 295
rect 13 294 14 295
rect 12 294 13 295
rect 11 294 12 295
rect 10 294 11 295
rect 9 294 10 295
rect 8 294 9 295
rect 7 294 8 295
rect 6 294 7 295
rect 5 294 6 295
rect 4 294 5 295
rect 3 294 4 295
rect 480 295 481 296
rect 479 295 480 296
rect 478 295 479 296
rect 477 295 478 296
rect 476 295 477 296
rect 475 295 476 296
rect 474 295 475 296
rect 473 295 474 296
rect 472 295 473 296
rect 471 295 472 296
rect 470 295 471 296
rect 469 295 470 296
rect 468 295 469 296
rect 467 295 468 296
rect 466 295 467 296
rect 465 295 466 296
rect 464 295 465 296
rect 463 295 464 296
rect 462 295 463 296
rect 461 295 462 296
rect 460 295 461 296
rect 417 295 418 296
rect 416 295 417 296
rect 415 295 416 296
rect 414 295 415 296
rect 275 295 276 296
rect 274 295 275 296
rect 273 295 274 296
rect 272 295 273 296
rect 271 295 272 296
rect 270 295 271 296
rect 269 295 270 296
rect 268 295 269 296
rect 267 295 268 296
rect 266 295 267 296
rect 265 295 266 296
rect 264 295 265 296
rect 263 295 264 296
rect 262 295 263 296
rect 261 295 262 296
rect 260 295 261 296
rect 259 295 260 296
rect 258 295 259 296
rect 257 295 258 296
rect 256 295 257 296
rect 255 295 256 296
rect 254 295 255 296
rect 253 295 254 296
rect 252 295 253 296
rect 251 295 252 296
rect 250 295 251 296
rect 249 295 250 296
rect 248 295 249 296
rect 247 295 248 296
rect 246 295 247 296
rect 245 295 246 296
rect 244 295 245 296
rect 243 295 244 296
rect 242 295 243 296
rect 241 295 242 296
rect 240 295 241 296
rect 239 295 240 296
rect 238 295 239 296
rect 237 295 238 296
rect 236 295 237 296
rect 235 295 236 296
rect 234 295 235 296
rect 233 295 234 296
rect 232 295 233 296
rect 231 295 232 296
rect 230 295 231 296
rect 229 295 230 296
rect 228 295 229 296
rect 227 295 228 296
rect 226 295 227 296
rect 225 295 226 296
rect 224 295 225 296
rect 223 295 224 296
rect 222 295 223 296
rect 221 295 222 296
rect 220 295 221 296
rect 219 295 220 296
rect 218 295 219 296
rect 217 295 218 296
rect 216 295 217 296
rect 215 295 216 296
rect 214 295 215 296
rect 213 295 214 296
rect 212 295 213 296
rect 211 295 212 296
rect 187 295 188 296
rect 186 295 187 296
rect 185 295 186 296
rect 184 295 185 296
rect 183 295 184 296
rect 182 295 183 296
rect 181 295 182 296
rect 180 295 181 296
rect 179 295 180 296
rect 178 295 179 296
rect 177 295 178 296
rect 176 295 177 296
rect 175 295 176 296
rect 174 295 175 296
rect 173 295 174 296
rect 172 295 173 296
rect 171 295 172 296
rect 170 295 171 296
rect 169 295 170 296
rect 168 295 169 296
rect 167 295 168 296
rect 166 295 167 296
rect 165 295 166 296
rect 164 295 165 296
rect 163 295 164 296
rect 162 295 163 296
rect 161 295 162 296
rect 160 295 161 296
rect 159 295 160 296
rect 158 295 159 296
rect 157 295 158 296
rect 156 295 157 296
rect 155 295 156 296
rect 154 295 155 296
rect 153 295 154 296
rect 152 295 153 296
rect 151 295 152 296
rect 150 295 151 296
rect 149 295 150 296
rect 148 295 149 296
rect 147 295 148 296
rect 146 295 147 296
rect 145 295 146 296
rect 144 295 145 296
rect 143 295 144 296
rect 142 295 143 296
rect 141 295 142 296
rect 140 295 141 296
rect 139 295 140 296
rect 120 295 121 296
rect 119 295 120 296
rect 118 295 119 296
rect 117 295 118 296
rect 116 295 117 296
rect 115 295 116 296
rect 114 295 115 296
rect 113 295 114 296
rect 112 295 113 296
rect 111 295 112 296
rect 110 295 111 296
rect 109 295 110 296
rect 108 295 109 296
rect 107 295 108 296
rect 106 295 107 296
rect 105 295 106 296
rect 104 295 105 296
rect 103 295 104 296
rect 102 295 103 296
rect 101 295 102 296
rect 100 295 101 296
rect 99 295 100 296
rect 98 295 99 296
rect 97 295 98 296
rect 96 295 97 296
rect 95 295 96 296
rect 94 295 95 296
rect 93 295 94 296
rect 92 295 93 296
rect 91 295 92 296
rect 90 295 91 296
rect 89 295 90 296
rect 88 295 89 296
rect 87 295 88 296
rect 86 295 87 296
rect 85 295 86 296
rect 84 295 85 296
rect 68 295 69 296
rect 67 295 68 296
rect 66 295 67 296
rect 65 295 66 296
rect 64 295 65 296
rect 63 295 64 296
rect 62 295 63 296
rect 61 295 62 296
rect 60 295 61 296
rect 59 295 60 296
rect 58 295 59 296
rect 57 295 58 296
rect 56 295 57 296
rect 55 295 56 296
rect 54 295 55 296
rect 53 295 54 296
rect 52 295 53 296
rect 51 295 52 296
rect 50 295 51 296
rect 49 295 50 296
rect 48 295 49 296
rect 47 295 48 296
rect 46 295 47 296
rect 45 295 46 296
rect 44 295 45 296
rect 43 295 44 296
rect 42 295 43 296
rect 41 295 42 296
rect 40 295 41 296
rect 39 295 40 296
rect 29 295 30 296
rect 28 295 29 296
rect 27 295 28 296
rect 26 295 27 296
rect 25 295 26 296
rect 24 295 25 296
rect 23 295 24 296
rect 22 295 23 296
rect 21 295 22 296
rect 20 295 21 296
rect 19 295 20 296
rect 18 295 19 296
rect 17 295 18 296
rect 16 295 17 296
rect 15 295 16 296
rect 14 295 15 296
rect 13 295 14 296
rect 12 295 13 296
rect 11 295 12 296
rect 10 295 11 296
rect 9 295 10 296
rect 8 295 9 296
rect 7 295 8 296
rect 6 295 7 296
rect 5 295 6 296
rect 4 295 5 296
rect 3 295 4 296
rect 480 296 481 297
rect 479 296 480 297
rect 478 296 479 297
rect 477 296 478 297
rect 476 296 477 297
rect 475 296 476 297
rect 474 296 475 297
rect 473 296 474 297
rect 472 296 473 297
rect 471 296 472 297
rect 470 296 471 297
rect 469 296 470 297
rect 468 296 469 297
rect 467 296 468 297
rect 466 296 467 297
rect 465 296 466 297
rect 464 296 465 297
rect 463 296 464 297
rect 462 296 463 297
rect 461 296 462 297
rect 460 296 461 297
rect 417 296 418 297
rect 416 296 417 297
rect 415 296 416 297
rect 414 296 415 297
rect 273 296 274 297
rect 272 296 273 297
rect 271 296 272 297
rect 270 296 271 297
rect 269 296 270 297
rect 268 296 269 297
rect 267 296 268 297
rect 266 296 267 297
rect 265 296 266 297
rect 264 296 265 297
rect 263 296 264 297
rect 262 296 263 297
rect 261 296 262 297
rect 260 296 261 297
rect 259 296 260 297
rect 258 296 259 297
rect 257 296 258 297
rect 256 296 257 297
rect 255 296 256 297
rect 254 296 255 297
rect 253 296 254 297
rect 252 296 253 297
rect 251 296 252 297
rect 250 296 251 297
rect 249 296 250 297
rect 248 296 249 297
rect 247 296 248 297
rect 246 296 247 297
rect 245 296 246 297
rect 244 296 245 297
rect 243 296 244 297
rect 242 296 243 297
rect 241 296 242 297
rect 240 296 241 297
rect 239 296 240 297
rect 238 296 239 297
rect 237 296 238 297
rect 236 296 237 297
rect 235 296 236 297
rect 234 296 235 297
rect 233 296 234 297
rect 232 296 233 297
rect 231 296 232 297
rect 230 296 231 297
rect 229 296 230 297
rect 228 296 229 297
rect 227 296 228 297
rect 226 296 227 297
rect 225 296 226 297
rect 224 296 225 297
rect 223 296 224 297
rect 222 296 223 297
rect 221 296 222 297
rect 220 296 221 297
rect 219 296 220 297
rect 218 296 219 297
rect 217 296 218 297
rect 216 296 217 297
rect 215 296 216 297
rect 214 296 215 297
rect 213 296 214 297
rect 212 296 213 297
rect 211 296 212 297
rect 186 296 187 297
rect 185 296 186 297
rect 184 296 185 297
rect 183 296 184 297
rect 182 296 183 297
rect 181 296 182 297
rect 180 296 181 297
rect 179 296 180 297
rect 178 296 179 297
rect 177 296 178 297
rect 176 296 177 297
rect 175 296 176 297
rect 174 296 175 297
rect 173 296 174 297
rect 172 296 173 297
rect 171 296 172 297
rect 170 296 171 297
rect 169 296 170 297
rect 168 296 169 297
rect 167 296 168 297
rect 166 296 167 297
rect 165 296 166 297
rect 164 296 165 297
rect 163 296 164 297
rect 162 296 163 297
rect 161 296 162 297
rect 160 296 161 297
rect 159 296 160 297
rect 158 296 159 297
rect 157 296 158 297
rect 156 296 157 297
rect 155 296 156 297
rect 154 296 155 297
rect 153 296 154 297
rect 152 296 153 297
rect 151 296 152 297
rect 150 296 151 297
rect 149 296 150 297
rect 148 296 149 297
rect 147 296 148 297
rect 146 296 147 297
rect 145 296 146 297
rect 144 296 145 297
rect 143 296 144 297
rect 142 296 143 297
rect 141 296 142 297
rect 140 296 141 297
rect 120 296 121 297
rect 119 296 120 297
rect 118 296 119 297
rect 117 296 118 297
rect 116 296 117 297
rect 115 296 116 297
rect 114 296 115 297
rect 113 296 114 297
rect 112 296 113 297
rect 111 296 112 297
rect 110 296 111 297
rect 109 296 110 297
rect 108 296 109 297
rect 107 296 108 297
rect 106 296 107 297
rect 105 296 106 297
rect 104 296 105 297
rect 103 296 104 297
rect 102 296 103 297
rect 101 296 102 297
rect 100 296 101 297
rect 99 296 100 297
rect 98 296 99 297
rect 97 296 98 297
rect 96 296 97 297
rect 95 296 96 297
rect 94 296 95 297
rect 93 296 94 297
rect 92 296 93 297
rect 91 296 92 297
rect 90 296 91 297
rect 89 296 90 297
rect 88 296 89 297
rect 87 296 88 297
rect 86 296 87 297
rect 85 296 86 297
rect 84 296 85 297
rect 68 296 69 297
rect 67 296 68 297
rect 66 296 67 297
rect 65 296 66 297
rect 64 296 65 297
rect 63 296 64 297
rect 62 296 63 297
rect 61 296 62 297
rect 60 296 61 297
rect 59 296 60 297
rect 58 296 59 297
rect 57 296 58 297
rect 56 296 57 297
rect 55 296 56 297
rect 54 296 55 297
rect 53 296 54 297
rect 52 296 53 297
rect 51 296 52 297
rect 50 296 51 297
rect 49 296 50 297
rect 48 296 49 297
rect 47 296 48 297
rect 46 296 47 297
rect 45 296 46 297
rect 44 296 45 297
rect 43 296 44 297
rect 42 296 43 297
rect 41 296 42 297
rect 40 296 41 297
rect 39 296 40 297
rect 29 296 30 297
rect 28 296 29 297
rect 27 296 28 297
rect 26 296 27 297
rect 25 296 26 297
rect 24 296 25 297
rect 23 296 24 297
rect 22 296 23 297
rect 21 296 22 297
rect 20 296 21 297
rect 19 296 20 297
rect 18 296 19 297
rect 17 296 18 297
rect 16 296 17 297
rect 15 296 16 297
rect 14 296 15 297
rect 13 296 14 297
rect 12 296 13 297
rect 11 296 12 297
rect 10 296 11 297
rect 9 296 10 297
rect 8 296 9 297
rect 7 296 8 297
rect 6 296 7 297
rect 5 296 6 297
rect 4 296 5 297
rect 480 297 481 298
rect 460 297 461 298
rect 417 297 418 298
rect 416 297 417 298
rect 415 297 416 298
rect 414 297 415 298
rect 272 297 273 298
rect 271 297 272 298
rect 270 297 271 298
rect 269 297 270 298
rect 268 297 269 298
rect 267 297 268 298
rect 266 297 267 298
rect 265 297 266 298
rect 264 297 265 298
rect 263 297 264 298
rect 262 297 263 298
rect 261 297 262 298
rect 260 297 261 298
rect 259 297 260 298
rect 258 297 259 298
rect 257 297 258 298
rect 256 297 257 298
rect 255 297 256 298
rect 254 297 255 298
rect 253 297 254 298
rect 252 297 253 298
rect 251 297 252 298
rect 250 297 251 298
rect 249 297 250 298
rect 248 297 249 298
rect 247 297 248 298
rect 246 297 247 298
rect 245 297 246 298
rect 244 297 245 298
rect 243 297 244 298
rect 242 297 243 298
rect 241 297 242 298
rect 240 297 241 298
rect 239 297 240 298
rect 238 297 239 298
rect 237 297 238 298
rect 236 297 237 298
rect 235 297 236 298
rect 234 297 235 298
rect 233 297 234 298
rect 232 297 233 298
rect 231 297 232 298
rect 230 297 231 298
rect 229 297 230 298
rect 228 297 229 298
rect 227 297 228 298
rect 226 297 227 298
rect 225 297 226 298
rect 224 297 225 298
rect 223 297 224 298
rect 222 297 223 298
rect 221 297 222 298
rect 220 297 221 298
rect 219 297 220 298
rect 218 297 219 298
rect 217 297 218 298
rect 216 297 217 298
rect 215 297 216 298
rect 214 297 215 298
rect 213 297 214 298
rect 212 297 213 298
rect 211 297 212 298
rect 210 297 211 298
rect 185 297 186 298
rect 184 297 185 298
rect 183 297 184 298
rect 182 297 183 298
rect 181 297 182 298
rect 180 297 181 298
rect 179 297 180 298
rect 178 297 179 298
rect 177 297 178 298
rect 176 297 177 298
rect 175 297 176 298
rect 174 297 175 298
rect 173 297 174 298
rect 172 297 173 298
rect 171 297 172 298
rect 170 297 171 298
rect 169 297 170 298
rect 168 297 169 298
rect 167 297 168 298
rect 166 297 167 298
rect 165 297 166 298
rect 164 297 165 298
rect 163 297 164 298
rect 162 297 163 298
rect 161 297 162 298
rect 160 297 161 298
rect 159 297 160 298
rect 158 297 159 298
rect 157 297 158 298
rect 156 297 157 298
rect 155 297 156 298
rect 154 297 155 298
rect 153 297 154 298
rect 152 297 153 298
rect 151 297 152 298
rect 150 297 151 298
rect 149 297 150 298
rect 148 297 149 298
rect 147 297 148 298
rect 146 297 147 298
rect 145 297 146 298
rect 144 297 145 298
rect 143 297 144 298
rect 142 297 143 298
rect 141 297 142 298
rect 120 297 121 298
rect 119 297 120 298
rect 118 297 119 298
rect 117 297 118 298
rect 116 297 117 298
rect 115 297 116 298
rect 114 297 115 298
rect 113 297 114 298
rect 112 297 113 298
rect 111 297 112 298
rect 110 297 111 298
rect 109 297 110 298
rect 108 297 109 298
rect 107 297 108 298
rect 106 297 107 298
rect 105 297 106 298
rect 104 297 105 298
rect 103 297 104 298
rect 102 297 103 298
rect 101 297 102 298
rect 100 297 101 298
rect 99 297 100 298
rect 98 297 99 298
rect 97 297 98 298
rect 96 297 97 298
rect 95 297 96 298
rect 94 297 95 298
rect 93 297 94 298
rect 92 297 93 298
rect 91 297 92 298
rect 90 297 91 298
rect 89 297 90 298
rect 88 297 89 298
rect 87 297 88 298
rect 86 297 87 298
rect 85 297 86 298
rect 84 297 85 298
rect 68 297 69 298
rect 67 297 68 298
rect 66 297 67 298
rect 65 297 66 298
rect 64 297 65 298
rect 63 297 64 298
rect 62 297 63 298
rect 61 297 62 298
rect 60 297 61 298
rect 59 297 60 298
rect 58 297 59 298
rect 57 297 58 298
rect 56 297 57 298
rect 55 297 56 298
rect 54 297 55 298
rect 53 297 54 298
rect 52 297 53 298
rect 51 297 52 298
rect 50 297 51 298
rect 49 297 50 298
rect 48 297 49 298
rect 47 297 48 298
rect 46 297 47 298
rect 45 297 46 298
rect 44 297 45 298
rect 43 297 44 298
rect 42 297 43 298
rect 41 297 42 298
rect 40 297 41 298
rect 30 297 31 298
rect 29 297 30 298
rect 28 297 29 298
rect 27 297 28 298
rect 26 297 27 298
rect 25 297 26 298
rect 24 297 25 298
rect 23 297 24 298
rect 22 297 23 298
rect 21 297 22 298
rect 20 297 21 298
rect 19 297 20 298
rect 18 297 19 298
rect 17 297 18 298
rect 16 297 17 298
rect 15 297 16 298
rect 14 297 15 298
rect 13 297 14 298
rect 12 297 13 298
rect 11 297 12 298
rect 10 297 11 298
rect 9 297 10 298
rect 8 297 9 298
rect 7 297 8 298
rect 6 297 7 298
rect 5 297 6 298
rect 4 297 5 298
rect 480 298 481 299
rect 460 298 461 299
rect 417 298 418 299
rect 416 298 417 299
rect 415 298 416 299
rect 414 298 415 299
rect 271 298 272 299
rect 270 298 271 299
rect 269 298 270 299
rect 268 298 269 299
rect 267 298 268 299
rect 266 298 267 299
rect 265 298 266 299
rect 264 298 265 299
rect 263 298 264 299
rect 262 298 263 299
rect 261 298 262 299
rect 260 298 261 299
rect 259 298 260 299
rect 258 298 259 299
rect 257 298 258 299
rect 256 298 257 299
rect 255 298 256 299
rect 254 298 255 299
rect 253 298 254 299
rect 252 298 253 299
rect 251 298 252 299
rect 250 298 251 299
rect 249 298 250 299
rect 248 298 249 299
rect 247 298 248 299
rect 246 298 247 299
rect 245 298 246 299
rect 244 298 245 299
rect 243 298 244 299
rect 242 298 243 299
rect 241 298 242 299
rect 240 298 241 299
rect 239 298 240 299
rect 238 298 239 299
rect 237 298 238 299
rect 236 298 237 299
rect 235 298 236 299
rect 234 298 235 299
rect 233 298 234 299
rect 232 298 233 299
rect 231 298 232 299
rect 230 298 231 299
rect 229 298 230 299
rect 228 298 229 299
rect 227 298 228 299
rect 226 298 227 299
rect 225 298 226 299
rect 224 298 225 299
rect 223 298 224 299
rect 222 298 223 299
rect 221 298 222 299
rect 220 298 221 299
rect 219 298 220 299
rect 218 298 219 299
rect 217 298 218 299
rect 216 298 217 299
rect 215 298 216 299
rect 214 298 215 299
rect 213 298 214 299
rect 212 298 213 299
rect 211 298 212 299
rect 210 298 211 299
rect 209 298 210 299
rect 184 298 185 299
rect 183 298 184 299
rect 182 298 183 299
rect 181 298 182 299
rect 180 298 181 299
rect 179 298 180 299
rect 178 298 179 299
rect 177 298 178 299
rect 176 298 177 299
rect 175 298 176 299
rect 174 298 175 299
rect 173 298 174 299
rect 172 298 173 299
rect 171 298 172 299
rect 170 298 171 299
rect 169 298 170 299
rect 168 298 169 299
rect 167 298 168 299
rect 166 298 167 299
rect 165 298 166 299
rect 164 298 165 299
rect 163 298 164 299
rect 162 298 163 299
rect 161 298 162 299
rect 160 298 161 299
rect 159 298 160 299
rect 158 298 159 299
rect 157 298 158 299
rect 156 298 157 299
rect 155 298 156 299
rect 154 298 155 299
rect 153 298 154 299
rect 152 298 153 299
rect 151 298 152 299
rect 150 298 151 299
rect 149 298 150 299
rect 148 298 149 299
rect 147 298 148 299
rect 146 298 147 299
rect 145 298 146 299
rect 144 298 145 299
rect 143 298 144 299
rect 142 298 143 299
rect 121 298 122 299
rect 120 298 121 299
rect 119 298 120 299
rect 118 298 119 299
rect 117 298 118 299
rect 116 298 117 299
rect 115 298 116 299
rect 114 298 115 299
rect 113 298 114 299
rect 112 298 113 299
rect 111 298 112 299
rect 110 298 111 299
rect 109 298 110 299
rect 108 298 109 299
rect 107 298 108 299
rect 106 298 107 299
rect 105 298 106 299
rect 104 298 105 299
rect 103 298 104 299
rect 102 298 103 299
rect 101 298 102 299
rect 100 298 101 299
rect 99 298 100 299
rect 98 298 99 299
rect 97 298 98 299
rect 96 298 97 299
rect 95 298 96 299
rect 94 298 95 299
rect 93 298 94 299
rect 92 298 93 299
rect 91 298 92 299
rect 90 298 91 299
rect 89 298 90 299
rect 88 298 89 299
rect 87 298 88 299
rect 86 298 87 299
rect 85 298 86 299
rect 68 298 69 299
rect 67 298 68 299
rect 66 298 67 299
rect 65 298 66 299
rect 64 298 65 299
rect 63 298 64 299
rect 62 298 63 299
rect 61 298 62 299
rect 60 298 61 299
rect 59 298 60 299
rect 58 298 59 299
rect 57 298 58 299
rect 56 298 57 299
rect 55 298 56 299
rect 54 298 55 299
rect 53 298 54 299
rect 52 298 53 299
rect 51 298 52 299
rect 50 298 51 299
rect 49 298 50 299
rect 48 298 49 299
rect 47 298 48 299
rect 46 298 47 299
rect 45 298 46 299
rect 44 298 45 299
rect 43 298 44 299
rect 42 298 43 299
rect 41 298 42 299
rect 40 298 41 299
rect 30 298 31 299
rect 29 298 30 299
rect 28 298 29 299
rect 27 298 28 299
rect 26 298 27 299
rect 25 298 26 299
rect 24 298 25 299
rect 23 298 24 299
rect 22 298 23 299
rect 21 298 22 299
rect 20 298 21 299
rect 19 298 20 299
rect 18 298 19 299
rect 17 298 18 299
rect 16 298 17 299
rect 15 298 16 299
rect 14 298 15 299
rect 13 298 14 299
rect 12 298 13 299
rect 11 298 12 299
rect 10 298 11 299
rect 9 298 10 299
rect 8 298 9 299
rect 7 298 8 299
rect 6 298 7 299
rect 5 298 6 299
rect 4 298 5 299
rect 480 299 481 300
rect 460 299 461 300
rect 417 299 418 300
rect 416 299 417 300
rect 415 299 416 300
rect 414 299 415 300
rect 270 299 271 300
rect 269 299 270 300
rect 268 299 269 300
rect 267 299 268 300
rect 266 299 267 300
rect 265 299 266 300
rect 264 299 265 300
rect 263 299 264 300
rect 262 299 263 300
rect 261 299 262 300
rect 260 299 261 300
rect 259 299 260 300
rect 258 299 259 300
rect 257 299 258 300
rect 256 299 257 300
rect 255 299 256 300
rect 254 299 255 300
rect 253 299 254 300
rect 252 299 253 300
rect 251 299 252 300
rect 250 299 251 300
rect 249 299 250 300
rect 248 299 249 300
rect 247 299 248 300
rect 246 299 247 300
rect 245 299 246 300
rect 244 299 245 300
rect 243 299 244 300
rect 242 299 243 300
rect 241 299 242 300
rect 240 299 241 300
rect 239 299 240 300
rect 238 299 239 300
rect 237 299 238 300
rect 236 299 237 300
rect 235 299 236 300
rect 234 299 235 300
rect 233 299 234 300
rect 232 299 233 300
rect 231 299 232 300
rect 230 299 231 300
rect 229 299 230 300
rect 228 299 229 300
rect 227 299 228 300
rect 226 299 227 300
rect 225 299 226 300
rect 224 299 225 300
rect 223 299 224 300
rect 222 299 223 300
rect 221 299 222 300
rect 220 299 221 300
rect 219 299 220 300
rect 218 299 219 300
rect 217 299 218 300
rect 216 299 217 300
rect 215 299 216 300
rect 214 299 215 300
rect 213 299 214 300
rect 212 299 213 300
rect 211 299 212 300
rect 210 299 211 300
rect 209 299 210 300
rect 182 299 183 300
rect 181 299 182 300
rect 180 299 181 300
rect 179 299 180 300
rect 178 299 179 300
rect 177 299 178 300
rect 176 299 177 300
rect 175 299 176 300
rect 174 299 175 300
rect 173 299 174 300
rect 172 299 173 300
rect 171 299 172 300
rect 170 299 171 300
rect 169 299 170 300
rect 168 299 169 300
rect 167 299 168 300
rect 166 299 167 300
rect 165 299 166 300
rect 164 299 165 300
rect 163 299 164 300
rect 162 299 163 300
rect 161 299 162 300
rect 160 299 161 300
rect 159 299 160 300
rect 158 299 159 300
rect 157 299 158 300
rect 156 299 157 300
rect 155 299 156 300
rect 154 299 155 300
rect 153 299 154 300
rect 152 299 153 300
rect 151 299 152 300
rect 150 299 151 300
rect 149 299 150 300
rect 148 299 149 300
rect 147 299 148 300
rect 146 299 147 300
rect 145 299 146 300
rect 144 299 145 300
rect 143 299 144 300
rect 121 299 122 300
rect 120 299 121 300
rect 119 299 120 300
rect 118 299 119 300
rect 117 299 118 300
rect 116 299 117 300
rect 115 299 116 300
rect 114 299 115 300
rect 113 299 114 300
rect 112 299 113 300
rect 111 299 112 300
rect 110 299 111 300
rect 109 299 110 300
rect 108 299 109 300
rect 107 299 108 300
rect 106 299 107 300
rect 105 299 106 300
rect 104 299 105 300
rect 103 299 104 300
rect 102 299 103 300
rect 101 299 102 300
rect 100 299 101 300
rect 99 299 100 300
rect 98 299 99 300
rect 97 299 98 300
rect 96 299 97 300
rect 95 299 96 300
rect 94 299 95 300
rect 93 299 94 300
rect 92 299 93 300
rect 91 299 92 300
rect 90 299 91 300
rect 89 299 90 300
rect 88 299 89 300
rect 87 299 88 300
rect 86 299 87 300
rect 85 299 86 300
rect 69 299 70 300
rect 68 299 69 300
rect 67 299 68 300
rect 66 299 67 300
rect 65 299 66 300
rect 64 299 65 300
rect 63 299 64 300
rect 62 299 63 300
rect 61 299 62 300
rect 60 299 61 300
rect 59 299 60 300
rect 58 299 59 300
rect 57 299 58 300
rect 56 299 57 300
rect 55 299 56 300
rect 54 299 55 300
rect 53 299 54 300
rect 52 299 53 300
rect 51 299 52 300
rect 50 299 51 300
rect 49 299 50 300
rect 48 299 49 300
rect 47 299 48 300
rect 46 299 47 300
rect 45 299 46 300
rect 44 299 45 300
rect 43 299 44 300
rect 42 299 43 300
rect 41 299 42 300
rect 40 299 41 300
rect 30 299 31 300
rect 29 299 30 300
rect 28 299 29 300
rect 27 299 28 300
rect 26 299 27 300
rect 25 299 26 300
rect 24 299 25 300
rect 23 299 24 300
rect 22 299 23 300
rect 21 299 22 300
rect 20 299 21 300
rect 19 299 20 300
rect 18 299 19 300
rect 17 299 18 300
rect 16 299 17 300
rect 15 299 16 300
rect 14 299 15 300
rect 13 299 14 300
rect 12 299 13 300
rect 11 299 12 300
rect 10 299 11 300
rect 9 299 10 300
rect 8 299 9 300
rect 7 299 8 300
rect 6 299 7 300
rect 5 299 6 300
rect 461 300 462 301
rect 460 300 461 301
rect 417 300 418 301
rect 416 300 417 301
rect 415 300 416 301
rect 414 300 415 301
rect 269 300 270 301
rect 268 300 269 301
rect 267 300 268 301
rect 266 300 267 301
rect 265 300 266 301
rect 264 300 265 301
rect 263 300 264 301
rect 262 300 263 301
rect 261 300 262 301
rect 260 300 261 301
rect 259 300 260 301
rect 258 300 259 301
rect 257 300 258 301
rect 256 300 257 301
rect 255 300 256 301
rect 254 300 255 301
rect 253 300 254 301
rect 252 300 253 301
rect 251 300 252 301
rect 250 300 251 301
rect 249 300 250 301
rect 248 300 249 301
rect 247 300 248 301
rect 246 300 247 301
rect 245 300 246 301
rect 244 300 245 301
rect 243 300 244 301
rect 242 300 243 301
rect 241 300 242 301
rect 240 300 241 301
rect 239 300 240 301
rect 238 300 239 301
rect 237 300 238 301
rect 236 300 237 301
rect 235 300 236 301
rect 234 300 235 301
rect 233 300 234 301
rect 232 300 233 301
rect 231 300 232 301
rect 230 300 231 301
rect 229 300 230 301
rect 228 300 229 301
rect 227 300 228 301
rect 226 300 227 301
rect 225 300 226 301
rect 224 300 225 301
rect 223 300 224 301
rect 222 300 223 301
rect 221 300 222 301
rect 220 300 221 301
rect 219 300 220 301
rect 218 300 219 301
rect 217 300 218 301
rect 216 300 217 301
rect 215 300 216 301
rect 214 300 215 301
rect 213 300 214 301
rect 212 300 213 301
rect 211 300 212 301
rect 210 300 211 301
rect 209 300 210 301
rect 208 300 209 301
rect 181 300 182 301
rect 180 300 181 301
rect 179 300 180 301
rect 178 300 179 301
rect 177 300 178 301
rect 176 300 177 301
rect 175 300 176 301
rect 174 300 175 301
rect 173 300 174 301
rect 172 300 173 301
rect 171 300 172 301
rect 170 300 171 301
rect 169 300 170 301
rect 168 300 169 301
rect 167 300 168 301
rect 166 300 167 301
rect 165 300 166 301
rect 164 300 165 301
rect 163 300 164 301
rect 162 300 163 301
rect 161 300 162 301
rect 160 300 161 301
rect 159 300 160 301
rect 158 300 159 301
rect 157 300 158 301
rect 156 300 157 301
rect 155 300 156 301
rect 154 300 155 301
rect 153 300 154 301
rect 152 300 153 301
rect 151 300 152 301
rect 150 300 151 301
rect 149 300 150 301
rect 148 300 149 301
rect 147 300 148 301
rect 146 300 147 301
rect 145 300 146 301
rect 144 300 145 301
rect 121 300 122 301
rect 120 300 121 301
rect 119 300 120 301
rect 118 300 119 301
rect 117 300 118 301
rect 116 300 117 301
rect 115 300 116 301
rect 114 300 115 301
rect 113 300 114 301
rect 112 300 113 301
rect 111 300 112 301
rect 110 300 111 301
rect 109 300 110 301
rect 108 300 109 301
rect 107 300 108 301
rect 106 300 107 301
rect 105 300 106 301
rect 104 300 105 301
rect 103 300 104 301
rect 102 300 103 301
rect 101 300 102 301
rect 100 300 101 301
rect 99 300 100 301
rect 98 300 99 301
rect 97 300 98 301
rect 96 300 97 301
rect 95 300 96 301
rect 94 300 95 301
rect 93 300 94 301
rect 92 300 93 301
rect 91 300 92 301
rect 90 300 91 301
rect 89 300 90 301
rect 88 300 89 301
rect 87 300 88 301
rect 86 300 87 301
rect 85 300 86 301
rect 69 300 70 301
rect 68 300 69 301
rect 67 300 68 301
rect 66 300 67 301
rect 65 300 66 301
rect 64 300 65 301
rect 63 300 64 301
rect 62 300 63 301
rect 61 300 62 301
rect 60 300 61 301
rect 59 300 60 301
rect 58 300 59 301
rect 57 300 58 301
rect 56 300 57 301
rect 55 300 56 301
rect 54 300 55 301
rect 53 300 54 301
rect 52 300 53 301
rect 51 300 52 301
rect 50 300 51 301
rect 49 300 50 301
rect 48 300 49 301
rect 47 300 48 301
rect 46 300 47 301
rect 45 300 46 301
rect 44 300 45 301
rect 43 300 44 301
rect 42 300 43 301
rect 41 300 42 301
rect 40 300 41 301
rect 30 300 31 301
rect 29 300 30 301
rect 28 300 29 301
rect 27 300 28 301
rect 26 300 27 301
rect 25 300 26 301
rect 24 300 25 301
rect 23 300 24 301
rect 22 300 23 301
rect 21 300 22 301
rect 20 300 21 301
rect 19 300 20 301
rect 18 300 19 301
rect 17 300 18 301
rect 16 300 17 301
rect 15 300 16 301
rect 14 300 15 301
rect 13 300 14 301
rect 12 300 13 301
rect 11 300 12 301
rect 10 300 11 301
rect 9 300 10 301
rect 8 300 9 301
rect 7 300 8 301
rect 6 300 7 301
rect 5 300 6 301
rect 462 301 463 302
rect 461 301 462 302
rect 460 301 461 302
rect 417 301 418 302
rect 416 301 417 302
rect 415 301 416 302
rect 414 301 415 302
rect 268 301 269 302
rect 267 301 268 302
rect 266 301 267 302
rect 265 301 266 302
rect 264 301 265 302
rect 263 301 264 302
rect 262 301 263 302
rect 261 301 262 302
rect 260 301 261 302
rect 259 301 260 302
rect 258 301 259 302
rect 257 301 258 302
rect 256 301 257 302
rect 255 301 256 302
rect 254 301 255 302
rect 253 301 254 302
rect 252 301 253 302
rect 251 301 252 302
rect 250 301 251 302
rect 249 301 250 302
rect 248 301 249 302
rect 247 301 248 302
rect 246 301 247 302
rect 245 301 246 302
rect 244 301 245 302
rect 243 301 244 302
rect 242 301 243 302
rect 241 301 242 302
rect 240 301 241 302
rect 239 301 240 302
rect 238 301 239 302
rect 237 301 238 302
rect 236 301 237 302
rect 235 301 236 302
rect 234 301 235 302
rect 233 301 234 302
rect 232 301 233 302
rect 231 301 232 302
rect 230 301 231 302
rect 229 301 230 302
rect 228 301 229 302
rect 227 301 228 302
rect 226 301 227 302
rect 225 301 226 302
rect 224 301 225 302
rect 223 301 224 302
rect 222 301 223 302
rect 221 301 222 302
rect 220 301 221 302
rect 219 301 220 302
rect 218 301 219 302
rect 217 301 218 302
rect 216 301 217 302
rect 215 301 216 302
rect 214 301 215 302
rect 213 301 214 302
rect 212 301 213 302
rect 211 301 212 302
rect 210 301 211 302
rect 209 301 210 302
rect 208 301 209 302
rect 207 301 208 302
rect 180 301 181 302
rect 179 301 180 302
rect 178 301 179 302
rect 177 301 178 302
rect 176 301 177 302
rect 175 301 176 302
rect 174 301 175 302
rect 173 301 174 302
rect 172 301 173 302
rect 171 301 172 302
rect 170 301 171 302
rect 169 301 170 302
rect 168 301 169 302
rect 167 301 168 302
rect 166 301 167 302
rect 165 301 166 302
rect 164 301 165 302
rect 163 301 164 302
rect 162 301 163 302
rect 161 301 162 302
rect 160 301 161 302
rect 159 301 160 302
rect 158 301 159 302
rect 157 301 158 302
rect 156 301 157 302
rect 155 301 156 302
rect 154 301 155 302
rect 153 301 154 302
rect 152 301 153 302
rect 151 301 152 302
rect 150 301 151 302
rect 149 301 150 302
rect 148 301 149 302
rect 147 301 148 302
rect 146 301 147 302
rect 122 301 123 302
rect 121 301 122 302
rect 120 301 121 302
rect 119 301 120 302
rect 118 301 119 302
rect 117 301 118 302
rect 116 301 117 302
rect 115 301 116 302
rect 114 301 115 302
rect 113 301 114 302
rect 112 301 113 302
rect 111 301 112 302
rect 110 301 111 302
rect 109 301 110 302
rect 108 301 109 302
rect 107 301 108 302
rect 106 301 107 302
rect 105 301 106 302
rect 104 301 105 302
rect 103 301 104 302
rect 102 301 103 302
rect 101 301 102 302
rect 100 301 101 302
rect 99 301 100 302
rect 98 301 99 302
rect 97 301 98 302
rect 96 301 97 302
rect 95 301 96 302
rect 94 301 95 302
rect 93 301 94 302
rect 92 301 93 302
rect 91 301 92 302
rect 90 301 91 302
rect 89 301 90 302
rect 88 301 89 302
rect 87 301 88 302
rect 86 301 87 302
rect 85 301 86 302
rect 69 301 70 302
rect 68 301 69 302
rect 67 301 68 302
rect 66 301 67 302
rect 65 301 66 302
rect 64 301 65 302
rect 63 301 64 302
rect 62 301 63 302
rect 61 301 62 302
rect 60 301 61 302
rect 59 301 60 302
rect 58 301 59 302
rect 57 301 58 302
rect 56 301 57 302
rect 55 301 56 302
rect 54 301 55 302
rect 53 301 54 302
rect 52 301 53 302
rect 51 301 52 302
rect 50 301 51 302
rect 49 301 50 302
rect 48 301 49 302
rect 47 301 48 302
rect 46 301 47 302
rect 45 301 46 302
rect 44 301 45 302
rect 43 301 44 302
rect 42 301 43 302
rect 41 301 42 302
rect 30 301 31 302
rect 29 301 30 302
rect 28 301 29 302
rect 27 301 28 302
rect 26 301 27 302
rect 25 301 26 302
rect 24 301 25 302
rect 23 301 24 302
rect 22 301 23 302
rect 21 301 22 302
rect 20 301 21 302
rect 19 301 20 302
rect 18 301 19 302
rect 17 301 18 302
rect 16 301 17 302
rect 15 301 16 302
rect 14 301 15 302
rect 13 301 14 302
rect 12 301 13 302
rect 11 301 12 302
rect 10 301 11 302
rect 9 301 10 302
rect 8 301 9 302
rect 7 301 8 302
rect 6 301 7 302
rect 5 301 6 302
rect 464 302 465 303
rect 463 302 464 303
rect 462 302 463 303
rect 461 302 462 303
rect 460 302 461 303
rect 459 302 460 303
rect 439 302 440 303
rect 438 302 439 303
rect 417 302 418 303
rect 416 302 417 303
rect 415 302 416 303
rect 414 302 415 303
rect 396 302 397 303
rect 395 302 396 303
rect 266 302 267 303
rect 265 302 266 303
rect 264 302 265 303
rect 263 302 264 303
rect 262 302 263 303
rect 261 302 262 303
rect 260 302 261 303
rect 259 302 260 303
rect 258 302 259 303
rect 257 302 258 303
rect 256 302 257 303
rect 255 302 256 303
rect 254 302 255 303
rect 253 302 254 303
rect 252 302 253 303
rect 251 302 252 303
rect 250 302 251 303
rect 249 302 250 303
rect 248 302 249 303
rect 247 302 248 303
rect 246 302 247 303
rect 245 302 246 303
rect 244 302 245 303
rect 243 302 244 303
rect 242 302 243 303
rect 241 302 242 303
rect 240 302 241 303
rect 239 302 240 303
rect 238 302 239 303
rect 237 302 238 303
rect 236 302 237 303
rect 235 302 236 303
rect 234 302 235 303
rect 233 302 234 303
rect 232 302 233 303
rect 231 302 232 303
rect 230 302 231 303
rect 229 302 230 303
rect 228 302 229 303
rect 227 302 228 303
rect 226 302 227 303
rect 225 302 226 303
rect 224 302 225 303
rect 223 302 224 303
rect 222 302 223 303
rect 221 302 222 303
rect 220 302 221 303
rect 219 302 220 303
rect 218 302 219 303
rect 217 302 218 303
rect 216 302 217 303
rect 215 302 216 303
rect 214 302 215 303
rect 213 302 214 303
rect 212 302 213 303
rect 211 302 212 303
rect 210 302 211 303
rect 209 302 210 303
rect 208 302 209 303
rect 207 302 208 303
rect 178 302 179 303
rect 177 302 178 303
rect 176 302 177 303
rect 175 302 176 303
rect 174 302 175 303
rect 173 302 174 303
rect 172 302 173 303
rect 171 302 172 303
rect 170 302 171 303
rect 169 302 170 303
rect 168 302 169 303
rect 167 302 168 303
rect 166 302 167 303
rect 165 302 166 303
rect 164 302 165 303
rect 163 302 164 303
rect 162 302 163 303
rect 161 302 162 303
rect 160 302 161 303
rect 159 302 160 303
rect 158 302 159 303
rect 157 302 158 303
rect 156 302 157 303
rect 155 302 156 303
rect 154 302 155 303
rect 153 302 154 303
rect 152 302 153 303
rect 151 302 152 303
rect 150 302 151 303
rect 149 302 150 303
rect 148 302 149 303
rect 147 302 148 303
rect 122 302 123 303
rect 121 302 122 303
rect 120 302 121 303
rect 119 302 120 303
rect 118 302 119 303
rect 117 302 118 303
rect 116 302 117 303
rect 115 302 116 303
rect 114 302 115 303
rect 113 302 114 303
rect 112 302 113 303
rect 111 302 112 303
rect 110 302 111 303
rect 109 302 110 303
rect 108 302 109 303
rect 107 302 108 303
rect 106 302 107 303
rect 105 302 106 303
rect 104 302 105 303
rect 103 302 104 303
rect 102 302 103 303
rect 101 302 102 303
rect 100 302 101 303
rect 99 302 100 303
rect 98 302 99 303
rect 97 302 98 303
rect 96 302 97 303
rect 95 302 96 303
rect 94 302 95 303
rect 93 302 94 303
rect 92 302 93 303
rect 91 302 92 303
rect 90 302 91 303
rect 89 302 90 303
rect 88 302 89 303
rect 87 302 88 303
rect 86 302 87 303
rect 69 302 70 303
rect 68 302 69 303
rect 67 302 68 303
rect 66 302 67 303
rect 65 302 66 303
rect 64 302 65 303
rect 63 302 64 303
rect 62 302 63 303
rect 61 302 62 303
rect 60 302 61 303
rect 59 302 60 303
rect 58 302 59 303
rect 57 302 58 303
rect 56 302 57 303
rect 55 302 56 303
rect 54 302 55 303
rect 53 302 54 303
rect 52 302 53 303
rect 51 302 52 303
rect 50 302 51 303
rect 49 302 50 303
rect 48 302 49 303
rect 47 302 48 303
rect 46 302 47 303
rect 45 302 46 303
rect 44 302 45 303
rect 43 302 44 303
rect 42 302 43 303
rect 41 302 42 303
rect 30 302 31 303
rect 29 302 30 303
rect 28 302 29 303
rect 27 302 28 303
rect 26 302 27 303
rect 25 302 26 303
rect 24 302 25 303
rect 23 302 24 303
rect 22 302 23 303
rect 21 302 22 303
rect 20 302 21 303
rect 19 302 20 303
rect 18 302 19 303
rect 17 302 18 303
rect 16 302 17 303
rect 15 302 16 303
rect 14 302 15 303
rect 13 302 14 303
rect 12 302 13 303
rect 11 302 12 303
rect 10 302 11 303
rect 9 302 10 303
rect 8 302 9 303
rect 7 302 8 303
rect 6 302 7 303
rect 464 303 465 304
rect 463 303 464 304
rect 462 303 463 304
rect 461 303 462 304
rect 460 303 461 304
rect 459 303 460 304
rect 439 303 440 304
rect 438 303 439 304
rect 437 303 438 304
rect 417 303 418 304
rect 416 303 417 304
rect 415 303 416 304
rect 414 303 415 304
rect 397 303 398 304
rect 396 303 397 304
rect 395 303 396 304
rect 265 303 266 304
rect 264 303 265 304
rect 263 303 264 304
rect 262 303 263 304
rect 261 303 262 304
rect 260 303 261 304
rect 259 303 260 304
rect 258 303 259 304
rect 257 303 258 304
rect 256 303 257 304
rect 255 303 256 304
rect 254 303 255 304
rect 253 303 254 304
rect 252 303 253 304
rect 251 303 252 304
rect 250 303 251 304
rect 249 303 250 304
rect 248 303 249 304
rect 247 303 248 304
rect 246 303 247 304
rect 245 303 246 304
rect 244 303 245 304
rect 243 303 244 304
rect 242 303 243 304
rect 241 303 242 304
rect 240 303 241 304
rect 239 303 240 304
rect 238 303 239 304
rect 237 303 238 304
rect 236 303 237 304
rect 235 303 236 304
rect 234 303 235 304
rect 233 303 234 304
rect 232 303 233 304
rect 231 303 232 304
rect 230 303 231 304
rect 229 303 230 304
rect 228 303 229 304
rect 227 303 228 304
rect 226 303 227 304
rect 225 303 226 304
rect 224 303 225 304
rect 223 303 224 304
rect 222 303 223 304
rect 221 303 222 304
rect 220 303 221 304
rect 219 303 220 304
rect 218 303 219 304
rect 217 303 218 304
rect 216 303 217 304
rect 215 303 216 304
rect 214 303 215 304
rect 213 303 214 304
rect 212 303 213 304
rect 211 303 212 304
rect 210 303 211 304
rect 209 303 210 304
rect 208 303 209 304
rect 207 303 208 304
rect 206 303 207 304
rect 177 303 178 304
rect 176 303 177 304
rect 175 303 176 304
rect 174 303 175 304
rect 173 303 174 304
rect 172 303 173 304
rect 171 303 172 304
rect 170 303 171 304
rect 169 303 170 304
rect 168 303 169 304
rect 167 303 168 304
rect 166 303 167 304
rect 165 303 166 304
rect 164 303 165 304
rect 163 303 164 304
rect 162 303 163 304
rect 161 303 162 304
rect 160 303 161 304
rect 159 303 160 304
rect 158 303 159 304
rect 157 303 158 304
rect 156 303 157 304
rect 155 303 156 304
rect 154 303 155 304
rect 153 303 154 304
rect 152 303 153 304
rect 151 303 152 304
rect 150 303 151 304
rect 149 303 150 304
rect 123 303 124 304
rect 122 303 123 304
rect 121 303 122 304
rect 120 303 121 304
rect 119 303 120 304
rect 118 303 119 304
rect 117 303 118 304
rect 116 303 117 304
rect 115 303 116 304
rect 114 303 115 304
rect 113 303 114 304
rect 112 303 113 304
rect 111 303 112 304
rect 110 303 111 304
rect 109 303 110 304
rect 108 303 109 304
rect 107 303 108 304
rect 106 303 107 304
rect 105 303 106 304
rect 104 303 105 304
rect 103 303 104 304
rect 102 303 103 304
rect 101 303 102 304
rect 100 303 101 304
rect 99 303 100 304
rect 98 303 99 304
rect 97 303 98 304
rect 96 303 97 304
rect 95 303 96 304
rect 94 303 95 304
rect 93 303 94 304
rect 92 303 93 304
rect 91 303 92 304
rect 90 303 91 304
rect 89 303 90 304
rect 88 303 89 304
rect 87 303 88 304
rect 86 303 87 304
rect 70 303 71 304
rect 69 303 70 304
rect 68 303 69 304
rect 67 303 68 304
rect 66 303 67 304
rect 65 303 66 304
rect 64 303 65 304
rect 63 303 64 304
rect 62 303 63 304
rect 61 303 62 304
rect 60 303 61 304
rect 59 303 60 304
rect 58 303 59 304
rect 57 303 58 304
rect 56 303 57 304
rect 55 303 56 304
rect 54 303 55 304
rect 53 303 54 304
rect 52 303 53 304
rect 51 303 52 304
rect 50 303 51 304
rect 49 303 50 304
rect 48 303 49 304
rect 47 303 48 304
rect 46 303 47 304
rect 45 303 46 304
rect 44 303 45 304
rect 43 303 44 304
rect 42 303 43 304
rect 41 303 42 304
rect 31 303 32 304
rect 30 303 31 304
rect 29 303 30 304
rect 28 303 29 304
rect 27 303 28 304
rect 26 303 27 304
rect 25 303 26 304
rect 24 303 25 304
rect 23 303 24 304
rect 22 303 23 304
rect 21 303 22 304
rect 20 303 21 304
rect 19 303 20 304
rect 18 303 19 304
rect 17 303 18 304
rect 16 303 17 304
rect 15 303 16 304
rect 14 303 15 304
rect 13 303 14 304
rect 12 303 13 304
rect 11 303 12 304
rect 10 303 11 304
rect 9 303 10 304
rect 8 303 9 304
rect 7 303 8 304
rect 6 303 7 304
rect 439 304 440 305
rect 438 304 439 305
rect 437 304 438 305
rect 417 304 418 305
rect 416 304 417 305
rect 415 304 416 305
rect 414 304 415 305
rect 397 304 398 305
rect 396 304 397 305
rect 395 304 396 305
rect 264 304 265 305
rect 263 304 264 305
rect 262 304 263 305
rect 261 304 262 305
rect 260 304 261 305
rect 259 304 260 305
rect 258 304 259 305
rect 257 304 258 305
rect 256 304 257 305
rect 255 304 256 305
rect 254 304 255 305
rect 253 304 254 305
rect 252 304 253 305
rect 251 304 252 305
rect 250 304 251 305
rect 249 304 250 305
rect 248 304 249 305
rect 247 304 248 305
rect 246 304 247 305
rect 245 304 246 305
rect 244 304 245 305
rect 243 304 244 305
rect 242 304 243 305
rect 241 304 242 305
rect 240 304 241 305
rect 239 304 240 305
rect 238 304 239 305
rect 237 304 238 305
rect 236 304 237 305
rect 235 304 236 305
rect 234 304 235 305
rect 233 304 234 305
rect 232 304 233 305
rect 231 304 232 305
rect 230 304 231 305
rect 229 304 230 305
rect 228 304 229 305
rect 227 304 228 305
rect 226 304 227 305
rect 225 304 226 305
rect 224 304 225 305
rect 223 304 224 305
rect 222 304 223 305
rect 221 304 222 305
rect 220 304 221 305
rect 219 304 220 305
rect 218 304 219 305
rect 217 304 218 305
rect 216 304 217 305
rect 215 304 216 305
rect 214 304 215 305
rect 213 304 214 305
rect 212 304 213 305
rect 211 304 212 305
rect 210 304 211 305
rect 209 304 210 305
rect 208 304 209 305
rect 207 304 208 305
rect 206 304 207 305
rect 205 304 206 305
rect 175 304 176 305
rect 174 304 175 305
rect 173 304 174 305
rect 172 304 173 305
rect 171 304 172 305
rect 170 304 171 305
rect 169 304 170 305
rect 168 304 169 305
rect 167 304 168 305
rect 166 304 167 305
rect 165 304 166 305
rect 164 304 165 305
rect 163 304 164 305
rect 162 304 163 305
rect 161 304 162 305
rect 160 304 161 305
rect 159 304 160 305
rect 158 304 159 305
rect 157 304 158 305
rect 156 304 157 305
rect 155 304 156 305
rect 154 304 155 305
rect 153 304 154 305
rect 152 304 153 305
rect 151 304 152 305
rect 123 304 124 305
rect 122 304 123 305
rect 121 304 122 305
rect 120 304 121 305
rect 119 304 120 305
rect 118 304 119 305
rect 117 304 118 305
rect 116 304 117 305
rect 115 304 116 305
rect 114 304 115 305
rect 113 304 114 305
rect 112 304 113 305
rect 111 304 112 305
rect 110 304 111 305
rect 109 304 110 305
rect 108 304 109 305
rect 107 304 108 305
rect 106 304 107 305
rect 105 304 106 305
rect 104 304 105 305
rect 103 304 104 305
rect 102 304 103 305
rect 101 304 102 305
rect 100 304 101 305
rect 99 304 100 305
rect 98 304 99 305
rect 97 304 98 305
rect 96 304 97 305
rect 95 304 96 305
rect 94 304 95 305
rect 93 304 94 305
rect 92 304 93 305
rect 91 304 92 305
rect 90 304 91 305
rect 89 304 90 305
rect 88 304 89 305
rect 87 304 88 305
rect 86 304 87 305
rect 70 304 71 305
rect 69 304 70 305
rect 68 304 69 305
rect 67 304 68 305
rect 66 304 67 305
rect 65 304 66 305
rect 64 304 65 305
rect 63 304 64 305
rect 62 304 63 305
rect 61 304 62 305
rect 60 304 61 305
rect 59 304 60 305
rect 58 304 59 305
rect 57 304 58 305
rect 56 304 57 305
rect 55 304 56 305
rect 54 304 55 305
rect 53 304 54 305
rect 52 304 53 305
rect 51 304 52 305
rect 50 304 51 305
rect 49 304 50 305
rect 48 304 49 305
rect 47 304 48 305
rect 46 304 47 305
rect 45 304 46 305
rect 44 304 45 305
rect 43 304 44 305
rect 42 304 43 305
rect 31 304 32 305
rect 30 304 31 305
rect 29 304 30 305
rect 28 304 29 305
rect 27 304 28 305
rect 26 304 27 305
rect 25 304 26 305
rect 24 304 25 305
rect 23 304 24 305
rect 22 304 23 305
rect 21 304 22 305
rect 20 304 21 305
rect 19 304 20 305
rect 18 304 19 305
rect 17 304 18 305
rect 16 304 17 305
rect 15 304 16 305
rect 14 304 15 305
rect 13 304 14 305
rect 12 304 13 305
rect 11 304 12 305
rect 10 304 11 305
rect 9 304 10 305
rect 8 304 9 305
rect 7 304 8 305
rect 439 305 440 306
rect 438 305 439 306
rect 437 305 438 306
rect 417 305 418 306
rect 416 305 417 306
rect 415 305 416 306
rect 414 305 415 306
rect 397 305 398 306
rect 396 305 397 306
rect 395 305 396 306
rect 262 305 263 306
rect 261 305 262 306
rect 260 305 261 306
rect 259 305 260 306
rect 258 305 259 306
rect 257 305 258 306
rect 256 305 257 306
rect 255 305 256 306
rect 254 305 255 306
rect 253 305 254 306
rect 252 305 253 306
rect 251 305 252 306
rect 250 305 251 306
rect 249 305 250 306
rect 248 305 249 306
rect 247 305 248 306
rect 246 305 247 306
rect 245 305 246 306
rect 244 305 245 306
rect 243 305 244 306
rect 242 305 243 306
rect 241 305 242 306
rect 240 305 241 306
rect 239 305 240 306
rect 238 305 239 306
rect 237 305 238 306
rect 236 305 237 306
rect 235 305 236 306
rect 234 305 235 306
rect 233 305 234 306
rect 232 305 233 306
rect 231 305 232 306
rect 230 305 231 306
rect 229 305 230 306
rect 228 305 229 306
rect 227 305 228 306
rect 226 305 227 306
rect 225 305 226 306
rect 224 305 225 306
rect 223 305 224 306
rect 222 305 223 306
rect 221 305 222 306
rect 220 305 221 306
rect 219 305 220 306
rect 218 305 219 306
rect 217 305 218 306
rect 216 305 217 306
rect 215 305 216 306
rect 214 305 215 306
rect 213 305 214 306
rect 212 305 213 306
rect 211 305 212 306
rect 210 305 211 306
rect 209 305 210 306
rect 208 305 209 306
rect 207 305 208 306
rect 206 305 207 306
rect 205 305 206 306
rect 204 305 205 306
rect 173 305 174 306
rect 172 305 173 306
rect 171 305 172 306
rect 170 305 171 306
rect 169 305 170 306
rect 168 305 169 306
rect 167 305 168 306
rect 166 305 167 306
rect 165 305 166 306
rect 164 305 165 306
rect 163 305 164 306
rect 162 305 163 306
rect 161 305 162 306
rect 160 305 161 306
rect 159 305 160 306
rect 158 305 159 306
rect 157 305 158 306
rect 156 305 157 306
rect 155 305 156 306
rect 154 305 155 306
rect 153 305 154 306
rect 124 305 125 306
rect 123 305 124 306
rect 122 305 123 306
rect 121 305 122 306
rect 120 305 121 306
rect 119 305 120 306
rect 118 305 119 306
rect 117 305 118 306
rect 116 305 117 306
rect 115 305 116 306
rect 114 305 115 306
rect 113 305 114 306
rect 112 305 113 306
rect 111 305 112 306
rect 110 305 111 306
rect 109 305 110 306
rect 108 305 109 306
rect 107 305 108 306
rect 106 305 107 306
rect 105 305 106 306
rect 104 305 105 306
rect 103 305 104 306
rect 102 305 103 306
rect 101 305 102 306
rect 100 305 101 306
rect 99 305 100 306
rect 98 305 99 306
rect 97 305 98 306
rect 96 305 97 306
rect 95 305 96 306
rect 94 305 95 306
rect 93 305 94 306
rect 92 305 93 306
rect 91 305 92 306
rect 90 305 91 306
rect 89 305 90 306
rect 88 305 89 306
rect 87 305 88 306
rect 70 305 71 306
rect 69 305 70 306
rect 68 305 69 306
rect 67 305 68 306
rect 66 305 67 306
rect 65 305 66 306
rect 64 305 65 306
rect 63 305 64 306
rect 62 305 63 306
rect 61 305 62 306
rect 60 305 61 306
rect 59 305 60 306
rect 58 305 59 306
rect 57 305 58 306
rect 56 305 57 306
rect 55 305 56 306
rect 54 305 55 306
rect 53 305 54 306
rect 52 305 53 306
rect 51 305 52 306
rect 50 305 51 306
rect 49 305 50 306
rect 48 305 49 306
rect 47 305 48 306
rect 46 305 47 306
rect 45 305 46 306
rect 44 305 45 306
rect 43 305 44 306
rect 42 305 43 306
rect 31 305 32 306
rect 30 305 31 306
rect 29 305 30 306
rect 28 305 29 306
rect 27 305 28 306
rect 26 305 27 306
rect 25 305 26 306
rect 24 305 25 306
rect 23 305 24 306
rect 22 305 23 306
rect 21 305 22 306
rect 20 305 21 306
rect 19 305 20 306
rect 18 305 19 306
rect 17 305 18 306
rect 16 305 17 306
rect 15 305 16 306
rect 14 305 15 306
rect 13 305 14 306
rect 12 305 13 306
rect 11 305 12 306
rect 10 305 11 306
rect 9 305 10 306
rect 8 305 9 306
rect 7 305 8 306
rect 439 306 440 307
rect 438 306 439 307
rect 437 306 438 307
rect 417 306 418 307
rect 416 306 417 307
rect 415 306 416 307
rect 414 306 415 307
rect 397 306 398 307
rect 396 306 397 307
rect 395 306 396 307
rect 261 306 262 307
rect 260 306 261 307
rect 259 306 260 307
rect 258 306 259 307
rect 257 306 258 307
rect 256 306 257 307
rect 255 306 256 307
rect 254 306 255 307
rect 253 306 254 307
rect 252 306 253 307
rect 251 306 252 307
rect 250 306 251 307
rect 249 306 250 307
rect 248 306 249 307
rect 247 306 248 307
rect 246 306 247 307
rect 245 306 246 307
rect 244 306 245 307
rect 243 306 244 307
rect 242 306 243 307
rect 241 306 242 307
rect 240 306 241 307
rect 239 306 240 307
rect 238 306 239 307
rect 237 306 238 307
rect 236 306 237 307
rect 235 306 236 307
rect 234 306 235 307
rect 233 306 234 307
rect 232 306 233 307
rect 231 306 232 307
rect 230 306 231 307
rect 229 306 230 307
rect 228 306 229 307
rect 227 306 228 307
rect 226 306 227 307
rect 225 306 226 307
rect 224 306 225 307
rect 223 306 224 307
rect 222 306 223 307
rect 221 306 222 307
rect 220 306 221 307
rect 219 306 220 307
rect 218 306 219 307
rect 217 306 218 307
rect 216 306 217 307
rect 215 306 216 307
rect 214 306 215 307
rect 213 306 214 307
rect 212 306 213 307
rect 211 306 212 307
rect 210 306 211 307
rect 209 306 210 307
rect 208 306 209 307
rect 207 306 208 307
rect 206 306 207 307
rect 205 306 206 307
rect 204 306 205 307
rect 203 306 204 307
rect 170 306 171 307
rect 169 306 170 307
rect 168 306 169 307
rect 167 306 168 307
rect 166 306 167 307
rect 165 306 166 307
rect 164 306 165 307
rect 163 306 164 307
rect 162 306 163 307
rect 161 306 162 307
rect 160 306 161 307
rect 159 306 160 307
rect 158 306 159 307
rect 157 306 158 307
rect 156 306 157 307
rect 125 306 126 307
rect 124 306 125 307
rect 123 306 124 307
rect 122 306 123 307
rect 121 306 122 307
rect 120 306 121 307
rect 119 306 120 307
rect 118 306 119 307
rect 117 306 118 307
rect 116 306 117 307
rect 115 306 116 307
rect 114 306 115 307
rect 113 306 114 307
rect 112 306 113 307
rect 111 306 112 307
rect 110 306 111 307
rect 109 306 110 307
rect 108 306 109 307
rect 107 306 108 307
rect 106 306 107 307
rect 105 306 106 307
rect 104 306 105 307
rect 103 306 104 307
rect 102 306 103 307
rect 101 306 102 307
rect 100 306 101 307
rect 99 306 100 307
rect 98 306 99 307
rect 97 306 98 307
rect 96 306 97 307
rect 95 306 96 307
rect 94 306 95 307
rect 93 306 94 307
rect 92 306 93 307
rect 91 306 92 307
rect 90 306 91 307
rect 89 306 90 307
rect 88 306 89 307
rect 87 306 88 307
rect 71 306 72 307
rect 70 306 71 307
rect 69 306 70 307
rect 68 306 69 307
rect 67 306 68 307
rect 66 306 67 307
rect 65 306 66 307
rect 64 306 65 307
rect 63 306 64 307
rect 62 306 63 307
rect 61 306 62 307
rect 60 306 61 307
rect 59 306 60 307
rect 58 306 59 307
rect 57 306 58 307
rect 56 306 57 307
rect 55 306 56 307
rect 54 306 55 307
rect 53 306 54 307
rect 52 306 53 307
rect 51 306 52 307
rect 50 306 51 307
rect 49 306 50 307
rect 48 306 49 307
rect 47 306 48 307
rect 46 306 47 307
rect 45 306 46 307
rect 44 306 45 307
rect 43 306 44 307
rect 42 306 43 307
rect 31 306 32 307
rect 30 306 31 307
rect 29 306 30 307
rect 28 306 29 307
rect 27 306 28 307
rect 26 306 27 307
rect 25 306 26 307
rect 24 306 25 307
rect 23 306 24 307
rect 22 306 23 307
rect 21 306 22 307
rect 20 306 21 307
rect 19 306 20 307
rect 18 306 19 307
rect 17 306 18 307
rect 16 306 17 307
rect 15 306 16 307
rect 14 306 15 307
rect 13 306 14 307
rect 12 306 13 307
rect 11 306 12 307
rect 10 306 11 307
rect 9 306 10 307
rect 8 306 9 307
rect 439 307 440 308
rect 438 307 439 308
rect 437 307 438 308
rect 436 307 437 308
rect 417 307 418 308
rect 416 307 417 308
rect 415 307 416 308
rect 414 307 415 308
rect 399 307 400 308
rect 398 307 399 308
rect 397 307 398 308
rect 396 307 397 308
rect 395 307 396 308
rect 259 307 260 308
rect 258 307 259 308
rect 257 307 258 308
rect 256 307 257 308
rect 255 307 256 308
rect 254 307 255 308
rect 253 307 254 308
rect 252 307 253 308
rect 251 307 252 308
rect 250 307 251 308
rect 249 307 250 308
rect 248 307 249 308
rect 247 307 248 308
rect 246 307 247 308
rect 245 307 246 308
rect 244 307 245 308
rect 243 307 244 308
rect 242 307 243 308
rect 241 307 242 308
rect 240 307 241 308
rect 239 307 240 308
rect 238 307 239 308
rect 237 307 238 308
rect 236 307 237 308
rect 235 307 236 308
rect 234 307 235 308
rect 233 307 234 308
rect 232 307 233 308
rect 231 307 232 308
rect 230 307 231 308
rect 229 307 230 308
rect 228 307 229 308
rect 227 307 228 308
rect 226 307 227 308
rect 225 307 226 308
rect 224 307 225 308
rect 223 307 224 308
rect 222 307 223 308
rect 221 307 222 308
rect 220 307 221 308
rect 219 307 220 308
rect 218 307 219 308
rect 217 307 218 308
rect 216 307 217 308
rect 215 307 216 308
rect 214 307 215 308
rect 213 307 214 308
rect 212 307 213 308
rect 211 307 212 308
rect 210 307 211 308
rect 209 307 210 308
rect 208 307 209 308
rect 207 307 208 308
rect 206 307 207 308
rect 205 307 206 308
rect 204 307 205 308
rect 203 307 204 308
rect 164 307 165 308
rect 163 307 164 308
rect 162 307 163 308
rect 125 307 126 308
rect 124 307 125 308
rect 123 307 124 308
rect 122 307 123 308
rect 121 307 122 308
rect 120 307 121 308
rect 119 307 120 308
rect 118 307 119 308
rect 117 307 118 308
rect 116 307 117 308
rect 115 307 116 308
rect 114 307 115 308
rect 113 307 114 308
rect 112 307 113 308
rect 111 307 112 308
rect 110 307 111 308
rect 109 307 110 308
rect 108 307 109 308
rect 107 307 108 308
rect 106 307 107 308
rect 105 307 106 308
rect 104 307 105 308
rect 103 307 104 308
rect 102 307 103 308
rect 101 307 102 308
rect 100 307 101 308
rect 99 307 100 308
rect 98 307 99 308
rect 97 307 98 308
rect 96 307 97 308
rect 95 307 96 308
rect 94 307 95 308
rect 93 307 94 308
rect 92 307 93 308
rect 91 307 92 308
rect 90 307 91 308
rect 89 307 90 308
rect 88 307 89 308
rect 71 307 72 308
rect 70 307 71 308
rect 69 307 70 308
rect 68 307 69 308
rect 67 307 68 308
rect 66 307 67 308
rect 65 307 66 308
rect 64 307 65 308
rect 63 307 64 308
rect 62 307 63 308
rect 61 307 62 308
rect 60 307 61 308
rect 59 307 60 308
rect 58 307 59 308
rect 57 307 58 308
rect 56 307 57 308
rect 55 307 56 308
rect 54 307 55 308
rect 53 307 54 308
rect 52 307 53 308
rect 51 307 52 308
rect 50 307 51 308
rect 49 307 50 308
rect 48 307 49 308
rect 47 307 48 308
rect 46 307 47 308
rect 45 307 46 308
rect 44 307 45 308
rect 43 307 44 308
rect 32 307 33 308
rect 31 307 32 308
rect 30 307 31 308
rect 29 307 30 308
rect 28 307 29 308
rect 27 307 28 308
rect 26 307 27 308
rect 25 307 26 308
rect 24 307 25 308
rect 23 307 24 308
rect 22 307 23 308
rect 21 307 22 308
rect 20 307 21 308
rect 19 307 20 308
rect 18 307 19 308
rect 17 307 18 308
rect 16 307 17 308
rect 15 307 16 308
rect 14 307 15 308
rect 13 307 14 308
rect 12 307 13 308
rect 11 307 12 308
rect 10 307 11 308
rect 9 307 10 308
rect 8 307 9 308
rect 439 308 440 309
rect 438 308 439 309
rect 437 308 438 309
rect 436 308 437 309
rect 435 308 436 309
rect 434 308 435 309
rect 433 308 434 309
rect 432 308 433 309
rect 431 308 432 309
rect 430 308 431 309
rect 429 308 430 309
rect 428 308 429 309
rect 427 308 428 309
rect 426 308 427 309
rect 425 308 426 309
rect 424 308 425 309
rect 423 308 424 309
rect 422 308 423 309
rect 421 308 422 309
rect 420 308 421 309
rect 419 308 420 309
rect 418 308 419 309
rect 417 308 418 309
rect 416 308 417 309
rect 415 308 416 309
rect 414 308 415 309
rect 413 308 414 309
rect 412 308 413 309
rect 411 308 412 309
rect 410 308 411 309
rect 409 308 410 309
rect 408 308 409 309
rect 407 308 408 309
rect 406 308 407 309
rect 405 308 406 309
rect 404 308 405 309
rect 403 308 404 309
rect 402 308 403 309
rect 401 308 402 309
rect 400 308 401 309
rect 399 308 400 309
rect 398 308 399 309
rect 397 308 398 309
rect 396 308 397 309
rect 395 308 396 309
rect 258 308 259 309
rect 257 308 258 309
rect 256 308 257 309
rect 255 308 256 309
rect 254 308 255 309
rect 253 308 254 309
rect 252 308 253 309
rect 251 308 252 309
rect 250 308 251 309
rect 249 308 250 309
rect 248 308 249 309
rect 247 308 248 309
rect 246 308 247 309
rect 245 308 246 309
rect 244 308 245 309
rect 243 308 244 309
rect 242 308 243 309
rect 241 308 242 309
rect 240 308 241 309
rect 239 308 240 309
rect 238 308 239 309
rect 237 308 238 309
rect 236 308 237 309
rect 235 308 236 309
rect 234 308 235 309
rect 233 308 234 309
rect 232 308 233 309
rect 231 308 232 309
rect 230 308 231 309
rect 229 308 230 309
rect 228 308 229 309
rect 227 308 228 309
rect 226 308 227 309
rect 225 308 226 309
rect 224 308 225 309
rect 223 308 224 309
rect 222 308 223 309
rect 221 308 222 309
rect 220 308 221 309
rect 219 308 220 309
rect 218 308 219 309
rect 217 308 218 309
rect 216 308 217 309
rect 215 308 216 309
rect 214 308 215 309
rect 213 308 214 309
rect 212 308 213 309
rect 211 308 212 309
rect 210 308 211 309
rect 209 308 210 309
rect 208 308 209 309
rect 207 308 208 309
rect 206 308 207 309
rect 205 308 206 309
rect 204 308 205 309
rect 203 308 204 309
rect 202 308 203 309
rect 126 308 127 309
rect 125 308 126 309
rect 124 308 125 309
rect 123 308 124 309
rect 122 308 123 309
rect 121 308 122 309
rect 120 308 121 309
rect 119 308 120 309
rect 118 308 119 309
rect 117 308 118 309
rect 116 308 117 309
rect 115 308 116 309
rect 114 308 115 309
rect 113 308 114 309
rect 112 308 113 309
rect 111 308 112 309
rect 110 308 111 309
rect 109 308 110 309
rect 108 308 109 309
rect 107 308 108 309
rect 106 308 107 309
rect 105 308 106 309
rect 104 308 105 309
rect 103 308 104 309
rect 102 308 103 309
rect 101 308 102 309
rect 100 308 101 309
rect 99 308 100 309
rect 98 308 99 309
rect 97 308 98 309
rect 96 308 97 309
rect 95 308 96 309
rect 94 308 95 309
rect 93 308 94 309
rect 92 308 93 309
rect 91 308 92 309
rect 90 308 91 309
rect 89 308 90 309
rect 88 308 89 309
rect 72 308 73 309
rect 71 308 72 309
rect 70 308 71 309
rect 69 308 70 309
rect 68 308 69 309
rect 67 308 68 309
rect 66 308 67 309
rect 65 308 66 309
rect 64 308 65 309
rect 63 308 64 309
rect 62 308 63 309
rect 61 308 62 309
rect 60 308 61 309
rect 59 308 60 309
rect 58 308 59 309
rect 57 308 58 309
rect 56 308 57 309
rect 55 308 56 309
rect 54 308 55 309
rect 53 308 54 309
rect 52 308 53 309
rect 51 308 52 309
rect 50 308 51 309
rect 49 308 50 309
rect 48 308 49 309
rect 47 308 48 309
rect 46 308 47 309
rect 45 308 46 309
rect 44 308 45 309
rect 43 308 44 309
rect 32 308 33 309
rect 31 308 32 309
rect 30 308 31 309
rect 29 308 30 309
rect 28 308 29 309
rect 27 308 28 309
rect 26 308 27 309
rect 25 308 26 309
rect 24 308 25 309
rect 23 308 24 309
rect 22 308 23 309
rect 21 308 22 309
rect 20 308 21 309
rect 19 308 20 309
rect 18 308 19 309
rect 17 308 18 309
rect 16 308 17 309
rect 15 308 16 309
rect 14 308 15 309
rect 13 308 14 309
rect 12 308 13 309
rect 11 308 12 309
rect 10 308 11 309
rect 9 308 10 309
rect 439 309 440 310
rect 438 309 439 310
rect 437 309 438 310
rect 436 309 437 310
rect 435 309 436 310
rect 434 309 435 310
rect 433 309 434 310
rect 432 309 433 310
rect 431 309 432 310
rect 430 309 431 310
rect 429 309 430 310
rect 428 309 429 310
rect 427 309 428 310
rect 426 309 427 310
rect 425 309 426 310
rect 424 309 425 310
rect 423 309 424 310
rect 422 309 423 310
rect 421 309 422 310
rect 420 309 421 310
rect 419 309 420 310
rect 418 309 419 310
rect 417 309 418 310
rect 416 309 417 310
rect 415 309 416 310
rect 414 309 415 310
rect 413 309 414 310
rect 412 309 413 310
rect 411 309 412 310
rect 410 309 411 310
rect 409 309 410 310
rect 408 309 409 310
rect 407 309 408 310
rect 406 309 407 310
rect 405 309 406 310
rect 404 309 405 310
rect 403 309 404 310
rect 402 309 403 310
rect 401 309 402 310
rect 400 309 401 310
rect 399 309 400 310
rect 398 309 399 310
rect 397 309 398 310
rect 396 309 397 310
rect 395 309 396 310
rect 256 309 257 310
rect 255 309 256 310
rect 254 309 255 310
rect 253 309 254 310
rect 252 309 253 310
rect 251 309 252 310
rect 250 309 251 310
rect 249 309 250 310
rect 248 309 249 310
rect 247 309 248 310
rect 246 309 247 310
rect 245 309 246 310
rect 244 309 245 310
rect 243 309 244 310
rect 242 309 243 310
rect 241 309 242 310
rect 240 309 241 310
rect 239 309 240 310
rect 238 309 239 310
rect 237 309 238 310
rect 236 309 237 310
rect 235 309 236 310
rect 234 309 235 310
rect 233 309 234 310
rect 232 309 233 310
rect 231 309 232 310
rect 230 309 231 310
rect 229 309 230 310
rect 228 309 229 310
rect 227 309 228 310
rect 226 309 227 310
rect 225 309 226 310
rect 224 309 225 310
rect 223 309 224 310
rect 222 309 223 310
rect 221 309 222 310
rect 220 309 221 310
rect 219 309 220 310
rect 218 309 219 310
rect 217 309 218 310
rect 216 309 217 310
rect 215 309 216 310
rect 214 309 215 310
rect 213 309 214 310
rect 212 309 213 310
rect 211 309 212 310
rect 210 309 211 310
rect 209 309 210 310
rect 208 309 209 310
rect 207 309 208 310
rect 206 309 207 310
rect 205 309 206 310
rect 204 309 205 310
rect 203 309 204 310
rect 202 309 203 310
rect 201 309 202 310
rect 127 309 128 310
rect 126 309 127 310
rect 125 309 126 310
rect 124 309 125 310
rect 123 309 124 310
rect 122 309 123 310
rect 121 309 122 310
rect 120 309 121 310
rect 119 309 120 310
rect 118 309 119 310
rect 117 309 118 310
rect 116 309 117 310
rect 115 309 116 310
rect 114 309 115 310
rect 113 309 114 310
rect 112 309 113 310
rect 111 309 112 310
rect 110 309 111 310
rect 109 309 110 310
rect 108 309 109 310
rect 107 309 108 310
rect 106 309 107 310
rect 105 309 106 310
rect 104 309 105 310
rect 103 309 104 310
rect 102 309 103 310
rect 101 309 102 310
rect 100 309 101 310
rect 99 309 100 310
rect 98 309 99 310
rect 97 309 98 310
rect 96 309 97 310
rect 95 309 96 310
rect 94 309 95 310
rect 93 309 94 310
rect 92 309 93 310
rect 91 309 92 310
rect 90 309 91 310
rect 89 309 90 310
rect 72 309 73 310
rect 71 309 72 310
rect 70 309 71 310
rect 69 309 70 310
rect 68 309 69 310
rect 67 309 68 310
rect 66 309 67 310
rect 65 309 66 310
rect 64 309 65 310
rect 63 309 64 310
rect 62 309 63 310
rect 61 309 62 310
rect 60 309 61 310
rect 59 309 60 310
rect 58 309 59 310
rect 57 309 58 310
rect 56 309 57 310
rect 55 309 56 310
rect 54 309 55 310
rect 53 309 54 310
rect 52 309 53 310
rect 51 309 52 310
rect 50 309 51 310
rect 49 309 50 310
rect 48 309 49 310
rect 47 309 48 310
rect 46 309 47 310
rect 45 309 46 310
rect 44 309 45 310
rect 43 309 44 310
rect 32 309 33 310
rect 31 309 32 310
rect 30 309 31 310
rect 29 309 30 310
rect 28 309 29 310
rect 27 309 28 310
rect 26 309 27 310
rect 25 309 26 310
rect 24 309 25 310
rect 23 309 24 310
rect 22 309 23 310
rect 21 309 22 310
rect 20 309 21 310
rect 19 309 20 310
rect 18 309 19 310
rect 17 309 18 310
rect 16 309 17 310
rect 15 309 16 310
rect 14 309 15 310
rect 13 309 14 310
rect 12 309 13 310
rect 11 309 12 310
rect 10 309 11 310
rect 439 310 440 311
rect 438 310 439 311
rect 437 310 438 311
rect 436 310 437 311
rect 435 310 436 311
rect 434 310 435 311
rect 433 310 434 311
rect 432 310 433 311
rect 431 310 432 311
rect 430 310 431 311
rect 429 310 430 311
rect 428 310 429 311
rect 427 310 428 311
rect 426 310 427 311
rect 425 310 426 311
rect 424 310 425 311
rect 423 310 424 311
rect 422 310 423 311
rect 421 310 422 311
rect 420 310 421 311
rect 419 310 420 311
rect 418 310 419 311
rect 417 310 418 311
rect 416 310 417 311
rect 415 310 416 311
rect 414 310 415 311
rect 413 310 414 311
rect 412 310 413 311
rect 411 310 412 311
rect 410 310 411 311
rect 409 310 410 311
rect 408 310 409 311
rect 407 310 408 311
rect 406 310 407 311
rect 405 310 406 311
rect 404 310 405 311
rect 403 310 404 311
rect 402 310 403 311
rect 401 310 402 311
rect 400 310 401 311
rect 399 310 400 311
rect 398 310 399 311
rect 397 310 398 311
rect 396 310 397 311
rect 395 310 396 311
rect 254 310 255 311
rect 253 310 254 311
rect 252 310 253 311
rect 251 310 252 311
rect 250 310 251 311
rect 249 310 250 311
rect 248 310 249 311
rect 247 310 248 311
rect 246 310 247 311
rect 245 310 246 311
rect 244 310 245 311
rect 243 310 244 311
rect 242 310 243 311
rect 241 310 242 311
rect 240 310 241 311
rect 239 310 240 311
rect 238 310 239 311
rect 237 310 238 311
rect 236 310 237 311
rect 235 310 236 311
rect 234 310 235 311
rect 233 310 234 311
rect 232 310 233 311
rect 231 310 232 311
rect 230 310 231 311
rect 229 310 230 311
rect 228 310 229 311
rect 227 310 228 311
rect 226 310 227 311
rect 225 310 226 311
rect 224 310 225 311
rect 223 310 224 311
rect 222 310 223 311
rect 221 310 222 311
rect 220 310 221 311
rect 219 310 220 311
rect 218 310 219 311
rect 217 310 218 311
rect 216 310 217 311
rect 215 310 216 311
rect 214 310 215 311
rect 213 310 214 311
rect 212 310 213 311
rect 211 310 212 311
rect 210 310 211 311
rect 209 310 210 311
rect 208 310 209 311
rect 207 310 208 311
rect 206 310 207 311
rect 205 310 206 311
rect 204 310 205 311
rect 203 310 204 311
rect 202 310 203 311
rect 201 310 202 311
rect 200 310 201 311
rect 128 310 129 311
rect 127 310 128 311
rect 126 310 127 311
rect 125 310 126 311
rect 124 310 125 311
rect 123 310 124 311
rect 122 310 123 311
rect 121 310 122 311
rect 120 310 121 311
rect 119 310 120 311
rect 118 310 119 311
rect 117 310 118 311
rect 116 310 117 311
rect 115 310 116 311
rect 114 310 115 311
rect 113 310 114 311
rect 112 310 113 311
rect 111 310 112 311
rect 110 310 111 311
rect 109 310 110 311
rect 108 310 109 311
rect 107 310 108 311
rect 106 310 107 311
rect 105 310 106 311
rect 104 310 105 311
rect 103 310 104 311
rect 102 310 103 311
rect 101 310 102 311
rect 100 310 101 311
rect 99 310 100 311
rect 98 310 99 311
rect 97 310 98 311
rect 96 310 97 311
rect 95 310 96 311
rect 94 310 95 311
rect 93 310 94 311
rect 92 310 93 311
rect 91 310 92 311
rect 90 310 91 311
rect 89 310 90 311
rect 72 310 73 311
rect 71 310 72 311
rect 70 310 71 311
rect 69 310 70 311
rect 68 310 69 311
rect 67 310 68 311
rect 66 310 67 311
rect 65 310 66 311
rect 64 310 65 311
rect 63 310 64 311
rect 62 310 63 311
rect 61 310 62 311
rect 60 310 61 311
rect 59 310 60 311
rect 58 310 59 311
rect 57 310 58 311
rect 56 310 57 311
rect 55 310 56 311
rect 54 310 55 311
rect 53 310 54 311
rect 52 310 53 311
rect 51 310 52 311
rect 50 310 51 311
rect 49 310 50 311
rect 48 310 49 311
rect 47 310 48 311
rect 46 310 47 311
rect 45 310 46 311
rect 44 310 45 311
rect 32 310 33 311
rect 31 310 32 311
rect 30 310 31 311
rect 29 310 30 311
rect 28 310 29 311
rect 27 310 28 311
rect 26 310 27 311
rect 25 310 26 311
rect 24 310 25 311
rect 23 310 24 311
rect 22 310 23 311
rect 21 310 22 311
rect 20 310 21 311
rect 19 310 20 311
rect 18 310 19 311
rect 17 310 18 311
rect 16 310 17 311
rect 15 310 16 311
rect 14 310 15 311
rect 13 310 14 311
rect 12 310 13 311
rect 11 310 12 311
rect 10 310 11 311
rect 439 311 440 312
rect 438 311 439 312
rect 437 311 438 312
rect 436 311 437 312
rect 435 311 436 312
rect 434 311 435 312
rect 433 311 434 312
rect 432 311 433 312
rect 431 311 432 312
rect 430 311 431 312
rect 429 311 430 312
rect 428 311 429 312
rect 427 311 428 312
rect 426 311 427 312
rect 425 311 426 312
rect 424 311 425 312
rect 423 311 424 312
rect 422 311 423 312
rect 421 311 422 312
rect 420 311 421 312
rect 419 311 420 312
rect 418 311 419 312
rect 417 311 418 312
rect 416 311 417 312
rect 415 311 416 312
rect 414 311 415 312
rect 413 311 414 312
rect 412 311 413 312
rect 411 311 412 312
rect 410 311 411 312
rect 409 311 410 312
rect 408 311 409 312
rect 407 311 408 312
rect 406 311 407 312
rect 405 311 406 312
rect 404 311 405 312
rect 403 311 404 312
rect 402 311 403 312
rect 401 311 402 312
rect 400 311 401 312
rect 399 311 400 312
rect 398 311 399 312
rect 397 311 398 312
rect 396 311 397 312
rect 395 311 396 312
rect 253 311 254 312
rect 252 311 253 312
rect 251 311 252 312
rect 250 311 251 312
rect 249 311 250 312
rect 248 311 249 312
rect 247 311 248 312
rect 246 311 247 312
rect 245 311 246 312
rect 244 311 245 312
rect 243 311 244 312
rect 242 311 243 312
rect 241 311 242 312
rect 240 311 241 312
rect 239 311 240 312
rect 238 311 239 312
rect 237 311 238 312
rect 236 311 237 312
rect 235 311 236 312
rect 234 311 235 312
rect 233 311 234 312
rect 232 311 233 312
rect 231 311 232 312
rect 230 311 231 312
rect 229 311 230 312
rect 228 311 229 312
rect 227 311 228 312
rect 226 311 227 312
rect 225 311 226 312
rect 224 311 225 312
rect 223 311 224 312
rect 222 311 223 312
rect 221 311 222 312
rect 220 311 221 312
rect 219 311 220 312
rect 218 311 219 312
rect 217 311 218 312
rect 216 311 217 312
rect 215 311 216 312
rect 214 311 215 312
rect 213 311 214 312
rect 212 311 213 312
rect 211 311 212 312
rect 210 311 211 312
rect 209 311 210 312
rect 208 311 209 312
rect 207 311 208 312
rect 206 311 207 312
rect 205 311 206 312
rect 204 311 205 312
rect 203 311 204 312
rect 202 311 203 312
rect 201 311 202 312
rect 200 311 201 312
rect 199 311 200 312
rect 129 311 130 312
rect 128 311 129 312
rect 127 311 128 312
rect 126 311 127 312
rect 125 311 126 312
rect 124 311 125 312
rect 123 311 124 312
rect 122 311 123 312
rect 121 311 122 312
rect 120 311 121 312
rect 119 311 120 312
rect 118 311 119 312
rect 117 311 118 312
rect 116 311 117 312
rect 115 311 116 312
rect 114 311 115 312
rect 113 311 114 312
rect 112 311 113 312
rect 111 311 112 312
rect 110 311 111 312
rect 109 311 110 312
rect 108 311 109 312
rect 107 311 108 312
rect 106 311 107 312
rect 105 311 106 312
rect 104 311 105 312
rect 103 311 104 312
rect 102 311 103 312
rect 101 311 102 312
rect 100 311 101 312
rect 99 311 100 312
rect 98 311 99 312
rect 97 311 98 312
rect 96 311 97 312
rect 95 311 96 312
rect 94 311 95 312
rect 93 311 94 312
rect 92 311 93 312
rect 91 311 92 312
rect 90 311 91 312
rect 73 311 74 312
rect 72 311 73 312
rect 71 311 72 312
rect 70 311 71 312
rect 69 311 70 312
rect 68 311 69 312
rect 67 311 68 312
rect 66 311 67 312
rect 65 311 66 312
rect 64 311 65 312
rect 63 311 64 312
rect 62 311 63 312
rect 61 311 62 312
rect 60 311 61 312
rect 59 311 60 312
rect 58 311 59 312
rect 57 311 58 312
rect 56 311 57 312
rect 55 311 56 312
rect 54 311 55 312
rect 53 311 54 312
rect 52 311 53 312
rect 51 311 52 312
rect 50 311 51 312
rect 49 311 50 312
rect 48 311 49 312
rect 47 311 48 312
rect 46 311 47 312
rect 45 311 46 312
rect 44 311 45 312
rect 33 311 34 312
rect 32 311 33 312
rect 31 311 32 312
rect 30 311 31 312
rect 29 311 30 312
rect 28 311 29 312
rect 27 311 28 312
rect 26 311 27 312
rect 25 311 26 312
rect 24 311 25 312
rect 23 311 24 312
rect 22 311 23 312
rect 21 311 22 312
rect 20 311 21 312
rect 19 311 20 312
rect 18 311 19 312
rect 17 311 18 312
rect 16 311 17 312
rect 15 311 16 312
rect 14 311 15 312
rect 13 311 14 312
rect 12 311 13 312
rect 11 311 12 312
rect 460 312 461 313
rect 439 312 440 313
rect 438 312 439 313
rect 437 312 438 313
rect 436 312 437 313
rect 435 312 436 313
rect 434 312 435 313
rect 433 312 434 313
rect 432 312 433 313
rect 431 312 432 313
rect 430 312 431 313
rect 429 312 430 313
rect 428 312 429 313
rect 427 312 428 313
rect 426 312 427 313
rect 425 312 426 313
rect 424 312 425 313
rect 423 312 424 313
rect 422 312 423 313
rect 421 312 422 313
rect 420 312 421 313
rect 419 312 420 313
rect 418 312 419 313
rect 417 312 418 313
rect 416 312 417 313
rect 415 312 416 313
rect 414 312 415 313
rect 413 312 414 313
rect 412 312 413 313
rect 411 312 412 313
rect 410 312 411 313
rect 409 312 410 313
rect 408 312 409 313
rect 407 312 408 313
rect 406 312 407 313
rect 405 312 406 313
rect 404 312 405 313
rect 403 312 404 313
rect 402 312 403 313
rect 401 312 402 313
rect 400 312 401 313
rect 399 312 400 313
rect 398 312 399 313
rect 397 312 398 313
rect 396 312 397 313
rect 395 312 396 313
rect 251 312 252 313
rect 250 312 251 313
rect 249 312 250 313
rect 248 312 249 313
rect 247 312 248 313
rect 246 312 247 313
rect 245 312 246 313
rect 244 312 245 313
rect 243 312 244 313
rect 242 312 243 313
rect 241 312 242 313
rect 240 312 241 313
rect 239 312 240 313
rect 238 312 239 313
rect 237 312 238 313
rect 236 312 237 313
rect 235 312 236 313
rect 234 312 235 313
rect 233 312 234 313
rect 232 312 233 313
rect 231 312 232 313
rect 230 312 231 313
rect 229 312 230 313
rect 228 312 229 313
rect 227 312 228 313
rect 226 312 227 313
rect 225 312 226 313
rect 224 312 225 313
rect 223 312 224 313
rect 222 312 223 313
rect 221 312 222 313
rect 220 312 221 313
rect 219 312 220 313
rect 218 312 219 313
rect 217 312 218 313
rect 216 312 217 313
rect 215 312 216 313
rect 214 312 215 313
rect 213 312 214 313
rect 212 312 213 313
rect 211 312 212 313
rect 210 312 211 313
rect 209 312 210 313
rect 208 312 209 313
rect 207 312 208 313
rect 206 312 207 313
rect 205 312 206 313
rect 204 312 205 313
rect 203 312 204 313
rect 202 312 203 313
rect 201 312 202 313
rect 200 312 201 313
rect 199 312 200 313
rect 198 312 199 313
rect 130 312 131 313
rect 129 312 130 313
rect 128 312 129 313
rect 127 312 128 313
rect 126 312 127 313
rect 125 312 126 313
rect 124 312 125 313
rect 123 312 124 313
rect 122 312 123 313
rect 121 312 122 313
rect 120 312 121 313
rect 119 312 120 313
rect 118 312 119 313
rect 117 312 118 313
rect 116 312 117 313
rect 115 312 116 313
rect 114 312 115 313
rect 113 312 114 313
rect 112 312 113 313
rect 111 312 112 313
rect 110 312 111 313
rect 109 312 110 313
rect 108 312 109 313
rect 107 312 108 313
rect 106 312 107 313
rect 105 312 106 313
rect 104 312 105 313
rect 103 312 104 313
rect 102 312 103 313
rect 101 312 102 313
rect 100 312 101 313
rect 99 312 100 313
rect 98 312 99 313
rect 97 312 98 313
rect 96 312 97 313
rect 95 312 96 313
rect 94 312 95 313
rect 93 312 94 313
rect 92 312 93 313
rect 91 312 92 313
rect 73 312 74 313
rect 72 312 73 313
rect 71 312 72 313
rect 70 312 71 313
rect 69 312 70 313
rect 68 312 69 313
rect 67 312 68 313
rect 66 312 67 313
rect 65 312 66 313
rect 64 312 65 313
rect 63 312 64 313
rect 62 312 63 313
rect 61 312 62 313
rect 60 312 61 313
rect 59 312 60 313
rect 58 312 59 313
rect 57 312 58 313
rect 56 312 57 313
rect 55 312 56 313
rect 54 312 55 313
rect 53 312 54 313
rect 52 312 53 313
rect 51 312 52 313
rect 50 312 51 313
rect 49 312 50 313
rect 48 312 49 313
rect 47 312 48 313
rect 46 312 47 313
rect 45 312 46 313
rect 44 312 45 313
rect 33 312 34 313
rect 32 312 33 313
rect 31 312 32 313
rect 30 312 31 313
rect 29 312 30 313
rect 28 312 29 313
rect 27 312 28 313
rect 26 312 27 313
rect 25 312 26 313
rect 24 312 25 313
rect 23 312 24 313
rect 22 312 23 313
rect 21 312 22 313
rect 20 312 21 313
rect 19 312 20 313
rect 18 312 19 313
rect 17 312 18 313
rect 16 312 17 313
rect 15 312 16 313
rect 14 312 15 313
rect 13 312 14 313
rect 12 312 13 313
rect 460 313 461 314
rect 439 313 440 314
rect 438 313 439 314
rect 437 313 438 314
rect 436 313 437 314
rect 435 313 436 314
rect 434 313 435 314
rect 433 313 434 314
rect 432 313 433 314
rect 431 313 432 314
rect 430 313 431 314
rect 429 313 430 314
rect 428 313 429 314
rect 427 313 428 314
rect 426 313 427 314
rect 425 313 426 314
rect 424 313 425 314
rect 423 313 424 314
rect 422 313 423 314
rect 421 313 422 314
rect 420 313 421 314
rect 419 313 420 314
rect 418 313 419 314
rect 417 313 418 314
rect 416 313 417 314
rect 415 313 416 314
rect 414 313 415 314
rect 413 313 414 314
rect 412 313 413 314
rect 411 313 412 314
rect 410 313 411 314
rect 409 313 410 314
rect 408 313 409 314
rect 407 313 408 314
rect 406 313 407 314
rect 405 313 406 314
rect 404 313 405 314
rect 403 313 404 314
rect 402 313 403 314
rect 401 313 402 314
rect 400 313 401 314
rect 399 313 400 314
rect 398 313 399 314
rect 397 313 398 314
rect 396 313 397 314
rect 395 313 396 314
rect 249 313 250 314
rect 248 313 249 314
rect 247 313 248 314
rect 246 313 247 314
rect 245 313 246 314
rect 244 313 245 314
rect 243 313 244 314
rect 242 313 243 314
rect 241 313 242 314
rect 240 313 241 314
rect 239 313 240 314
rect 238 313 239 314
rect 237 313 238 314
rect 236 313 237 314
rect 235 313 236 314
rect 234 313 235 314
rect 233 313 234 314
rect 232 313 233 314
rect 231 313 232 314
rect 230 313 231 314
rect 229 313 230 314
rect 228 313 229 314
rect 227 313 228 314
rect 226 313 227 314
rect 225 313 226 314
rect 224 313 225 314
rect 223 313 224 314
rect 222 313 223 314
rect 221 313 222 314
rect 220 313 221 314
rect 219 313 220 314
rect 218 313 219 314
rect 217 313 218 314
rect 216 313 217 314
rect 215 313 216 314
rect 214 313 215 314
rect 213 313 214 314
rect 212 313 213 314
rect 211 313 212 314
rect 210 313 211 314
rect 209 313 210 314
rect 208 313 209 314
rect 207 313 208 314
rect 206 313 207 314
rect 205 313 206 314
rect 204 313 205 314
rect 203 313 204 314
rect 202 313 203 314
rect 201 313 202 314
rect 200 313 201 314
rect 199 313 200 314
rect 198 313 199 314
rect 197 313 198 314
rect 131 313 132 314
rect 130 313 131 314
rect 129 313 130 314
rect 128 313 129 314
rect 127 313 128 314
rect 126 313 127 314
rect 125 313 126 314
rect 124 313 125 314
rect 123 313 124 314
rect 122 313 123 314
rect 121 313 122 314
rect 120 313 121 314
rect 119 313 120 314
rect 118 313 119 314
rect 117 313 118 314
rect 116 313 117 314
rect 115 313 116 314
rect 114 313 115 314
rect 113 313 114 314
rect 112 313 113 314
rect 111 313 112 314
rect 110 313 111 314
rect 109 313 110 314
rect 108 313 109 314
rect 107 313 108 314
rect 106 313 107 314
rect 105 313 106 314
rect 104 313 105 314
rect 103 313 104 314
rect 102 313 103 314
rect 101 313 102 314
rect 100 313 101 314
rect 99 313 100 314
rect 98 313 99 314
rect 97 313 98 314
rect 96 313 97 314
rect 95 313 96 314
rect 94 313 95 314
rect 93 313 94 314
rect 92 313 93 314
rect 91 313 92 314
rect 74 313 75 314
rect 73 313 74 314
rect 72 313 73 314
rect 71 313 72 314
rect 70 313 71 314
rect 69 313 70 314
rect 68 313 69 314
rect 67 313 68 314
rect 66 313 67 314
rect 65 313 66 314
rect 64 313 65 314
rect 63 313 64 314
rect 62 313 63 314
rect 61 313 62 314
rect 60 313 61 314
rect 59 313 60 314
rect 58 313 59 314
rect 57 313 58 314
rect 56 313 57 314
rect 55 313 56 314
rect 54 313 55 314
rect 53 313 54 314
rect 52 313 53 314
rect 51 313 52 314
rect 50 313 51 314
rect 49 313 50 314
rect 48 313 49 314
rect 47 313 48 314
rect 46 313 47 314
rect 45 313 46 314
rect 33 313 34 314
rect 32 313 33 314
rect 31 313 32 314
rect 30 313 31 314
rect 29 313 30 314
rect 28 313 29 314
rect 27 313 28 314
rect 26 313 27 314
rect 25 313 26 314
rect 24 313 25 314
rect 23 313 24 314
rect 22 313 23 314
rect 21 313 22 314
rect 20 313 21 314
rect 19 313 20 314
rect 18 313 19 314
rect 17 313 18 314
rect 16 313 17 314
rect 15 313 16 314
rect 14 313 15 314
rect 13 313 14 314
rect 12 313 13 314
rect 461 314 462 315
rect 460 314 461 315
rect 439 314 440 315
rect 438 314 439 315
rect 437 314 438 315
rect 436 314 437 315
rect 435 314 436 315
rect 434 314 435 315
rect 433 314 434 315
rect 432 314 433 315
rect 431 314 432 315
rect 430 314 431 315
rect 429 314 430 315
rect 428 314 429 315
rect 427 314 428 315
rect 426 314 427 315
rect 425 314 426 315
rect 424 314 425 315
rect 423 314 424 315
rect 422 314 423 315
rect 421 314 422 315
rect 420 314 421 315
rect 419 314 420 315
rect 418 314 419 315
rect 417 314 418 315
rect 416 314 417 315
rect 415 314 416 315
rect 414 314 415 315
rect 413 314 414 315
rect 412 314 413 315
rect 411 314 412 315
rect 410 314 411 315
rect 409 314 410 315
rect 408 314 409 315
rect 407 314 408 315
rect 406 314 407 315
rect 405 314 406 315
rect 404 314 405 315
rect 403 314 404 315
rect 402 314 403 315
rect 401 314 402 315
rect 400 314 401 315
rect 399 314 400 315
rect 398 314 399 315
rect 397 314 398 315
rect 396 314 397 315
rect 395 314 396 315
rect 247 314 248 315
rect 246 314 247 315
rect 245 314 246 315
rect 244 314 245 315
rect 243 314 244 315
rect 242 314 243 315
rect 241 314 242 315
rect 240 314 241 315
rect 239 314 240 315
rect 238 314 239 315
rect 237 314 238 315
rect 236 314 237 315
rect 235 314 236 315
rect 234 314 235 315
rect 233 314 234 315
rect 232 314 233 315
rect 231 314 232 315
rect 230 314 231 315
rect 229 314 230 315
rect 228 314 229 315
rect 227 314 228 315
rect 226 314 227 315
rect 225 314 226 315
rect 224 314 225 315
rect 223 314 224 315
rect 222 314 223 315
rect 221 314 222 315
rect 220 314 221 315
rect 219 314 220 315
rect 218 314 219 315
rect 217 314 218 315
rect 216 314 217 315
rect 215 314 216 315
rect 214 314 215 315
rect 213 314 214 315
rect 212 314 213 315
rect 211 314 212 315
rect 210 314 211 315
rect 209 314 210 315
rect 208 314 209 315
rect 207 314 208 315
rect 206 314 207 315
rect 205 314 206 315
rect 204 314 205 315
rect 203 314 204 315
rect 202 314 203 315
rect 201 314 202 315
rect 200 314 201 315
rect 199 314 200 315
rect 198 314 199 315
rect 197 314 198 315
rect 196 314 197 315
rect 132 314 133 315
rect 131 314 132 315
rect 130 314 131 315
rect 129 314 130 315
rect 128 314 129 315
rect 127 314 128 315
rect 126 314 127 315
rect 125 314 126 315
rect 124 314 125 315
rect 123 314 124 315
rect 122 314 123 315
rect 121 314 122 315
rect 120 314 121 315
rect 119 314 120 315
rect 118 314 119 315
rect 117 314 118 315
rect 116 314 117 315
rect 115 314 116 315
rect 114 314 115 315
rect 113 314 114 315
rect 112 314 113 315
rect 111 314 112 315
rect 110 314 111 315
rect 109 314 110 315
rect 108 314 109 315
rect 107 314 108 315
rect 106 314 107 315
rect 105 314 106 315
rect 104 314 105 315
rect 103 314 104 315
rect 102 314 103 315
rect 101 314 102 315
rect 100 314 101 315
rect 99 314 100 315
rect 98 314 99 315
rect 97 314 98 315
rect 96 314 97 315
rect 95 314 96 315
rect 94 314 95 315
rect 93 314 94 315
rect 92 314 93 315
rect 74 314 75 315
rect 73 314 74 315
rect 72 314 73 315
rect 71 314 72 315
rect 70 314 71 315
rect 69 314 70 315
rect 68 314 69 315
rect 67 314 68 315
rect 66 314 67 315
rect 65 314 66 315
rect 64 314 65 315
rect 63 314 64 315
rect 62 314 63 315
rect 61 314 62 315
rect 60 314 61 315
rect 59 314 60 315
rect 58 314 59 315
rect 57 314 58 315
rect 56 314 57 315
rect 55 314 56 315
rect 54 314 55 315
rect 53 314 54 315
rect 52 314 53 315
rect 51 314 52 315
rect 50 314 51 315
rect 49 314 50 315
rect 48 314 49 315
rect 47 314 48 315
rect 46 314 47 315
rect 45 314 46 315
rect 33 314 34 315
rect 32 314 33 315
rect 31 314 32 315
rect 30 314 31 315
rect 29 314 30 315
rect 28 314 29 315
rect 27 314 28 315
rect 26 314 27 315
rect 25 314 26 315
rect 24 314 25 315
rect 23 314 24 315
rect 22 314 23 315
rect 21 314 22 315
rect 20 314 21 315
rect 19 314 20 315
rect 18 314 19 315
rect 17 314 18 315
rect 16 314 17 315
rect 15 314 16 315
rect 14 314 15 315
rect 13 314 14 315
rect 463 315 464 316
rect 462 315 463 316
rect 461 315 462 316
rect 460 315 461 316
rect 439 315 440 316
rect 438 315 439 316
rect 437 315 438 316
rect 436 315 437 316
rect 435 315 436 316
rect 434 315 435 316
rect 433 315 434 316
rect 432 315 433 316
rect 431 315 432 316
rect 430 315 431 316
rect 429 315 430 316
rect 428 315 429 316
rect 427 315 428 316
rect 426 315 427 316
rect 425 315 426 316
rect 424 315 425 316
rect 423 315 424 316
rect 422 315 423 316
rect 421 315 422 316
rect 420 315 421 316
rect 419 315 420 316
rect 418 315 419 316
rect 417 315 418 316
rect 416 315 417 316
rect 415 315 416 316
rect 414 315 415 316
rect 413 315 414 316
rect 412 315 413 316
rect 411 315 412 316
rect 410 315 411 316
rect 409 315 410 316
rect 408 315 409 316
rect 407 315 408 316
rect 406 315 407 316
rect 405 315 406 316
rect 404 315 405 316
rect 403 315 404 316
rect 402 315 403 316
rect 401 315 402 316
rect 400 315 401 316
rect 399 315 400 316
rect 398 315 399 316
rect 397 315 398 316
rect 396 315 397 316
rect 395 315 396 316
rect 245 315 246 316
rect 244 315 245 316
rect 243 315 244 316
rect 242 315 243 316
rect 241 315 242 316
rect 240 315 241 316
rect 239 315 240 316
rect 238 315 239 316
rect 237 315 238 316
rect 236 315 237 316
rect 235 315 236 316
rect 234 315 235 316
rect 233 315 234 316
rect 232 315 233 316
rect 231 315 232 316
rect 230 315 231 316
rect 229 315 230 316
rect 228 315 229 316
rect 227 315 228 316
rect 226 315 227 316
rect 225 315 226 316
rect 224 315 225 316
rect 223 315 224 316
rect 222 315 223 316
rect 221 315 222 316
rect 220 315 221 316
rect 219 315 220 316
rect 218 315 219 316
rect 217 315 218 316
rect 216 315 217 316
rect 215 315 216 316
rect 214 315 215 316
rect 213 315 214 316
rect 212 315 213 316
rect 211 315 212 316
rect 210 315 211 316
rect 209 315 210 316
rect 208 315 209 316
rect 207 315 208 316
rect 206 315 207 316
rect 205 315 206 316
rect 204 315 205 316
rect 203 315 204 316
rect 202 315 203 316
rect 201 315 202 316
rect 200 315 201 316
rect 199 315 200 316
rect 198 315 199 316
rect 197 315 198 316
rect 196 315 197 316
rect 195 315 196 316
rect 133 315 134 316
rect 132 315 133 316
rect 131 315 132 316
rect 130 315 131 316
rect 129 315 130 316
rect 128 315 129 316
rect 127 315 128 316
rect 126 315 127 316
rect 125 315 126 316
rect 124 315 125 316
rect 123 315 124 316
rect 122 315 123 316
rect 121 315 122 316
rect 120 315 121 316
rect 119 315 120 316
rect 118 315 119 316
rect 117 315 118 316
rect 116 315 117 316
rect 115 315 116 316
rect 114 315 115 316
rect 113 315 114 316
rect 112 315 113 316
rect 111 315 112 316
rect 110 315 111 316
rect 109 315 110 316
rect 108 315 109 316
rect 107 315 108 316
rect 106 315 107 316
rect 105 315 106 316
rect 104 315 105 316
rect 103 315 104 316
rect 102 315 103 316
rect 101 315 102 316
rect 100 315 101 316
rect 99 315 100 316
rect 98 315 99 316
rect 97 315 98 316
rect 96 315 97 316
rect 95 315 96 316
rect 94 315 95 316
rect 93 315 94 316
rect 92 315 93 316
rect 75 315 76 316
rect 74 315 75 316
rect 73 315 74 316
rect 72 315 73 316
rect 71 315 72 316
rect 70 315 71 316
rect 69 315 70 316
rect 68 315 69 316
rect 67 315 68 316
rect 66 315 67 316
rect 65 315 66 316
rect 64 315 65 316
rect 63 315 64 316
rect 62 315 63 316
rect 61 315 62 316
rect 60 315 61 316
rect 59 315 60 316
rect 58 315 59 316
rect 57 315 58 316
rect 56 315 57 316
rect 55 315 56 316
rect 54 315 55 316
rect 53 315 54 316
rect 52 315 53 316
rect 51 315 52 316
rect 50 315 51 316
rect 49 315 50 316
rect 48 315 49 316
rect 47 315 48 316
rect 46 315 47 316
rect 45 315 46 316
rect 34 315 35 316
rect 33 315 34 316
rect 32 315 33 316
rect 31 315 32 316
rect 30 315 31 316
rect 29 315 30 316
rect 28 315 29 316
rect 27 315 28 316
rect 26 315 27 316
rect 25 315 26 316
rect 24 315 25 316
rect 23 315 24 316
rect 22 315 23 316
rect 21 315 22 316
rect 20 315 21 316
rect 19 315 20 316
rect 18 315 19 316
rect 17 315 18 316
rect 16 315 17 316
rect 15 315 16 316
rect 14 315 15 316
rect 13 315 14 316
rect 465 316 466 317
rect 464 316 465 317
rect 463 316 464 317
rect 462 316 463 317
rect 461 316 462 317
rect 460 316 461 317
rect 439 316 440 317
rect 438 316 439 317
rect 437 316 438 317
rect 436 316 437 317
rect 435 316 436 317
rect 434 316 435 317
rect 433 316 434 317
rect 432 316 433 317
rect 431 316 432 317
rect 430 316 431 317
rect 429 316 430 317
rect 428 316 429 317
rect 427 316 428 317
rect 426 316 427 317
rect 425 316 426 317
rect 424 316 425 317
rect 423 316 424 317
rect 422 316 423 317
rect 421 316 422 317
rect 420 316 421 317
rect 419 316 420 317
rect 418 316 419 317
rect 417 316 418 317
rect 416 316 417 317
rect 415 316 416 317
rect 414 316 415 317
rect 413 316 414 317
rect 412 316 413 317
rect 411 316 412 317
rect 410 316 411 317
rect 409 316 410 317
rect 408 316 409 317
rect 407 316 408 317
rect 406 316 407 317
rect 405 316 406 317
rect 404 316 405 317
rect 403 316 404 317
rect 402 316 403 317
rect 401 316 402 317
rect 400 316 401 317
rect 399 316 400 317
rect 398 316 399 317
rect 397 316 398 317
rect 396 316 397 317
rect 395 316 396 317
rect 242 316 243 317
rect 241 316 242 317
rect 240 316 241 317
rect 239 316 240 317
rect 238 316 239 317
rect 237 316 238 317
rect 236 316 237 317
rect 235 316 236 317
rect 234 316 235 317
rect 233 316 234 317
rect 232 316 233 317
rect 231 316 232 317
rect 230 316 231 317
rect 229 316 230 317
rect 228 316 229 317
rect 227 316 228 317
rect 226 316 227 317
rect 225 316 226 317
rect 224 316 225 317
rect 223 316 224 317
rect 222 316 223 317
rect 221 316 222 317
rect 220 316 221 317
rect 219 316 220 317
rect 218 316 219 317
rect 217 316 218 317
rect 216 316 217 317
rect 215 316 216 317
rect 214 316 215 317
rect 213 316 214 317
rect 212 316 213 317
rect 211 316 212 317
rect 210 316 211 317
rect 209 316 210 317
rect 208 316 209 317
rect 207 316 208 317
rect 206 316 207 317
rect 205 316 206 317
rect 204 316 205 317
rect 203 316 204 317
rect 202 316 203 317
rect 201 316 202 317
rect 200 316 201 317
rect 199 316 200 317
rect 198 316 199 317
rect 197 316 198 317
rect 196 316 197 317
rect 195 316 196 317
rect 194 316 195 317
rect 134 316 135 317
rect 133 316 134 317
rect 132 316 133 317
rect 131 316 132 317
rect 130 316 131 317
rect 129 316 130 317
rect 128 316 129 317
rect 127 316 128 317
rect 126 316 127 317
rect 125 316 126 317
rect 124 316 125 317
rect 123 316 124 317
rect 122 316 123 317
rect 121 316 122 317
rect 120 316 121 317
rect 119 316 120 317
rect 118 316 119 317
rect 117 316 118 317
rect 116 316 117 317
rect 115 316 116 317
rect 114 316 115 317
rect 113 316 114 317
rect 112 316 113 317
rect 111 316 112 317
rect 110 316 111 317
rect 109 316 110 317
rect 108 316 109 317
rect 107 316 108 317
rect 106 316 107 317
rect 105 316 106 317
rect 104 316 105 317
rect 103 316 104 317
rect 102 316 103 317
rect 101 316 102 317
rect 100 316 101 317
rect 99 316 100 317
rect 98 316 99 317
rect 97 316 98 317
rect 96 316 97 317
rect 95 316 96 317
rect 94 316 95 317
rect 93 316 94 317
rect 75 316 76 317
rect 74 316 75 317
rect 73 316 74 317
rect 72 316 73 317
rect 71 316 72 317
rect 70 316 71 317
rect 69 316 70 317
rect 68 316 69 317
rect 67 316 68 317
rect 66 316 67 317
rect 65 316 66 317
rect 64 316 65 317
rect 63 316 64 317
rect 62 316 63 317
rect 61 316 62 317
rect 60 316 61 317
rect 59 316 60 317
rect 58 316 59 317
rect 57 316 58 317
rect 56 316 57 317
rect 55 316 56 317
rect 54 316 55 317
rect 53 316 54 317
rect 52 316 53 317
rect 51 316 52 317
rect 50 316 51 317
rect 49 316 50 317
rect 48 316 49 317
rect 47 316 48 317
rect 46 316 47 317
rect 34 316 35 317
rect 33 316 34 317
rect 32 316 33 317
rect 31 316 32 317
rect 30 316 31 317
rect 29 316 30 317
rect 28 316 29 317
rect 27 316 28 317
rect 26 316 27 317
rect 25 316 26 317
rect 24 316 25 317
rect 23 316 24 317
rect 22 316 23 317
rect 21 316 22 317
rect 20 316 21 317
rect 19 316 20 317
rect 18 316 19 317
rect 17 316 18 317
rect 16 316 17 317
rect 15 316 16 317
rect 14 316 15 317
rect 480 317 481 318
rect 466 317 467 318
rect 465 317 466 318
rect 464 317 465 318
rect 463 317 464 318
rect 462 317 463 318
rect 461 317 462 318
rect 460 317 461 318
rect 439 317 440 318
rect 438 317 439 318
rect 437 317 438 318
rect 436 317 437 318
rect 435 317 436 318
rect 434 317 435 318
rect 433 317 434 318
rect 432 317 433 318
rect 431 317 432 318
rect 430 317 431 318
rect 429 317 430 318
rect 428 317 429 318
rect 427 317 428 318
rect 426 317 427 318
rect 425 317 426 318
rect 424 317 425 318
rect 423 317 424 318
rect 422 317 423 318
rect 421 317 422 318
rect 420 317 421 318
rect 419 317 420 318
rect 418 317 419 318
rect 417 317 418 318
rect 416 317 417 318
rect 415 317 416 318
rect 414 317 415 318
rect 413 317 414 318
rect 412 317 413 318
rect 411 317 412 318
rect 410 317 411 318
rect 409 317 410 318
rect 408 317 409 318
rect 407 317 408 318
rect 406 317 407 318
rect 405 317 406 318
rect 404 317 405 318
rect 403 317 404 318
rect 402 317 403 318
rect 401 317 402 318
rect 400 317 401 318
rect 399 317 400 318
rect 398 317 399 318
rect 397 317 398 318
rect 396 317 397 318
rect 395 317 396 318
rect 240 317 241 318
rect 239 317 240 318
rect 238 317 239 318
rect 237 317 238 318
rect 236 317 237 318
rect 235 317 236 318
rect 234 317 235 318
rect 233 317 234 318
rect 232 317 233 318
rect 231 317 232 318
rect 230 317 231 318
rect 229 317 230 318
rect 228 317 229 318
rect 227 317 228 318
rect 226 317 227 318
rect 225 317 226 318
rect 224 317 225 318
rect 223 317 224 318
rect 222 317 223 318
rect 221 317 222 318
rect 220 317 221 318
rect 219 317 220 318
rect 218 317 219 318
rect 217 317 218 318
rect 216 317 217 318
rect 215 317 216 318
rect 214 317 215 318
rect 213 317 214 318
rect 212 317 213 318
rect 211 317 212 318
rect 210 317 211 318
rect 209 317 210 318
rect 208 317 209 318
rect 207 317 208 318
rect 206 317 207 318
rect 205 317 206 318
rect 204 317 205 318
rect 203 317 204 318
rect 202 317 203 318
rect 201 317 202 318
rect 200 317 201 318
rect 199 317 200 318
rect 198 317 199 318
rect 197 317 198 318
rect 196 317 197 318
rect 195 317 196 318
rect 194 317 195 318
rect 193 317 194 318
rect 136 317 137 318
rect 135 317 136 318
rect 134 317 135 318
rect 133 317 134 318
rect 132 317 133 318
rect 131 317 132 318
rect 130 317 131 318
rect 129 317 130 318
rect 128 317 129 318
rect 127 317 128 318
rect 126 317 127 318
rect 125 317 126 318
rect 124 317 125 318
rect 123 317 124 318
rect 122 317 123 318
rect 121 317 122 318
rect 120 317 121 318
rect 119 317 120 318
rect 118 317 119 318
rect 117 317 118 318
rect 116 317 117 318
rect 115 317 116 318
rect 114 317 115 318
rect 113 317 114 318
rect 112 317 113 318
rect 111 317 112 318
rect 110 317 111 318
rect 109 317 110 318
rect 108 317 109 318
rect 107 317 108 318
rect 106 317 107 318
rect 105 317 106 318
rect 104 317 105 318
rect 103 317 104 318
rect 102 317 103 318
rect 101 317 102 318
rect 100 317 101 318
rect 99 317 100 318
rect 98 317 99 318
rect 97 317 98 318
rect 96 317 97 318
rect 95 317 96 318
rect 94 317 95 318
rect 76 317 77 318
rect 75 317 76 318
rect 74 317 75 318
rect 73 317 74 318
rect 72 317 73 318
rect 71 317 72 318
rect 70 317 71 318
rect 69 317 70 318
rect 68 317 69 318
rect 67 317 68 318
rect 66 317 67 318
rect 65 317 66 318
rect 64 317 65 318
rect 63 317 64 318
rect 62 317 63 318
rect 61 317 62 318
rect 60 317 61 318
rect 59 317 60 318
rect 58 317 59 318
rect 57 317 58 318
rect 56 317 57 318
rect 55 317 56 318
rect 54 317 55 318
rect 53 317 54 318
rect 52 317 53 318
rect 51 317 52 318
rect 50 317 51 318
rect 49 317 50 318
rect 48 317 49 318
rect 47 317 48 318
rect 46 317 47 318
rect 34 317 35 318
rect 33 317 34 318
rect 32 317 33 318
rect 31 317 32 318
rect 30 317 31 318
rect 29 317 30 318
rect 28 317 29 318
rect 27 317 28 318
rect 26 317 27 318
rect 25 317 26 318
rect 24 317 25 318
rect 23 317 24 318
rect 22 317 23 318
rect 21 317 22 318
rect 20 317 21 318
rect 19 317 20 318
rect 18 317 19 318
rect 17 317 18 318
rect 16 317 17 318
rect 15 317 16 318
rect 480 318 481 319
rect 468 318 469 319
rect 467 318 468 319
rect 466 318 467 319
rect 465 318 466 319
rect 464 318 465 319
rect 463 318 464 319
rect 462 318 463 319
rect 461 318 462 319
rect 460 318 461 319
rect 439 318 440 319
rect 438 318 439 319
rect 437 318 438 319
rect 436 318 437 319
rect 398 318 399 319
rect 397 318 398 319
rect 396 318 397 319
rect 395 318 396 319
rect 237 318 238 319
rect 236 318 237 319
rect 235 318 236 319
rect 234 318 235 319
rect 233 318 234 319
rect 232 318 233 319
rect 231 318 232 319
rect 230 318 231 319
rect 229 318 230 319
rect 228 318 229 319
rect 227 318 228 319
rect 226 318 227 319
rect 225 318 226 319
rect 224 318 225 319
rect 223 318 224 319
rect 222 318 223 319
rect 221 318 222 319
rect 220 318 221 319
rect 219 318 220 319
rect 218 318 219 319
rect 217 318 218 319
rect 216 318 217 319
rect 215 318 216 319
rect 214 318 215 319
rect 213 318 214 319
rect 212 318 213 319
rect 211 318 212 319
rect 210 318 211 319
rect 209 318 210 319
rect 208 318 209 319
rect 207 318 208 319
rect 206 318 207 319
rect 205 318 206 319
rect 204 318 205 319
rect 203 318 204 319
rect 202 318 203 319
rect 201 318 202 319
rect 200 318 201 319
rect 199 318 200 319
rect 198 318 199 319
rect 197 318 198 319
rect 196 318 197 319
rect 195 318 196 319
rect 194 318 195 319
rect 193 318 194 319
rect 192 318 193 319
rect 137 318 138 319
rect 136 318 137 319
rect 135 318 136 319
rect 134 318 135 319
rect 133 318 134 319
rect 132 318 133 319
rect 131 318 132 319
rect 130 318 131 319
rect 129 318 130 319
rect 128 318 129 319
rect 127 318 128 319
rect 126 318 127 319
rect 125 318 126 319
rect 124 318 125 319
rect 123 318 124 319
rect 122 318 123 319
rect 121 318 122 319
rect 120 318 121 319
rect 119 318 120 319
rect 118 318 119 319
rect 117 318 118 319
rect 116 318 117 319
rect 115 318 116 319
rect 114 318 115 319
rect 113 318 114 319
rect 112 318 113 319
rect 111 318 112 319
rect 110 318 111 319
rect 109 318 110 319
rect 108 318 109 319
rect 107 318 108 319
rect 106 318 107 319
rect 105 318 106 319
rect 104 318 105 319
rect 103 318 104 319
rect 102 318 103 319
rect 101 318 102 319
rect 100 318 101 319
rect 99 318 100 319
rect 98 318 99 319
rect 97 318 98 319
rect 96 318 97 319
rect 95 318 96 319
rect 94 318 95 319
rect 76 318 77 319
rect 75 318 76 319
rect 74 318 75 319
rect 73 318 74 319
rect 72 318 73 319
rect 71 318 72 319
rect 70 318 71 319
rect 69 318 70 319
rect 68 318 69 319
rect 67 318 68 319
rect 66 318 67 319
rect 65 318 66 319
rect 64 318 65 319
rect 63 318 64 319
rect 62 318 63 319
rect 61 318 62 319
rect 60 318 61 319
rect 59 318 60 319
rect 58 318 59 319
rect 57 318 58 319
rect 56 318 57 319
rect 55 318 56 319
rect 54 318 55 319
rect 53 318 54 319
rect 52 318 53 319
rect 51 318 52 319
rect 50 318 51 319
rect 49 318 50 319
rect 48 318 49 319
rect 47 318 48 319
rect 46 318 47 319
rect 35 318 36 319
rect 34 318 35 319
rect 33 318 34 319
rect 32 318 33 319
rect 31 318 32 319
rect 30 318 31 319
rect 29 318 30 319
rect 28 318 29 319
rect 27 318 28 319
rect 26 318 27 319
rect 25 318 26 319
rect 24 318 25 319
rect 23 318 24 319
rect 22 318 23 319
rect 21 318 22 319
rect 20 318 21 319
rect 19 318 20 319
rect 18 318 19 319
rect 17 318 18 319
rect 16 318 17 319
rect 480 319 481 320
rect 479 319 480 320
rect 470 319 471 320
rect 469 319 470 320
rect 468 319 469 320
rect 467 319 468 320
rect 466 319 467 320
rect 465 319 466 320
rect 464 319 465 320
rect 463 319 464 320
rect 462 319 463 320
rect 461 319 462 320
rect 460 319 461 320
rect 439 319 440 320
rect 438 319 439 320
rect 437 319 438 320
rect 397 319 398 320
rect 396 319 397 320
rect 395 319 396 320
rect 234 319 235 320
rect 233 319 234 320
rect 232 319 233 320
rect 231 319 232 320
rect 230 319 231 320
rect 229 319 230 320
rect 228 319 229 320
rect 227 319 228 320
rect 226 319 227 320
rect 225 319 226 320
rect 224 319 225 320
rect 223 319 224 320
rect 222 319 223 320
rect 221 319 222 320
rect 220 319 221 320
rect 219 319 220 320
rect 218 319 219 320
rect 217 319 218 320
rect 216 319 217 320
rect 215 319 216 320
rect 214 319 215 320
rect 213 319 214 320
rect 212 319 213 320
rect 211 319 212 320
rect 210 319 211 320
rect 209 319 210 320
rect 208 319 209 320
rect 207 319 208 320
rect 206 319 207 320
rect 205 319 206 320
rect 204 319 205 320
rect 203 319 204 320
rect 202 319 203 320
rect 201 319 202 320
rect 200 319 201 320
rect 199 319 200 320
rect 198 319 199 320
rect 197 319 198 320
rect 196 319 197 320
rect 195 319 196 320
rect 194 319 195 320
rect 193 319 194 320
rect 192 319 193 320
rect 191 319 192 320
rect 138 319 139 320
rect 137 319 138 320
rect 136 319 137 320
rect 135 319 136 320
rect 134 319 135 320
rect 133 319 134 320
rect 132 319 133 320
rect 131 319 132 320
rect 130 319 131 320
rect 129 319 130 320
rect 128 319 129 320
rect 127 319 128 320
rect 126 319 127 320
rect 125 319 126 320
rect 124 319 125 320
rect 123 319 124 320
rect 122 319 123 320
rect 121 319 122 320
rect 120 319 121 320
rect 119 319 120 320
rect 118 319 119 320
rect 117 319 118 320
rect 116 319 117 320
rect 115 319 116 320
rect 114 319 115 320
rect 113 319 114 320
rect 112 319 113 320
rect 111 319 112 320
rect 110 319 111 320
rect 109 319 110 320
rect 108 319 109 320
rect 107 319 108 320
rect 106 319 107 320
rect 105 319 106 320
rect 104 319 105 320
rect 103 319 104 320
rect 102 319 103 320
rect 101 319 102 320
rect 100 319 101 320
rect 99 319 100 320
rect 98 319 99 320
rect 97 319 98 320
rect 96 319 97 320
rect 95 319 96 320
rect 77 319 78 320
rect 76 319 77 320
rect 75 319 76 320
rect 74 319 75 320
rect 73 319 74 320
rect 72 319 73 320
rect 71 319 72 320
rect 70 319 71 320
rect 69 319 70 320
rect 68 319 69 320
rect 67 319 68 320
rect 66 319 67 320
rect 65 319 66 320
rect 64 319 65 320
rect 63 319 64 320
rect 62 319 63 320
rect 61 319 62 320
rect 60 319 61 320
rect 59 319 60 320
rect 58 319 59 320
rect 57 319 58 320
rect 56 319 57 320
rect 55 319 56 320
rect 54 319 55 320
rect 53 319 54 320
rect 52 319 53 320
rect 51 319 52 320
rect 50 319 51 320
rect 49 319 50 320
rect 48 319 49 320
rect 47 319 48 320
rect 35 319 36 320
rect 34 319 35 320
rect 33 319 34 320
rect 32 319 33 320
rect 31 319 32 320
rect 30 319 31 320
rect 29 319 30 320
rect 28 319 29 320
rect 27 319 28 320
rect 26 319 27 320
rect 25 319 26 320
rect 24 319 25 320
rect 23 319 24 320
rect 22 319 23 320
rect 21 319 22 320
rect 20 319 21 320
rect 19 319 20 320
rect 18 319 19 320
rect 17 319 18 320
rect 16 319 17 320
rect 480 320 481 321
rect 479 320 480 321
rect 478 320 479 321
rect 477 320 478 321
rect 476 320 477 321
rect 475 320 476 321
rect 474 320 475 321
rect 473 320 474 321
rect 472 320 473 321
rect 471 320 472 321
rect 470 320 471 321
rect 469 320 470 321
rect 468 320 469 321
rect 467 320 468 321
rect 466 320 467 321
rect 465 320 466 321
rect 464 320 465 321
rect 460 320 461 321
rect 439 320 440 321
rect 438 320 439 321
rect 437 320 438 321
rect 397 320 398 321
rect 396 320 397 321
rect 395 320 396 321
rect 230 320 231 321
rect 229 320 230 321
rect 228 320 229 321
rect 227 320 228 321
rect 226 320 227 321
rect 225 320 226 321
rect 224 320 225 321
rect 223 320 224 321
rect 222 320 223 321
rect 221 320 222 321
rect 220 320 221 321
rect 219 320 220 321
rect 218 320 219 321
rect 217 320 218 321
rect 216 320 217 321
rect 215 320 216 321
rect 214 320 215 321
rect 213 320 214 321
rect 212 320 213 321
rect 211 320 212 321
rect 210 320 211 321
rect 209 320 210 321
rect 208 320 209 321
rect 207 320 208 321
rect 206 320 207 321
rect 205 320 206 321
rect 204 320 205 321
rect 203 320 204 321
rect 202 320 203 321
rect 201 320 202 321
rect 200 320 201 321
rect 199 320 200 321
rect 198 320 199 321
rect 197 320 198 321
rect 196 320 197 321
rect 195 320 196 321
rect 194 320 195 321
rect 193 320 194 321
rect 192 320 193 321
rect 191 320 192 321
rect 190 320 191 321
rect 140 320 141 321
rect 139 320 140 321
rect 138 320 139 321
rect 137 320 138 321
rect 136 320 137 321
rect 135 320 136 321
rect 134 320 135 321
rect 133 320 134 321
rect 132 320 133 321
rect 131 320 132 321
rect 130 320 131 321
rect 129 320 130 321
rect 128 320 129 321
rect 127 320 128 321
rect 126 320 127 321
rect 125 320 126 321
rect 124 320 125 321
rect 123 320 124 321
rect 122 320 123 321
rect 121 320 122 321
rect 120 320 121 321
rect 119 320 120 321
rect 118 320 119 321
rect 117 320 118 321
rect 116 320 117 321
rect 115 320 116 321
rect 114 320 115 321
rect 113 320 114 321
rect 112 320 113 321
rect 111 320 112 321
rect 110 320 111 321
rect 109 320 110 321
rect 108 320 109 321
rect 107 320 108 321
rect 106 320 107 321
rect 105 320 106 321
rect 104 320 105 321
rect 103 320 104 321
rect 102 320 103 321
rect 101 320 102 321
rect 100 320 101 321
rect 99 320 100 321
rect 98 320 99 321
rect 97 320 98 321
rect 96 320 97 321
rect 77 320 78 321
rect 76 320 77 321
rect 75 320 76 321
rect 74 320 75 321
rect 73 320 74 321
rect 72 320 73 321
rect 71 320 72 321
rect 70 320 71 321
rect 69 320 70 321
rect 68 320 69 321
rect 67 320 68 321
rect 66 320 67 321
rect 65 320 66 321
rect 64 320 65 321
rect 63 320 64 321
rect 62 320 63 321
rect 61 320 62 321
rect 60 320 61 321
rect 59 320 60 321
rect 58 320 59 321
rect 57 320 58 321
rect 56 320 57 321
rect 55 320 56 321
rect 54 320 55 321
rect 53 320 54 321
rect 52 320 53 321
rect 51 320 52 321
rect 50 320 51 321
rect 49 320 50 321
rect 48 320 49 321
rect 47 320 48 321
rect 35 320 36 321
rect 34 320 35 321
rect 33 320 34 321
rect 32 320 33 321
rect 31 320 32 321
rect 30 320 31 321
rect 29 320 30 321
rect 28 320 29 321
rect 27 320 28 321
rect 26 320 27 321
rect 25 320 26 321
rect 24 320 25 321
rect 23 320 24 321
rect 22 320 23 321
rect 21 320 22 321
rect 20 320 21 321
rect 19 320 20 321
rect 18 320 19 321
rect 17 320 18 321
rect 480 321 481 322
rect 479 321 480 322
rect 478 321 479 322
rect 477 321 478 322
rect 476 321 477 322
rect 475 321 476 322
rect 474 321 475 322
rect 473 321 474 322
rect 472 321 473 322
rect 471 321 472 322
rect 470 321 471 322
rect 469 321 470 322
rect 468 321 469 322
rect 467 321 468 322
rect 466 321 467 322
rect 460 321 461 322
rect 439 321 440 322
rect 438 321 439 322
rect 437 321 438 322
rect 397 321 398 322
rect 396 321 397 322
rect 395 321 396 322
rect 226 321 227 322
rect 225 321 226 322
rect 224 321 225 322
rect 223 321 224 322
rect 222 321 223 322
rect 221 321 222 322
rect 220 321 221 322
rect 219 321 220 322
rect 218 321 219 322
rect 217 321 218 322
rect 216 321 217 322
rect 215 321 216 322
rect 214 321 215 322
rect 213 321 214 322
rect 212 321 213 322
rect 211 321 212 322
rect 210 321 211 322
rect 209 321 210 322
rect 208 321 209 322
rect 207 321 208 322
rect 206 321 207 322
rect 205 321 206 322
rect 204 321 205 322
rect 203 321 204 322
rect 202 321 203 322
rect 201 321 202 322
rect 200 321 201 322
rect 199 321 200 322
rect 198 321 199 322
rect 197 321 198 322
rect 196 321 197 322
rect 195 321 196 322
rect 194 321 195 322
rect 193 321 194 322
rect 142 321 143 322
rect 141 321 142 322
rect 140 321 141 322
rect 139 321 140 322
rect 138 321 139 322
rect 137 321 138 322
rect 136 321 137 322
rect 135 321 136 322
rect 134 321 135 322
rect 133 321 134 322
rect 132 321 133 322
rect 131 321 132 322
rect 130 321 131 322
rect 129 321 130 322
rect 128 321 129 322
rect 127 321 128 322
rect 126 321 127 322
rect 125 321 126 322
rect 124 321 125 322
rect 123 321 124 322
rect 122 321 123 322
rect 121 321 122 322
rect 120 321 121 322
rect 119 321 120 322
rect 118 321 119 322
rect 117 321 118 322
rect 116 321 117 322
rect 115 321 116 322
rect 114 321 115 322
rect 113 321 114 322
rect 112 321 113 322
rect 111 321 112 322
rect 110 321 111 322
rect 109 321 110 322
rect 108 321 109 322
rect 107 321 108 322
rect 106 321 107 322
rect 105 321 106 322
rect 104 321 105 322
rect 103 321 104 322
rect 102 321 103 322
rect 101 321 102 322
rect 100 321 101 322
rect 99 321 100 322
rect 98 321 99 322
rect 97 321 98 322
rect 78 321 79 322
rect 77 321 78 322
rect 76 321 77 322
rect 75 321 76 322
rect 74 321 75 322
rect 73 321 74 322
rect 72 321 73 322
rect 71 321 72 322
rect 70 321 71 322
rect 69 321 70 322
rect 68 321 69 322
rect 67 321 68 322
rect 66 321 67 322
rect 65 321 66 322
rect 64 321 65 322
rect 63 321 64 322
rect 62 321 63 322
rect 61 321 62 322
rect 60 321 61 322
rect 59 321 60 322
rect 58 321 59 322
rect 57 321 58 322
rect 56 321 57 322
rect 55 321 56 322
rect 54 321 55 322
rect 53 321 54 322
rect 52 321 53 322
rect 51 321 52 322
rect 50 321 51 322
rect 49 321 50 322
rect 48 321 49 322
rect 47 321 48 322
rect 35 321 36 322
rect 34 321 35 322
rect 33 321 34 322
rect 32 321 33 322
rect 31 321 32 322
rect 30 321 31 322
rect 29 321 30 322
rect 28 321 29 322
rect 27 321 28 322
rect 26 321 27 322
rect 25 321 26 322
rect 24 321 25 322
rect 23 321 24 322
rect 22 321 23 322
rect 21 321 22 322
rect 20 321 21 322
rect 19 321 20 322
rect 18 321 19 322
rect 480 322 481 323
rect 479 322 480 323
rect 478 322 479 323
rect 477 322 478 323
rect 476 322 477 323
rect 475 322 476 323
rect 474 322 475 323
rect 473 322 474 323
rect 472 322 473 323
rect 471 322 472 323
rect 470 322 471 323
rect 469 322 470 323
rect 468 322 469 323
rect 439 322 440 323
rect 438 322 439 323
rect 437 322 438 323
rect 397 322 398 323
rect 396 322 397 323
rect 395 322 396 323
rect 219 322 220 323
rect 218 322 219 323
rect 217 322 218 323
rect 216 322 217 323
rect 215 322 216 323
rect 214 322 215 323
rect 213 322 214 323
rect 212 322 213 323
rect 211 322 212 323
rect 210 322 211 323
rect 209 322 210 323
rect 208 322 209 323
rect 207 322 208 323
rect 206 322 207 323
rect 205 322 206 323
rect 204 322 205 323
rect 203 322 204 323
rect 202 322 203 323
rect 201 322 202 323
rect 200 322 201 323
rect 143 322 144 323
rect 142 322 143 323
rect 141 322 142 323
rect 140 322 141 323
rect 139 322 140 323
rect 138 322 139 323
rect 137 322 138 323
rect 136 322 137 323
rect 135 322 136 323
rect 134 322 135 323
rect 133 322 134 323
rect 132 322 133 323
rect 131 322 132 323
rect 130 322 131 323
rect 129 322 130 323
rect 128 322 129 323
rect 127 322 128 323
rect 126 322 127 323
rect 125 322 126 323
rect 124 322 125 323
rect 123 322 124 323
rect 122 322 123 323
rect 121 322 122 323
rect 120 322 121 323
rect 119 322 120 323
rect 118 322 119 323
rect 117 322 118 323
rect 116 322 117 323
rect 115 322 116 323
rect 114 322 115 323
rect 113 322 114 323
rect 112 322 113 323
rect 111 322 112 323
rect 110 322 111 323
rect 109 322 110 323
rect 108 322 109 323
rect 107 322 108 323
rect 106 322 107 323
rect 105 322 106 323
rect 104 322 105 323
rect 103 322 104 323
rect 102 322 103 323
rect 101 322 102 323
rect 100 322 101 323
rect 99 322 100 323
rect 98 322 99 323
rect 97 322 98 323
rect 79 322 80 323
rect 78 322 79 323
rect 77 322 78 323
rect 76 322 77 323
rect 75 322 76 323
rect 74 322 75 323
rect 73 322 74 323
rect 72 322 73 323
rect 71 322 72 323
rect 70 322 71 323
rect 69 322 70 323
rect 68 322 69 323
rect 67 322 68 323
rect 66 322 67 323
rect 65 322 66 323
rect 64 322 65 323
rect 63 322 64 323
rect 62 322 63 323
rect 61 322 62 323
rect 60 322 61 323
rect 59 322 60 323
rect 58 322 59 323
rect 57 322 58 323
rect 56 322 57 323
rect 55 322 56 323
rect 54 322 55 323
rect 53 322 54 323
rect 52 322 53 323
rect 51 322 52 323
rect 50 322 51 323
rect 49 322 50 323
rect 48 322 49 323
rect 36 322 37 323
rect 35 322 36 323
rect 34 322 35 323
rect 33 322 34 323
rect 32 322 33 323
rect 31 322 32 323
rect 30 322 31 323
rect 29 322 30 323
rect 28 322 29 323
rect 27 322 28 323
rect 26 322 27 323
rect 25 322 26 323
rect 24 322 25 323
rect 23 322 24 323
rect 22 322 23 323
rect 21 322 22 323
rect 20 322 21 323
rect 19 322 20 323
rect 18 322 19 323
rect 480 323 481 324
rect 479 323 480 324
rect 478 323 479 324
rect 477 323 478 324
rect 476 323 477 324
rect 475 323 476 324
rect 474 323 475 324
rect 473 323 474 324
rect 472 323 473 324
rect 471 323 472 324
rect 470 323 471 324
rect 469 323 470 324
rect 145 323 146 324
rect 144 323 145 324
rect 143 323 144 324
rect 142 323 143 324
rect 141 323 142 324
rect 140 323 141 324
rect 139 323 140 324
rect 138 323 139 324
rect 137 323 138 324
rect 136 323 137 324
rect 135 323 136 324
rect 134 323 135 324
rect 133 323 134 324
rect 132 323 133 324
rect 131 323 132 324
rect 130 323 131 324
rect 129 323 130 324
rect 128 323 129 324
rect 127 323 128 324
rect 126 323 127 324
rect 125 323 126 324
rect 124 323 125 324
rect 123 323 124 324
rect 122 323 123 324
rect 121 323 122 324
rect 120 323 121 324
rect 119 323 120 324
rect 118 323 119 324
rect 117 323 118 324
rect 116 323 117 324
rect 115 323 116 324
rect 114 323 115 324
rect 113 323 114 324
rect 112 323 113 324
rect 111 323 112 324
rect 110 323 111 324
rect 109 323 110 324
rect 108 323 109 324
rect 107 323 108 324
rect 106 323 107 324
rect 105 323 106 324
rect 104 323 105 324
rect 103 323 104 324
rect 102 323 103 324
rect 101 323 102 324
rect 100 323 101 324
rect 99 323 100 324
rect 98 323 99 324
rect 79 323 80 324
rect 78 323 79 324
rect 77 323 78 324
rect 76 323 77 324
rect 75 323 76 324
rect 74 323 75 324
rect 73 323 74 324
rect 72 323 73 324
rect 71 323 72 324
rect 70 323 71 324
rect 69 323 70 324
rect 68 323 69 324
rect 67 323 68 324
rect 66 323 67 324
rect 65 323 66 324
rect 64 323 65 324
rect 63 323 64 324
rect 62 323 63 324
rect 61 323 62 324
rect 60 323 61 324
rect 59 323 60 324
rect 58 323 59 324
rect 57 323 58 324
rect 56 323 57 324
rect 55 323 56 324
rect 54 323 55 324
rect 53 323 54 324
rect 52 323 53 324
rect 51 323 52 324
rect 50 323 51 324
rect 49 323 50 324
rect 48 323 49 324
rect 36 323 37 324
rect 35 323 36 324
rect 34 323 35 324
rect 33 323 34 324
rect 32 323 33 324
rect 31 323 32 324
rect 30 323 31 324
rect 29 323 30 324
rect 28 323 29 324
rect 27 323 28 324
rect 26 323 27 324
rect 25 323 26 324
rect 24 323 25 324
rect 23 323 24 324
rect 22 323 23 324
rect 21 323 22 324
rect 20 323 21 324
rect 19 323 20 324
rect 480 324 481 325
rect 479 324 480 325
rect 478 324 479 325
rect 477 324 478 325
rect 476 324 477 325
rect 475 324 476 325
rect 474 324 475 325
rect 473 324 474 325
rect 472 324 473 325
rect 471 324 472 325
rect 470 324 471 325
rect 469 324 470 325
rect 468 324 469 325
rect 147 324 148 325
rect 146 324 147 325
rect 145 324 146 325
rect 144 324 145 325
rect 143 324 144 325
rect 142 324 143 325
rect 141 324 142 325
rect 140 324 141 325
rect 139 324 140 325
rect 138 324 139 325
rect 137 324 138 325
rect 136 324 137 325
rect 135 324 136 325
rect 134 324 135 325
rect 133 324 134 325
rect 132 324 133 325
rect 131 324 132 325
rect 130 324 131 325
rect 129 324 130 325
rect 128 324 129 325
rect 127 324 128 325
rect 126 324 127 325
rect 125 324 126 325
rect 124 324 125 325
rect 123 324 124 325
rect 122 324 123 325
rect 121 324 122 325
rect 120 324 121 325
rect 119 324 120 325
rect 118 324 119 325
rect 117 324 118 325
rect 116 324 117 325
rect 115 324 116 325
rect 114 324 115 325
rect 113 324 114 325
rect 112 324 113 325
rect 111 324 112 325
rect 110 324 111 325
rect 109 324 110 325
rect 108 324 109 325
rect 107 324 108 325
rect 106 324 107 325
rect 105 324 106 325
rect 104 324 105 325
rect 103 324 104 325
rect 102 324 103 325
rect 101 324 102 325
rect 100 324 101 325
rect 99 324 100 325
rect 80 324 81 325
rect 79 324 80 325
rect 78 324 79 325
rect 77 324 78 325
rect 76 324 77 325
rect 75 324 76 325
rect 74 324 75 325
rect 73 324 74 325
rect 72 324 73 325
rect 71 324 72 325
rect 70 324 71 325
rect 69 324 70 325
rect 68 324 69 325
rect 67 324 68 325
rect 66 324 67 325
rect 65 324 66 325
rect 64 324 65 325
rect 63 324 64 325
rect 62 324 63 325
rect 61 324 62 325
rect 60 324 61 325
rect 59 324 60 325
rect 58 324 59 325
rect 57 324 58 325
rect 56 324 57 325
rect 55 324 56 325
rect 54 324 55 325
rect 53 324 54 325
rect 52 324 53 325
rect 51 324 52 325
rect 50 324 51 325
rect 49 324 50 325
rect 48 324 49 325
rect 36 324 37 325
rect 35 324 36 325
rect 34 324 35 325
rect 33 324 34 325
rect 32 324 33 325
rect 31 324 32 325
rect 30 324 31 325
rect 29 324 30 325
rect 28 324 29 325
rect 27 324 28 325
rect 26 324 27 325
rect 25 324 26 325
rect 24 324 25 325
rect 23 324 24 325
rect 22 324 23 325
rect 21 324 22 325
rect 20 324 21 325
rect 480 325 481 326
rect 469 325 470 326
rect 468 325 469 326
rect 467 325 468 326
rect 466 325 467 326
rect 460 325 461 326
rect 149 325 150 326
rect 148 325 149 326
rect 147 325 148 326
rect 146 325 147 326
rect 145 325 146 326
rect 144 325 145 326
rect 143 325 144 326
rect 142 325 143 326
rect 141 325 142 326
rect 140 325 141 326
rect 139 325 140 326
rect 138 325 139 326
rect 137 325 138 326
rect 136 325 137 326
rect 135 325 136 326
rect 134 325 135 326
rect 133 325 134 326
rect 132 325 133 326
rect 131 325 132 326
rect 130 325 131 326
rect 129 325 130 326
rect 128 325 129 326
rect 127 325 128 326
rect 126 325 127 326
rect 125 325 126 326
rect 124 325 125 326
rect 123 325 124 326
rect 122 325 123 326
rect 121 325 122 326
rect 120 325 121 326
rect 119 325 120 326
rect 118 325 119 326
rect 117 325 118 326
rect 116 325 117 326
rect 115 325 116 326
rect 114 325 115 326
rect 113 325 114 326
rect 112 325 113 326
rect 111 325 112 326
rect 110 325 111 326
rect 109 325 110 326
rect 108 325 109 326
rect 107 325 108 326
rect 106 325 107 326
rect 105 325 106 326
rect 104 325 105 326
rect 103 325 104 326
rect 102 325 103 326
rect 101 325 102 326
rect 100 325 101 326
rect 80 325 81 326
rect 79 325 80 326
rect 78 325 79 326
rect 77 325 78 326
rect 76 325 77 326
rect 75 325 76 326
rect 74 325 75 326
rect 73 325 74 326
rect 72 325 73 326
rect 71 325 72 326
rect 70 325 71 326
rect 69 325 70 326
rect 68 325 69 326
rect 67 325 68 326
rect 66 325 67 326
rect 65 325 66 326
rect 64 325 65 326
rect 63 325 64 326
rect 62 325 63 326
rect 61 325 62 326
rect 60 325 61 326
rect 59 325 60 326
rect 58 325 59 326
rect 57 325 58 326
rect 56 325 57 326
rect 55 325 56 326
rect 54 325 55 326
rect 53 325 54 326
rect 52 325 53 326
rect 51 325 52 326
rect 50 325 51 326
rect 49 325 50 326
rect 37 325 38 326
rect 36 325 37 326
rect 35 325 36 326
rect 34 325 35 326
rect 33 325 34 326
rect 32 325 33 326
rect 31 325 32 326
rect 30 325 31 326
rect 29 325 30 326
rect 28 325 29 326
rect 27 325 28 326
rect 26 325 27 326
rect 25 325 26 326
rect 24 325 25 326
rect 23 325 24 326
rect 22 325 23 326
rect 21 325 22 326
rect 480 326 481 327
rect 467 326 468 327
rect 466 326 467 327
rect 465 326 466 327
rect 464 326 465 327
rect 460 326 461 327
rect 151 326 152 327
rect 150 326 151 327
rect 149 326 150 327
rect 148 326 149 327
rect 147 326 148 327
rect 146 326 147 327
rect 145 326 146 327
rect 144 326 145 327
rect 143 326 144 327
rect 142 326 143 327
rect 141 326 142 327
rect 140 326 141 327
rect 139 326 140 327
rect 138 326 139 327
rect 137 326 138 327
rect 136 326 137 327
rect 135 326 136 327
rect 134 326 135 327
rect 133 326 134 327
rect 132 326 133 327
rect 131 326 132 327
rect 130 326 131 327
rect 129 326 130 327
rect 128 326 129 327
rect 127 326 128 327
rect 126 326 127 327
rect 125 326 126 327
rect 124 326 125 327
rect 123 326 124 327
rect 122 326 123 327
rect 121 326 122 327
rect 120 326 121 327
rect 119 326 120 327
rect 118 326 119 327
rect 117 326 118 327
rect 116 326 117 327
rect 115 326 116 327
rect 114 326 115 327
rect 113 326 114 327
rect 112 326 113 327
rect 111 326 112 327
rect 110 326 111 327
rect 109 326 110 327
rect 108 326 109 327
rect 107 326 108 327
rect 106 326 107 327
rect 105 326 106 327
rect 104 326 105 327
rect 103 326 104 327
rect 102 326 103 327
rect 101 326 102 327
rect 100 326 101 327
rect 81 326 82 327
rect 80 326 81 327
rect 79 326 80 327
rect 78 326 79 327
rect 77 326 78 327
rect 76 326 77 327
rect 75 326 76 327
rect 74 326 75 327
rect 73 326 74 327
rect 72 326 73 327
rect 71 326 72 327
rect 70 326 71 327
rect 69 326 70 327
rect 68 326 69 327
rect 67 326 68 327
rect 66 326 67 327
rect 65 326 66 327
rect 64 326 65 327
rect 63 326 64 327
rect 62 326 63 327
rect 61 326 62 327
rect 60 326 61 327
rect 59 326 60 327
rect 58 326 59 327
rect 57 326 58 327
rect 56 326 57 327
rect 55 326 56 327
rect 54 326 55 327
rect 53 326 54 327
rect 52 326 53 327
rect 51 326 52 327
rect 50 326 51 327
rect 49 326 50 327
rect 37 326 38 327
rect 36 326 37 327
rect 35 326 36 327
rect 34 326 35 327
rect 33 326 34 327
rect 32 326 33 327
rect 31 326 32 327
rect 30 326 31 327
rect 29 326 30 327
rect 28 326 29 327
rect 27 326 28 327
rect 26 326 27 327
rect 25 326 26 327
rect 24 326 25 327
rect 23 326 24 327
rect 22 326 23 327
rect 480 327 481 328
rect 465 327 466 328
rect 464 327 465 328
rect 463 327 464 328
rect 462 327 463 328
rect 461 327 462 328
rect 460 327 461 328
rect 153 327 154 328
rect 152 327 153 328
rect 151 327 152 328
rect 150 327 151 328
rect 149 327 150 328
rect 148 327 149 328
rect 147 327 148 328
rect 146 327 147 328
rect 145 327 146 328
rect 144 327 145 328
rect 143 327 144 328
rect 142 327 143 328
rect 141 327 142 328
rect 140 327 141 328
rect 139 327 140 328
rect 138 327 139 328
rect 137 327 138 328
rect 136 327 137 328
rect 135 327 136 328
rect 134 327 135 328
rect 133 327 134 328
rect 132 327 133 328
rect 131 327 132 328
rect 130 327 131 328
rect 129 327 130 328
rect 128 327 129 328
rect 127 327 128 328
rect 126 327 127 328
rect 125 327 126 328
rect 124 327 125 328
rect 123 327 124 328
rect 122 327 123 328
rect 121 327 122 328
rect 120 327 121 328
rect 119 327 120 328
rect 118 327 119 328
rect 117 327 118 328
rect 116 327 117 328
rect 115 327 116 328
rect 114 327 115 328
rect 113 327 114 328
rect 112 327 113 328
rect 111 327 112 328
rect 110 327 111 328
rect 109 327 110 328
rect 108 327 109 328
rect 107 327 108 328
rect 106 327 107 328
rect 105 327 106 328
rect 104 327 105 328
rect 103 327 104 328
rect 102 327 103 328
rect 101 327 102 328
rect 82 327 83 328
rect 81 327 82 328
rect 80 327 81 328
rect 79 327 80 328
rect 78 327 79 328
rect 77 327 78 328
rect 76 327 77 328
rect 75 327 76 328
rect 74 327 75 328
rect 73 327 74 328
rect 72 327 73 328
rect 71 327 72 328
rect 70 327 71 328
rect 69 327 70 328
rect 68 327 69 328
rect 67 327 68 328
rect 66 327 67 328
rect 65 327 66 328
rect 64 327 65 328
rect 63 327 64 328
rect 62 327 63 328
rect 61 327 62 328
rect 60 327 61 328
rect 59 327 60 328
rect 58 327 59 328
rect 57 327 58 328
rect 56 327 57 328
rect 55 327 56 328
rect 54 327 55 328
rect 53 327 54 328
rect 52 327 53 328
rect 51 327 52 328
rect 50 327 51 328
rect 37 327 38 328
rect 36 327 37 328
rect 35 327 36 328
rect 34 327 35 328
rect 33 327 34 328
rect 32 327 33 328
rect 31 327 32 328
rect 30 327 31 328
rect 29 327 30 328
rect 28 327 29 328
rect 27 327 28 328
rect 26 327 27 328
rect 25 327 26 328
rect 24 327 25 328
rect 23 327 24 328
rect 22 327 23 328
rect 463 328 464 329
rect 462 328 463 329
rect 461 328 462 329
rect 460 328 461 329
rect 156 328 157 329
rect 155 328 156 329
rect 154 328 155 329
rect 153 328 154 329
rect 152 328 153 329
rect 151 328 152 329
rect 150 328 151 329
rect 149 328 150 329
rect 148 328 149 329
rect 147 328 148 329
rect 146 328 147 329
rect 145 328 146 329
rect 144 328 145 329
rect 143 328 144 329
rect 142 328 143 329
rect 141 328 142 329
rect 140 328 141 329
rect 139 328 140 329
rect 138 328 139 329
rect 137 328 138 329
rect 136 328 137 329
rect 135 328 136 329
rect 134 328 135 329
rect 133 328 134 329
rect 132 328 133 329
rect 131 328 132 329
rect 130 328 131 329
rect 129 328 130 329
rect 128 328 129 329
rect 127 328 128 329
rect 126 328 127 329
rect 125 328 126 329
rect 124 328 125 329
rect 123 328 124 329
rect 122 328 123 329
rect 121 328 122 329
rect 120 328 121 329
rect 119 328 120 329
rect 118 328 119 329
rect 117 328 118 329
rect 116 328 117 329
rect 115 328 116 329
rect 114 328 115 329
rect 113 328 114 329
rect 112 328 113 329
rect 111 328 112 329
rect 110 328 111 329
rect 109 328 110 329
rect 108 328 109 329
rect 107 328 108 329
rect 106 328 107 329
rect 105 328 106 329
rect 104 328 105 329
rect 103 328 104 329
rect 102 328 103 329
rect 82 328 83 329
rect 81 328 82 329
rect 80 328 81 329
rect 79 328 80 329
rect 78 328 79 329
rect 77 328 78 329
rect 76 328 77 329
rect 75 328 76 329
rect 74 328 75 329
rect 73 328 74 329
rect 72 328 73 329
rect 71 328 72 329
rect 70 328 71 329
rect 69 328 70 329
rect 68 328 69 329
rect 67 328 68 329
rect 66 328 67 329
rect 65 328 66 329
rect 64 328 65 329
rect 63 328 64 329
rect 62 328 63 329
rect 61 328 62 329
rect 60 328 61 329
rect 59 328 60 329
rect 58 328 59 329
rect 57 328 58 329
rect 56 328 57 329
rect 55 328 56 329
rect 54 328 55 329
rect 53 328 54 329
rect 52 328 53 329
rect 51 328 52 329
rect 50 328 51 329
rect 38 328 39 329
rect 37 328 38 329
rect 36 328 37 329
rect 35 328 36 329
rect 34 328 35 329
rect 33 328 34 329
rect 32 328 33 329
rect 31 328 32 329
rect 30 328 31 329
rect 29 328 30 329
rect 28 328 29 329
rect 27 328 28 329
rect 26 328 27 329
rect 25 328 26 329
rect 24 328 25 329
rect 23 328 24 329
rect 462 329 463 330
rect 461 329 462 330
rect 460 329 461 330
rect 158 329 159 330
rect 157 329 158 330
rect 156 329 157 330
rect 155 329 156 330
rect 154 329 155 330
rect 153 329 154 330
rect 152 329 153 330
rect 151 329 152 330
rect 150 329 151 330
rect 149 329 150 330
rect 148 329 149 330
rect 147 329 148 330
rect 146 329 147 330
rect 145 329 146 330
rect 144 329 145 330
rect 143 329 144 330
rect 142 329 143 330
rect 141 329 142 330
rect 140 329 141 330
rect 139 329 140 330
rect 138 329 139 330
rect 137 329 138 330
rect 136 329 137 330
rect 135 329 136 330
rect 134 329 135 330
rect 133 329 134 330
rect 132 329 133 330
rect 131 329 132 330
rect 130 329 131 330
rect 129 329 130 330
rect 128 329 129 330
rect 127 329 128 330
rect 126 329 127 330
rect 125 329 126 330
rect 124 329 125 330
rect 123 329 124 330
rect 122 329 123 330
rect 121 329 122 330
rect 120 329 121 330
rect 119 329 120 330
rect 118 329 119 330
rect 117 329 118 330
rect 116 329 117 330
rect 115 329 116 330
rect 114 329 115 330
rect 113 329 114 330
rect 112 329 113 330
rect 111 329 112 330
rect 110 329 111 330
rect 109 329 110 330
rect 108 329 109 330
rect 107 329 108 330
rect 106 329 107 330
rect 105 329 106 330
rect 104 329 105 330
rect 103 329 104 330
rect 83 329 84 330
rect 82 329 83 330
rect 81 329 82 330
rect 80 329 81 330
rect 79 329 80 330
rect 78 329 79 330
rect 77 329 78 330
rect 76 329 77 330
rect 75 329 76 330
rect 74 329 75 330
rect 73 329 74 330
rect 72 329 73 330
rect 71 329 72 330
rect 70 329 71 330
rect 69 329 70 330
rect 68 329 69 330
rect 67 329 68 330
rect 66 329 67 330
rect 65 329 66 330
rect 64 329 65 330
rect 63 329 64 330
rect 62 329 63 330
rect 61 329 62 330
rect 60 329 61 330
rect 59 329 60 330
rect 58 329 59 330
rect 57 329 58 330
rect 56 329 57 330
rect 55 329 56 330
rect 54 329 55 330
rect 53 329 54 330
rect 52 329 53 330
rect 51 329 52 330
rect 50 329 51 330
rect 38 329 39 330
rect 37 329 38 330
rect 36 329 37 330
rect 35 329 36 330
rect 34 329 35 330
rect 33 329 34 330
rect 32 329 33 330
rect 31 329 32 330
rect 30 329 31 330
rect 29 329 30 330
rect 28 329 29 330
rect 27 329 28 330
rect 26 329 27 330
rect 25 329 26 330
rect 24 329 25 330
rect 461 330 462 331
rect 460 330 461 331
rect 161 330 162 331
rect 160 330 161 331
rect 159 330 160 331
rect 158 330 159 331
rect 157 330 158 331
rect 156 330 157 331
rect 155 330 156 331
rect 154 330 155 331
rect 153 330 154 331
rect 152 330 153 331
rect 151 330 152 331
rect 150 330 151 331
rect 149 330 150 331
rect 148 330 149 331
rect 147 330 148 331
rect 146 330 147 331
rect 145 330 146 331
rect 144 330 145 331
rect 143 330 144 331
rect 142 330 143 331
rect 141 330 142 331
rect 140 330 141 331
rect 139 330 140 331
rect 138 330 139 331
rect 137 330 138 331
rect 136 330 137 331
rect 135 330 136 331
rect 134 330 135 331
rect 133 330 134 331
rect 132 330 133 331
rect 131 330 132 331
rect 130 330 131 331
rect 129 330 130 331
rect 128 330 129 331
rect 127 330 128 331
rect 126 330 127 331
rect 125 330 126 331
rect 124 330 125 331
rect 123 330 124 331
rect 122 330 123 331
rect 121 330 122 331
rect 120 330 121 331
rect 119 330 120 331
rect 118 330 119 331
rect 117 330 118 331
rect 116 330 117 331
rect 115 330 116 331
rect 114 330 115 331
rect 113 330 114 331
rect 112 330 113 331
rect 111 330 112 331
rect 110 330 111 331
rect 109 330 110 331
rect 108 330 109 331
rect 107 330 108 331
rect 106 330 107 331
rect 105 330 106 331
rect 104 330 105 331
rect 84 330 85 331
rect 83 330 84 331
rect 82 330 83 331
rect 81 330 82 331
rect 80 330 81 331
rect 79 330 80 331
rect 78 330 79 331
rect 77 330 78 331
rect 76 330 77 331
rect 75 330 76 331
rect 74 330 75 331
rect 73 330 74 331
rect 72 330 73 331
rect 71 330 72 331
rect 70 330 71 331
rect 69 330 70 331
rect 68 330 69 331
rect 67 330 68 331
rect 66 330 67 331
rect 65 330 66 331
rect 64 330 65 331
rect 63 330 64 331
rect 62 330 63 331
rect 61 330 62 331
rect 60 330 61 331
rect 59 330 60 331
rect 58 330 59 331
rect 57 330 58 331
rect 56 330 57 331
rect 55 330 56 331
rect 54 330 55 331
rect 53 330 54 331
rect 52 330 53 331
rect 51 330 52 331
rect 39 330 40 331
rect 38 330 39 331
rect 37 330 38 331
rect 36 330 37 331
rect 35 330 36 331
rect 34 330 35 331
rect 33 330 34 331
rect 32 330 33 331
rect 31 330 32 331
rect 30 330 31 331
rect 29 330 30 331
rect 28 330 29 331
rect 27 330 28 331
rect 26 330 27 331
rect 25 330 26 331
rect 460 331 461 332
rect 439 331 440 332
rect 438 331 439 332
rect 437 331 438 332
rect 164 331 165 332
rect 163 331 164 332
rect 162 331 163 332
rect 161 331 162 332
rect 160 331 161 332
rect 159 331 160 332
rect 158 331 159 332
rect 157 331 158 332
rect 156 331 157 332
rect 155 331 156 332
rect 154 331 155 332
rect 153 331 154 332
rect 152 331 153 332
rect 151 331 152 332
rect 150 331 151 332
rect 149 331 150 332
rect 148 331 149 332
rect 147 331 148 332
rect 146 331 147 332
rect 145 331 146 332
rect 144 331 145 332
rect 143 331 144 332
rect 142 331 143 332
rect 141 331 142 332
rect 140 331 141 332
rect 139 331 140 332
rect 138 331 139 332
rect 137 331 138 332
rect 136 331 137 332
rect 135 331 136 332
rect 134 331 135 332
rect 133 331 134 332
rect 132 331 133 332
rect 131 331 132 332
rect 130 331 131 332
rect 129 331 130 332
rect 128 331 129 332
rect 127 331 128 332
rect 126 331 127 332
rect 125 331 126 332
rect 124 331 125 332
rect 123 331 124 332
rect 122 331 123 332
rect 121 331 122 332
rect 120 331 121 332
rect 119 331 120 332
rect 118 331 119 332
rect 117 331 118 332
rect 116 331 117 332
rect 115 331 116 332
rect 114 331 115 332
rect 113 331 114 332
rect 112 331 113 332
rect 111 331 112 332
rect 110 331 111 332
rect 109 331 110 332
rect 108 331 109 332
rect 107 331 108 332
rect 106 331 107 332
rect 105 331 106 332
rect 104 331 105 332
rect 84 331 85 332
rect 83 331 84 332
rect 82 331 83 332
rect 81 331 82 332
rect 80 331 81 332
rect 79 331 80 332
rect 78 331 79 332
rect 77 331 78 332
rect 76 331 77 332
rect 75 331 76 332
rect 74 331 75 332
rect 73 331 74 332
rect 72 331 73 332
rect 71 331 72 332
rect 70 331 71 332
rect 69 331 70 332
rect 68 331 69 332
rect 67 331 68 332
rect 66 331 67 332
rect 65 331 66 332
rect 64 331 65 332
rect 63 331 64 332
rect 62 331 63 332
rect 61 331 62 332
rect 60 331 61 332
rect 59 331 60 332
rect 58 331 59 332
rect 57 331 58 332
rect 56 331 57 332
rect 55 331 56 332
rect 54 331 55 332
rect 53 331 54 332
rect 52 331 53 332
rect 51 331 52 332
rect 39 331 40 332
rect 38 331 39 332
rect 37 331 38 332
rect 36 331 37 332
rect 35 331 36 332
rect 34 331 35 332
rect 33 331 34 332
rect 32 331 33 332
rect 31 331 32 332
rect 30 331 31 332
rect 29 331 30 332
rect 28 331 29 332
rect 27 331 28 332
rect 26 331 27 332
rect 460 332 461 333
rect 439 332 440 333
rect 438 332 439 333
rect 437 332 438 333
rect 397 332 398 333
rect 396 332 397 333
rect 395 332 396 333
rect 167 332 168 333
rect 166 332 167 333
rect 165 332 166 333
rect 164 332 165 333
rect 163 332 164 333
rect 162 332 163 333
rect 161 332 162 333
rect 160 332 161 333
rect 159 332 160 333
rect 158 332 159 333
rect 157 332 158 333
rect 156 332 157 333
rect 155 332 156 333
rect 154 332 155 333
rect 153 332 154 333
rect 152 332 153 333
rect 151 332 152 333
rect 150 332 151 333
rect 149 332 150 333
rect 148 332 149 333
rect 147 332 148 333
rect 146 332 147 333
rect 145 332 146 333
rect 144 332 145 333
rect 143 332 144 333
rect 142 332 143 333
rect 141 332 142 333
rect 140 332 141 333
rect 139 332 140 333
rect 138 332 139 333
rect 137 332 138 333
rect 136 332 137 333
rect 135 332 136 333
rect 134 332 135 333
rect 133 332 134 333
rect 132 332 133 333
rect 131 332 132 333
rect 130 332 131 333
rect 129 332 130 333
rect 128 332 129 333
rect 127 332 128 333
rect 126 332 127 333
rect 125 332 126 333
rect 124 332 125 333
rect 123 332 124 333
rect 122 332 123 333
rect 121 332 122 333
rect 120 332 121 333
rect 119 332 120 333
rect 118 332 119 333
rect 117 332 118 333
rect 116 332 117 333
rect 115 332 116 333
rect 114 332 115 333
rect 113 332 114 333
rect 112 332 113 333
rect 111 332 112 333
rect 110 332 111 333
rect 109 332 110 333
rect 108 332 109 333
rect 107 332 108 333
rect 106 332 107 333
rect 105 332 106 333
rect 85 332 86 333
rect 84 332 85 333
rect 83 332 84 333
rect 82 332 83 333
rect 81 332 82 333
rect 80 332 81 333
rect 79 332 80 333
rect 78 332 79 333
rect 77 332 78 333
rect 76 332 77 333
rect 75 332 76 333
rect 74 332 75 333
rect 73 332 74 333
rect 72 332 73 333
rect 71 332 72 333
rect 70 332 71 333
rect 69 332 70 333
rect 68 332 69 333
rect 67 332 68 333
rect 66 332 67 333
rect 65 332 66 333
rect 64 332 65 333
rect 63 332 64 333
rect 62 332 63 333
rect 61 332 62 333
rect 60 332 61 333
rect 59 332 60 333
rect 58 332 59 333
rect 57 332 58 333
rect 56 332 57 333
rect 55 332 56 333
rect 54 332 55 333
rect 53 332 54 333
rect 52 332 53 333
rect 51 332 52 333
rect 39 332 40 333
rect 38 332 39 333
rect 37 332 38 333
rect 36 332 37 333
rect 35 332 36 333
rect 34 332 35 333
rect 33 332 34 333
rect 32 332 33 333
rect 31 332 32 333
rect 30 332 31 333
rect 29 332 30 333
rect 28 332 29 333
rect 27 332 28 333
rect 439 333 440 334
rect 438 333 439 334
rect 437 333 438 334
rect 397 333 398 334
rect 396 333 397 334
rect 395 333 396 334
rect 170 333 171 334
rect 169 333 170 334
rect 168 333 169 334
rect 167 333 168 334
rect 166 333 167 334
rect 165 333 166 334
rect 164 333 165 334
rect 163 333 164 334
rect 162 333 163 334
rect 161 333 162 334
rect 160 333 161 334
rect 159 333 160 334
rect 158 333 159 334
rect 157 333 158 334
rect 156 333 157 334
rect 155 333 156 334
rect 154 333 155 334
rect 153 333 154 334
rect 152 333 153 334
rect 151 333 152 334
rect 150 333 151 334
rect 149 333 150 334
rect 148 333 149 334
rect 147 333 148 334
rect 146 333 147 334
rect 145 333 146 334
rect 144 333 145 334
rect 143 333 144 334
rect 142 333 143 334
rect 141 333 142 334
rect 140 333 141 334
rect 139 333 140 334
rect 138 333 139 334
rect 137 333 138 334
rect 136 333 137 334
rect 135 333 136 334
rect 134 333 135 334
rect 133 333 134 334
rect 132 333 133 334
rect 131 333 132 334
rect 130 333 131 334
rect 129 333 130 334
rect 128 333 129 334
rect 127 333 128 334
rect 126 333 127 334
rect 125 333 126 334
rect 124 333 125 334
rect 123 333 124 334
rect 122 333 123 334
rect 121 333 122 334
rect 120 333 121 334
rect 119 333 120 334
rect 118 333 119 334
rect 117 333 118 334
rect 116 333 117 334
rect 115 333 116 334
rect 114 333 115 334
rect 113 333 114 334
rect 112 333 113 334
rect 111 333 112 334
rect 110 333 111 334
rect 109 333 110 334
rect 108 333 109 334
rect 107 333 108 334
rect 106 333 107 334
rect 86 333 87 334
rect 85 333 86 334
rect 84 333 85 334
rect 83 333 84 334
rect 82 333 83 334
rect 81 333 82 334
rect 80 333 81 334
rect 79 333 80 334
rect 78 333 79 334
rect 77 333 78 334
rect 76 333 77 334
rect 75 333 76 334
rect 74 333 75 334
rect 73 333 74 334
rect 72 333 73 334
rect 71 333 72 334
rect 70 333 71 334
rect 69 333 70 334
rect 68 333 69 334
rect 67 333 68 334
rect 66 333 67 334
rect 65 333 66 334
rect 64 333 65 334
rect 63 333 64 334
rect 62 333 63 334
rect 61 333 62 334
rect 60 333 61 334
rect 59 333 60 334
rect 58 333 59 334
rect 57 333 58 334
rect 56 333 57 334
rect 55 333 56 334
rect 54 333 55 334
rect 53 333 54 334
rect 52 333 53 334
rect 40 333 41 334
rect 39 333 40 334
rect 38 333 39 334
rect 37 333 38 334
rect 36 333 37 334
rect 35 333 36 334
rect 34 333 35 334
rect 33 333 34 334
rect 32 333 33 334
rect 31 333 32 334
rect 30 333 31 334
rect 29 333 30 334
rect 28 333 29 334
rect 439 334 440 335
rect 438 334 439 335
rect 437 334 438 335
rect 397 334 398 335
rect 396 334 397 335
rect 395 334 396 335
rect 174 334 175 335
rect 173 334 174 335
rect 172 334 173 335
rect 171 334 172 335
rect 170 334 171 335
rect 169 334 170 335
rect 168 334 169 335
rect 167 334 168 335
rect 166 334 167 335
rect 165 334 166 335
rect 164 334 165 335
rect 163 334 164 335
rect 162 334 163 335
rect 161 334 162 335
rect 160 334 161 335
rect 159 334 160 335
rect 158 334 159 335
rect 157 334 158 335
rect 156 334 157 335
rect 155 334 156 335
rect 154 334 155 335
rect 153 334 154 335
rect 152 334 153 335
rect 151 334 152 335
rect 150 334 151 335
rect 149 334 150 335
rect 148 334 149 335
rect 147 334 148 335
rect 146 334 147 335
rect 145 334 146 335
rect 144 334 145 335
rect 143 334 144 335
rect 142 334 143 335
rect 141 334 142 335
rect 140 334 141 335
rect 139 334 140 335
rect 138 334 139 335
rect 137 334 138 335
rect 136 334 137 335
rect 135 334 136 335
rect 134 334 135 335
rect 133 334 134 335
rect 132 334 133 335
rect 131 334 132 335
rect 130 334 131 335
rect 129 334 130 335
rect 128 334 129 335
rect 127 334 128 335
rect 126 334 127 335
rect 125 334 126 335
rect 124 334 125 335
rect 123 334 124 335
rect 122 334 123 335
rect 121 334 122 335
rect 120 334 121 335
rect 119 334 120 335
rect 118 334 119 335
rect 117 334 118 335
rect 116 334 117 335
rect 115 334 116 335
rect 114 334 115 335
rect 113 334 114 335
rect 112 334 113 335
rect 111 334 112 335
rect 110 334 111 335
rect 109 334 110 335
rect 108 334 109 335
rect 107 334 108 335
rect 87 334 88 335
rect 86 334 87 335
rect 85 334 86 335
rect 84 334 85 335
rect 83 334 84 335
rect 82 334 83 335
rect 81 334 82 335
rect 80 334 81 335
rect 79 334 80 335
rect 78 334 79 335
rect 77 334 78 335
rect 76 334 77 335
rect 75 334 76 335
rect 74 334 75 335
rect 73 334 74 335
rect 72 334 73 335
rect 71 334 72 335
rect 70 334 71 335
rect 69 334 70 335
rect 68 334 69 335
rect 67 334 68 335
rect 66 334 67 335
rect 65 334 66 335
rect 64 334 65 335
rect 63 334 64 335
rect 62 334 63 335
rect 61 334 62 335
rect 60 334 61 335
rect 59 334 60 335
rect 58 334 59 335
rect 57 334 58 335
rect 56 334 57 335
rect 55 334 56 335
rect 54 334 55 335
rect 53 334 54 335
rect 52 334 53 335
rect 40 334 41 335
rect 39 334 40 335
rect 38 334 39 335
rect 37 334 38 335
rect 36 334 37 335
rect 35 334 36 335
rect 34 334 35 335
rect 33 334 34 335
rect 32 334 33 335
rect 31 334 32 335
rect 30 334 31 335
rect 29 334 30 335
rect 439 335 440 336
rect 438 335 439 336
rect 437 335 438 336
rect 397 335 398 336
rect 396 335 397 336
rect 395 335 396 336
rect 178 335 179 336
rect 177 335 178 336
rect 176 335 177 336
rect 175 335 176 336
rect 174 335 175 336
rect 173 335 174 336
rect 172 335 173 336
rect 171 335 172 336
rect 170 335 171 336
rect 169 335 170 336
rect 168 335 169 336
rect 167 335 168 336
rect 166 335 167 336
rect 165 335 166 336
rect 164 335 165 336
rect 163 335 164 336
rect 162 335 163 336
rect 161 335 162 336
rect 160 335 161 336
rect 159 335 160 336
rect 158 335 159 336
rect 157 335 158 336
rect 156 335 157 336
rect 155 335 156 336
rect 154 335 155 336
rect 153 335 154 336
rect 152 335 153 336
rect 151 335 152 336
rect 150 335 151 336
rect 149 335 150 336
rect 148 335 149 336
rect 147 335 148 336
rect 146 335 147 336
rect 145 335 146 336
rect 144 335 145 336
rect 143 335 144 336
rect 142 335 143 336
rect 141 335 142 336
rect 140 335 141 336
rect 139 335 140 336
rect 138 335 139 336
rect 137 335 138 336
rect 136 335 137 336
rect 135 335 136 336
rect 134 335 135 336
rect 133 335 134 336
rect 132 335 133 336
rect 131 335 132 336
rect 130 335 131 336
rect 129 335 130 336
rect 128 335 129 336
rect 127 335 128 336
rect 126 335 127 336
rect 125 335 126 336
rect 124 335 125 336
rect 123 335 124 336
rect 122 335 123 336
rect 121 335 122 336
rect 120 335 121 336
rect 119 335 120 336
rect 118 335 119 336
rect 117 335 118 336
rect 116 335 117 336
rect 115 335 116 336
rect 114 335 115 336
rect 113 335 114 336
rect 112 335 113 336
rect 111 335 112 336
rect 110 335 111 336
rect 109 335 110 336
rect 108 335 109 336
rect 87 335 88 336
rect 86 335 87 336
rect 85 335 86 336
rect 84 335 85 336
rect 83 335 84 336
rect 82 335 83 336
rect 81 335 82 336
rect 80 335 81 336
rect 79 335 80 336
rect 78 335 79 336
rect 77 335 78 336
rect 76 335 77 336
rect 75 335 76 336
rect 74 335 75 336
rect 73 335 74 336
rect 72 335 73 336
rect 71 335 72 336
rect 70 335 71 336
rect 69 335 70 336
rect 68 335 69 336
rect 67 335 68 336
rect 66 335 67 336
rect 65 335 66 336
rect 64 335 65 336
rect 63 335 64 336
rect 62 335 63 336
rect 61 335 62 336
rect 60 335 61 336
rect 59 335 60 336
rect 58 335 59 336
rect 57 335 58 336
rect 56 335 57 336
rect 55 335 56 336
rect 54 335 55 336
rect 53 335 54 336
rect 40 335 41 336
rect 39 335 40 336
rect 38 335 39 336
rect 37 335 38 336
rect 36 335 37 336
rect 35 335 36 336
rect 34 335 35 336
rect 33 335 34 336
rect 32 335 33 336
rect 31 335 32 336
rect 30 335 31 336
rect 439 336 440 337
rect 438 336 439 337
rect 437 336 438 337
rect 436 336 437 337
rect 398 336 399 337
rect 397 336 398 337
rect 396 336 397 337
rect 395 336 396 337
rect 177 336 178 337
rect 176 336 177 337
rect 175 336 176 337
rect 174 336 175 337
rect 173 336 174 337
rect 172 336 173 337
rect 171 336 172 337
rect 170 336 171 337
rect 169 336 170 337
rect 168 336 169 337
rect 167 336 168 337
rect 166 336 167 337
rect 165 336 166 337
rect 164 336 165 337
rect 163 336 164 337
rect 162 336 163 337
rect 161 336 162 337
rect 160 336 161 337
rect 159 336 160 337
rect 158 336 159 337
rect 157 336 158 337
rect 156 336 157 337
rect 155 336 156 337
rect 154 336 155 337
rect 153 336 154 337
rect 152 336 153 337
rect 151 336 152 337
rect 150 336 151 337
rect 149 336 150 337
rect 148 336 149 337
rect 147 336 148 337
rect 146 336 147 337
rect 145 336 146 337
rect 144 336 145 337
rect 143 336 144 337
rect 142 336 143 337
rect 141 336 142 337
rect 140 336 141 337
rect 139 336 140 337
rect 138 336 139 337
rect 137 336 138 337
rect 136 336 137 337
rect 135 336 136 337
rect 134 336 135 337
rect 133 336 134 337
rect 132 336 133 337
rect 131 336 132 337
rect 130 336 131 337
rect 129 336 130 337
rect 128 336 129 337
rect 127 336 128 337
rect 126 336 127 337
rect 125 336 126 337
rect 124 336 125 337
rect 123 336 124 337
rect 122 336 123 337
rect 121 336 122 337
rect 120 336 121 337
rect 119 336 120 337
rect 118 336 119 337
rect 117 336 118 337
rect 116 336 117 337
rect 115 336 116 337
rect 114 336 115 337
rect 113 336 114 337
rect 112 336 113 337
rect 111 336 112 337
rect 110 336 111 337
rect 109 336 110 337
rect 88 336 89 337
rect 87 336 88 337
rect 86 336 87 337
rect 85 336 86 337
rect 84 336 85 337
rect 83 336 84 337
rect 82 336 83 337
rect 81 336 82 337
rect 80 336 81 337
rect 79 336 80 337
rect 78 336 79 337
rect 77 336 78 337
rect 76 336 77 337
rect 75 336 76 337
rect 74 336 75 337
rect 73 336 74 337
rect 72 336 73 337
rect 71 336 72 337
rect 70 336 71 337
rect 69 336 70 337
rect 68 336 69 337
rect 67 336 68 337
rect 66 336 67 337
rect 65 336 66 337
rect 64 336 65 337
rect 63 336 64 337
rect 62 336 63 337
rect 61 336 62 337
rect 60 336 61 337
rect 59 336 60 337
rect 58 336 59 337
rect 57 336 58 337
rect 56 336 57 337
rect 55 336 56 337
rect 54 336 55 337
rect 53 336 54 337
rect 41 336 42 337
rect 40 336 41 337
rect 39 336 40 337
rect 38 336 39 337
rect 37 336 38 337
rect 36 336 37 337
rect 35 336 36 337
rect 34 336 35 337
rect 33 336 34 337
rect 32 336 33 337
rect 31 336 32 337
rect 439 337 440 338
rect 438 337 439 338
rect 437 337 438 338
rect 436 337 437 338
rect 435 337 436 338
rect 434 337 435 338
rect 433 337 434 338
rect 432 337 433 338
rect 431 337 432 338
rect 430 337 431 338
rect 429 337 430 338
rect 428 337 429 338
rect 427 337 428 338
rect 426 337 427 338
rect 425 337 426 338
rect 424 337 425 338
rect 423 337 424 338
rect 422 337 423 338
rect 421 337 422 338
rect 420 337 421 338
rect 419 337 420 338
rect 418 337 419 338
rect 417 337 418 338
rect 416 337 417 338
rect 415 337 416 338
rect 414 337 415 338
rect 413 337 414 338
rect 412 337 413 338
rect 411 337 412 338
rect 410 337 411 338
rect 409 337 410 338
rect 408 337 409 338
rect 407 337 408 338
rect 406 337 407 338
rect 405 337 406 338
rect 404 337 405 338
rect 403 337 404 338
rect 402 337 403 338
rect 401 337 402 338
rect 400 337 401 338
rect 399 337 400 338
rect 398 337 399 338
rect 397 337 398 338
rect 396 337 397 338
rect 395 337 396 338
rect 176 337 177 338
rect 175 337 176 338
rect 174 337 175 338
rect 173 337 174 338
rect 172 337 173 338
rect 171 337 172 338
rect 170 337 171 338
rect 169 337 170 338
rect 168 337 169 338
rect 167 337 168 338
rect 166 337 167 338
rect 165 337 166 338
rect 164 337 165 338
rect 163 337 164 338
rect 162 337 163 338
rect 161 337 162 338
rect 160 337 161 338
rect 159 337 160 338
rect 158 337 159 338
rect 157 337 158 338
rect 156 337 157 338
rect 155 337 156 338
rect 154 337 155 338
rect 153 337 154 338
rect 152 337 153 338
rect 151 337 152 338
rect 150 337 151 338
rect 149 337 150 338
rect 148 337 149 338
rect 147 337 148 338
rect 146 337 147 338
rect 145 337 146 338
rect 144 337 145 338
rect 143 337 144 338
rect 142 337 143 338
rect 141 337 142 338
rect 140 337 141 338
rect 139 337 140 338
rect 138 337 139 338
rect 137 337 138 338
rect 136 337 137 338
rect 135 337 136 338
rect 134 337 135 338
rect 133 337 134 338
rect 132 337 133 338
rect 131 337 132 338
rect 130 337 131 338
rect 129 337 130 338
rect 128 337 129 338
rect 127 337 128 338
rect 126 337 127 338
rect 125 337 126 338
rect 124 337 125 338
rect 123 337 124 338
rect 122 337 123 338
rect 121 337 122 338
rect 120 337 121 338
rect 119 337 120 338
rect 118 337 119 338
rect 117 337 118 338
rect 116 337 117 338
rect 115 337 116 338
rect 114 337 115 338
rect 113 337 114 338
rect 112 337 113 338
rect 111 337 112 338
rect 110 337 111 338
rect 89 337 90 338
rect 88 337 89 338
rect 87 337 88 338
rect 86 337 87 338
rect 85 337 86 338
rect 84 337 85 338
rect 83 337 84 338
rect 82 337 83 338
rect 81 337 82 338
rect 80 337 81 338
rect 79 337 80 338
rect 78 337 79 338
rect 77 337 78 338
rect 76 337 77 338
rect 75 337 76 338
rect 74 337 75 338
rect 73 337 74 338
rect 72 337 73 338
rect 71 337 72 338
rect 70 337 71 338
rect 69 337 70 338
rect 68 337 69 338
rect 67 337 68 338
rect 66 337 67 338
rect 65 337 66 338
rect 64 337 65 338
rect 63 337 64 338
rect 62 337 63 338
rect 61 337 62 338
rect 60 337 61 338
rect 59 337 60 338
rect 58 337 59 338
rect 57 337 58 338
rect 56 337 57 338
rect 55 337 56 338
rect 54 337 55 338
rect 53 337 54 338
rect 41 337 42 338
rect 40 337 41 338
rect 39 337 40 338
rect 38 337 39 338
rect 37 337 38 338
rect 36 337 37 338
rect 35 337 36 338
rect 34 337 35 338
rect 33 337 34 338
rect 32 337 33 338
rect 439 338 440 339
rect 438 338 439 339
rect 437 338 438 339
rect 436 338 437 339
rect 435 338 436 339
rect 434 338 435 339
rect 433 338 434 339
rect 432 338 433 339
rect 431 338 432 339
rect 430 338 431 339
rect 429 338 430 339
rect 428 338 429 339
rect 427 338 428 339
rect 426 338 427 339
rect 425 338 426 339
rect 424 338 425 339
rect 423 338 424 339
rect 422 338 423 339
rect 421 338 422 339
rect 420 338 421 339
rect 419 338 420 339
rect 418 338 419 339
rect 417 338 418 339
rect 416 338 417 339
rect 415 338 416 339
rect 414 338 415 339
rect 413 338 414 339
rect 412 338 413 339
rect 411 338 412 339
rect 410 338 411 339
rect 409 338 410 339
rect 408 338 409 339
rect 407 338 408 339
rect 406 338 407 339
rect 405 338 406 339
rect 404 338 405 339
rect 403 338 404 339
rect 402 338 403 339
rect 401 338 402 339
rect 400 338 401 339
rect 399 338 400 339
rect 398 338 399 339
rect 397 338 398 339
rect 396 338 397 339
rect 395 338 396 339
rect 175 338 176 339
rect 174 338 175 339
rect 173 338 174 339
rect 172 338 173 339
rect 171 338 172 339
rect 170 338 171 339
rect 169 338 170 339
rect 168 338 169 339
rect 167 338 168 339
rect 166 338 167 339
rect 165 338 166 339
rect 164 338 165 339
rect 163 338 164 339
rect 162 338 163 339
rect 161 338 162 339
rect 160 338 161 339
rect 159 338 160 339
rect 158 338 159 339
rect 157 338 158 339
rect 156 338 157 339
rect 155 338 156 339
rect 154 338 155 339
rect 153 338 154 339
rect 152 338 153 339
rect 151 338 152 339
rect 150 338 151 339
rect 149 338 150 339
rect 148 338 149 339
rect 147 338 148 339
rect 146 338 147 339
rect 145 338 146 339
rect 144 338 145 339
rect 143 338 144 339
rect 142 338 143 339
rect 141 338 142 339
rect 140 338 141 339
rect 139 338 140 339
rect 138 338 139 339
rect 137 338 138 339
rect 136 338 137 339
rect 135 338 136 339
rect 134 338 135 339
rect 133 338 134 339
rect 132 338 133 339
rect 131 338 132 339
rect 130 338 131 339
rect 129 338 130 339
rect 128 338 129 339
rect 127 338 128 339
rect 126 338 127 339
rect 125 338 126 339
rect 124 338 125 339
rect 123 338 124 339
rect 122 338 123 339
rect 121 338 122 339
rect 120 338 121 339
rect 119 338 120 339
rect 118 338 119 339
rect 117 338 118 339
rect 116 338 117 339
rect 115 338 116 339
rect 114 338 115 339
rect 113 338 114 339
rect 112 338 113 339
rect 111 338 112 339
rect 90 338 91 339
rect 89 338 90 339
rect 88 338 89 339
rect 87 338 88 339
rect 86 338 87 339
rect 85 338 86 339
rect 84 338 85 339
rect 83 338 84 339
rect 82 338 83 339
rect 81 338 82 339
rect 80 338 81 339
rect 79 338 80 339
rect 78 338 79 339
rect 77 338 78 339
rect 76 338 77 339
rect 75 338 76 339
rect 74 338 75 339
rect 73 338 74 339
rect 72 338 73 339
rect 71 338 72 339
rect 70 338 71 339
rect 69 338 70 339
rect 68 338 69 339
rect 67 338 68 339
rect 66 338 67 339
rect 65 338 66 339
rect 64 338 65 339
rect 63 338 64 339
rect 62 338 63 339
rect 61 338 62 339
rect 60 338 61 339
rect 59 338 60 339
rect 58 338 59 339
rect 57 338 58 339
rect 56 338 57 339
rect 55 338 56 339
rect 54 338 55 339
rect 42 338 43 339
rect 41 338 42 339
rect 40 338 41 339
rect 39 338 40 339
rect 38 338 39 339
rect 37 338 38 339
rect 36 338 37 339
rect 35 338 36 339
rect 34 338 35 339
rect 33 338 34 339
rect 439 339 440 340
rect 438 339 439 340
rect 437 339 438 340
rect 436 339 437 340
rect 435 339 436 340
rect 434 339 435 340
rect 433 339 434 340
rect 432 339 433 340
rect 431 339 432 340
rect 430 339 431 340
rect 429 339 430 340
rect 428 339 429 340
rect 427 339 428 340
rect 426 339 427 340
rect 425 339 426 340
rect 424 339 425 340
rect 423 339 424 340
rect 422 339 423 340
rect 421 339 422 340
rect 420 339 421 340
rect 419 339 420 340
rect 418 339 419 340
rect 417 339 418 340
rect 416 339 417 340
rect 415 339 416 340
rect 414 339 415 340
rect 413 339 414 340
rect 412 339 413 340
rect 411 339 412 340
rect 410 339 411 340
rect 409 339 410 340
rect 408 339 409 340
rect 407 339 408 340
rect 406 339 407 340
rect 405 339 406 340
rect 404 339 405 340
rect 403 339 404 340
rect 402 339 403 340
rect 401 339 402 340
rect 400 339 401 340
rect 399 339 400 340
rect 398 339 399 340
rect 397 339 398 340
rect 396 339 397 340
rect 395 339 396 340
rect 174 339 175 340
rect 173 339 174 340
rect 172 339 173 340
rect 171 339 172 340
rect 170 339 171 340
rect 169 339 170 340
rect 168 339 169 340
rect 167 339 168 340
rect 166 339 167 340
rect 165 339 166 340
rect 164 339 165 340
rect 163 339 164 340
rect 162 339 163 340
rect 161 339 162 340
rect 160 339 161 340
rect 159 339 160 340
rect 158 339 159 340
rect 157 339 158 340
rect 156 339 157 340
rect 155 339 156 340
rect 154 339 155 340
rect 153 339 154 340
rect 152 339 153 340
rect 151 339 152 340
rect 150 339 151 340
rect 149 339 150 340
rect 148 339 149 340
rect 147 339 148 340
rect 146 339 147 340
rect 145 339 146 340
rect 144 339 145 340
rect 143 339 144 340
rect 142 339 143 340
rect 141 339 142 340
rect 140 339 141 340
rect 139 339 140 340
rect 138 339 139 340
rect 137 339 138 340
rect 136 339 137 340
rect 135 339 136 340
rect 134 339 135 340
rect 133 339 134 340
rect 132 339 133 340
rect 131 339 132 340
rect 130 339 131 340
rect 129 339 130 340
rect 128 339 129 340
rect 127 339 128 340
rect 126 339 127 340
rect 125 339 126 340
rect 124 339 125 340
rect 123 339 124 340
rect 122 339 123 340
rect 121 339 122 340
rect 120 339 121 340
rect 119 339 120 340
rect 118 339 119 340
rect 117 339 118 340
rect 116 339 117 340
rect 115 339 116 340
rect 114 339 115 340
rect 113 339 114 340
rect 112 339 113 340
rect 91 339 92 340
rect 90 339 91 340
rect 89 339 90 340
rect 88 339 89 340
rect 87 339 88 340
rect 86 339 87 340
rect 85 339 86 340
rect 84 339 85 340
rect 83 339 84 340
rect 82 339 83 340
rect 81 339 82 340
rect 80 339 81 340
rect 79 339 80 340
rect 78 339 79 340
rect 77 339 78 340
rect 76 339 77 340
rect 75 339 76 340
rect 74 339 75 340
rect 73 339 74 340
rect 72 339 73 340
rect 71 339 72 340
rect 70 339 71 340
rect 69 339 70 340
rect 68 339 69 340
rect 67 339 68 340
rect 66 339 67 340
rect 65 339 66 340
rect 64 339 65 340
rect 63 339 64 340
rect 62 339 63 340
rect 61 339 62 340
rect 60 339 61 340
rect 59 339 60 340
rect 58 339 59 340
rect 57 339 58 340
rect 56 339 57 340
rect 55 339 56 340
rect 54 339 55 340
rect 42 339 43 340
rect 41 339 42 340
rect 40 339 41 340
rect 39 339 40 340
rect 38 339 39 340
rect 37 339 38 340
rect 36 339 37 340
rect 35 339 36 340
rect 34 339 35 340
rect 439 340 440 341
rect 438 340 439 341
rect 437 340 438 341
rect 436 340 437 341
rect 435 340 436 341
rect 434 340 435 341
rect 433 340 434 341
rect 432 340 433 341
rect 431 340 432 341
rect 430 340 431 341
rect 429 340 430 341
rect 428 340 429 341
rect 427 340 428 341
rect 426 340 427 341
rect 425 340 426 341
rect 424 340 425 341
rect 423 340 424 341
rect 422 340 423 341
rect 421 340 422 341
rect 420 340 421 341
rect 419 340 420 341
rect 418 340 419 341
rect 417 340 418 341
rect 416 340 417 341
rect 415 340 416 341
rect 414 340 415 341
rect 413 340 414 341
rect 412 340 413 341
rect 411 340 412 341
rect 410 340 411 341
rect 409 340 410 341
rect 408 340 409 341
rect 407 340 408 341
rect 406 340 407 341
rect 405 340 406 341
rect 404 340 405 341
rect 403 340 404 341
rect 402 340 403 341
rect 401 340 402 341
rect 400 340 401 341
rect 399 340 400 341
rect 398 340 399 341
rect 397 340 398 341
rect 396 340 397 341
rect 395 340 396 341
rect 172 340 173 341
rect 171 340 172 341
rect 170 340 171 341
rect 169 340 170 341
rect 168 340 169 341
rect 167 340 168 341
rect 166 340 167 341
rect 165 340 166 341
rect 164 340 165 341
rect 163 340 164 341
rect 162 340 163 341
rect 161 340 162 341
rect 160 340 161 341
rect 159 340 160 341
rect 158 340 159 341
rect 157 340 158 341
rect 156 340 157 341
rect 155 340 156 341
rect 154 340 155 341
rect 153 340 154 341
rect 152 340 153 341
rect 151 340 152 341
rect 150 340 151 341
rect 149 340 150 341
rect 148 340 149 341
rect 147 340 148 341
rect 146 340 147 341
rect 145 340 146 341
rect 144 340 145 341
rect 143 340 144 341
rect 142 340 143 341
rect 141 340 142 341
rect 140 340 141 341
rect 139 340 140 341
rect 138 340 139 341
rect 137 340 138 341
rect 136 340 137 341
rect 135 340 136 341
rect 134 340 135 341
rect 133 340 134 341
rect 132 340 133 341
rect 131 340 132 341
rect 130 340 131 341
rect 129 340 130 341
rect 128 340 129 341
rect 127 340 128 341
rect 126 340 127 341
rect 125 340 126 341
rect 124 340 125 341
rect 123 340 124 341
rect 122 340 123 341
rect 121 340 122 341
rect 120 340 121 341
rect 119 340 120 341
rect 118 340 119 341
rect 117 340 118 341
rect 116 340 117 341
rect 115 340 116 341
rect 114 340 115 341
rect 113 340 114 341
rect 91 340 92 341
rect 90 340 91 341
rect 89 340 90 341
rect 88 340 89 341
rect 87 340 88 341
rect 86 340 87 341
rect 85 340 86 341
rect 84 340 85 341
rect 83 340 84 341
rect 82 340 83 341
rect 81 340 82 341
rect 80 340 81 341
rect 79 340 80 341
rect 78 340 79 341
rect 77 340 78 341
rect 76 340 77 341
rect 75 340 76 341
rect 74 340 75 341
rect 73 340 74 341
rect 72 340 73 341
rect 71 340 72 341
rect 70 340 71 341
rect 69 340 70 341
rect 68 340 69 341
rect 67 340 68 341
rect 66 340 67 341
rect 65 340 66 341
rect 64 340 65 341
rect 63 340 64 341
rect 62 340 63 341
rect 61 340 62 341
rect 60 340 61 341
rect 59 340 60 341
rect 58 340 59 341
rect 57 340 58 341
rect 56 340 57 341
rect 55 340 56 341
rect 43 340 44 341
rect 42 340 43 341
rect 41 340 42 341
rect 40 340 41 341
rect 39 340 40 341
rect 38 340 39 341
rect 37 340 38 341
rect 36 340 37 341
rect 35 340 36 341
rect 439 341 440 342
rect 438 341 439 342
rect 437 341 438 342
rect 436 341 437 342
rect 435 341 436 342
rect 434 341 435 342
rect 433 341 434 342
rect 432 341 433 342
rect 431 341 432 342
rect 430 341 431 342
rect 429 341 430 342
rect 428 341 429 342
rect 427 341 428 342
rect 426 341 427 342
rect 425 341 426 342
rect 424 341 425 342
rect 423 341 424 342
rect 422 341 423 342
rect 421 341 422 342
rect 420 341 421 342
rect 419 341 420 342
rect 418 341 419 342
rect 417 341 418 342
rect 416 341 417 342
rect 415 341 416 342
rect 414 341 415 342
rect 413 341 414 342
rect 412 341 413 342
rect 411 341 412 342
rect 410 341 411 342
rect 409 341 410 342
rect 408 341 409 342
rect 407 341 408 342
rect 406 341 407 342
rect 405 341 406 342
rect 404 341 405 342
rect 403 341 404 342
rect 402 341 403 342
rect 401 341 402 342
rect 400 341 401 342
rect 399 341 400 342
rect 398 341 399 342
rect 397 341 398 342
rect 396 341 397 342
rect 395 341 396 342
rect 170 341 171 342
rect 169 341 170 342
rect 168 341 169 342
rect 167 341 168 342
rect 166 341 167 342
rect 165 341 166 342
rect 164 341 165 342
rect 163 341 164 342
rect 162 341 163 342
rect 161 341 162 342
rect 160 341 161 342
rect 159 341 160 342
rect 158 341 159 342
rect 157 341 158 342
rect 156 341 157 342
rect 155 341 156 342
rect 154 341 155 342
rect 153 341 154 342
rect 152 341 153 342
rect 151 341 152 342
rect 150 341 151 342
rect 149 341 150 342
rect 148 341 149 342
rect 147 341 148 342
rect 146 341 147 342
rect 145 341 146 342
rect 144 341 145 342
rect 143 341 144 342
rect 142 341 143 342
rect 141 341 142 342
rect 140 341 141 342
rect 139 341 140 342
rect 138 341 139 342
rect 137 341 138 342
rect 136 341 137 342
rect 135 341 136 342
rect 134 341 135 342
rect 133 341 134 342
rect 132 341 133 342
rect 131 341 132 342
rect 130 341 131 342
rect 129 341 130 342
rect 128 341 129 342
rect 127 341 128 342
rect 126 341 127 342
rect 125 341 126 342
rect 124 341 125 342
rect 123 341 124 342
rect 122 341 123 342
rect 121 341 122 342
rect 120 341 121 342
rect 119 341 120 342
rect 118 341 119 342
rect 117 341 118 342
rect 116 341 117 342
rect 115 341 116 342
rect 114 341 115 342
rect 92 341 93 342
rect 91 341 92 342
rect 90 341 91 342
rect 89 341 90 342
rect 88 341 89 342
rect 87 341 88 342
rect 86 341 87 342
rect 85 341 86 342
rect 84 341 85 342
rect 83 341 84 342
rect 82 341 83 342
rect 81 341 82 342
rect 80 341 81 342
rect 79 341 80 342
rect 78 341 79 342
rect 77 341 78 342
rect 76 341 77 342
rect 75 341 76 342
rect 74 341 75 342
rect 73 341 74 342
rect 72 341 73 342
rect 71 341 72 342
rect 70 341 71 342
rect 69 341 70 342
rect 68 341 69 342
rect 67 341 68 342
rect 66 341 67 342
rect 65 341 66 342
rect 64 341 65 342
rect 63 341 64 342
rect 62 341 63 342
rect 61 341 62 342
rect 60 341 61 342
rect 59 341 60 342
rect 58 341 59 342
rect 57 341 58 342
rect 56 341 57 342
rect 55 341 56 342
rect 43 341 44 342
rect 42 341 43 342
rect 41 341 42 342
rect 40 341 41 342
rect 39 341 40 342
rect 38 341 39 342
rect 37 341 38 342
rect 439 342 440 343
rect 438 342 439 343
rect 437 342 438 343
rect 436 342 437 343
rect 435 342 436 343
rect 434 342 435 343
rect 433 342 434 343
rect 432 342 433 343
rect 431 342 432 343
rect 430 342 431 343
rect 429 342 430 343
rect 428 342 429 343
rect 427 342 428 343
rect 426 342 427 343
rect 425 342 426 343
rect 424 342 425 343
rect 423 342 424 343
rect 422 342 423 343
rect 421 342 422 343
rect 420 342 421 343
rect 419 342 420 343
rect 418 342 419 343
rect 417 342 418 343
rect 416 342 417 343
rect 415 342 416 343
rect 414 342 415 343
rect 413 342 414 343
rect 412 342 413 343
rect 411 342 412 343
rect 410 342 411 343
rect 409 342 410 343
rect 408 342 409 343
rect 407 342 408 343
rect 406 342 407 343
rect 405 342 406 343
rect 404 342 405 343
rect 403 342 404 343
rect 402 342 403 343
rect 401 342 402 343
rect 400 342 401 343
rect 399 342 400 343
rect 398 342 399 343
rect 397 342 398 343
rect 396 342 397 343
rect 395 342 396 343
rect 168 342 169 343
rect 167 342 168 343
rect 166 342 167 343
rect 165 342 166 343
rect 164 342 165 343
rect 163 342 164 343
rect 162 342 163 343
rect 161 342 162 343
rect 160 342 161 343
rect 159 342 160 343
rect 158 342 159 343
rect 157 342 158 343
rect 156 342 157 343
rect 155 342 156 343
rect 154 342 155 343
rect 153 342 154 343
rect 152 342 153 343
rect 151 342 152 343
rect 150 342 151 343
rect 149 342 150 343
rect 148 342 149 343
rect 147 342 148 343
rect 146 342 147 343
rect 145 342 146 343
rect 144 342 145 343
rect 143 342 144 343
rect 142 342 143 343
rect 141 342 142 343
rect 140 342 141 343
rect 139 342 140 343
rect 138 342 139 343
rect 137 342 138 343
rect 136 342 137 343
rect 135 342 136 343
rect 134 342 135 343
rect 133 342 134 343
rect 132 342 133 343
rect 131 342 132 343
rect 130 342 131 343
rect 129 342 130 343
rect 128 342 129 343
rect 127 342 128 343
rect 126 342 127 343
rect 125 342 126 343
rect 124 342 125 343
rect 123 342 124 343
rect 122 342 123 343
rect 121 342 122 343
rect 120 342 121 343
rect 119 342 120 343
rect 118 342 119 343
rect 117 342 118 343
rect 116 342 117 343
rect 115 342 116 343
rect 93 342 94 343
rect 92 342 93 343
rect 91 342 92 343
rect 90 342 91 343
rect 89 342 90 343
rect 88 342 89 343
rect 87 342 88 343
rect 86 342 87 343
rect 85 342 86 343
rect 84 342 85 343
rect 83 342 84 343
rect 82 342 83 343
rect 81 342 82 343
rect 80 342 81 343
rect 79 342 80 343
rect 78 342 79 343
rect 77 342 78 343
rect 76 342 77 343
rect 75 342 76 343
rect 74 342 75 343
rect 73 342 74 343
rect 72 342 73 343
rect 71 342 72 343
rect 70 342 71 343
rect 69 342 70 343
rect 68 342 69 343
rect 67 342 68 343
rect 66 342 67 343
rect 65 342 66 343
rect 64 342 65 343
rect 63 342 64 343
rect 62 342 63 343
rect 61 342 62 343
rect 60 342 61 343
rect 59 342 60 343
rect 58 342 59 343
rect 57 342 58 343
rect 56 342 57 343
rect 55 342 56 343
rect 44 342 45 343
rect 43 342 44 343
rect 42 342 43 343
rect 41 342 42 343
rect 40 342 41 343
rect 39 342 40 343
rect 38 342 39 343
rect 439 343 440 344
rect 438 343 439 344
rect 437 343 438 344
rect 436 343 437 344
rect 435 343 436 344
rect 434 343 435 344
rect 433 343 434 344
rect 432 343 433 344
rect 431 343 432 344
rect 430 343 431 344
rect 429 343 430 344
rect 428 343 429 344
rect 427 343 428 344
rect 426 343 427 344
rect 425 343 426 344
rect 424 343 425 344
rect 423 343 424 344
rect 422 343 423 344
rect 421 343 422 344
rect 420 343 421 344
rect 419 343 420 344
rect 418 343 419 344
rect 417 343 418 344
rect 416 343 417 344
rect 415 343 416 344
rect 414 343 415 344
rect 413 343 414 344
rect 412 343 413 344
rect 411 343 412 344
rect 410 343 411 344
rect 409 343 410 344
rect 408 343 409 344
rect 407 343 408 344
rect 406 343 407 344
rect 405 343 406 344
rect 404 343 405 344
rect 403 343 404 344
rect 402 343 403 344
rect 401 343 402 344
rect 400 343 401 344
rect 399 343 400 344
rect 398 343 399 344
rect 397 343 398 344
rect 396 343 397 344
rect 395 343 396 344
rect 166 343 167 344
rect 165 343 166 344
rect 164 343 165 344
rect 163 343 164 344
rect 162 343 163 344
rect 161 343 162 344
rect 160 343 161 344
rect 159 343 160 344
rect 158 343 159 344
rect 157 343 158 344
rect 156 343 157 344
rect 155 343 156 344
rect 154 343 155 344
rect 153 343 154 344
rect 152 343 153 344
rect 151 343 152 344
rect 150 343 151 344
rect 149 343 150 344
rect 148 343 149 344
rect 147 343 148 344
rect 146 343 147 344
rect 145 343 146 344
rect 144 343 145 344
rect 143 343 144 344
rect 142 343 143 344
rect 141 343 142 344
rect 140 343 141 344
rect 139 343 140 344
rect 138 343 139 344
rect 137 343 138 344
rect 136 343 137 344
rect 135 343 136 344
rect 134 343 135 344
rect 133 343 134 344
rect 132 343 133 344
rect 131 343 132 344
rect 130 343 131 344
rect 129 343 130 344
rect 128 343 129 344
rect 127 343 128 344
rect 126 343 127 344
rect 125 343 126 344
rect 124 343 125 344
rect 123 343 124 344
rect 122 343 123 344
rect 121 343 122 344
rect 120 343 121 344
rect 119 343 120 344
rect 118 343 119 344
rect 117 343 118 344
rect 94 343 95 344
rect 93 343 94 344
rect 92 343 93 344
rect 91 343 92 344
rect 90 343 91 344
rect 89 343 90 344
rect 88 343 89 344
rect 87 343 88 344
rect 86 343 87 344
rect 85 343 86 344
rect 84 343 85 344
rect 83 343 84 344
rect 82 343 83 344
rect 81 343 82 344
rect 80 343 81 344
rect 79 343 80 344
rect 78 343 79 344
rect 77 343 78 344
rect 76 343 77 344
rect 75 343 76 344
rect 74 343 75 344
rect 73 343 74 344
rect 72 343 73 344
rect 71 343 72 344
rect 70 343 71 344
rect 69 343 70 344
rect 68 343 69 344
rect 67 343 68 344
rect 66 343 67 344
rect 65 343 66 344
rect 64 343 65 344
rect 63 343 64 344
rect 62 343 63 344
rect 61 343 62 344
rect 60 343 61 344
rect 59 343 60 344
rect 58 343 59 344
rect 57 343 58 344
rect 56 343 57 344
rect 44 343 45 344
rect 43 343 44 344
rect 42 343 43 344
rect 41 343 42 344
rect 40 343 41 344
rect 439 344 440 345
rect 438 344 439 345
rect 437 344 438 345
rect 436 344 437 345
rect 435 344 436 345
rect 434 344 435 345
rect 433 344 434 345
rect 432 344 433 345
rect 431 344 432 345
rect 430 344 431 345
rect 429 344 430 345
rect 428 344 429 345
rect 427 344 428 345
rect 426 344 427 345
rect 425 344 426 345
rect 424 344 425 345
rect 423 344 424 345
rect 422 344 423 345
rect 421 344 422 345
rect 420 344 421 345
rect 419 344 420 345
rect 418 344 419 345
rect 417 344 418 345
rect 416 344 417 345
rect 415 344 416 345
rect 414 344 415 345
rect 413 344 414 345
rect 412 344 413 345
rect 411 344 412 345
rect 410 344 411 345
rect 409 344 410 345
rect 408 344 409 345
rect 407 344 408 345
rect 406 344 407 345
rect 405 344 406 345
rect 404 344 405 345
rect 403 344 404 345
rect 402 344 403 345
rect 401 344 402 345
rect 400 344 401 345
rect 399 344 400 345
rect 398 344 399 345
rect 397 344 398 345
rect 396 344 397 345
rect 395 344 396 345
rect 163 344 164 345
rect 162 344 163 345
rect 161 344 162 345
rect 160 344 161 345
rect 159 344 160 345
rect 158 344 159 345
rect 157 344 158 345
rect 156 344 157 345
rect 155 344 156 345
rect 154 344 155 345
rect 153 344 154 345
rect 152 344 153 345
rect 151 344 152 345
rect 150 344 151 345
rect 149 344 150 345
rect 148 344 149 345
rect 147 344 148 345
rect 146 344 147 345
rect 145 344 146 345
rect 144 344 145 345
rect 143 344 144 345
rect 142 344 143 345
rect 141 344 142 345
rect 140 344 141 345
rect 139 344 140 345
rect 138 344 139 345
rect 137 344 138 345
rect 136 344 137 345
rect 135 344 136 345
rect 134 344 135 345
rect 133 344 134 345
rect 132 344 133 345
rect 131 344 132 345
rect 130 344 131 345
rect 129 344 130 345
rect 128 344 129 345
rect 127 344 128 345
rect 126 344 127 345
rect 125 344 126 345
rect 124 344 125 345
rect 123 344 124 345
rect 122 344 123 345
rect 121 344 122 345
rect 120 344 121 345
rect 119 344 120 345
rect 118 344 119 345
rect 95 344 96 345
rect 94 344 95 345
rect 93 344 94 345
rect 92 344 93 345
rect 91 344 92 345
rect 90 344 91 345
rect 89 344 90 345
rect 88 344 89 345
rect 87 344 88 345
rect 86 344 87 345
rect 85 344 86 345
rect 84 344 85 345
rect 83 344 84 345
rect 82 344 83 345
rect 81 344 82 345
rect 80 344 81 345
rect 79 344 80 345
rect 78 344 79 345
rect 77 344 78 345
rect 76 344 77 345
rect 75 344 76 345
rect 74 344 75 345
rect 73 344 74 345
rect 72 344 73 345
rect 71 344 72 345
rect 70 344 71 345
rect 69 344 70 345
rect 68 344 69 345
rect 67 344 68 345
rect 66 344 67 345
rect 65 344 66 345
rect 64 344 65 345
rect 63 344 64 345
rect 62 344 63 345
rect 61 344 62 345
rect 60 344 61 345
rect 59 344 60 345
rect 58 344 59 345
rect 57 344 58 345
rect 56 344 57 345
rect 45 344 46 345
rect 44 344 45 345
rect 43 344 44 345
rect 439 345 440 346
rect 438 345 439 346
rect 437 345 438 346
rect 436 345 437 346
rect 435 345 436 346
rect 434 345 435 346
rect 433 345 434 346
rect 432 345 433 346
rect 431 345 432 346
rect 430 345 431 346
rect 429 345 430 346
rect 428 345 429 346
rect 427 345 428 346
rect 426 345 427 346
rect 425 345 426 346
rect 424 345 425 346
rect 423 345 424 346
rect 422 345 423 346
rect 421 345 422 346
rect 420 345 421 346
rect 419 345 420 346
rect 418 345 419 346
rect 417 345 418 346
rect 416 345 417 346
rect 415 345 416 346
rect 414 345 415 346
rect 413 345 414 346
rect 412 345 413 346
rect 411 345 412 346
rect 410 345 411 346
rect 409 345 410 346
rect 408 345 409 346
rect 407 345 408 346
rect 406 345 407 346
rect 405 345 406 346
rect 404 345 405 346
rect 403 345 404 346
rect 402 345 403 346
rect 401 345 402 346
rect 400 345 401 346
rect 399 345 400 346
rect 398 345 399 346
rect 397 345 398 346
rect 396 345 397 346
rect 395 345 396 346
rect 160 345 161 346
rect 159 345 160 346
rect 158 345 159 346
rect 157 345 158 346
rect 156 345 157 346
rect 155 345 156 346
rect 154 345 155 346
rect 153 345 154 346
rect 152 345 153 346
rect 151 345 152 346
rect 150 345 151 346
rect 149 345 150 346
rect 148 345 149 346
rect 147 345 148 346
rect 146 345 147 346
rect 145 345 146 346
rect 144 345 145 346
rect 143 345 144 346
rect 142 345 143 346
rect 141 345 142 346
rect 140 345 141 346
rect 139 345 140 346
rect 138 345 139 346
rect 137 345 138 346
rect 136 345 137 346
rect 135 345 136 346
rect 134 345 135 346
rect 133 345 134 346
rect 132 345 133 346
rect 131 345 132 346
rect 130 345 131 346
rect 129 345 130 346
rect 128 345 129 346
rect 127 345 128 346
rect 126 345 127 346
rect 125 345 126 346
rect 124 345 125 346
rect 123 345 124 346
rect 122 345 123 346
rect 121 345 122 346
rect 96 345 97 346
rect 95 345 96 346
rect 94 345 95 346
rect 93 345 94 346
rect 92 345 93 346
rect 91 345 92 346
rect 90 345 91 346
rect 89 345 90 346
rect 88 345 89 346
rect 87 345 88 346
rect 86 345 87 346
rect 85 345 86 346
rect 84 345 85 346
rect 83 345 84 346
rect 82 345 83 346
rect 81 345 82 346
rect 80 345 81 346
rect 79 345 80 346
rect 78 345 79 346
rect 77 345 78 346
rect 76 345 77 346
rect 75 345 76 346
rect 74 345 75 346
rect 73 345 74 346
rect 72 345 73 346
rect 71 345 72 346
rect 70 345 71 346
rect 69 345 70 346
rect 68 345 69 346
rect 67 345 68 346
rect 66 345 67 346
rect 65 345 66 346
rect 64 345 65 346
rect 63 345 64 346
rect 62 345 63 346
rect 61 345 62 346
rect 60 345 61 346
rect 59 345 60 346
rect 58 345 59 346
rect 57 345 58 346
rect 439 346 440 347
rect 438 346 439 347
rect 437 346 438 347
rect 436 346 437 347
rect 435 346 436 347
rect 434 346 435 347
rect 433 346 434 347
rect 432 346 433 347
rect 431 346 432 347
rect 430 346 431 347
rect 429 346 430 347
rect 428 346 429 347
rect 427 346 428 347
rect 426 346 427 347
rect 425 346 426 347
rect 424 346 425 347
rect 423 346 424 347
rect 422 346 423 347
rect 421 346 422 347
rect 420 346 421 347
rect 419 346 420 347
rect 418 346 419 347
rect 417 346 418 347
rect 416 346 417 347
rect 415 346 416 347
rect 414 346 415 347
rect 413 346 414 347
rect 412 346 413 347
rect 411 346 412 347
rect 410 346 411 347
rect 409 346 410 347
rect 408 346 409 347
rect 407 346 408 347
rect 406 346 407 347
rect 405 346 406 347
rect 404 346 405 347
rect 403 346 404 347
rect 402 346 403 347
rect 401 346 402 347
rect 400 346 401 347
rect 399 346 400 347
rect 398 346 399 347
rect 397 346 398 347
rect 396 346 397 347
rect 395 346 396 347
rect 156 346 157 347
rect 155 346 156 347
rect 154 346 155 347
rect 153 346 154 347
rect 152 346 153 347
rect 151 346 152 347
rect 150 346 151 347
rect 149 346 150 347
rect 148 346 149 347
rect 147 346 148 347
rect 146 346 147 347
rect 145 346 146 347
rect 144 346 145 347
rect 143 346 144 347
rect 142 346 143 347
rect 141 346 142 347
rect 140 346 141 347
rect 139 346 140 347
rect 138 346 139 347
rect 137 346 138 347
rect 136 346 137 347
rect 135 346 136 347
rect 134 346 135 347
rect 133 346 134 347
rect 132 346 133 347
rect 131 346 132 347
rect 130 346 131 347
rect 129 346 130 347
rect 128 346 129 347
rect 127 346 128 347
rect 126 346 127 347
rect 125 346 126 347
rect 124 346 125 347
rect 97 346 98 347
rect 96 346 97 347
rect 95 346 96 347
rect 94 346 95 347
rect 93 346 94 347
rect 92 346 93 347
rect 91 346 92 347
rect 90 346 91 347
rect 89 346 90 347
rect 88 346 89 347
rect 87 346 88 347
rect 86 346 87 347
rect 85 346 86 347
rect 84 346 85 347
rect 83 346 84 347
rect 82 346 83 347
rect 81 346 82 347
rect 80 346 81 347
rect 79 346 80 347
rect 78 346 79 347
rect 77 346 78 347
rect 76 346 77 347
rect 75 346 76 347
rect 74 346 75 347
rect 73 346 74 347
rect 72 346 73 347
rect 71 346 72 347
rect 70 346 71 347
rect 69 346 70 347
rect 68 346 69 347
rect 67 346 68 347
rect 66 346 67 347
rect 65 346 66 347
rect 64 346 65 347
rect 63 346 64 347
rect 62 346 63 347
rect 61 346 62 347
rect 60 346 61 347
rect 59 346 60 347
rect 58 346 59 347
rect 57 346 58 347
rect 439 347 440 348
rect 438 347 439 348
rect 437 347 438 348
rect 436 347 437 348
rect 418 347 419 348
rect 417 347 418 348
rect 416 347 417 348
rect 415 347 416 348
rect 397 347 398 348
rect 396 347 397 348
rect 395 347 396 348
rect 150 347 151 348
rect 149 347 150 348
rect 148 347 149 348
rect 147 347 148 348
rect 146 347 147 348
rect 145 347 146 348
rect 144 347 145 348
rect 143 347 144 348
rect 142 347 143 348
rect 141 347 142 348
rect 140 347 141 348
rect 139 347 140 348
rect 138 347 139 348
rect 137 347 138 348
rect 136 347 137 348
rect 135 347 136 348
rect 134 347 135 348
rect 133 347 134 348
rect 132 347 133 348
rect 131 347 132 348
rect 130 347 131 348
rect 129 347 130 348
rect 98 347 99 348
rect 97 347 98 348
rect 96 347 97 348
rect 95 347 96 348
rect 94 347 95 348
rect 93 347 94 348
rect 92 347 93 348
rect 91 347 92 348
rect 90 347 91 348
rect 89 347 90 348
rect 88 347 89 348
rect 87 347 88 348
rect 86 347 87 348
rect 85 347 86 348
rect 84 347 85 348
rect 83 347 84 348
rect 82 347 83 348
rect 81 347 82 348
rect 80 347 81 348
rect 79 347 80 348
rect 78 347 79 348
rect 77 347 78 348
rect 76 347 77 348
rect 75 347 76 348
rect 74 347 75 348
rect 73 347 74 348
rect 72 347 73 348
rect 71 347 72 348
rect 70 347 71 348
rect 69 347 70 348
rect 68 347 69 348
rect 67 347 68 348
rect 66 347 67 348
rect 65 347 66 348
rect 64 347 65 348
rect 63 347 64 348
rect 62 347 63 348
rect 61 347 62 348
rect 60 347 61 348
rect 59 347 60 348
rect 58 347 59 348
rect 439 348 440 349
rect 438 348 439 349
rect 437 348 438 349
rect 436 348 437 349
rect 418 348 419 349
rect 417 348 418 349
rect 416 348 417 349
rect 415 348 416 349
rect 397 348 398 349
rect 396 348 397 349
rect 395 348 396 349
rect 99 348 100 349
rect 98 348 99 349
rect 97 348 98 349
rect 96 348 97 349
rect 95 348 96 349
rect 94 348 95 349
rect 93 348 94 349
rect 92 348 93 349
rect 91 348 92 349
rect 90 348 91 349
rect 89 348 90 349
rect 88 348 89 349
rect 87 348 88 349
rect 86 348 87 349
rect 85 348 86 349
rect 84 348 85 349
rect 83 348 84 349
rect 82 348 83 349
rect 81 348 82 349
rect 80 348 81 349
rect 79 348 80 349
rect 78 348 79 349
rect 77 348 78 349
rect 76 348 77 349
rect 75 348 76 349
rect 74 348 75 349
rect 73 348 74 349
rect 72 348 73 349
rect 71 348 72 349
rect 70 348 71 349
rect 69 348 70 349
rect 68 348 69 349
rect 67 348 68 349
rect 66 348 67 349
rect 65 348 66 349
rect 64 348 65 349
rect 63 348 64 349
rect 62 348 63 349
rect 61 348 62 349
rect 60 348 61 349
rect 59 348 60 349
rect 58 348 59 349
rect 439 349 440 350
rect 438 349 439 350
rect 437 349 438 350
rect 418 349 419 350
rect 417 349 418 350
rect 416 349 417 350
rect 415 349 416 350
rect 397 349 398 350
rect 396 349 397 350
rect 395 349 396 350
rect 100 349 101 350
rect 99 349 100 350
rect 98 349 99 350
rect 97 349 98 350
rect 96 349 97 350
rect 95 349 96 350
rect 94 349 95 350
rect 93 349 94 350
rect 92 349 93 350
rect 91 349 92 350
rect 90 349 91 350
rect 89 349 90 350
rect 88 349 89 350
rect 87 349 88 350
rect 86 349 87 350
rect 85 349 86 350
rect 84 349 85 350
rect 83 349 84 350
rect 82 349 83 350
rect 81 349 82 350
rect 80 349 81 350
rect 79 349 80 350
rect 78 349 79 350
rect 77 349 78 350
rect 76 349 77 350
rect 75 349 76 350
rect 74 349 75 350
rect 73 349 74 350
rect 72 349 73 350
rect 71 349 72 350
rect 70 349 71 350
rect 69 349 70 350
rect 68 349 69 350
rect 67 349 68 350
rect 66 349 67 350
rect 65 349 66 350
rect 64 349 65 350
rect 63 349 64 350
rect 62 349 63 350
rect 61 349 62 350
rect 60 349 61 350
rect 59 349 60 350
rect 58 349 59 350
rect 439 350 440 351
rect 438 350 439 351
rect 437 350 438 351
rect 418 350 419 351
rect 417 350 418 351
rect 416 350 417 351
rect 415 350 416 351
rect 397 350 398 351
rect 396 350 397 351
rect 395 350 396 351
rect 101 350 102 351
rect 100 350 101 351
rect 99 350 100 351
rect 98 350 99 351
rect 97 350 98 351
rect 96 350 97 351
rect 95 350 96 351
rect 94 350 95 351
rect 93 350 94 351
rect 92 350 93 351
rect 91 350 92 351
rect 90 350 91 351
rect 89 350 90 351
rect 88 350 89 351
rect 87 350 88 351
rect 86 350 87 351
rect 85 350 86 351
rect 84 350 85 351
rect 83 350 84 351
rect 82 350 83 351
rect 81 350 82 351
rect 80 350 81 351
rect 79 350 80 351
rect 78 350 79 351
rect 77 350 78 351
rect 76 350 77 351
rect 75 350 76 351
rect 74 350 75 351
rect 73 350 74 351
rect 72 350 73 351
rect 71 350 72 351
rect 70 350 71 351
rect 69 350 70 351
rect 68 350 69 351
rect 67 350 68 351
rect 66 350 67 351
rect 65 350 66 351
rect 64 350 65 351
rect 63 350 64 351
rect 62 350 63 351
rect 61 350 62 351
rect 60 350 61 351
rect 59 350 60 351
rect 439 351 440 352
rect 438 351 439 352
rect 437 351 438 352
rect 418 351 419 352
rect 417 351 418 352
rect 416 351 417 352
rect 415 351 416 352
rect 397 351 398 352
rect 396 351 397 352
rect 395 351 396 352
rect 103 351 104 352
rect 102 351 103 352
rect 101 351 102 352
rect 100 351 101 352
rect 99 351 100 352
rect 98 351 99 352
rect 97 351 98 352
rect 96 351 97 352
rect 95 351 96 352
rect 94 351 95 352
rect 93 351 94 352
rect 92 351 93 352
rect 91 351 92 352
rect 90 351 91 352
rect 89 351 90 352
rect 88 351 89 352
rect 87 351 88 352
rect 86 351 87 352
rect 85 351 86 352
rect 84 351 85 352
rect 83 351 84 352
rect 82 351 83 352
rect 81 351 82 352
rect 80 351 81 352
rect 79 351 80 352
rect 78 351 79 352
rect 77 351 78 352
rect 76 351 77 352
rect 75 351 76 352
rect 74 351 75 352
rect 73 351 74 352
rect 72 351 73 352
rect 71 351 72 352
rect 70 351 71 352
rect 69 351 70 352
rect 68 351 69 352
rect 67 351 68 352
rect 66 351 67 352
rect 65 351 66 352
rect 64 351 65 352
rect 63 351 64 352
rect 62 351 63 352
rect 61 351 62 352
rect 60 351 61 352
rect 439 352 440 353
rect 438 352 439 353
rect 437 352 438 353
rect 418 352 419 353
rect 417 352 418 353
rect 416 352 417 353
rect 415 352 416 353
rect 397 352 398 353
rect 396 352 397 353
rect 395 352 396 353
rect 104 352 105 353
rect 103 352 104 353
rect 102 352 103 353
rect 101 352 102 353
rect 100 352 101 353
rect 99 352 100 353
rect 98 352 99 353
rect 97 352 98 353
rect 96 352 97 353
rect 95 352 96 353
rect 94 352 95 353
rect 93 352 94 353
rect 92 352 93 353
rect 91 352 92 353
rect 90 352 91 353
rect 89 352 90 353
rect 88 352 89 353
rect 87 352 88 353
rect 86 352 87 353
rect 85 352 86 353
rect 84 352 85 353
rect 83 352 84 353
rect 82 352 83 353
rect 81 352 82 353
rect 80 352 81 353
rect 79 352 80 353
rect 78 352 79 353
rect 77 352 78 353
rect 76 352 77 353
rect 75 352 76 353
rect 74 352 75 353
rect 73 352 74 353
rect 72 352 73 353
rect 71 352 72 353
rect 70 352 71 353
rect 69 352 70 353
rect 68 352 69 353
rect 67 352 68 353
rect 66 352 67 353
rect 65 352 66 353
rect 64 352 65 353
rect 63 352 64 353
rect 62 352 63 353
rect 61 352 62 353
rect 439 353 440 354
rect 438 353 439 354
rect 437 353 438 354
rect 418 353 419 354
rect 417 353 418 354
rect 416 353 417 354
rect 415 353 416 354
rect 397 353 398 354
rect 396 353 397 354
rect 395 353 396 354
rect 105 353 106 354
rect 104 353 105 354
rect 103 353 104 354
rect 102 353 103 354
rect 101 353 102 354
rect 100 353 101 354
rect 99 353 100 354
rect 98 353 99 354
rect 97 353 98 354
rect 96 353 97 354
rect 95 353 96 354
rect 94 353 95 354
rect 93 353 94 354
rect 92 353 93 354
rect 91 353 92 354
rect 90 353 91 354
rect 89 353 90 354
rect 88 353 89 354
rect 87 353 88 354
rect 86 353 87 354
rect 85 353 86 354
rect 84 353 85 354
rect 83 353 84 354
rect 82 353 83 354
rect 81 353 82 354
rect 80 353 81 354
rect 79 353 80 354
rect 78 353 79 354
rect 77 353 78 354
rect 76 353 77 354
rect 75 353 76 354
rect 74 353 75 354
rect 73 353 74 354
rect 72 353 73 354
rect 71 353 72 354
rect 70 353 71 354
rect 69 353 70 354
rect 68 353 69 354
rect 67 353 68 354
rect 66 353 67 354
rect 65 353 66 354
rect 64 353 65 354
rect 63 353 64 354
rect 62 353 63 354
rect 61 353 62 354
rect 439 354 440 355
rect 438 354 439 355
rect 437 354 438 355
rect 418 354 419 355
rect 417 354 418 355
rect 416 354 417 355
rect 415 354 416 355
rect 397 354 398 355
rect 396 354 397 355
rect 395 354 396 355
rect 107 354 108 355
rect 106 354 107 355
rect 105 354 106 355
rect 104 354 105 355
rect 103 354 104 355
rect 102 354 103 355
rect 101 354 102 355
rect 100 354 101 355
rect 99 354 100 355
rect 98 354 99 355
rect 97 354 98 355
rect 96 354 97 355
rect 95 354 96 355
rect 94 354 95 355
rect 93 354 94 355
rect 92 354 93 355
rect 91 354 92 355
rect 90 354 91 355
rect 89 354 90 355
rect 88 354 89 355
rect 87 354 88 355
rect 86 354 87 355
rect 85 354 86 355
rect 84 354 85 355
rect 83 354 84 355
rect 82 354 83 355
rect 81 354 82 355
rect 80 354 81 355
rect 79 354 80 355
rect 78 354 79 355
rect 77 354 78 355
rect 76 354 77 355
rect 75 354 76 355
rect 74 354 75 355
rect 73 354 74 355
rect 72 354 73 355
rect 71 354 72 355
rect 70 354 71 355
rect 69 354 70 355
rect 68 354 69 355
rect 67 354 68 355
rect 66 354 67 355
rect 65 354 66 355
rect 64 354 65 355
rect 63 354 64 355
rect 439 355 440 356
rect 438 355 439 356
rect 437 355 438 356
rect 418 355 419 356
rect 417 355 418 356
rect 416 355 417 356
rect 415 355 416 356
rect 397 355 398 356
rect 396 355 397 356
rect 395 355 396 356
rect 108 355 109 356
rect 107 355 108 356
rect 106 355 107 356
rect 105 355 106 356
rect 104 355 105 356
rect 103 355 104 356
rect 102 355 103 356
rect 101 355 102 356
rect 100 355 101 356
rect 99 355 100 356
rect 98 355 99 356
rect 97 355 98 356
rect 96 355 97 356
rect 95 355 96 356
rect 94 355 95 356
rect 93 355 94 356
rect 92 355 93 356
rect 91 355 92 356
rect 90 355 91 356
rect 89 355 90 356
rect 88 355 89 356
rect 87 355 88 356
rect 86 355 87 356
rect 85 355 86 356
rect 84 355 85 356
rect 83 355 84 356
rect 82 355 83 356
rect 81 355 82 356
rect 80 355 81 356
rect 79 355 80 356
rect 78 355 79 356
rect 77 355 78 356
rect 76 355 77 356
rect 75 355 76 356
rect 74 355 75 356
rect 73 355 74 356
rect 72 355 73 356
rect 71 355 72 356
rect 70 355 71 356
rect 69 355 70 356
rect 68 355 69 356
rect 67 355 68 356
rect 66 355 67 356
rect 65 355 66 356
rect 64 355 65 356
rect 439 356 440 357
rect 438 356 439 357
rect 437 356 438 357
rect 418 356 419 357
rect 417 356 418 357
rect 416 356 417 357
rect 415 356 416 357
rect 398 356 399 357
rect 397 356 398 357
rect 396 356 397 357
rect 395 356 396 357
rect 110 356 111 357
rect 109 356 110 357
rect 108 356 109 357
rect 107 356 108 357
rect 106 356 107 357
rect 105 356 106 357
rect 104 356 105 357
rect 103 356 104 357
rect 102 356 103 357
rect 101 356 102 357
rect 100 356 101 357
rect 99 356 100 357
rect 98 356 99 357
rect 97 356 98 357
rect 96 356 97 357
rect 95 356 96 357
rect 94 356 95 357
rect 93 356 94 357
rect 92 356 93 357
rect 91 356 92 357
rect 90 356 91 357
rect 89 356 90 357
rect 88 356 89 357
rect 87 356 88 357
rect 86 356 87 357
rect 85 356 86 357
rect 84 356 85 357
rect 83 356 84 357
rect 82 356 83 357
rect 81 356 82 357
rect 80 356 81 357
rect 79 356 80 357
rect 78 356 79 357
rect 77 356 78 357
rect 76 356 77 357
rect 75 356 76 357
rect 74 356 75 357
rect 73 356 74 357
rect 72 356 73 357
rect 71 356 72 357
rect 70 356 71 357
rect 69 356 70 357
rect 68 356 69 357
rect 67 356 68 357
rect 66 356 67 357
rect 65 356 66 357
rect 439 357 440 358
rect 438 357 439 358
rect 437 357 438 358
rect 419 357 420 358
rect 418 357 419 358
rect 417 357 418 358
rect 416 357 417 358
rect 415 357 416 358
rect 414 357 415 358
rect 398 357 399 358
rect 397 357 398 358
rect 396 357 397 358
rect 395 357 396 358
rect 111 357 112 358
rect 110 357 111 358
rect 109 357 110 358
rect 108 357 109 358
rect 107 357 108 358
rect 106 357 107 358
rect 105 357 106 358
rect 104 357 105 358
rect 103 357 104 358
rect 102 357 103 358
rect 101 357 102 358
rect 100 357 101 358
rect 99 357 100 358
rect 98 357 99 358
rect 97 357 98 358
rect 96 357 97 358
rect 95 357 96 358
rect 94 357 95 358
rect 93 357 94 358
rect 92 357 93 358
rect 91 357 92 358
rect 90 357 91 358
rect 89 357 90 358
rect 88 357 89 358
rect 87 357 88 358
rect 86 357 87 358
rect 85 357 86 358
rect 84 357 85 358
rect 83 357 84 358
rect 82 357 83 358
rect 81 357 82 358
rect 80 357 81 358
rect 79 357 80 358
rect 78 357 79 358
rect 77 357 78 358
rect 76 357 77 358
rect 75 357 76 358
rect 74 357 75 358
rect 73 357 74 358
rect 72 357 73 358
rect 71 357 72 358
rect 70 357 71 358
rect 69 357 70 358
rect 68 357 69 358
rect 67 357 68 358
rect 439 358 440 359
rect 438 358 439 359
rect 437 358 438 359
rect 422 358 423 359
rect 421 358 422 359
rect 420 358 421 359
rect 419 358 420 359
rect 418 358 419 359
rect 417 358 418 359
rect 416 358 417 359
rect 415 358 416 359
rect 414 358 415 359
rect 413 358 414 359
rect 412 358 413 359
rect 411 358 412 359
rect 398 358 399 359
rect 397 358 398 359
rect 396 358 397 359
rect 395 358 396 359
rect 113 358 114 359
rect 112 358 113 359
rect 111 358 112 359
rect 110 358 111 359
rect 109 358 110 359
rect 108 358 109 359
rect 107 358 108 359
rect 106 358 107 359
rect 105 358 106 359
rect 104 358 105 359
rect 103 358 104 359
rect 102 358 103 359
rect 101 358 102 359
rect 100 358 101 359
rect 99 358 100 359
rect 98 358 99 359
rect 97 358 98 359
rect 96 358 97 359
rect 95 358 96 359
rect 94 358 95 359
rect 93 358 94 359
rect 92 358 93 359
rect 91 358 92 359
rect 90 358 91 359
rect 89 358 90 359
rect 88 358 89 359
rect 87 358 88 359
rect 86 358 87 359
rect 85 358 86 359
rect 84 358 85 359
rect 83 358 84 359
rect 82 358 83 359
rect 81 358 82 359
rect 80 358 81 359
rect 79 358 80 359
rect 78 358 79 359
rect 77 358 78 359
rect 76 358 77 359
rect 75 358 76 359
rect 74 358 75 359
rect 73 358 74 359
rect 72 358 73 359
rect 71 358 72 359
rect 70 358 71 359
rect 69 358 70 359
rect 439 359 440 360
rect 438 359 439 360
rect 437 359 438 360
rect 436 359 437 360
rect 423 359 424 360
rect 422 359 423 360
rect 421 359 422 360
rect 420 359 421 360
rect 419 359 420 360
rect 418 359 419 360
rect 417 359 418 360
rect 416 359 417 360
rect 415 359 416 360
rect 414 359 415 360
rect 413 359 414 360
rect 412 359 413 360
rect 411 359 412 360
rect 410 359 411 360
rect 399 359 400 360
rect 398 359 399 360
rect 397 359 398 360
rect 396 359 397 360
rect 395 359 396 360
rect 115 359 116 360
rect 114 359 115 360
rect 113 359 114 360
rect 112 359 113 360
rect 111 359 112 360
rect 110 359 111 360
rect 109 359 110 360
rect 108 359 109 360
rect 107 359 108 360
rect 106 359 107 360
rect 105 359 106 360
rect 104 359 105 360
rect 103 359 104 360
rect 102 359 103 360
rect 101 359 102 360
rect 100 359 101 360
rect 99 359 100 360
rect 98 359 99 360
rect 97 359 98 360
rect 96 359 97 360
rect 95 359 96 360
rect 94 359 95 360
rect 93 359 94 360
rect 92 359 93 360
rect 91 359 92 360
rect 90 359 91 360
rect 89 359 90 360
rect 88 359 89 360
rect 87 359 88 360
rect 86 359 87 360
rect 85 359 86 360
rect 84 359 85 360
rect 83 359 84 360
rect 82 359 83 360
rect 81 359 82 360
rect 80 359 81 360
rect 79 359 80 360
rect 78 359 79 360
rect 77 359 78 360
rect 76 359 77 360
rect 75 359 76 360
rect 74 359 75 360
rect 73 359 74 360
rect 72 359 73 360
rect 71 359 72 360
rect 439 360 440 361
rect 438 360 439 361
rect 437 360 438 361
rect 436 360 437 361
rect 423 360 424 361
rect 422 360 423 361
rect 421 360 422 361
rect 420 360 421 361
rect 419 360 420 361
rect 418 360 419 361
rect 417 360 418 361
rect 416 360 417 361
rect 415 360 416 361
rect 414 360 415 361
rect 413 360 414 361
rect 412 360 413 361
rect 411 360 412 361
rect 410 360 411 361
rect 400 360 401 361
rect 399 360 400 361
rect 398 360 399 361
rect 397 360 398 361
rect 396 360 397 361
rect 395 360 396 361
rect 117 360 118 361
rect 116 360 117 361
rect 115 360 116 361
rect 114 360 115 361
rect 113 360 114 361
rect 112 360 113 361
rect 111 360 112 361
rect 110 360 111 361
rect 109 360 110 361
rect 108 360 109 361
rect 107 360 108 361
rect 106 360 107 361
rect 105 360 106 361
rect 104 360 105 361
rect 103 360 104 361
rect 102 360 103 361
rect 101 360 102 361
rect 100 360 101 361
rect 99 360 100 361
rect 98 360 99 361
rect 97 360 98 361
rect 96 360 97 361
rect 95 360 96 361
rect 94 360 95 361
rect 93 360 94 361
rect 92 360 93 361
rect 91 360 92 361
rect 90 360 91 361
rect 89 360 90 361
rect 88 360 89 361
rect 87 360 88 361
rect 86 360 87 361
rect 85 360 86 361
rect 84 360 85 361
rect 83 360 84 361
rect 82 360 83 361
rect 81 360 82 361
rect 80 360 81 361
rect 79 360 80 361
rect 78 360 79 361
rect 77 360 78 361
rect 76 360 77 361
rect 75 360 76 361
rect 74 360 75 361
rect 73 360 74 361
rect 439 361 440 362
rect 438 361 439 362
rect 437 361 438 362
rect 436 361 437 362
rect 435 361 436 362
rect 402 361 403 362
rect 401 361 402 362
rect 400 361 401 362
rect 399 361 400 362
rect 398 361 399 362
rect 397 361 398 362
rect 396 361 397 362
rect 395 361 396 362
rect 116 361 117 362
rect 115 361 116 362
rect 114 361 115 362
rect 113 361 114 362
rect 112 361 113 362
rect 111 361 112 362
rect 110 361 111 362
rect 109 361 110 362
rect 108 361 109 362
rect 107 361 108 362
rect 106 361 107 362
rect 105 361 106 362
rect 104 361 105 362
rect 103 361 104 362
rect 102 361 103 362
rect 101 361 102 362
rect 100 361 101 362
rect 99 361 100 362
rect 98 361 99 362
rect 97 361 98 362
rect 96 361 97 362
rect 95 361 96 362
rect 94 361 95 362
rect 93 361 94 362
rect 92 361 93 362
rect 91 361 92 362
rect 90 361 91 362
rect 89 361 90 362
rect 88 361 89 362
rect 87 361 88 362
rect 86 361 87 362
rect 85 361 86 362
rect 84 361 85 362
rect 83 361 84 362
rect 82 361 83 362
rect 81 361 82 362
rect 80 361 81 362
rect 79 361 80 362
rect 78 361 79 362
rect 77 361 78 362
rect 76 361 77 362
rect 439 362 440 363
rect 438 362 439 363
rect 437 362 438 363
rect 436 362 437 363
rect 435 362 436 363
rect 434 362 435 363
rect 405 362 406 363
rect 404 362 405 363
rect 403 362 404 363
rect 402 362 403 363
rect 401 362 402 363
rect 400 362 401 363
rect 399 362 400 363
rect 398 362 399 363
rect 397 362 398 363
rect 396 362 397 363
rect 395 362 396 363
rect 114 362 115 363
rect 113 362 114 363
rect 112 362 113 363
rect 111 362 112 363
rect 110 362 111 363
rect 109 362 110 363
rect 108 362 109 363
rect 107 362 108 363
rect 106 362 107 363
rect 105 362 106 363
rect 104 362 105 363
rect 103 362 104 363
rect 102 362 103 363
rect 101 362 102 363
rect 100 362 101 363
rect 99 362 100 363
rect 98 362 99 363
rect 97 362 98 363
rect 96 362 97 363
rect 95 362 96 363
rect 94 362 95 363
rect 93 362 94 363
rect 92 362 93 363
rect 91 362 92 363
rect 90 362 91 363
rect 89 362 90 363
rect 88 362 89 363
rect 87 362 88 363
rect 86 362 87 363
rect 85 362 86 363
rect 84 362 85 363
rect 83 362 84 363
rect 82 362 83 363
rect 81 362 82 363
rect 80 362 81 363
rect 439 363 440 364
rect 438 363 439 364
rect 437 363 438 364
rect 436 363 437 364
rect 435 363 436 364
rect 434 363 435 364
rect 433 363 434 364
rect 405 363 406 364
rect 404 363 405 364
rect 403 363 404 364
rect 402 363 403 364
rect 401 363 402 364
rect 400 363 401 364
rect 399 363 400 364
rect 398 363 399 364
rect 397 363 398 364
rect 396 363 397 364
rect 395 363 396 364
rect 111 363 112 364
rect 110 363 111 364
rect 109 363 110 364
rect 108 363 109 364
rect 107 363 108 364
rect 106 363 107 364
rect 105 363 106 364
rect 104 363 105 364
rect 103 363 104 364
rect 102 363 103 364
rect 101 363 102 364
rect 100 363 101 364
rect 99 363 100 364
rect 98 363 99 364
rect 97 363 98 364
rect 96 363 97 364
rect 95 363 96 364
rect 94 363 95 364
rect 93 363 94 364
rect 92 363 93 364
rect 91 363 92 364
rect 90 363 91 364
rect 89 363 90 364
rect 88 363 89 364
rect 87 363 88 364
rect 86 363 87 364
rect 85 363 86 364
rect 84 363 85 364
rect 439 364 440 365
rect 438 364 439 365
rect 437 364 438 365
rect 436 364 437 365
rect 435 364 436 365
rect 434 364 435 365
rect 433 364 434 365
rect 432 364 433 365
rect 431 364 432 365
rect 405 364 406 365
rect 404 364 405 365
rect 403 364 404 365
rect 402 364 403 365
rect 401 364 402 365
rect 400 364 401 365
rect 399 364 400 365
rect 398 364 399 365
rect 397 364 398 365
rect 105 364 106 365
rect 104 364 105 365
rect 103 364 104 365
rect 102 364 103 365
rect 101 364 102 365
rect 100 364 101 365
rect 99 364 100 365
rect 98 364 99 365
rect 97 364 98 365
rect 96 364 97 365
rect 95 364 96 365
rect 94 364 95 365
rect 93 364 94 365
rect 92 364 93 365
rect 91 364 92 365
rect 439 365 440 366
rect 438 365 439 366
rect 437 365 438 366
rect 436 365 437 366
rect 435 365 436 366
rect 434 365 435 366
rect 433 365 434 366
rect 432 365 433 366
rect 431 365 432 366
rect 430 365 431 366
rect 429 365 430 366
rect 438 366 439 367
rect 437 366 438 367
rect 436 366 437 367
rect 435 366 436 367
rect 434 366 435 367
rect 433 366 434 367
rect 432 366 433 367
rect 431 366 432 367
rect 430 366 431 367
rect 429 366 430 367
rect 428 366 429 367
rect 433 367 434 368
rect 432 367 433 368
rect 431 367 432 368
rect 430 367 431 368
rect 429 367 430 368
rect 428 367 429 368
rect 439 374 440 375
rect 438 374 439 375
rect 439 375 440 376
rect 438 375 439 376
rect 437 375 438 376
rect 397 375 398 376
rect 396 375 397 376
rect 395 375 396 376
rect 439 376 440 377
rect 438 376 439 377
rect 437 376 438 377
rect 397 376 398 377
rect 396 376 397 377
rect 395 376 396 377
rect 439 377 440 378
rect 438 377 439 378
rect 437 377 438 378
rect 397 377 398 378
rect 396 377 397 378
rect 395 377 396 378
rect 439 378 440 379
rect 438 378 439 379
rect 437 378 438 379
rect 397 378 398 379
rect 396 378 397 379
rect 395 378 396 379
rect 439 379 440 380
rect 438 379 439 380
rect 437 379 438 380
rect 436 379 437 380
rect 398 379 399 380
rect 397 379 398 380
rect 396 379 397 380
rect 395 379 396 380
rect 439 380 440 381
rect 438 380 439 381
rect 437 380 438 381
rect 436 380 437 381
rect 435 380 436 381
rect 434 380 435 381
rect 433 380 434 381
rect 432 380 433 381
rect 431 380 432 381
rect 430 380 431 381
rect 429 380 430 381
rect 428 380 429 381
rect 427 380 428 381
rect 426 380 427 381
rect 425 380 426 381
rect 424 380 425 381
rect 423 380 424 381
rect 422 380 423 381
rect 421 380 422 381
rect 420 380 421 381
rect 419 380 420 381
rect 418 380 419 381
rect 417 380 418 381
rect 416 380 417 381
rect 415 380 416 381
rect 414 380 415 381
rect 413 380 414 381
rect 412 380 413 381
rect 411 380 412 381
rect 410 380 411 381
rect 409 380 410 381
rect 408 380 409 381
rect 407 380 408 381
rect 406 380 407 381
rect 405 380 406 381
rect 404 380 405 381
rect 403 380 404 381
rect 402 380 403 381
rect 401 380 402 381
rect 400 380 401 381
rect 399 380 400 381
rect 398 380 399 381
rect 397 380 398 381
rect 396 380 397 381
rect 395 380 396 381
rect 439 381 440 382
rect 438 381 439 382
rect 437 381 438 382
rect 436 381 437 382
rect 435 381 436 382
rect 434 381 435 382
rect 433 381 434 382
rect 432 381 433 382
rect 431 381 432 382
rect 430 381 431 382
rect 429 381 430 382
rect 428 381 429 382
rect 427 381 428 382
rect 426 381 427 382
rect 425 381 426 382
rect 424 381 425 382
rect 423 381 424 382
rect 422 381 423 382
rect 421 381 422 382
rect 420 381 421 382
rect 419 381 420 382
rect 418 381 419 382
rect 417 381 418 382
rect 416 381 417 382
rect 415 381 416 382
rect 414 381 415 382
rect 413 381 414 382
rect 412 381 413 382
rect 411 381 412 382
rect 410 381 411 382
rect 409 381 410 382
rect 408 381 409 382
rect 407 381 408 382
rect 406 381 407 382
rect 405 381 406 382
rect 404 381 405 382
rect 403 381 404 382
rect 402 381 403 382
rect 401 381 402 382
rect 400 381 401 382
rect 399 381 400 382
rect 398 381 399 382
rect 397 381 398 382
rect 396 381 397 382
rect 395 381 396 382
rect 439 382 440 383
rect 438 382 439 383
rect 437 382 438 383
rect 436 382 437 383
rect 435 382 436 383
rect 434 382 435 383
rect 433 382 434 383
rect 432 382 433 383
rect 431 382 432 383
rect 430 382 431 383
rect 429 382 430 383
rect 428 382 429 383
rect 427 382 428 383
rect 426 382 427 383
rect 425 382 426 383
rect 424 382 425 383
rect 423 382 424 383
rect 422 382 423 383
rect 421 382 422 383
rect 420 382 421 383
rect 419 382 420 383
rect 418 382 419 383
rect 417 382 418 383
rect 416 382 417 383
rect 415 382 416 383
rect 414 382 415 383
rect 413 382 414 383
rect 412 382 413 383
rect 411 382 412 383
rect 410 382 411 383
rect 409 382 410 383
rect 408 382 409 383
rect 407 382 408 383
rect 406 382 407 383
rect 405 382 406 383
rect 404 382 405 383
rect 403 382 404 383
rect 402 382 403 383
rect 401 382 402 383
rect 400 382 401 383
rect 399 382 400 383
rect 398 382 399 383
rect 397 382 398 383
rect 396 382 397 383
rect 395 382 396 383
rect 439 383 440 384
rect 438 383 439 384
rect 437 383 438 384
rect 436 383 437 384
rect 435 383 436 384
rect 434 383 435 384
rect 433 383 434 384
rect 432 383 433 384
rect 431 383 432 384
rect 430 383 431 384
rect 429 383 430 384
rect 428 383 429 384
rect 427 383 428 384
rect 426 383 427 384
rect 425 383 426 384
rect 424 383 425 384
rect 423 383 424 384
rect 422 383 423 384
rect 421 383 422 384
rect 420 383 421 384
rect 419 383 420 384
rect 418 383 419 384
rect 417 383 418 384
rect 416 383 417 384
rect 415 383 416 384
rect 414 383 415 384
rect 413 383 414 384
rect 412 383 413 384
rect 411 383 412 384
rect 410 383 411 384
rect 409 383 410 384
rect 408 383 409 384
rect 407 383 408 384
rect 406 383 407 384
rect 405 383 406 384
rect 404 383 405 384
rect 403 383 404 384
rect 402 383 403 384
rect 401 383 402 384
rect 400 383 401 384
rect 399 383 400 384
rect 398 383 399 384
rect 397 383 398 384
rect 396 383 397 384
rect 395 383 396 384
rect 439 384 440 385
rect 438 384 439 385
rect 437 384 438 385
rect 436 384 437 385
rect 435 384 436 385
rect 434 384 435 385
rect 433 384 434 385
rect 432 384 433 385
rect 431 384 432 385
rect 430 384 431 385
rect 429 384 430 385
rect 428 384 429 385
rect 427 384 428 385
rect 426 384 427 385
rect 425 384 426 385
rect 424 384 425 385
rect 423 384 424 385
rect 422 384 423 385
rect 421 384 422 385
rect 420 384 421 385
rect 419 384 420 385
rect 418 384 419 385
rect 417 384 418 385
rect 416 384 417 385
rect 415 384 416 385
rect 414 384 415 385
rect 413 384 414 385
rect 412 384 413 385
rect 411 384 412 385
rect 410 384 411 385
rect 409 384 410 385
rect 408 384 409 385
rect 407 384 408 385
rect 406 384 407 385
rect 405 384 406 385
rect 404 384 405 385
rect 403 384 404 385
rect 402 384 403 385
rect 401 384 402 385
rect 400 384 401 385
rect 399 384 400 385
rect 398 384 399 385
rect 397 384 398 385
rect 396 384 397 385
rect 395 384 396 385
rect 439 385 440 386
rect 438 385 439 386
rect 437 385 438 386
rect 436 385 437 386
rect 435 385 436 386
rect 434 385 435 386
rect 433 385 434 386
rect 432 385 433 386
rect 431 385 432 386
rect 430 385 431 386
rect 429 385 430 386
rect 428 385 429 386
rect 427 385 428 386
rect 426 385 427 386
rect 425 385 426 386
rect 424 385 425 386
rect 423 385 424 386
rect 422 385 423 386
rect 421 385 422 386
rect 420 385 421 386
rect 419 385 420 386
rect 418 385 419 386
rect 417 385 418 386
rect 416 385 417 386
rect 415 385 416 386
rect 414 385 415 386
rect 413 385 414 386
rect 412 385 413 386
rect 411 385 412 386
rect 410 385 411 386
rect 409 385 410 386
rect 408 385 409 386
rect 407 385 408 386
rect 406 385 407 386
rect 405 385 406 386
rect 404 385 405 386
rect 403 385 404 386
rect 402 385 403 386
rect 401 385 402 386
rect 400 385 401 386
rect 399 385 400 386
rect 398 385 399 386
rect 397 385 398 386
rect 396 385 397 386
rect 395 385 396 386
rect 439 386 440 387
rect 438 386 439 387
rect 437 386 438 387
rect 436 386 437 387
rect 435 386 436 387
rect 434 386 435 387
rect 433 386 434 387
rect 432 386 433 387
rect 431 386 432 387
rect 430 386 431 387
rect 429 386 430 387
rect 428 386 429 387
rect 427 386 428 387
rect 426 386 427 387
rect 425 386 426 387
rect 424 386 425 387
rect 423 386 424 387
rect 422 386 423 387
rect 421 386 422 387
rect 420 386 421 387
rect 419 386 420 387
rect 418 386 419 387
rect 417 386 418 387
rect 416 386 417 387
rect 415 386 416 387
rect 414 386 415 387
rect 413 386 414 387
rect 412 386 413 387
rect 411 386 412 387
rect 410 386 411 387
rect 409 386 410 387
rect 408 386 409 387
rect 407 386 408 387
rect 406 386 407 387
rect 405 386 406 387
rect 404 386 405 387
rect 403 386 404 387
rect 402 386 403 387
rect 401 386 402 387
rect 400 386 401 387
rect 399 386 400 387
rect 398 386 399 387
rect 397 386 398 387
rect 396 386 397 387
rect 395 386 396 387
rect 439 387 440 388
rect 438 387 439 388
rect 437 387 438 388
rect 436 387 437 388
rect 435 387 436 388
rect 434 387 435 388
rect 433 387 434 388
rect 432 387 433 388
rect 431 387 432 388
rect 430 387 431 388
rect 429 387 430 388
rect 428 387 429 388
rect 427 387 428 388
rect 426 387 427 388
rect 425 387 426 388
rect 424 387 425 388
rect 423 387 424 388
rect 422 387 423 388
rect 421 387 422 388
rect 420 387 421 388
rect 419 387 420 388
rect 418 387 419 388
rect 417 387 418 388
rect 416 387 417 388
rect 415 387 416 388
rect 414 387 415 388
rect 413 387 414 388
rect 412 387 413 388
rect 411 387 412 388
rect 410 387 411 388
rect 409 387 410 388
rect 408 387 409 388
rect 407 387 408 388
rect 406 387 407 388
rect 405 387 406 388
rect 404 387 405 388
rect 403 387 404 388
rect 402 387 403 388
rect 401 387 402 388
rect 400 387 401 388
rect 399 387 400 388
rect 398 387 399 388
rect 397 387 398 388
rect 396 387 397 388
rect 395 387 396 388
rect 439 388 440 389
rect 438 388 439 389
rect 437 388 438 389
rect 436 388 437 389
rect 435 388 436 389
rect 434 388 435 389
rect 433 388 434 389
rect 432 388 433 389
rect 431 388 432 389
rect 430 388 431 389
rect 429 388 430 389
rect 428 388 429 389
rect 427 388 428 389
rect 426 388 427 389
rect 425 388 426 389
rect 424 388 425 389
rect 423 388 424 389
rect 422 388 423 389
rect 421 388 422 389
rect 420 388 421 389
rect 419 388 420 389
rect 418 388 419 389
rect 417 388 418 389
rect 416 388 417 389
rect 415 388 416 389
rect 414 388 415 389
rect 413 388 414 389
rect 412 388 413 389
rect 411 388 412 389
rect 410 388 411 389
rect 409 388 410 389
rect 408 388 409 389
rect 407 388 408 389
rect 406 388 407 389
rect 405 388 406 389
rect 404 388 405 389
rect 403 388 404 389
rect 402 388 403 389
rect 401 388 402 389
rect 400 388 401 389
rect 399 388 400 389
rect 398 388 399 389
rect 397 388 398 389
rect 396 388 397 389
rect 395 388 396 389
rect 439 389 440 390
rect 438 389 439 390
rect 437 389 438 390
rect 436 389 437 390
rect 435 389 436 390
rect 434 389 435 390
rect 433 389 434 390
rect 432 389 433 390
rect 431 389 432 390
rect 430 389 431 390
rect 429 389 430 390
rect 428 389 429 390
rect 427 389 428 390
rect 426 389 427 390
rect 425 389 426 390
rect 424 389 425 390
rect 423 389 424 390
rect 422 389 423 390
rect 421 389 422 390
rect 420 389 421 390
rect 419 389 420 390
rect 418 389 419 390
rect 417 389 418 390
rect 416 389 417 390
rect 415 389 416 390
rect 414 389 415 390
rect 413 389 414 390
rect 412 389 413 390
rect 411 389 412 390
rect 410 389 411 390
rect 409 389 410 390
rect 408 389 409 390
rect 407 389 408 390
rect 406 389 407 390
rect 405 389 406 390
rect 404 389 405 390
rect 403 389 404 390
rect 402 389 403 390
rect 401 389 402 390
rect 400 389 401 390
rect 399 389 400 390
rect 398 389 399 390
rect 397 389 398 390
rect 396 389 397 390
rect 395 389 396 390
rect 439 390 440 391
rect 438 390 439 391
rect 437 390 438 391
rect 436 390 437 391
rect 435 390 436 391
rect 418 390 419 391
rect 417 390 418 391
rect 416 390 417 391
rect 415 390 416 391
rect 398 390 399 391
rect 397 390 398 391
rect 396 390 397 391
rect 395 390 396 391
rect 439 391 440 392
rect 438 391 439 392
rect 437 391 438 392
rect 436 391 437 392
rect 418 391 419 392
rect 417 391 418 392
rect 416 391 417 392
rect 415 391 416 392
rect 397 391 398 392
rect 396 391 397 392
rect 395 391 396 392
rect 439 392 440 393
rect 438 392 439 393
rect 437 392 438 393
rect 418 392 419 393
rect 417 392 418 393
rect 416 392 417 393
rect 415 392 416 393
rect 397 392 398 393
rect 396 392 397 393
rect 395 392 396 393
rect 439 393 440 394
rect 438 393 439 394
rect 437 393 438 394
rect 418 393 419 394
rect 417 393 418 394
rect 416 393 417 394
rect 415 393 416 394
rect 397 393 398 394
rect 396 393 397 394
rect 395 393 396 394
rect 439 394 440 395
rect 438 394 439 395
rect 437 394 438 395
rect 418 394 419 395
rect 417 394 418 395
rect 416 394 417 395
rect 415 394 416 395
rect 397 394 398 395
rect 396 394 397 395
rect 395 394 396 395
rect 439 395 440 396
rect 438 395 439 396
rect 437 395 438 396
rect 418 395 419 396
rect 417 395 418 396
rect 416 395 417 396
rect 415 395 416 396
rect 397 395 398 396
rect 396 395 397 396
rect 395 395 396 396
rect 439 396 440 397
rect 438 396 439 397
rect 437 396 438 397
rect 418 396 419 397
rect 417 396 418 397
rect 416 396 417 397
rect 415 396 416 397
rect 397 396 398 397
rect 396 396 397 397
rect 395 396 396 397
rect 439 397 440 398
rect 438 397 439 398
rect 437 397 438 398
rect 418 397 419 398
rect 417 397 418 398
rect 416 397 417 398
rect 415 397 416 398
rect 397 397 398 398
rect 396 397 397 398
rect 395 397 396 398
rect 439 398 440 399
rect 438 398 439 399
rect 437 398 438 399
rect 418 398 419 399
rect 417 398 418 399
rect 416 398 417 399
rect 415 398 416 399
rect 397 398 398 399
rect 396 398 397 399
rect 395 398 396 399
rect 439 399 440 400
rect 438 399 439 400
rect 437 399 438 400
rect 418 399 419 400
rect 417 399 418 400
rect 416 399 417 400
rect 415 399 416 400
rect 398 399 399 400
rect 397 399 398 400
rect 396 399 397 400
rect 395 399 396 400
rect 439 400 440 401
rect 438 400 439 401
rect 437 400 438 401
rect 419 400 420 401
rect 418 400 419 401
rect 417 400 418 401
rect 416 400 417 401
rect 415 400 416 401
rect 414 400 415 401
rect 398 400 399 401
rect 397 400 398 401
rect 396 400 397 401
rect 395 400 396 401
rect 439 401 440 402
rect 438 401 439 402
rect 437 401 438 402
rect 421 401 422 402
rect 420 401 421 402
rect 419 401 420 402
rect 418 401 419 402
rect 417 401 418 402
rect 416 401 417 402
rect 415 401 416 402
rect 414 401 415 402
rect 413 401 414 402
rect 412 401 413 402
rect 398 401 399 402
rect 397 401 398 402
rect 396 401 397 402
rect 395 401 396 402
rect 439 402 440 403
rect 438 402 439 403
rect 437 402 438 403
rect 436 402 437 403
rect 423 402 424 403
rect 422 402 423 403
rect 421 402 422 403
rect 420 402 421 403
rect 419 402 420 403
rect 418 402 419 403
rect 417 402 418 403
rect 416 402 417 403
rect 415 402 416 403
rect 414 402 415 403
rect 413 402 414 403
rect 412 402 413 403
rect 411 402 412 403
rect 410 402 411 403
rect 399 402 400 403
rect 398 402 399 403
rect 397 402 398 403
rect 396 402 397 403
rect 395 402 396 403
rect 439 403 440 404
rect 438 403 439 404
rect 437 403 438 404
rect 436 403 437 404
rect 423 403 424 404
rect 422 403 423 404
rect 421 403 422 404
rect 420 403 421 404
rect 419 403 420 404
rect 418 403 419 404
rect 417 403 418 404
rect 416 403 417 404
rect 415 403 416 404
rect 414 403 415 404
rect 413 403 414 404
rect 412 403 413 404
rect 411 403 412 404
rect 410 403 411 404
rect 400 403 401 404
rect 399 403 400 404
rect 398 403 399 404
rect 397 403 398 404
rect 396 403 397 404
rect 395 403 396 404
rect 439 404 440 405
rect 438 404 439 405
rect 437 404 438 405
rect 436 404 437 405
rect 435 404 436 405
rect 423 404 424 405
rect 422 404 423 405
rect 421 404 422 405
rect 420 404 421 405
rect 419 404 420 405
rect 418 404 419 405
rect 417 404 418 405
rect 416 404 417 405
rect 415 404 416 405
rect 414 404 415 405
rect 413 404 414 405
rect 412 404 413 405
rect 411 404 412 405
rect 410 404 411 405
rect 402 404 403 405
rect 401 404 402 405
rect 400 404 401 405
rect 399 404 400 405
rect 398 404 399 405
rect 397 404 398 405
rect 396 404 397 405
rect 395 404 396 405
rect 439 405 440 406
rect 438 405 439 406
rect 437 405 438 406
rect 436 405 437 406
rect 435 405 436 406
rect 434 405 435 406
rect 405 405 406 406
rect 404 405 405 406
rect 403 405 404 406
rect 402 405 403 406
rect 401 405 402 406
rect 400 405 401 406
rect 399 405 400 406
rect 398 405 399 406
rect 397 405 398 406
rect 396 405 397 406
rect 395 405 396 406
rect 439 406 440 407
rect 438 406 439 407
rect 437 406 438 407
rect 436 406 437 407
rect 435 406 436 407
rect 434 406 435 407
rect 433 406 434 407
rect 405 406 406 407
rect 404 406 405 407
rect 403 406 404 407
rect 402 406 403 407
rect 401 406 402 407
rect 400 406 401 407
rect 399 406 400 407
rect 398 406 399 407
rect 397 406 398 407
rect 396 406 397 407
rect 395 406 396 407
rect 439 407 440 408
rect 438 407 439 408
rect 437 407 438 408
rect 436 407 437 408
rect 435 407 436 408
rect 434 407 435 408
rect 433 407 434 408
rect 432 407 433 408
rect 431 407 432 408
rect 405 407 406 408
rect 404 407 405 408
rect 403 407 404 408
rect 402 407 403 408
rect 401 407 402 408
rect 400 407 401 408
rect 399 407 400 408
rect 398 407 399 408
rect 397 407 398 408
rect 396 407 397 408
rect 395 407 396 408
rect 439 408 440 409
rect 438 408 439 409
rect 437 408 438 409
rect 436 408 437 409
rect 435 408 436 409
rect 434 408 435 409
rect 433 408 434 409
rect 432 408 433 409
rect 431 408 432 409
rect 430 408 431 409
rect 429 408 430 409
rect 438 409 439 410
rect 437 409 438 410
rect 436 409 437 410
rect 435 409 436 410
rect 434 409 435 410
rect 433 409 434 410
rect 432 409 433 410
rect 431 409 432 410
rect 430 409 431 410
rect 429 409 430 410
rect 428 409 429 410
rect 434 410 435 411
rect 433 410 434 411
rect 432 410 433 411
rect 431 410 432 411
rect 430 410 431 411
rect 429 410 430 411
rect 428 410 429 411
rect 429 411 430 412
rect 428 411 429 412
<< metal3 >>
rect 441 4 442 5
rect 440 4 441 5
rect 399 4 400 5
rect 398 4 399 5
rect 397 4 398 5
rect 441 5 442 6
rect 440 5 441 6
rect 439 5 440 6
rect 399 5 400 6
rect 398 5 399 6
rect 397 5 398 6
rect 441 6 442 7
rect 440 6 441 7
rect 439 6 440 7
rect 399 6 400 7
rect 398 6 399 7
rect 397 6 398 7
rect 441 7 442 8
rect 440 7 441 8
rect 439 7 440 8
rect 399 7 400 8
rect 398 7 399 8
rect 397 7 398 8
rect 441 8 442 9
rect 440 8 441 9
rect 439 8 440 9
rect 400 8 401 9
rect 399 8 400 9
rect 398 8 399 9
rect 397 8 398 9
rect 441 9 442 10
rect 440 9 441 10
rect 439 9 440 10
rect 438 9 439 10
rect 437 9 438 10
rect 401 9 402 10
rect 400 9 401 10
rect 399 9 400 10
rect 398 9 399 10
rect 397 9 398 10
rect 441 10 442 11
rect 440 10 441 11
rect 439 10 440 11
rect 438 10 439 11
rect 437 10 438 11
rect 436 10 437 11
rect 435 10 436 11
rect 434 10 435 11
rect 433 10 434 11
rect 432 10 433 11
rect 431 10 432 11
rect 430 10 431 11
rect 429 10 430 11
rect 428 10 429 11
rect 427 10 428 11
rect 426 10 427 11
rect 425 10 426 11
rect 424 10 425 11
rect 423 10 424 11
rect 422 10 423 11
rect 421 10 422 11
rect 420 10 421 11
rect 419 10 420 11
rect 418 10 419 11
rect 417 10 418 11
rect 416 10 417 11
rect 415 10 416 11
rect 414 10 415 11
rect 413 10 414 11
rect 412 10 413 11
rect 411 10 412 11
rect 410 10 411 11
rect 409 10 410 11
rect 408 10 409 11
rect 407 10 408 11
rect 406 10 407 11
rect 405 10 406 11
rect 404 10 405 11
rect 403 10 404 11
rect 402 10 403 11
rect 401 10 402 11
rect 400 10 401 11
rect 399 10 400 11
rect 398 10 399 11
rect 397 10 398 11
rect 441 11 442 12
rect 440 11 441 12
rect 439 11 440 12
rect 438 11 439 12
rect 437 11 438 12
rect 436 11 437 12
rect 435 11 436 12
rect 434 11 435 12
rect 433 11 434 12
rect 432 11 433 12
rect 431 11 432 12
rect 430 11 431 12
rect 429 11 430 12
rect 428 11 429 12
rect 427 11 428 12
rect 426 11 427 12
rect 425 11 426 12
rect 424 11 425 12
rect 423 11 424 12
rect 422 11 423 12
rect 421 11 422 12
rect 420 11 421 12
rect 419 11 420 12
rect 418 11 419 12
rect 417 11 418 12
rect 416 11 417 12
rect 415 11 416 12
rect 414 11 415 12
rect 413 11 414 12
rect 412 11 413 12
rect 411 11 412 12
rect 410 11 411 12
rect 409 11 410 12
rect 408 11 409 12
rect 407 11 408 12
rect 406 11 407 12
rect 405 11 406 12
rect 404 11 405 12
rect 403 11 404 12
rect 402 11 403 12
rect 401 11 402 12
rect 400 11 401 12
rect 399 11 400 12
rect 398 11 399 12
rect 397 11 398 12
rect 441 12 442 13
rect 440 12 441 13
rect 439 12 440 13
rect 438 12 439 13
rect 437 12 438 13
rect 436 12 437 13
rect 435 12 436 13
rect 434 12 435 13
rect 433 12 434 13
rect 432 12 433 13
rect 431 12 432 13
rect 430 12 431 13
rect 429 12 430 13
rect 428 12 429 13
rect 427 12 428 13
rect 426 12 427 13
rect 425 12 426 13
rect 424 12 425 13
rect 423 12 424 13
rect 422 12 423 13
rect 421 12 422 13
rect 420 12 421 13
rect 419 12 420 13
rect 418 12 419 13
rect 417 12 418 13
rect 416 12 417 13
rect 415 12 416 13
rect 414 12 415 13
rect 413 12 414 13
rect 412 12 413 13
rect 411 12 412 13
rect 410 12 411 13
rect 409 12 410 13
rect 408 12 409 13
rect 407 12 408 13
rect 406 12 407 13
rect 405 12 406 13
rect 404 12 405 13
rect 403 12 404 13
rect 402 12 403 13
rect 401 12 402 13
rect 400 12 401 13
rect 399 12 400 13
rect 398 12 399 13
rect 397 12 398 13
rect 441 13 442 14
rect 440 13 441 14
rect 439 13 440 14
rect 438 13 439 14
rect 437 13 438 14
rect 436 13 437 14
rect 435 13 436 14
rect 434 13 435 14
rect 433 13 434 14
rect 432 13 433 14
rect 431 13 432 14
rect 430 13 431 14
rect 429 13 430 14
rect 428 13 429 14
rect 427 13 428 14
rect 426 13 427 14
rect 425 13 426 14
rect 424 13 425 14
rect 423 13 424 14
rect 422 13 423 14
rect 421 13 422 14
rect 420 13 421 14
rect 419 13 420 14
rect 418 13 419 14
rect 417 13 418 14
rect 416 13 417 14
rect 415 13 416 14
rect 414 13 415 14
rect 413 13 414 14
rect 412 13 413 14
rect 411 13 412 14
rect 410 13 411 14
rect 409 13 410 14
rect 408 13 409 14
rect 407 13 408 14
rect 406 13 407 14
rect 405 13 406 14
rect 404 13 405 14
rect 403 13 404 14
rect 402 13 403 14
rect 401 13 402 14
rect 400 13 401 14
rect 399 13 400 14
rect 398 13 399 14
rect 397 13 398 14
rect 441 14 442 15
rect 440 14 441 15
rect 439 14 440 15
rect 438 14 439 15
rect 437 14 438 15
rect 436 14 437 15
rect 435 14 436 15
rect 434 14 435 15
rect 433 14 434 15
rect 432 14 433 15
rect 431 14 432 15
rect 430 14 431 15
rect 429 14 430 15
rect 428 14 429 15
rect 427 14 428 15
rect 426 14 427 15
rect 425 14 426 15
rect 424 14 425 15
rect 423 14 424 15
rect 422 14 423 15
rect 421 14 422 15
rect 420 14 421 15
rect 419 14 420 15
rect 418 14 419 15
rect 417 14 418 15
rect 416 14 417 15
rect 415 14 416 15
rect 414 14 415 15
rect 413 14 414 15
rect 412 14 413 15
rect 411 14 412 15
rect 410 14 411 15
rect 409 14 410 15
rect 408 14 409 15
rect 407 14 408 15
rect 406 14 407 15
rect 405 14 406 15
rect 404 14 405 15
rect 403 14 404 15
rect 402 14 403 15
rect 401 14 402 15
rect 400 14 401 15
rect 399 14 400 15
rect 398 14 399 15
rect 397 14 398 15
rect 441 15 442 16
rect 440 15 441 16
rect 439 15 440 16
rect 438 15 439 16
rect 437 15 438 16
rect 436 15 437 16
rect 435 15 436 16
rect 434 15 435 16
rect 433 15 434 16
rect 432 15 433 16
rect 431 15 432 16
rect 430 15 431 16
rect 429 15 430 16
rect 428 15 429 16
rect 427 15 428 16
rect 426 15 427 16
rect 425 15 426 16
rect 424 15 425 16
rect 423 15 424 16
rect 422 15 423 16
rect 421 15 422 16
rect 420 15 421 16
rect 419 15 420 16
rect 418 15 419 16
rect 417 15 418 16
rect 416 15 417 16
rect 415 15 416 16
rect 414 15 415 16
rect 413 15 414 16
rect 412 15 413 16
rect 411 15 412 16
rect 410 15 411 16
rect 409 15 410 16
rect 408 15 409 16
rect 407 15 408 16
rect 406 15 407 16
rect 405 15 406 16
rect 404 15 405 16
rect 403 15 404 16
rect 402 15 403 16
rect 401 15 402 16
rect 400 15 401 16
rect 399 15 400 16
rect 398 15 399 16
rect 397 15 398 16
rect 441 16 442 17
rect 440 16 441 17
rect 439 16 440 17
rect 438 16 439 17
rect 437 16 438 17
rect 436 16 437 17
rect 435 16 436 17
rect 434 16 435 17
rect 433 16 434 17
rect 432 16 433 17
rect 431 16 432 17
rect 430 16 431 17
rect 429 16 430 17
rect 428 16 429 17
rect 427 16 428 17
rect 426 16 427 17
rect 425 16 426 17
rect 424 16 425 17
rect 423 16 424 17
rect 422 16 423 17
rect 421 16 422 17
rect 420 16 421 17
rect 419 16 420 17
rect 418 16 419 17
rect 417 16 418 17
rect 416 16 417 17
rect 415 16 416 17
rect 414 16 415 17
rect 413 16 414 17
rect 412 16 413 17
rect 411 16 412 17
rect 410 16 411 17
rect 409 16 410 17
rect 408 16 409 17
rect 407 16 408 17
rect 406 16 407 17
rect 405 16 406 17
rect 404 16 405 17
rect 403 16 404 17
rect 402 16 403 17
rect 401 16 402 17
rect 400 16 401 17
rect 399 16 400 17
rect 398 16 399 17
rect 397 16 398 17
rect 441 17 442 18
rect 440 17 441 18
rect 439 17 440 18
rect 438 17 439 18
rect 437 17 438 18
rect 436 17 437 18
rect 435 17 436 18
rect 434 17 435 18
rect 433 17 434 18
rect 432 17 433 18
rect 431 17 432 18
rect 430 17 431 18
rect 429 17 430 18
rect 428 17 429 18
rect 427 17 428 18
rect 426 17 427 18
rect 425 17 426 18
rect 424 17 425 18
rect 423 17 424 18
rect 422 17 423 18
rect 421 17 422 18
rect 420 17 421 18
rect 419 17 420 18
rect 418 17 419 18
rect 417 17 418 18
rect 416 17 417 18
rect 415 17 416 18
rect 414 17 415 18
rect 413 17 414 18
rect 412 17 413 18
rect 411 17 412 18
rect 410 17 411 18
rect 409 17 410 18
rect 408 17 409 18
rect 407 17 408 18
rect 406 17 407 18
rect 405 17 406 18
rect 404 17 405 18
rect 403 17 404 18
rect 402 17 403 18
rect 401 17 402 18
rect 400 17 401 18
rect 399 17 400 18
rect 398 17 399 18
rect 397 17 398 18
rect 441 18 442 19
rect 440 18 441 19
rect 439 18 440 19
rect 438 18 439 19
rect 437 18 438 19
rect 436 18 437 19
rect 435 18 436 19
rect 434 18 435 19
rect 433 18 434 19
rect 432 18 433 19
rect 431 18 432 19
rect 430 18 431 19
rect 429 18 430 19
rect 428 18 429 19
rect 427 18 428 19
rect 426 18 427 19
rect 425 18 426 19
rect 424 18 425 19
rect 423 18 424 19
rect 422 18 423 19
rect 421 18 422 19
rect 420 18 421 19
rect 419 18 420 19
rect 418 18 419 19
rect 417 18 418 19
rect 416 18 417 19
rect 415 18 416 19
rect 414 18 415 19
rect 413 18 414 19
rect 412 18 413 19
rect 411 18 412 19
rect 410 18 411 19
rect 409 18 410 19
rect 408 18 409 19
rect 407 18 408 19
rect 406 18 407 19
rect 405 18 406 19
rect 404 18 405 19
rect 403 18 404 19
rect 402 18 403 19
rect 401 18 402 19
rect 400 18 401 19
rect 399 18 400 19
rect 398 18 399 19
rect 397 18 398 19
rect 441 19 442 20
rect 440 19 441 20
rect 439 19 440 20
rect 438 19 439 20
rect 437 19 438 20
rect 420 19 421 20
rect 419 19 420 20
rect 418 19 419 20
rect 401 19 402 20
rect 400 19 401 20
rect 399 19 400 20
rect 398 19 399 20
rect 397 19 398 20
rect 441 20 442 21
rect 440 20 441 21
rect 439 20 440 21
rect 438 20 439 21
rect 420 20 421 21
rect 419 20 420 21
rect 418 20 419 21
rect 417 20 418 21
rect 400 20 401 21
rect 399 20 400 21
rect 398 20 399 21
rect 397 20 398 21
rect 441 21 442 22
rect 440 21 441 22
rect 439 21 440 22
rect 421 21 422 22
rect 420 21 421 22
rect 419 21 420 22
rect 418 21 419 22
rect 417 21 418 22
rect 399 21 400 22
rect 398 21 399 22
rect 397 21 398 22
rect 441 22 442 23
rect 440 22 441 23
rect 439 22 440 23
rect 422 22 423 23
rect 421 22 422 23
rect 420 22 421 23
rect 419 22 420 23
rect 418 22 419 23
rect 417 22 418 23
rect 416 22 417 23
rect 399 22 400 23
rect 398 22 399 23
rect 397 22 398 23
rect 441 23 442 24
rect 440 23 441 24
rect 439 23 440 24
rect 423 23 424 24
rect 422 23 423 24
rect 421 23 422 24
rect 420 23 421 24
rect 419 23 420 24
rect 418 23 419 24
rect 417 23 418 24
rect 416 23 417 24
rect 415 23 416 24
rect 399 23 400 24
rect 398 23 399 24
rect 397 23 398 24
rect 441 24 442 25
rect 440 24 441 25
rect 439 24 440 25
rect 425 24 426 25
rect 424 24 425 25
rect 423 24 424 25
rect 422 24 423 25
rect 421 24 422 25
rect 420 24 421 25
rect 419 24 420 25
rect 418 24 419 25
rect 417 24 418 25
rect 416 24 417 25
rect 415 24 416 25
rect 414 24 415 25
rect 399 24 400 25
rect 398 24 399 25
rect 397 24 398 25
rect 426 25 427 26
rect 425 25 426 26
rect 424 25 425 26
rect 423 25 424 26
rect 422 25 423 26
rect 421 25 422 26
rect 420 25 421 26
rect 419 25 420 26
rect 418 25 419 26
rect 417 25 418 26
rect 416 25 417 26
rect 415 25 416 26
rect 414 25 415 26
rect 413 25 414 26
rect 428 26 429 27
rect 427 26 428 27
rect 426 26 427 27
rect 425 26 426 27
rect 424 26 425 27
rect 423 26 424 27
rect 422 26 423 27
rect 421 26 422 27
rect 420 26 421 27
rect 419 26 420 27
rect 418 26 419 27
rect 417 26 418 27
rect 416 26 417 27
rect 415 26 416 27
rect 414 26 415 27
rect 413 26 414 27
rect 412 26 413 27
rect 429 27 430 28
rect 428 27 429 28
rect 427 27 428 28
rect 426 27 427 28
rect 425 27 426 28
rect 424 27 425 28
rect 423 27 424 28
rect 422 27 423 28
rect 421 27 422 28
rect 420 27 421 28
rect 419 27 420 28
rect 418 27 419 28
rect 417 27 418 28
rect 416 27 417 28
rect 415 27 416 28
rect 414 27 415 28
rect 413 27 414 28
rect 412 27 413 28
rect 411 27 412 28
rect 431 28 432 29
rect 430 28 431 29
rect 429 28 430 29
rect 428 28 429 29
rect 427 28 428 29
rect 426 28 427 29
rect 425 28 426 29
rect 424 28 425 29
rect 423 28 424 29
rect 422 28 423 29
rect 421 28 422 29
rect 420 28 421 29
rect 419 28 420 29
rect 418 28 419 29
rect 417 28 418 29
rect 416 28 417 29
rect 415 28 416 29
rect 413 28 414 29
rect 412 28 413 29
rect 411 28 412 29
rect 410 28 411 29
rect 432 29 433 30
rect 431 29 432 30
rect 430 29 431 30
rect 429 29 430 30
rect 428 29 429 30
rect 427 29 428 30
rect 426 29 427 30
rect 425 29 426 30
rect 424 29 425 30
rect 423 29 424 30
rect 422 29 423 30
rect 421 29 422 30
rect 420 29 421 30
rect 419 29 420 30
rect 418 29 419 30
rect 417 29 418 30
rect 412 29 413 30
rect 411 29 412 30
rect 410 29 411 30
rect 409 29 410 30
rect 433 30 434 31
rect 432 30 433 31
rect 431 30 432 31
rect 430 30 431 31
rect 429 30 430 31
rect 428 30 429 31
rect 427 30 428 31
rect 426 30 427 31
rect 425 30 426 31
rect 424 30 425 31
rect 423 30 424 31
rect 422 30 423 31
rect 421 30 422 31
rect 420 30 421 31
rect 419 30 420 31
rect 418 30 419 31
rect 411 30 412 31
rect 410 30 411 31
rect 409 30 410 31
rect 408 30 409 31
rect 435 31 436 32
rect 434 31 435 32
rect 433 31 434 32
rect 432 31 433 32
rect 431 31 432 32
rect 430 31 431 32
rect 429 31 430 32
rect 428 31 429 32
rect 427 31 428 32
rect 426 31 427 32
rect 425 31 426 32
rect 424 31 425 32
rect 423 31 424 32
rect 422 31 423 32
rect 421 31 422 32
rect 420 31 421 32
rect 419 31 420 32
rect 410 31 411 32
rect 409 31 410 32
rect 408 31 409 32
rect 407 31 408 32
rect 406 31 407 32
rect 399 31 400 32
rect 398 31 399 32
rect 397 31 398 32
rect 436 32 437 33
rect 435 32 436 33
rect 434 32 435 33
rect 433 32 434 33
rect 432 32 433 33
rect 431 32 432 33
rect 430 32 431 33
rect 429 32 430 33
rect 428 32 429 33
rect 427 32 428 33
rect 426 32 427 33
rect 425 32 426 33
rect 424 32 425 33
rect 423 32 424 33
rect 422 32 423 33
rect 421 32 422 33
rect 409 32 410 33
rect 408 32 409 33
rect 407 32 408 33
rect 406 32 407 33
rect 405 32 406 33
rect 399 32 400 33
rect 398 32 399 33
rect 397 32 398 33
rect 438 33 439 34
rect 437 33 438 34
rect 436 33 437 34
rect 435 33 436 34
rect 434 33 435 34
rect 433 33 434 34
rect 432 33 433 34
rect 431 33 432 34
rect 430 33 431 34
rect 429 33 430 34
rect 428 33 429 34
rect 427 33 428 34
rect 426 33 427 34
rect 425 33 426 34
rect 424 33 425 34
rect 423 33 424 34
rect 422 33 423 34
rect 408 33 409 34
rect 407 33 408 34
rect 406 33 407 34
rect 405 33 406 34
rect 404 33 405 34
rect 399 33 400 34
rect 398 33 399 34
rect 397 33 398 34
rect 439 34 440 35
rect 438 34 439 35
rect 437 34 438 35
rect 436 34 437 35
rect 435 34 436 35
rect 434 34 435 35
rect 433 34 434 35
rect 432 34 433 35
rect 431 34 432 35
rect 430 34 431 35
rect 429 34 430 35
rect 428 34 429 35
rect 427 34 428 35
rect 426 34 427 35
rect 425 34 426 35
rect 424 34 425 35
rect 407 34 408 35
rect 406 34 407 35
rect 405 34 406 35
rect 404 34 405 35
rect 403 34 404 35
rect 402 34 403 35
rect 399 34 400 35
rect 398 34 399 35
rect 397 34 398 35
rect 441 35 442 36
rect 440 35 441 36
rect 439 35 440 36
rect 438 35 439 36
rect 437 35 438 36
rect 436 35 437 36
rect 435 35 436 36
rect 434 35 435 36
rect 433 35 434 36
rect 432 35 433 36
rect 431 35 432 36
rect 430 35 431 36
rect 429 35 430 36
rect 428 35 429 36
rect 427 35 428 36
rect 426 35 427 36
rect 425 35 426 36
rect 406 35 407 36
rect 405 35 406 36
rect 404 35 405 36
rect 403 35 404 36
rect 402 35 403 36
rect 401 35 402 36
rect 400 35 401 36
rect 399 35 400 36
rect 398 35 399 36
rect 397 35 398 36
rect 441 36 442 37
rect 440 36 441 37
rect 439 36 440 37
rect 438 36 439 37
rect 437 36 438 37
rect 436 36 437 37
rect 435 36 436 37
rect 434 36 435 37
rect 433 36 434 37
rect 432 36 433 37
rect 431 36 432 37
rect 430 36 431 37
rect 429 36 430 37
rect 428 36 429 37
rect 427 36 428 37
rect 426 36 427 37
rect 405 36 406 37
rect 404 36 405 37
rect 403 36 404 37
rect 402 36 403 37
rect 401 36 402 37
rect 400 36 401 37
rect 399 36 400 37
rect 398 36 399 37
rect 397 36 398 37
rect 441 37 442 38
rect 440 37 441 38
rect 439 37 440 38
rect 438 37 439 38
rect 437 37 438 38
rect 436 37 437 38
rect 435 37 436 38
rect 434 37 435 38
rect 433 37 434 38
rect 432 37 433 38
rect 431 37 432 38
rect 430 37 431 38
rect 429 37 430 38
rect 428 37 429 38
rect 404 37 405 38
rect 403 37 404 38
rect 402 37 403 38
rect 401 37 402 38
rect 400 37 401 38
rect 399 37 400 38
rect 398 37 399 38
rect 397 37 398 38
rect 441 38 442 39
rect 440 38 441 39
rect 439 38 440 39
rect 438 38 439 39
rect 437 38 438 39
rect 436 38 437 39
rect 435 38 436 39
rect 434 38 435 39
rect 433 38 434 39
rect 432 38 433 39
rect 431 38 432 39
rect 430 38 431 39
rect 429 38 430 39
rect 403 38 404 39
rect 402 38 403 39
rect 401 38 402 39
rect 400 38 401 39
rect 399 38 400 39
rect 398 38 399 39
rect 397 38 398 39
rect 441 39 442 40
rect 440 39 441 40
rect 439 39 440 40
rect 438 39 439 40
rect 437 39 438 40
rect 436 39 437 40
rect 435 39 436 40
rect 434 39 435 40
rect 433 39 434 40
rect 432 39 433 40
rect 431 39 432 40
rect 430 39 431 40
rect 402 39 403 40
rect 401 39 402 40
rect 400 39 401 40
rect 399 39 400 40
rect 398 39 399 40
rect 397 39 398 40
rect 441 40 442 41
rect 440 40 441 41
rect 439 40 440 41
rect 438 40 439 41
rect 437 40 438 41
rect 436 40 437 41
rect 435 40 436 41
rect 434 40 435 41
rect 433 40 434 41
rect 432 40 433 41
rect 402 40 403 41
rect 401 40 402 41
rect 400 40 401 41
rect 399 40 400 41
rect 398 40 399 41
rect 397 40 398 41
rect 441 41 442 42
rect 440 41 441 42
rect 439 41 440 42
rect 438 41 439 42
rect 437 41 438 42
rect 436 41 437 42
rect 435 41 436 42
rect 434 41 435 42
rect 433 41 434 42
rect 401 41 402 42
rect 400 41 401 42
rect 399 41 400 42
rect 398 41 399 42
rect 397 41 398 42
rect 441 42 442 43
rect 440 42 441 43
rect 439 42 440 43
rect 438 42 439 43
rect 437 42 438 43
rect 436 42 437 43
rect 435 42 436 43
rect 434 42 435 43
rect 400 42 401 43
rect 399 42 400 43
rect 398 42 399 43
rect 397 42 398 43
rect 441 43 442 44
rect 440 43 441 44
rect 439 43 440 44
rect 438 43 439 44
rect 437 43 438 44
rect 436 43 437 44
rect 435 43 436 44
rect 400 43 401 44
rect 399 43 400 44
rect 398 43 399 44
rect 397 43 398 44
rect 441 44 442 45
rect 440 44 441 45
rect 439 44 440 45
rect 438 44 439 45
rect 437 44 438 45
rect 400 44 401 45
rect 399 44 400 45
rect 398 44 399 45
rect 397 44 398 45
rect 441 45 442 46
rect 440 45 441 46
rect 439 45 440 46
rect 438 45 439 46
rect 437 45 438 46
rect 399 45 400 46
rect 398 45 399 46
rect 397 45 398 46
rect 441 46 442 47
rect 440 46 441 47
rect 439 46 440 47
rect 438 46 439 47
rect 399 46 400 47
rect 398 46 399 47
rect 397 46 398 47
rect 441 47 442 48
rect 440 47 441 48
rect 439 47 440 48
rect 399 47 400 48
rect 398 47 399 48
rect 397 47 398 48
rect 441 48 442 49
rect 440 48 441 49
rect 439 48 440 49
rect 399 48 400 49
rect 398 48 399 49
rect 397 48 398 49
rect 441 49 442 50
rect 440 49 441 50
rect 439 49 440 50
rect 93 51 94 52
rect 92 51 93 52
rect 91 51 92 52
rect 90 51 91 52
rect 89 51 90 52
rect 88 51 89 52
rect 95 52 96 53
rect 94 52 95 53
rect 93 52 94 53
rect 92 52 93 53
rect 91 52 92 53
rect 90 52 91 53
rect 89 52 90 53
rect 88 52 89 53
rect 87 52 88 53
rect 86 52 87 53
rect 96 53 97 54
rect 95 53 96 54
rect 94 53 95 54
rect 93 53 94 54
rect 92 53 93 54
rect 91 53 92 54
rect 90 53 91 54
rect 89 53 90 54
rect 88 53 89 54
rect 87 53 88 54
rect 86 53 87 54
rect 85 53 86 54
rect 398 54 399 55
rect 397 54 398 55
rect 96 54 97 55
rect 95 54 96 55
rect 94 54 95 55
rect 93 54 94 55
rect 92 54 93 55
rect 91 54 92 55
rect 90 54 91 55
rect 89 54 90 55
rect 88 54 89 55
rect 87 54 88 55
rect 86 54 87 55
rect 85 54 86 55
rect 84 54 85 55
rect 399 55 400 56
rect 398 55 399 56
rect 397 55 398 56
rect 97 55 98 56
rect 96 55 97 56
rect 95 55 96 56
rect 94 55 95 56
rect 93 55 94 56
rect 92 55 93 56
rect 91 55 92 56
rect 90 55 91 56
rect 89 55 90 56
rect 88 55 89 56
rect 87 55 88 56
rect 86 55 87 56
rect 85 55 86 56
rect 84 55 85 56
rect 83 55 84 56
rect 399 56 400 57
rect 398 56 399 57
rect 397 56 398 57
rect 97 56 98 57
rect 96 56 97 57
rect 95 56 96 57
rect 94 56 95 57
rect 93 56 94 57
rect 92 56 93 57
rect 91 56 92 57
rect 90 56 91 57
rect 89 56 90 57
rect 88 56 89 57
rect 87 56 88 57
rect 86 56 87 57
rect 85 56 86 57
rect 84 56 85 57
rect 83 56 84 57
rect 82 56 83 57
rect 399 57 400 58
rect 398 57 399 58
rect 397 57 398 58
rect 97 57 98 58
rect 96 57 97 58
rect 95 57 96 58
rect 94 57 95 58
rect 93 57 94 58
rect 92 57 93 58
rect 91 57 92 58
rect 90 57 91 58
rect 89 57 90 58
rect 88 57 89 58
rect 87 57 88 58
rect 86 57 87 58
rect 85 57 86 58
rect 84 57 85 58
rect 83 57 84 58
rect 82 57 83 58
rect 81 57 82 58
rect 400 58 401 59
rect 399 58 400 59
rect 398 58 399 59
rect 397 58 398 59
rect 109 58 110 59
rect 96 58 97 59
rect 95 58 96 59
rect 94 58 95 59
rect 93 58 94 59
rect 92 58 93 59
rect 91 58 92 59
rect 90 58 91 59
rect 89 58 90 59
rect 88 58 89 59
rect 87 58 88 59
rect 86 58 87 59
rect 85 58 86 59
rect 84 58 85 59
rect 83 58 84 59
rect 82 58 83 59
rect 81 58 82 59
rect 80 58 81 59
rect 401 59 402 60
rect 400 59 401 60
rect 399 59 400 60
rect 398 59 399 60
rect 397 59 398 60
rect 112 59 113 60
rect 111 59 112 60
rect 110 59 111 60
rect 109 59 110 60
rect 108 59 109 60
rect 107 59 108 60
rect 106 59 107 60
rect 96 59 97 60
rect 95 59 96 60
rect 94 59 95 60
rect 93 59 94 60
rect 92 59 93 60
rect 91 59 92 60
rect 90 59 91 60
rect 89 59 90 60
rect 88 59 89 60
rect 87 59 88 60
rect 86 59 87 60
rect 85 59 86 60
rect 84 59 85 60
rect 83 59 84 60
rect 82 59 83 60
rect 81 59 82 60
rect 80 59 81 60
rect 402 60 403 61
rect 401 60 402 61
rect 400 60 401 61
rect 399 60 400 61
rect 398 60 399 61
rect 397 60 398 61
rect 114 60 115 61
rect 113 60 114 61
rect 112 60 113 61
rect 111 60 112 61
rect 110 60 111 61
rect 109 60 110 61
rect 108 60 109 61
rect 107 60 108 61
rect 106 60 107 61
rect 105 60 106 61
rect 104 60 105 61
rect 96 60 97 61
rect 95 60 96 61
rect 94 60 95 61
rect 93 60 94 61
rect 92 60 93 61
rect 91 60 92 61
rect 90 60 91 61
rect 89 60 90 61
rect 88 60 89 61
rect 87 60 88 61
rect 86 60 87 61
rect 85 60 86 61
rect 84 60 85 61
rect 83 60 84 61
rect 82 60 83 61
rect 81 60 82 61
rect 80 60 81 61
rect 79 60 80 61
rect 404 61 405 62
rect 403 61 404 62
rect 402 61 403 62
rect 401 61 402 62
rect 400 61 401 62
rect 399 61 400 62
rect 398 61 399 62
rect 397 61 398 62
rect 116 61 117 62
rect 115 61 116 62
rect 114 61 115 62
rect 113 61 114 62
rect 112 61 113 62
rect 111 61 112 62
rect 110 61 111 62
rect 109 61 110 62
rect 108 61 109 62
rect 107 61 108 62
rect 106 61 107 62
rect 105 61 106 62
rect 104 61 105 62
rect 103 61 104 62
rect 96 61 97 62
rect 95 61 96 62
rect 94 61 95 62
rect 93 61 94 62
rect 92 61 93 62
rect 91 61 92 62
rect 90 61 91 62
rect 89 61 90 62
rect 88 61 89 62
rect 87 61 88 62
rect 86 61 87 62
rect 85 61 86 62
rect 84 61 85 62
rect 83 61 84 62
rect 82 61 83 62
rect 81 61 82 62
rect 80 61 81 62
rect 79 61 80 62
rect 78 61 79 62
rect 406 62 407 63
rect 405 62 406 63
rect 404 62 405 63
rect 403 62 404 63
rect 402 62 403 63
rect 401 62 402 63
rect 400 62 401 63
rect 399 62 400 63
rect 398 62 399 63
rect 397 62 398 63
rect 118 62 119 63
rect 117 62 118 63
rect 116 62 117 63
rect 115 62 116 63
rect 114 62 115 63
rect 113 62 114 63
rect 112 62 113 63
rect 111 62 112 63
rect 110 62 111 63
rect 109 62 110 63
rect 108 62 109 63
rect 107 62 108 63
rect 106 62 107 63
rect 105 62 106 63
rect 104 62 105 63
rect 103 62 104 63
rect 102 62 103 63
rect 95 62 96 63
rect 94 62 95 63
rect 93 62 94 63
rect 92 62 93 63
rect 91 62 92 63
rect 90 62 91 63
rect 89 62 90 63
rect 88 62 89 63
rect 87 62 88 63
rect 86 62 87 63
rect 85 62 86 63
rect 84 62 85 63
rect 83 62 84 63
rect 82 62 83 63
rect 81 62 82 63
rect 80 62 81 63
rect 79 62 80 63
rect 78 62 79 63
rect 407 63 408 64
rect 406 63 407 64
rect 405 63 406 64
rect 404 63 405 64
rect 403 63 404 64
rect 402 63 403 64
rect 401 63 402 64
rect 400 63 401 64
rect 399 63 400 64
rect 398 63 399 64
rect 397 63 398 64
rect 119 63 120 64
rect 118 63 119 64
rect 117 63 118 64
rect 116 63 117 64
rect 115 63 116 64
rect 114 63 115 64
rect 113 63 114 64
rect 112 63 113 64
rect 111 63 112 64
rect 110 63 111 64
rect 109 63 110 64
rect 108 63 109 64
rect 107 63 108 64
rect 106 63 107 64
rect 105 63 106 64
rect 104 63 105 64
rect 103 63 104 64
rect 102 63 103 64
rect 101 63 102 64
rect 95 63 96 64
rect 94 63 95 64
rect 93 63 94 64
rect 92 63 93 64
rect 91 63 92 64
rect 90 63 91 64
rect 89 63 90 64
rect 88 63 89 64
rect 87 63 88 64
rect 86 63 87 64
rect 85 63 86 64
rect 84 63 85 64
rect 83 63 84 64
rect 82 63 83 64
rect 81 63 82 64
rect 80 63 81 64
rect 79 63 80 64
rect 78 63 79 64
rect 77 63 78 64
rect 409 64 410 65
rect 408 64 409 65
rect 407 64 408 65
rect 406 64 407 65
rect 405 64 406 65
rect 404 64 405 65
rect 403 64 404 65
rect 402 64 403 65
rect 401 64 402 65
rect 400 64 401 65
rect 399 64 400 65
rect 398 64 399 65
rect 397 64 398 65
rect 120 64 121 65
rect 119 64 120 65
rect 118 64 119 65
rect 117 64 118 65
rect 116 64 117 65
rect 115 64 116 65
rect 114 64 115 65
rect 113 64 114 65
rect 112 64 113 65
rect 111 64 112 65
rect 110 64 111 65
rect 109 64 110 65
rect 108 64 109 65
rect 107 64 108 65
rect 106 64 107 65
rect 105 64 106 65
rect 104 64 105 65
rect 103 64 104 65
rect 102 64 103 65
rect 101 64 102 65
rect 100 64 101 65
rect 95 64 96 65
rect 94 64 95 65
rect 93 64 94 65
rect 92 64 93 65
rect 91 64 92 65
rect 90 64 91 65
rect 89 64 90 65
rect 88 64 89 65
rect 87 64 88 65
rect 86 64 87 65
rect 85 64 86 65
rect 84 64 85 65
rect 83 64 84 65
rect 82 64 83 65
rect 81 64 82 65
rect 80 64 81 65
rect 79 64 80 65
rect 78 64 79 65
rect 77 64 78 65
rect 441 65 442 66
rect 440 65 441 66
rect 411 65 412 66
rect 410 65 411 66
rect 409 65 410 66
rect 408 65 409 66
rect 407 65 408 66
rect 406 65 407 66
rect 405 65 406 66
rect 404 65 405 66
rect 403 65 404 66
rect 402 65 403 66
rect 401 65 402 66
rect 400 65 401 66
rect 399 65 400 66
rect 398 65 399 66
rect 397 65 398 66
rect 121 65 122 66
rect 120 65 121 66
rect 119 65 120 66
rect 118 65 119 66
rect 117 65 118 66
rect 116 65 117 66
rect 115 65 116 66
rect 114 65 115 66
rect 113 65 114 66
rect 112 65 113 66
rect 111 65 112 66
rect 110 65 111 66
rect 109 65 110 66
rect 108 65 109 66
rect 107 65 108 66
rect 106 65 107 66
rect 105 65 106 66
rect 104 65 105 66
rect 103 65 104 66
rect 102 65 103 66
rect 101 65 102 66
rect 100 65 101 66
rect 99 65 100 66
rect 94 65 95 66
rect 93 65 94 66
rect 92 65 93 66
rect 91 65 92 66
rect 90 65 91 66
rect 89 65 90 66
rect 88 65 89 66
rect 87 65 88 66
rect 86 65 87 66
rect 85 65 86 66
rect 84 65 85 66
rect 83 65 84 66
rect 82 65 83 66
rect 81 65 82 66
rect 80 65 81 66
rect 79 65 80 66
rect 78 65 79 66
rect 77 65 78 66
rect 76 65 77 66
rect 441 66 442 67
rect 440 66 441 67
rect 439 66 440 67
rect 413 66 414 67
rect 412 66 413 67
rect 411 66 412 67
rect 410 66 411 67
rect 409 66 410 67
rect 408 66 409 67
rect 407 66 408 67
rect 406 66 407 67
rect 405 66 406 67
rect 404 66 405 67
rect 403 66 404 67
rect 402 66 403 67
rect 401 66 402 67
rect 400 66 401 67
rect 399 66 400 67
rect 398 66 399 67
rect 397 66 398 67
rect 122 66 123 67
rect 121 66 122 67
rect 120 66 121 67
rect 119 66 120 67
rect 118 66 119 67
rect 117 66 118 67
rect 116 66 117 67
rect 115 66 116 67
rect 114 66 115 67
rect 113 66 114 67
rect 112 66 113 67
rect 111 66 112 67
rect 110 66 111 67
rect 109 66 110 67
rect 108 66 109 67
rect 107 66 108 67
rect 106 66 107 67
rect 105 66 106 67
rect 104 66 105 67
rect 103 66 104 67
rect 102 66 103 67
rect 101 66 102 67
rect 100 66 101 67
rect 99 66 100 67
rect 98 66 99 67
rect 94 66 95 67
rect 93 66 94 67
rect 92 66 93 67
rect 91 66 92 67
rect 90 66 91 67
rect 89 66 90 67
rect 88 66 89 67
rect 87 66 88 67
rect 86 66 87 67
rect 85 66 86 67
rect 84 66 85 67
rect 83 66 84 67
rect 82 66 83 67
rect 81 66 82 67
rect 80 66 81 67
rect 79 66 80 67
rect 78 66 79 67
rect 77 66 78 67
rect 76 66 77 67
rect 75 66 76 67
rect 441 67 442 68
rect 440 67 441 68
rect 439 67 440 68
rect 414 67 415 68
rect 413 67 414 68
rect 412 67 413 68
rect 411 67 412 68
rect 410 67 411 68
rect 409 67 410 68
rect 408 67 409 68
rect 407 67 408 68
rect 406 67 407 68
rect 405 67 406 68
rect 404 67 405 68
rect 403 67 404 68
rect 402 67 403 68
rect 401 67 402 68
rect 400 67 401 68
rect 399 67 400 68
rect 398 67 399 68
rect 397 67 398 68
rect 123 67 124 68
rect 122 67 123 68
rect 121 67 122 68
rect 120 67 121 68
rect 119 67 120 68
rect 118 67 119 68
rect 117 67 118 68
rect 116 67 117 68
rect 115 67 116 68
rect 114 67 115 68
rect 113 67 114 68
rect 112 67 113 68
rect 111 67 112 68
rect 110 67 111 68
rect 109 67 110 68
rect 108 67 109 68
rect 107 67 108 68
rect 106 67 107 68
rect 105 67 106 68
rect 104 67 105 68
rect 103 67 104 68
rect 102 67 103 68
rect 101 67 102 68
rect 100 67 101 68
rect 99 67 100 68
rect 98 67 99 68
rect 97 67 98 68
rect 93 67 94 68
rect 92 67 93 68
rect 91 67 92 68
rect 90 67 91 68
rect 89 67 90 68
rect 88 67 89 68
rect 87 67 88 68
rect 86 67 87 68
rect 85 67 86 68
rect 84 67 85 68
rect 83 67 84 68
rect 82 67 83 68
rect 81 67 82 68
rect 80 67 81 68
rect 79 67 80 68
rect 78 67 79 68
rect 77 67 78 68
rect 76 67 77 68
rect 75 67 76 68
rect 441 68 442 69
rect 440 68 441 69
rect 439 68 440 69
rect 416 68 417 69
rect 415 68 416 69
rect 414 68 415 69
rect 413 68 414 69
rect 412 68 413 69
rect 411 68 412 69
rect 410 68 411 69
rect 409 68 410 69
rect 408 68 409 69
rect 407 68 408 69
rect 406 68 407 69
rect 405 68 406 69
rect 404 68 405 69
rect 403 68 404 69
rect 402 68 403 69
rect 401 68 402 69
rect 400 68 401 69
rect 399 68 400 69
rect 398 68 399 69
rect 397 68 398 69
rect 124 68 125 69
rect 123 68 124 69
rect 122 68 123 69
rect 121 68 122 69
rect 120 68 121 69
rect 119 68 120 69
rect 118 68 119 69
rect 117 68 118 69
rect 116 68 117 69
rect 115 68 116 69
rect 114 68 115 69
rect 113 68 114 69
rect 112 68 113 69
rect 111 68 112 69
rect 110 68 111 69
rect 109 68 110 69
rect 108 68 109 69
rect 107 68 108 69
rect 106 68 107 69
rect 105 68 106 69
rect 104 68 105 69
rect 103 68 104 69
rect 102 68 103 69
rect 101 68 102 69
rect 100 68 101 69
rect 99 68 100 69
rect 98 68 99 69
rect 97 68 98 69
rect 96 68 97 69
rect 93 68 94 69
rect 92 68 93 69
rect 91 68 92 69
rect 90 68 91 69
rect 89 68 90 69
rect 88 68 89 69
rect 87 68 88 69
rect 86 68 87 69
rect 85 68 86 69
rect 84 68 85 69
rect 83 68 84 69
rect 82 68 83 69
rect 81 68 82 69
rect 80 68 81 69
rect 79 68 80 69
rect 78 68 79 69
rect 77 68 78 69
rect 76 68 77 69
rect 75 68 76 69
rect 74 68 75 69
rect 441 69 442 70
rect 440 69 441 70
rect 439 69 440 70
rect 418 69 419 70
rect 417 69 418 70
rect 416 69 417 70
rect 415 69 416 70
rect 414 69 415 70
rect 413 69 414 70
rect 412 69 413 70
rect 411 69 412 70
rect 410 69 411 70
rect 409 69 410 70
rect 408 69 409 70
rect 407 69 408 70
rect 406 69 407 70
rect 405 69 406 70
rect 404 69 405 70
rect 403 69 404 70
rect 402 69 403 70
rect 401 69 402 70
rect 400 69 401 70
rect 399 69 400 70
rect 398 69 399 70
rect 397 69 398 70
rect 125 69 126 70
rect 124 69 125 70
rect 123 69 124 70
rect 122 69 123 70
rect 121 69 122 70
rect 120 69 121 70
rect 119 69 120 70
rect 118 69 119 70
rect 117 69 118 70
rect 116 69 117 70
rect 115 69 116 70
rect 114 69 115 70
rect 113 69 114 70
rect 112 69 113 70
rect 111 69 112 70
rect 110 69 111 70
rect 109 69 110 70
rect 108 69 109 70
rect 107 69 108 70
rect 106 69 107 70
rect 105 69 106 70
rect 104 69 105 70
rect 103 69 104 70
rect 102 69 103 70
rect 101 69 102 70
rect 100 69 101 70
rect 99 69 100 70
rect 98 69 99 70
rect 97 69 98 70
rect 96 69 97 70
rect 95 69 96 70
rect 92 69 93 70
rect 91 69 92 70
rect 90 69 91 70
rect 89 69 90 70
rect 88 69 89 70
rect 87 69 88 70
rect 86 69 87 70
rect 85 69 86 70
rect 84 69 85 70
rect 83 69 84 70
rect 82 69 83 70
rect 81 69 82 70
rect 80 69 81 70
rect 79 69 80 70
rect 78 69 79 70
rect 77 69 78 70
rect 76 69 77 70
rect 75 69 76 70
rect 74 69 75 70
rect 441 70 442 71
rect 440 70 441 71
rect 439 70 440 71
rect 438 70 439 71
rect 420 70 421 71
rect 419 70 420 71
rect 418 70 419 71
rect 417 70 418 71
rect 416 70 417 71
rect 415 70 416 71
rect 414 70 415 71
rect 413 70 414 71
rect 412 70 413 71
rect 411 70 412 71
rect 410 70 411 71
rect 409 70 410 71
rect 408 70 409 71
rect 407 70 408 71
rect 406 70 407 71
rect 405 70 406 71
rect 404 70 405 71
rect 403 70 404 71
rect 402 70 403 71
rect 400 70 401 71
rect 399 70 400 71
rect 398 70 399 71
rect 397 70 398 71
rect 125 70 126 71
rect 124 70 125 71
rect 123 70 124 71
rect 122 70 123 71
rect 121 70 122 71
rect 120 70 121 71
rect 119 70 120 71
rect 118 70 119 71
rect 117 70 118 71
rect 116 70 117 71
rect 115 70 116 71
rect 114 70 115 71
rect 113 70 114 71
rect 112 70 113 71
rect 111 70 112 71
rect 110 70 111 71
rect 109 70 110 71
rect 108 70 109 71
rect 107 70 108 71
rect 106 70 107 71
rect 105 70 106 71
rect 104 70 105 71
rect 103 70 104 71
rect 102 70 103 71
rect 101 70 102 71
rect 100 70 101 71
rect 99 70 100 71
rect 98 70 99 71
rect 97 70 98 71
rect 96 70 97 71
rect 95 70 96 71
rect 94 70 95 71
rect 92 70 93 71
rect 91 70 92 71
rect 90 70 91 71
rect 89 70 90 71
rect 88 70 89 71
rect 87 70 88 71
rect 86 70 87 71
rect 85 70 86 71
rect 84 70 85 71
rect 83 70 84 71
rect 82 70 83 71
rect 81 70 82 71
rect 80 70 81 71
rect 79 70 80 71
rect 78 70 79 71
rect 77 70 78 71
rect 76 70 77 71
rect 75 70 76 71
rect 74 70 75 71
rect 441 71 442 72
rect 440 71 441 72
rect 439 71 440 72
rect 438 71 439 72
rect 437 71 438 72
rect 436 71 437 72
rect 435 71 436 72
rect 434 71 435 72
rect 433 71 434 72
rect 432 71 433 72
rect 431 71 432 72
rect 430 71 431 72
rect 429 71 430 72
rect 428 71 429 72
rect 427 71 428 72
rect 426 71 427 72
rect 425 71 426 72
rect 424 71 425 72
rect 423 71 424 72
rect 422 71 423 72
rect 421 71 422 72
rect 420 71 421 72
rect 419 71 420 72
rect 418 71 419 72
rect 417 71 418 72
rect 416 71 417 72
rect 415 71 416 72
rect 414 71 415 72
rect 413 71 414 72
rect 412 71 413 72
rect 411 71 412 72
rect 410 71 411 72
rect 409 71 410 72
rect 408 71 409 72
rect 407 71 408 72
rect 406 71 407 72
rect 405 71 406 72
rect 404 71 405 72
rect 399 71 400 72
rect 398 71 399 72
rect 397 71 398 72
rect 126 71 127 72
rect 125 71 126 72
rect 124 71 125 72
rect 123 71 124 72
rect 122 71 123 72
rect 121 71 122 72
rect 120 71 121 72
rect 119 71 120 72
rect 118 71 119 72
rect 117 71 118 72
rect 116 71 117 72
rect 115 71 116 72
rect 114 71 115 72
rect 113 71 114 72
rect 112 71 113 72
rect 111 71 112 72
rect 110 71 111 72
rect 109 71 110 72
rect 108 71 109 72
rect 107 71 108 72
rect 106 71 107 72
rect 105 71 106 72
rect 104 71 105 72
rect 103 71 104 72
rect 102 71 103 72
rect 101 71 102 72
rect 100 71 101 72
rect 99 71 100 72
rect 98 71 99 72
rect 97 71 98 72
rect 96 71 97 72
rect 95 71 96 72
rect 94 71 95 72
rect 93 71 94 72
rect 91 71 92 72
rect 90 71 91 72
rect 89 71 90 72
rect 88 71 89 72
rect 87 71 88 72
rect 86 71 87 72
rect 85 71 86 72
rect 84 71 85 72
rect 83 71 84 72
rect 82 71 83 72
rect 81 71 82 72
rect 80 71 81 72
rect 79 71 80 72
rect 78 71 79 72
rect 77 71 78 72
rect 76 71 77 72
rect 75 71 76 72
rect 74 71 75 72
rect 73 71 74 72
rect 441 72 442 73
rect 440 72 441 73
rect 439 72 440 73
rect 438 72 439 73
rect 437 72 438 73
rect 436 72 437 73
rect 435 72 436 73
rect 434 72 435 73
rect 433 72 434 73
rect 432 72 433 73
rect 431 72 432 73
rect 430 72 431 73
rect 429 72 430 73
rect 428 72 429 73
rect 427 72 428 73
rect 426 72 427 73
rect 425 72 426 73
rect 424 72 425 73
rect 423 72 424 73
rect 422 72 423 73
rect 421 72 422 73
rect 420 72 421 73
rect 419 72 420 73
rect 418 72 419 73
rect 417 72 418 73
rect 416 72 417 73
rect 415 72 416 73
rect 414 72 415 73
rect 413 72 414 73
rect 412 72 413 73
rect 411 72 412 73
rect 410 72 411 73
rect 409 72 410 73
rect 408 72 409 73
rect 407 72 408 73
rect 406 72 407 73
rect 399 72 400 73
rect 398 72 399 73
rect 397 72 398 73
rect 126 72 127 73
rect 125 72 126 73
rect 124 72 125 73
rect 123 72 124 73
rect 122 72 123 73
rect 121 72 122 73
rect 120 72 121 73
rect 119 72 120 73
rect 118 72 119 73
rect 117 72 118 73
rect 116 72 117 73
rect 115 72 116 73
rect 114 72 115 73
rect 113 72 114 73
rect 112 72 113 73
rect 111 72 112 73
rect 110 72 111 73
rect 109 72 110 73
rect 108 72 109 73
rect 107 72 108 73
rect 106 72 107 73
rect 105 72 106 73
rect 104 72 105 73
rect 103 72 104 73
rect 102 72 103 73
rect 101 72 102 73
rect 100 72 101 73
rect 99 72 100 73
rect 98 72 99 73
rect 97 72 98 73
rect 96 72 97 73
rect 95 72 96 73
rect 94 72 95 73
rect 93 72 94 73
rect 92 72 93 73
rect 91 72 92 73
rect 90 72 91 73
rect 89 72 90 73
rect 88 72 89 73
rect 87 72 88 73
rect 86 72 87 73
rect 85 72 86 73
rect 84 72 85 73
rect 83 72 84 73
rect 82 72 83 73
rect 81 72 82 73
rect 80 72 81 73
rect 79 72 80 73
rect 78 72 79 73
rect 77 72 78 73
rect 76 72 77 73
rect 75 72 76 73
rect 74 72 75 73
rect 73 72 74 73
rect 441 73 442 74
rect 440 73 441 74
rect 439 73 440 74
rect 438 73 439 74
rect 437 73 438 74
rect 436 73 437 74
rect 435 73 436 74
rect 434 73 435 74
rect 433 73 434 74
rect 432 73 433 74
rect 431 73 432 74
rect 430 73 431 74
rect 429 73 430 74
rect 428 73 429 74
rect 427 73 428 74
rect 426 73 427 74
rect 425 73 426 74
rect 424 73 425 74
rect 423 73 424 74
rect 422 73 423 74
rect 421 73 422 74
rect 420 73 421 74
rect 419 73 420 74
rect 418 73 419 74
rect 417 73 418 74
rect 416 73 417 74
rect 415 73 416 74
rect 414 73 415 74
rect 413 73 414 74
rect 412 73 413 74
rect 411 73 412 74
rect 410 73 411 74
rect 409 73 410 74
rect 408 73 409 74
rect 399 73 400 74
rect 398 73 399 74
rect 397 73 398 74
rect 141 73 142 74
rect 140 73 141 74
rect 139 73 140 74
rect 138 73 139 74
rect 137 73 138 74
rect 136 73 137 74
rect 126 73 127 74
rect 125 73 126 74
rect 124 73 125 74
rect 123 73 124 74
rect 122 73 123 74
rect 121 73 122 74
rect 120 73 121 74
rect 119 73 120 74
rect 118 73 119 74
rect 117 73 118 74
rect 116 73 117 74
rect 115 73 116 74
rect 114 73 115 74
rect 113 73 114 74
rect 112 73 113 74
rect 111 73 112 74
rect 110 73 111 74
rect 109 73 110 74
rect 108 73 109 74
rect 107 73 108 74
rect 106 73 107 74
rect 105 73 106 74
rect 104 73 105 74
rect 103 73 104 74
rect 102 73 103 74
rect 101 73 102 74
rect 100 73 101 74
rect 99 73 100 74
rect 98 73 99 74
rect 97 73 98 74
rect 96 73 97 74
rect 95 73 96 74
rect 94 73 95 74
rect 93 73 94 74
rect 92 73 93 74
rect 91 73 92 74
rect 90 73 91 74
rect 89 73 90 74
rect 88 73 89 74
rect 87 73 88 74
rect 86 73 87 74
rect 85 73 86 74
rect 84 73 85 74
rect 83 73 84 74
rect 82 73 83 74
rect 81 73 82 74
rect 80 73 81 74
rect 79 73 80 74
rect 78 73 79 74
rect 77 73 78 74
rect 76 73 77 74
rect 75 73 76 74
rect 74 73 75 74
rect 73 73 74 74
rect 72 73 73 74
rect 441 74 442 75
rect 440 74 441 75
rect 439 74 440 75
rect 438 74 439 75
rect 437 74 438 75
rect 436 74 437 75
rect 435 74 436 75
rect 434 74 435 75
rect 433 74 434 75
rect 432 74 433 75
rect 431 74 432 75
rect 430 74 431 75
rect 429 74 430 75
rect 428 74 429 75
rect 427 74 428 75
rect 426 74 427 75
rect 425 74 426 75
rect 424 74 425 75
rect 423 74 424 75
rect 422 74 423 75
rect 421 74 422 75
rect 420 74 421 75
rect 419 74 420 75
rect 418 74 419 75
rect 417 74 418 75
rect 416 74 417 75
rect 415 74 416 75
rect 414 74 415 75
rect 413 74 414 75
rect 412 74 413 75
rect 411 74 412 75
rect 410 74 411 75
rect 144 74 145 75
rect 143 74 144 75
rect 142 74 143 75
rect 141 74 142 75
rect 140 74 141 75
rect 139 74 140 75
rect 138 74 139 75
rect 137 74 138 75
rect 136 74 137 75
rect 135 74 136 75
rect 134 74 135 75
rect 126 74 127 75
rect 125 74 126 75
rect 124 74 125 75
rect 123 74 124 75
rect 122 74 123 75
rect 121 74 122 75
rect 120 74 121 75
rect 119 74 120 75
rect 118 74 119 75
rect 117 74 118 75
rect 116 74 117 75
rect 115 74 116 75
rect 114 74 115 75
rect 113 74 114 75
rect 112 74 113 75
rect 111 74 112 75
rect 110 74 111 75
rect 109 74 110 75
rect 108 74 109 75
rect 107 74 108 75
rect 106 74 107 75
rect 105 74 106 75
rect 104 74 105 75
rect 103 74 104 75
rect 102 74 103 75
rect 101 74 102 75
rect 100 74 101 75
rect 99 74 100 75
rect 98 74 99 75
rect 97 74 98 75
rect 96 74 97 75
rect 95 74 96 75
rect 94 74 95 75
rect 93 74 94 75
rect 92 74 93 75
rect 91 74 92 75
rect 90 74 91 75
rect 89 74 90 75
rect 88 74 89 75
rect 87 74 88 75
rect 86 74 87 75
rect 85 74 86 75
rect 84 74 85 75
rect 83 74 84 75
rect 82 74 83 75
rect 81 74 82 75
rect 80 74 81 75
rect 79 74 80 75
rect 78 74 79 75
rect 77 74 78 75
rect 76 74 77 75
rect 75 74 76 75
rect 74 74 75 75
rect 73 74 74 75
rect 72 74 73 75
rect 441 75 442 76
rect 440 75 441 76
rect 439 75 440 76
rect 438 75 439 76
rect 437 75 438 76
rect 436 75 437 76
rect 435 75 436 76
rect 434 75 435 76
rect 433 75 434 76
rect 432 75 433 76
rect 431 75 432 76
rect 430 75 431 76
rect 429 75 430 76
rect 428 75 429 76
rect 427 75 428 76
rect 426 75 427 76
rect 425 75 426 76
rect 424 75 425 76
rect 423 75 424 76
rect 422 75 423 76
rect 421 75 422 76
rect 420 75 421 76
rect 419 75 420 76
rect 418 75 419 76
rect 417 75 418 76
rect 416 75 417 76
rect 415 75 416 76
rect 414 75 415 76
rect 413 75 414 76
rect 412 75 413 76
rect 146 75 147 76
rect 145 75 146 76
rect 144 75 145 76
rect 143 75 144 76
rect 142 75 143 76
rect 141 75 142 76
rect 140 75 141 76
rect 139 75 140 76
rect 138 75 139 76
rect 137 75 138 76
rect 136 75 137 76
rect 135 75 136 76
rect 134 75 135 76
rect 126 75 127 76
rect 125 75 126 76
rect 124 75 125 76
rect 123 75 124 76
rect 122 75 123 76
rect 121 75 122 76
rect 120 75 121 76
rect 119 75 120 76
rect 118 75 119 76
rect 117 75 118 76
rect 116 75 117 76
rect 115 75 116 76
rect 114 75 115 76
rect 113 75 114 76
rect 112 75 113 76
rect 111 75 112 76
rect 110 75 111 76
rect 109 75 110 76
rect 108 75 109 76
rect 107 75 108 76
rect 106 75 107 76
rect 105 75 106 76
rect 104 75 105 76
rect 103 75 104 76
rect 102 75 103 76
rect 101 75 102 76
rect 100 75 101 76
rect 99 75 100 76
rect 98 75 99 76
rect 97 75 98 76
rect 96 75 97 76
rect 95 75 96 76
rect 94 75 95 76
rect 93 75 94 76
rect 92 75 93 76
rect 91 75 92 76
rect 90 75 91 76
rect 89 75 90 76
rect 88 75 89 76
rect 87 75 88 76
rect 86 75 87 76
rect 85 75 86 76
rect 84 75 85 76
rect 83 75 84 76
rect 82 75 83 76
rect 81 75 82 76
rect 80 75 81 76
rect 79 75 80 76
rect 78 75 79 76
rect 77 75 78 76
rect 76 75 77 76
rect 75 75 76 76
rect 74 75 75 76
rect 73 75 74 76
rect 72 75 73 76
rect 71 75 72 76
rect 441 76 442 77
rect 440 76 441 77
rect 439 76 440 77
rect 438 76 439 77
rect 437 76 438 77
rect 436 76 437 77
rect 435 76 436 77
rect 434 76 435 77
rect 433 76 434 77
rect 432 76 433 77
rect 431 76 432 77
rect 430 76 431 77
rect 429 76 430 77
rect 428 76 429 77
rect 427 76 428 77
rect 426 76 427 77
rect 425 76 426 77
rect 424 76 425 77
rect 423 76 424 77
rect 422 76 423 77
rect 421 76 422 77
rect 420 76 421 77
rect 419 76 420 77
rect 418 76 419 77
rect 417 76 418 77
rect 416 76 417 77
rect 415 76 416 77
rect 414 76 415 77
rect 148 76 149 77
rect 147 76 148 77
rect 146 76 147 77
rect 145 76 146 77
rect 144 76 145 77
rect 143 76 144 77
rect 142 76 143 77
rect 141 76 142 77
rect 140 76 141 77
rect 139 76 140 77
rect 138 76 139 77
rect 137 76 138 77
rect 136 76 137 77
rect 135 76 136 77
rect 134 76 135 77
rect 133 76 134 77
rect 127 76 128 77
rect 126 76 127 77
rect 125 76 126 77
rect 124 76 125 77
rect 123 76 124 77
rect 122 76 123 77
rect 121 76 122 77
rect 120 76 121 77
rect 119 76 120 77
rect 118 76 119 77
rect 117 76 118 77
rect 116 76 117 77
rect 115 76 116 77
rect 114 76 115 77
rect 113 76 114 77
rect 112 76 113 77
rect 111 76 112 77
rect 110 76 111 77
rect 109 76 110 77
rect 108 76 109 77
rect 107 76 108 77
rect 106 76 107 77
rect 105 76 106 77
rect 104 76 105 77
rect 103 76 104 77
rect 102 76 103 77
rect 101 76 102 77
rect 100 76 101 77
rect 99 76 100 77
rect 98 76 99 77
rect 97 76 98 77
rect 96 76 97 77
rect 95 76 96 77
rect 94 76 95 77
rect 93 76 94 77
rect 92 76 93 77
rect 91 76 92 77
rect 90 76 91 77
rect 89 76 90 77
rect 88 76 89 77
rect 87 76 88 77
rect 86 76 87 77
rect 85 76 86 77
rect 84 76 85 77
rect 83 76 84 77
rect 82 76 83 77
rect 81 76 82 77
rect 80 76 81 77
rect 79 76 80 77
rect 78 76 79 77
rect 77 76 78 77
rect 76 76 77 77
rect 75 76 76 77
rect 74 76 75 77
rect 73 76 74 77
rect 72 76 73 77
rect 71 76 72 77
rect 441 77 442 78
rect 440 77 441 78
rect 439 77 440 78
rect 438 77 439 78
rect 437 77 438 78
rect 436 77 437 78
rect 435 77 436 78
rect 434 77 435 78
rect 433 77 434 78
rect 432 77 433 78
rect 431 77 432 78
rect 430 77 431 78
rect 429 77 430 78
rect 428 77 429 78
rect 427 77 428 78
rect 426 77 427 78
rect 425 77 426 78
rect 424 77 425 78
rect 423 77 424 78
rect 422 77 423 78
rect 421 77 422 78
rect 420 77 421 78
rect 419 77 420 78
rect 418 77 419 78
rect 417 77 418 78
rect 416 77 417 78
rect 149 77 150 78
rect 148 77 149 78
rect 147 77 148 78
rect 146 77 147 78
rect 145 77 146 78
rect 144 77 145 78
rect 143 77 144 78
rect 142 77 143 78
rect 141 77 142 78
rect 140 77 141 78
rect 139 77 140 78
rect 138 77 139 78
rect 137 77 138 78
rect 136 77 137 78
rect 135 77 136 78
rect 134 77 135 78
rect 133 77 134 78
rect 126 77 127 78
rect 125 77 126 78
rect 124 77 125 78
rect 123 77 124 78
rect 122 77 123 78
rect 121 77 122 78
rect 120 77 121 78
rect 119 77 120 78
rect 118 77 119 78
rect 117 77 118 78
rect 116 77 117 78
rect 115 77 116 78
rect 114 77 115 78
rect 113 77 114 78
rect 112 77 113 78
rect 111 77 112 78
rect 110 77 111 78
rect 109 77 110 78
rect 108 77 109 78
rect 107 77 108 78
rect 106 77 107 78
rect 105 77 106 78
rect 104 77 105 78
rect 103 77 104 78
rect 102 77 103 78
rect 101 77 102 78
rect 100 77 101 78
rect 99 77 100 78
rect 98 77 99 78
rect 97 77 98 78
rect 96 77 97 78
rect 95 77 96 78
rect 94 77 95 78
rect 93 77 94 78
rect 92 77 93 78
rect 91 77 92 78
rect 90 77 91 78
rect 89 77 90 78
rect 88 77 89 78
rect 87 77 88 78
rect 86 77 87 78
rect 85 77 86 78
rect 84 77 85 78
rect 83 77 84 78
rect 82 77 83 78
rect 81 77 82 78
rect 80 77 81 78
rect 79 77 80 78
rect 78 77 79 78
rect 77 77 78 78
rect 76 77 77 78
rect 75 77 76 78
rect 74 77 75 78
rect 73 77 74 78
rect 72 77 73 78
rect 71 77 72 78
rect 70 77 71 78
rect 441 78 442 79
rect 440 78 441 79
rect 439 78 440 79
rect 438 78 439 79
rect 437 78 438 79
rect 436 78 437 79
rect 435 78 436 79
rect 434 78 435 79
rect 433 78 434 79
rect 432 78 433 79
rect 431 78 432 79
rect 430 78 431 79
rect 429 78 430 79
rect 428 78 429 79
rect 427 78 428 79
rect 426 78 427 79
rect 425 78 426 79
rect 424 78 425 79
rect 423 78 424 79
rect 422 78 423 79
rect 421 78 422 79
rect 420 78 421 79
rect 419 78 420 79
rect 418 78 419 79
rect 151 78 152 79
rect 150 78 151 79
rect 149 78 150 79
rect 148 78 149 79
rect 147 78 148 79
rect 146 78 147 79
rect 145 78 146 79
rect 144 78 145 79
rect 143 78 144 79
rect 142 78 143 79
rect 141 78 142 79
rect 140 78 141 79
rect 139 78 140 79
rect 138 78 139 79
rect 137 78 138 79
rect 136 78 137 79
rect 135 78 136 79
rect 134 78 135 79
rect 133 78 134 79
rect 126 78 127 79
rect 125 78 126 79
rect 124 78 125 79
rect 123 78 124 79
rect 122 78 123 79
rect 121 78 122 79
rect 120 78 121 79
rect 119 78 120 79
rect 118 78 119 79
rect 117 78 118 79
rect 116 78 117 79
rect 115 78 116 79
rect 114 78 115 79
rect 113 78 114 79
rect 112 78 113 79
rect 111 78 112 79
rect 110 78 111 79
rect 109 78 110 79
rect 108 78 109 79
rect 107 78 108 79
rect 106 78 107 79
rect 105 78 106 79
rect 104 78 105 79
rect 103 78 104 79
rect 102 78 103 79
rect 101 78 102 79
rect 100 78 101 79
rect 99 78 100 79
rect 98 78 99 79
rect 97 78 98 79
rect 96 78 97 79
rect 95 78 96 79
rect 94 78 95 79
rect 93 78 94 79
rect 92 78 93 79
rect 91 78 92 79
rect 90 78 91 79
rect 89 78 90 79
rect 88 78 89 79
rect 87 78 88 79
rect 86 78 87 79
rect 85 78 86 79
rect 84 78 85 79
rect 83 78 84 79
rect 82 78 83 79
rect 81 78 82 79
rect 80 78 81 79
rect 79 78 80 79
rect 78 78 79 79
rect 77 78 78 79
rect 76 78 77 79
rect 75 78 76 79
rect 74 78 75 79
rect 73 78 74 79
rect 72 78 73 79
rect 71 78 72 79
rect 70 78 71 79
rect 441 79 442 80
rect 440 79 441 80
rect 439 79 440 80
rect 438 79 439 80
rect 437 79 438 80
rect 436 79 437 80
rect 435 79 436 80
rect 434 79 435 80
rect 433 79 434 80
rect 432 79 433 80
rect 431 79 432 80
rect 430 79 431 80
rect 429 79 430 80
rect 428 79 429 80
rect 427 79 428 80
rect 426 79 427 80
rect 425 79 426 80
rect 424 79 425 80
rect 423 79 424 80
rect 422 79 423 80
rect 421 79 422 80
rect 420 79 421 80
rect 419 79 420 80
rect 418 79 419 80
rect 417 79 418 80
rect 152 79 153 80
rect 151 79 152 80
rect 150 79 151 80
rect 149 79 150 80
rect 148 79 149 80
rect 147 79 148 80
rect 146 79 147 80
rect 145 79 146 80
rect 144 79 145 80
rect 143 79 144 80
rect 142 79 143 80
rect 141 79 142 80
rect 140 79 141 80
rect 139 79 140 80
rect 138 79 139 80
rect 137 79 138 80
rect 136 79 137 80
rect 135 79 136 80
rect 134 79 135 80
rect 133 79 134 80
rect 126 79 127 80
rect 125 79 126 80
rect 124 79 125 80
rect 123 79 124 80
rect 122 79 123 80
rect 121 79 122 80
rect 120 79 121 80
rect 119 79 120 80
rect 118 79 119 80
rect 117 79 118 80
rect 116 79 117 80
rect 115 79 116 80
rect 114 79 115 80
rect 113 79 114 80
rect 112 79 113 80
rect 111 79 112 80
rect 110 79 111 80
rect 109 79 110 80
rect 108 79 109 80
rect 107 79 108 80
rect 106 79 107 80
rect 105 79 106 80
rect 104 79 105 80
rect 103 79 104 80
rect 102 79 103 80
rect 101 79 102 80
rect 100 79 101 80
rect 99 79 100 80
rect 98 79 99 80
rect 97 79 98 80
rect 96 79 97 80
rect 95 79 96 80
rect 94 79 95 80
rect 93 79 94 80
rect 92 79 93 80
rect 91 79 92 80
rect 90 79 91 80
rect 89 79 90 80
rect 88 79 89 80
rect 87 79 88 80
rect 86 79 87 80
rect 85 79 86 80
rect 84 79 85 80
rect 83 79 84 80
rect 82 79 83 80
rect 81 79 82 80
rect 80 79 81 80
rect 79 79 80 80
rect 78 79 79 80
rect 77 79 78 80
rect 76 79 77 80
rect 75 79 76 80
rect 74 79 75 80
rect 73 79 74 80
rect 72 79 73 80
rect 71 79 72 80
rect 70 79 71 80
rect 69 79 70 80
rect 441 80 442 81
rect 440 80 441 81
rect 439 80 440 81
rect 438 80 439 81
rect 437 80 438 81
rect 436 80 437 81
rect 435 80 436 81
rect 434 80 435 81
rect 433 80 434 81
rect 432 80 433 81
rect 431 80 432 81
rect 430 80 431 81
rect 429 80 430 81
rect 428 80 429 81
rect 427 80 428 81
rect 426 80 427 81
rect 425 80 426 81
rect 424 80 425 81
rect 423 80 424 81
rect 422 80 423 81
rect 421 80 422 81
rect 420 80 421 81
rect 419 80 420 81
rect 418 80 419 81
rect 417 80 418 81
rect 416 80 417 81
rect 415 80 416 81
rect 154 80 155 81
rect 153 80 154 81
rect 152 80 153 81
rect 151 80 152 81
rect 150 80 151 81
rect 149 80 150 81
rect 148 80 149 81
rect 147 80 148 81
rect 146 80 147 81
rect 145 80 146 81
rect 144 80 145 81
rect 143 80 144 81
rect 142 80 143 81
rect 141 80 142 81
rect 140 80 141 81
rect 139 80 140 81
rect 138 80 139 81
rect 137 80 138 81
rect 136 80 137 81
rect 135 80 136 81
rect 134 80 135 81
rect 133 80 134 81
rect 126 80 127 81
rect 125 80 126 81
rect 124 80 125 81
rect 123 80 124 81
rect 122 80 123 81
rect 121 80 122 81
rect 120 80 121 81
rect 119 80 120 81
rect 118 80 119 81
rect 117 80 118 81
rect 116 80 117 81
rect 115 80 116 81
rect 114 80 115 81
rect 113 80 114 81
rect 112 80 113 81
rect 111 80 112 81
rect 110 80 111 81
rect 109 80 110 81
rect 108 80 109 81
rect 107 80 108 81
rect 106 80 107 81
rect 105 80 106 81
rect 104 80 105 81
rect 103 80 104 81
rect 102 80 103 81
rect 101 80 102 81
rect 100 80 101 81
rect 99 80 100 81
rect 98 80 99 81
rect 97 80 98 81
rect 96 80 97 81
rect 95 80 96 81
rect 94 80 95 81
rect 93 80 94 81
rect 92 80 93 81
rect 91 80 92 81
rect 90 80 91 81
rect 89 80 90 81
rect 88 80 89 81
rect 87 80 88 81
rect 86 80 87 81
rect 85 80 86 81
rect 84 80 85 81
rect 83 80 84 81
rect 82 80 83 81
rect 81 80 82 81
rect 80 80 81 81
rect 79 80 80 81
rect 78 80 79 81
rect 77 80 78 81
rect 76 80 77 81
rect 75 80 76 81
rect 74 80 75 81
rect 73 80 74 81
rect 72 80 73 81
rect 71 80 72 81
rect 70 80 71 81
rect 69 80 70 81
rect 441 81 442 82
rect 440 81 441 82
rect 439 81 440 82
rect 438 81 439 82
rect 419 81 420 82
rect 418 81 419 82
rect 417 81 418 82
rect 416 81 417 82
rect 415 81 416 82
rect 414 81 415 82
rect 413 81 414 82
rect 156 81 157 82
rect 155 81 156 82
rect 154 81 155 82
rect 153 81 154 82
rect 152 81 153 82
rect 151 81 152 82
rect 150 81 151 82
rect 149 81 150 82
rect 148 81 149 82
rect 147 81 148 82
rect 146 81 147 82
rect 145 81 146 82
rect 144 81 145 82
rect 143 81 144 82
rect 142 81 143 82
rect 141 81 142 82
rect 140 81 141 82
rect 139 81 140 82
rect 138 81 139 82
rect 137 81 138 82
rect 136 81 137 82
rect 135 81 136 82
rect 134 81 135 82
rect 133 81 134 82
rect 126 81 127 82
rect 125 81 126 82
rect 124 81 125 82
rect 123 81 124 82
rect 122 81 123 82
rect 121 81 122 82
rect 120 81 121 82
rect 119 81 120 82
rect 118 81 119 82
rect 117 81 118 82
rect 116 81 117 82
rect 115 81 116 82
rect 114 81 115 82
rect 113 81 114 82
rect 112 81 113 82
rect 111 81 112 82
rect 110 81 111 82
rect 109 81 110 82
rect 108 81 109 82
rect 107 81 108 82
rect 106 81 107 82
rect 105 81 106 82
rect 104 81 105 82
rect 103 81 104 82
rect 102 81 103 82
rect 101 81 102 82
rect 100 81 101 82
rect 99 81 100 82
rect 98 81 99 82
rect 97 81 98 82
rect 96 81 97 82
rect 95 81 96 82
rect 94 81 95 82
rect 93 81 94 82
rect 92 81 93 82
rect 91 81 92 82
rect 90 81 91 82
rect 89 81 90 82
rect 88 81 89 82
rect 87 81 88 82
rect 86 81 87 82
rect 85 81 86 82
rect 84 81 85 82
rect 83 81 84 82
rect 82 81 83 82
rect 81 81 82 82
rect 80 81 81 82
rect 79 81 80 82
rect 78 81 79 82
rect 77 81 78 82
rect 76 81 77 82
rect 75 81 76 82
rect 74 81 75 82
rect 73 81 74 82
rect 72 81 73 82
rect 71 81 72 82
rect 70 81 71 82
rect 69 81 70 82
rect 68 81 69 82
rect 441 82 442 83
rect 440 82 441 83
rect 439 82 440 83
rect 417 82 418 83
rect 416 82 417 83
rect 415 82 416 83
rect 414 82 415 83
rect 413 82 414 83
rect 412 82 413 83
rect 411 82 412 83
rect 399 82 400 83
rect 398 82 399 83
rect 397 82 398 83
rect 159 82 160 83
rect 158 82 159 83
rect 157 82 158 83
rect 156 82 157 83
rect 155 82 156 83
rect 154 82 155 83
rect 153 82 154 83
rect 152 82 153 83
rect 151 82 152 83
rect 150 82 151 83
rect 149 82 150 83
rect 148 82 149 83
rect 147 82 148 83
rect 146 82 147 83
rect 145 82 146 83
rect 144 82 145 83
rect 143 82 144 83
rect 142 82 143 83
rect 141 82 142 83
rect 140 82 141 83
rect 139 82 140 83
rect 138 82 139 83
rect 137 82 138 83
rect 136 82 137 83
rect 135 82 136 83
rect 134 82 135 83
rect 133 82 134 83
rect 126 82 127 83
rect 125 82 126 83
rect 124 82 125 83
rect 123 82 124 83
rect 122 82 123 83
rect 121 82 122 83
rect 120 82 121 83
rect 119 82 120 83
rect 118 82 119 83
rect 117 82 118 83
rect 116 82 117 83
rect 115 82 116 83
rect 114 82 115 83
rect 113 82 114 83
rect 112 82 113 83
rect 111 82 112 83
rect 110 82 111 83
rect 109 82 110 83
rect 108 82 109 83
rect 107 82 108 83
rect 106 82 107 83
rect 105 82 106 83
rect 104 82 105 83
rect 103 82 104 83
rect 102 82 103 83
rect 101 82 102 83
rect 100 82 101 83
rect 99 82 100 83
rect 98 82 99 83
rect 97 82 98 83
rect 96 82 97 83
rect 95 82 96 83
rect 94 82 95 83
rect 93 82 94 83
rect 92 82 93 83
rect 91 82 92 83
rect 90 82 91 83
rect 89 82 90 83
rect 88 82 89 83
rect 87 82 88 83
rect 86 82 87 83
rect 85 82 86 83
rect 84 82 85 83
rect 83 82 84 83
rect 82 82 83 83
rect 81 82 82 83
rect 80 82 81 83
rect 79 82 80 83
rect 78 82 79 83
rect 77 82 78 83
rect 76 82 77 83
rect 75 82 76 83
rect 74 82 75 83
rect 73 82 74 83
rect 72 82 73 83
rect 71 82 72 83
rect 70 82 71 83
rect 69 82 70 83
rect 68 82 69 83
rect 67 82 68 83
rect 462 83 463 84
rect 441 83 442 84
rect 440 83 441 84
rect 439 83 440 84
rect 415 83 416 84
rect 414 83 415 84
rect 413 83 414 84
rect 412 83 413 84
rect 411 83 412 84
rect 410 83 411 84
rect 409 83 410 84
rect 399 83 400 84
rect 398 83 399 84
rect 397 83 398 84
rect 161 83 162 84
rect 160 83 161 84
rect 159 83 160 84
rect 158 83 159 84
rect 157 83 158 84
rect 156 83 157 84
rect 155 83 156 84
rect 154 83 155 84
rect 153 83 154 84
rect 152 83 153 84
rect 151 83 152 84
rect 150 83 151 84
rect 149 83 150 84
rect 148 83 149 84
rect 147 83 148 84
rect 146 83 147 84
rect 145 83 146 84
rect 144 83 145 84
rect 143 83 144 84
rect 142 83 143 84
rect 141 83 142 84
rect 140 83 141 84
rect 139 83 140 84
rect 138 83 139 84
rect 137 83 138 84
rect 136 83 137 84
rect 135 83 136 84
rect 134 83 135 84
rect 133 83 134 84
rect 126 83 127 84
rect 125 83 126 84
rect 124 83 125 84
rect 123 83 124 84
rect 122 83 123 84
rect 121 83 122 84
rect 120 83 121 84
rect 119 83 120 84
rect 118 83 119 84
rect 117 83 118 84
rect 116 83 117 84
rect 115 83 116 84
rect 114 83 115 84
rect 113 83 114 84
rect 112 83 113 84
rect 111 83 112 84
rect 110 83 111 84
rect 109 83 110 84
rect 108 83 109 84
rect 107 83 108 84
rect 106 83 107 84
rect 105 83 106 84
rect 104 83 105 84
rect 103 83 104 84
rect 102 83 103 84
rect 101 83 102 84
rect 100 83 101 84
rect 99 83 100 84
rect 98 83 99 84
rect 97 83 98 84
rect 96 83 97 84
rect 95 83 96 84
rect 94 83 95 84
rect 93 83 94 84
rect 92 83 93 84
rect 91 83 92 84
rect 90 83 91 84
rect 89 83 90 84
rect 88 83 89 84
rect 87 83 88 84
rect 86 83 87 84
rect 85 83 86 84
rect 84 83 85 84
rect 83 83 84 84
rect 82 83 83 84
rect 81 83 82 84
rect 80 83 81 84
rect 79 83 80 84
rect 78 83 79 84
rect 77 83 78 84
rect 76 83 77 84
rect 75 83 76 84
rect 74 83 75 84
rect 73 83 74 84
rect 72 83 73 84
rect 71 83 72 84
rect 70 83 71 84
rect 69 83 70 84
rect 68 83 69 84
rect 67 83 68 84
rect 462 84 463 85
rect 441 84 442 85
rect 440 84 441 85
rect 439 84 440 85
rect 413 84 414 85
rect 412 84 413 85
rect 411 84 412 85
rect 410 84 411 85
rect 409 84 410 85
rect 408 84 409 85
rect 407 84 408 85
rect 399 84 400 85
rect 398 84 399 85
rect 397 84 398 85
rect 163 84 164 85
rect 162 84 163 85
rect 161 84 162 85
rect 160 84 161 85
rect 159 84 160 85
rect 158 84 159 85
rect 157 84 158 85
rect 156 84 157 85
rect 155 84 156 85
rect 154 84 155 85
rect 153 84 154 85
rect 152 84 153 85
rect 151 84 152 85
rect 150 84 151 85
rect 149 84 150 85
rect 148 84 149 85
rect 147 84 148 85
rect 146 84 147 85
rect 145 84 146 85
rect 144 84 145 85
rect 143 84 144 85
rect 142 84 143 85
rect 141 84 142 85
rect 140 84 141 85
rect 139 84 140 85
rect 138 84 139 85
rect 137 84 138 85
rect 136 84 137 85
rect 135 84 136 85
rect 134 84 135 85
rect 133 84 134 85
rect 126 84 127 85
rect 125 84 126 85
rect 124 84 125 85
rect 123 84 124 85
rect 122 84 123 85
rect 121 84 122 85
rect 120 84 121 85
rect 119 84 120 85
rect 118 84 119 85
rect 117 84 118 85
rect 116 84 117 85
rect 115 84 116 85
rect 114 84 115 85
rect 113 84 114 85
rect 112 84 113 85
rect 111 84 112 85
rect 110 84 111 85
rect 109 84 110 85
rect 108 84 109 85
rect 107 84 108 85
rect 106 84 107 85
rect 105 84 106 85
rect 104 84 105 85
rect 103 84 104 85
rect 102 84 103 85
rect 101 84 102 85
rect 100 84 101 85
rect 99 84 100 85
rect 98 84 99 85
rect 97 84 98 85
rect 96 84 97 85
rect 95 84 96 85
rect 94 84 95 85
rect 93 84 94 85
rect 92 84 93 85
rect 91 84 92 85
rect 90 84 91 85
rect 89 84 90 85
rect 88 84 89 85
rect 87 84 88 85
rect 86 84 87 85
rect 85 84 86 85
rect 84 84 85 85
rect 83 84 84 85
rect 82 84 83 85
rect 81 84 82 85
rect 80 84 81 85
rect 79 84 80 85
rect 78 84 79 85
rect 77 84 78 85
rect 76 84 77 85
rect 75 84 76 85
rect 74 84 75 85
rect 73 84 74 85
rect 72 84 73 85
rect 71 84 72 85
rect 70 84 71 85
rect 69 84 70 85
rect 68 84 69 85
rect 67 84 68 85
rect 66 84 67 85
rect 463 85 464 86
rect 462 85 463 86
rect 441 85 442 86
rect 440 85 441 86
rect 439 85 440 86
rect 412 85 413 86
rect 411 85 412 86
rect 410 85 411 86
rect 409 85 410 86
rect 408 85 409 86
rect 407 85 408 86
rect 406 85 407 86
rect 405 85 406 86
rect 399 85 400 86
rect 398 85 399 86
rect 397 85 398 86
rect 227 85 228 86
rect 226 85 227 86
rect 225 85 226 86
rect 224 85 225 86
rect 223 85 224 86
rect 222 85 223 86
rect 221 85 222 86
rect 220 85 221 86
rect 219 85 220 86
rect 218 85 219 86
rect 217 85 218 86
rect 216 85 217 86
rect 215 85 216 86
rect 214 85 215 86
rect 213 85 214 86
rect 212 85 213 86
rect 211 85 212 86
rect 164 85 165 86
rect 163 85 164 86
rect 162 85 163 86
rect 161 85 162 86
rect 160 85 161 86
rect 159 85 160 86
rect 158 85 159 86
rect 157 85 158 86
rect 156 85 157 86
rect 155 85 156 86
rect 154 85 155 86
rect 153 85 154 86
rect 152 85 153 86
rect 151 85 152 86
rect 150 85 151 86
rect 149 85 150 86
rect 148 85 149 86
rect 147 85 148 86
rect 146 85 147 86
rect 145 85 146 86
rect 144 85 145 86
rect 143 85 144 86
rect 142 85 143 86
rect 141 85 142 86
rect 140 85 141 86
rect 139 85 140 86
rect 138 85 139 86
rect 137 85 138 86
rect 136 85 137 86
rect 135 85 136 86
rect 134 85 135 86
rect 133 85 134 86
rect 126 85 127 86
rect 125 85 126 86
rect 124 85 125 86
rect 123 85 124 86
rect 122 85 123 86
rect 121 85 122 86
rect 120 85 121 86
rect 119 85 120 86
rect 118 85 119 86
rect 117 85 118 86
rect 116 85 117 86
rect 115 85 116 86
rect 114 85 115 86
rect 113 85 114 86
rect 112 85 113 86
rect 111 85 112 86
rect 110 85 111 86
rect 109 85 110 86
rect 108 85 109 86
rect 107 85 108 86
rect 106 85 107 86
rect 105 85 106 86
rect 104 85 105 86
rect 103 85 104 86
rect 102 85 103 86
rect 101 85 102 86
rect 100 85 101 86
rect 99 85 100 86
rect 98 85 99 86
rect 97 85 98 86
rect 96 85 97 86
rect 95 85 96 86
rect 94 85 95 86
rect 93 85 94 86
rect 92 85 93 86
rect 91 85 92 86
rect 90 85 91 86
rect 89 85 90 86
rect 88 85 89 86
rect 87 85 88 86
rect 86 85 87 86
rect 85 85 86 86
rect 84 85 85 86
rect 83 85 84 86
rect 82 85 83 86
rect 81 85 82 86
rect 80 85 81 86
rect 79 85 80 86
rect 78 85 79 86
rect 77 85 78 86
rect 76 85 77 86
rect 75 85 76 86
rect 74 85 75 86
rect 73 85 74 86
rect 72 85 73 86
rect 71 85 72 86
rect 70 85 71 86
rect 69 85 70 86
rect 68 85 69 86
rect 67 85 68 86
rect 66 85 67 86
rect 478 86 479 87
rect 477 86 478 87
rect 476 86 477 87
rect 475 86 476 87
rect 474 86 475 87
rect 473 86 474 87
rect 472 86 473 87
rect 471 86 472 87
rect 470 86 471 87
rect 469 86 470 87
rect 468 86 469 87
rect 467 86 468 87
rect 466 86 467 87
rect 465 86 466 87
rect 464 86 465 87
rect 463 86 464 87
rect 462 86 463 87
rect 441 86 442 87
rect 440 86 441 87
rect 410 86 411 87
rect 409 86 410 87
rect 408 86 409 87
rect 407 86 408 87
rect 406 86 407 87
rect 405 86 406 87
rect 404 86 405 87
rect 403 86 404 87
rect 402 86 403 87
rect 401 86 402 87
rect 400 86 401 87
rect 399 86 400 87
rect 398 86 399 87
rect 397 86 398 87
rect 233 86 234 87
rect 232 86 233 87
rect 231 86 232 87
rect 230 86 231 87
rect 229 86 230 87
rect 228 86 229 87
rect 227 86 228 87
rect 226 86 227 87
rect 225 86 226 87
rect 224 86 225 87
rect 223 86 224 87
rect 222 86 223 87
rect 221 86 222 87
rect 220 86 221 87
rect 219 86 220 87
rect 218 86 219 87
rect 217 86 218 87
rect 216 86 217 87
rect 215 86 216 87
rect 214 86 215 87
rect 213 86 214 87
rect 212 86 213 87
rect 211 86 212 87
rect 210 86 211 87
rect 209 86 210 87
rect 208 86 209 87
rect 207 86 208 87
rect 206 86 207 87
rect 164 86 165 87
rect 163 86 164 87
rect 162 86 163 87
rect 161 86 162 87
rect 160 86 161 87
rect 159 86 160 87
rect 158 86 159 87
rect 157 86 158 87
rect 156 86 157 87
rect 155 86 156 87
rect 154 86 155 87
rect 153 86 154 87
rect 152 86 153 87
rect 151 86 152 87
rect 150 86 151 87
rect 149 86 150 87
rect 148 86 149 87
rect 147 86 148 87
rect 146 86 147 87
rect 145 86 146 87
rect 144 86 145 87
rect 143 86 144 87
rect 142 86 143 87
rect 141 86 142 87
rect 140 86 141 87
rect 139 86 140 87
rect 138 86 139 87
rect 137 86 138 87
rect 136 86 137 87
rect 135 86 136 87
rect 134 86 135 87
rect 133 86 134 87
rect 132 86 133 87
rect 125 86 126 87
rect 124 86 125 87
rect 123 86 124 87
rect 122 86 123 87
rect 121 86 122 87
rect 120 86 121 87
rect 119 86 120 87
rect 118 86 119 87
rect 117 86 118 87
rect 116 86 117 87
rect 115 86 116 87
rect 114 86 115 87
rect 113 86 114 87
rect 112 86 113 87
rect 111 86 112 87
rect 110 86 111 87
rect 109 86 110 87
rect 108 86 109 87
rect 107 86 108 87
rect 106 86 107 87
rect 105 86 106 87
rect 104 86 105 87
rect 103 86 104 87
rect 102 86 103 87
rect 101 86 102 87
rect 100 86 101 87
rect 99 86 100 87
rect 98 86 99 87
rect 97 86 98 87
rect 96 86 97 87
rect 95 86 96 87
rect 94 86 95 87
rect 93 86 94 87
rect 92 86 93 87
rect 91 86 92 87
rect 90 86 91 87
rect 89 86 90 87
rect 88 86 89 87
rect 87 86 88 87
rect 86 86 87 87
rect 85 86 86 87
rect 84 86 85 87
rect 83 86 84 87
rect 82 86 83 87
rect 81 86 82 87
rect 80 86 81 87
rect 79 86 80 87
rect 78 86 79 87
rect 77 86 78 87
rect 76 86 77 87
rect 75 86 76 87
rect 74 86 75 87
rect 73 86 74 87
rect 72 86 73 87
rect 71 86 72 87
rect 70 86 71 87
rect 69 86 70 87
rect 68 86 69 87
rect 67 86 68 87
rect 66 86 67 87
rect 65 86 66 87
rect 480 87 481 88
rect 479 87 480 88
rect 478 87 479 88
rect 477 87 478 88
rect 476 87 477 88
rect 475 87 476 88
rect 474 87 475 88
rect 473 87 474 88
rect 472 87 473 88
rect 471 87 472 88
rect 470 87 471 88
rect 469 87 470 88
rect 468 87 469 88
rect 467 87 468 88
rect 466 87 467 88
rect 465 87 466 88
rect 464 87 465 88
rect 463 87 464 88
rect 462 87 463 88
rect 441 87 442 88
rect 440 87 441 88
rect 408 87 409 88
rect 407 87 408 88
rect 406 87 407 88
rect 405 87 406 88
rect 404 87 405 88
rect 403 87 404 88
rect 402 87 403 88
rect 401 87 402 88
rect 400 87 401 88
rect 399 87 400 88
rect 398 87 399 88
rect 397 87 398 88
rect 237 87 238 88
rect 236 87 237 88
rect 235 87 236 88
rect 234 87 235 88
rect 233 87 234 88
rect 232 87 233 88
rect 231 87 232 88
rect 230 87 231 88
rect 229 87 230 88
rect 228 87 229 88
rect 227 87 228 88
rect 226 87 227 88
rect 225 87 226 88
rect 224 87 225 88
rect 223 87 224 88
rect 222 87 223 88
rect 221 87 222 88
rect 220 87 221 88
rect 219 87 220 88
rect 218 87 219 88
rect 217 87 218 88
rect 216 87 217 88
rect 215 87 216 88
rect 214 87 215 88
rect 213 87 214 88
rect 212 87 213 88
rect 211 87 212 88
rect 210 87 211 88
rect 209 87 210 88
rect 208 87 209 88
rect 207 87 208 88
rect 206 87 207 88
rect 205 87 206 88
rect 204 87 205 88
rect 203 87 204 88
rect 202 87 203 88
rect 164 87 165 88
rect 163 87 164 88
rect 162 87 163 88
rect 161 87 162 88
rect 160 87 161 88
rect 159 87 160 88
rect 158 87 159 88
rect 157 87 158 88
rect 156 87 157 88
rect 155 87 156 88
rect 154 87 155 88
rect 153 87 154 88
rect 152 87 153 88
rect 151 87 152 88
rect 150 87 151 88
rect 149 87 150 88
rect 148 87 149 88
rect 147 87 148 88
rect 146 87 147 88
rect 145 87 146 88
rect 144 87 145 88
rect 143 87 144 88
rect 142 87 143 88
rect 141 87 142 88
rect 140 87 141 88
rect 139 87 140 88
rect 138 87 139 88
rect 137 87 138 88
rect 136 87 137 88
rect 135 87 136 88
rect 134 87 135 88
rect 133 87 134 88
rect 132 87 133 88
rect 125 87 126 88
rect 124 87 125 88
rect 123 87 124 88
rect 122 87 123 88
rect 121 87 122 88
rect 120 87 121 88
rect 119 87 120 88
rect 118 87 119 88
rect 117 87 118 88
rect 116 87 117 88
rect 115 87 116 88
rect 114 87 115 88
rect 113 87 114 88
rect 112 87 113 88
rect 111 87 112 88
rect 110 87 111 88
rect 109 87 110 88
rect 108 87 109 88
rect 107 87 108 88
rect 106 87 107 88
rect 105 87 106 88
rect 104 87 105 88
rect 103 87 104 88
rect 102 87 103 88
rect 101 87 102 88
rect 100 87 101 88
rect 99 87 100 88
rect 98 87 99 88
rect 97 87 98 88
rect 96 87 97 88
rect 95 87 96 88
rect 94 87 95 88
rect 93 87 94 88
rect 92 87 93 88
rect 91 87 92 88
rect 90 87 91 88
rect 89 87 90 88
rect 88 87 89 88
rect 87 87 88 88
rect 86 87 87 88
rect 85 87 86 88
rect 84 87 85 88
rect 83 87 84 88
rect 82 87 83 88
rect 81 87 82 88
rect 80 87 81 88
rect 79 87 80 88
rect 78 87 79 88
rect 77 87 78 88
rect 76 87 77 88
rect 75 87 76 88
rect 74 87 75 88
rect 73 87 74 88
rect 72 87 73 88
rect 71 87 72 88
rect 70 87 71 88
rect 69 87 70 88
rect 68 87 69 88
rect 67 87 68 88
rect 66 87 67 88
rect 65 87 66 88
rect 64 87 65 88
rect 481 88 482 89
rect 480 88 481 89
rect 479 88 480 89
rect 478 88 479 89
rect 477 88 478 89
rect 476 88 477 89
rect 475 88 476 89
rect 474 88 475 89
rect 473 88 474 89
rect 472 88 473 89
rect 471 88 472 89
rect 470 88 471 89
rect 469 88 470 89
rect 468 88 469 89
rect 467 88 468 89
rect 466 88 467 89
rect 465 88 466 89
rect 464 88 465 89
rect 463 88 464 89
rect 462 88 463 89
rect 407 88 408 89
rect 406 88 407 89
rect 405 88 406 89
rect 404 88 405 89
rect 403 88 404 89
rect 402 88 403 89
rect 401 88 402 89
rect 400 88 401 89
rect 399 88 400 89
rect 398 88 399 89
rect 397 88 398 89
rect 240 88 241 89
rect 239 88 240 89
rect 238 88 239 89
rect 237 88 238 89
rect 236 88 237 89
rect 235 88 236 89
rect 234 88 235 89
rect 233 88 234 89
rect 232 88 233 89
rect 231 88 232 89
rect 230 88 231 89
rect 229 88 230 89
rect 228 88 229 89
rect 227 88 228 89
rect 226 88 227 89
rect 225 88 226 89
rect 224 88 225 89
rect 223 88 224 89
rect 222 88 223 89
rect 221 88 222 89
rect 220 88 221 89
rect 219 88 220 89
rect 218 88 219 89
rect 217 88 218 89
rect 216 88 217 89
rect 215 88 216 89
rect 214 88 215 89
rect 213 88 214 89
rect 212 88 213 89
rect 211 88 212 89
rect 210 88 211 89
rect 209 88 210 89
rect 208 88 209 89
rect 207 88 208 89
rect 206 88 207 89
rect 205 88 206 89
rect 204 88 205 89
rect 203 88 204 89
rect 202 88 203 89
rect 201 88 202 89
rect 200 88 201 89
rect 164 88 165 89
rect 163 88 164 89
rect 162 88 163 89
rect 161 88 162 89
rect 160 88 161 89
rect 159 88 160 89
rect 158 88 159 89
rect 157 88 158 89
rect 156 88 157 89
rect 155 88 156 89
rect 154 88 155 89
rect 153 88 154 89
rect 152 88 153 89
rect 151 88 152 89
rect 150 88 151 89
rect 149 88 150 89
rect 148 88 149 89
rect 147 88 148 89
rect 146 88 147 89
rect 145 88 146 89
rect 144 88 145 89
rect 143 88 144 89
rect 142 88 143 89
rect 141 88 142 89
rect 140 88 141 89
rect 139 88 140 89
rect 138 88 139 89
rect 137 88 138 89
rect 136 88 137 89
rect 135 88 136 89
rect 134 88 135 89
rect 133 88 134 89
rect 132 88 133 89
rect 125 88 126 89
rect 124 88 125 89
rect 123 88 124 89
rect 122 88 123 89
rect 121 88 122 89
rect 120 88 121 89
rect 119 88 120 89
rect 118 88 119 89
rect 117 88 118 89
rect 116 88 117 89
rect 115 88 116 89
rect 114 88 115 89
rect 113 88 114 89
rect 112 88 113 89
rect 111 88 112 89
rect 110 88 111 89
rect 109 88 110 89
rect 108 88 109 89
rect 107 88 108 89
rect 106 88 107 89
rect 105 88 106 89
rect 104 88 105 89
rect 103 88 104 89
rect 102 88 103 89
rect 101 88 102 89
rect 100 88 101 89
rect 99 88 100 89
rect 98 88 99 89
rect 97 88 98 89
rect 96 88 97 89
rect 95 88 96 89
rect 94 88 95 89
rect 93 88 94 89
rect 92 88 93 89
rect 91 88 92 89
rect 90 88 91 89
rect 89 88 90 89
rect 88 88 89 89
rect 87 88 88 89
rect 86 88 87 89
rect 85 88 86 89
rect 84 88 85 89
rect 83 88 84 89
rect 82 88 83 89
rect 81 88 82 89
rect 80 88 81 89
rect 79 88 80 89
rect 78 88 79 89
rect 77 88 78 89
rect 76 88 77 89
rect 75 88 76 89
rect 74 88 75 89
rect 73 88 74 89
rect 72 88 73 89
rect 71 88 72 89
rect 70 88 71 89
rect 69 88 70 89
rect 68 88 69 89
rect 67 88 68 89
rect 66 88 67 89
rect 65 88 66 89
rect 64 88 65 89
rect 482 89 483 90
rect 481 89 482 90
rect 480 89 481 90
rect 479 89 480 90
rect 478 89 479 90
rect 477 89 478 90
rect 476 89 477 90
rect 475 89 476 90
rect 474 89 475 90
rect 473 89 474 90
rect 472 89 473 90
rect 471 89 472 90
rect 470 89 471 90
rect 469 89 470 90
rect 468 89 469 90
rect 467 89 468 90
rect 466 89 467 90
rect 465 89 466 90
rect 464 89 465 90
rect 463 89 464 90
rect 462 89 463 90
rect 405 89 406 90
rect 404 89 405 90
rect 403 89 404 90
rect 402 89 403 90
rect 401 89 402 90
rect 400 89 401 90
rect 399 89 400 90
rect 398 89 399 90
rect 397 89 398 90
rect 243 89 244 90
rect 242 89 243 90
rect 241 89 242 90
rect 240 89 241 90
rect 239 89 240 90
rect 238 89 239 90
rect 237 89 238 90
rect 236 89 237 90
rect 235 89 236 90
rect 234 89 235 90
rect 233 89 234 90
rect 232 89 233 90
rect 231 89 232 90
rect 230 89 231 90
rect 229 89 230 90
rect 228 89 229 90
rect 227 89 228 90
rect 226 89 227 90
rect 225 89 226 90
rect 224 89 225 90
rect 223 89 224 90
rect 222 89 223 90
rect 221 89 222 90
rect 220 89 221 90
rect 219 89 220 90
rect 218 89 219 90
rect 217 89 218 90
rect 216 89 217 90
rect 215 89 216 90
rect 214 89 215 90
rect 213 89 214 90
rect 212 89 213 90
rect 211 89 212 90
rect 210 89 211 90
rect 209 89 210 90
rect 208 89 209 90
rect 207 89 208 90
rect 206 89 207 90
rect 205 89 206 90
rect 204 89 205 90
rect 203 89 204 90
rect 202 89 203 90
rect 201 89 202 90
rect 200 89 201 90
rect 199 89 200 90
rect 198 89 199 90
rect 164 89 165 90
rect 163 89 164 90
rect 162 89 163 90
rect 161 89 162 90
rect 160 89 161 90
rect 159 89 160 90
rect 158 89 159 90
rect 157 89 158 90
rect 156 89 157 90
rect 155 89 156 90
rect 154 89 155 90
rect 153 89 154 90
rect 152 89 153 90
rect 151 89 152 90
rect 150 89 151 90
rect 149 89 150 90
rect 148 89 149 90
rect 147 89 148 90
rect 146 89 147 90
rect 145 89 146 90
rect 144 89 145 90
rect 143 89 144 90
rect 142 89 143 90
rect 141 89 142 90
rect 140 89 141 90
rect 139 89 140 90
rect 138 89 139 90
rect 137 89 138 90
rect 136 89 137 90
rect 135 89 136 90
rect 134 89 135 90
rect 133 89 134 90
rect 132 89 133 90
rect 125 89 126 90
rect 124 89 125 90
rect 123 89 124 90
rect 122 89 123 90
rect 121 89 122 90
rect 120 89 121 90
rect 119 89 120 90
rect 118 89 119 90
rect 117 89 118 90
rect 116 89 117 90
rect 115 89 116 90
rect 114 89 115 90
rect 113 89 114 90
rect 112 89 113 90
rect 111 89 112 90
rect 110 89 111 90
rect 109 89 110 90
rect 108 89 109 90
rect 107 89 108 90
rect 106 89 107 90
rect 105 89 106 90
rect 104 89 105 90
rect 103 89 104 90
rect 102 89 103 90
rect 101 89 102 90
rect 100 89 101 90
rect 99 89 100 90
rect 98 89 99 90
rect 97 89 98 90
rect 96 89 97 90
rect 95 89 96 90
rect 94 89 95 90
rect 93 89 94 90
rect 92 89 93 90
rect 91 89 92 90
rect 90 89 91 90
rect 89 89 90 90
rect 88 89 89 90
rect 87 89 88 90
rect 86 89 87 90
rect 85 89 86 90
rect 84 89 85 90
rect 83 89 84 90
rect 82 89 83 90
rect 81 89 82 90
rect 80 89 81 90
rect 79 89 80 90
rect 78 89 79 90
rect 77 89 78 90
rect 76 89 77 90
rect 75 89 76 90
rect 74 89 75 90
rect 73 89 74 90
rect 72 89 73 90
rect 71 89 72 90
rect 70 89 71 90
rect 69 89 70 90
rect 68 89 69 90
rect 67 89 68 90
rect 66 89 67 90
rect 65 89 66 90
rect 64 89 65 90
rect 63 89 64 90
rect 483 90 484 91
rect 482 90 483 91
rect 481 90 482 91
rect 480 90 481 91
rect 479 90 480 91
rect 478 90 479 91
rect 477 90 478 91
rect 476 90 477 91
rect 475 90 476 91
rect 464 90 465 91
rect 463 90 464 91
rect 462 90 463 91
rect 403 90 404 91
rect 402 90 403 91
rect 401 90 402 91
rect 400 90 401 91
rect 399 90 400 91
rect 398 90 399 91
rect 397 90 398 91
rect 245 90 246 91
rect 244 90 245 91
rect 243 90 244 91
rect 242 90 243 91
rect 241 90 242 91
rect 240 90 241 91
rect 239 90 240 91
rect 238 90 239 91
rect 237 90 238 91
rect 236 90 237 91
rect 235 90 236 91
rect 234 90 235 91
rect 233 90 234 91
rect 232 90 233 91
rect 231 90 232 91
rect 230 90 231 91
rect 229 90 230 91
rect 228 90 229 91
rect 227 90 228 91
rect 226 90 227 91
rect 225 90 226 91
rect 224 90 225 91
rect 223 90 224 91
rect 222 90 223 91
rect 221 90 222 91
rect 220 90 221 91
rect 219 90 220 91
rect 218 90 219 91
rect 217 90 218 91
rect 216 90 217 91
rect 215 90 216 91
rect 214 90 215 91
rect 213 90 214 91
rect 212 90 213 91
rect 211 90 212 91
rect 210 90 211 91
rect 209 90 210 91
rect 208 90 209 91
rect 207 90 208 91
rect 206 90 207 91
rect 205 90 206 91
rect 204 90 205 91
rect 203 90 204 91
rect 202 90 203 91
rect 201 90 202 91
rect 200 90 201 91
rect 199 90 200 91
rect 198 90 199 91
rect 197 90 198 91
rect 196 90 197 91
rect 164 90 165 91
rect 163 90 164 91
rect 162 90 163 91
rect 161 90 162 91
rect 160 90 161 91
rect 159 90 160 91
rect 158 90 159 91
rect 157 90 158 91
rect 156 90 157 91
rect 155 90 156 91
rect 154 90 155 91
rect 153 90 154 91
rect 152 90 153 91
rect 151 90 152 91
rect 150 90 151 91
rect 149 90 150 91
rect 148 90 149 91
rect 147 90 148 91
rect 146 90 147 91
rect 145 90 146 91
rect 144 90 145 91
rect 143 90 144 91
rect 142 90 143 91
rect 141 90 142 91
rect 140 90 141 91
rect 139 90 140 91
rect 138 90 139 91
rect 137 90 138 91
rect 136 90 137 91
rect 135 90 136 91
rect 134 90 135 91
rect 133 90 134 91
rect 132 90 133 91
rect 125 90 126 91
rect 124 90 125 91
rect 123 90 124 91
rect 122 90 123 91
rect 121 90 122 91
rect 120 90 121 91
rect 119 90 120 91
rect 118 90 119 91
rect 117 90 118 91
rect 116 90 117 91
rect 115 90 116 91
rect 114 90 115 91
rect 113 90 114 91
rect 112 90 113 91
rect 111 90 112 91
rect 110 90 111 91
rect 109 90 110 91
rect 108 90 109 91
rect 107 90 108 91
rect 106 90 107 91
rect 105 90 106 91
rect 104 90 105 91
rect 103 90 104 91
rect 102 90 103 91
rect 101 90 102 91
rect 100 90 101 91
rect 99 90 100 91
rect 98 90 99 91
rect 97 90 98 91
rect 96 90 97 91
rect 95 90 96 91
rect 94 90 95 91
rect 93 90 94 91
rect 92 90 93 91
rect 91 90 92 91
rect 90 90 91 91
rect 89 90 90 91
rect 88 90 89 91
rect 87 90 88 91
rect 86 90 87 91
rect 85 90 86 91
rect 84 90 85 91
rect 83 90 84 91
rect 82 90 83 91
rect 81 90 82 91
rect 80 90 81 91
rect 79 90 80 91
rect 78 90 79 91
rect 77 90 78 91
rect 76 90 77 91
rect 75 90 76 91
rect 74 90 75 91
rect 73 90 74 91
rect 72 90 73 91
rect 71 90 72 91
rect 70 90 71 91
rect 69 90 70 91
rect 68 90 69 91
rect 67 90 68 91
rect 66 90 67 91
rect 65 90 66 91
rect 64 90 65 91
rect 63 90 64 91
rect 62 90 63 91
rect 483 91 484 92
rect 482 91 483 92
rect 481 91 482 92
rect 480 91 481 92
rect 479 91 480 92
rect 462 91 463 92
rect 402 91 403 92
rect 401 91 402 92
rect 400 91 401 92
rect 399 91 400 92
rect 398 91 399 92
rect 397 91 398 92
rect 248 91 249 92
rect 247 91 248 92
rect 246 91 247 92
rect 245 91 246 92
rect 244 91 245 92
rect 243 91 244 92
rect 242 91 243 92
rect 241 91 242 92
rect 240 91 241 92
rect 239 91 240 92
rect 238 91 239 92
rect 237 91 238 92
rect 236 91 237 92
rect 235 91 236 92
rect 234 91 235 92
rect 233 91 234 92
rect 232 91 233 92
rect 231 91 232 92
rect 230 91 231 92
rect 229 91 230 92
rect 228 91 229 92
rect 227 91 228 92
rect 226 91 227 92
rect 225 91 226 92
rect 224 91 225 92
rect 223 91 224 92
rect 222 91 223 92
rect 221 91 222 92
rect 220 91 221 92
rect 219 91 220 92
rect 218 91 219 92
rect 217 91 218 92
rect 216 91 217 92
rect 215 91 216 92
rect 214 91 215 92
rect 213 91 214 92
rect 212 91 213 92
rect 211 91 212 92
rect 210 91 211 92
rect 209 91 210 92
rect 208 91 209 92
rect 207 91 208 92
rect 206 91 207 92
rect 205 91 206 92
rect 204 91 205 92
rect 203 91 204 92
rect 202 91 203 92
rect 201 91 202 92
rect 200 91 201 92
rect 199 91 200 92
rect 198 91 199 92
rect 197 91 198 92
rect 196 91 197 92
rect 195 91 196 92
rect 194 91 195 92
rect 164 91 165 92
rect 163 91 164 92
rect 162 91 163 92
rect 161 91 162 92
rect 160 91 161 92
rect 159 91 160 92
rect 158 91 159 92
rect 157 91 158 92
rect 156 91 157 92
rect 155 91 156 92
rect 154 91 155 92
rect 153 91 154 92
rect 152 91 153 92
rect 151 91 152 92
rect 150 91 151 92
rect 149 91 150 92
rect 148 91 149 92
rect 147 91 148 92
rect 146 91 147 92
rect 145 91 146 92
rect 144 91 145 92
rect 143 91 144 92
rect 142 91 143 92
rect 141 91 142 92
rect 140 91 141 92
rect 139 91 140 92
rect 138 91 139 92
rect 137 91 138 92
rect 136 91 137 92
rect 135 91 136 92
rect 134 91 135 92
rect 133 91 134 92
rect 132 91 133 92
rect 125 91 126 92
rect 124 91 125 92
rect 123 91 124 92
rect 122 91 123 92
rect 121 91 122 92
rect 120 91 121 92
rect 119 91 120 92
rect 118 91 119 92
rect 117 91 118 92
rect 116 91 117 92
rect 115 91 116 92
rect 114 91 115 92
rect 113 91 114 92
rect 112 91 113 92
rect 111 91 112 92
rect 110 91 111 92
rect 109 91 110 92
rect 108 91 109 92
rect 107 91 108 92
rect 106 91 107 92
rect 105 91 106 92
rect 104 91 105 92
rect 103 91 104 92
rect 102 91 103 92
rect 101 91 102 92
rect 100 91 101 92
rect 99 91 100 92
rect 98 91 99 92
rect 97 91 98 92
rect 96 91 97 92
rect 95 91 96 92
rect 94 91 95 92
rect 93 91 94 92
rect 92 91 93 92
rect 91 91 92 92
rect 90 91 91 92
rect 89 91 90 92
rect 88 91 89 92
rect 87 91 88 92
rect 86 91 87 92
rect 85 91 86 92
rect 84 91 85 92
rect 83 91 84 92
rect 82 91 83 92
rect 81 91 82 92
rect 80 91 81 92
rect 79 91 80 92
rect 78 91 79 92
rect 77 91 78 92
rect 76 91 77 92
rect 75 91 76 92
rect 74 91 75 92
rect 73 91 74 92
rect 72 91 73 92
rect 71 91 72 92
rect 70 91 71 92
rect 69 91 70 92
rect 68 91 69 92
rect 67 91 68 92
rect 66 91 67 92
rect 65 91 66 92
rect 64 91 65 92
rect 63 91 64 92
rect 62 91 63 92
rect 483 92 484 93
rect 482 92 483 93
rect 481 92 482 93
rect 480 92 481 93
rect 462 92 463 93
rect 401 92 402 93
rect 400 92 401 93
rect 399 92 400 93
rect 398 92 399 93
rect 397 92 398 93
rect 250 92 251 93
rect 249 92 250 93
rect 248 92 249 93
rect 247 92 248 93
rect 246 92 247 93
rect 245 92 246 93
rect 244 92 245 93
rect 243 92 244 93
rect 242 92 243 93
rect 241 92 242 93
rect 240 92 241 93
rect 239 92 240 93
rect 238 92 239 93
rect 237 92 238 93
rect 236 92 237 93
rect 235 92 236 93
rect 234 92 235 93
rect 233 92 234 93
rect 232 92 233 93
rect 231 92 232 93
rect 230 92 231 93
rect 229 92 230 93
rect 228 92 229 93
rect 227 92 228 93
rect 226 92 227 93
rect 225 92 226 93
rect 224 92 225 93
rect 223 92 224 93
rect 222 92 223 93
rect 221 92 222 93
rect 220 92 221 93
rect 219 92 220 93
rect 218 92 219 93
rect 217 92 218 93
rect 216 92 217 93
rect 215 92 216 93
rect 214 92 215 93
rect 213 92 214 93
rect 212 92 213 93
rect 211 92 212 93
rect 210 92 211 93
rect 209 92 210 93
rect 208 92 209 93
rect 207 92 208 93
rect 206 92 207 93
rect 205 92 206 93
rect 204 92 205 93
rect 203 92 204 93
rect 202 92 203 93
rect 201 92 202 93
rect 200 92 201 93
rect 199 92 200 93
rect 198 92 199 93
rect 197 92 198 93
rect 196 92 197 93
rect 195 92 196 93
rect 194 92 195 93
rect 193 92 194 93
rect 192 92 193 93
rect 163 92 164 93
rect 162 92 163 93
rect 161 92 162 93
rect 160 92 161 93
rect 159 92 160 93
rect 158 92 159 93
rect 157 92 158 93
rect 156 92 157 93
rect 155 92 156 93
rect 154 92 155 93
rect 153 92 154 93
rect 152 92 153 93
rect 151 92 152 93
rect 150 92 151 93
rect 149 92 150 93
rect 148 92 149 93
rect 147 92 148 93
rect 146 92 147 93
rect 145 92 146 93
rect 144 92 145 93
rect 143 92 144 93
rect 142 92 143 93
rect 141 92 142 93
rect 140 92 141 93
rect 139 92 140 93
rect 138 92 139 93
rect 137 92 138 93
rect 136 92 137 93
rect 135 92 136 93
rect 134 92 135 93
rect 133 92 134 93
rect 132 92 133 93
rect 125 92 126 93
rect 124 92 125 93
rect 123 92 124 93
rect 122 92 123 93
rect 121 92 122 93
rect 120 92 121 93
rect 119 92 120 93
rect 118 92 119 93
rect 117 92 118 93
rect 116 92 117 93
rect 115 92 116 93
rect 114 92 115 93
rect 113 92 114 93
rect 112 92 113 93
rect 111 92 112 93
rect 110 92 111 93
rect 109 92 110 93
rect 108 92 109 93
rect 107 92 108 93
rect 106 92 107 93
rect 105 92 106 93
rect 104 92 105 93
rect 103 92 104 93
rect 102 92 103 93
rect 101 92 102 93
rect 100 92 101 93
rect 99 92 100 93
rect 98 92 99 93
rect 97 92 98 93
rect 96 92 97 93
rect 95 92 96 93
rect 94 92 95 93
rect 93 92 94 93
rect 92 92 93 93
rect 91 92 92 93
rect 90 92 91 93
rect 89 92 90 93
rect 88 92 89 93
rect 87 92 88 93
rect 86 92 87 93
rect 85 92 86 93
rect 84 92 85 93
rect 83 92 84 93
rect 82 92 83 93
rect 81 92 82 93
rect 80 92 81 93
rect 79 92 80 93
rect 78 92 79 93
rect 77 92 78 93
rect 76 92 77 93
rect 75 92 76 93
rect 74 92 75 93
rect 73 92 74 93
rect 72 92 73 93
rect 71 92 72 93
rect 70 92 71 93
rect 69 92 70 93
rect 68 92 69 93
rect 67 92 68 93
rect 66 92 67 93
rect 65 92 66 93
rect 64 92 65 93
rect 63 92 64 93
rect 62 92 63 93
rect 61 92 62 93
rect 483 93 484 94
rect 482 93 483 94
rect 481 93 482 94
rect 400 93 401 94
rect 399 93 400 94
rect 398 93 399 94
rect 397 93 398 94
rect 252 93 253 94
rect 251 93 252 94
rect 250 93 251 94
rect 249 93 250 94
rect 248 93 249 94
rect 247 93 248 94
rect 246 93 247 94
rect 245 93 246 94
rect 244 93 245 94
rect 243 93 244 94
rect 242 93 243 94
rect 241 93 242 94
rect 240 93 241 94
rect 239 93 240 94
rect 238 93 239 94
rect 237 93 238 94
rect 236 93 237 94
rect 235 93 236 94
rect 234 93 235 94
rect 233 93 234 94
rect 232 93 233 94
rect 231 93 232 94
rect 230 93 231 94
rect 229 93 230 94
rect 228 93 229 94
rect 227 93 228 94
rect 226 93 227 94
rect 225 93 226 94
rect 224 93 225 94
rect 223 93 224 94
rect 222 93 223 94
rect 221 93 222 94
rect 220 93 221 94
rect 219 93 220 94
rect 218 93 219 94
rect 217 93 218 94
rect 216 93 217 94
rect 215 93 216 94
rect 214 93 215 94
rect 213 93 214 94
rect 212 93 213 94
rect 211 93 212 94
rect 210 93 211 94
rect 209 93 210 94
rect 208 93 209 94
rect 207 93 208 94
rect 206 93 207 94
rect 205 93 206 94
rect 204 93 205 94
rect 203 93 204 94
rect 202 93 203 94
rect 201 93 202 94
rect 200 93 201 94
rect 199 93 200 94
rect 198 93 199 94
rect 197 93 198 94
rect 196 93 197 94
rect 195 93 196 94
rect 194 93 195 94
rect 193 93 194 94
rect 192 93 193 94
rect 191 93 192 94
rect 163 93 164 94
rect 162 93 163 94
rect 161 93 162 94
rect 160 93 161 94
rect 159 93 160 94
rect 158 93 159 94
rect 157 93 158 94
rect 156 93 157 94
rect 155 93 156 94
rect 154 93 155 94
rect 153 93 154 94
rect 152 93 153 94
rect 151 93 152 94
rect 150 93 151 94
rect 149 93 150 94
rect 148 93 149 94
rect 147 93 148 94
rect 146 93 147 94
rect 145 93 146 94
rect 144 93 145 94
rect 143 93 144 94
rect 142 93 143 94
rect 141 93 142 94
rect 140 93 141 94
rect 139 93 140 94
rect 138 93 139 94
rect 137 93 138 94
rect 136 93 137 94
rect 135 93 136 94
rect 134 93 135 94
rect 133 93 134 94
rect 132 93 133 94
rect 125 93 126 94
rect 124 93 125 94
rect 123 93 124 94
rect 122 93 123 94
rect 121 93 122 94
rect 120 93 121 94
rect 119 93 120 94
rect 118 93 119 94
rect 117 93 118 94
rect 116 93 117 94
rect 115 93 116 94
rect 114 93 115 94
rect 113 93 114 94
rect 112 93 113 94
rect 111 93 112 94
rect 110 93 111 94
rect 109 93 110 94
rect 108 93 109 94
rect 107 93 108 94
rect 106 93 107 94
rect 105 93 106 94
rect 104 93 105 94
rect 103 93 104 94
rect 102 93 103 94
rect 101 93 102 94
rect 100 93 101 94
rect 99 93 100 94
rect 98 93 99 94
rect 97 93 98 94
rect 96 93 97 94
rect 95 93 96 94
rect 94 93 95 94
rect 93 93 94 94
rect 92 93 93 94
rect 91 93 92 94
rect 90 93 91 94
rect 89 93 90 94
rect 88 93 89 94
rect 87 93 88 94
rect 86 93 87 94
rect 85 93 86 94
rect 84 93 85 94
rect 83 93 84 94
rect 82 93 83 94
rect 81 93 82 94
rect 80 93 81 94
rect 79 93 80 94
rect 78 93 79 94
rect 77 93 78 94
rect 76 93 77 94
rect 75 93 76 94
rect 74 93 75 94
rect 73 93 74 94
rect 72 93 73 94
rect 71 93 72 94
rect 70 93 71 94
rect 69 93 70 94
rect 68 93 69 94
rect 67 93 68 94
rect 66 93 67 94
rect 65 93 66 94
rect 64 93 65 94
rect 63 93 64 94
rect 62 93 63 94
rect 61 93 62 94
rect 60 93 61 94
rect 483 94 484 95
rect 482 94 483 95
rect 481 94 482 95
rect 400 94 401 95
rect 399 94 400 95
rect 398 94 399 95
rect 397 94 398 95
rect 254 94 255 95
rect 253 94 254 95
rect 252 94 253 95
rect 251 94 252 95
rect 250 94 251 95
rect 249 94 250 95
rect 248 94 249 95
rect 247 94 248 95
rect 246 94 247 95
rect 245 94 246 95
rect 244 94 245 95
rect 243 94 244 95
rect 242 94 243 95
rect 241 94 242 95
rect 240 94 241 95
rect 239 94 240 95
rect 238 94 239 95
rect 237 94 238 95
rect 236 94 237 95
rect 235 94 236 95
rect 234 94 235 95
rect 233 94 234 95
rect 232 94 233 95
rect 231 94 232 95
rect 230 94 231 95
rect 229 94 230 95
rect 228 94 229 95
rect 227 94 228 95
rect 226 94 227 95
rect 225 94 226 95
rect 224 94 225 95
rect 223 94 224 95
rect 222 94 223 95
rect 221 94 222 95
rect 220 94 221 95
rect 219 94 220 95
rect 218 94 219 95
rect 217 94 218 95
rect 216 94 217 95
rect 215 94 216 95
rect 214 94 215 95
rect 213 94 214 95
rect 212 94 213 95
rect 211 94 212 95
rect 210 94 211 95
rect 209 94 210 95
rect 208 94 209 95
rect 207 94 208 95
rect 206 94 207 95
rect 205 94 206 95
rect 204 94 205 95
rect 203 94 204 95
rect 202 94 203 95
rect 201 94 202 95
rect 200 94 201 95
rect 199 94 200 95
rect 198 94 199 95
rect 197 94 198 95
rect 196 94 197 95
rect 195 94 196 95
rect 194 94 195 95
rect 193 94 194 95
rect 192 94 193 95
rect 191 94 192 95
rect 190 94 191 95
rect 189 94 190 95
rect 163 94 164 95
rect 162 94 163 95
rect 161 94 162 95
rect 160 94 161 95
rect 159 94 160 95
rect 158 94 159 95
rect 157 94 158 95
rect 156 94 157 95
rect 155 94 156 95
rect 154 94 155 95
rect 153 94 154 95
rect 152 94 153 95
rect 151 94 152 95
rect 150 94 151 95
rect 149 94 150 95
rect 148 94 149 95
rect 147 94 148 95
rect 146 94 147 95
rect 145 94 146 95
rect 144 94 145 95
rect 143 94 144 95
rect 142 94 143 95
rect 141 94 142 95
rect 140 94 141 95
rect 139 94 140 95
rect 138 94 139 95
rect 137 94 138 95
rect 136 94 137 95
rect 135 94 136 95
rect 134 94 135 95
rect 133 94 134 95
rect 132 94 133 95
rect 124 94 125 95
rect 123 94 124 95
rect 122 94 123 95
rect 121 94 122 95
rect 120 94 121 95
rect 119 94 120 95
rect 118 94 119 95
rect 117 94 118 95
rect 116 94 117 95
rect 115 94 116 95
rect 114 94 115 95
rect 113 94 114 95
rect 112 94 113 95
rect 111 94 112 95
rect 110 94 111 95
rect 109 94 110 95
rect 108 94 109 95
rect 107 94 108 95
rect 106 94 107 95
rect 105 94 106 95
rect 104 94 105 95
rect 103 94 104 95
rect 102 94 103 95
rect 101 94 102 95
rect 100 94 101 95
rect 99 94 100 95
rect 98 94 99 95
rect 97 94 98 95
rect 96 94 97 95
rect 95 94 96 95
rect 94 94 95 95
rect 93 94 94 95
rect 92 94 93 95
rect 91 94 92 95
rect 90 94 91 95
rect 89 94 90 95
rect 88 94 89 95
rect 87 94 88 95
rect 86 94 87 95
rect 85 94 86 95
rect 84 94 85 95
rect 83 94 84 95
rect 82 94 83 95
rect 81 94 82 95
rect 80 94 81 95
rect 79 94 80 95
rect 78 94 79 95
rect 77 94 78 95
rect 76 94 77 95
rect 75 94 76 95
rect 74 94 75 95
rect 73 94 74 95
rect 72 94 73 95
rect 71 94 72 95
rect 70 94 71 95
rect 69 94 70 95
rect 68 94 69 95
rect 67 94 68 95
rect 66 94 67 95
rect 65 94 66 95
rect 64 94 65 95
rect 63 94 64 95
rect 62 94 63 95
rect 61 94 62 95
rect 60 94 61 95
rect 483 95 484 96
rect 482 95 483 96
rect 399 95 400 96
rect 398 95 399 96
rect 397 95 398 96
rect 256 95 257 96
rect 255 95 256 96
rect 254 95 255 96
rect 253 95 254 96
rect 252 95 253 96
rect 251 95 252 96
rect 250 95 251 96
rect 249 95 250 96
rect 248 95 249 96
rect 247 95 248 96
rect 246 95 247 96
rect 245 95 246 96
rect 244 95 245 96
rect 243 95 244 96
rect 242 95 243 96
rect 241 95 242 96
rect 240 95 241 96
rect 239 95 240 96
rect 238 95 239 96
rect 237 95 238 96
rect 236 95 237 96
rect 235 95 236 96
rect 234 95 235 96
rect 233 95 234 96
rect 232 95 233 96
rect 231 95 232 96
rect 230 95 231 96
rect 229 95 230 96
rect 228 95 229 96
rect 227 95 228 96
rect 226 95 227 96
rect 225 95 226 96
rect 224 95 225 96
rect 223 95 224 96
rect 222 95 223 96
rect 221 95 222 96
rect 220 95 221 96
rect 219 95 220 96
rect 218 95 219 96
rect 217 95 218 96
rect 216 95 217 96
rect 215 95 216 96
rect 214 95 215 96
rect 213 95 214 96
rect 212 95 213 96
rect 211 95 212 96
rect 210 95 211 96
rect 209 95 210 96
rect 208 95 209 96
rect 207 95 208 96
rect 206 95 207 96
rect 205 95 206 96
rect 204 95 205 96
rect 203 95 204 96
rect 202 95 203 96
rect 201 95 202 96
rect 200 95 201 96
rect 199 95 200 96
rect 198 95 199 96
rect 197 95 198 96
rect 196 95 197 96
rect 195 95 196 96
rect 194 95 195 96
rect 193 95 194 96
rect 192 95 193 96
rect 191 95 192 96
rect 190 95 191 96
rect 189 95 190 96
rect 188 95 189 96
rect 162 95 163 96
rect 161 95 162 96
rect 160 95 161 96
rect 159 95 160 96
rect 158 95 159 96
rect 157 95 158 96
rect 156 95 157 96
rect 155 95 156 96
rect 154 95 155 96
rect 153 95 154 96
rect 152 95 153 96
rect 151 95 152 96
rect 150 95 151 96
rect 149 95 150 96
rect 148 95 149 96
rect 147 95 148 96
rect 146 95 147 96
rect 145 95 146 96
rect 144 95 145 96
rect 143 95 144 96
rect 142 95 143 96
rect 141 95 142 96
rect 140 95 141 96
rect 139 95 140 96
rect 138 95 139 96
rect 137 95 138 96
rect 136 95 137 96
rect 135 95 136 96
rect 134 95 135 96
rect 133 95 134 96
rect 132 95 133 96
rect 131 95 132 96
rect 124 95 125 96
rect 123 95 124 96
rect 122 95 123 96
rect 121 95 122 96
rect 120 95 121 96
rect 119 95 120 96
rect 118 95 119 96
rect 117 95 118 96
rect 116 95 117 96
rect 115 95 116 96
rect 114 95 115 96
rect 113 95 114 96
rect 112 95 113 96
rect 111 95 112 96
rect 110 95 111 96
rect 109 95 110 96
rect 108 95 109 96
rect 107 95 108 96
rect 106 95 107 96
rect 105 95 106 96
rect 104 95 105 96
rect 103 95 104 96
rect 102 95 103 96
rect 101 95 102 96
rect 100 95 101 96
rect 99 95 100 96
rect 98 95 99 96
rect 97 95 98 96
rect 96 95 97 96
rect 95 95 96 96
rect 94 95 95 96
rect 93 95 94 96
rect 92 95 93 96
rect 91 95 92 96
rect 90 95 91 96
rect 89 95 90 96
rect 88 95 89 96
rect 87 95 88 96
rect 86 95 87 96
rect 85 95 86 96
rect 84 95 85 96
rect 83 95 84 96
rect 82 95 83 96
rect 81 95 82 96
rect 80 95 81 96
rect 79 95 80 96
rect 78 95 79 96
rect 77 95 78 96
rect 76 95 77 96
rect 75 95 76 96
rect 74 95 75 96
rect 73 95 74 96
rect 72 95 73 96
rect 71 95 72 96
rect 70 95 71 96
rect 69 95 70 96
rect 68 95 69 96
rect 67 95 68 96
rect 66 95 67 96
rect 65 95 66 96
rect 64 95 65 96
rect 63 95 64 96
rect 62 95 63 96
rect 61 95 62 96
rect 60 95 61 96
rect 59 95 60 96
rect 483 96 484 97
rect 482 96 483 97
rect 399 96 400 97
rect 398 96 399 97
rect 397 96 398 97
rect 257 96 258 97
rect 256 96 257 97
rect 255 96 256 97
rect 254 96 255 97
rect 253 96 254 97
rect 252 96 253 97
rect 251 96 252 97
rect 250 96 251 97
rect 249 96 250 97
rect 248 96 249 97
rect 247 96 248 97
rect 246 96 247 97
rect 245 96 246 97
rect 244 96 245 97
rect 243 96 244 97
rect 242 96 243 97
rect 241 96 242 97
rect 240 96 241 97
rect 239 96 240 97
rect 238 96 239 97
rect 237 96 238 97
rect 236 96 237 97
rect 235 96 236 97
rect 234 96 235 97
rect 233 96 234 97
rect 232 96 233 97
rect 231 96 232 97
rect 230 96 231 97
rect 229 96 230 97
rect 228 96 229 97
rect 227 96 228 97
rect 226 96 227 97
rect 225 96 226 97
rect 224 96 225 97
rect 223 96 224 97
rect 222 96 223 97
rect 221 96 222 97
rect 220 96 221 97
rect 219 96 220 97
rect 218 96 219 97
rect 217 96 218 97
rect 216 96 217 97
rect 215 96 216 97
rect 214 96 215 97
rect 213 96 214 97
rect 212 96 213 97
rect 211 96 212 97
rect 210 96 211 97
rect 209 96 210 97
rect 208 96 209 97
rect 207 96 208 97
rect 206 96 207 97
rect 205 96 206 97
rect 204 96 205 97
rect 203 96 204 97
rect 202 96 203 97
rect 201 96 202 97
rect 200 96 201 97
rect 199 96 200 97
rect 198 96 199 97
rect 197 96 198 97
rect 196 96 197 97
rect 195 96 196 97
rect 194 96 195 97
rect 193 96 194 97
rect 192 96 193 97
rect 191 96 192 97
rect 190 96 191 97
rect 189 96 190 97
rect 188 96 189 97
rect 187 96 188 97
rect 162 96 163 97
rect 161 96 162 97
rect 160 96 161 97
rect 159 96 160 97
rect 158 96 159 97
rect 157 96 158 97
rect 156 96 157 97
rect 155 96 156 97
rect 154 96 155 97
rect 153 96 154 97
rect 152 96 153 97
rect 151 96 152 97
rect 150 96 151 97
rect 149 96 150 97
rect 148 96 149 97
rect 147 96 148 97
rect 146 96 147 97
rect 145 96 146 97
rect 144 96 145 97
rect 143 96 144 97
rect 142 96 143 97
rect 141 96 142 97
rect 140 96 141 97
rect 139 96 140 97
rect 138 96 139 97
rect 137 96 138 97
rect 136 96 137 97
rect 135 96 136 97
rect 134 96 135 97
rect 133 96 134 97
rect 132 96 133 97
rect 131 96 132 97
rect 124 96 125 97
rect 123 96 124 97
rect 122 96 123 97
rect 121 96 122 97
rect 120 96 121 97
rect 119 96 120 97
rect 118 96 119 97
rect 117 96 118 97
rect 116 96 117 97
rect 115 96 116 97
rect 114 96 115 97
rect 113 96 114 97
rect 112 96 113 97
rect 111 96 112 97
rect 110 96 111 97
rect 109 96 110 97
rect 108 96 109 97
rect 107 96 108 97
rect 106 96 107 97
rect 105 96 106 97
rect 104 96 105 97
rect 103 96 104 97
rect 102 96 103 97
rect 101 96 102 97
rect 100 96 101 97
rect 99 96 100 97
rect 98 96 99 97
rect 97 96 98 97
rect 96 96 97 97
rect 95 96 96 97
rect 94 96 95 97
rect 93 96 94 97
rect 92 96 93 97
rect 91 96 92 97
rect 90 96 91 97
rect 89 96 90 97
rect 88 96 89 97
rect 87 96 88 97
rect 86 96 87 97
rect 85 96 86 97
rect 84 96 85 97
rect 83 96 84 97
rect 82 96 83 97
rect 81 96 82 97
rect 80 96 81 97
rect 79 96 80 97
rect 78 96 79 97
rect 77 96 78 97
rect 76 96 77 97
rect 75 96 76 97
rect 74 96 75 97
rect 73 96 74 97
rect 72 96 73 97
rect 71 96 72 97
rect 70 96 71 97
rect 69 96 70 97
rect 68 96 69 97
rect 67 96 68 97
rect 66 96 67 97
rect 65 96 66 97
rect 64 96 65 97
rect 63 96 64 97
rect 62 96 63 97
rect 61 96 62 97
rect 60 96 61 97
rect 59 96 60 97
rect 58 96 59 97
rect 483 97 484 98
rect 482 97 483 98
rect 481 97 482 98
rect 399 97 400 98
rect 398 97 399 98
rect 397 97 398 98
rect 259 97 260 98
rect 258 97 259 98
rect 257 97 258 98
rect 256 97 257 98
rect 255 97 256 98
rect 254 97 255 98
rect 253 97 254 98
rect 252 97 253 98
rect 251 97 252 98
rect 250 97 251 98
rect 249 97 250 98
rect 248 97 249 98
rect 247 97 248 98
rect 246 97 247 98
rect 245 97 246 98
rect 244 97 245 98
rect 243 97 244 98
rect 242 97 243 98
rect 241 97 242 98
rect 240 97 241 98
rect 239 97 240 98
rect 238 97 239 98
rect 237 97 238 98
rect 236 97 237 98
rect 235 97 236 98
rect 234 97 235 98
rect 233 97 234 98
rect 232 97 233 98
rect 231 97 232 98
rect 230 97 231 98
rect 229 97 230 98
rect 228 97 229 98
rect 227 97 228 98
rect 226 97 227 98
rect 225 97 226 98
rect 224 97 225 98
rect 223 97 224 98
rect 222 97 223 98
rect 221 97 222 98
rect 220 97 221 98
rect 219 97 220 98
rect 218 97 219 98
rect 217 97 218 98
rect 216 97 217 98
rect 215 97 216 98
rect 214 97 215 98
rect 213 97 214 98
rect 212 97 213 98
rect 211 97 212 98
rect 210 97 211 98
rect 209 97 210 98
rect 208 97 209 98
rect 207 97 208 98
rect 206 97 207 98
rect 205 97 206 98
rect 204 97 205 98
rect 203 97 204 98
rect 202 97 203 98
rect 201 97 202 98
rect 200 97 201 98
rect 199 97 200 98
rect 198 97 199 98
rect 197 97 198 98
rect 196 97 197 98
rect 195 97 196 98
rect 194 97 195 98
rect 193 97 194 98
rect 192 97 193 98
rect 191 97 192 98
rect 190 97 191 98
rect 189 97 190 98
rect 188 97 189 98
rect 187 97 188 98
rect 186 97 187 98
rect 162 97 163 98
rect 161 97 162 98
rect 160 97 161 98
rect 159 97 160 98
rect 158 97 159 98
rect 157 97 158 98
rect 156 97 157 98
rect 155 97 156 98
rect 154 97 155 98
rect 153 97 154 98
rect 152 97 153 98
rect 151 97 152 98
rect 150 97 151 98
rect 149 97 150 98
rect 148 97 149 98
rect 147 97 148 98
rect 146 97 147 98
rect 145 97 146 98
rect 144 97 145 98
rect 143 97 144 98
rect 142 97 143 98
rect 141 97 142 98
rect 140 97 141 98
rect 139 97 140 98
rect 138 97 139 98
rect 137 97 138 98
rect 136 97 137 98
rect 135 97 136 98
rect 134 97 135 98
rect 133 97 134 98
rect 132 97 133 98
rect 131 97 132 98
rect 124 97 125 98
rect 123 97 124 98
rect 122 97 123 98
rect 121 97 122 98
rect 120 97 121 98
rect 119 97 120 98
rect 118 97 119 98
rect 117 97 118 98
rect 116 97 117 98
rect 115 97 116 98
rect 114 97 115 98
rect 113 97 114 98
rect 112 97 113 98
rect 111 97 112 98
rect 110 97 111 98
rect 109 97 110 98
rect 108 97 109 98
rect 107 97 108 98
rect 106 97 107 98
rect 105 97 106 98
rect 104 97 105 98
rect 103 97 104 98
rect 102 97 103 98
rect 101 97 102 98
rect 100 97 101 98
rect 99 97 100 98
rect 98 97 99 98
rect 97 97 98 98
rect 96 97 97 98
rect 95 97 96 98
rect 94 97 95 98
rect 93 97 94 98
rect 92 97 93 98
rect 91 97 92 98
rect 90 97 91 98
rect 89 97 90 98
rect 88 97 89 98
rect 87 97 88 98
rect 86 97 87 98
rect 85 97 86 98
rect 84 97 85 98
rect 83 97 84 98
rect 82 97 83 98
rect 81 97 82 98
rect 80 97 81 98
rect 79 97 80 98
rect 78 97 79 98
rect 77 97 78 98
rect 76 97 77 98
rect 75 97 76 98
rect 74 97 75 98
rect 73 97 74 98
rect 72 97 73 98
rect 71 97 72 98
rect 70 97 71 98
rect 69 97 70 98
rect 68 97 69 98
rect 67 97 68 98
rect 66 97 67 98
rect 65 97 66 98
rect 64 97 65 98
rect 63 97 64 98
rect 62 97 63 98
rect 61 97 62 98
rect 60 97 61 98
rect 59 97 60 98
rect 58 97 59 98
rect 57 97 58 98
rect 482 98 483 99
rect 481 98 482 99
rect 462 98 463 99
rect 261 98 262 99
rect 260 98 261 99
rect 259 98 260 99
rect 258 98 259 99
rect 257 98 258 99
rect 256 98 257 99
rect 255 98 256 99
rect 254 98 255 99
rect 253 98 254 99
rect 252 98 253 99
rect 251 98 252 99
rect 250 98 251 99
rect 249 98 250 99
rect 248 98 249 99
rect 247 98 248 99
rect 246 98 247 99
rect 245 98 246 99
rect 244 98 245 99
rect 243 98 244 99
rect 242 98 243 99
rect 241 98 242 99
rect 240 98 241 99
rect 239 98 240 99
rect 238 98 239 99
rect 237 98 238 99
rect 236 98 237 99
rect 235 98 236 99
rect 234 98 235 99
rect 233 98 234 99
rect 232 98 233 99
rect 231 98 232 99
rect 230 98 231 99
rect 229 98 230 99
rect 228 98 229 99
rect 227 98 228 99
rect 226 98 227 99
rect 225 98 226 99
rect 224 98 225 99
rect 223 98 224 99
rect 222 98 223 99
rect 221 98 222 99
rect 220 98 221 99
rect 219 98 220 99
rect 218 98 219 99
rect 217 98 218 99
rect 216 98 217 99
rect 215 98 216 99
rect 214 98 215 99
rect 213 98 214 99
rect 212 98 213 99
rect 211 98 212 99
rect 210 98 211 99
rect 209 98 210 99
rect 208 98 209 99
rect 207 98 208 99
rect 206 98 207 99
rect 205 98 206 99
rect 204 98 205 99
rect 203 98 204 99
rect 202 98 203 99
rect 201 98 202 99
rect 200 98 201 99
rect 199 98 200 99
rect 198 98 199 99
rect 197 98 198 99
rect 196 98 197 99
rect 195 98 196 99
rect 194 98 195 99
rect 193 98 194 99
rect 192 98 193 99
rect 191 98 192 99
rect 190 98 191 99
rect 189 98 190 99
rect 188 98 189 99
rect 187 98 188 99
rect 186 98 187 99
rect 185 98 186 99
rect 161 98 162 99
rect 160 98 161 99
rect 159 98 160 99
rect 158 98 159 99
rect 157 98 158 99
rect 156 98 157 99
rect 155 98 156 99
rect 154 98 155 99
rect 153 98 154 99
rect 152 98 153 99
rect 151 98 152 99
rect 150 98 151 99
rect 149 98 150 99
rect 148 98 149 99
rect 147 98 148 99
rect 146 98 147 99
rect 145 98 146 99
rect 144 98 145 99
rect 143 98 144 99
rect 142 98 143 99
rect 141 98 142 99
rect 140 98 141 99
rect 139 98 140 99
rect 138 98 139 99
rect 137 98 138 99
rect 136 98 137 99
rect 135 98 136 99
rect 134 98 135 99
rect 133 98 134 99
rect 132 98 133 99
rect 131 98 132 99
rect 123 98 124 99
rect 122 98 123 99
rect 121 98 122 99
rect 120 98 121 99
rect 119 98 120 99
rect 118 98 119 99
rect 117 98 118 99
rect 116 98 117 99
rect 115 98 116 99
rect 114 98 115 99
rect 113 98 114 99
rect 112 98 113 99
rect 111 98 112 99
rect 110 98 111 99
rect 109 98 110 99
rect 108 98 109 99
rect 107 98 108 99
rect 106 98 107 99
rect 105 98 106 99
rect 104 98 105 99
rect 103 98 104 99
rect 102 98 103 99
rect 101 98 102 99
rect 100 98 101 99
rect 99 98 100 99
rect 98 98 99 99
rect 97 98 98 99
rect 96 98 97 99
rect 95 98 96 99
rect 94 98 95 99
rect 93 98 94 99
rect 92 98 93 99
rect 91 98 92 99
rect 90 98 91 99
rect 89 98 90 99
rect 88 98 89 99
rect 87 98 88 99
rect 86 98 87 99
rect 85 98 86 99
rect 84 98 85 99
rect 83 98 84 99
rect 82 98 83 99
rect 81 98 82 99
rect 80 98 81 99
rect 79 98 80 99
rect 78 98 79 99
rect 77 98 78 99
rect 76 98 77 99
rect 75 98 76 99
rect 74 98 75 99
rect 73 98 74 99
rect 72 98 73 99
rect 71 98 72 99
rect 70 98 71 99
rect 69 98 70 99
rect 68 98 69 99
rect 67 98 68 99
rect 66 98 67 99
rect 65 98 66 99
rect 64 98 65 99
rect 63 98 64 99
rect 62 98 63 99
rect 61 98 62 99
rect 60 98 61 99
rect 59 98 60 99
rect 58 98 59 99
rect 57 98 58 99
rect 56 98 57 99
rect 482 99 483 100
rect 481 99 482 100
rect 480 99 481 100
rect 462 99 463 100
rect 262 99 263 100
rect 261 99 262 100
rect 260 99 261 100
rect 259 99 260 100
rect 258 99 259 100
rect 257 99 258 100
rect 256 99 257 100
rect 255 99 256 100
rect 254 99 255 100
rect 253 99 254 100
rect 252 99 253 100
rect 251 99 252 100
rect 250 99 251 100
rect 249 99 250 100
rect 248 99 249 100
rect 247 99 248 100
rect 246 99 247 100
rect 245 99 246 100
rect 244 99 245 100
rect 243 99 244 100
rect 242 99 243 100
rect 241 99 242 100
rect 240 99 241 100
rect 239 99 240 100
rect 238 99 239 100
rect 237 99 238 100
rect 236 99 237 100
rect 235 99 236 100
rect 234 99 235 100
rect 233 99 234 100
rect 232 99 233 100
rect 231 99 232 100
rect 230 99 231 100
rect 229 99 230 100
rect 228 99 229 100
rect 227 99 228 100
rect 226 99 227 100
rect 225 99 226 100
rect 224 99 225 100
rect 223 99 224 100
rect 222 99 223 100
rect 221 99 222 100
rect 220 99 221 100
rect 219 99 220 100
rect 218 99 219 100
rect 217 99 218 100
rect 216 99 217 100
rect 215 99 216 100
rect 214 99 215 100
rect 213 99 214 100
rect 212 99 213 100
rect 211 99 212 100
rect 210 99 211 100
rect 209 99 210 100
rect 208 99 209 100
rect 207 99 208 100
rect 206 99 207 100
rect 205 99 206 100
rect 204 99 205 100
rect 203 99 204 100
rect 202 99 203 100
rect 201 99 202 100
rect 200 99 201 100
rect 199 99 200 100
rect 198 99 199 100
rect 197 99 198 100
rect 196 99 197 100
rect 195 99 196 100
rect 194 99 195 100
rect 193 99 194 100
rect 192 99 193 100
rect 191 99 192 100
rect 190 99 191 100
rect 189 99 190 100
rect 188 99 189 100
rect 187 99 188 100
rect 186 99 187 100
rect 185 99 186 100
rect 184 99 185 100
rect 161 99 162 100
rect 160 99 161 100
rect 159 99 160 100
rect 158 99 159 100
rect 157 99 158 100
rect 156 99 157 100
rect 155 99 156 100
rect 154 99 155 100
rect 153 99 154 100
rect 152 99 153 100
rect 151 99 152 100
rect 150 99 151 100
rect 149 99 150 100
rect 148 99 149 100
rect 147 99 148 100
rect 146 99 147 100
rect 145 99 146 100
rect 144 99 145 100
rect 143 99 144 100
rect 142 99 143 100
rect 141 99 142 100
rect 140 99 141 100
rect 139 99 140 100
rect 138 99 139 100
rect 137 99 138 100
rect 136 99 137 100
rect 135 99 136 100
rect 134 99 135 100
rect 133 99 134 100
rect 132 99 133 100
rect 131 99 132 100
rect 123 99 124 100
rect 122 99 123 100
rect 121 99 122 100
rect 120 99 121 100
rect 119 99 120 100
rect 118 99 119 100
rect 117 99 118 100
rect 116 99 117 100
rect 115 99 116 100
rect 114 99 115 100
rect 113 99 114 100
rect 112 99 113 100
rect 111 99 112 100
rect 110 99 111 100
rect 109 99 110 100
rect 108 99 109 100
rect 107 99 108 100
rect 106 99 107 100
rect 105 99 106 100
rect 104 99 105 100
rect 103 99 104 100
rect 102 99 103 100
rect 101 99 102 100
rect 100 99 101 100
rect 99 99 100 100
rect 98 99 99 100
rect 97 99 98 100
rect 96 99 97 100
rect 95 99 96 100
rect 94 99 95 100
rect 93 99 94 100
rect 92 99 93 100
rect 91 99 92 100
rect 90 99 91 100
rect 89 99 90 100
rect 88 99 89 100
rect 87 99 88 100
rect 86 99 87 100
rect 85 99 86 100
rect 84 99 85 100
rect 83 99 84 100
rect 82 99 83 100
rect 81 99 82 100
rect 80 99 81 100
rect 79 99 80 100
rect 78 99 79 100
rect 77 99 78 100
rect 74 99 75 100
rect 73 99 74 100
rect 72 99 73 100
rect 71 99 72 100
rect 70 99 71 100
rect 69 99 70 100
rect 68 99 69 100
rect 67 99 68 100
rect 66 99 67 100
rect 65 99 66 100
rect 64 99 65 100
rect 63 99 64 100
rect 62 99 63 100
rect 61 99 62 100
rect 60 99 61 100
rect 59 99 60 100
rect 58 99 59 100
rect 57 99 58 100
rect 56 99 57 100
rect 55 99 56 100
rect 481 100 482 101
rect 480 100 481 101
rect 479 100 480 101
rect 463 100 464 101
rect 462 100 463 101
rect 264 100 265 101
rect 263 100 264 101
rect 262 100 263 101
rect 261 100 262 101
rect 260 100 261 101
rect 259 100 260 101
rect 258 100 259 101
rect 257 100 258 101
rect 256 100 257 101
rect 255 100 256 101
rect 254 100 255 101
rect 253 100 254 101
rect 252 100 253 101
rect 251 100 252 101
rect 250 100 251 101
rect 249 100 250 101
rect 248 100 249 101
rect 247 100 248 101
rect 246 100 247 101
rect 245 100 246 101
rect 244 100 245 101
rect 243 100 244 101
rect 242 100 243 101
rect 241 100 242 101
rect 240 100 241 101
rect 239 100 240 101
rect 238 100 239 101
rect 237 100 238 101
rect 236 100 237 101
rect 235 100 236 101
rect 234 100 235 101
rect 233 100 234 101
rect 232 100 233 101
rect 231 100 232 101
rect 230 100 231 101
rect 229 100 230 101
rect 228 100 229 101
rect 227 100 228 101
rect 226 100 227 101
rect 225 100 226 101
rect 224 100 225 101
rect 223 100 224 101
rect 222 100 223 101
rect 221 100 222 101
rect 220 100 221 101
rect 219 100 220 101
rect 218 100 219 101
rect 217 100 218 101
rect 216 100 217 101
rect 215 100 216 101
rect 214 100 215 101
rect 213 100 214 101
rect 212 100 213 101
rect 211 100 212 101
rect 210 100 211 101
rect 209 100 210 101
rect 208 100 209 101
rect 207 100 208 101
rect 206 100 207 101
rect 205 100 206 101
rect 204 100 205 101
rect 203 100 204 101
rect 202 100 203 101
rect 201 100 202 101
rect 200 100 201 101
rect 199 100 200 101
rect 198 100 199 101
rect 197 100 198 101
rect 196 100 197 101
rect 195 100 196 101
rect 194 100 195 101
rect 193 100 194 101
rect 192 100 193 101
rect 191 100 192 101
rect 190 100 191 101
rect 189 100 190 101
rect 188 100 189 101
rect 187 100 188 101
rect 186 100 187 101
rect 185 100 186 101
rect 184 100 185 101
rect 183 100 184 101
rect 161 100 162 101
rect 160 100 161 101
rect 159 100 160 101
rect 158 100 159 101
rect 157 100 158 101
rect 156 100 157 101
rect 155 100 156 101
rect 154 100 155 101
rect 153 100 154 101
rect 152 100 153 101
rect 151 100 152 101
rect 150 100 151 101
rect 149 100 150 101
rect 148 100 149 101
rect 147 100 148 101
rect 146 100 147 101
rect 145 100 146 101
rect 144 100 145 101
rect 143 100 144 101
rect 142 100 143 101
rect 141 100 142 101
rect 140 100 141 101
rect 139 100 140 101
rect 138 100 139 101
rect 137 100 138 101
rect 136 100 137 101
rect 135 100 136 101
rect 134 100 135 101
rect 133 100 134 101
rect 132 100 133 101
rect 131 100 132 101
rect 123 100 124 101
rect 122 100 123 101
rect 121 100 122 101
rect 120 100 121 101
rect 119 100 120 101
rect 118 100 119 101
rect 117 100 118 101
rect 116 100 117 101
rect 115 100 116 101
rect 114 100 115 101
rect 113 100 114 101
rect 112 100 113 101
rect 111 100 112 101
rect 110 100 111 101
rect 109 100 110 101
rect 108 100 109 101
rect 107 100 108 101
rect 106 100 107 101
rect 105 100 106 101
rect 104 100 105 101
rect 103 100 104 101
rect 102 100 103 101
rect 101 100 102 101
rect 100 100 101 101
rect 99 100 100 101
rect 98 100 99 101
rect 97 100 98 101
rect 96 100 97 101
rect 95 100 96 101
rect 94 100 95 101
rect 93 100 94 101
rect 92 100 93 101
rect 91 100 92 101
rect 90 100 91 101
rect 89 100 90 101
rect 88 100 89 101
rect 87 100 88 101
rect 86 100 87 101
rect 85 100 86 101
rect 84 100 85 101
rect 83 100 84 101
rect 82 100 83 101
rect 81 100 82 101
rect 80 100 81 101
rect 79 100 80 101
rect 78 100 79 101
rect 77 100 78 101
rect 73 100 74 101
rect 72 100 73 101
rect 71 100 72 101
rect 70 100 71 101
rect 69 100 70 101
rect 68 100 69 101
rect 67 100 68 101
rect 66 100 67 101
rect 65 100 66 101
rect 64 100 65 101
rect 63 100 64 101
rect 62 100 63 101
rect 61 100 62 101
rect 60 100 61 101
rect 59 100 60 101
rect 58 100 59 101
rect 57 100 58 101
rect 56 100 57 101
rect 55 100 56 101
rect 54 100 55 101
rect 480 101 481 102
rect 479 101 480 102
rect 478 101 479 102
rect 477 101 478 102
rect 476 101 477 102
rect 475 101 476 102
rect 474 101 475 102
rect 473 101 474 102
rect 472 101 473 102
rect 471 101 472 102
rect 470 101 471 102
rect 469 101 470 102
rect 468 101 469 102
rect 467 101 468 102
rect 466 101 467 102
rect 465 101 466 102
rect 464 101 465 102
rect 463 101 464 102
rect 462 101 463 102
rect 265 101 266 102
rect 264 101 265 102
rect 263 101 264 102
rect 262 101 263 102
rect 261 101 262 102
rect 260 101 261 102
rect 259 101 260 102
rect 258 101 259 102
rect 257 101 258 102
rect 256 101 257 102
rect 255 101 256 102
rect 254 101 255 102
rect 253 101 254 102
rect 252 101 253 102
rect 251 101 252 102
rect 250 101 251 102
rect 249 101 250 102
rect 248 101 249 102
rect 247 101 248 102
rect 246 101 247 102
rect 245 101 246 102
rect 244 101 245 102
rect 243 101 244 102
rect 242 101 243 102
rect 241 101 242 102
rect 240 101 241 102
rect 239 101 240 102
rect 238 101 239 102
rect 237 101 238 102
rect 236 101 237 102
rect 235 101 236 102
rect 234 101 235 102
rect 233 101 234 102
rect 232 101 233 102
rect 231 101 232 102
rect 230 101 231 102
rect 229 101 230 102
rect 228 101 229 102
rect 227 101 228 102
rect 226 101 227 102
rect 225 101 226 102
rect 224 101 225 102
rect 223 101 224 102
rect 222 101 223 102
rect 221 101 222 102
rect 220 101 221 102
rect 219 101 220 102
rect 218 101 219 102
rect 217 101 218 102
rect 216 101 217 102
rect 215 101 216 102
rect 214 101 215 102
rect 213 101 214 102
rect 212 101 213 102
rect 211 101 212 102
rect 210 101 211 102
rect 209 101 210 102
rect 208 101 209 102
rect 207 101 208 102
rect 206 101 207 102
rect 205 101 206 102
rect 204 101 205 102
rect 203 101 204 102
rect 202 101 203 102
rect 201 101 202 102
rect 200 101 201 102
rect 199 101 200 102
rect 198 101 199 102
rect 197 101 198 102
rect 196 101 197 102
rect 195 101 196 102
rect 194 101 195 102
rect 193 101 194 102
rect 192 101 193 102
rect 191 101 192 102
rect 190 101 191 102
rect 189 101 190 102
rect 188 101 189 102
rect 187 101 188 102
rect 186 101 187 102
rect 185 101 186 102
rect 184 101 185 102
rect 183 101 184 102
rect 182 101 183 102
rect 160 101 161 102
rect 159 101 160 102
rect 158 101 159 102
rect 157 101 158 102
rect 156 101 157 102
rect 155 101 156 102
rect 154 101 155 102
rect 153 101 154 102
rect 152 101 153 102
rect 151 101 152 102
rect 150 101 151 102
rect 149 101 150 102
rect 148 101 149 102
rect 147 101 148 102
rect 146 101 147 102
rect 145 101 146 102
rect 144 101 145 102
rect 143 101 144 102
rect 142 101 143 102
rect 141 101 142 102
rect 140 101 141 102
rect 139 101 140 102
rect 138 101 139 102
rect 137 101 138 102
rect 136 101 137 102
rect 135 101 136 102
rect 134 101 135 102
rect 133 101 134 102
rect 132 101 133 102
rect 131 101 132 102
rect 130 101 131 102
rect 122 101 123 102
rect 121 101 122 102
rect 120 101 121 102
rect 119 101 120 102
rect 118 101 119 102
rect 117 101 118 102
rect 116 101 117 102
rect 115 101 116 102
rect 114 101 115 102
rect 113 101 114 102
rect 112 101 113 102
rect 111 101 112 102
rect 110 101 111 102
rect 109 101 110 102
rect 108 101 109 102
rect 107 101 108 102
rect 106 101 107 102
rect 105 101 106 102
rect 104 101 105 102
rect 103 101 104 102
rect 102 101 103 102
rect 101 101 102 102
rect 100 101 101 102
rect 99 101 100 102
rect 98 101 99 102
rect 97 101 98 102
rect 96 101 97 102
rect 95 101 96 102
rect 94 101 95 102
rect 93 101 94 102
rect 92 101 93 102
rect 91 101 92 102
rect 90 101 91 102
rect 89 101 90 102
rect 88 101 89 102
rect 87 101 88 102
rect 86 101 87 102
rect 85 101 86 102
rect 84 101 85 102
rect 83 101 84 102
rect 82 101 83 102
rect 81 101 82 102
rect 80 101 81 102
rect 79 101 80 102
rect 78 101 79 102
rect 77 101 78 102
rect 76 101 77 102
rect 72 101 73 102
rect 71 101 72 102
rect 70 101 71 102
rect 69 101 70 102
rect 68 101 69 102
rect 67 101 68 102
rect 66 101 67 102
rect 65 101 66 102
rect 64 101 65 102
rect 63 101 64 102
rect 62 101 63 102
rect 61 101 62 102
rect 60 101 61 102
rect 59 101 60 102
rect 58 101 59 102
rect 57 101 58 102
rect 56 101 57 102
rect 55 101 56 102
rect 54 101 55 102
rect 53 101 54 102
rect 478 102 479 103
rect 477 102 478 103
rect 476 102 477 103
rect 475 102 476 103
rect 474 102 475 103
rect 473 102 474 103
rect 472 102 473 103
rect 471 102 472 103
rect 470 102 471 103
rect 469 102 470 103
rect 468 102 469 103
rect 467 102 468 103
rect 466 102 467 103
rect 465 102 466 103
rect 464 102 465 103
rect 463 102 464 103
rect 462 102 463 103
rect 266 102 267 103
rect 265 102 266 103
rect 264 102 265 103
rect 263 102 264 103
rect 262 102 263 103
rect 261 102 262 103
rect 260 102 261 103
rect 259 102 260 103
rect 258 102 259 103
rect 257 102 258 103
rect 256 102 257 103
rect 255 102 256 103
rect 254 102 255 103
rect 253 102 254 103
rect 252 102 253 103
rect 251 102 252 103
rect 250 102 251 103
rect 249 102 250 103
rect 248 102 249 103
rect 247 102 248 103
rect 246 102 247 103
rect 245 102 246 103
rect 244 102 245 103
rect 243 102 244 103
rect 242 102 243 103
rect 241 102 242 103
rect 240 102 241 103
rect 239 102 240 103
rect 238 102 239 103
rect 237 102 238 103
rect 236 102 237 103
rect 235 102 236 103
rect 234 102 235 103
rect 233 102 234 103
rect 232 102 233 103
rect 231 102 232 103
rect 230 102 231 103
rect 229 102 230 103
rect 228 102 229 103
rect 227 102 228 103
rect 226 102 227 103
rect 225 102 226 103
rect 224 102 225 103
rect 223 102 224 103
rect 222 102 223 103
rect 221 102 222 103
rect 220 102 221 103
rect 219 102 220 103
rect 218 102 219 103
rect 217 102 218 103
rect 216 102 217 103
rect 215 102 216 103
rect 214 102 215 103
rect 213 102 214 103
rect 212 102 213 103
rect 211 102 212 103
rect 210 102 211 103
rect 209 102 210 103
rect 208 102 209 103
rect 207 102 208 103
rect 206 102 207 103
rect 205 102 206 103
rect 204 102 205 103
rect 203 102 204 103
rect 202 102 203 103
rect 201 102 202 103
rect 200 102 201 103
rect 199 102 200 103
rect 198 102 199 103
rect 197 102 198 103
rect 196 102 197 103
rect 195 102 196 103
rect 194 102 195 103
rect 193 102 194 103
rect 192 102 193 103
rect 191 102 192 103
rect 190 102 191 103
rect 189 102 190 103
rect 188 102 189 103
rect 187 102 188 103
rect 186 102 187 103
rect 185 102 186 103
rect 184 102 185 103
rect 183 102 184 103
rect 182 102 183 103
rect 181 102 182 103
rect 160 102 161 103
rect 159 102 160 103
rect 158 102 159 103
rect 157 102 158 103
rect 156 102 157 103
rect 155 102 156 103
rect 154 102 155 103
rect 153 102 154 103
rect 152 102 153 103
rect 151 102 152 103
rect 150 102 151 103
rect 149 102 150 103
rect 148 102 149 103
rect 147 102 148 103
rect 146 102 147 103
rect 145 102 146 103
rect 144 102 145 103
rect 143 102 144 103
rect 142 102 143 103
rect 141 102 142 103
rect 140 102 141 103
rect 139 102 140 103
rect 138 102 139 103
rect 137 102 138 103
rect 136 102 137 103
rect 135 102 136 103
rect 134 102 135 103
rect 133 102 134 103
rect 132 102 133 103
rect 131 102 132 103
rect 130 102 131 103
rect 121 102 122 103
rect 120 102 121 103
rect 119 102 120 103
rect 118 102 119 103
rect 117 102 118 103
rect 116 102 117 103
rect 115 102 116 103
rect 114 102 115 103
rect 113 102 114 103
rect 112 102 113 103
rect 111 102 112 103
rect 110 102 111 103
rect 109 102 110 103
rect 108 102 109 103
rect 107 102 108 103
rect 106 102 107 103
rect 105 102 106 103
rect 104 102 105 103
rect 103 102 104 103
rect 102 102 103 103
rect 101 102 102 103
rect 100 102 101 103
rect 99 102 100 103
rect 98 102 99 103
rect 97 102 98 103
rect 96 102 97 103
rect 95 102 96 103
rect 94 102 95 103
rect 93 102 94 103
rect 92 102 93 103
rect 91 102 92 103
rect 90 102 91 103
rect 89 102 90 103
rect 88 102 89 103
rect 87 102 88 103
rect 86 102 87 103
rect 85 102 86 103
rect 84 102 85 103
rect 83 102 84 103
rect 82 102 83 103
rect 81 102 82 103
rect 80 102 81 103
rect 79 102 80 103
rect 78 102 79 103
rect 77 102 78 103
rect 76 102 77 103
rect 71 102 72 103
rect 70 102 71 103
rect 69 102 70 103
rect 68 102 69 103
rect 67 102 68 103
rect 66 102 67 103
rect 65 102 66 103
rect 64 102 65 103
rect 63 102 64 103
rect 62 102 63 103
rect 61 102 62 103
rect 60 102 61 103
rect 59 102 60 103
rect 58 102 59 103
rect 57 102 58 103
rect 56 102 57 103
rect 55 102 56 103
rect 54 102 55 103
rect 53 102 54 103
rect 52 102 53 103
rect 465 103 466 104
rect 464 103 465 104
rect 463 103 464 104
rect 462 103 463 104
rect 267 103 268 104
rect 266 103 267 104
rect 265 103 266 104
rect 264 103 265 104
rect 263 103 264 104
rect 262 103 263 104
rect 261 103 262 104
rect 260 103 261 104
rect 259 103 260 104
rect 258 103 259 104
rect 257 103 258 104
rect 256 103 257 104
rect 255 103 256 104
rect 254 103 255 104
rect 253 103 254 104
rect 252 103 253 104
rect 251 103 252 104
rect 250 103 251 104
rect 249 103 250 104
rect 248 103 249 104
rect 247 103 248 104
rect 246 103 247 104
rect 245 103 246 104
rect 244 103 245 104
rect 243 103 244 104
rect 242 103 243 104
rect 241 103 242 104
rect 240 103 241 104
rect 239 103 240 104
rect 238 103 239 104
rect 237 103 238 104
rect 236 103 237 104
rect 235 103 236 104
rect 234 103 235 104
rect 233 103 234 104
rect 232 103 233 104
rect 231 103 232 104
rect 230 103 231 104
rect 229 103 230 104
rect 228 103 229 104
rect 227 103 228 104
rect 226 103 227 104
rect 225 103 226 104
rect 224 103 225 104
rect 223 103 224 104
rect 222 103 223 104
rect 221 103 222 104
rect 220 103 221 104
rect 219 103 220 104
rect 218 103 219 104
rect 217 103 218 104
rect 216 103 217 104
rect 215 103 216 104
rect 214 103 215 104
rect 213 103 214 104
rect 212 103 213 104
rect 211 103 212 104
rect 210 103 211 104
rect 209 103 210 104
rect 208 103 209 104
rect 207 103 208 104
rect 206 103 207 104
rect 205 103 206 104
rect 204 103 205 104
rect 203 103 204 104
rect 202 103 203 104
rect 201 103 202 104
rect 200 103 201 104
rect 199 103 200 104
rect 198 103 199 104
rect 197 103 198 104
rect 196 103 197 104
rect 195 103 196 104
rect 194 103 195 104
rect 193 103 194 104
rect 192 103 193 104
rect 191 103 192 104
rect 190 103 191 104
rect 189 103 190 104
rect 188 103 189 104
rect 187 103 188 104
rect 186 103 187 104
rect 185 103 186 104
rect 184 103 185 104
rect 183 103 184 104
rect 182 103 183 104
rect 181 103 182 104
rect 160 103 161 104
rect 159 103 160 104
rect 158 103 159 104
rect 157 103 158 104
rect 156 103 157 104
rect 155 103 156 104
rect 154 103 155 104
rect 153 103 154 104
rect 152 103 153 104
rect 151 103 152 104
rect 150 103 151 104
rect 149 103 150 104
rect 148 103 149 104
rect 147 103 148 104
rect 146 103 147 104
rect 145 103 146 104
rect 144 103 145 104
rect 143 103 144 104
rect 142 103 143 104
rect 141 103 142 104
rect 140 103 141 104
rect 139 103 140 104
rect 138 103 139 104
rect 137 103 138 104
rect 136 103 137 104
rect 135 103 136 104
rect 134 103 135 104
rect 133 103 134 104
rect 132 103 133 104
rect 131 103 132 104
rect 130 103 131 104
rect 120 103 121 104
rect 119 103 120 104
rect 118 103 119 104
rect 117 103 118 104
rect 116 103 117 104
rect 115 103 116 104
rect 114 103 115 104
rect 113 103 114 104
rect 112 103 113 104
rect 111 103 112 104
rect 110 103 111 104
rect 109 103 110 104
rect 108 103 109 104
rect 107 103 108 104
rect 106 103 107 104
rect 105 103 106 104
rect 104 103 105 104
rect 103 103 104 104
rect 102 103 103 104
rect 101 103 102 104
rect 100 103 101 104
rect 99 103 100 104
rect 98 103 99 104
rect 97 103 98 104
rect 96 103 97 104
rect 95 103 96 104
rect 94 103 95 104
rect 93 103 94 104
rect 92 103 93 104
rect 91 103 92 104
rect 90 103 91 104
rect 89 103 90 104
rect 88 103 89 104
rect 87 103 88 104
rect 86 103 87 104
rect 85 103 86 104
rect 84 103 85 104
rect 83 103 84 104
rect 82 103 83 104
rect 81 103 82 104
rect 80 103 81 104
rect 79 103 80 104
rect 78 103 79 104
rect 77 103 78 104
rect 76 103 77 104
rect 71 103 72 104
rect 70 103 71 104
rect 69 103 70 104
rect 68 103 69 104
rect 67 103 68 104
rect 66 103 67 104
rect 65 103 66 104
rect 64 103 65 104
rect 63 103 64 104
rect 62 103 63 104
rect 61 103 62 104
rect 60 103 61 104
rect 59 103 60 104
rect 58 103 59 104
rect 57 103 58 104
rect 56 103 57 104
rect 55 103 56 104
rect 54 103 55 104
rect 53 103 54 104
rect 52 103 53 104
rect 51 103 52 104
rect 463 104 464 105
rect 462 104 463 105
rect 399 104 400 105
rect 398 104 399 105
rect 397 104 398 105
rect 269 104 270 105
rect 268 104 269 105
rect 267 104 268 105
rect 266 104 267 105
rect 265 104 266 105
rect 264 104 265 105
rect 263 104 264 105
rect 262 104 263 105
rect 261 104 262 105
rect 260 104 261 105
rect 259 104 260 105
rect 258 104 259 105
rect 257 104 258 105
rect 256 104 257 105
rect 255 104 256 105
rect 254 104 255 105
rect 253 104 254 105
rect 252 104 253 105
rect 251 104 252 105
rect 250 104 251 105
rect 249 104 250 105
rect 248 104 249 105
rect 247 104 248 105
rect 246 104 247 105
rect 245 104 246 105
rect 244 104 245 105
rect 243 104 244 105
rect 242 104 243 105
rect 241 104 242 105
rect 240 104 241 105
rect 239 104 240 105
rect 238 104 239 105
rect 237 104 238 105
rect 236 104 237 105
rect 235 104 236 105
rect 234 104 235 105
rect 233 104 234 105
rect 232 104 233 105
rect 231 104 232 105
rect 230 104 231 105
rect 229 104 230 105
rect 228 104 229 105
rect 227 104 228 105
rect 226 104 227 105
rect 225 104 226 105
rect 224 104 225 105
rect 223 104 224 105
rect 222 104 223 105
rect 221 104 222 105
rect 220 104 221 105
rect 219 104 220 105
rect 218 104 219 105
rect 217 104 218 105
rect 216 104 217 105
rect 215 104 216 105
rect 214 104 215 105
rect 213 104 214 105
rect 212 104 213 105
rect 211 104 212 105
rect 210 104 211 105
rect 209 104 210 105
rect 208 104 209 105
rect 207 104 208 105
rect 206 104 207 105
rect 205 104 206 105
rect 204 104 205 105
rect 203 104 204 105
rect 202 104 203 105
rect 201 104 202 105
rect 200 104 201 105
rect 199 104 200 105
rect 198 104 199 105
rect 197 104 198 105
rect 196 104 197 105
rect 195 104 196 105
rect 194 104 195 105
rect 193 104 194 105
rect 192 104 193 105
rect 191 104 192 105
rect 190 104 191 105
rect 189 104 190 105
rect 188 104 189 105
rect 187 104 188 105
rect 186 104 187 105
rect 185 104 186 105
rect 184 104 185 105
rect 183 104 184 105
rect 182 104 183 105
rect 181 104 182 105
rect 180 104 181 105
rect 159 104 160 105
rect 158 104 159 105
rect 157 104 158 105
rect 156 104 157 105
rect 155 104 156 105
rect 154 104 155 105
rect 153 104 154 105
rect 152 104 153 105
rect 151 104 152 105
rect 150 104 151 105
rect 149 104 150 105
rect 148 104 149 105
rect 147 104 148 105
rect 146 104 147 105
rect 145 104 146 105
rect 144 104 145 105
rect 143 104 144 105
rect 142 104 143 105
rect 141 104 142 105
rect 140 104 141 105
rect 139 104 140 105
rect 138 104 139 105
rect 137 104 138 105
rect 136 104 137 105
rect 135 104 136 105
rect 134 104 135 105
rect 133 104 134 105
rect 132 104 133 105
rect 131 104 132 105
rect 130 104 131 105
rect 119 104 120 105
rect 118 104 119 105
rect 117 104 118 105
rect 116 104 117 105
rect 115 104 116 105
rect 114 104 115 105
rect 113 104 114 105
rect 112 104 113 105
rect 111 104 112 105
rect 110 104 111 105
rect 109 104 110 105
rect 108 104 109 105
rect 107 104 108 105
rect 106 104 107 105
rect 105 104 106 105
rect 104 104 105 105
rect 103 104 104 105
rect 102 104 103 105
rect 101 104 102 105
rect 100 104 101 105
rect 99 104 100 105
rect 98 104 99 105
rect 97 104 98 105
rect 96 104 97 105
rect 95 104 96 105
rect 94 104 95 105
rect 93 104 94 105
rect 92 104 93 105
rect 91 104 92 105
rect 90 104 91 105
rect 89 104 90 105
rect 88 104 89 105
rect 87 104 88 105
rect 86 104 87 105
rect 85 104 86 105
rect 84 104 85 105
rect 83 104 84 105
rect 82 104 83 105
rect 81 104 82 105
rect 80 104 81 105
rect 79 104 80 105
rect 78 104 79 105
rect 77 104 78 105
rect 76 104 77 105
rect 70 104 71 105
rect 69 104 70 105
rect 68 104 69 105
rect 67 104 68 105
rect 66 104 67 105
rect 65 104 66 105
rect 64 104 65 105
rect 63 104 64 105
rect 62 104 63 105
rect 61 104 62 105
rect 60 104 61 105
rect 59 104 60 105
rect 58 104 59 105
rect 57 104 58 105
rect 56 104 57 105
rect 55 104 56 105
rect 54 104 55 105
rect 53 104 54 105
rect 52 104 53 105
rect 51 104 52 105
rect 50 104 51 105
rect 462 105 463 106
rect 399 105 400 106
rect 398 105 399 106
rect 397 105 398 106
rect 270 105 271 106
rect 269 105 270 106
rect 268 105 269 106
rect 267 105 268 106
rect 266 105 267 106
rect 265 105 266 106
rect 264 105 265 106
rect 263 105 264 106
rect 262 105 263 106
rect 261 105 262 106
rect 260 105 261 106
rect 259 105 260 106
rect 258 105 259 106
rect 257 105 258 106
rect 256 105 257 106
rect 255 105 256 106
rect 254 105 255 106
rect 253 105 254 106
rect 252 105 253 106
rect 251 105 252 106
rect 250 105 251 106
rect 249 105 250 106
rect 248 105 249 106
rect 247 105 248 106
rect 246 105 247 106
rect 245 105 246 106
rect 244 105 245 106
rect 243 105 244 106
rect 242 105 243 106
rect 241 105 242 106
rect 240 105 241 106
rect 239 105 240 106
rect 238 105 239 106
rect 237 105 238 106
rect 236 105 237 106
rect 235 105 236 106
rect 234 105 235 106
rect 233 105 234 106
rect 232 105 233 106
rect 231 105 232 106
rect 230 105 231 106
rect 229 105 230 106
rect 228 105 229 106
rect 227 105 228 106
rect 226 105 227 106
rect 225 105 226 106
rect 224 105 225 106
rect 223 105 224 106
rect 222 105 223 106
rect 221 105 222 106
rect 220 105 221 106
rect 219 105 220 106
rect 218 105 219 106
rect 217 105 218 106
rect 216 105 217 106
rect 215 105 216 106
rect 214 105 215 106
rect 213 105 214 106
rect 212 105 213 106
rect 211 105 212 106
rect 210 105 211 106
rect 209 105 210 106
rect 208 105 209 106
rect 207 105 208 106
rect 206 105 207 106
rect 205 105 206 106
rect 204 105 205 106
rect 203 105 204 106
rect 202 105 203 106
rect 201 105 202 106
rect 200 105 201 106
rect 199 105 200 106
rect 198 105 199 106
rect 197 105 198 106
rect 196 105 197 106
rect 195 105 196 106
rect 194 105 195 106
rect 193 105 194 106
rect 192 105 193 106
rect 191 105 192 106
rect 190 105 191 106
rect 189 105 190 106
rect 188 105 189 106
rect 187 105 188 106
rect 186 105 187 106
rect 185 105 186 106
rect 184 105 185 106
rect 183 105 184 106
rect 182 105 183 106
rect 181 105 182 106
rect 180 105 181 106
rect 179 105 180 106
rect 159 105 160 106
rect 158 105 159 106
rect 157 105 158 106
rect 156 105 157 106
rect 155 105 156 106
rect 154 105 155 106
rect 153 105 154 106
rect 152 105 153 106
rect 151 105 152 106
rect 150 105 151 106
rect 149 105 150 106
rect 148 105 149 106
rect 147 105 148 106
rect 146 105 147 106
rect 145 105 146 106
rect 144 105 145 106
rect 143 105 144 106
rect 142 105 143 106
rect 141 105 142 106
rect 140 105 141 106
rect 139 105 140 106
rect 138 105 139 106
rect 137 105 138 106
rect 136 105 137 106
rect 135 105 136 106
rect 134 105 135 106
rect 133 105 134 106
rect 132 105 133 106
rect 131 105 132 106
rect 130 105 131 106
rect 129 105 130 106
rect 118 105 119 106
rect 117 105 118 106
rect 116 105 117 106
rect 115 105 116 106
rect 114 105 115 106
rect 113 105 114 106
rect 112 105 113 106
rect 111 105 112 106
rect 110 105 111 106
rect 109 105 110 106
rect 108 105 109 106
rect 107 105 108 106
rect 106 105 107 106
rect 105 105 106 106
rect 104 105 105 106
rect 103 105 104 106
rect 102 105 103 106
rect 101 105 102 106
rect 100 105 101 106
rect 99 105 100 106
rect 98 105 99 106
rect 97 105 98 106
rect 96 105 97 106
rect 95 105 96 106
rect 94 105 95 106
rect 93 105 94 106
rect 92 105 93 106
rect 91 105 92 106
rect 90 105 91 106
rect 89 105 90 106
rect 88 105 89 106
rect 87 105 88 106
rect 86 105 87 106
rect 85 105 86 106
rect 84 105 85 106
rect 83 105 84 106
rect 82 105 83 106
rect 81 105 82 106
rect 80 105 81 106
rect 79 105 80 106
rect 78 105 79 106
rect 77 105 78 106
rect 76 105 77 106
rect 70 105 71 106
rect 69 105 70 106
rect 68 105 69 106
rect 67 105 68 106
rect 66 105 67 106
rect 65 105 66 106
rect 64 105 65 106
rect 63 105 64 106
rect 62 105 63 106
rect 61 105 62 106
rect 60 105 61 106
rect 59 105 60 106
rect 58 105 59 106
rect 57 105 58 106
rect 56 105 57 106
rect 55 105 56 106
rect 54 105 55 106
rect 53 105 54 106
rect 52 105 53 106
rect 51 105 52 106
rect 50 105 51 106
rect 49 105 50 106
rect 399 106 400 107
rect 398 106 399 107
rect 397 106 398 107
rect 271 106 272 107
rect 270 106 271 107
rect 269 106 270 107
rect 268 106 269 107
rect 267 106 268 107
rect 266 106 267 107
rect 265 106 266 107
rect 264 106 265 107
rect 263 106 264 107
rect 262 106 263 107
rect 261 106 262 107
rect 260 106 261 107
rect 259 106 260 107
rect 258 106 259 107
rect 257 106 258 107
rect 256 106 257 107
rect 255 106 256 107
rect 254 106 255 107
rect 253 106 254 107
rect 252 106 253 107
rect 251 106 252 107
rect 250 106 251 107
rect 249 106 250 107
rect 248 106 249 107
rect 247 106 248 107
rect 246 106 247 107
rect 245 106 246 107
rect 244 106 245 107
rect 243 106 244 107
rect 242 106 243 107
rect 241 106 242 107
rect 240 106 241 107
rect 239 106 240 107
rect 238 106 239 107
rect 237 106 238 107
rect 236 106 237 107
rect 235 106 236 107
rect 234 106 235 107
rect 233 106 234 107
rect 232 106 233 107
rect 231 106 232 107
rect 230 106 231 107
rect 229 106 230 107
rect 228 106 229 107
rect 227 106 228 107
rect 226 106 227 107
rect 225 106 226 107
rect 224 106 225 107
rect 223 106 224 107
rect 222 106 223 107
rect 221 106 222 107
rect 220 106 221 107
rect 219 106 220 107
rect 218 106 219 107
rect 217 106 218 107
rect 216 106 217 107
rect 215 106 216 107
rect 214 106 215 107
rect 213 106 214 107
rect 212 106 213 107
rect 211 106 212 107
rect 210 106 211 107
rect 209 106 210 107
rect 208 106 209 107
rect 207 106 208 107
rect 206 106 207 107
rect 205 106 206 107
rect 204 106 205 107
rect 203 106 204 107
rect 202 106 203 107
rect 201 106 202 107
rect 200 106 201 107
rect 199 106 200 107
rect 198 106 199 107
rect 197 106 198 107
rect 196 106 197 107
rect 195 106 196 107
rect 194 106 195 107
rect 193 106 194 107
rect 192 106 193 107
rect 191 106 192 107
rect 190 106 191 107
rect 189 106 190 107
rect 188 106 189 107
rect 187 106 188 107
rect 186 106 187 107
rect 185 106 186 107
rect 184 106 185 107
rect 183 106 184 107
rect 182 106 183 107
rect 181 106 182 107
rect 180 106 181 107
rect 179 106 180 107
rect 159 106 160 107
rect 158 106 159 107
rect 157 106 158 107
rect 156 106 157 107
rect 155 106 156 107
rect 154 106 155 107
rect 153 106 154 107
rect 152 106 153 107
rect 151 106 152 107
rect 150 106 151 107
rect 149 106 150 107
rect 148 106 149 107
rect 147 106 148 107
rect 146 106 147 107
rect 145 106 146 107
rect 144 106 145 107
rect 143 106 144 107
rect 142 106 143 107
rect 141 106 142 107
rect 140 106 141 107
rect 139 106 140 107
rect 138 106 139 107
rect 137 106 138 107
rect 136 106 137 107
rect 135 106 136 107
rect 134 106 135 107
rect 133 106 134 107
rect 132 106 133 107
rect 131 106 132 107
rect 130 106 131 107
rect 129 106 130 107
rect 118 106 119 107
rect 117 106 118 107
rect 116 106 117 107
rect 115 106 116 107
rect 114 106 115 107
rect 113 106 114 107
rect 112 106 113 107
rect 111 106 112 107
rect 110 106 111 107
rect 109 106 110 107
rect 108 106 109 107
rect 107 106 108 107
rect 106 106 107 107
rect 105 106 106 107
rect 104 106 105 107
rect 103 106 104 107
rect 102 106 103 107
rect 101 106 102 107
rect 100 106 101 107
rect 99 106 100 107
rect 98 106 99 107
rect 97 106 98 107
rect 96 106 97 107
rect 95 106 96 107
rect 94 106 95 107
rect 93 106 94 107
rect 92 106 93 107
rect 91 106 92 107
rect 90 106 91 107
rect 89 106 90 107
rect 88 106 89 107
rect 87 106 88 107
rect 86 106 87 107
rect 85 106 86 107
rect 84 106 85 107
rect 83 106 84 107
rect 82 106 83 107
rect 81 106 82 107
rect 80 106 81 107
rect 79 106 80 107
rect 78 106 79 107
rect 77 106 78 107
rect 76 106 77 107
rect 75 106 76 107
rect 69 106 70 107
rect 68 106 69 107
rect 67 106 68 107
rect 66 106 67 107
rect 65 106 66 107
rect 64 106 65 107
rect 63 106 64 107
rect 62 106 63 107
rect 61 106 62 107
rect 60 106 61 107
rect 59 106 60 107
rect 58 106 59 107
rect 57 106 58 107
rect 56 106 57 107
rect 55 106 56 107
rect 54 106 55 107
rect 53 106 54 107
rect 52 106 53 107
rect 51 106 52 107
rect 50 106 51 107
rect 49 106 50 107
rect 48 106 49 107
rect 399 107 400 108
rect 398 107 399 108
rect 397 107 398 108
rect 272 107 273 108
rect 271 107 272 108
rect 270 107 271 108
rect 269 107 270 108
rect 268 107 269 108
rect 267 107 268 108
rect 266 107 267 108
rect 265 107 266 108
rect 264 107 265 108
rect 263 107 264 108
rect 262 107 263 108
rect 261 107 262 108
rect 260 107 261 108
rect 259 107 260 108
rect 258 107 259 108
rect 257 107 258 108
rect 256 107 257 108
rect 255 107 256 108
rect 254 107 255 108
rect 253 107 254 108
rect 252 107 253 108
rect 251 107 252 108
rect 250 107 251 108
rect 249 107 250 108
rect 248 107 249 108
rect 247 107 248 108
rect 246 107 247 108
rect 245 107 246 108
rect 244 107 245 108
rect 243 107 244 108
rect 242 107 243 108
rect 241 107 242 108
rect 240 107 241 108
rect 239 107 240 108
rect 238 107 239 108
rect 237 107 238 108
rect 236 107 237 108
rect 235 107 236 108
rect 234 107 235 108
rect 233 107 234 108
rect 232 107 233 108
rect 231 107 232 108
rect 230 107 231 108
rect 229 107 230 108
rect 228 107 229 108
rect 227 107 228 108
rect 226 107 227 108
rect 225 107 226 108
rect 224 107 225 108
rect 223 107 224 108
rect 222 107 223 108
rect 221 107 222 108
rect 220 107 221 108
rect 219 107 220 108
rect 218 107 219 108
rect 217 107 218 108
rect 216 107 217 108
rect 215 107 216 108
rect 214 107 215 108
rect 213 107 214 108
rect 212 107 213 108
rect 211 107 212 108
rect 210 107 211 108
rect 209 107 210 108
rect 208 107 209 108
rect 207 107 208 108
rect 206 107 207 108
rect 205 107 206 108
rect 204 107 205 108
rect 203 107 204 108
rect 202 107 203 108
rect 201 107 202 108
rect 200 107 201 108
rect 199 107 200 108
rect 198 107 199 108
rect 197 107 198 108
rect 196 107 197 108
rect 195 107 196 108
rect 194 107 195 108
rect 193 107 194 108
rect 192 107 193 108
rect 191 107 192 108
rect 190 107 191 108
rect 189 107 190 108
rect 188 107 189 108
rect 187 107 188 108
rect 186 107 187 108
rect 185 107 186 108
rect 184 107 185 108
rect 183 107 184 108
rect 182 107 183 108
rect 181 107 182 108
rect 180 107 181 108
rect 179 107 180 108
rect 178 107 179 108
rect 158 107 159 108
rect 157 107 158 108
rect 156 107 157 108
rect 155 107 156 108
rect 154 107 155 108
rect 153 107 154 108
rect 152 107 153 108
rect 151 107 152 108
rect 150 107 151 108
rect 149 107 150 108
rect 148 107 149 108
rect 147 107 148 108
rect 146 107 147 108
rect 145 107 146 108
rect 144 107 145 108
rect 143 107 144 108
rect 142 107 143 108
rect 141 107 142 108
rect 140 107 141 108
rect 139 107 140 108
rect 138 107 139 108
rect 137 107 138 108
rect 136 107 137 108
rect 135 107 136 108
rect 134 107 135 108
rect 133 107 134 108
rect 132 107 133 108
rect 131 107 132 108
rect 130 107 131 108
rect 129 107 130 108
rect 117 107 118 108
rect 116 107 117 108
rect 115 107 116 108
rect 114 107 115 108
rect 113 107 114 108
rect 112 107 113 108
rect 111 107 112 108
rect 110 107 111 108
rect 109 107 110 108
rect 108 107 109 108
rect 107 107 108 108
rect 106 107 107 108
rect 105 107 106 108
rect 104 107 105 108
rect 103 107 104 108
rect 102 107 103 108
rect 101 107 102 108
rect 100 107 101 108
rect 99 107 100 108
rect 98 107 99 108
rect 97 107 98 108
rect 96 107 97 108
rect 95 107 96 108
rect 94 107 95 108
rect 93 107 94 108
rect 92 107 93 108
rect 91 107 92 108
rect 90 107 91 108
rect 89 107 90 108
rect 88 107 89 108
rect 87 107 88 108
rect 86 107 87 108
rect 85 107 86 108
rect 84 107 85 108
rect 83 107 84 108
rect 82 107 83 108
rect 81 107 82 108
rect 80 107 81 108
rect 79 107 80 108
rect 78 107 79 108
rect 77 107 78 108
rect 76 107 77 108
rect 75 107 76 108
rect 69 107 70 108
rect 68 107 69 108
rect 67 107 68 108
rect 66 107 67 108
rect 65 107 66 108
rect 64 107 65 108
rect 63 107 64 108
rect 62 107 63 108
rect 61 107 62 108
rect 60 107 61 108
rect 59 107 60 108
rect 58 107 59 108
rect 57 107 58 108
rect 56 107 57 108
rect 55 107 56 108
rect 54 107 55 108
rect 53 107 54 108
rect 52 107 53 108
rect 51 107 52 108
rect 50 107 51 108
rect 49 107 50 108
rect 48 107 49 108
rect 47 107 48 108
rect 46 107 47 108
rect 400 108 401 109
rect 399 108 400 109
rect 398 108 399 109
rect 397 108 398 109
rect 273 108 274 109
rect 272 108 273 109
rect 271 108 272 109
rect 270 108 271 109
rect 269 108 270 109
rect 268 108 269 109
rect 267 108 268 109
rect 266 108 267 109
rect 265 108 266 109
rect 264 108 265 109
rect 263 108 264 109
rect 262 108 263 109
rect 261 108 262 109
rect 260 108 261 109
rect 259 108 260 109
rect 258 108 259 109
rect 257 108 258 109
rect 256 108 257 109
rect 255 108 256 109
rect 254 108 255 109
rect 253 108 254 109
rect 252 108 253 109
rect 251 108 252 109
rect 250 108 251 109
rect 249 108 250 109
rect 248 108 249 109
rect 247 108 248 109
rect 246 108 247 109
rect 245 108 246 109
rect 244 108 245 109
rect 243 108 244 109
rect 242 108 243 109
rect 241 108 242 109
rect 240 108 241 109
rect 239 108 240 109
rect 238 108 239 109
rect 237 108 238 109
rect 236 108 237 109
rect 235 108 236 109
rect 234 108 235 109
rect 233 108 234 109
rect 232 108 233 109
rect 231 108 232 109
rect 230 108 231 109
rect 229 108 230 109
rect 228 108 229 109
rect 227 108 228 109
rect 226 108 227 109
rect 225 108 226 109
rect 224 108 225 109
rect 223 108 224 109
rect 222 108 223 109
rect 221 108 222 109
rect 220 108 221 109
rect 219 108 220 109
rect 218 108 219 109
rect 217 108 218 109
rect 216 108 217 109
rect 215 108 216 109
rect 214 108 215 109
rect 213 108 214 109
rect 212 108 213 109
rect 211 108 212 109
rect 210 108 211 109
rect 209 108 210 109
rect 208 108 209 109
rect 207 108 208 109
rect 206 108 207 109
rect 205 108 206 109
rect 204 108 205 109
rect 203 108 204 109
rect 202 108 203 109
rect 201 108 202 109
rect 200 108 201 109
rect 199 108 200 109
rect 198 108 199 109
rect 197 108 198 109
rect 196 108 197 109
rect 195 108 196 109
rect 194 108 195 109
rect 193 108 194 109
rect 192 108 193 109
rect 191 108 192 109
rect 190 108 191 109
rect 189 108 190 109
rect 188 108 189 109
rect 187 108 188 109
rect 186 108 187 109
rect 185 108 186 109
rect 184 108 185 109
rect 183 108 184 109
rect 182 108 183 109
rect 181 108 182 109
rect 180 108 181 109
rect 179 108 180 109
rect 178 108 179 109
rect 177 108 178 109
rect 158 108 159 109
rect 157 108 158 109
rect 156 108 157 109
rect 155 108 156 109
rect 154 108 155 109
rect 153 108 154 109
rect 152 108 153 109
rect 151 108 152 109
rect 150 108 151 109
rect 149 108 150 109
rect 148 108 149 109
rect 147 108 148 109
rect 146 108 147 109
rect 145 108 146 109
rect 144 108 145 109
rect 143 108 144 109
rect 142 108 143 109
rect 141 108 142 109
rect 140 108 141 109
rect 139 108 140 109
rect 138 108 139 109
rect 137 108 138 109
rect 136 108 137 109
rect 135 108 136 109
rect 134 108 135 109
rect 133 108 134 109
rect 132 108 133 109
rect 131 108 132 109
rect 130 108 131 109
rect 129 108 130 109
rect 128 108 129 109
rect 117 108 118 109
rect 116 108 117 109
rect 115 108 116 109
rect 114 108 115 109
rect 113 108 114 109
rect 112 108 113 109
rect 111 108 112 109
rect 110 108 111 109
rect 109 108 110 109
rect 108 108 109 109
rect 107 108 108 109
rect 106 108 107 109
rect 105 108 106 109
rect 104 108 105 109
rect 103 108 104 109
rect 102 108 103 109
rect 101 108 102 109
rect 100 108 101 109
rect 99 108 100 109
rect 98 108 99 109
rect 97 108 98 109
rect 96 108 97 109
rect 95 108 96 109
rect 94 108 95 109
rect 93 108 94 109
rect 92 108 93 109
rect 91 108 92 109
rect 90 108 91 109
rect 89 108 90 109
rect 88 108 89 109
rect 87 108 88 109
rect 86 108 87 109
rect 85 108 86 109
rect 84 108 85 109
rect 83 108 84 109
rect 82 108 83 109
rect 81 108 82 109
rect 80 108 81 109
rect 79 108 80 109
rect 68 108 69 109
rect 67 108 68 109
rect 66 108 67 109
rect 65 108 66 109
rect 64 108 65 109
rect 63 108 64 109
rect 62 108 63 109
rect 61 108 62 109
rect 60 108 61 109
rect 59 108 60 109
rect 58 108 59 109
rect 57 108 58 109
rect 56 108 57 109
rect 55 108 56 109
rect 54 108 55 109
rect 53 108 54 109
rect 52 108 53 109
rect 51 108 52 109
rect 50 108 51 109
rect 49 108 50 109
rect 48 108 49 109
rect 47 108 48 109
rect 46 108 47 109
rect 45 108 46 109
rect 425 109 426 110
rect 424 109 425 110
rect 423 109 424 110
rect 422 109 423 110
rect 421 109 422 110
rect 420 109 421 110
rect 419 109 420 110
rect 418 109 419 110
rect 417 109 418 110
rect 416 109 417 110
rect 415 109 416 110
rect 414 109 415 110
rect 413 109 414 110
rect 412 109 413 110
rect 411 109 412 110
rect 410 109 411 110
rect 409 109 410 110
rect 408 109 409 110
rect 407 109 408 110
rect 406 109 407 110
rect 405 109 406 110
rect 404 109 405 110
rect 403 109 404 110
rect 402 109 403 110
rect 401 109 402 110
rect 400 109 401 110
rect 399 109 400 110
rect 398 109 399 110
rect 397 109 398 110
rect 274 109 275 110
rect 273 109 274 110
rect 272 109 273 110
rect 271 109 272 110
rect 270 109 271 110
rect 269 109 270 110
rect 268 109 269 110
rect 267 109 268 110
rect 266 109 267 110
rect 265 109 266 110
rect 264 109 265 110
rect 263 109 264 110
rect 262 109 263 110
rect 261 109 262 110
rect 260 109 261 110
rect 259 109 260 110
rect 258 109 259 110
rect 257 109 258 110
rect 256 109 257 110
rect 255 109 256 110
rect 254 109 255 110
rect 253 109 254 110
rect 252 109 253 110
rect 251 109 252 110
rect 250 109 251 110
rect 249 109 250 110
rect 248 109 249 110
rect 247 109 248 110
rect 246 109 247 110
rect 245 109 246 110
rect 244 109 245 110
rect 243 109 244 110
rect 242 109 243 110
rect 241 109 242 110
rect 240 109 241 110
rect 239 109 240 110
rect 238 109 239 110
rect 237 109 238 110
rect 236 109 237 110
rect 235 109 236 110
rect 234 109 235 110
rect 233 109 234 110
rect 232 109 233 110
rect 231 109 232 110
rect 230 109 231 110
rect 229 109 230 110
rect 228 109 229 110
rect 227 109 228 110
rect 226 109 227 110
rect 225 109 226 110
rect 224 109 225 110
rect 223 109 224 110
rect 222 109 223 110
rect 221 109 222 110
rect 220 109 221 110
rect 219 109 220 110
rect 218 109 219 110
rect 217 109 218 110
rect 216 109 217 110
rect 215 109 216 110
rect 214 109 215 110
rect 213 109 214 110
rect 212 109 213 110
rect 211 109 212 110
rect 210 109 211 110
rect 209 109 210 110
rect 208 109 209 110
rect 207 109 208 110
rect 206 109 207 110
rect 205 109 206 110
rect 204 109 205 110
rect 203 109 204 110
rect 202 109 203 110
rect 201 109 202 110
rect 200 109 201 110
rect 199 109 200 110
rect 198 109 199 110
rect 197 109 198 110
rect 196 109 197 110
rect 195 109 196 110
rect 194 109 195 110
rect 193 109 194 110
rect 192 109 193 110
rect 191 109 192 110
rect 190 109 191 110
rect 189 109 190 110
rect 188 109 189 110
rect 187 109 188 110
rect 186 109 187 110
rect 185 109 186 110
rect 184 109 185 110
rect 183 109 184 110
rect 182 109 183 110
rect 181 109 182 110
rect 180 109 181 110
rect 179 109 180 110
rect 178 109 179 110
rect 177 109 178 110
rect 158 109 159 110
rect 157 109 158 110
rect 156 109 157 110
rect 155 109 156 110
rect 154 109 155 110
rect 153 109 154 110
rect 152 109 153 110
rect 151 109 152 110
rect 150 109 151 110
rect 149 109 150 110
rect 148 109 149 110
rect 147 109 148 110
rect 146 109 147 110
rect 145 109 146 110
rect 144 109 145 110
rect 143 109 144 110
rect 142 109 143 110
rect 141 109 142 110
rect 140 109 141 110
rect 139 109 140 110
rect 138 109 139 110
rect 137 109 138 110
rect 136 109 137 110
rect 135 109 136 110
rect 134 109 135 110
rect 133 109 134 110
rect 132 109 133 110
rect 131 109 132 110
rect 130 109 131 110
rect 129 109 130 110
rect 128 109 129 110
rect 118 109 119 110
rect 117 109 118 110
rect 116 109 117 110
rect 115 109 116 110
rect 114 109 115 110
rect 113 109 114 110
rect 112 109 113 110
rect 111 109 112 110
rect 110 109 111 110
rect 109 109 110 110
rect 108 109 109 110
rect 107 109 108 110
rect 106 109 107 110
rect 105 109 106 110
rect 104 109 105 110
rect 103 109 104 110
rect 102 109 103 110
rect 101 109 102 110
rect 100 109 101 110
rect 99 109 100 110
rect 98 109 99 110
rect 97 109 98 110
rect 96 109 97 110
rect 95 109 96 110
rect 94 109 95 110
rect 93 109 94 110
rect 92 109 93 110
rect 91 109 92 110
rect 90 109 91 110
rect 89 109 90 110
rect 88 109 89 110
rect 87 109 88 110
rect 86 109 87 110
rect 85 109 86 110
rect 84 109 85 110
rect 83 109 84 110
rect 82 109 83 110
rect 67 109 68 110
rect 66 109 67 110
rect 65 109 66 110
rect 64 109 65 110
rect 63 109 64 110
rect 62 109 63 110
rect 61 109 62 110
rect 60 109 61 110
rect 59 109 60 110
rect 58 109 59 110
rect 57 109 58 110
rect 56 109 57 110
rect 55 109 56 110
rect 54 109 55 110
rect 53 109 54 110
rect 52 109 53 110
rect 51 109 52 110
rect 50 109 51 110
rect 49 109 50 110
rect 48 109 49 110
rect 47 109 48 110
rect 46 109 47 110
rect 45 109 46 110
rect 44 109 45 110
rect 43 109 44 110
rect 431 110 432 111
rect 430 110 431 111
rect 429 110 430 111
rect 428 110 429 111
rect 427 110 428 111
rect 426 110 427 111
rect 425 110 426 111
rect 424 110 425 111
rect 423 110 424 111
rect 422 110 423 111
rect 421 110 422 111
rect 420 110 421 111
rect 419 110 420 111
rect 418 110 419 111
rect 417 110 418 111
rect 416 110 417 111
rect 415 110 416 111
rect 414 110 415 111
rect 413 110 414 111
rect 412 110 413 111
rect 411 110 412 111
rect 410 110 411 111
rect 409 110 410 111
rect 408 110 409 111
rect 407 110 408 111
rect 406 110 407 111
rect 405 110 406 111
rect 404 110 405 111
rect 403 110 404 111
rect 402 110 403 111
rect 401 110 402 111
rect 400 110 401 111
rect 399 110 400 111
rect 398 110 399 111
rect 397 110 398 111
rect 275 110 276 111
rect 274 110 275 111
rect 273 110 274 111
rect 272 110 273 111
rect 271 110 272 111
rect 270 110 271 111
rect 269 110 270 111
rect 268 110 269 111
rect 267 110 268 111
rect 266 110 267 111
rect 265 110 266 111
rect 264 110 265 111
rect 263 110 264 111
rect 262 110 263 111
rect 261 110 262 111
rect 260 110 261 111
rect 259 110 260 111
rect 258 110 259 111
rect 257 110 258 111
rect 256 110 257 111
rect 255 110 256 111
rect 254 110 255 111
rect 253 110 254 111
rect 252 110 253 111
rect 251 110 252 111
rect 250 110 251 111
rect 249 110 250 111
rect 248 110 249 111
rect 247 110 248 111
rect 246 110 247 111
rect 245 110 246 111
rect 244 110 245 111
rect 243 110 244 111
rect 242 110 243 111
rect 241 110 242 111
rect 240 110 241 111
rect 239 110 240 111
rect 238 110 239 111
rect 237 110 238 111
rect 236 110 237 111
rect 235 110 236 111
rect 234 110 235 111
rect 233 110 234 111
rect 232 110 233 111
rect 231 110 232 111
rect 230 110 231 111
rect 229 110 230 111
rect 228 110 229 111
rect 227 110 228 111
rect 226 110 227 111
rect 225 110 226 111
rect 224 110 225 111
rect 223 110 224 111
rect 222 110 223 111
rect 221 110 222 111
rect 220 110 221 111
rect 219 110 220 111
rect 218 110 219 111
rect 217 110 218 111
rect 216 110 217 111
rect 215 110 216 111
rect 214 110 215 111
rect 213 110 214 111
rect 212 110 213 111
rect 211 110 212 111
rect 210 110 211 111
rect 209 110 210 111
rect 208 110 209 111
rect 207 110 208 111
rect 206 110 207 111
rect 205 110 206 111
rect 204 110 205 111
rect 203 110 204 111
rect 202 110 203 111
rect 201 110 202 111
rect 200 110 201 111
rect 199 110 200 111
rect 198 110 199 111
rect 197 110 198 111
rect 196 110 197 111
rect 195 110 196 111
rect 194 110 195 111
rect 193 110 194 111
rect 192 110 193 111
rect 191 110 192 111
rect 190 110 191 111
rect 189 110 190 111
rect 188 110 189 111
rect 187 110 188 111
rect 186 110 187 111
rect 185 110 186 111
rect 184 110 185 111
rect 183 110 184 111
rect 182 110 183 111
rect 181 110 182 111
rect 180 110 181 111
rect 179 110 180 111
rect 178 110 179 111
rect 177 110 178 111
rect 176 110 177 111
rect 157 110 158 111
rect 156 110 157 111
rect 155 110 156 111
rect 154 110 155 111
rect 153 110 154 111
rect 152 110 153 111
rect 151 110 152 111
rect 150 110 151 111
rect 149 110 150 111
rect 148 110 149 111
rect 147 110 148 111
rect 146 110 147 111
rect 145 110 146 111
rect 144 110 145 111
rect 143 110 144 111
rect 142 110 143 111
rect 141 110 142 111
rect 140 110 141 111
rect 139 110 140 111
rect 138 110 139 111
rect 137 110 138 111
rect 136 110 137 111
rect 135 110 136 111
rect 134 110 135 111
rect 133 110 134 111
rect 132 110 133 111
rect 131 110 132 111
rect 130 110 131 111
rect 129 110 130 111
rect 128 110 129 111
rect 118 110 119 111
rect 117 110 118 111
rect 116 110 117 111
rect 115 110 116 111
rect 114 110 115 111
rect 113 110 114 111
rect 112 110 113 111
rect 111 110 112 111
rect 110 110 111 111
rect 109 110 110 111
rect 108 110 109 111
rect 107 110 108 111
rect 106 110 107 111
rect 105 110 106 111
rect 104 110 105 111
rect 103 110 104 111
rect 102 110 103 111
rect 101 110 102 111
rect 100 110 101 111
rect 99 110 100 111
rect 98 110 99 111
rect 97 110 98 111
rect 96 110 97 111
rect 95 110 96 111
rect 94 110 95 111
rect 93 110 94 111
rect 92 110 93 111
rect 91 110 92 111
rect 90 110 91 111
rect 89 110 90 111
rect 88 110 89 111
rect 87 110 88 111
rect 86 110 87 111
rect 85 110 86 111
rect 84 110 85 111
rect 83 110 84 111
rect 67 110 68 111
rect 66 110 67 111
rect 65 110 66 111
rect 64 110 65 111
rect 63 110 64 111
rect 62 110 63 111
rect 61 110 62 111
rect 60 110 61 111
rect 59 110 60 111
rect 58 110 59 111
rect 57 110 58 111
rect 56 110 57 111
rect 55 110 56 111
rect 54 110 55 111
rect 53 110 54 111
rect 52 110 53 111
rect 51 110 52 111
rect 50 110 51 111
rect 49 110 50 111
rect 48 110 49 111
rect 47 110 48 111
rect 46 110 47 111
rect 45 110 46 111
rect 44 110 45 111
rect 43 110 44 111
rect 42 110 43 111
rect 434 111 435 112
rect 433 111 434 112
rect 432 111 433 112
rect 431 111 432 112
rect 430 111 431 112
rect 429 111 430 112
rect 428 111 429 112
rect 427 111 428 112
rect 426 111 427 112
rect 425 111 426 112
rect 424 111 425 112
rect 423 111 424 112
rect 422 111 423 112
rect 421 111 422 112
rect 420 111 421 112
rect 419 111 420 112
rect 418 111 419 112
rect 417 111 418 112
rect 416 111 417 112
rect 415 111 416 112
rect 414 111 415 112
rect 413 111 414 112
rect 412 111 413 112
rect 411 111 412 112
rect 410 111 411 112
rect 409 111 410 112
rect 408 111 409 112
rect 407 111 408 112
rect 406 111 407 112
rect 405 111 406 112
rect 404 111 405 112
rect 403 111 404 112
rect 402 111 403 112
rect 401 111 402 112
rect 400 111 401 112
rect 399 111 400 112
rect 398 111 399 112
rect 397 111 398 112
rect 276 111 277 112
rect 275 111 276 112
rect 274 111 275 112
rect 273 111 274 112
rect 272 111 273 112
rect 271 111 272 112
rect 270 111 271 112
rect 269 111 270 112
rect 268 111 269 112
rect 267 111 268 112
rect 266 111 267 112
rect 265 111 266 112
rect 264 111 265 112
rect 263 111 264 112
rect 262 111 263 112
rect 261 111 262 112
rect 260 111 261 112
rect 259 111 260 112
rect 258 111 259 112
rect 257 111 258 112
rect 256 111 257 112
rect 255 111 256 112
rect 254 111 255 112
rect 253 111 254 112
rect 252 111 253 112
rect 251 111 252 112
rect 250 111 251 112
rect 249 111 250 112
rect 248 111 249 112
rect 247 111 248 112
rect 246 111 247 112
rect 245 111 246 112
rect 244 111 245 112
rect 243 111 244 112
rect 242 111 243 112
rect 241 111 242 112
rect 240 111 241 112
rect 239 111 240 112
rect 238 111 239 112
rect 237 111 238 112
rect 236 111 237 112
rect 235 111 236 112
rect 234 111 235 112
rect 233 111 234 112
rect 232 111 233 112
rect 231 111 232 112
rect 230 111 231 112
rect 229 111 230 112
rect 228 111 229 112
rect 227 111 228 112
rect 226 111 227 112
rect 225 111 226 112
rect 224 111 225 112
rect 223 111 224 112
rect 222 111 223 112
rect 221 111 222 112
rect 220 111 221 112
rect 219 111 220 112
rect 218 111 219 112
rect 217 111 218 112
rect 216 111 217 112
rect 215 111 216 112
rect 214 111 215 112
rect 213 111 214 112
rect 212 111 213 112
rect 211 111 212 112
rect 210 111 211 112
rect 209 111 210 112
rect 208 111 209 112
rect 207 111 208 112
rect 206 111 207 112
rect 205 111 206 112
rect 204 111 205 112
rect 203 111 204 112
rect 202 111 203 112
rect 201 111 202 112
rect 200 111 201 112
rect 199 111 200 112
rect 198 111 199 112
rect 197 111 198 112
rect 196 111 197 112
rect 195 111 196 112
rect 194 111 195 112
rect 193 111 194 112
rect 192 111 193 112
rect 191 111 192 112
rect 190 111 191 112
rect 189 111 190 112
rect 188 111 189 112
rect 187 111 188 112
rect 186 111 187 112
rect 185 111 186 112
rect 184 111 185 112
rect 183 111 184 112
rect 182 111 183 112
rect 181 111 182 112
rect 180 111 181 112
rect 179 111 180 112
rect 178 111 179 112
rect 177 111 178 112
rect 176 111 177 112
rect 157 111 158 112
rect 156 111 157 112
rect 155 111 156 112
rect 154 111 155 112
rect 153 111 154 112
rect 152 111 153 112
rect 151 111 152 112
rect 150 111 151 112
rect 149 111 150 112
rect 148 111 149 112
rect 147 111 148 112
rect 146 111 147 112
rect 145 111 146 112
rect 144 111 145 112
rect 143 111 144 112
rect 142 111 143 112
rect 141 111 142 112
rect 140 111 141 112
rect 139 111 140 112
rect 138 111 139 112
rect 137 111 138 112
rect 136 111 137 112
rect 135 111 136 112
rect 134 111 135 112
rect 133 111 134 112
rect 132 111 133 112
rect 131 111 132 112
rect 130 111 131 112
rect 129 111 130 112
rect 128 111 129 112
rect 127 111 128 112
rect 119 111 120 112
rect 118 111 119 112
rect 117 111 118 112
rect 116 111 117 112
rect 115 111 116 112
rect 114 111 115 112
rect 113 111 114 112
rect 112 111 113 112
rect 111 111 112 112
rect 110 111 111 112
rect 109 111 110 112
rect 108 111 109 112
rect 107 111 108 112
rect 106 111 107 112
rect 105 111 106 112
rect 104 111 105 112
rect 103 111 104 112
rect 102 111 103 112
rect 101 111 102 112
rect 100 111 101 112
rect 99 111 100 112
rect 98 111 99 112
rect 97 111 98 112
rect 96 111 97 112
rect 95 111 96 112
rect 94 111 95 112
rect 93 111 94 112
rect 92 111 93 112
rect 91 111 92 112
rect 90 111 91 112
rect 89 111 90 112
rect 88 111 89 112
rect 87 111 88 112
rect 86 111 87 112
rect 85 111 86 112
rect 84 111 85 112
rect 66 111 67 112
rect 65 111 66 112
rect 64 111 65 112
rect 63 111 64 112
rect 62 111 63 112
rect 61 111 62 112
rect 60 111 61 112
rect 59 111 60 112
rect 58 111 59 112
rect 57 111 58 112
rect 56 111 57 112
rect 55 111 56 112
rect 54 111 55 112
rect 53 111 54 112
rect 52 111 53 112
rect 51 111 52 112
rect 50 111 51 112
rect 49 111 50 112
rect 48 111 49 112
rect 47 111 48 112
rect 46 111 47 112
rect 45 111 46 112
rect 44 111 45 112
rect 43 111 44 112
rect 42 111 43 112
rect 41 111 42 112
rect 40 111 41 112
rect 436 112 437 113
rect 435 112 436 113
rect 434 112 435 113
rect 433 112 434 113
rect 432 112 433 113
rect 431 112 432 113
rect 430 112 431 113
rect 429 112 430 113
rect 428 112 429 113
rect 427 112 428 113
rect 426 112 427 113
rect 425 112 426 113
rect 424 112 425 113
rect 423 112 424 113
rect 422 112 423 113
rect 421 112 422 113
rect 420 112 421 113
rect 419 112 420 113
rect 418 112 419 113
rect 417 112 418 113
rect 416 112 417 113
rect 415 112 416 113
rect 414 112 415 113
rect 413 112 414 113
rect 412 112 413 113
rect 411 112 412 113
rect 410 112 411 113
rect 409 112 410 113
rect 408 112 409 113
rect 407 112 408 113
rect 406 112 407 113
rect 405 112 406 113
rect 404 112 405 113
rect 403 112 404 113
rect 402 112 403 113
rect 401 112 402 113
rect 400 112 401 113
rect 399 112 400 113
rect 398 112 399 113
rect 397 112 398 113
rect 277 112 278 113
rect 276 112 277 113
rect 275 112 276 113
rect 274 112 275 113
rect 273 112 274 113
rect 272 112 273 113
rect 271 112 272 113
rect 270 112 271 113
rect 269 112 270 113
rect 268 112 269 113
rect 267 112 268 113
rect 266 112 267 113
rect 265 112 266 113
rect 264 112 265 113
rect 263 112 264 113
rect 262 112 263 113
rect 261 112 262 113
rect 260 112 261 113
rect 259 112 260 113
rect 258 112 259 113
rect 257 112 258 113
rect 256 112 257 113
rect 255 112 256 113
rect 254 112 255 113
rect 253 112 254 113
rect 252 112 253 113
rect 251 112 252 113
rect 250 112 251 113
rect 249 112 250 113
rect 248 112 249 113
rect 247 112 248 113
rect 246 112 247 113
rect 245 112 246 113
rect 244 112 245 113
rect 243 112 244 113
rect 242 112 243 113
rect 241 112 242 113
rect 240 112 241 113
rect 239 112 240 113
rect 238 112 239 113
rect 237 112 238 113
rect 236 112 237 113
rect 235 112 236 113
rect 234 112 235 113
rect 233 112 234 113
rect 232 112 233 113
rect 231 112 232 113
rect 230 112 231 113
rect 229 112 230 113
rect 228 112 229 113
rect 227 112 228 113
rect 226 112 227 113
rect 225 112 226 113
rect 224 112 225 113
rect 223 112 224 113
rect 222 112 223 113
rect 221 112 222 113
rect 220 112 221 113
rect 219 112 220 113
rect 218 112 219 113
rect 217 112 218 113
rect 216 112 217 113
rect 215 112 216 113
rect 214 112 215 113
rect 213 112 214 113
rect 212 112 213 113
rect 211 112 212 113
rect 210 112 211 113
rect 209 112 210 113
rect 208 112 209 113
rect 207 112 208 113
rect 206 112 207 113
rect 205 112 206 113
rect 204 112 205 113
rect 203 112 204 113
rect 202 112 203 113
rect 201 112 202 113
rect 200 112 201 113
rect 199 112 200 113
rect 198 112 199 113
rect 197 112 198 113
rect 196 112 197 113
rect 195 112 196 113
rect 194 112 195 113
rect 193 112 194 113
rect 192 112 193 113
rect 191 112 192 113
rect 190 112 191 113
rect 189 112 190 113
rect 188 112 189 113
rect 187 112 188 113
rect 186 112 187 113
rect 185 112 186 113
rect 184 112 185 113
rect 183 112 184 113
rect 182 112 183 113
rect 181 112 182 113
rect 180 112 181 113
rect 179 112 180 113
rect 178 112 179 113
rect 177 112 178 113
rect 176 112 177 113
rect 175 112 176 113
rect 157 112 158 113
rect 156 112 157 113
rect 155 112 156 113
rect 154 112 155 113
rect 153 112 154 113
rect 152 112 153 113
rect 151 112 152 113
rect 150 112 151 113
rect 149 112 150 113
rect 148 112 149 113
rect 147 112 148 113
rect 146 112 147 113
rect 145 112 146 113
rect 144 112 145 113
rect 143 112 144 113
rect 142 112 143 113
rect 141 112 142 113
rect 140 112 141 113
rect 139 112 140 113
rect 138 112 139 113
rect 137 112 138 113
rect 136 112 137 113
rect 135 112 136 113
rect 134 112 135 113
rect 133 112 134 113
rect 132 112 133 113
rect 131 112 132 113
rect 130 112 131 113
rect 129 112 130 113
rect 128 112 129 113
rect 127 112 128 113
rect 120 112 121 113
rect 119 112 120 113
rect 118 112 119 113
rect 117 112 118 113
rect 116 112 117 113
rect 115 112 116 113
rect 114 112 115 113
rect 113 112 114 113
rect 112 112 113 113
rect 111 112 112 113
rect 110 112 111 113
rect 109 112 110 113
rect 108 112 109 113
rect 107 112 108 113
rect 106 112 107 113
rect 105 112 106 113
rect 104 112 105 113
rect 103 112 104 113
rect 102 112 103 113
rect 101 112 102 113
rect 100 112 101 113
rect 99 112 100 113
rect 98 112 99 113
rect 97 112 98 113
rect 96 112 97 113
rect 95 112 96 113
rect 94 112 95 113
rect 93 112 94 113
rect 92 112 93 113
rect 91 112 92 113
rect 90 112 91 113
rect 89 112 90 113
rect 88 112 89 113
rect 87 112 88 113
rect 86 112 87 113
rect 85 112 86 113
rect 84 112 85 113
rect 66 112 67 113
rect 65 112 66 113
rect 64 112 65 113
rect 63 112 64 113
rect 62 112 63 113
rect 61 112 62 113
rect 60 112 61 113
rect 59 112 60 113
rect 58 112 59 113
rect 57 112 58 113
rect 56 112 57 113
rect 55 112 56 113
rect 54 112 55 113
rect 53 112 54 113
rect 52 112 53 113
rect 51 112 52 113
rect 50 112 51 113
rect 49 112 50 113
rect 48 112 49 113
rect 47 112 48 113
rect 46 112 47 113
rect 45 112 46 113
rect 44 112 45 113
rect 43 112 44 113
rect 42 112 43 113
rect 41 112 42 113
rect 40 112 41 113
rect 39 112 40 113
rect 482 113 483 114
rect 462 113 463 114
rect 437 113 438 114
rect 436 113 437 114
rect 435 113 436 114
rect 434 113 435 114
rect 433 113 434 114
rect 432 113 433 114
rect 431 113 432 114
rect 430 113 431 114
rect 429 113 430 114
rect 428 113 429 114
rect 427 113 428 114
rect 426 113 427 114
rect 425 113 426 114
rect 424 113 425 114
rect 423 113 424 114
rect 422 113 423 114
rect 421 113 422 114
rect 420 113 421 114
rect 419 113 420 114
rect 418 113 419 114
rect 417 113 418 114
rect 416 113 417 114
rect 415 113 416 114
rect 414 113 415 114
rect 413 113 414 114
rect 412 113 413 114
rect 411 113 412 114
rect 410 113 411 114
rect 409 113 410 114
rect 408 113 409 114
rect 407 113 408 114
rect 406 113 407 114
rect 405 113 406 114
rect 404 113 405 114
rect 403 113 404 114
rect 402 113 403 114
rect 401 113 402 114
rect 400 113 401 114
rect 399 113 400 114
rect 398 113 399 114
rect 397 113 398 114
rect 278 113 279 114
rect 277 113 278 114
rect 276 113 277 114
rect 275 113 276 114
rect 274 113 275 114
rect 273 113 274 114
rect 272 113 273 114
rect 271 113 272 114
rect 270 113 271 114
rect 269 113 270 114
rect 268 113 269 114
rect 267 113 268 114
rect 266 113 267 114
rect 265 113 266 114
rect 264 113 265 114
rect 263 113 264 114
rect 262 113 263 114
rect 261 113 262 114
rect 260 113 261 114
rect 259 113 260 114
rect 258 113 259 114
rect 257 113 258 114
rect 256 113 257 114
rect 255 113 256 114
rect 254 113 255 114
rect 253 113 254 114
rect 252 113 253 114
rect 251 113 252 114
rect 250 113 251 114
rect 249 113 250 114
rect 248 113 249 114
rect 247 113 248 114
rect 246 113 247 114
rect 245 113 246 114
rect 244 113 245 114
rect 243 113 244 114
rect 242 113 243 114
rect 241 113 242 114
rect 240 113 241 114
rect 239 113 240 114
rect 238 113 239 114
rect 237 113 238 114
rect 236 113 237 114
rect 235 113 236 114
rect 234 113 235 114
rect 233 113 234 114
rect 232 113 233 114
rect 231 113 232 114
rect 230 113 231 114
rect 229 113 230 114
rect 228 113 229 114
rect 227 113 228 114
rect 226 113 227 114
rect 225 113 226 114
rect 224 113 225 114
rect 223 113 224 114
rect 222 113 223 114
rect 221 113 222 114
rect 220 113 221 114
rect 219 113 220 114
rect 218 113 219 114
rect 217 113 218 114
rect 216 113 217 114
rect 215 113 216 114
rect 214 113 215 114
rect 213 113 214 114
rect 212 113 213 114
rect 211 113 212 114
rect 210 113 211 114
rect 209 113 210 114
rect 208 113 209 114
rect 207 113 208 114
rect 206 113 207 114
rect 205 113 206 114
rect 204 113 205 114
rect 203 113 204 114
rect 202 113 203 114
rect 201 113 202 114
rect 200 113 201 114
rect 199 113 200 114
rect 198 113 199 114
rect 197 113 198 114
rect 196 113 197 114
rect 195 113 196 114
rect 194 113 195 114
rect 193 113 194 114
rect 192 113 193 114
rect 191 113 192 114
rect 190 113 191 114
rect 189 113 190 114
rect 188 113 189 114
rect 187 113 188 114
rect 186 113 187 114
rect 185 113 186 114
rect 184 113 185 114
rect 183 113 184 114
rect 182 113 183 114
rect 181 113 182 114
rect 180 113 181 114
rect 179 113 180 114
rect 178 113 179 114
rect 177 113 178 114
rect 176 113 177 114
rect 175 113 176 114
rect 157 113 158 114
rect 156 113 157 114
rect 155 113 156 114
rect 154 113 155 114
rect 153 113 154 114
rect 152 113 153 114
rect 151 113 152 114
rect 150 113 151 114
rect 149 113 150 114
rect 148 113 149 114
rect 147 113 148 114
rect 146 113 147 114
rect 145 113 146 114
rect 144 113 145 114
rect 143 113 144 114
rect 142 113 143 114
rect 141 113 142 114
rect 140 113 141 114
rect 139 113 140 114
rect 138 113 139 114
rect 137 113 138 114
rect 136 113 137 114
rect 135 113 136 114
rect 134 113 135 114
rect 133 113 134 114
rect 132 113 133 114
rect 131 113 132 114
rect 130 113 131 114
rect 129 113 130 114
rect 128 113 129 114
rect 127 113 128 114
rect 126 113 127 114
rect 125 113 126 114
rect 122 113 123 114
rect 121 113 122 114
rect 120 113 121 114
rect 119 113 120 114
rect 118 113 119 114
rect 117 113 118 114
rect 116 113 117 114
rect 115 113 116 114
rect 114 113 115 114
rect 113 113 114 114
rect 112 113 113 114
rect 111 113 112 114
rect 110 113 111 114
rect 109 113 110 114
rect 108 113 109 114
rect 107 113 108 114
rect 106 113 107 114
rect 105 113 106 114
rect 104 113 105 114
rect 103 113 104 114
rect 102 113 103 114
rect 101 113 102 114
rect 100 113 101 114
rect 99 113 100 114
rect 98 113 99 114
rect 97 113 98 114
rect 96 113 97 114
rect 95 113 96 114
rect 94 113 95 114
rect 93 113 94 114
rect 92 113 93 114
rect 91 113 92 114
rect 90 113 91 114
rect 89 113 90 114
rect 88 113 89 114
rect 87 113 88 114
rect 86 113 87 114
rect 85 113 86 114
rect 84 113 85 114
rect 83 113 84 114
rect 65 113 66 114
rect 64 113 65 114
rect 63 113 64 114
rect 62 113 63 114
rect 61 113 62 114
rect 60 113 61 114
rect 59 113 60 114
rect 58 113 59 114
rect 57 113 58 114
rect 56 113 57 114
rect 55 113 56 114
rect 54 113 55 114
rect 53 113 54 114
rect 52 113 53 114
rect 51 113 52 114
rect 50 113 51 114
rect 49 113 50 114
rect 48 113 49 114
rect 47 113 48 114
rect 46 113 47 114
rect 45 113 46 114
rect 44 113 45 114
rect 43 113 44 114
rect 42 113 43 114
rect 41 113 42 114
rect 40 113 41 114
rect 39 113 40 114
rect 38 113 39 114
rect 482 114 483 115
rect 462 114 463 115
rect 438 114 439 115
rect 437 114 438 115
rect 436 114 437 115
rect 435 114 436 115
rect 434 114 435 115
rect 433 114 434 115
rect 432 114 433 115
rect 431 114 432 115
rect 430 114 431 115
rect 429 114 430 115
rect 428 114 429 115
rect 427 114 428 115
rect 426 114 427 115
rect 425 114 426 115
rect 424 114 425 115
rect 423 114 424 115
rect 422 114 423 115
rect 421 114 422 115
rect 420 114 421 115
rect 419 114 420 115
rect 418 114 419 115
rect 417 114 418 115
rect 416 114 417 115
rect 415 114 416 115
rect 414 114 415 115
rect 413 114 414 115
rect 412 114 413 115
rect 411 114 412 115
rect 410 114 411 115
rect 409 114 410 115
rect 408 114 409 115
rect 407 114 408 115
rect 406 114 407 115
rect 405 114 406 115
rect 404 114 405 115
rect 403 114 404 115
rect 402 114 403 115
rect 401 114 402 115
rect 400 114 401 115
rect 399 114 400 115
rect 398 114 399 115
rect 397 114 398 115
rect 279 114 280 115
rect 278 114 279 115
rect 277 114 278 115
rect 276 114 277 115
rect 275 114 276 115
rect 274 114 275 115
rect 273 114 274 115
rect 272 114 273 115
rect 271 114 272 115
rect 270 114 271 115
rect 269 114 270 115
rect 268 114 269 115
rect 267 114 268 115
rect 266 114 267 115
rect 265 114 266 115
rect 264 114 265 115
rect 263 114 264 115
rect 262 114 263 115
rect 261 114 262 115
rect 260 114 261 115
rect 259 114 260 115
rect 258 114 259 115
rect 257 114 258 115
rect 256 114 257 115
rect 255 114 256 115
rect 254 114 255 115
rect 253 114 254 115
rect 252 114 253 115
rect 251 114 252 115
rect 250 114 251 115
rect 249 114 250 115
rect 248 114 249 115
rect 247 114 248 115
rect 246 114 247 115
rect 245 114 246 115
rect 244 114 245 115
rect 243 114 244 115
rect 242 114 243 115
rect 241 114 242 115
rect 240 114 241 115
rect 239 114 240 115
rect 238 114 239 115
rect 237 114 238 115
rect 236 114 237 115
rect 235 114 236 115
rect 234 114 235 115
rect 233 114 234 115
rect 232 114 233 115
rect 231 114 232 115
rect 230 114 231 115
rect 229 114 230 115
rect 228 114 229 115
rect 227 114 228 115
rect 226 114 227 115
rect 225 114 226 115
rect 224 114 225 115
rect 223 114 224 115
rect 222 114 223 115
rect 221 114 222 115
rect 220 114 221 115
rect 219 114 220 115
rect 218 114 219 115
rect 217 114 218 115
rect 216 114 217 115
rect 215 114 216 115
rect 214 114 215 115
rect 213 114 214 115
rect 212 114 213 115
rect 211 114 212 115
rect 210 114 211 115
rect 209 114 210 115
rect 208 114 209 115
rect 207 114 208 115
rect 206 114 207 115
rect 205 114 206 115
rect 204 114 205 115
rect 203 114 204 115
rect 202 114 203 115
rect 201 114 202 115
rect 200 114 201 115
rect 199 114 200 115
rect 198 114 199 115
rect 197 114 198 115
rect 196 114 197 115
rect 195 114 196 115
rect 194 114 195 115
rect 193 114 194 115
rect 192 114 193 115
rect 191 114 192 115
rect 190 114 191 115
rect 189 114 190 115
rect 188 114 189 115
rect 187 114 188 115
rect 186 114 187 115
rect 185 114 186 115
rect 184 114 185 115
rect 183 114 184 115
rect 182 114 183 115
rect 181 114 182 115
rect 180 114 181 115
rect 179 114 180 115
rect 178 114 179 115
rect 177 114 178 115
rect 176 114 177 115
rect 175 114 176 115
rect 174 114 175 115
rect 156 114 157 115
rect 155 114 156 115
rect 154 114 155 115
rect 153 114 154 115
rect 152 114 153 115
rect 151 114 152 115
rect 150 114 151 115
rect 149 114 150 115
rect 148 114 149 115
rect 147 114 148 115
rect 146 114 147 115
rect 145 114 146 115
rect 144 114 145 115
rect 143 114 144 115
rect 142 114 143 115
rect 141 114 142 115
rect 140 114 141 115
rect 139 114 140 115
rect 138 114 139 115
rect 137 114 138 115
rect 136 114 137 115
rect 135 114 136 115
rect 134 114 135 115
rect 133 114 134 115
rect 132 114 133 115
rect 131 114 132 115
rect 130 114 131 115
rect 129 114 130 115
rect 128 114 129 115
rect 127 114 128 115
rect 126 114 127 115
rect 125 114 126 115
rect 124 114 125 115
rect 123 114 124 115
rect 122 114 123 115
rect 121 114 122 115
rect 120 114 121 115
rect 119 114 120 115
rect 118 114 119 115
rect 117 114 118 115
rect 116 114 117 115
rect 115 114 116 115
rect 114 114 115 115
rect 113 114 114 115
rect 112 114 113 115
rect 111 114 112 115
rect 110 114 111 115
rect 109 114 110 115
rect 108 114 109 115
rect 107 114 108 115
rect 106 114 107 115
rect 105 114 106 115
rect 104 114 105 115
rect 103 114 104 115
rect 102 114 103 115
rect 101 114 102 115
rect 100 114 101 115
rect 99 114 100 115
rect 98 114 99 115
rect 97 114 98 115
rect 96 114 97 115
rect 95 114 96 115
rect 94 114 95 115
rect 93 114 94 115
rect 92 114 93 115
rect 91 114 92 115
rect 90 114 91 115
rect 89 114 90 115
rect 88 114 89 115
rect 87 114 88 115
rect 86 114 87 115
rect 85 114 86 115
rect 84 114 85 115
rect 83 114 84 115
rect 82 114 83 115
rect 81 114 82 115
rect 65 114 66 115
rect 64 114 65 115
rect 63 114 64 115
rect 62 114 63 115
rect 61 114 62 115
rect 60 114 61 115
rect 59 114 60 115
rect 58 114 59 115
rect 57 114 58 115
rect 56 114 57 115
rect 55 114 56 115
rect 54 114 55 115
rect 53 114 54 115
rect 52 114 53 115
rect 51 114 52 115
rect 50 114 51 115
rect 49 114 50 115
rect 48 114 49 115
rect 47 114 48 115
rect 46 114 47 115
rect 45 114 46 115
rect 44 114 45 115
rect 43 114 44 115
rect 42 114 43 115
rect 41 114 42 115
rect 40 114 41 115
rect 39 114 40 115
rect 38 114 39 115
rect 37 114 38 115
rect 482 115 483 116
rect 481 115 482 116
rect 463 115 464 116
rect 462 115 463 116
rect 439 115 440 116
rect 438 115 439 116
rect 437 115 438 116
rect 436 115 437 116
rect 435 115 436 116
rect 434 115 435 116
rect 433 115 434 116
rect 432 115 433 116
rect 431 115 432 116
rect 430 115 431 116
rect 429 115 430 116
rect 428 115 429 116
rect 427 115 428 116
rect 426 115 427 116
rect 425 115 426 116
rect 424 115 425 116
rect 423 115 424 116
rect 422 115 423 116
rect 421 115 422 116
rect 420 115 421 116
rect 419 115 420 116
rect 418 115 419 116
rect 417 115 418 116
rect 416 115 417 116
rect 415 115 416 116
rect 414 115 415 116
rect 413 115 414 116
rect 412 115 413 116
rect 411 115 412 116
rect 410 115 411 116
rect 409 115 410 116
rect 408 115 409 116
rect 407 115 408 116
rect 406 115 407 116
rect 405 115 406 116
rect 404 115 405 116
rect 403 115 404 116
rect 402 115 403 116
rect 401 115 402 116
rect 400 115 401 116
rect 399 115 400 116
rect 398 115 399 116
rect 397 115 398 116
rect 267 115 268 116
rect 266 115 267 116
rect 265 115 266 116
rect 264 115 265 116
rect 263 115 264 116
rect 262 115 263 116
rect 261 115 262 116
rect 260 115 261 116
rect 259 115 260 116
rect 258 115 259 116
rect 257 115 258 116
rect 256 115 257 116
rect 255 115 256 116
rect 254 115 255 116
rect 253 115 254 116
rect 252 115 253 116
rect 251 115 252 116
rect 250 115 251 116
rect 249 115 250 116
rect 248 115 249 116
rect 247 115 248 116
rect 246 115 247 116
rect 245 115 246 116
rect 244 115 245 116
rect 243 115 244 116
rect 242 115 243 116
rect 241 115 242 116
rect 240 115 241 116
rect 239 115 240 116
rect 238 115 239 116
rect 237 115 238 116
rect 236 115 237 116
rect 235 115 236 116
rect 234 115 235 116
rect 233 115 234 116
rect 232 115 233 116
rect 231 115 232 116
rect 230 115 231 116
rect 229 115 230 116
rect 228 115 229 116
rect 227 115 228 116
rect 226 115 227 116
rect 225 115 226 116
rect 224 115 225 116
rect 223 115 224 116
rect 222 115 223 116
rect 221 115 222 116
rect 220 115 221 116
rect 219 115 220 116
rect 218 115 219 116
rect 217 115 218 116
rect 216 115 217 116
rect 215 115 216 116
rect 214 115 215 116
rect 213 115 214 116
rect 212 115 213 116
rect 211 115 212 116
rect 210 115 211 116
rect 209 115 210 116
rect 208 115 209 116
rect 207 115 208 116
rect 206 115 207 116
rect 205 115 206 116
rect 204 115 205 116
rect 203 115 204 116
rect 202 115 203 116
rect 201 115 202 116
rect 200 115 201 116
rect 199 115 200 116
rect 198 115 199 116
rect 197 115 198 116
rect 196 115 197 116
rect 195 115 196 116
rect 194 115 195 116
rect 193 115 194 116
rect 192 115 193 116
rect 191 115 192 116
rect 190 115 191 116
rect 189 115 190 116
rect 188 115 189 116
rect 187 115 188 116
rect 186 115 187 116
rect 185 115 186 116
rect 184 115 185 116
rect 183 115 184 116
rect 182 115 183 116
rect 181 115 182 116
rect 180 115 181 116
rect 179 115 180 116
rect 178 115 179 116
rect 177 115 178 116
rect 176 115 177 116
rect 175 115 176 116
rect 174 115 175 116
rect 156 115 157 116
rect 155 115 156 116
rect 154 115 155 116
rect 153 115 154 116
rect 152 115 153 116
rect 151 115 152 116
rect 150 115 151 116
rect 149 115 150 116
rect 148 115 149 116
rect 147 115 148 116
rect 146 115 147 116
rect 145 115 146 116
rect 144 115 145 116
rect 143 115 144 116
rect 142 115 143 116
rect 141 115 142 116
rect 140 115 141 116
rect 139 115 140 116
rect 138 115 139 116
rect 137 115 138 116
rect 136 115 137 116
rect 135 115 136 116
rect 134 115 135 116
rect 133 115 134 116
rect 132 115 133 116
rect 131 115 132 116
rect 130 115 131 116
rect 129 115 130 116
rect 128 115 129 116
rect 127 115 128 116
rect 126 115 127 116
rect 125 115 126 116
rect 124 115 125 116
rect 123 115 124 116
rect 122 115 123 116
rect 121 115 122 116
rect 120 115 121 116
rect 119 115 120 116
rect 118 115 119 116
rect 117 115 118 116
rect 116 115 117 116
rect 115 115 116 116
rect 114 115 115 116
rect 113 115 114 116
rect 112 115 113 116
rect 111 115 112 116
rect 110 115 111 116
rect 109 115 110 116
rect 108 115 109 116
rect 107 115 108 116
rect 106 115 107 116
rect 105 115 106 116
rect 104 115 105 116
rect 103 115 104 116
rect 102 115 103 116
rect 101 115 102 116
rect 100 115 101 116
rect 99 115 100 116
rect 98 115 99 116
rect 97 115 98 116
rect 96 115 97 116
rect 95 115 96 116
rect 94 115 95 116
rect 93 115 94 116
rect 92 115 93 116
rect 91 115 92 116
rect 90 115 91 116
rect 89 115 90 116
rect 88 115 89 116
rect 87 115 88 116
rect 86 115 87 116
rect 85 115 86 116
rect 84 115 85 116
rect 83 115 84 116
rect 82 115 83 116
rect 81 115 82 116
rect 80 115 81 116
rect 79 115 80 116
rect 65 115 66 116
rect 64 115 65 116
rect 63 115 64 116
rect 62 115 63 116
rect 61 115 62 116
rect 60 115 61 116
rect 59 115 60 116
rect 58 115 59 116
rect 57 115 58 116
rect 56 115 57 116
rect 55 115 56 116
rect 54 115 55 116
rect 53 115 54 116
rect 52 115 53 116
rect 51 115 52 116
rect 50 115 51 116
rect 49 115 50 116
rect 48 115 49 116
rect 47 115 48 116
rect 46 115 47 116
rect 45 115 46 116
rect 44 115 45 116
rect 43 115 44 116
rect 42 115 43 116
rect 41 115 42 116
rect 40 115 41 116
rect 39 115 40 116
rect 38 115 39 116
rect 37 115 38 116
rect 36 115 37 116
rect 482 116 483 117
rect 481 116 482 117
rect 480 116 481 117
rect 479 116 480 117
rect 478 116 479 117
rect 477 116 478 117
rect 476 116 477 117
rect 475 116 476 117
rect 474 116 475 117
rect 473 116 474 117
rect 472 116 473 117
rect 471 116 472 117
rect 470 116 471 117
rect 469 116 470 117
rect 468 116 469 117
rect 467 116 468 117
rect 466 116 467 117
rect 465 116 466 117
rect 464 116 465 117
rect 463 116 464 117
rect 462 116 463 117
rect 440 116 441 117
rect 439 116 440 117
rect 438 116 439 117
rect 437 116 438 117
rect 436 116 437 117
rect 435 116 436 117
rect 434 116 435 117
rect 433 116 434 117
rect 432 116 433 117
rect 431 116 432 117
rect 430 116 431 117
rect 429 116 430 117
rect 428 116 429 117
rect 427 116 428 117
rect 426 116 427 117
rect 425 116 426 117
rect 424 116 425 117
rect 423 116 424 117
rect 422 116 423 117
rect 421 116 422 117
rect 420 116 421 117
rect 419 116 420 117
rect 418 116 419 117
rect 417 116 418 117
rect 416 116 417 117
rect 415 116 416 117
rect 414 116 415 117
rect 413 116 414 117
rect 412 116 413 117
rect 411 116 412 117
rect 410 116 411 117
rect 409 116 410 117
rect 408 116 409 117
rect 407 116 408 117
rect 406 116 407 117
rect 405 116 406 117
rect 404 116 405 117
rect 403 116 404 117
rect 402 116 403 117
rect 401 116 402 117
rect 400 116 401 117
rect 399 116 400 117
rect 398 116 399 117
rect 397 116 398 117
rect 259 116 260 117
rect 258 116 259 117
rect 257 116 258 117
rect 256 116 257 117
rect 255 116 256 117
rect 254 116 255 117
rect 253 116 254 117
rect 252 116 253 117
rect 251 116 252 117
rect 250 116 251 117
rect 249 116 250 117
rect 248 116 249 117
rect 247 116 248 117
rect 246 116 247 117
rect 245 116 246 117
rect 244 116 245 117
rect 243 116 244 117
rect 242 116 243 117
rect 241 116 242 117
rect 240 116 241 117
rect 239 116 240 117
rect 238 116 239 117
rect 237 116 238 117
rect 236 116 237 117
rect 235 116 236 117
rect 234 116 235 117
rect 233 116 234 117
rect 232 116 233 117
rect 231 116 232 117
rect 230 116 231 117
rect 229 116 230 117
rect 228 116 229 117
rect 227 116 228 117
rect 226 116 227 117
rect 225 116 226 117
rect 224 116 225 117
rect 223 116 224 117
rect 222 116 223 117
rect 221 116 222 117
rect 220 116 221 117
rect 219 116 220 117
rect 218 116 219 117
rect 217 116 218 117
rect 216 116 217 117
rect 215 116 216 117
rect 214 116 215 117
rect 213 116 214 117
rect 212 116 213 117
rect 211 116 212 117
rect 210 116 211 117
rect 209 116 210 117
rect 208 116 209 117
rect 207 116 208 117
rect 206 116 207 117
rect 205 116 206 117
rect 204 116 205 117
rect 203 116 204 117
rect 202 116 203 117
rect 201 116 202 117
rect 200 116 201 117
rect 199 116 200 117
rect 198 116 199 117
rect 197 116 198 117
rect 196 116 197 117
rect 195 116 196 117
rect 194 116 195 117
rect 193 116 194 117
rect 192 116 193 117
rect 191 116 192 117
rect 190 116 191 117
rect 189 116 190 117
rect 188 116 189 117
rect 187 116 188 117
rect 186 116 187 117
rect 185 116 186 117
rect 184 116 185 117
rect 183 116 184 117
rect 182 116 183 117
rect 181 116 182 117
rect 180 116 181 117
rect 179 116 180 117
rect 178 116 179 117
rect 177 116 178 117
rect 176 116 177 117
rect 175 116 176 117
rect 174 116 175 117
rect 173 116 174 117
rect 155 116 156 117
rect 154 116 155 117
rect 153 116 154 117
rect 152 116 153 117
rect 151 116 152 117
rect 150 116 151 117
rect 149 116 150 117
rect 148 116 149 117
rect 147 116 148 117
rect 146 116 147 117
rect 145 116 146 117
rect 144 116 145 117
rect 143 116 144 117
rect 142 116 143 117
rect 141 116 142 117
rect 140 116 141 117
rect 139 116 140 117
rect 138 116 139 117
rect 137 116 138 117
rect 136 116 137 117
rect 135 116 136 117
rect 134 116 135 117
rect 133 116 134 117
rect 132 116 133 117
rect 131 116 132 117
rect 130 116 131 117
rect 129 116 130 117
rect 128 116 129 117
rect 127 116 128 117
rect 126 116 127 117
rect 125 116 126 117
rect 124 116 125 117
rect 123 116 124 117
rect 122 116 123 117
rect 121 116 122 117
rect 120 116 121 117
rect 119 116 120 117
rect 118 116 119 117
rect 117 116 118 117
rect 116 116 117 117
rect 115 116 116 117
rect 114 116 115 117
rect 113 116 114 117
rect 112 116 113 117
rect 111 116 112 117
rect 110 116 111 117
rect 109 116 110 117
rect 108 116 109 117
rect 107 116 108 117
rect 106 116 107 117
rect 105 116 106 117
rect 104 116 105 117
rect 103 116 104 117
rect 102 116 103 117
rect 101 116 102 117
rect 100 116 101 117
rect 99 116 100 117
rect 98 116 99 117
rect 97 116 98 117
rect 96 116 97 117
rect 95 116 96 117
rect 94 116 95 117
rect 93 116 94 117
rect 92 116 93 117
rect 91 116 92 117
rect 90 116 91 117
rect 89 116 90 117
rect 88 116 89 117
rect 87 116 88 117
rect 86 116 87 117
rect 85 116 86 117
rect 84 116 85 117
rect 83 116 84 117
rect 82 116 83 117
rect 81 116 82 117
rect 80 116 81 117
rect 79 116 80 117
rect 78 116 79 117
rect 77 116 78 117
rect 64 116 65 117
rect 63 116 64 117
rect 62 116 63 117
rect 61 116 62 117
rect 60 116 61 117
rect 59 116 60 117
rect 58 116 59 117
rect 57 116 58 117
rect 56 116 57 117
rect 55 116 56 117
rect 54 116 55 117
rect 53 116 54 117
rect 52 116 53 117
rect 51 116 52 117
rect 50 116 51 117
rect 49 116 50 117
rect 48 116 49 117
rect 47 116 48 117
rect 46 116 47 117
rect 45 116 46 117
rect 44 116 45 117
rect 43 116 44 117
rect 42 116 43 117
rect 41 116 42 117
rect 40 116 41 117
rect 39 116 40 117
rect 38 116 39 117
rect 37 116 38 117
rect 36 116 37 117
rect 35 116 36 117
rect 482 117 483 118
rect 481 117 482 118
rect 480 117 481 118
rect 479 117 480 118
rect 478 117 479 118
rect 477 117 478 118
rect 476 117 477 118
rect 475 117 476 118
rect 474 117 475 118
rect 473 117 474 118
rect 472 117 473 118
rect 471 117 472 118
rect 470 117 471 118
rect 469 117 470 118
rect 468 117 469 118
rect 467 117 468 118
rect 466 117 467 118
rect 465 117 466 118
rect 464 117 465 118
rect 463 117 464 118
rect 462 117 463 118
rect 440 117 441 118
rect 439 117 440 118
rect 438 117 439 118
rect 437 117 438 118
rect 436 117 437 118
rect 435 117 436 118
rect 434 117 435 118
rect 433 117 434 118
rect 432 117 433 118
rect 431 117 432 118
rect 430 117 431 118
rect 429 117 430 118
rect 428 117 429 118
rect 427 117 428 118
rect 426 117 427 118
rect 425 117 426 118
rect 424 117 425 118
rect 423 117 424 118
rect 422 117 423 118
rect 421 117 422 118
rect 420 117 421 118
rect 419 117 420 118
rect 418 117 419 118
rect 417 117 418 118
rect 416 117 417 118
rect 415 117 416 118
rect 414 117 415 118
rect 413 117 414 118
rect 412 117 413 118
rect 411 117 412 118
rect 410 117 411 118
rect 409 117 410 118
rect 408 117 409 118
rect 407 117 408 118
rect 406 117 407 118
rect 405 117 406 118
rect 404 117 405 118
rect 403 117 404 118
rect 402 117 403 118
rect 401 117 402 118
rect 400 117 401 118
rect 399 117 400 118
rect 398 117 399 118
rect 397 117 398 118
rect 255 117 256 118
rect 254 117 255 118
rect 253 117 254 118
rect 252 117 253 118
rect 251 117 252 118
rect 250 117 251 118
rect 249 117 250 118
rect 248 117 249 118
rect 247 117 248 118
rect 246 117 247 118
rect 245 117 246 118
rect 244 117 245 118
rect 243 117 244 118
rect 242 117 243 118
rect 241 117 242 118
rect 240 117 241 118
rect 239 117 240 118
rect 238 117 239 118
rect 237 117 238 118
rect 236 117 237 118
rect 235 117 236 118
rect 234 117 235 118
rect 233 117 234 118
rect 232 117 233 118
rect 231 117 232 118
rect 230 117 231 118
rect 229 117 230 118
rect 228 117 229 118
rect 227 117 228 118
rect 226 117 227 118
rect 225 117 226 118
rect 224 117 225 118
rect 223 117 224 118
rect 222 117 223 118
rect 221 117 222 118
rect 220 117 221 118
rect 219 117 220 118
rect 218 117 219 118
rect 217 117 218 118
rect 216 117 217 118
rect 215 117 216 118
rect 214 117 215 118
rect 213 117 214 118
rect 212 117 213 118
rect 211 117 212 118
rect 210 117 211 118
rect 209 117 210 118
rect 208 117 209 118
rect 207 117 208 118
rect 206 117 207 118
rect 205 117 206 118
rect 204 117 205 118
rect 203 117 204 118
rect 202 117 203 118
rect 201 117 202 118
rect 200 117 201 118
rect 199 117 200 118
rect 198 117 199 118
rect 197 117 198 118
rect 196 117 197 118
rect 195 117 196 118
rect 194 117 195 118
rect 193 117 194 118
rect 192 117 193 118
rect 191 117 192 118
rect 190 117 191 118
rect 189 117 190 118
rect 188 117 189 118
rect 187 117 188 118
rect 186 117 187 118
rect 185 117 186 118
rect 184 117 185 118
rect 183 117 184 118
rect 182 117 183 118
rect 181 117 182 118
rect 180 117 181 118
rect 179 117 180 118
rect 178 117 179 118
rect 177 117 178 118
rect 176 117 177 118
rect 175 117 176 118
rect 174 117 175 118
rect 173 117 174 118
rect 155 117 156 118
rect 154 117 155 118
rect 153 117 154 118
rect 152 117 153 118
rect 151 117 152 118
rect 150 117 151 118
rect 149 117 150 118
rect 148 117 149 118
rect 147 117 148 118
rect 146 117 147 118
rect 145 117 146 118
rect 144 117 145 118
rect 143 117 144 118
rect 142 117 143 118
rect 141 117 142 118
rect 140 117 141 118
rect 139 117 140 118
rect 138 117 139 118
rect 137 117 138 118
rect 136 117 137 118
rect 135 117 136 118
rect 134 117 135 118
rect 133 117 134 118
rect 132 117 133 118
rect 131 117 132 118
rect 130 117 131 118
rect 129 117 130 118
rect 128 117 129 118
rect 127 117 128 118
rect 126 117 127 118
rect 125 117 126 118
rect 124 117 125 118
rect 123 117 124 118
rect 122 117 123 118
rect 121 117 122 118
rect 120 117 121 118
rect 119 117 120 118
rect 118 117 119 118
rect 117 117 118 118
rect 116 117 117 118
rect 115 117 116 118
rect 114 117 115 118
rect 113 117 114 118
rect 112 117 113 118
rect 111 117 112 118
rect 110 117 111 118
rect 109 117 110 118
rect 108 117 109 118
rect 107 117 108 118
rect 106 117 107 118
rect 105 117 106 118
rect 104 117 105 118
rect 103 117 104 118
rect 102 117 103 118
rect 101 117 102 118
rect 100 117 101 118
rect 99 117 100 118
rect 98 117 99 118
rect 97 117 98 118
rect 96 117 97 118
rect 95 117 96 118
rect 94 117 95 118
rect 93 117 94 118
rect 92 117 93 118
rect 91 117 92 118
rect 90 117 91 118
rect 89 117 90 118
rect 88 117 89 118
rect 87 117 88 118
rect 86 117 87 118
rect 85 117 86 118
rect 84 117 85 118
rect 83 117 84 118
rect 82 117 83 118
rect 81 117 82 118
rect 80 117 81 118
rect 79 117 80 118
rect 78 117 79 118
rect 77 117 78 118
rect 76 117 77 118
rect 64 117 65 118
rect 63 117 64 118
rect 62 117 63 118
rect 61 117 62 118
rect 60 117 61 118
rect 59 117 60 118
rect 58 117 59 118
rect 57 117 58 118
rect 56 117 57 118
rect 55 117 56 118
rect 54 117 55 118
rect 53 117 54 118
rect 52 117 53 118
rect 51 117 52 118
rect 50 117 51 118
rect 49 117 50 118
rect 48 117 49 118
rect 47 117 48 118
rect 46 117 47 118
rect 45 117 46 118
rect 44 117 45 118
rect 43 117 44 118
rect 42 117 43 118
rect 41 117 42 118
rect 40 117 41 118
rect 39 117 40 118
rect 38 117 39 118
rect 37 117 38 118
rect 36 117 37 118
rect 35 117 36 118
rect 34 117 35 118
rect 482 118 483 119
rect 481 118 482 119
rect 480 118 481 119
rect 467 118 468 119
rect 466 118 467 119
rect 465 118 466 119
rect 464 118 465 119
rect 463 118 464 119
rect 462 118 463 119
rect 441 118 442 119
rect 440 118 441 119
rect 439 118 440 119
rect 438 118 439 119
rect 437 118 438 119
rect 436 118 437 119
rect 435 118 436 119
rect 434 118 435 119
rect 433 118 434 119
rect 432 118 433 119
rect 431 118 432 119
rect 430 118 431 119
rect 429 118 430 119
rect 428 118 429 119
rect 427 118 428 119
rect 426 118 427 119
rect 425 118 426 119
rect 424 118 425 119
rect 423 118 424 119
rect 422 118 423 119
rect 421 118 422 119
rect 420 118 421 119
rect 419 118 420 119
rect 418 118 419 119
rect 417 118 418 119
rect 416 118 417 119
rect 415 118 416 119
rect 414 118 415 119
rect 413 118 414 119
rect 412 118 413 119
rect 411 118 412 119
rect 410 118 411 119
rect 409 118 410 119
rect 408 118 409 119
rect 407 118 408 119
rect 406 118 407 119
rect 405 118 406 119
rect 404 118 405 119
rect 403 118 404 119
rect 402 118 403 119
rect 401 118 402 119
rect 400 118 401 119
rect 399 118 400 119
rect 398 118 399 119
rect 397 118 398 119
rect 251 118 252 119
rect 250 118 251 119
rect 249 118 250 119
rect 248 118 249 119
rect 247 118 248 119
rect 246 118 247 119
rect 245 118 246 119
rect 244 118 245 119
rect 243 118 244 119
rect 242 118 243 119
rect 241 118 242 119
rect 240 118 241 119
rect 239 118 240 119
rect 238 118 239 119
rect 237 118 238 119
rect 236 118 237 119
rect 235 118 236 119
rect 234 118 235 119
rect 233 118 234 119
rect 232 118 233 119
rect 231 118 232 119
rect 230 118 231 119
rect 229 118 230 119
rect 228 118 229 119
rect 227 118 228 119
rect 226 118 227 119
rect 225 118 226 119
rect 224 118 225 119
rect 223 118 224 119
rect 222 118 223 119
rect 221 118 222 119
rect 220 118 221 119
rect 219 118 220 119
rect 218 118 219 119
rect 217 118 218 119
rect 216 118 217 119
rect 215 118 216 119
rect 214 118 215 119
rect 213 118 214 119
rect 212 118 213 119
rect 211 118 212 119
rect 210 118 211 119
rect 209 118 210 119
rect 208 118 209 119
rect 207 118 208 119
rect 206 118 207 119
rect 205 118 206 119
rect 204 118 205 119
rect 203 118 204 119
rect 202 118 203 119
rect 201 118 202 119
rect 200 118 201 119
rect 199 118 200 119
rect 198 118 199 119
rect 197 118 198 119
rect 196 118 197 119
rect 195 118 196 119
rect 194 118 195 119
rect 193 118 194 119
rect 192 118 193 119
rect 191 118 192 119
rect 190 118 191 119
rect 189 118 190 119
rect 188 118 189 119
rect 187 118 188 119
rect 186 118 187 119
rect 185 118 186 119
rect 184 118 185 119
rect 183 118 184 119
rect 182 118 183 119
rect 181 118 182 119
rect 180 118 181 119
rect 179 118 180 119
rect 178 118 179 119
rect 177 118 178 119
rect 176 118 177 119
rect 175 118 176 119
rect 174 118 175 119
rect 173 118 174 119
rect 172 118 173 119
rect 155 118 156 119
rect 154 118 155 119
rect 153 118 154 119
rect 152 118 153 119
rect 151 118 152 119
rect 150 118 151 119
rect 149 118 150 119
rect 148 118 149 119
rect 147 118 148 119
rect 146 118 147 119
rect 145 118 146 119
rect 144 118 145 119
rect 143 118 144 119
rect 142 118 143 119
rect 141 118 142 119
rect 140 118 141 119
rect 139 118 140 119
rect 138 118 139 119
rect 137 118 138 119
rect 136 118 137 119
rect 135 118 136 119
rect 134 118 135 119
rect 133 118 134 119
rect 132 118 133 119
rect 131 118 132 119
rect 130 118 131 119
rect 129 118 130 119
rect 128 118 129 119
rect 127 118 128 119
rect 126 118 127 119
rect 125 118 126 119
rect 124 118 125 119
rect 123 118 124 119
rect 122 118 123 119
rect 121 118 122 119
rect 120 118 121 119
rect 119 118 120 119
rect 118 118 119 119
rect 117 118 118 119
rect 116 118 117 119
rect 115 118 116 119
rect 114 118 115 119
rect 113 118 114 119
rect 112 118 113 119
rect 111 118 112 119
rect 110 118 111 119
rect 109 118 110 119
rect 108 118 109 119
rect 107 118 108 119
rect 106 118 107 119
rect 105 118 106 119
rect 104 118 105 119
rect 103 118 104 119
rect 102 118 103 119
rect 101 118 102 119
rect 100 118 101 119
rect 99 118 100 119
rect 98 118 99 119
rect 97 118 98 119
rect 96 118 97 119
rect 95 118 96 119
rect 94 118 95 119
rect 93 118 94 119
rect 92 118 93 119
rect 91 118 92 119
rect 90 118 91 119
rect 89 118 90 119
rect 88 118 89 119
rect 87 118 88 119
rect 86 118 87 119
rect 85 118 86 119
rect 84 118 85 119
rect 83 118 84 119
rect 82 118 83 119
rect 81 118 82 119
rect 80 118 81 119
rect 79 118 80 119
rect 78 118 79 119
rect 77 118 78 119
rect 76 118 77 119
rect 75 118 76 119
rect 64 118 65 119
rect 63 118 64 119
rect 62 118 63 119
rect 61 118 62 119
rect 60 118 61 119
rect 59 118 60 119
rect 58 118 59 119
rect 57 118 58 119
rect 56 118 57 119
rect 55 118 56 119
rect 54 118 55 119
rect 53 118 54 119
rect 52 118 53 119
rect 51 118 52 119
rect 50 118 51 119
rect 49 118 50 119
rect 48 118 49 119
rect 47 118 48 119
rect 46 118 47 119
rect 45 118 46 119
rect 44 118 45 119
rect 43 118 44 119
rect 42 118 43 119
rect 41 118 42 119
rect 40 118 41 119
rect 39 118 40 119
rect 38 118 39 119
rect 37 118 38 119
rect 36 118 37 119
rect 35 118 36 119
rect 34 118 35 119
rect 482 119 483 120
rect 468 119 469 120
rect 467 119 468 120
rect 466 119 467 120
rect 465 119 466 120
rect 464 119 465 120
rect 463 119 464 120
rect 462 119 463 120
rect 441 119 442 120
rect 440 119 441 120
rect 439 119 440 120
rect 438 119 439 120
rect 437 119 438 120
rect 436 119 437 120
rect 435 119 436 120
rect 434 119 435 120
rect 433 119 434 120
rect 432 119 433 120
rect 431 119 432 120
rect 430 119 431 120
rect 429 119 430 120
rect 428 119 429 120
rect 401 119 402 120
rect 400 119 401 120
rect 399 119 400 120
rect 398 119 399 120
rect 397 119 398 120
rect 248 119 249 120
rect 247 119 248 120
rect 246 119 247 120
rect 245 119 246 120
rect 244 119 245 120
rect 243 119 244 120
rect 242 119 243 120
rect 241 119 242 120
rect 240 119 241 120
rect 239 119 240 120
rect 238 119 239 120
rect 237 119 238 120
rect 236 119 237 120
rect 235 119 236 120
rect 234 119 235 120
rect 233 119 234 120
rect 232 119 233 120
rect 231 119 232 120
rect 230 119 231 120
rect 229 119 230 120
rect 228 119 229 120
rect 227 119 228 120
rect 226 119 227 120
rect 225 119 226 120
rect 224 119 225 120
rect 223 119 224 120
rect 222 119 223 120
rect 221 119 222 120
rect 220 119 221 120
rect 219 119 220 120
rect 218 119 219 120
rect 217 119 218 120
rect 216 119 217 120
rect 215 119 216 120
rect 214 119 215 120
rect 213 119 214 120
rect 212 119 213 120
rect 211 119 212 120
rect 210 119 211 120
rect 209 119 210 120
rect 208 119 209 120
rect 207 119 208 120
rect 206 119 207 120
rect 205 119 206 120
rect 204 119 205 120
rect 203 119 204 120
rect 202 119 203 120
rect 201 119 202 120
rect 200 119 201 120
rect 199 119 200 120
rect 198 119 199 120
rect 197 119 198 120
rect 196 119 197 120
rect 195 119 196 120
rect 194 119 195 120
rect 193 119 194 120
rect 192 119 193 120
rect 191 119 192 120
rect 190 119 191 120
rect 189 119 190 120
rect 188 119 189 120
rect 187 119 188 120
rect 186 119 187 120
rect 185 119 186 120
rect 184 119 185 120
rect 183 119 184 120
rect 182 119 183 120
rect 181 119 182 120
rect 180 119 181 120
rect 179 119 180 120
rect 178 119 179 120
rect 177 119 178 120
rect 176 119 177 120
rect 175 119 176 120
rect 174 119 175 120
rect 173 119 174 120
rect 172 119 173 120
rect 154 119 155 120
rect 153 119 154 120
rect 152 119 153 120
rect 151 119 152 120
rect 150 119 151 120
rect 149 119 150 120
rect 148 119 149 120
rect 147 119 148 120
rect 146 119 147 120
rect 145 119 146 120
rect 144 119 145 120
rect 143 119 144 120
rect 142 119 143 120
rect 141 119 142 120
rect 140 119 141 120
rect 139 119 140 120
rect 138 119 139 120
rect 137 119 138 120
rect 136 119 137 120
rect 135 119 136 120
rect 134 119 135 120
rect 133 119 134 120
rect 132 119 133 120
rect 131 119 132 120
rect 130 119 131 120
rect 129 119 130 120
rect 128 119 129 120
rect 127 119 128 120
rect 126 119 127 120
rect 125 119 126 120
rect 124 119 125 120
rect 123 119 124 120
rect 122 119 123 120
rect 121 119 122 120
rect 120 119 121 120
rect 119 119 120 120
rect 118 119 119 120
rect 117 119 118 120
rect 116 119 117 120
rect 115 119 116 120
rect 114 119 115 120
rect 113 119 114 120
rect 112 119 113 120
rect 111 119 112 120
rect 110 119 111 120
rect 109 119 110 120
rect 108 119 109 120
rect 107 119 108 120
rect 106 119 107 120
rect 105 119 106 120
rect 104 119 105 120
rect 103 119 104 120
rect 102 119 103 120
rect 101 119 102 120
rect 100 119 101 120
rect 99 119 100 120
rect 98 119 99 120
rect 97 119 98 120
rect 96 119 97 120
rect 95 119 96 120
rect 94 119 95 120
rect 93 119 94 120
rect 92 119 93 120
rect 91 119 92 120
rect 90 119 91 120
rect 89 119 90 120
rect 88 119 89 120
rect 87 119 88 120
rect 86 119 87 120
rect 85 119 86 120
rect 84 119 85 120
rect 83 119 84 120
rect 82 119 83 120
rect 81 119 82 120
rect 80 119 81 120
rect 79 119 80 120
rect 78 119 79 120
rect 77 119 78 120
rect 76 119 77 120
rect 75 119 76 120
rect 74 119 75 120
rect 73 119 74 120
rect 64 119 65 120
rect 63 119 64 120
rect 62 119 63 120
rect 61 119 62 120
rect 60 119 61 120
rect 59 119 60 120
rect 58 119 59 120
rect 57 119 58 120
rect 56 119 57 120
rect 55 119 56 120
rect 54 119 55 120
rect 53 119 54 120
rect 52 119 53 120
rect 51 119 52 120
rect 50 119 51 120
rect 49 119 50 120
rect 48 119 49 120
rect 47 119 48 120
rect 46 119 47 120
rect 45 119 46 120
rect 44 119 45 120
rect 43 119 44 120
rect 42 119 43 120
rect 41 119 42 120
rect 40 119 41 120
rect 39 119 40 120
rect 38 119 39 120
rect 37 119 38 120
rect 36 119 37 120
rect 35 119 36 120
rect 34 119 35 120
rect 33 119 34 120
rect 482 120 483 121
rect 469 120 470 121
rect 468 120 469 121
rect 467 120 468 121
rect 466 120 467 121
rect 465 120 466 121
rect 464 120 465 121
rect 463 120 464 121
rect 441 120 442 121
rect 440 120 441 121
rect 439 120 440 121
rect 438 120 439 121
rect 437 120 438 121
rect 436 120 437 121
rect 435 120 436 121
rect 434 120 435 121
rect 433 120 434 121
rect 432 120 433 121
rect 400 120 401 121
rect 399 120 400 121
rect 398 120 399 121
rect 397 120 398 121
rect 246 120 247 121
rect 245 120 246 121
rect 244 120 245 121
rect 243 120 244 121
rect 242 120 243 121
rect 241 120 242 121
rect 240 120 241 121
rect 239 120 240 121
rect 238 120 239 121
rect 237 120 238 121
rect 236 120 237 121
rect 235 120 236 121
rect 234 120 235 121
rect 233 120 234 121
rect 232 120 233 121
rect 231 120 232 121
rect 230 120 231 121
rect 229 120 230 121
rect 228 120 229 121
rect 227 120 228 121
rect 226 120 227 121
rect 225 120 226 121
rect 224 120 225 121
rect 223 120 224 121
rect 222 120 223 121
rect 221 120 222 121
rect 220 120 221 121
rect 219 120 220 121
rect 218 120 219 121
rect 217 120 218 121
rect 216 120 217 121
rect 215 120 216 121
rect 214 120 215 121
rect 213 120 214 121
rect 212 120 213 121
rect 211 120 212 121
rect 210 120 211 121
rect 209 120 210 121
rect 208 120 209 121
rect 207 120 208 121
rect 206 120 207 121
rect 205 120 206 121
rect 204 120 205 121
rect 203 120 204 121
rect 202 120 203 121
rect 201 120 202 121
rect 200 120 201 121
rect 199 120 200 121
rect 198 120 199 121
rect 197 120 198 121
rect 196 120 197 121
rect 195 120 196 121
rect 194 120 195 121
rect 193 120 194 121
rect 192 120 193 121
rect 191 120 192 121
rect 190 120 191 121
rect 189 120 190 121
rect 188 120 189 121
rect 187 120 188 121
rect 186 120 187 121
rect 185 120 186 121
rect 184 120 185 121
rect 183 120 184 121
rect 182 120 183 121
rect 181 120 182 121
rect 180 120 181 121
rect 179 120 180 121
rect 178 120 179 121
rect 177 120 178 121
rect 176 120 177 121
rect 175 120 176 121
rect 174 120 175 121
rect 173 120 174 121
rect 172 120 173 121
rect 154 120 155 121
rect 153 120 154 121
rect 152 120 153 121
rect 151 120 152 121
rect 150 120 151 121
rect 149 120 150 121
rect 148 120 149 121
rect 147 120 148 121
rect 146 120 147 121
rect 145 120 146 121
rect 144 120 145 121
rect 143 120 144 121
rect 142 120 143 121
rect 141 120 142 121
rect 140 120 141 121
rect 139 120 140 121
rect 138 120 139 121
rect 137 120 138 121
rect 136 120 137 121
rect 135 120 136 121
rect 134 120 135 121
rect 133 120 134 121
rect 132 120 133 121
rect 131 120 132 121
rect 130 120 131 121
rect 129 120 130 121
rect 128 120 129 121
rect 127 120 128 121
rect 126 120 127 121
rect 125 120 126 121
rect 124 120 125 121
rect 123 120 124 121
rect 122 120 123 121
rect 121 120 122 121
rect 120 120 121 121
rect 119 120 120 121
rect 118 120 119 121
rect 117 120 118 121
rect 116 120 117 121
rect 115 120 116 121
rect 114 120 115 121
rect 113 120 114 121
rect 112 120 113 121
rect 111 120 112 121
rect 110 120 111 121
rect 109 120 110 121
rect 108 120 109 121
rect 107 120 108 121
rect 106 120 107 121
rect 105 120 106 121
rect 104 120 105 121
rect 103 120 104 121
rect 102 120 103 121
rect 101 120 102 121
rect 100 120 101 121
rect 99 120 100 121
rect 98 120 99 121
rect 97 120 98 121
rect 96 120 97 121
rect 95 120 96 121
rect 94 120 95 121
rect 93 120 94 121
rect 92 120 93 121
rect 91 120 92 121
rect 90 120 91 121
rect 89 120 90 121
rect 88 120 89 121
rect 87 120 88 121
rect 86 120 87 121
rect 85 120 86 121
rect 84 120 85 121
rect 83 120 84 121
rect 82 120 83 121
rect 81 120 82 121
rect 80 120 81 121
rect 79 120 80 121
rect 78 120 79 121
rect 77 120 78 121
rect 76 120 77 121
rect 75 120 76 121
rect 74 120 75 121
rect 73 120 74 121
rect 72 120 73 121
rect 63 120 64 121
rect 62 120 63 121
rect 61 120 62 121
rect 60 120 61 121
rect 59 120 60 121
rect 58 120 59 121
rect 57 120 58 121
rect 56 120 57 121
rect 55 120 56 121
rect 54 120 55 121
rect 53 120 54 121
rect 52 120 53 121
rect 51 120 52 121
rect 50 120 51 121
rect 49 120 50 121
rect 48 120 49 121
rect 47 120 48 121
rect 46 120 47 121
rect 45 120 46 121
rect 44 120 45 121
rect 43 120 44 121
rect 42 120 43 121
rect 41 120 42 121
rect 40 120 41 121
rect 39 120 40 121
rect 38 120 39 121
rect 37 120 38 121
rect 36 120 37 121
rect 35 120 36 121
rect 34 120 35 121
rect 33 120 34 121
rect 482 121 483 122
rect 470 121 471 122
rect 469 121 470 122
rect 468 121 469 122
rect 467 121 468 122
rect 466 121 467 122
rect 465 121 466 122
rect 464 121 465 122
rect 442 121 443 122
rect 441 121 442 122
rect 440 121 441 122
rect 439 121 440 122
rect 438 121 439 122
rect 437 121 438 122
rect 436 121 437 122
rect 435 121 436 122
rect 434 121 435 122
rect 399 121 400 122
rect 398 121 399 122
rect 397 121 398 122
rect 244 121 245 122
rect 243 121 244 122
rect 242 121 243 122
rect 241 121 242 122
rect 240 121 241 122
rect 239 121 240 122
rect 238 121 239 122
rect 237 121 238 122
rect 236 121 237 122
rect 235 121 236 122
rect 234 121 235 122
rect 233 121 234 122
rect 232 121 233 122
rect 231 121 232 122
rect 230 121 231 122
rect 229 121 230 122
rect 228 121 229 122
rect 227 121 228 122
rect 226 121 227 122
rect 225 121 226 122
rect 224 121 225 122
rect 223 121 224 122
rect 222 121 223 122
rect 221 121 222 122
rect 220 121 221 122
rect 219 121 220 122
rect 218 121 219 122
rect 217 121 218 122
rect 216 121 217 122
rect 215 121 216 122
rect 214 121 215 122
rect 213 121 214 122
rect 212 121 213 122
rect 211 121 212 122
rect 210 121 211 122
rect 209 121 210 122
rect 208 121 209 122
rect 207 121 208 122
rect 206 121 207 122
rect 205 121 206 122
rect 204 121 205 122
rect 203 121 204 122
rect 202 121 203 122
rect 201 121 202 122
rect 200 121 201 122
rect 199 121 200 122
rect 198 121 199 122
rect 197 121 198 122
rect 196 121 197 122
rect 195 121 196 122
rect 194 121 195 122
rect 193 121 194 122
rect 192 121 193 122
rect 191 121 192 122
rect 190 121 191 122
rect 189 121 190 122
rect 188 121 189 122
rect 187 121 188 122
rect 186 121 187 122
rect 185 121 186 122
rect 184 121 185 122
rect 183 121 184 122
rect 182 121 183 122
rect 181 121 182 122
rect 180 121 181 122
rect 179 121 180 122
rect 178 121 179 122
rect 177 121 178 122
rect 176 121 177 122
rect 175 121 176 122
rect 174 121 175 122
rect 173 121 174 122
rect 172 121 173 122
rect 171 121 172 122
rect 154 121 155 122
rect 153 121 154 122
rect 152 121 153 122
rect 151 121 152 122
rect 150 121 151 122
rect 149 121 150 122
rect 148 121 149 122
rect 147 121 148 122
rect 146 121 147 122
rect 145 121 146 122
rect 144 121 145 122
rect 143 121 144 122
rect 142 121 143 122
rect 141 121 142 122
rect 140 121 141 122
rect 139 121 140 122
rect 138 121 139 122
rect 137 121 138 122
rect 136 121 137 122
rect 135 121 136 122
rect 134 121 135 122
rect 133 121 134 122
rect 132 121 133 122
rect 131 121 132 122
rect 130 121 131 122
rect 129 121 130 122
rect 128 121 129 122
rect 127 121 128 122
rect 126 121 127 122
rect 125 121 126 122
rect 124 121 125 122
rect 123 121 124 122
rect 122 121 123 122
rect 121 121 122 122
rect 120 121 121 122
rect 119 121 120 122
rect 118 121 119 122
rect 117 121 118 122
rect 116 121 117 122
rect 115 121 116 122
rect 114 121 115 122
rect 113 121 114 122
rect 112 121 113 122
rect 111 121 112 122
rect 110 121 111 122
rect 109 121 110 122
rect 108 121 109 122
rect 107 121 108 122
rect 106 121 107 122
rect 105 121 106 122
rect 104 121 105 122
rect 103 121 104 122
rect 102 121 103 122
rect 101 121 102 122
rect 100 121 101 122
rect 99 121 100 122
rect 98 121 99 122
rect 97 121 98 122
rect 96 121 97 122
rect 95 121 96 122
rect 94 121 95 122
rect 93 121 94 122
rect 92 121 93 122
rect 91 121 92 122
rect 90 121 91 122
rect 89 121 90 122
rect 88 121 89 122
rect 87 121 88 122
rect 86 121 87 122
rect 85 121 86 122
rect 84 121 85 122
rect 83 121 84 122
rect 82 121 83 122
rect 81 121 82 122
rect 80 121 81 122
rect 79 121 80 122
rect 78 121 79 122
rect 77 121 78 122
rect 76 121 77 122
rect 75 121 76 122
rect 74 121 75 122
rect 73 121 74 122
rect 72 121 73 122
rect 71 121 72 122
rect 63 121 64 122
rect 62 121 63 122
rect 61 121 62 122
rect 60 121 61 122
rect 59 121 60 122
rect 58 121 59 122
rect 57 121 58 122
rect 56 121 57 122
rect 55 121 56 122
rect 54 121 55 122
rect 53 121 54 122
rect 52 121 53 122
rect 51 121 52 122
rect 50 121 51 122
rect 49 121 50 122
rect 48 121 49 122
rect 47 121 48 122
rect 46 121 47 122
rect 45 121 46 122
rect 44 121 45 122
rect 43 121 44 122
rect 42 121 43 122
rect 41 121 42 122
rect 40 121 41 122
rect 39 121 40 122
rect 38 121 39 122
rect 37 121 38 122
rect 36 121 37 122
rect 35 121 36 122
rect 34 121 35 122
rect 33 121 34 122
rect 32 121 33 122
rect 471 122 472 123
rect 470 122 471 123
rect 469 122 470 123
rect 468 122 469 123
rect 467 122 468 123
rect 466 122 467 123
rect 465 122 466 123
rect 442 122 443 123
rect 441 122 442 123
rect 440 122 441 123
rect 439 122 440 123
rect 438 122 439 123
rect 437 122 438 123
rect 436 122 437 123
rect 435 122 436 123
rect 399 122 400 123
rect 398 122 399 123
rect 397 122 398 123
rect 242 122 243 123
rect 241 122 242 123
rect 240 122 241 123
rect 239 122 240 123
rect 238 122 239 123
rect 237 122 238 123
rect 236 122 237 123
rect 235 122 236 123
rect 234 122 235 123
rect 233 122 234 123
rect 232 122 233 123
rect 231 122 232 123
rect 230 122 231 123
rect 229 122 230 123
rect 228 122 229 123
rect 227 122 228 123
rect 226 122 227 123
rect 225 122 226 123
rect 224 122 225 123
rect 223 122 224 123
rect 222 122 223 123
rect 221 122 222 123
rect 220 122 221 123
rect 219 122 220 123
rect 218 122 219 123
rect 217 122 218 123
rect 216 122 217 123
rect 215 122 216 123
rect 214 122 215 123
rect 213 122 214 123
rect 212 122 213 123
rect 211 122 212 123
rect 210 122 211 123
rect 209 122 210 123
rect 208 122 209 123
rect 207 122 208 123
rect 206 122 207 123
rect 205 122 206 123
rect 204 122 205 123
rect 203 122 204 123
rect 202 122 203 123
rect 201 122 202 123
rect 200 122 201 123
rect 199 122 200 123
rect 198 122 199 123
rect 197 122 198 123
rect 196 122 197 123
rect 195 122 196 123
rect 194 122 195 123
rect 193 122 194 123
rect 192 122 193 123
rect 191 122 192 123
rect 190 122 191 123
rect 189 122 190 123
rect 188 122 189 123
rect 187 122 188 123
rect 186 122 187 123
rect 185 122 186 123
rect 184 122 185 123
rect 183 122 184 123
rect 182 122 183 123
rect 181 122 182 123
rect 180 122 181 123
rect 179 122 180 123
rect 178 122 179 123
rect 177 122 178 123
rect 176 122 177 123
rect 175 122 176 123
rect 174 122 175 123
rect 173 122 174 123
rect 172 122 173 123
rect 171 122 172 123
rect 153 122 154 123
rect 152 122 153 123
rect 151 122 152 123
rect 150 122 151 123
rect 149 122 150 123
rect 148 122 149 123
rect 147 122 148 123
rect 146 122 147 123
rect 145 122 146 123
rect 144 122 145 123
rect 143 122 144 123
rect 142 122 143 123
rect 141 122 142 123
rect 140 122 141 123
rect 139 122 140 123
rect 138 122 139 123
rect 137 122 138 123
rect 136 122 137 123
rect 135 122 136 123
rect 134 122 135 123
rect 133 122 134 123
rect 132 122 133 123
rect 131 122 132 123
rect 130 122 131 123
rect 129 122 130 123
rect 128 122 129 123
rect 127 122 128 123
rect 126 122 127 123
rect 125 122 126 123
rect 124 122 125 123
rect 123 122 124 123
rect 122 122 123 123
rect 121 122 122 123
rect 120 122 121 123
rect 119 122 120 123
rect 118 122 119 123
rect 117 122 118 123
rect 116 122 117 123
rect 115 122 116 123
rect 114 122 115 123
rect 113 122 114 123
rect 112 122 113 123
rect 111 122 112 123
rect 110 122 111 123
rect 109 122 110 123
rect 108 122 109 123
rect 107 122 108 123
rect 106 122 107 123
rect 105 122 106 123
rect 104 122 105 123
rect 103 122 104 123
rect 102 122 103 123
rect 101 122 102 123
rect 100 122 101 123
rect 99 122 100 123
rect 98 122 99 123
rect 97 122 98 123
rect 96 122 97 123
rect 95 122 96 123
rect 94 122 95 123
rect 93 122 94 123
rect 92 122 93 123
rect 91 122 92 123
rect 90 122 91 123
rect 89 122 90 123
rect 88 122 89 123
rect 87 122 88 123
rect 86 122 87 123
rect 85 122 86 123
rect 84 122 85 123
rect 83 122 84 123
rect 82 122 83 123
rect 81 122 82 123
rect 80 122 81 123
rect 79 122 80 123
rect 78 122 79 123
rect 77 122 78 123
rect 76 122 77 123
rect 75 122 76 123
rect 74 122 75 123
rect 73 122 74 123
rect 72 122 73 123
rect 71 122 72 123
rect 63 122 64 123
rect 62 122 63 123
rect 61 122 62 123
rect 60 122 61 123
rect 59 122 60 123
rect 58 122 59 123
rect 57 122 58 123
rect 56 122 57 123
rect 55 122 56 123
rect 54 122 55 123
rect 53 122 54 123
rect 52 122 53 123
rect 51 122 52 123
rect 50 122 51 123
rect 49 122 50 123
rect 48 122 49 123
rect 47 122 48 123
rect 46 122 47 123
rect 45 122 46 123
rect 44 122 45 123
rect 43 122 44 123
rect 42 122 43 123
rect 41 122 42 123
rect 40 122 41 123
rect 39 122 40 123
rect 38 122 39 123
rect 37 122 38 123
rect 36 122 37 123
rect 35 122 36 123
rect 34 122 35 123
rect 33 122 34 123
rect 32 122 33 123
rect 473 123 474 124
rect 472 123 473 124
rect 471 123 472 124
rect 470 123 471 124
rect 469 123 470 124
rect 468 123 469 124
rect 467 123 468 124
rect 466 123 467 124
rect 442 123 443 124
rect 441 123 442 124
rect 440 123 441 124
rect 439 123 440 124
rect 438 123 439 124
rect 437 123 438 124
rect 436 123 437 124
rect 399 123 400 124
rect 398 123 399 124
rect 397 123 398 124
rect 240 123 241 124
rect 239 123 240 124
rect 238 123 239 124
rect 237 123 238 124
rect 236 123 237 124
rect 235 123 236 124
rect 234 123 235 124
rect 233 123 234 124
rect 232 123 233 124
rect 231 123 232 124
rect 230 123 231 124
rect 229 123 230 124
rect 228 123 229 124
rect 227 123 228 124
rect 226 123 227 124
rect 225 123 226 124
rect 224 123 225 124
rect 223 123 224 124
rect 222 123 223 124
rect 221 123 222 124
rect 220 123 221 124
rect 219 123 220 124
rect 218 123 219 124
rect 217 123 218 124
rect 216 123 217 124
rect 215 123 216 124
rect 214 123 215 124
rect 213 123 214 124
rect 212 123 213 124
rect 211 123 212 124
rect 210 123 211 124
rect 209 123 210 124
rect 208 123 209 124
rect 207 123 208 124
rect 206 123 207 124
rect 205 123 206 124
rect 204 123 205 124
rect 203 123 204 124
rect 202 123 203 124
rect 201 123 202 124
rect 200 123 201 124
rect 199 123 200 124
rect 198 123 199 124
rect 197 123 198 124
rect 196 123 197 124
rect 195 123 196 124
rect 194 123 195 124
rect 193 123 194 124
rect 192 123 193 124
rect 191 123 192 124
rect 190 123 191 124
rect 189 123 190 124
rect 188 123 189 124
rect 187 123 188 124
rect 186 123 187 124
rect 185 123 186 124
rect 184 123 185 124
rect 183 123 184 124
rect 182 123 183 124
rect 181 123 182 124
rect 180 123 181 124
rect 179 123 180 124
rect 178 123 179 124
rect 177 123 178 124
rect 176 123 177 124
rect 175 123 176 124
rect 174 123 175 124
rect 173 123 174 124
rect 172 123 173 124
rect 171 123 172 124
rect 170 123 171 124
rect 153 123 154 124
rect 152 123 153 124
rect 151 123 152 124
rect 150 123 151 124
rect 149 123 150 124
rect 148 123 149 124
rect 147 123 148 124
rect 146 123 147 124
rect 145 123 146 124
rect 144 123 145 124
rect 143 123 144 124
rect 142 123 143 124
rect 141 123 142 124
rect 140 123 141 124
rect 139 123 140 124
rect 138 123 139 124
rect 137 123 138 124
rect 136 123 137 124
rect 135 123 136 124
rect 134 123 135 124
rect 133 123 134 124
rect 132 123 133 124
rect 131 123 132 124
rect 130 123 131 124
rect 129 123 130 124
rect 128 123 129 124
rect 127 123 128 124
rect 126 123 127 124
rect 125 123 126 124
rect 124 123 125 124
rect 123 123 124 124
rect 122 123 123 124
rect 121 123 122 124
rect 120 123 121 124
rect 119 123 120 124
rect 118 123 119 124
rect 117 123 118 124
rect 116 123 117 124
rect 115 123 116 124
rect 114 123 115 124
rect 113 123 114 124
rect 112 123 113 124
rect 111 123 112 124
rect 110 123 111 124
rect 109 123 110 124
rect 108 123 109 124
rect 107 123 108 124
rect 106 123 107 124
rect 105 123 106 124
rect 104 123 105 124
rect 103 123 104 124
rect 102 123 103 124
rect 101 123 102 124
rect 100 123 101 124
rect 99 123 100 124
rect 98 123 99 124
rect 97 123 98 124
rect 96 123 97 124
rect 95 123 96 124
rect 94 123 95 124
rect 93 123 94 124
rect 92 123 93 124
rect 91 123 92 124
rect 90 123 91 124
rect 89 123 90 124
rect 88 123 89 124
rect 87 123 88 124
rect 86 123 87 124
rect 85 123 86 124
rect 84 123 85 124
rect 83 123 84 124
rect 82 123 83 124
rect 81 123 82 124
rect 80 123 81 124
rect 79 123 80 124
rect 78 123 79 124
rect 77 123 78 124
rect 76 123 77 124
rect 75 123 76 124
rect 74 123 75 124
rect 73 123 74 124
rect 72 123 73 124
rect 71 123 72 124
rect 70 123 71 124
rect 62 123 63 124
rect 61 123 62 124
rect 60 123 61 124
rect 59 123 60 124
rect 58 123 59 124
rect 57 123 58 124
rect 56 123 57 124
rect 55 123 56 124
rect 54 123 55 124
rect 53 123 54 124
rect 52 123 53 124
rect 51 123 52 124
rect 50 123 51 124
rect 49 123 50 124
rect 48 123 49 124
rect 47 123 48 124
rect 46 123 47 124
rect 45 123 46 124
rect 44 123 45 124
rect 43 123 44 124
rect 42 123 43 124
rect 41 123 42 124
rect 40 123 41 124
rect 39 123 40 124
rect 38 123 39 124
rect 37 123 38 124
rect 36 123 37 124
rect 35 123 36 124
rect 34 123 35 124
rect 33 123 34 124
rect 32 123 33 124
rect 474 124 475 125
rect 473 124 474 125
rect 472 124 473 125
rect 471 124 472 125
rect 470 124 471 125
rect 469 124 470 125
rect 468 124 469 125
rect 442 124 443 125
rect 441 124 442 125
rect 440 124 441 125
rect 439 124 440 125
rect 438 124 439 125
rect 437 124 438 125
rect 398 124 399 125
rect 397 124 398 125
rect 239 124 240 125
rect 238 124 239 125
rect 237 124 238 125
rect 236 124 237 125
rect 235 124 236 125
rect 234 124 235 125
rect 233 124 234 125
rect 232 124 233 125
rect 231 124 232 125
rect 230 124 231 125
rect 229 124 230 125
rect 228 124 229 125
rect 227 124 228 125
rect 226 124 227 125
rect 225 124 226 125
rect 224 124 225 125
rect 223 124 224 125
rect 222 124 223 125
rect 221 124 222 125
rect 220 124 221 125
rect 219 124 220 125
rect 218 124 219 125
rect 217 124 218 125
rect 216 124 217 125
rect 215 124 216 125
rect 214 124 215 125
rect 213 124 214 125
rect 212 124 213 125
rect 211 124 212 125
rect 210 124 211 125
rect 209 124 210 125
rect 208 124 209 125
rect 207 124 208 125
rect 206 124 207 125
rect 205 124 206 125
rect 204 124 205 125
rect 203 124 204 125
rect 202 124 203 125
rect 201 124 202 125
rect 200 124 201 125
rect 199 124 200 125
rect 198 124 199 125
rect 197 124 198 125
rect 196 124 197 125
rect 195 124 196 125
rect 194 124 195 125
rect 193 124 194 125
rect 192 124 193 125
rect 191 124 192 125
rect 190 124 191 125
rect 189 124 190 125
rect 188 124 189 125
rect 187 124 188 125
rect 186 124 187 125
rect 185 124 186 125
rect 184 124 185 125
rect 183 124 184 125
rect 182 124 183 125
rect 181 124 182 125
rect 180 124 181 125
rect 179 124 180 125
rect 178 124 179 125
rect 177 124 178 125
rect 176 124 177 125
rect 175 124 176 125
rect 174 124 175 125
rect 173 124 174 125
rect 172 124 173 125
rect 171 124 172 125
rect 170 124 171 125
rect 153 124 154 125
rect 152 124 153 125
rect 151 124 152 125
rect 150 124 151 125
rect 149 124 150 125
rect 148 124 149 125
rect 147 124 148 125
rect 146 124 147 125
rect 145 124 146 125
rect 144 124 145 125
rect 143 124 144 125
rect 142 124 143 125
rect 141 124 142 125
rect 140 124 141 125
rect 139 124 140 125
rect 138 124 139 125
rect 137 124 138 125
rect 136 124 137 125
rect 135 124 136 125
rect 134 124 135 125
rect 133 124 134 125
rect 132 124 133 125
rect 131 124 132 125
rect 130 124 131 125
rect 129 124 130 125
rect 128 124 129 125
rect 127 124 128 125
rect 126 124 127 125
rect 125 124 126 125
rect 124 124 125 125
rect 123 124 124 125
rect 122 124 123 125
rect 121 124 122 125
rect 120 124 121 125
rect 119 124 120 125
rect 118 124 119 125
rect 117 124 118 125
rect 116 124 117 125
rect 115 124 116 125
rect 114 124 115 125
rect 113 124 114 125
rect 112 124 113 125
rect 111 124 112 125
rect 110 124 111 125
rect 109 124 110 125
rect 108 124 109 125
rect 107 124 108 125
rect 106 124 107 125
rect 105 124 106 125
rect 104 124 105 125
rect 103 124 104 125
rect 102 124 103 125
rect 101 124 102 125
rect 100 124 101 125
rect 99 124 100 125
rect 98 124 99 125
rect 97 124 98 125
rect 96 124 97 125
rect 95 124 96 125
rect 94 124 95 125
rect 93 124 94 125
rect 92 124 93 125
rect 91 124 92 125
rect 90 124 91 125
rect 89 124 90 125
rect 88 124 89 125
rect 87 124 88 125
rect 86 124 87 125
rect 85 124 86 125
rect 84 124 85 125
rect 83 124 84 125
rect 82 124 83 125
rect 81 124 82 125
rect 80 124 81 125
rect 79 124 80 125
rect 78 124 79 125
rect 77 124 78 125
rect 76 124 77 125
rect 75 124 76 125
rect 74 124 75 125
rect 73 124 74 125
rect 72 124 73 125
rect 71 124 72 125
rect 70 124 71 125
rect 69 124 70 125
rect 62 124 63 125
rect 61 124 62 125
rect 60 124 61 125
rect 59 124 60 125
rect 58 124 59 125
rect 57 124 58 125
rect 56 124 57 125
rect 55 124 56 125
rect 54 124 55 125
rect 53 124 54 125
rect 52 124 53 125
rect 51 124 52 125
rect 50 124 51 125
rect 49 124 50 125
rect 48 124 49 125
rect 47 124 48 125
rect 46 124 47 125
rect 45 124 46 125
rect 44 124 45 125
rect 43 124 44 125
rect 42 124 43 125
rect 41 124 42 125
rect 40 124 41 125
rect 39 124 40 125
rect 38 124 39 125
rect 37 124 38 125
rect 36 124 37 125
rect 35 124 36 125
rect 34 124 35 125
rect 33 124 34 125
rect 32 124 33 125
rect 31 124 32 125
rect 475 125 476 126
rect 474 125 475 126
rect 473 125 474 126
rect 472 125 473 126
rect 471 125 472 126
rect 470 125 471 126
rect 469 125 470 126
rect 442 125 443 126
rect 441 125 442 126
rect 440 125 441 126
rect 439 125 440 126
rect 438 125 439 126
rect 437 125 438 126
rect 292 125 293 126
rect 291 125 292 126
rect 290 125 291 126
rect 289 125 290 126
rect 288 125 289 126
rect 287 125 288 126
rect 286 125 287 126
rect 285 125 286 126
rect 284 125 285 126
rect 283 125 284 126
rect 237 125 238 126
rect 236 125 237 126
rect 235 125 236 126
rect 234 125 235 126
rect 233 125 234 126
rect 232 125 233 126
rect 231 125 232 126
rect 230 125 231 126
rect 229 125 230 126
rect 228 125 229 126
rect 227 125 228 126
rect 226 125 227 126
rect 225 125 226 126
rect 224 125 225 126
rect 223 125 224 126
rect 222 125 223 126
rect 221 125 222 126
rect 220 125 221 126
rect 219 125 220 126
rect 218 125 219 126
rect 217 125 218 126
rect 216 125 217 126
rect 215 125 216 126
rect 214 125 215 126
rect 213 125 214 126
rect 212 125 213 126
rect 211 125 212 126
rect 210 125 211 126
rect 209 125 210 126
rect 208 125 209 126
rect 207 125 208 126
rect 206 125 207 126
rect 205 125 206 126
rect 204 125 205 126
rect 203 125 204 126
rect 202 125 203 126
rect 201 125 202 126
rect 200 125 201 126
rect 199 125 200 126
rect 198 125 199 126
rect 197 125 198 126
rect 196 125 197 126
rect 195 125 196 126
rect 194 125 195 126
rect 193 125 194 126
rect 192 125 193 126
rect 191 125 192 126
rect 190 125 191 126
rect 189 125 190 126
rect 188 125 189 126
rect 187 125 188 126
rect 186 125 187 126
rect 185 125 186 126
rect 184 125 185 126
rect 183 125 184 126
rect 182 125 183 126
rect 181 125 182 126
rect 180 125 181 126
rect 179 125 180 126
rect 178 125 179 126
rect 177 125 178 126
rect 176 125 177 126
rect 175 125 176 126
rect 174 125 175 126
rect 173 125 174 126
rect 172 125 173 126
rect 171 125 172 126
rect 170 125 171 126
rect 169 125 170 126
rect 152 125 153 126
rect 151 125 152 126
rect 150 125 151 126
rect 149 125 150 126
rect 148 125 149 126
rect 147 125 148 126
rect 146 125 147 126
rect 145 125 146 126
rect 144 125 145 126
rect 143 125 144 126
rect 142 125 143 126
rect 141 125 142 126
rect 140 125 141 126
rect 139 125 140 126
rect 138 125 139 126
rect 137 125 138 126
rect 136 125 137 126
rect 135 125 136 126
rect 134 125 135 126
rect 133 125 134 126
rect 132 125 133 126
rect 131 125 132 126
rect 130 125 131 126
rect 129 125 130 126
rect 128 125 129 126
rect 127 125 128 126
rect 126 125 127 126
rect 125 125 126 126
rect 124 125 125 126
rect 123 125 124 126
rect 122 125 123 126
rect 121 125 122 126
rect 120 125 121 126
rect 119 125 120 126
rect 118 125 119 126
rect 117 125 118 126
rect 116 125 117 126
rect 115 125 116 126
rect 114 125 115 126
rect 113 125 114 126
rect 112 125 113 126
rect 111 125 112 126
rect 110 125 111 126
rect 109 125 110 126
rect 108 125 109 126
rect 107 125 108 126
rect 106 125 107 126
rect 105 125 106 126
rect 104 125 105 126
rect 103 125 104 126
rect 102 125 103 126
rect 101 125 102 126
rect 100 125 101 126
rect 99 125 100 126
rect 98 125 99 126
rect 97 125 98 126
rect 96 125 97 126
rect 95 125 96 126
rect 94 125 95 126
rect 93 125 94 126
rect 92 125 93 126
rect 91 125 92 126
rect 90 125 91 126
rect 89 125 90 126
rect 88 125 89 126
rect 87 125 88 126
rect 86 125 87 126
rect 85 125 86 126
rect 84 125 85 126
rect 83 125 84 126
rect 82 125 83 126
rect 81 125 82 126
rect 80 125 81 126
rect 79 125 80 126
rect 78 125 79 126
rect 77 125 78 126
rect 76 125 77 126
rect 75 125 76 126
rect 74 125 75 126
rect 73 125 74 126
rect 72 125 73 126
rect 71 125 72 126
rect 70 125 71 126
rect 69 125 70 126
rect 62 125 63 126
rect 61 125 62 126
rect 60 125 61 126
rect 59 125 60 126
rect 58 125 59 126
rect 57 125 58 126
rect 56 125 57 126
rect 55 125 56 126
rect 54 125 55 126
rect 53 125 54 126
rect 52 125 53 126
rect 51 125 52 126
rect 50 125 51 126
rect 49 125 50 126
rect 48 125 49 126
rect 47 125 48 126
rect 46 125 47 126
rect 45 125 46 126
rect 44 125 45 126
rect 43 125 44 126
rect 42 125 43 126
rect 41 125 42 126
rect 40 125 41 126
rect 39 125 40 126
rect 38 125 39 126
rect 37 125 38 126
rect 36 125 37 126
rect 35 125 36 126
rect 34 125 35 126
rect 33 125 34 126
rect 32 125 33 126
rect 31 125 32 126
rect 476 126 477 127
rect 475 126 476 127
rect 474 126 475 127
rect 473 126 474 127
rect 472 126 473 127
rect 471 126 472 127
rect 470 126 471 127
rect 442 126 443 127
rect 441 126 442 127
rect 440 126 441 127
rect 439 126 440 127
rect 438 126 439 127
rect 295 126 296 127
rect 294 126 295 127
rect 293 126 294 127
rect 292 126 293 127
rect 291 126 292 127
rect 290 126 291 127
rect 289 126 290 127
rect 288 126 289 127
rect 287 126 288 127
rect 286 126 287 127
rect 285 126 286 127
rect 284 126 285 127
rect 283 126 284 127
rect 282 126 283 127
rect 281 126 282 127
rect 280 126 281 127
rect 279 126 280 127
rect 278 126 279 127
rect 236 126 237 127
rect 235 126 236 127
rect 234 126 235 127
rect 233 126 234 127
rect 232 126 233 127
rect 231 126 232 127
rect 230 126 231 127
rect 229 126 230 127
rect 228 126 229 127
rect 227 126 228 127
rect 226 126 227 127
rect 225 126 226 127
rect 224 126 225 127
rect 223 126 224 127
rect 222 126 223 127
rect 221 126 222 127
rect 220 126 221 127
rect 219 126 220 127
rect 218 126 219 127
rect 217 126 218 127
rect 216 126 217 127
rect 215 126 216 127
rect 214 126 215 127
rect 213 126 214 127
rect 212 126 213 127
rect 211 126 212 127
rect 210 126 211 127
rect 209 126 210 127
rect 208 126 209 127
rect 207 126 208 127
rect 206 126 207 127
rect 205 126 206 127
rect 204 126 205 127
rect 203 126 204 127
rect 202 126 203 127
rect 201 126 202 127
rect 200 126 201 127
rect 199 126 200 127
rect 198 126 199 127
rect 197 126 198 127
rect 196 126 197 127
rect 195 126 196 127
rect 194 126 195 127
rect 193 126 194 127
rect 192 126 193 127
rect 191 126 192 127
rect 190 126 191 127
rect 189 126 190 127
rect 188 126 189 127
rect 187 126 188 127
rect 186 126 187 127
rect 185 126 186 127
rect 184 126 185 127
rect 183 126 184 127
rect 182 126 183 127
rect 181 126 182 127
rect 180 126 181 127
rect 179 126 180 127
rect 178 126 179 127
rect 177 126 178 127
rect 176 126 177 127
rect 175 126 176 127
rect 174 126 175 127
rect 173 126 174 127
rect 172 126 173 127
rect 171 126 172 127
rect 170 126 171 127
rect 169 126 170 127
rect 152 126 153 127
rect 151 126 152 127
rect 150 126 151 127
rect 149 126 150 127
rect 148 126 149 127
rect 147 126 148 127
rect 146 126 147 127
rect 145 126 146 127
rect 144 126 145 127
rect 143 126 144 127
rect 142 126 143 127
rect 141 126 142 127
rect 140 126 141 127
rect 139 126 140 127
rect 138 126 139 127
rect 137 126 138 127
rect 136 126 137 127
rect 135 126 136 127
rect 134 126 135 127
rect 133 126 134 127
rect 132 126 133 127
rect 131 126 132 127
rect 130 126 131 127
rect 129 126 130 127
rect 128 126 129 127
rect 127 126 128 127
rect 126 126 127 127
rect 125 126 126 127
rect 124 126 125 127
rect 123 126 124 127
rect 122 126 123 127
rect 121 126 122 127
rect 120 126 121 127
rect 119 126 120 127
rect 118 126 119 127
rect 117 126 118 127
rect 116 126 117 127
rect 115 126 116 127
rect 114 126 115 127
rect 113 126 114 127
rect 112 126 113 127
rect 111 126 112 127
rect 110 126 111 127
rect 109 126 110 127
rect 108 126 109 127
rect 107 126 108 127
rect 106 126 107 127
rect 105 126 106 127
rect 104 126 105 127
rect 103 126 104 127
rect 102 126 103 127
rect 101 126 102 127
rect 100 126 101 127
rect 99 126 100 127
rect 98 126 99 127
rect 97 126 98 127
rect 96 126 97 127
rect 95 126 96 127
rect 94 126 95 127
rect 93 126 94 127
rect 92 126 93 127
rect 91 126 92 127
rect 90 126 91 127
rect 89 126 90 127
rect 88 126 89 127
rect 87 126 88 127
rect 86 126 87 127
rect 85 126 86 127
rect 84 126 85 127
rect 83 126 84 127
rect 82 126 83 127
rect 81 126 82 127
rect 80 126 81 127
rect 79 126 80 127
rect 78 126 79 127
rect 77 126 78 127
rect 76 126 77 127
rect 75 126 76 127
rect 74 126 75 127
rect 73 126 74 127
rect 72 126 73 127
rect 71 126 72 127
rect 70 126 71 127
rect 69 126 70 127
rect 68 126 69 127
rect 62 126 63 127
rect 61 126 62 127
rect 60 126 61 127
rect 59 126 60 127
rect 58 126 59 127
rect 57 126 58 127
rect 56 126 57 127
rect 55 126 56 127
rect 54 126 55 127
rect 53 126 54 127
rect 52 126 53 127
rect 51 126 52 127
rect 50 126 51 127
rect 49 126 50 127
rect 48 126 49 127
rect 47 126 48 127
rect 46 126 47 127
rect 45 126 46 127
rect 44 126 45 127
rect 43 126 44 127
rect 42 126 43 127
rect 41 126 42 127
rect 40 126 41 127
rect 39 126 40 127
rect 38 126 39 127
rect 37 126 38 127
rect 36 126 37 127
rect 35 126 36 127
rect 34 126 35 127
rect 33 126 34 127
rect 32 126 33 127
rect 31 126 32 127
rect 477 127 478 128
rect 476 127 477 128
rect 475 127 476 128
rect 474 127 475 128
rect 473 127 474 128
rect 472 127 473 128
rect 471 127 472 128
rect 442 127 443 128
rect 441 127 442 128
rect 440 127 441 128
rect 439 127 440 128
rect 438 127 439 128
rect 297 127 298 128
rect 296 127 297 128
rect 295 127 296 128
rect 294 127 295 128
rect 293 127 294 128
rect 292 127 293 128
rect 291 127 292 128
rect 290 127 291 128
rect 289 127 290 128
rect 288 127 289 128
rect 287 127 288 128
rect 286 127 287 128
rect 285 127 286 128
rect 284 127 285 128
rect 283 127 284 128
rect 282 127 283 128
rect 281 127 282 128
rect 280 127 281 128
rect 279 127 280 128
rect 278 127 279 128
rect 277 127 278 128
rect 276 127 277 128
rect 275 127 276 128
rect 274 127 275 128
rect 235 127 236 128
rect 234 127 235 128
rect 233 127 234 128
rect 232 127 233 128
rect 231 127 232 128
rect 230 127 231 128
rect 229 127 230 128
rect 228 127 229 128
rect 227 127 228 128
rect 226 127 227 128
rect 225 127 226 128
rect 224 127 225 128
rect 223 127 224 128
rect 222 127 223 128
rect 221 127 222 128
rect 220 127 221 128
rect 219 127 220 128
rect 218 127 219 128
rect 217 127 218 128
rect 216 127 217 128
rect 215 127 216 128
rect 214 127 215 128
rect 213 127 214 128
rect 212 127 213 128
rect 211 127 212 128
rect 210 127 211 128
rect 209 127 210 128
rect 208 127 209 128
rect 207 127 208 128
rect 206 127 207 128
rect 205 127 206 128
rect 204 127 205 128
rect 203 127 204 128
rect 202 127 203 128
rect 201 127 202 128
rect 200 127 201 128
rect 199 127 200 128
rect 198 127 199 128
rect 197 127 198 128
rect 196 127 197 128
rect 195 127 196 128
rect 194 127 195 128
rect 193 127 194 128
rect 192 127 193 128
rect 191 127 192 128
rect 190 127 191 128
rect 189 127 190 128
rect 188 127 189 128
rect 187 127 188 128
rect 186 127 187 128
rect 185 127 186 128
rect 184 127 185 128
rect 183 127 184 128
rect 182 127 183 128
rect 181 127 182 128
rect 180 127 181 128
rect 179 127 180 128
rect 178 127 179 128
rect 177 127 178 128
rect 176 127 177 128
rect 175 127 176 128
rect 174 127 175 128
rect 173 127 174 128
rect 172 127 173 128
rect 171 127 172 128
rect 170 127 171 128
rect 169 127 170 128
rect 151 127 152 128
rect 150 127 151 128
rect 149 127 150 128
rect 148 127 149 128
rect 147 127 148 128
rect 146 127 147 128
rect 145 127 146 128
rect 144 127 145 128
rect 143 127 144 128
rect 142 127 143 128
rect 141 127 142 128
rect 140 127 141 128
rect 139 127 140 128
rect 138 127 139 128
rect 137 127 138 128
rect 136 127 137 128
rect 135 127 136 128
rect 134 127 135 128
rect 133 127 134 128
rect 132 127 133 128
rect 131 127 132 128
rect 130 127 131 128
rect 129 127 130 128
rect 128 127 129 128
rect 127 127 128 128
rect 126 127 127 128
rect 125 127 126 128
rect 124 127 125 128
rect 123 127 124 128
rect 122 127 123 128
rect 121 127 122 128
rect 120 127 121 128
rect 119 127 120 128
rect 118 127 119 128
rect 117 127 118 128
rect 116 127 117 128
rect 115 127 116 128
rect 114 127 115 128
rect 113 127 114 128
rect 112 127 113 128
rect 111 127 112 128
rect 110 127 111 128
rect 109 127 110 128
rect 108 127 109 128
rect 107 127 108 128
rect 106 127 107 128
rect 105 127 106 128
rect 104 127 105 128
rect 103 127 104 128
rect 102 127 103 128
rect 101 127 102 128
rect 100 127 101 128
rect 99 127 100 128
rect 98 127 99 128
rect 97 127 98 128
rect 96 127 97 128
rect 95 127 96 128
rect 94 127 95 128
rect 93 127 94 128
rect 92 127 93 128
rect 91 127 92 128
rect 90 127 91 128
rect 89 127 90 128
rect 88 127 89 128
rect 87 127 88 128
rect 86 127 87 128
rect 85 127 86 128
rect 84 127 85 128
rect 83 127 84 128
rect 82 127 83 128
rect 81 127 82 128
rect 80 127 81 128
rect 79 127 80 128
rect 78 127 79 128
rect 77 127 78 128
rect 76 127 77 128
rect 75 127 76 128
rect 74 127 75 128
rect 73 127 74 128
rect 72 127 73 128
rect 71 127 72 128
rect 70 127 71 128
rect 69 127 70 128
rect 68 127 69 128
rect 61 127 62 128
rect 60 127 61 128
rect 59 127 60 128
rect 58 127 59 128
rect 57 127 58 128
rect 56 127 57 128
rect 55 127 56 128
rect 54 127 55 128
rect 53 127 54 128
rect 52 127 53 128
rect 51 127 52 128
rect 50 127 51 128
rect 49 127 50 128
rect 48 127 49 128
rect 47 127 48 128
rect 46 127 47 128
rect 45 127 46 128
rect 44 127 45 128
rect 43 127 44 128
rect 42 127 43 128
rect 41 127 42 128
rect 40 127 41 128
rect 39 127 40 128
rect 38 127 39 128
rect 37 127 38 128
rect 36 127 37 128
rect 35 127 36 128
rect 34 127 35 128
rect 33 127 34 128
rect 32 127 33 128
rect 31 127 32 128
rect 479 128 480 129
rect 478 128 479 129
rect 477 128 478 129
rect 476 128 477 129
rect 475 128 476 129
rect 474 128 475 129
rect 473 128 474 129
rect 472 128 473 129
rect 462 128 463 129
rect 442 128 443 129
rect 441 128 442 129
rect 440 128 441 129
rect 439 128 440 129
rect 438 128 439 129
rect 299 128 300 129
rect 298 128 299 129
rect 297 128 298 129
rect 296 128 297 129
rect 295 128 296 129
rect 294 128 295 129
rect 293 128 294 129
rect 292 128 293 129
rect 291 128 292 129
rect 290 128 291 129
rect 289 128 290 129
rect 288 128 289 129
rect 287 128 288 129
rect 286 128 287 129
rect 285 128 286 129
rect 284 128 285 129
rect 283 128 284 129
rect 282 128 283 129
rect 281 128 282 129
rect 280 128 281 129
rect 279 128 280 129
rect 278 128 279 129
rect 277 128 278 129
rect 276 128 277 129
rect 275 128 276 129
rect 274 128 275 129
rect 273 128 274 129
rect 272 128 273 129
rect 271 128 272 129
rect 234 128 235 129
rect 233 128 234 129
rect 232 128 233 129
rect 231 128 232 129
rect 230 128 231 129
rect 229 128 230 129
rect 228 128 229 129
rect 227 128 228 129
rect 226 128 227 129
rect 225 128 226 129
rect 224 128 225 129
rect 223 128 224 129
rect 222 128 223 129
rect 221 128 222 129
rect 220 128 221 129
rect 219 128 220 129
rect 218 128 219 129
rect 217 128 218 129
rect 216 128 217 129
rect 215 128 216 129
rect 214 128 215 129
rect 213 128 214 129
rect 212 128 213 129
rect 211 128 212 129
rect 210 128 211 129
rect 209 128 210 129
rect 208 128 209 129
rect 207 128 208 129
rect 206 128 207 129
rect 205 128 206 129
rect 204 128 205 129
rect 203 128 204 129
rect 202 128 203 129
rect 201 128 202 129
rect 200 128 201 129
rect 199 128 200 129
rect 198 128 199 129
rect 197 128 198 129
rect 196 128 197 129
rect 195 128 196 129
rect 194 128 195 129
rect 193 128 194 129
rect 192 128 193 129
rect 191 128 192 129
rect 190 128 191 129
rect 189 128 190 129
rect 188 128 189 129
rect 187 128 188 129
rect 186 128 187 129
rect 185 128 186 129
rect 184 128 185 129
rect 183 128 184 129
rect 182 128 183 129
rect 181 128 182 129
rect 180 128 181 129
rect 179 128 180 129
rect 178 128 179 129
rect 177 128 178 129
rect 176 128 177 129
rect 175 128 176 129
rect 174 128 175 129
rect 173 128 174 129
rect 172 128 173 129
rect 171 128 172 129
rect 170 128 171 129
rect 169 128 170 129
rect 168 128 169 129
rect 151 128 152 129
rect 150 128 151 129
rect 149 128 150 129
rect 148 128 149 129
rect 147 128 148 129
rect 146 128 147 129
rect 145 128 146 129
rect 144 128 145 129
rect 143 128 144 129
rect 142 128 143 129
rect 141 128 142 129
rect 140 128 141 129
rect 139 128 140 129
rect 138 128 139 129
rect 137 128 138 129
rect 136 128 137 129
rect 135 128 136 129
rect 134 128 135 129
rect 133 128 134 129
rect 132 128 133 129
rect 131 128 132 129
rect 130 128 131 129
rect 129 128 130 129
rect 128 128 129 129
rect 127 128 128 129
rect 126 128 127 129
rect 125 128 126 129
rect 124 128 125 129
rect 123 128 124 129
rect 122 128 123 129
rect 121 128 122 129
rect 120 128 121 129
rect 119 128 120 129
rect 118 128 119 129
rect 117 128 118 129
rect 116 128 117 129
rect 115 128 116 129
rect 114 128 115 129
rect 113 128 114 129
rect 112 128 113 129
rect 111 128 112 129
rect 110 128 111 129
rect 109 128 110 129
rect 108 128 109 129
rect 107 128 108 129
rect 106 128 107 129
rect 105 128 106 129
rect 104 128 105 129
rect 103 128 104 129
rect 102 128 103 129
rect 101 128 102 129
rect 100 128 101 129
rect 99 128 100 129
rect 98 128 99 129
rect 97 128 98 129
rect 96 128 97 129
rect 95 128 96 129
rect 94 128 95 129
rect 93 128 94 129
rect 92 128 93 129
rect 91 128 92 129
rect 90 128 91 129
rect 89 128 90 129
rect 88 128 89 129
rect 87 128 88 129
rect 86 128 87 129
rect 85 128 86 129
rect 84 128 85 129
rect 83 128 84 129
rect 82 128 83 129
rect 81 128 82 129
rect 80 128 81 129
rect 79 128 80 129
rect 78 128 79 129
rect 77 128 78 129
rect 76 128 77 129
rect 75 128 76 129
rect 74 128 75 129
rect 73 128 74 129
rect 72 128 73 129
rect 71 128 72 129
rect 70 128 71 129
rect 69 128 70 129
rect 68 128 69 129
rect 67 128 68 129
rect 61 128 62 129
rect 60 128 61 129
rect 59 128 60 129
rect 58 128 59 129
rect 57 128 58 129
rect 56 128 57 129
rect 55 128 56 129
rect 54 128 55 129
rect 53 128 54 129
rect 52 128 53 129
rect 51 128 52 129
rect 50 128 51 129
rect 49 128 50 129
rect 48 128 49 129
rect 47 128 48 129
rect 46 128 47 129
rect 45 128 46 129
rect 44 128 45 129
rect 43 128 44 129
rect 42 128 43 129
rect 41 128 42 129
rect 40 128 41 129
rect 39 128 40 129
rect 38 128 39 129
rect 37 128 38 129
rect 36 128 37 129
rect 35 128 36 129
rect 34 128 35 129
rect 33 128 34 129
rect 32 128 33 129
rect 31 128 32 129
rect 480 129 481 130
rect 479 129 480 130
rect 478 129 479 130
rect 477 129 478 130
rect 476 129 477 130
rect 475 129 476 130
rect 474 129 475 130
rect 473 129 474 130
rect 462 129 463 130
rect 442 129 443 130
rect 441 129 442 130
rect 440 129 441 130
rect 439 129 440 130
rect 438 129 439 130
rect 301 129 302 130
rect 300 129 301 130
rect 299 129 300 130
rect 298 129 299 130
rect 297 129 298 130
rect 296 129 297 130
rect 295 129 296 130
rect 294 129 295 130
rect 293 129 294 130
rect 292 129 293 130
rect 291 129 292 130
rect 290 129 291 130
rect 289 129 290 130
rect 288 129 289 130
rect 287 129 288 130
rect 286 129 287 130
rect 285 129 286 130
rect 284 129 285 130
rect 283 129 284 130
rect 282 129 283 130
rect 281 129 282 130
rect 280 129 281 130
rect 279 129 280 130
rect 278 129 279 130
rect 277 129 278 130
rect 276 129 277 130
rect 275 129 276 130
rect 274 129 275 130
rect 273 129 274 130
rect 272 129 273 130
rect 271 129 272 130
rect 270 129 271 130
rect 269 129 270 130
rect 268 129 269 130
rect 233 129 234 130
rect 232 129 233 130
rect 231 129 232 130
rect 230 129 231 130
rect 229 129 230 130
rect 228 129 229 130
rect 227 129 228 130
rect 226 129 227 130
rect 225 129 226 130
rect 224 129 225 130
rect 223 129 224 130
rect 222 129 223 130
rect 221 129 222 130
rect 220 129 221 130
rect 219 129 220 130
rect 218 129 219 130
rect 217 129 218 130
rect 216 129 217 130
rect 215 129 216 130
rect 214 129 215 130
rect 213 129 214 130
rect 212 129 213 130
rect 211 129 212 130
rect 210 129 211 130
rect 209 129 210 130
rect 208 129 209 130
rect 207 129 208 130
rect 206 129 207 130
rect 205 129 206 130
rect 204 129 205 130
rect 203 129 204 130
rect 202 129 203 130
rect 201 129 202 130
rect 200 129 201 130
rect 199 129 200 130
rect 198 129 199 130
rect 197 129 198 130
rect 196 129 197 130
rect 195 129 196 130
rect 194 129 195 130
rect 193 129 194 130
rect 192 129 193 130
rect 191 129 192 130
rect 190 129 191 130
rect 189 129 190 130
rect 188 129 189 130
rect 187 129 188 130
rect 186 129 187 130
rect 185 129 186 130
rect 184 129 185 130
rect 183 129 184 130
rect 182 129 183 130
rect 181 129 182 130
rect 180 129 181 130
rect 179 129 180 130
rect 178 129 179 130
rect 177 129 178 130
rect 176 129 177 130
rect 175 129 176 130
rect 174 129 175 130
rect 173 129 174 130
rect 172 129 173 130
rect 171 129 172 130
rect 170 129 171 130
rect 169 129 170 130
rect 168 129 169 130
rect 150 129 151 130
rect 149 129 150 130
rect 148 129 149 130
rect 147 129 148 130
rect 146 129 147 130
rect 145 129 146 130
rect 144 129 145 130
rect 143 129 144 130
rect 142 129 143 130
rect 141 129 142 130
rect 140 129 141 130
rect 139 129 140 130
rect 138 129 139 130
rect 137 129 138 130
rect 136 129 137 130
rect 135 129 136 130
rect 134 129 135 130
rect 133 129 134 130
rect 132 129 133 130
rect 131 129 132 130
rect 130 129 131 130
rect 129 129 130 130
rect 128 129 129 130
rect 127 129 128 130
rect 126 129 127 130
rect 125 129 126 130
rect 124 129 125 130
rect 123 129 124 130
rect 122 129 123 130
rect 121 129 122 130
rect 120 129 121 130
rect 119 129 120 130
rect 118 129 119 130
rect 117 129 118 130
rect 116 129 117 130
rect 115 129 116 130
rect 114 129 115 130
rect 113 129 114 130
rect 112 129 113 130
rect 111 129 112 130
rect 110 129 111 130
rect 109 129 110 130
rect 108 129 109 130
rect 107 129 108 130
rect 106 129 107 130
rect 105 129 106 130
rect 104 129 105 130
rect 103 129 104 130
rect 102 129 103 130
rect 101 129 102 130
rect 100 129 101 130
rect 99 129 100 130
rect 98 129 99 130
rect 97 129 98 130
rect 96 129 97 130
rect 95 129 96 130
rect 94 129 95 130
rect 93 129 94 130
rect 92 129 93 130
rect 91 129 92 130
rect 90 129 91 130
rect 89 129 90 130
rect 88 129 89 130
rect 87 129 88 130
rect 86 129 87 130
rect 85 129 86 130
rect 84 129 85 130
rect 83 129 84 130
rect 82 129 83 130
rect 81 129 82 130
rect 80 129 81 130
rect 79 129 80 130
rect 78 129 79 130
rect 77 129 78 130
rect 76 129 77 130
rect 75 129 76 130
rect 74 129 75 130
rect 73 129 74 130
rect 72 129 73 130
rect 71 129 72 130
rect 70 129 71 130
rect 69 129 70 130
rect 68 129 69 130
rect 67 129 68 130
rect 61 129 62 130
rect 60 129 61 130
rect 59 129 60 130
rect 58 129 59 130
rect 57 129 58 130
rect 56 129 57 130
rect 55 129 56 130
rect 54 129 55 130
rect 53 129 54 130
rect 52 129 53 130
rect 51 129 52 130
rect 50 129 51 130
rect 49 129 50 130
rect 48 129 49 130
rect 47 129 48 130
rect 46 129 47 130
rect 45 129 46 130
rect 44 129 45 130
rect 43 129 44 130
rect 42 129 43 130
rect 41 129 42 130
rect 40 129 41 130
rect 39 129 40 130
rect 38 129 39 130
rect 37 129 38 130
rect 36 129 37 130
rect 35 129 36 130
rect 34 129 35 130
rect 33 129 34 130
rect 32 129 33 130
rect 481 130 482 131
rect 480 130 481 131
rect 479 130 480 131
rect 478 130 479 131
rect 477 130 478 131
rect 476 130 477 131
rect 475 130 476 131
rect 474 130 475 131
rect 462 130 463 131
rect 442 130 443 131
rect 441 130 442 131
rect 440 130 441 131
rect 439 130 440 131
rect 438 130 439 131
rect 302 130 303 131
rect 301 130 302 131
rect 300 130 301 131
rect 299 130 300 131
rect 298 130 299 131
rect 297 130 298 131
rect 296 130 297 131
rect 295 130 296 131
rect 294 130 295 131
rect 293 130 294 131
rect 292 130 293 131
rect 291 130 292 131
rect 290 130 291 131
rect 289 130 290 131
rect 288 130 289 131
rect 287 130 288 131
rect 286 130 287 131
rect 285 130 286 131
rect 284 130 285 131
rect 283 130 284 131
rect 282 130 283 131
rect 281 130 282 131
rect 280 130 281 131
rect 279 130 280 131
rect 278 130 279 131
rect 277 130 278 131
rect 276 130 277 131
rect 275 130 276 131
rect 274 130 275 131
rect 273 130 274 131
rect 272 130 273 131
rect 271 130 272 131
rect 270 130 271 131
rect 269 130 270 131
rect 268 130 269 131
rect 267 130 268 131
rect 266 130 267 131
rect 232 130 233 131
rect 231 130 232 131
rect 230 130 231 131
rect 229 130 230 131
rect 228 130 229 131
rect 227 130 228 131
rect 226 130 227 131
rect 225 130 226 131
rect 224 130 225 131
rect 223 130 224 131
rect 222 130 223 131
rect 221 130 222 131
rect 220 130 221 131
rect 219 130 220 131
rect 218 130 219 131
rect 217 130 218 131
rect 216 130 217 131
rect 215 130 216 131
rect 214 130 215 131
rect 213 130 214 131
rect 212 130 213 131
rect 211 130 212 131
rect 210 130 211 131
rect 209 130 210 131
rect 208 130 209 131
rect 207 130 208 131
rect 206 130 207 131
rect 205 130 206 131
rect 204 130 205 131
rect 203 130 204 131
rect 202 130 203 131
rect 201 130 202 131
rect 200 130 201 131
rect 199 130 200 131
rect 198 130 199 131
rect 197 130 198 131
rect 196 130 197 131
rect 195 130 196 131
rect 194 130 195 131
rect 193 130 194 131
rect 192 130 193 131
rect 191 130 192 131
rect 190 130 191 131
rect 189 130 190 131
rect 188 130 189 131
rect 187 130 188 131
rect 186 130 187 131
rect 185 130 186 131
rect 184 130 185 131
rect 183 130 184 131
rect 182 130 183 131
rect 181 130 182 131
rect 180 130 181 131
rect 179 130 180 131
rect 178 130 179 131
rect 177 130 178 131
rect 176 130 177 131
rect 175 130 176 131
rect 174 130 175 131
rect 173 130 174 131
rect 172 130 173 131
rect 171 130 172 131
rect 170 130 171 131
rect 169 130 170 131
rect 168 130 169 131
rect 167 130 168 131
rect 150 130 151 131
rect 149 130 150 131
rect 148 130 149 131
rect 147 130 148 131
rect 146 130 147 131
rect 145 130 146 131
rect 144 130 145 131
rect 143 130 144 131
rect 142 130 143 131
rect 141 130 142 131
rect 140 130 141 131
rect 139 130 140 131
rect 138 130 139 131
rect 137 130 138 131
rect 136 130 137 131
rect 135 130 136 131
rect 134 130 135 131
rect 133 130 134 131
rect 132 130 133 131
rect 131 130 132 131
rect 130 130 131 131
rect 129 130 130 131
rect 128 130 129 131
rect 127 130 128 131
rect 126 130 127 131
rect 125 130 126 131
rect 124 130 125 131
rect 123 130 124 131
rect 122 130 123 131
rect 121 130 122 131
rect 120 130 121 131
rect 119 130 120 131
rect 118 130 119 131
rect 117 130 118 131
rect 116 130 117 131
rect 115 130 116 131
rect 114 130 115 131
rect 113 130 114 131
rect 112 130 113 131
rect 111 130 112 131
rect 110 130 111 131
rect 109 130 110 131
rect 108 130 109 131
rect 107 130 108 131
rect 106 130 107 131
rect 105 130 106 131
rect 104 130 105 131
rect 103 130 104 131
rect 102 130 103 131
rect 101 130 102 131
rect 100 130 101 131
rect 99 130 100 131
rect 98 130 99 131
rect 97 130 98 131
rect 96 130 97 131
rect 95 130 96 131
rect 94 130 95 131
rect 93 130 94 131
rect 92 130 93 131
rect 91 130 92 131
rect 90 130 91 131
rect 89 130 90 131
rect 88 130 89 131
rect 87 130 88 131
rect 86 130 87 131
rect 85 130 86 131
rect 84 130 85 131
rect 83 130 84 131
rect 82 130 83 131
rect 81 130 82 131
rect 80 130 81 131
rect 79 130 80 131
rect 78 130 79 131
rect 77 130 78 131
rect 76 130 77 131
rect 75 130 76 131
rect 74 130 75 131
rect 73 130 74 131
rect 72 130 73 131
rect 71 130 72 131
rect 70 130 71 131
rect 69 130 70 131
rect 68 130 69 131
rect 67 130 68 131
rect 66 130 67 131
rect 61 130 62 131
rect 60 130 61 131
rect 59 130 60 131
rect 58 130 59 131
rect 57 130 58 131
rect 56 130 57 131
rect 55 130 56 131
rect 54 130 55 131
rect 53 130 54 131
rect 52 130 53 131
rect 51 130 52 131
rect 50 130 51 131
rect 49 130 50 131
rect 48 130 49 131
rect 47 130 48 131
rect 46 130 47 131
rect 45 130 46 131
rect 44 130 45 131
rect 43 130 44 131
rect 42 130 43 131
rect 41 130 42 131
rect 40 130 41 131
rect 39 130 40 131
rect 38 130 39 131
rect 37 130 38 131
rect 36 130 37 131
rect 35 130 36 131
rect 34 130 35 131
rect 33 130 34 131
rect 32 130 33 131
rect 482 131 483 132
rect 481 131 482 132
rect 480 131 481 132
rect 479 131 480 132
rect 478 131 479 132
rect 477 131 478 132
rect 476 131 477 132
rect 475 131 476 132
rect 464 131 465 132
rect 463 131 464 132
rect 462 131 463 132
rect 442 131 443 132
rect 441 131 442 132
rect 440 131 441 132
rect 439 131 440 132
rect 438 131 439 132
rect 304 131 305 132
rect 303 131 304 132
rect 302 131 303 132
rect 301 131 302 132
rect 300 131 301 132
rect 299 131 300 132
rect 298 131 299 132
rect 297 131 298 132
rect 296 131 297 132
rect 295 131 296 132
rect 294 131 295 132
rect 293 131 294 132
rect 292 131 293 132
rect 291 131 292 132
rect 290 131 291 132
rect 289 131 290 132
rect 288 131 289 132
rect 287 131 288 132
rect 286 131 287 132
rect 285 131 286 132
rect 284 131 285 132
rect 283 131 284 132
rect 282 131 283 132
rect 281 131 282 132
rect 280 131 281 132
rect 279 131 280 132
rect 278 131 279 132
rect 277 131 278 132
rect 276 131 277 132
rect 275 131 276 132
rect 274 131 275 132
rect 273 131 274 132
rect 272 131 273 132
rect 271 131 272 132
rect 270 131 271 132
rect 269 131 270 132
rect 268 131 269 132
rect 267 131 268 132
rect 266 131 267 132
rect 265 131 266 132
rect 264 131 265 132
rect 232 131 233 132
rect 231 131 232 132
rect 230 131 231 132
rect 229 131 230 132
rect 228 131 229 132
rect 227 131 228 132
rect 226 131 227 132
rect 225 131 226 132
rect 224 131 225 132
rect 223 131 224 132
rect 222 131 223 132
rect 221 131 222 132
rect 220 131 221 132
rect 219 131 220 132
rect 218 131 219 132
rect 217 131 218 132
rect 216 131 217 132
rect 215 131 216 132
rect 214 131 215 132
rect 213 131 214 132
rect 212 131 213 132
rect 211 131 212 132
rect 210 131 211 132
rect 209 131 210 132
rect 208 131 209 132
rect 207 131 208 132
rect 206 131 207 132
rect 205 131 206 132
rect 204 131 205 132
rect 203 131 204 132
rect 202 131 203 132
rect 201 131 202 132
rect 200 131 201 132
rect 199 131 200 132
rect 198 131 199 132
rect 197 131 198 132
rect 196 131 197 132
rect 195 131 196 132
rect 194 131 195 132
rect 193 131 194 132
rect 192 131 193 132
rect 191 131 192 132
rect 190 131 191 132
rect 189 131 190 132
rect 188 131 189 132
rect 187 131 188 132
rect 186 131 187 132
rect 185 131 186 132
rect 184 131 185 132
rect 183 131 184 132
rect 182 131 183 132
rect 181 131 182 132
rect 180 131 181 132
rect 179 131 180 132
rect 178 131 179 132
rect 177 131 178 132
rect 176 131 177 132
rect 175 131 176 132
rect 174 131 175 132
rect 173 131 174 132
rect 172 131 173 132
rect 171 131 172 132
rect 170 131 171 132
rect 169 131 170 132
rect 168 131 169 132
rect 167 131 168 132
rect 149 131 150 132
rect 148 131 149 132
rect 147 131 148 132
rect 146 131 147 132
rect 145 131 146 132
rect 144 131 145 132
rect 143 131 144 132
rect 142 131 143 132
rect 141 131 142 132
rect 140 131 141 132
rect 139 131 140 132
rect 138 131 139 132
rect 137 131 138 132
rect 136 131 137 132
rect 135 131 136 132
rect 134 131 135 132
rect 133 131 134 132
rect 132 131 133 132
rect 131 131 132 132
rect 130 131 131 132
rect 129 131 130 132
rect 128 131 129 132
rect 127 131 128 132
rect 126 131 127 132
rect 125 131 126 132
rect 124 131 125 132
rect 123 131 124 132
rect 122 131 123 132
rect 121 131 122 132
rect 120 131 121 132
rect 119 131 120 132
rect 118 131 119 132
rect 117 131 118 132
rect 116 131 117 132
rect 115 131 116 132
rect 114 131 115 132
rect 113 131 114 132
rect 112 131 113 132
rect 111 131 112 132
rect 110 131 111 132
rect 109 131 110 132
rect 108 131 109 132
rect 107 131 108 132
rect 106 131 107 132
rect 105 131 106 132
rect 104 131 105 132
rect 103 131 104 132
rect 102 131 103 132
rect 101 131 102 132
rect 100 131 101 132
rect 99 131 100 132
rect 98 131 99 132
rect 97 131 98 132
rect 96 131 97 132
rect 95 131 96 132
rect 94 131 95 132
rect 93 131 94 132
rect 92 131 93 132
rect 91 131 92 132
rect 90 131 91 132
rect 89 131 90 132
rect 88 131 89 132
rect 87 131 88 132
rect 86 131 87 132
rect 85 131 86 132
rect 84 131 85 132
rect 83 131 84 132
rect 82 131 83 132
rect 81 131 82 132
rect 80 131 81 132
rect 79 131 80 132
rect 78 131 79 132
rect 77 131 78 132
rect 76 131 77 132
rect 75 131 76 132
rect 74 131 75 132
rect 73 131 74 132
rect 72 131 73 132
rect 71 131 72 132
rect 70 131 71 132
rect 69 131 70 132
rect 68 131 69 132
rect 67 131 68 132
rect 66 131 67 132
rect 65 131 66 132
rect 61 131 62 132
rect 60 131 61 132
rect 59 131 60 132
rect 58 131 59 132
rect 57 131 58 132
rect 56 131 57 132
rect 55 131 56 132
rect 54 131 55 132
rect 53 131 54 132
rect 52 131 53 132
rect 51 131 52 132
rect 50 131 51 132
rect 49 131 50 132
rect 48 131 49 132
rect 47 131 48 132
rect 46 131 47 132
rect 45 131 46 132
rect 44 131 45 132
rect 43 131 44 132
rect 42 131 43 132
rect 41 131 42 132
rect 40 131 41 132
rect 39 131 40 132
rect 38 131 39 132
rect 37 131 38 132
rect 36 131 37 132
rect 35 131 36 132
rect 34 131 35 132
rect 33 131 34 132
rect 32 131 33 132
rect 483 132 484 133
rect 482 132 483 133
rect 481 132 482 133
rect 480 132 481 133
rect 479 132 480 133
rect 478 132 479 133
rect 477 132 478 133
rect 476 132 477 133
rect 475 132 476 133
rect 474 132 475 133
rect 473 132 474 133
rect 472 132 473 133
rect 471 132 472 133
rect 470 132 471 133
rect 469 132 470 133
rect 468 132 469 133
rect 467 132 468 133
rect 466 132 467 133
rect 465 132 466 133
rect 464 132 465 133
rect 463 132 464 133
rect 462 132 463 133
rect 442 132 443 133
rect 441 132 442 133
rect 440 132 441 133
rect 439 132 440 133
rect 438 132 439 133
rect 305 132 306 133
rect 304 132 305 133
rect 303 132 304 133
rect 302 132 303 133
rect 301 132 302 133
rect 300 132 301 133
rect 299 132 300 133
rect 298 132 299 133
rect 297 132 298 133
rect 296 132 297 133
rect 295 132 296 133
rect 294 132 295 133
rect 293 132 294 133
rect 292 132 293 133
rect 291 132 292 133
rect 290 132 291 133
rect 289 132 290 133
rect 288 132 289 133
rect 287 132 288 133
rect 286 132 287 133
rect 285 132 286 133
rect 284 132 285 133
rect 283 132 284 133
rect 282 132 283 133
rect 281 132 282 133
rect 280 132 281 133
rect 279 132 280 133
rect 278 132 279 133
rect 277 132 278 133
rect 276 132 277 133
rect 275 132 276 133
rect 274 132 275 133
rect 273 132 274 133
rect 272 132 273 133
rect 271 132 272 133
rect 270 132 271 133
rect 269 132 270 133
rect 268 132 269 133
rect 267 132 268 133
rect 266 132 267 133
rect 265 132 266 133
rect 264 132 265 133
rect 263 132 264 133
rect 262 132 263 133
rect 231 132 232 133
rect 230 132 231 133
rect 229 132 230 133
rect 228 132 229 133
rect 227 132 228 133
rect 226 132 227 133
rect 225 132 226 133
rect 224 132 225 133
rect 223 132 224 133
rect 222 132 223 133
rect 221 132 222 133
rect 220 132 221 133
rect 219 132 220 133
rect 218 132 219 133
rect 217 132 218 133
rect 216 132 217 133
rect 215 132 216 133
rect 214 132 215 133
rect 213 132 214 133
rect 212 132 213 133
rect 211 132 212 133
rect 210 132 211 133
rect 209 132 210 133
rect 208 132 209 133
rect 207 132 208 133
rect 206 132 207 133
rect 205 132 206 133
rect 204 132 205 133
rect 203 132 204 133
rect 202 132 203 133
rect 201 132 202 133
rect 200 132 201 133
rect 199 132 200 133
rect 198 132 199 133
rect 197 132 198 133
rect 196 132 197 133
rect 195 132 196 133
rect 194 132 195 133
rect 193 132 194 133
rect 192 132 193 133
rect 191 132 192 133
rect 190 132 191 133
rect 189 132 190 133
rect 188 132 189 133
rect 187 132 188 133
rect 186 132 187 133
rect 185 132 186 133
rect 184 132 185 133
rect 183 132 184 133
rect 182 132 183 133
rect 181 132 182 133
rect 180 132 181 133
rect 179 132 180 133
rect 178 132 179 133
rect 177 132 178 133
rect 176 132 177 133
rect 175 132 176 133
rect 174 132 175 133
rect 173 132 174 133
rect 172 132 173 133
rect 171 132 172 133
rect 170 132 171 133
rect 169 132 170 133
rect 168 132 169 133
rect 167 132 168 133
rect 166 132 167 133
rect 149 132 150 133
rect 148 132 149 133
rect 147 132 148 133
rect 146 132 147 133
rect 145 132 146 133
rect 144 132 145 133
rect 143 132 144 133
rect 142 132 143 133
rect 141 132 142 133
rect 140 132 141 133
rect 139 132 140 133
rect 138 132 139 133
rect 137 132 138 133
rect 136 132 137 133
rect 135 132 136 133
rect 134 132 135 133
rect 133 132 134 133
rect 132 132 133 133
rect 131 132 132 133
rect 130 132 131 133
rect 129 132 130 133
rect 128 132 129 133
rect 127 132 128 133
rect 126 132 127 133
rect 125 132 126 133
rect 124 132 125 133
rect 123 132 124 133
rect 122 132 123 133
rect 121 132 122 133
rect 120 132 121 133
rect 119 132 120 133
rect 118 132 119 133
rect 117 132 118 133
rect 116 132 117 133
rect 115 132 116 133
rect 114 132 115 133
rect 113 132 114 133
rect 112 132 113 133
rect 111 132 112 133
rect 110 132 111 133
rect 109 132 110 133
rect 108 132 109 133
rect 107 132 108 133
rect 106 132 107 133
rect 105 132 106 133
rect 104 132 105 133
rect 103 132 104 133
rect 102 132 103 133
rect 101 132 102 133
rect 100 132 101 133
rect 99 132 100 133
rect 98 132 99 133
rect 97 132 98 133
rect 96 132 97 133
rect 95 132 96 133
rect 94 132 95 133
rect 93 132 94 133
rect 92 132 93 133
rect 91 132 92 133
rect 90 132 91 133
rect 89 132 90 133
rect 88 132 89 133
rect 87 132 88 133
rect 86 132 87 133
rect 85 132 86 133
rect 84 132 85 133
rect 83 132 84 133
rect 82 132 83 133
rect 81 132 82 133
rect 80 132 81 133
rect 79 132 80 133
rect 78 132 79 133
rect 77 132 78 133
rect 76 132 77 133
rect 75 132 76 133
rect 74 132 75 133
rect 73 132 74 133
rect 72 132 73 133
rect 71 132 72 133
rect 70 132 71 133
rect 69 132 70 133
rect 68 132 69 133
rect 67 132 68 133
rect 66 132 67 133
rect 65 132 66 133
rect 60 132 61 133
rect 59 132 60 133
rect 58 132 59 133
rect 57 132 58 133
rect 56 132 57 133
rect 55 132 56 133
rect 54 132 55 133
rect 53 132 54 133
rect 52 132 53 133
rect 51 132 52 133
rect 50 132 51 133
rect 49 132 50 133
rect 48 132 49 133
rect 47 132 48 133
rect 46 132 47 133
rect 45 132 46 133
rect 44 132 45 133
rect 43 132 44 133
rect 42 132 43 133
rect 41 132 42 133
rect 40 132 41 133
rect 39 132 40 133
rect 38 132 39 133
rect 37 132 38 133
rect 36 132 37 133
rect 35 132 36 133
rect 34 132 35 133
rect 33 132 34 133
rect 483 133 484 134
rect 482 133 483 134
rect 481 133 482 134
rect 480 133 481 134
rect 479 133 480 134
rect 478 133 479 134
rect 477 133 478 134
rect 476 133 477 134
rect 475 133 476 134
rect 474 133 475 134
rect 473 133 474 134
rect 472 133 473 134
rect 471 133 472 134
rect 470 133 471 134
rect 469 133 470 134
rect 468 133 469 134
rect 467 133 468 134
rect 466 133 467 134
rect 465 133 466 134
rect 464 133 465 134
rect 463 133 464 134
rect 462 133 463 134
rect 442 133 443 134
rect 441 133 442 134
rect 440 133 441 134
rect 439 133 440 134
rect 438 133 439 134
rect 306 133 307 134
rect 305 133 306 134
rect 304 133 305 134
rect 303 133 304 134
rect 302 133 303 134
rect 301 133 302 134
rect 300 133 301 134
rect 299 133 300 134
rect 298 133 299 134
rect 297 133 298 134
rect 296 133 297 134
rect 295 133 296 134
rect 294 133 295 134
rect 293 133 294 134
rect 292 133 293 134
rect 291 133 292 134
rect 290 133 291 134
rect 289 133 290 134
rect 288 133 289 134
rect 287 133 288 134
rect 286 133 287 134
rect 285 133 286 134
rect 284 133 285 134
rect 283 133 284 134
rect 282 133 283 134
rect 281 133 282 134
rect 280 133 281 134
rect 279 133 280 134
rect 278 133 279 134
rect 277 133 278 134
rect 276 133 277 134
rect 275 133 276 134
rect 274 133 275 134
rect 273 133 274 134
rect 272 133 273 134
rect 271 133 272 134
rect 270 133 271 134
rect 269 133 270 134
rect 268 133 269 134
rect 267 133 268 134
rect 266 133 267 134
rect 265 133 266 134
rect 264 133 265 134
rect 263 133 264 134
rect 262 133 263 134
rect 261 133 262 134
rect 260 133 261 134
rect 230 133 231 134
rect 229 133 230 134
rect 228 133 229 134
rect 227 133 228 134
rect 226 133 227 134
rect 225 133 226 134
rect 224 133 225 134
rect 223 133 224 134
rect 222 133 223 134
rect 221 133 222 134
rect 220 133 221 134
rect 219 133 220 134
rect 218 133 219 134
rect 217 133 218 134
rect 216 133 217 134
rect 215 133 216 134
rect 214 133 215 134
rect 213 133 214 134
rect 212 133 213 134
rect 211 133 212 134
rect 210 133 211 134
rect 209 133 210 134
rect 208 133 209 134
rect 207 133 208 134
rect 206 133 207 134
rect 205 133 206 134
rect 204 133 205 134
rect 203 133 204 134
rect 202 133 203 134
rect 201 133 202 134
rect 200 133 201 134
rect 199 133 200 134
rect 198 133 199 134
rect 197 133 198 134
rect 196 133 197 134
rect 195 133 196 134
rect 194 133 195 134
rect 193 133 194 134
rect 192 133 193 134
rect 191 133 192 134
rect 190 133 191 134
rect 189 133 190 134
rect 188 133 189 134
rect 187 133 188 134
rect 186 133 187 134
rect 185 133 186 134
rect 184 133 185 134
rect 183 133 184 134
rect 182 133 183 134
rect 181 133 182 134
rect 180 133 181 134
rect 179 133 180 134
rect 178 133 179 134
rect 177 133 178 134
rect 176 133 177 134
rect 175 133 176 134
rect 174 133 175 134
rect 173 133 174 134
rect 172 133 173 134
rect 171 133 172 134
rect 170 133 171 134
rect 169 133 170 134
rect 168 133 169 134
rect 167 133 168 134
rect 166 133 167 134
rect 148 133 149 134
rect 147 133 148 134
rect 146 133 147 134
rect 145 133 146 134
rect 144 133 145 134
rect 143 133 144 134
rect 142 133 143 134
rect 141 133 142 134
rect 140 133 141 134
rect 139 133 140 134
rect 138 133 139 134
rect 137 133 138 134
rect 136 133 137 134
rect 135 133 136 134
rect 134 133 135 134
rect 133 133 134 134
rect 132 133 133 134
rect 131 133 132 134
rect 130 133 131 134
rect 129 133 130 134
rect 128 133 129 134
rect 127 133 128 134
rect 126 133 127 134
rect 125 133 126 134
rect 124 133 125 134
rect 123 133 124 134
rect 122 133 123 134
rect 121 133 122 134
rect 120 133 121 134
rect 119 133 120 134
rect 118 133 119 134
rect 117 133 118 134
rect 116 133 117 134
rect 115 133 116 134
rect 114 133 115 134
rect 113 133 114 134
rect 112 133 113 134
rect 111 133 112 134
rect 110 133 111 134
rect 109 133 110 134
rect 108 133 109 134
rect 107 133 108 134
rect 106 133 107 134
rect 105 133 106 134
rect 104 133 105 134
rect 103 133 104 134
rect 102 133 103 134
rect 101 133 102 134
rect 100 133 101 134
rect 99 133 100 134
rect 98 133 99 134
rect 97 133 98 134
rect 96 133 97 134
rect 95 133 96 134
rect 94 133 95 134
rect 93 133 94 134
rect 92 133 93 134
rect 91 133 92 134
rect 90 133 91 134
rect 89 133 90 134
rect 88 133 89 134
rect 87 133 88 134
rect 86 133 87 134
rect 85 133 86 134
rect 84 133 85 134
rect 83 133 84 134
rect 82 133 83 134
rect 81 133 82 134
rect 80 133 81 134
rect 79 133 80 134
rect 78 133 79 134
rect 77 133 78 134
rect 76 133 77 134
rect 75 133 76 134
rect 74 133 75 134
rect 73 133 74 134
rect 72 133 73 134
rect 71 133 72 134
rect 70 133 71 134
rect 69 133 70 134
rect 68 133 69 134
rect 67 133 68 134
rect 66 133 67 134
rect 65 133 66 134
rect 64 133 65 134
rect 60 133 61 134
rect 59 133 60 134
rect 58 133 59 134
rect 57 133 58 134
rect 56 133 57 134
rect 55 133 56 134
rect 54 133 55 134
rect 53 133 54 134
rect 52 133 53 134
rect 51 133 52 134
rect 50 133 51 134
rect 49 133 50 134
rect 48 133 49 134
rect 47 133 48 134
rect 46 133 47 134
rect 45 133 46 134
rect 44 133 45 134
rect 43 133 44 134
rect 42 133 43 134
rect 41 133 42 134
rect 40 133 41 134
rect 39 133 40 134
rect 38 133 39 134
rect 37 133 38 134
rect 36 133 37 134
rect 35 133 36 134
rect 34 133 35 134
rect 33 133 34 134
rect 463 134 464 135
rect 462 134 463 135
rect 442 134 443 135
rect 441 134 442 135
rect 440 134 441 135
rect 439 134 440 135
rect 438 134 439 135
rect 437 134 438 135
rect 398 134 399 135
rect 397 134 398 135
rect 308 134 309 135
rect 307 134 308 135
rect 306 134 307 135
rect 305 134 306 135
rect 304 134 305 135
rect 303 134 304 135
rect 302 134 303 135
rect 301 134 302 135
rect 300 134 301 135
rect 299 134 300 135
rect 298 134 299 135
rect 297 134 298 135
rect 296 134 297 135
rect 295 134 296 135
rect 294 134 295 135
rect 293 134 294 135
rect 292 134 293 135
rect 291 134 292 135
rect 290 134 291 135
rect 289 134 290 135
rect 288 134 289 135
rect 287 134 288 135
rect 286 134 287 135
rect 285 134 286 135
rect 284 134 285 135
rect 283 134 284 135
rect 282 134 283 135
rect 281 134 282 135
rect 280 134 281 135
rect 279 134 280 135
rect 278 134 279 135
rect 277 134 278 135
rect 276 134 277 135
rect 275 134 276 135
rect 274 134 275 135
rect 273 134 274 135
rect 272 134 273 135
rect 271 134 272 135
rect 270 134 271 135
rect 269 134 270 135
rect 268 134 269 135
rect 267 134 268 135
rect 266 134 267 135
rect 265 134 266 135
rect 264 134 265 135
rect 263 134 264 135
rect 262 134 263 135
rect 261 134 262 135
rect 260 134 261 135
rect 259 134 260 135
rect 229 134 230 135
rect 228 134 229 135
rect 227 134 228 135
rect 226 134 227 135
rect 225 134 226 135
rect 224 134 225 135
rect 223 134 224 135
rect 222 134 223 135
rect 221 134 222 135
rect 220 134 221 135
rect 219 134 220 135
rect 218 134 219 135
rect 217 134 218 135
rect 216 134 217 135
rect 215 134 216 135
rect 214 134 215 135
rect 213 134 214 135
rect 212 134 213 135
rect 211 134 212 135
rect 210 134 211 135
rect 209 134 210 135
rect 208 134 209 135
rect 207 134 208 135
rect 206 134 207 135
rect 205 134 206 135
rect 204 134 205 135
rect 203 134 204 135
rect 202 134 203 135
rect 201 134 202 135
rect 200 134 201 135
rect 199 134 200 135
rect 198 134 199 135
rect 197 134 198 135
rect 196 134 197 135
rect 195 134 196 135
rect 194 134 195 135
rect 193 134 194 135
rect 192 134 193 135
rect 191 134 192 135
rect 190 134 191 135
rect 189 134 190 135
rect 188 134 189 135
rect 187 134 188 135
rect 186 134 187 135
rect 185 134 186 135
rect 184 134 185 135
rect 183 134 184 135
rect 182 134 183 135
rect 181 134 182 135
rect 180 134 181 135
rect 179 134 180 135
rect 178 134 179 135
rect 177 134 178 135
rect 176 134 177 135
rect 175 134 176 135
rect 174 134 175 135
rect 173 134 174 135
rect 172 134 173 135
rect 171 134 172 135
rect 170 134 171 135
rect 169 134 170 135
rect 168 134 169 135
rect 167 134 168 135
rect 166 134 167 135
rect 148 134 149 135
rect 147 134 148 135
rect 146 134 147 135
rect 145 134 146 135
rect 144 134 145 135
rect 143 134 144 135
rect 142 134 143 135
rect 141 134 142 135
rect 140 134 141 135
rect 139 134 140 135
rect 138 134 139 135
rect 137 134 138 135
rect 136 134 137 135
rect 135 134 136 135
rect 134 134 135 135
rect 133 134 134 135
rect 132 134 133 135
rect 131 134 132 135
rect 130 134 131 135
rect 129 134 130 135
rect 128 134 129 135
rect 127 134 128 135
rect 126 134 127 135
rect 125 134 126 135
rect 124 134 125 135
rect 123 134 124 135
rect 122 134 123 135
rect 121 134 122 135
rect 120 134 121 135
rect 119 134 120 135
rect 118 134 119 135
rect 117 134 118 135
rect 116 134 117 135
rect 115 134 116 135
rect 114 134 115 135
rect 113 134 114 135
rect 112 134 113 135
rect 111 134 112 135
rect 110 134 111 135
rect 109 134 110 135
rect 108 134 109 135
rect 107 134 108 135
rect 106 134 107 135
rect 105 134 106 135
rect 104 134 105 135
rect 103 134 104 135
rect 102 134 103 135
rect 101 134 102 135
rect 100 134 101 135
rect 99 134 100 135
rect 98 134 99 135
rect 97 134 98 135
rect 96 134 97 135
rect 95 134 96 135
rect 94 134 95 135
rect 93 134 94 135
rect 92 134 93 135
rect 91 134 92 135
rect 90 134 91 135
rect 89 134 90 135
rect 88 134 89 135
rect 87 134 88 135
rect 86 134 87 135
rect 85 134 86 135
rect 84 134 85 135
rect 83 134 84 135
rect 82 134 83 135
rect 81 134 82 135
rect 80 134 81 135
rect 79 134 80 135
rect 78 134 79 135
rect 77 134 78 135
rect 76 134 77 135
rect 75 134 76 135
rect 74 134 75 135
rect 73 134 74 135
rect 72 134 73 135
rect 71 134 72 135
rect 70 134 71 135
rect 69 134 70 135
rect 68 134 69 135
rect 67 134 68 135
rect 66 134 67 135
rect 65 134 66 135
rect 64 134 65 135
rect 63 134 64 135
rect 60 134 61 135
rect 59 134 60 135
rect 58 134 59 135
rect 57 134 58 135
rect 56 134 57 135
rect 55 134 56 135
rect 54 134 55 135
rect 53 134 54 135
rect 52 134 53 135
rect 51 134 52 135
rect 50 134 51 135
rect 49 134 50 135
rect 48 134 49 135
rect 47 134 48 135
rect 46 134 47 135
rect 45 134 46 135
rect 44 134 45 135
rect 43 134 44 135
rect 42 134 43 135
rect 41 134 42 135
rect 40 134 41 135
rect 39 134 40 135
rect 38 134 39 135
rect 37 134 38 135
rect 36 134 37 135
rect 35 134 36 135
rect 34 134 35 135
rect 33 134 34 135
rect 462 135 463 136
rect 441 135 442 136
rect 440 135 441 136
rect 439 135 440 136
rect 438 135 439 136
rect 437 135 438 136
rect 399 135 400 136
rect 398 135 399 136
rect 397 135 398 136
rect 309 135 310 136
rect 308 135 309 136
rect 307 135 308 136
rect 306 135 307 136
rect 305 135 306 136
rect 304 135 305 136
rect 303 135 304 136
rect 302 135 303 136
rect 301 135 302 136
rect 300 135 301 136
rect 299 135 300 136
rect 298 135 299 136
rect 297 135 298 136
rect 296 135 297 136
rect 295 135 296 136
rect 294 135 295 136
rect 293 135 294 136
rect 292 135 293 136
rect 291 135 292 136
rect 290 135 291 136
rect 289 135 290 136
rect 288 135 289 136
rect 287 135 288 136
rect 286 135 287 136
rect 285 135 286 136
rect 284 135 285 136
rect 283 135 284 136
rect 282 135 283 136
rect 281 135 282 136
rect 280 135 281 136
rect 279 135 280 136
rect 278 135 279 136
rect 277 135 278 136
rect 276 135 277 136
rect 275 135 276 136
rect 274 135 275 136
rect 273 135 274 136
rect 272 135 273 136
rect 271 135 272 136
rect 270 135 271 136
rect 269 135 270 136
rect 268 135 269 136
rect 267 135 268 136
rect 266 135 267 136
rect 265 135 266 136
rect 264 135 265 136
rect 263 135 264 136
rect 262 135 263 136
rect 261 135 262 136
rect 260 135 261 136
rect 259 135 260 136
rect 258 135 259 136
rect 257 135 258 136
rect 229 135 230 136
rect 228 135 229 136
rect 227 135 228 136
rect 226 135 227 136
rect 225 135 226 136
rect 224 135 225 136
rect 223 135 224 136
rect 222 135 223 136
rect 221 135 222 136
rect 220 135 221 136
rect 219 135 220 136
rect 218 135 219 136
rect 217 135 218 136
rect 216 135 217 136
rect 215 135 216 136
rect 214 135 215 136
rect 213 135 214 136
rect 212 135 213 136
rect 211 135 212 136
rect 210 135 211 136
rect 209 135 210 136
rect 208 135 209 136
rect 207 135 208 136
rect 206 135 207 136
rect 205 135 206 136
rect 204 135 205 136
rect 203 135 204 136
rect 202 135 203 136
rect 201 135 202 136
rect 200 135 201 136
rect 199 135 200 136
rect 198 135 199 136
rect 197 135 198 136
rect 196 135 197 136
rect 195 135 196 136
rect 194 135 195 136
rect 193 135 194 136
rect 192 135 193 136
rect 191 135 192 136
rect 190 135 191 136
rect 189 135 190 136
rect 188 135 189 136
rect 187 135 188 136
rect 186 135 187 136
rect 185 135 186 136
rect 184 135 185 136
rect 183 135 184 136
rect 182 135 183 136
rect 181 135 182 136
rect 180 135 181 136
rect 179 135 180 136
rect 178 135 179 136
rect 177 135 178 136
rect 176 135 177 136
rect 175 135 176 136
rect 174 135 175 136
rect 173 135 174 136
rect 172 135 173 136
rect 171 135 172 136
rect 170 135 171 136
rect 169 135 170 136
rect 168 135 169 136
rect 167 135 168 136
rect 166 135 167 136
rect 165 135 166 136
rect 147 135 148 136
rect 146 135 147 136
rect 145 135 146 136
rect 144 135 145 136
rect 143 135 144 136
rect 142 135 143 136
rect 141 135 142 136
rect 140 135 141 136
rect 139 135 140 136
rect 138 135 139 136
rect 137 135 138 136
rect 136 135 137 136
rect 135 135 136 136
rect 134 135 135 136
rect 133 135 134 136
rect 132 135 133 136
rect 131 135 132 136
rect 130 135 131 136
rect 129 135 130 136
rect 128 135 129 136
rect 127 135 128 136
rect 126 135 127 136
rect 125 135 126 136
rect 124 135 125 136
rect 123 135 124 136
rect 122 135 123 136
rect 121 135 122 136
rect 120 135 121 136
rect 119 135 120 136
rect 118 135 119 136
rect 117 135 118 136
rect 116 135 117 136
rect 115 135 116 136
rect 114 135 115 136
rect 113 135 114 136
rect 112 135 113 136
rect 111 135 112 136
rect 110 135 111 136
rect 109 135 110 136
rect 108 135 109 136
rect 107 135 108 136
rect 106 135 107 136
rect 105 135 106 136
rect 104 135 105 136
rect 103 135 104 136
rect 102 135 103 136
rect 101 135 102 136
rect 100 135 101 136
rect 99 135 100 136
rect 98 135 99 136
rect 97 135 98 136
rect 96 135 97 136
rect 95 135 96 136
rect 94 135 95 136
rect 93 135 94 136
rect 92 135 93 136
rect 91 135 92 136
rect 90 135 91 136
rect 89 135 90 136
rect 88 135 89 136
rect 87 135 88 136
rect 86 135 87 136
rect 85 135 86 136
rect 84 135 85 136
rect 83 135 84 136
rect 82 135 83 136
rect 81 135 82 136
rect 80 135 81 136
rect 79 135 80 136
rect 78 135 79 136
rect 77 135 78 136
rect 76 135 77 136
rect 75 135 76 136
rect 74 135 75 136
rect 73 135 74 136
rect 72 135 73 136
rect 71 135 72 136
rect 70 135 71 136
rect 69 135 70 136
rect 68 135 69 136
rect 67 135 68 136
rect 66 135 67 136
rect 65 135 66 136
rect 64 135 65 136
rect 63 135 64 136
rect 60 135 61 136
rect 59 135 60 136
rect 58 135 59 136
rect 57 135 58 136
rect 56 135 57 136
rect 55 135 56 136
rect 54 135 55 136
rect 53 135 54 136
rect 52 135 53 136
rect 51 135 52 136
rect 50 135 51 136
rect 49 135 50 136
rect 48 135 49 136
rect 47 135 48 136
rect 46 135 47 136
rect 45 135 46 136
rect 44 135 45 136
rect 43 135 44 136
rect 42 135 43 136
rect 41 135 42 136
rect 40 135 41 136
rect 39 135 40 136
rect 38 135 39 136
rect 37 135 38 136
rect 36 135 37 136
rect 35 135 36 136
rect 34 135 35 136
rect 462 136 463 137
rect 441 136 442 137
rect 440 136 441 137
rect 439 136 440 137
rect 438 136 439 137
rect 437 136 438 137
rect 436 136 437 137
rect 399 136 400 137
rect 398 136 399 137
rect 397 136 398 137
rect 310 136 311 137
rect 309 136 310 137
rect 308 136 309 137
rect 307 136 308 137
rect 306 136 307 137
rect 305 136 306 137
rect 304 136 305 137
rect 303 136 304 137
rect 302 136 303 137
rect 301 136 302 137
rect 300 136 301 137
rect 299 136 300 137
rect 298 136 299 137
rect 297 136 298 137
rect 296 136 297 137
rect 295 136 296 137
rect 294 136 295 137
rect 293 136 294 137
rect 292 136 293 137
rect 291 136 292 137
rect 290 136 291 137
rect 289 136 290 137
rect 288 136 289 137
rect 287 136 288 137
rect 286 136 287 137
rect 285 136 286 137
rect 284 136 285 137
rect 283 136 284 137
rect 282 136 283 137
rect 281 136 282 137
rect 280 136 281 137
rect 279 136 280 137
rect 278 136 279 137
rect 277 136 278 137
rect 276 136 277 137
rect 275 136 276 137
rect 274 136 275 137
rect 273 136 274 137
rect 272 136 273 137
rect 271 136 272 137
rect 270 136 271 137
rect 269 136 270 137
rect 268 136 269 137
rect 267 136 268 137
rect 266 136 267 137
rect 265 136 266 137
rect 264 136 265 137
rect 263 136 264 137
rect 262 136 263 137
rect 261 136 262 137
rect 260 136 261 137
rect 259 136 260 137
rect 258 136 259 137
rect 257 136 258 137
rect 256 136 257 137
rect 228 136 229 137
rect 227 136 228 137
rect 226 136 227 137
rect 225 136 226 137
rect 224 136 225 137
rect 223 136 224 137
rect 222 136 223 137
rect 221 136 222 137
rect 220 136 221 137
rect 219 136 220 137
rect 218 136 219 137
rect 217 136 218 137
rect 216 136 217 137
rect 215 136 216 137
rect 214 136 215 137
rect 213 136 214 137
rect 212 136 213 137
rect 211 136 212 137
rect 210 136 211 137
rect 209 136 210 137
rect 208 136 209 137
rect 207 136 208 137
rect 206 136 207 137
rect 205 136 206 137
rect 204 136 205 137
rect 203 136 204 137
rect 202 136 203 137
rect 201 136 202 137
rect 200 136 201 137
rect 199 136 200 137
rect 198 136 199 137
rect 197 136 198 137
rect 196 136 197 137
rect 195 136 196 137
rect 194 136 195 137
rect 193 136 194 137
rect 192 136 193 137
rect 191 136 192 137
rect 190 136 191 137
rect 189 136 190 137
rect 188 136 189 137
rect 187 136 188 137
rect 186 136 187 137
rect 185 136 186 137
rect 184 136 185 137
rect 183 136 184 137
rect 182 136 183 137
rect 181 136 182 137
rect 180 136 181 137
rect 179 136 180 137
rect 178 136 179 137
rect 177 136 178 137
rect 176 136 177 137
rect 175 136 176 137
rect 174 136 175 137
rect 173 136 174 137
rect 172 136 173 137
rect 171 136 172 137
rect 170 136 171 137
rect 169 136 170 137
rect 168 136 169 137
rect 167 136 168 137
rect 166 136 167 137
rect 165 136 166 137
rect 147 136 148 137
rect 146 136 147 137
rect 145 136 146 137
rect 144 136 145 137
rect 143 136 144 137
rect 142 136 143 137
rect 141 136 142 137
rect 140 136 141 137
rect 139 136 140 137
rect 138 136 139 137
rect 137 136 138 137
rect 136 136 137 137
rect 135 136 136 137
rect 134 136 135 137
rect 133 136 134 137
rect 132 136 133 137
rect 131 136 132 137
rect 130 136 131 137
rect 129 136 130 137
rect 128 136 129 137
rect 127 136 128 137
rect 126 136 127 137
rect 125 136 126 137
rect 124 136 125 137
rect 123 136 124 137
rect 122 136 123 137
rect 121 136 122 137
rect 120 136 121 137
rect 119 136 120 137
rect 118 136 119 137
rect 117 136 118 137
rect 116 136 117 137
rect 115 136 116 137
rect 114 136 115 137
rect 113 136 114 137
rect 112 136 113 137
rect 111 136 112 137
rect 110 136 111 137
rect 109 136 110 137
rect 108 136 109 137
rect 107 136 108 137
rect 106 136 107 137
rect 105 136 106 137
rect 104 136 105 137
rect 103 136 104 137
rect 102 136 103 137
rect 101 136 102 137
rect 100 136 101 137
rect 99 136 100 137
rect 98 136 99 137
rect 97 136 98 137
rect 96 136 97 137
rect 95 136 96 137
rect 94 136 95 137
rect 93 136 94 137
rect 92 136 93 137
rect 91 136 92 137
rect 90 136 91 137
rect 89 136 90 137
rect 88 136 89 137
rect 87 136 88 137
rect 86 136 87 137
rect 85 136 86 137
rect 84 136 85 137
rect 83 136 84 137
rect 82 136 83 137
rect 81 136 82 137
rect 80 136 81 137
rect 79 136 80 137
rect 78 136 79 137
rect 77 136 78 137
rect 76 136 77 137
rect 75 136 76 137
rect 74 136 75 137
rect 73 136 74 137
rect 72 136 73 137
rect 71 136 72 137
rect 70 136 71 137
rect 69 136 70 137
rect 68 136 69 137
rect 67 136 68 137
rect 66 136 67 137
rect 65 136 66 137
rect 64 136 65 137
rect 63 136 64 137
rect 62 136 63 137
rect 60 136 61 137
rect 59 136 60 137
rect 58 136 59 137
rect 57 136 58 137
rect 56 136 57 137
rect 55 136 56 137
rect 54 136 55 137
rect 53 136 54 137
rect 52 136 53 137
rect 51 136 52 137
rect 50 136 51 137
rect 49 136 50 137
rect 48 136 49 137
rect 47 136 48 137
rect 46 136 47 137
rect 45 136 46 137
rect 44 136 45 137
rect 43 136 44 137
rect 42 136 43 137
rect 41 136 42 137
rect 40 136 41 137
rect 39 136 40 137
rect 38 136 39 137
rect 37 136 38 137
rect 36 136 37 137
rect 35 136 36 137
rect 441 137 442 138
rect 440 137 441 138
rect 439 137 440 138
rect 438 137 439 138
rect 437 137 438 138
rect 436 137 437 138
rect 435 137 436 138
rect 399 137 400 138
rect 398 137 399 138
rect 397 137 398 138
rect 311 137 312 138
rect 310 137 311 138
rect 309 137 310 138
rect 308 137 309 138
rect 307 137 308 138
rect 306 137 307 138
rect 305 137 306 138
rect 304 137 305 138
rect 303 137 304 138
rect 302 137 303 138
rect 301 137 302 138
rect 300 137 301 138
rect 299 137 300 138
rect 298 137 299 138
rect 297 137 298 138
rect 296 137 297 138
rect 295 137 296 138
rect 294 137 295 138
rect 293 137 294 138
rect 292 137 293 138
rect 291 137 292 138
rect 290 137 291 138
rect 289 137 290 138
rect 288 137 289 138
rect 287 137 288 138
rect 286 137 287 138
rect 285 137 286 138
rect 284 137 285 138
rect 283 137 284 138
rect 282 137 283 138
rect 281 137 282 138
rect 280 137 281 138
rect 279 137 280 138
rect 278 137 279 138
rect 277 137 278 138
rect 276 137 277 138
rect 275 137 276 138
rect 274 137 275 138
rect 273 137 274 138
rect 272 137 273 138
rect 271 137 272 138
rect 270 137 271 138
rect 269 137 270 138
rect 268 137 269 138
rect 267 137 268 138
rect 266 137 267 138
rect 265 137 266 138
rect 264 137 265 138
rect 263 137 264 138
rect 262 137 263 138
rect 261 137 262 138
rect 260 137 261 138
rect 259 137 260 138
rect 258 137 259 138
rect 257 137 258 138
rect 256 137 257 138
rect 255 137 256 138
rect 227 137 228 138
rect 226 137 227 138
rect 225 137 226 138
rect 224 137 225 138
rect 223 137 224 138
rect 222 137 223 138
rect 221 137 222 138
rect 220 137 221 138
rect 219 137 220 138
rect 218 137 219 138
rect 217 137 218 138
rect 216 137 217 138
rect 215 137 216 138
rect 214 137 215 138
rect 213 137 214 138
rect 212 137 213 138
rect 211 137 212 138
rect 210 137 211 138
rect 209 137 210 138
rect 208 137 209 138
rect 207 137 208 138
rect 206 137 207 138
rect 205 137 206 138
rect 204 137 205 138
rect 203 137 204 138
rect 202 137 203 138
rect 201 137 202 138
rect 200 137 201 138
rect 199 137 200 138
rect 198 137 199 138
rect 197 137 198 138
rect 196 137 197 138
rect 195 137 196 138
rect 194 137 195 138
rect 193 137 194 138
rect 192 137 193 138
rect 191 137 192 138
rect 190 137 191 138
rect 189 137 190 138
rect 188 137 189 138
rect 187 137 188 138
rect 186 137 187 138
rect 185 137 186 138
rect 184 137 185 138
rect 183 137 184 138
rect 182 137 183 138
rect 181 137 182 138
rect 180 137 181 138
rect 179 137 180 138
rect 178 137 179 138
rect 177 137 178 138
rect 176 137 177 138
rect 175 137 176 138
rect 174 137 175 138
rect 173 137 174 138
rect 172 137 173 138
rect 171 137 172 138
rect 170 137 171 138
rect 169 137 170 138
rect 168 137 169 138
rect 167 137 168 138
rect 166 137 167 138
rect 165 137 166 138
rect 164 137 165 138
rect 146 137 147 138
rect 145 137 146 138
rect 144 137 145 138
rect 143 137 144 138
rect 142 137 143 138
rect 141 137 142 138
rect 140 137 141 138
rect 139 137 140 138
rect 138 137 139 138
rect 137 137 138 138
rect 136 137 137 138
rect 135 137 136 138
rect 134 137 135 138
rect 133 137 134 138
rect 132 137 133 138
rect 131 137 132 138
rect 130 137 131 138
rect 129 137 130 138
rect 128 137 129 138
rect 127 137 128 138
rect 126 137 127 138
rect 125 137 126 138
rect 124 137 125 138
rect 123 137 124 138
rect 122 137 123 138
rect 121 137 122 138
rect 120 137 121 138
rect 119 137 120 138
rect 118 137 119 138
rect 117 137 118 138
rect 116 137 117 138
rect 115 137 116 138
rect 114 137 115 138
rect 113 137 114 138
rect 112 137 113 138
rect 111 137 112 138
rect 110 137 111 138
rect 109 137 110 138
rect 108 137 109 138
rect 107 137 108 138
rect 106 137 107 138
rect 105 137 106 138
rect 104 137 105 138
rect 103 137 104 138
rect 102 137 103 138
rect 101 137 102 138
rect 100 137 101 138
rect 99 137 100 138
rect 98 137 99 138
rect 97 137 98 138
rect 96 137 97 138
rect 95 137 96 138
rect 94 137 95 138
rect 93 137 94 138
rect 92 137 93 138
rect 91 137 92 138
rect 90 137 91 138
rect 89 137 90 138
rect 88 137 89 138
rect 87 137 88 138
rect 86 137 87 138
rect 85 137 86 138
rect 84 137 85 138
rect 83 137 84 138
rect 82 137 83 138
rect 81 137 82 138
rect 80 137 81 138
rect 79 137 80 138
rect 78 137 79 138
rect 77 137 78 138
rect 76 137 77 138
rect 75 137 76 138
rect 74 137 75 138
rect 73 137 74 138
rect 72 137 73 138
rect 71 137 72 138
rect 70 137 71 138
rect 69 137 70 138
rect 68 137 69 138
rect 67 137 68 138
rect 66 137 67 138
rect 65 137 66 138
rect 64 137 65 138
rect 63 137 64 138
rect 62 137 63 138
rect 61 137 62 138
rect 60 137 61 138
rect 59 137 60 138
rect 58 137 59 138
rect 57 137 58 138
rect 56 137 57 138
rect 55 137 56 138
rect 54 137 55 138
rect 53 137 54 138
rect 52 137 53 138
rect 51 137 52 138
rect 50 137 51 138
rect 49 137 50 138
rect 48 137 49 138
rect 47 137 48 138
rect 46 137 47 138
rect 45 137 46 138
rect 44 137 45 138
rect 43 137 44 138
rect 42 137 43 138
rect 41 137 42 138
rect 40 137 41 138
rect 39 137 40 138
rect 38 137 39 138
rect 37 137 38 138
rect 36 137 37 138
rect 35 137 36 138
rect 440 138 441 139
rect 439 138 440 139
rect 438 138 439 139
rect 437 138 438 139
rect 436 138 437 139
rect 435 138 436 139
rect 434 138 435 139
rect 400 138 401 139
rect 399 138 400 139
rect 398 138 399 139
rect 397 138 398 139
rect 312 138 313 139
rect 311 138 312 139
rect 310 138 311 139
rect 309 138 310 139
rect 308 138 309 139
rect 307 138 308 139
rect 306 138 307 139
rect 305 138 306 139
rect 304 138 305 139
rect 303 138 304 139
rect 302 138 303 139
rect 301 138 302 139
rect 300 138 301 139
rect 299 138 300 139
rect 298 138 299 139
rect 297 138 298 139
rect 296 138 297 139
rect 295 138 296 139
rect 294 138 295 139
rect 293 138 294 139
rect 292 138 293 139
rect 291 138 292 139
rect 290 138 291 139
rect 289 138 290 139
rect 288 138 289 139
rect 287 138 288 139
rect 286 138 287 139
rect 285 138 286 139
rect 284 138 285 139
rect 283 138 284 139
rect 282 138 283 139
rect 281 138 282 139
rect 280 138 281 139
rect 279 138 280 139
rect 278 138 279 139
rect 277 138 278 139
rect 276 138 277 139
rect 275 138 276 139
rect 274 138 275 139
rect 273 138 274 139
rect 272 138 273 139
rect 271 138 272 139
rect 270 138 271 139
rect 269 138 270 139
rect 268 138 269 139
rect 267 138 268 139
rect 266 138 267 139
rect 265 138 266 139
rect 264 138 265 139
rect 263 138 264 139
rect 262 138 263 139
rect 261 138 262 139
rect 260 138 261 139
rect 259 138 260 139
rect 258 138 259 139
rect 257 138 258 139
rect 256 138 257 139
rect 255 138 256 139
rect 254 138 255 139
rect 253 138 254 139
rect 227 138 228 139
rect 226 138 227 139
rect 225 138 226 139
rect 224 138 225 139
rect 223 138 224 139
rect 222 138 223 139
rect 221 138 222 139
rect 220 138 221 139
rect 219 138 220 139
rect 218 138 219 139
rect 217 138 218 139
rect 216 138 217 139
rect 215 138 216 139
rect 214 138 215 139
rect 213 138 214 139
rect 212 138 213 139
rect 211 138 212 139
rect 210 138 211 139
rect 209 138 210 139
rect 208 138 209 139
rect 207 138 208 139
rect 206 138 207 139
rect 205 138 206 139
rect 204 138 205 139
rect 203 138 204 139
rect 202 138 203 139
rect 201 138 202 139
rect 200 138 201 139
rect 199 138 200 139
rect 198 138 199 139
rect 197 138 198 139
rect 196 138 197 139
rect 195 138 196 139
rect 194 138 195 139
rect 193 138 194 139
rect 192 138 193 139
rect 191 138 192 139
rect 190 138 191 139
rect 189 138 190 139
rect 188 138 189 139
rect 187 138 188 139
rect 186 138 187 139
rect 185 138 186 139
rect 184 138 185 139
rect 183 138 184 139
rect 182 138 183 139
rect 181 138 182 139
rect 180 138 181 139
rect 179 138 180 139
rect 178 138 179 139
rect 177 138 178 139
rect 176 138 177 139
rect 175 138 176 139
rect 174 138 175 139
rect 173 138 174 139
rect 172 138 173 139
rect 171 138 172 139
rect 170 138 171 139
rect 169 138 170 139
rect 168 138 169 139
rect 167 138 168 139
rect 166 138 167 139
rect 165 138 166 139
rect 164 138 165 139
rect 145 138 146 139
rect 144 138 145 139
rect 143 138 144 139
rect 142 138 143 139
rect 141 138 142 139
rect 140 138 141 139
rect 139 138 140 139
rect 138 138 139 139
rect 137 138 138 139
rect 136 138 137 139
rect 135 138 136 139
rect 134 138 135 139
rect 133 138 134 139
rect 132 138 133 139
rect 131 138 132 139
rect 130 138 131 139
rect 129 138 130 139
rect 128 138 129 139
rect 127 138 128 139
rect 126 138 127 139
rect 125 138 126 139
rect 124 138 125 139
rect 123 138 124 139
rect 122 138 123 139
rect 121 138 122 139
rect 120 138 121 139
rect 119 138 120 139
rect 118 138 119 139
rect 117 138 118 139
rect 116 138 117 139
rect 115 138 116 139
rect 114 138 115 139
rect 113 138 114 139
rect 112 138 113 139
rect 111 138 112 139
rect 110 138 111 139
rect 109 138 110 139
rect 108 138 109 139
rect 107 138 108 139
rect 106 138 107 139
rect 105 138 106 139
rect 104 138 105 139
rect 103 138 104 139
rect 102 138 103 139
rect 101 138 102 139
rect 100 138 101 139
rect 99 138 100 139
rect 98 138 99 139
rect 97 138 98 139
rect 96 138 97 139
rect 95 138 96 139
rect 94 138 95 139
rect 93 138 94 139
rect 92 138 93 139
rect 91 138 92 139
rect 90 138 91 139
rect 89 138 90 139
rect 88 138 89 139
rect 87 138 88 139
rect 86 138 87 139
rect 85 138 86 139
rect 84 138 85 139
rect 83 138 84 139
rect 82 138 83 139
rect 81 138 82 139
rect 80 138 81 139
rect 79 138 80 139
rect 78 138 79 139
rect 77 138 78 139
rect 76 138 77 139
rect 75 138 76 139
rect 74 138 75 139
rect 73 138 74 139
rect 72 138 73 139
rect 71 138 72 139
rect 70 138 71 139
rect 69 138 70 139
rect 68 138 69 139
rect 67 138 68 139
rect 66 138 67 139
rect 65 138 66 139
rect 64 138 65 139
rect 63 138 64 139
rect 62 138 63 139
rect 61 138 62 139
rect 60 138 61 139
rect 59 138 60 139
rect 58 138 59 139
rect 57 138 58 139
rect 56 138 57 139
rect 55 138 56 139
rect 54 138 55 139
rect 53 138 54 139
rect 52 138 53 139
rect 51 138 52 139
rect 50 138 51 139
rect 49 138 50 139
rect 48 138 49 139
rect 47 138 48 139
rect 46 138 47 139
rect 45 138 46 139
rect 44 138 45 139
rect 43 138 44 139
rect 42 138 43 139
rect 41 138 42 139
rect 40 138 41 139
rect 39 138 40 139
rect 38 138 39 139
rect 37 138 38 139
rect 36 138 37 139
rect 440 139 441 140
rect 439 139 440 140
rect 438 139 439 140
rect 437 139 438 140
rect 436 139 437 140
rect 435 139 436 140
rect 434 139 435 140
rect 433 139 434 140
rect 432 139 433 140
rect 431 139 432 140
rect 401 139 402 140
rect 400 139 401 140
rect 399 139 400 140
rect 398 139 399 140
rect 397 139 398 140
rect 312 139 313 140
rect 311 139 312 140
rect 310 139 311 140
rect 309 139 310 140
rect 308 139 309 140
rect 307 139 308 140
rect 306 139 307 140
rect 305 139 306 140
rect 304 139 305 140
rect 303 139 304 140
rect 302 139 303 140
rect 301 139 302 140
rect 300 139 301 140
rect 299 139 300 140
rect 298 139 299 140
rect 297 139 298 140
rect 296 139 297 140
rect 295 139 296 140
rect 294 139 295 140
rect 293 139 294 140
rect 292 139 293 140
rect 291 139 292 140
rect 290 139 291 140
rect 289 139 290 140
rect 288 139 289 140
rect 287 139 288 140
rect 286 139 287 140
rect 285 139 286 140
rect 284 139 285 140
rect 283 139 284 140
rect 282 139 283 140
rect 281 139 282 140
rect 280 139 281 140
rect 279 139 280 140
rect 278 139 279 140
rect 277 139 278 140
rect 276 139 277 140
rect 275 139 276 140
rect 274 139 275 140
rect 273 139 274 140
rect 272 139 273 140
rect 271 139 272 140
rect 270 139 271 140
rect 269 139 270 140
rect 268 139 269 140
rect 267 139 268 140
rect 266 139 267 140
rect 265 139 266 140
rect 264 139 265 140
rect 263 139 264 140
rect 262 139 263 140
rect 261 139 262 140
rect 260 139 261 140
rect 259 139 260 140
rect 258 139 259 140
rect 257 139 258 140
rect 256 139 257 140
rect 255 139 256 140
rect 254 139 255 140
rect 253 139 254 140
rect 252 139 253 140
rect 226 139 227 140
rect 225 139 226 140
rect 224 139 225 140
rect 223 139 224 140
rect 222 139 223 140
rect 221 139 222 140
rect 220 139 221 140
rect 219 139 220 140
rect 218 139 219 140
rect 217 139 218 140
rect 216 139 217 140
rect 215 139 216 140
rect 214 139 215 140
rect 213 139 214 140
rect 212 139 213 140
rect 211 139 212 140
rect 210 139 211 140
rect 209 139 210 140
rect 208 139 209 140
rect 207 139 208 140
rect 206 139 207 140
rect 205 139 206 140
rect 204 139 205 140
rect 203 139 204 140
rect 202 139 203 140
rect 201 139 202 140
rect 200 139 201 140
rect 199 139 200 140
rect 198 139 199 140
rect 197 139 198 140
rect 196 139 197 140
rect 195 139 196 140
rect 194 139 195 140
rect 193 139 194 140
rect 192 139 193 140
rect 191 139 192 140
rect 190 139 191 140
rect 189 139 190 140
rect 188 139 189 140
rect 187 139 188 140
rect 186 139 187 140
rect 185 139 186 140
rect 184 139 185 140
rect 183 139 184 140
rect 182 139 183 140
rect 181 139 182 140
rect 180 139 181 140
rect 179 139 180 140
rect 178 139 179 140
rect 177 139 178 140
rect 176 139 177 140
rect 175 139 176 140
rect 174 139 175 140
rect 173 139 174 140
rect 172 139 173 140
rect 171 139 172 140
rect 170 139 171 140
rect 169 139 170 140
rect 168 139 169 140
rect 167 139 168 140
rect 166 139 167 140
rect 165 139 166 140
rect 164 139 165 140
rect 163 139 164 140
rect 145 139 146 140
rect 144 139 145 140
rect 143 139 144 140
rect 142 139 143 140
rect 141 139 142 140
rect 140 139 141 140
rect 139 139 140 140
rect 138 139 139 140
rect 137 139 138 140
rect 136 139 137 140
rect 135 139 136 140
rect 134 139 135 140
rect 133 139 134 140
rect 132 139 133 140
rect 131 139 132 140
rect 130 139 131 140
rect 129 139 130 140
rect 128 139 129 140
rect 127 139 128 140
rect 126 139 127 140
rect 125 139 126 140
rect 124 139 125 140
rect 123 139 124 140
rect 122 139 123 140
rect 121 139 122 140
rect 120 139 121 140
rect 119 139 120 140
rect 118 139 119 140
rect 117 139 118 140
rect 116 139 117 140
rect 115 139 116 140
rect 114 139 115 140
rect 113 139 114 140
rect 112 139 113 140
rect 111 139 112 140
rect 110 139 111 140
rect 109 139 110 140
rect 108 139 109 140
rect 107 139 108 140
rect 106 139 107 140
rect 105 139 106 140
rect 104 139 105 140
rect 103 139 104 140
rect 102 139 103 140
rect 101 139 102 140
rect 100 139 101 140
rect 99 139 100 140
rect 98 139 99 140
rect 97 139 98 140
rect 96 139 97 140
rect 95 139 96 140
rect 94 139 95 140
rect 93 139 94 140
rect 92 139 93 140
rect 91 139 92 140
rect 90 139 91 140
rect 89 139 90 140
rect 88 139 89 140
rect 87 139 88 140
rect 86 139 87 140
rect 85 139 86 140
rect 84 139 85 140
rect 83 139 84 140
rect 82 139 83 140
rect 81 139 82 140
rect 80 139 81 140
rect 79 139 80 140
rect 78 139 79 140
rect 77 139 78 140
rect 76 139 77 140
rect 75 139 76 140
rect 74 139 75 140
rect 73 139 74 140
rect 72 139 73 140
rect 71 139 72 140
rect 70 139 71 140
rect 69 139 70 140
rect 68 139 69 140
rect 67 139 68 140
rect 66 139 67 140
rect 65 139 66 140
rect 64 139 65 140
rect 63 139 64 140
rect 62 139 63 140
rect 61 139 62 140
rect 60 139 61 140
rect 59 139 60 140
rect 58 139 59 140
rect 57 139 58 140
rect 56 139 57 140
rect 55 139 56 140
rect 54 139 55 140
rect 53 139 54 140
rect 52 139 53 140
rect 51 139 52 140
rect 50 139 51 140
rect 49 139 50 140
rect 48 139 49 140
rect 47 139 48 140
rect 46 139 47 140
rect 45 139 46 140
rect 44 139 45 140
rect 43 139 44 140
rect 42 139 43 140
rect 41 139 42 140
rect 40 139 41 140
rect 39 139 40 140
rect 38 139 39 140
rect 37 139 38 140
rect 439 140 440 141
rect 438 140 439 141
rect 437 140 438 141
rect 436 140 437 141
rect 435 140 436 141
rect 434 140 435 141
rect 433 140 434 141
rect 432 140 433 141
rect 431 140 432 141
rect 430 140 431 141
rect 429 140 430 141
rect 428 140 429 141
rect 427 140 428 141
rect 426 140 427 141
rect 407 140 408 141
rect 406 140 407 141
rect 405 140 406 141
rect 404 140 405 141
rect 403 140 404 141
rect 402 140 403 141
rect 401 140 402 141
rect 400 140 401 141
rect 399 140 400 141
rect 398 140 399 141
rect 397 140 398 141
rect 313 140 314 141
rect 312 140 313 141
rect 311 140 312 141
rect 310 140 311 141
rect 309 140 310 141
rect 308 140 309 141
rect 307 140 308 141
rect 306 140 307 141
rect 305 140 306 141
rect 304 140 305 141
rect 303 140 304 141
rect 302 140 303 141
rect 301 140 302 141
rect 300 140 301 141
rect 299 140 300 141
rect 298 140 299 141
rect 297 140 298 141
rect 296 140 297 141
rect 295 140 296 141
rect 294 140 295 141
rect 293 140 294 141
rect 292 140 293 141
rect 291 140 292 141
rect 290 140 291 141
rect 289 140 290 141
rect 288 140 289 141
rect 287 140 288 141
rect 286 140 287 141
rect 285 140 286 141
rect 284 140 285 141
rect 283 140 284 141
rect 282 140 283 141
rect 281 140 282 141
rect 280 140 281 141
rect 279 140 280 141
rect 278 140 279 141
rect 277 140 278 141
rect 276 140 277 141
rect 275 140 276 141
rect 274 140 275 141
rect 273 140 274 141
rect 272 140 273 141
rect 271 140 272 141
rect 270 140 271 141
rect 269 140 270 141
rect 268 140 269 141
rect 267 140 268 141
rect 266 140 267 141
rect 265 140 266 141
rect 264 140 265 141
rect 263 140 264 141
rect 262 140 263 141
rect 261 140 262 141
rect 260 140 261 141
rect 259 140 260 141
rect 258 140 259 141
rect 257 140 258 141
rect 256 140 257 141
rect 255 140 256 141
rect 254 140 255 141
rect 253 140 254 141
rect 252 140 253 141
rect 251 140 252 141
rect 226 140 227 141
rect 225 140 226 141
rect 224 140 225 141
rect 223 140 224 141
rect 222 140 223 141
rect 221 140 222 141
rect 220 140 221 141
rect 219 140 220 141
rect 218 140 219 141
rect 217 140 218 141
rect 216 140 217 141
rect 215 140 216 141
rect 214 140 215 141
rect 213 140 214 141
rect 212 140 213 141
rect 211 140 212 141
rect 210 140 211 141
rect 209 140 210 141
rect 208 140 209 141
rect 207 140 208 141
rect 206 140 207 141
rect 205 140 206 141
rect 204 140 205 141
rect 203 140 204 141
rect 202 140 203 141
rect 201 140 202 141
rect 200 140 201 141
rect 199 140 200 141
rect 198 140 199 141
rect 197 140 198 141
rect 196 140 197 141
rect 195 140 196 141
rect 194 140 195 141
rect 193 140 194 141
rect 192 140 193 141
rect 191 140 192 141
rect 190 140 191 141
rect 189 140 190 141
rect 188 140 189 141
rect 187 140 188 141
rect 186 140 187 141
rect 185 140 186 141
rect 184 140 185 141
rect 183 140 184 141
rect 182 140 183 141
rect 181 140 182 141
rect 180 140 181 141
rect 179 140 180 141
rect 178 140 179 141
rect 177 140 178 141
rect 176 140 177 141
rect 175 140 176 141
rect 174 140 175 141
rect 173 140 174 141
rect 172 140 173 141
rect 171 140 172 141
rect 170 140 171 141
rect 169 140 170 141
rect 168 140 169 141
rect 167 140 168 141
rect 166 140 167 141
rect 165 140 166 141
rect 164 140 165 141
rect 163 140 164 141
rect 144 140 145 141
rect 143 140 144 141
rect 142 140 143 141
rect 141 140 142 141
rect 140 140 141 141
rect 139 140 140 141
rect 138 140 139 141
rect 137 140 138 141
rect 136 140 137 141
rect 135 140 136 141
rect 134 140 135 141
rect 133 140 134 141
rect 132 140 133 141
rect 131 140 132 141
rect 130 140 131 141
rect 129 140 130 141
rect 128 140 129 141
rect 127 140 128 141
rect 126 140 127 141
rect 125 140 126 141
rect 124 140 125 141
rect 123 140 124 141
rect 122 140 123 141
rect 121 140 122 141
rect 120 140 121 141
rect 119 140 120 141
rect 118 140 119 141
rect 117 140 118 141
rect 116 140 117 141
rect 115 140 116 141
rect 114 140 115 141
rect 113 140 114 141
rect 112 140 113 141
rect 111 140 112 141
rect 110 140 111 141
rect 109 140 110 141
rect 108 140 109 141
rect 107 140 108 141
rect 106 140 107 141
rect 105 140 106 141
rect 104 140 105 141
rect 103 140 104 141
rect 102 140 103 141
rect 101 140 102 141
rect 100 140 101 141
rect 99 140 100 141
rect 98 140 99 141
rect 97 140 98 141
rect 96 140 97 141
rect 95 140 96 141
rect 94 140 95 141
rect 93 140 94 141
rect 92 140 93 141
rect 91 140 92 141
rect 90 140 91 141
rect 89 140 90 141
rect 88 140 89 141
rect 87 140 88 141
rect 86 140 87 141
rect 85 140 86 141
rect 84 140 85 141
rect 83 140 84 141
rect 82 140 83 141
rect 81 140 82 141
rect 80 140 81 141
rect 79 140 80 141
rect 78 140 79 141
rect 77 140 78 141
rect 76 140 77 141
rect 75 140 76 141
rect 74 140 75 141
rect 73 140 74 141
rect 72 140 73 141
rect 71 140 72 141
rect 70 140 71 141
rect 69 140 70 141
rect 68 140 69 141
rect 67 140 68 141
rect 66 140 67 141
rect 65 140 66 141
rect 64 140 65 141
rect 63 140 64 141
rect 62 140 63 141
rect 61 140 62 141
rect 60 140 61 141
rect 59 140 60 141
rect 58 140 59 141
rect 57 140 58 141
rect 56 140 57 141
rect 55 140 56 141
rect 54 140 55 141
rect 53 140 54 141
rect 52 140 53 141
rect 51 140 52 141
rect 50 140 51 141
rect 49 140 50 141
rect 48 140 49 141
rect 47 140 48 141
rect 46 140 47 141
rect 45 140 46 141
rect 44 140 45 141
rect 43 140 44 141
rect 42 140 43 141
rect 41 140 42 141
rect 40 140 41 141
rect 39 140 40 141
rect 38 140 39 141
rect 438 141 439 142
rect 437 141 438 142
rect 436 141 437 142
rect 435 141 436 142
rect 434 141 435 142
rect 433 141 434 142
rect 432 141 433 142
rect 431 141 432 142
rect 430 141 431 142
rect 429 141 430 142
rect 428 141 429 142
rect 427 141 428 142
rect 426 141 427 142
rect 425 141 426 142
rect 424 141 425 142
rect 423 141 424 142
rect 422 141 423 142
rect 421 141 422 142
rect 420 141 421 142
rect 419 141 420 142
rect 418 141 419 142
rect 417 141 418 142
rect 416 141 417 142
rect 415 141 416 142
rect 414 141 415 142
rect 413 141 414 142
rect 412 141 413 142
rect 411 141 412 142
rect 410 141 411 142
rect 409 141 410 142
rect 408 141 409 142
rect 407 141 408 142
rect 406 141 407 142
rect 405 141 406 142
rect 404 141 405 142
rect 403 141 404 142
rect 402 141 403 142
rect 401 141 402 142
rect 400 141 401 142
rect 399 141 400 142
rect 398 141 399 142
rect 397 141 398 142
rect 314 141 315 142
rect 313 141 314 142
rect 312 141 313 142
rect 311 141 312 142
rect 310 141 311 142
rect 309 141 310 142
rect 308 141 309 142
rect 307 141 308 142
rect 306 141 307 142
rect 305 141 306 142
rect 304 141 305 142
rect 303 141 304 142
rect 302 141 303 142
rect 301 141 302 142
rect 300 141 301 142
rect 299 141 300 142
rect 298 141 299 142
rect 297 141 298 142
rect 296 141 297 142
rect 295 141 296 142
rect 294 141 295 142
rect 293 141 294 142
rect 292 141 293 142
rect 291 141 292 142
rect 290 141 291 142
rect 289 141 290 142
rect 288 141 289 142
rect 287 141 288 142
rect 286 141 287 142
rect 285 141 286 142
rect 284 141 285 142
rect 283 141 284 142
rect 282 141 283 142
rect 281 141 282 142
rect 280 141 281 142
rect 279 141 280 142
rect 278 141 279 142
rect 277 141 278 142
rect 276 141 277 142
rect 275 141 276 142
rect 274 141 275 142
rect 273 141 274 142
rect 272 141 273 142
rect 271 141 272 142
rect 270 141 271 142
rect 269 141 270 142
rect 268 141 269 142
rect 267 141 268 142
rect 266 141 267 142
rect 265 141 266 142
rect 264 141 265 142
rect 263 141 264 142
rect 262 141 263 142
rect 261 141 262 142
rect 260 141 261 142
rect 259 141 260 142
rect 258 141 259 142
rect 257 141 258 142
rect 256 141 257 142
rect 255 141 256 142
rect 254 141 255 142
rect 253 141 254 142
rect 252 141 253 142
rect 251 141 252 142
rect 250 141 251 142
rect 225 141 226 142
rect 224 141 225 142
rect 223 141 224 142
rect 222 141 223 142
rect 221 141 222 142
rect 220 141 221 142
rect 219 141 220 142
rect 218 141 219 142
rect 217 141 218 142
rect 216 141 217 142
rect 215 141 216 142
rect 214 141 215 142
rect 213 141 214 142
rect 212 141 213 142
rect 211 141 212 142
rect 210 141 211 142
rect 209 141 210 142
rect 208 141 209 142
rect 207 141 208 142
rect 206 141 207 142
rect 205 141 206 142
rect 204 141 205 142
rect 203 141 204 142
rect 202 141 203 142
rect 201 141 202 142
rect 200 141 201 142
rect 199 141 200 142
rect 198 141 199 142
rect 197 141 198 142
rect 196 141 197 142
rect 195 141 196 142
rect 194 141 195 142
rect 193 141 194 142
rect 192 141 193 142
rect 191 141 192 142
rect 190 141 191 142
rect 189 141 190 142
rect 188 141 189 142
rect 187 141 188 142
rect 186 141 187 142
rect 185 141 186 142
rect 184 141 185 142
rect 183 141 184 142
rect 182 141 183 142
rect 181 141 182 142
rect 180 141 181 142
rect 179 141 180 142
rect 178 141 179 142
rect 177 141 178 142
rect 176 141 177 142
rect 175 141 176 142
rect 174 141 175 142
rect 173 141 174 142
rect 172 141 173 142
rect 171 141 172 142
rect 170 141 171 142
rect 169 141 170 142
rect 168 141 169 142
rect 167 141 168 142
rect 166 141 167 142
rect 165 141 166 142
rect 164 141 165 142
rect 163 141 164 142
rect 162 141 163 142
rect 143 141 144 142
rect 142 141 143 142
rect 141 141 142 142
rect 140 141 141 142
rect 139 141 140 142
rect 138 141 139 142
rect 137 141 138 142
rect 136 141 137 142
rect 135 141 136 142
rect 134 141 135 142
rect 133 141 134 142
rect 132 141 133 142
rect 131 141 132 142
rect 130 141 131 142
rect 129 141 130 142
rect 128 141 129 142
rect 127 141 128 142
rect 126 141 127 142
rect 125 141 126 142
rect 124 141 125 142
rect 123 141 124 142
rect 122 141 123 142
rect 121 141 122 142
rect 120 141 121 142
rect 119 141 120 142
rect 118 141 119 142
rect 117 141 118 142
rect 116 141 117 142
rect 115 141 116 142
rect 114 141 115 142
rect 113 141 114 142
rect 112 141 113 142
rect 111 141 112 142
rect 110 141 111 142
rect 109 141 110 142
rect 108 141 109 142
rect 107 141 108 142
rect 106 141 107 142
rect 105 141 106 142
rect 104 141 105 142
rect 103 141 104 142
rect 102 141 103 142
rect 101 141 102 142
rect 100 141 101 142
rect 99 141 100 142
rect 98 141 99 142
rect 97 141 98 142
rect 96 141 97 142
rect 95 141 96 142
rect 94 141 95 142
rect 93 141 94 142
rect 92 141 93 142
rect 91 141 92 142
rect 90 141 91 142
rect 89 141 90 142
rect 88 141 89 142
rect 87 141 88 142
rect 86 141 87 142
rect 85 141 86 142
rect 84 141 85 142
rect 83 141 84 142
rect 82 141 83 142
rect 81 141 82 142
rect 80 141 81 142
rect 79 141 80 142
rect 78 141 79 142
rect 77 141 78 142
rect 76 141 77 142
rect 75 141 76 142
rect 74 141 75 142
rect 73 141 74 142
rect 72 141 73 142
rect 71 141 72 142
rect 70 141 71 142
rect 69 141 70 142
rect 68 141 69 142
rect 67 141 68 142
rect 66 141 67 142
rect 65 141 66 142
rect 64 141 65 142
rect 63 141 64 142
rect 62 141 63 142
rect 61 141 62 142
rect 60 141 61 142
rect 59 141 60 142
rect 58 141 59 142
rect 57 141 58 142
rect 56 141 57 142
rect 55 141 56 142
rect 54 141 55 142
rect 53 141 54 142
rect 52 141 53 142
rect 51 141 52 142
rect 50 141 51 142
rect 49 141 50 142
rect 48 141 49 142
rect 47 141 48 142
rect 46 141 47 142
rect 45 141 46 142
rect 44 141 45 142
rect 43 141 44 142
rect 42 141 43 142
rect 41 141 42 142
rect 40 141 41 142
rect 39 141 40 142
rect 437 142 438 143
rect 436 142 437 143
rect 435 142 436 143
rect 434 142 435 143
rect 433 142 434 143
rect 432 142 433 143
rect 431 142 432 143
rect 430 142 431 143
rect 429 142 430 143
rect 428 142 429 143
rect 427 142 428 143
rect 426 142 427 143
rect 425 142 426 143
rect 424 142 425 143
rect 423 142 424 143
rect 422 142 423 143
rect 421 142 422 143
rect 420 142 421 143
rect 419 142 420 143
rect 418 142 419 143
rect 417 142 418 143
rect 416 142 417 143
rect 415 142 416 143
rect 414 142 415 143
rect 413 142 414 143
rect 412 142 413 143
rect 411 142 412 143
rect 410 142 411 143
rect 409 142 410 143
rect 408 142 409 143
rect 407 142 408 143
rect 406 142 407 143
rect 405 142 406 143
rect 404 142 405 143
rect 403 142 404 143
rect 402 142 403 143
rect 401 142 402 143
rect 400 142 401 143
rect 399 142 400 143
rect 398 142 399 143
rect 397 142 398 143
rect 315 142 316 143
rect 314 142 315 143
rect 313 142 314 143
rect 312 142 313 143
rect 311 142 312 143
rect 310 142 311 143
rect 309 142 310 143
rect 308 142 309 143
rect 307 142 308 143
rect 306 142 307 143
rect 305 142 306 143
rect 304 142 305 143
rect 303 142 304 143
rect 302 142 303 143
rect 301 142 302 143
rect 300 142 301 143
rect 299 142 300 143
rect 298 142 299 143
rect 297 142 298 143
rect 296 142 297 143
rect 295 142 296 143
rect 294 142 295 143
rect 293 142 294 143
rect 292 142 293 143
rect 291 142 292 143
rect 290 142 291 143
rect 289 142 290 143
rect 288 142 289 143
rect 287 142 288 143
rect 286 142 287 143
rect 285 142 286 143
rect 284 142 285 143
rect 283 142 284 143
rect 282 142 283 143
rect 281 142 282 143
rect 280 142 281 143
rect 279 142 280 143
rect 278 142 279 143
rect 277 142 278 143
rect 276 142 277 143
rect 275 142 276 143
rect 274 142 275 143
rect 273 142 274 143
rect 272 142 273 143
rect 271 142 272 143
rect 270 142 271 143
rect 269 142 270 143
rect 268 142 269 143
rect 267 142 268 143
rect 266 142 267 143
rect 265 142 266 143
rect 264 142 265 143
rect 263 142 264 143
rect 262 142 263 143
rect 261 142 262 143
rect 260 142 261 143
rect 259 142 260 143
rect 258 142 259 143
rect 257 142 258 143
rect 256 142 257 143
rect 255 142 256 143
rect 254 142 255 143
rect 253 142 254 143
rect 252 142 253 143
rect 251 142 252 143
rect 250 142 251 143
rect 249 142 250 143
rect 225 142 226 143
rect 224 142 225 143
rect 223 142 224 143
rect 222 142 223 143
rect 221 142 222 143
rect 220 142 221 143
rect 219 142 220 143
rect 218 142 219 143
rect 217 142 218 143
rect 216 142 217 143
rect 215 142 216 143
rect 214 142 215 143
rect 213 142 214 143
rect 212 142 213 143
rect 211 142 212 143
rect 210 142 211 143
rect 209 142 210 143
rect 208 142 209 143
rect 207 142 208 143
rect 206 142 207 143
rect 205 142 206 143
rect 204 142 205 143
rect 203 142 204 143
rect 202 142 203 143
rect 201 142 202 143
rect 200 142 201 143
rect 199 142 200 143
rect 198 142 199 143
rect 197 142 198 143
rect 196 142 197 143
rect 195 142 196 143
rect 194 142 195 143
rect 193 142 194 143
rect 192 142 193 143
rect 191 142 192 143
rect 190 142 191 143
rect 189 142 190 143
rect 188 142 189 143
rect 187 142 188 143
rect 186 142 187 143
rect 185 142 186 143
rect 184 142 185 143
rect 183 142 184 143
rect 182 142 183 143
rect 181 142 182 143
rect 180 142 181 143
rect 179 142 180 143
rect 178 142 179 143
rect 177 142 178 143
rect 176 142 177 143
rect 175 142 176 143
rect 174 142 175 143
rect 173 142 174 143
rect 172 142 173 143
rect 171 142 172 143
rect 170 142 171 143
rect 169 142 170 143
rect 168 142 169 143
rect 167 142 168 143
rect 166 142 167 143
rect 165 142 166 143
rect 164 142 165 143
rect 163 142 164 143
rect 162 142 163 143
rect 142 142 143 143
rect 141 142 142 143
rect 140 142 141 143
rect 139 142 140 143
rect 138 142 139 143
rect 137 142 138 143
rect 136 142 137 143
rect 135 142 136 143
rect 134 142 135 143
rect 133 142 134 143
rect 132 142 133 143
rect 131 142 132 143
rect 130 142 131 143
rect 129 142 130 143
rect 128 142 129 143
rect 127 142 128 143
rect 126 142 127 143
rect 125 142 126 143
rect 124 142 125 143
rect 123 142 124 143
rect 122 142 123 143
rect 121 142 122 143
rect 120 142 121 143
rect 119 142 120 143
rect 118 142 119 143
rect 117 142 118 143
rect 116 142 117 143
rect 115 142 116 143
rect 114 142 115 143
rect 113 142 114 143
rect 112 142 113 143
rect 111 142 112 143
rect 110 142 111 143
rect 109 142 110 143
rect 108 142 109 143
rect 107 142 108 143
rect 106 142 107 143
rect 105 142 106 143
rect 104 142 105 143
rect 103 142 104 143
rect 102 142 103 143
rect 101 142 102 143
rect 100 142 101 143
rect 99 142 100 143
rect 98 142 99 143
rect 97 142 98 143
rect 96 142 97 143
rect 95 142 96 143
rect 94 142 95 143
rect 93 142 94 143
rect 92 142 93 143
rect 91 142 92 143
rect 90 142 91 143
rect 89 142 90 143
rect 88 142 89 143
rect 87 142 88 143
rect 86 142 87 143
rect 85 142 86 143
rect 84 142 85 143
rect 83 142 84 143
rect 82 142 83 143
rect 81 142 82 143
rect 80 142 81 143
rect 79 142 80 143
rect 78 142 79 143
rect 77 142 78 143
rect 76 142 77 143
rect 75 142 76 143
rect 74 142 75 143
rect 73 142 74 143
rect 72 142 73 143
rect 71 142 72 143
rect 70 142 71 143
rect 69 142 70 143
rect 68 142 69 143
rect 67 142 68 143
rect 66 142 67 143
rect 65 142 66 143
rect 64 142 65 143
rect 63 142 64 143
rect 62 142 63 143
rect 61 142 62 143
rect 60 142 61 143
rect 59 142 60 143
rect 58 142 59 143
rect 57 142 58 143
rect 56 142 57 143
rect 55 142 56 143
rect 54 142 55 143
rect 53 142 54 143
rect 52 142 53 143
rect 51 142 52 143
rect 50 142 51 143
rect 49 142 50 143
rect 48 142 49 143
rect 47 142 48 143
rect 46 142 47 143
rect 45 142 46 143
rect 44 142 45 143
rect 43 142 44 143
rect 42 142 43 143
rect 41 142 42 143
rect 40 142 41 143
rect 435 143 436 144
rect 434 143 435 144
rect 433 143 434 144
rect 432 143 433 144
rect 431 143 432 144
rect 430 143 431 144
rect 429 143 430 144
rect 428 143 429 144
rect 427 143 428 144
rect 426 143 427 144
rect 425 143 426 144
rect 424 143 425 144
rect 423 143 424 144
rect 422 143 423 144
rect 421 143 422 144
rect 420 143 421 144
rect 419 143 420 144
rect 418 143 419 144
rect 417 143 418 144
rect 416 143 417 144
rect 415 143 416 144
rect 414 143 415 144
rect 413 143 414 144
rect 412 143 413 144
rect 411 143 412 144
rect 410 143 411 144
rect 409 143 410 144
rect 408 143 409 144
rect 407 143 408 144
rect 406 143 407 144
rect 405 143 406 144
rect 404 143 405 144
rect 403 143 404 144
rect 402 143 403 144
rect 401 143 402 144
rect 400 143 401 144
rect 399 143 400 144
rect 398 143 399 144
rect 397 143 398 144
rect 315 143 316 144
rect 314 143 315 144
rect 313 143 314 144
rect 312 143 313 144
rect 311 143 312 144
rect 310 143 311 144
rect 309 143 310 144
rect 308 143 309 144
rect 307 143 308 144
rect 306 143 307 144
rect 305 143 306 144
rect 304 143 305 144
rect 303 143 304 144
rect 302 143 303 144
rect 301 143 302 144
rect 300 143 301 144
rect 299 143 300 144
rect 298 143 299 144
rect 297 143 298 144
rect 296 143 297 144
rect 295 143 296 144
rect 294 143 295 144
rect 293 143 294 144
rect 292 143 293 144
rect 291 143 292 144
rect 290 143 291 144
rect 289 143 290 144
rect 288 143 289 144
rect 287 143 288 144
rect 286 143 287 144
rect 285 143 286 144
rect 284 143 285 144
rect 283 143 284 144
rect 282 143 283 144
rect 281 143 282 144
rect 280 143 281 144
rect 279 143 280 144
rect 278 143 279 144
rect 277 143 278 144
rect 276 143 277 144
rect 275 143 276 144
rect 274 143 275 144
rect 273 143 274 144
rect 272 143 273 144
rect 271 143 272 144
rect 270 143 271 144
rect 269 143 270 144
rect 268 143 269 144
rect 267 143 268 144
rect 266 143 267 144
rect 265 143 266 144
rect 264 143 265 144
rect 263 143 264 144
rect 262 143 263 144
rect 261 143 262 144
rect 260 143 261 144
rect 259 143 260 144
rect 258 143 259 144
rect 257 143 258 144
rect 256 143 257 144
rect 255 143 256 144
rect 254 143 255 144
rect 253 143 254 144
rect 252 143 253 144
rect 251 143 252 144
rect 250 143 251 144
rect 249 143 250 144
rect 248 143 249 144
rect 224 143 225 144
rect 223 143 224 144
rect 222 143 223 144
rect 221 143 222 144
rect 220 143 221 144
rect 219 143 220 144
rect 218 143 219 144
rect 217 143 218 144
rect 216 143 217 144
rect 215 143 216 144
rect 214 143 215 144
rect 213 143 214 144
rect 212 143 213 144
rect 211 143 212 144
rect 210 143 211 144
rect 209 143 210 144
rect 208 143 209 144
rect 207 143 208 144
rect 206 143 207 144
rect 205 143 206 144
rect 204 143 205 144
rect 203 143 204 144
rect 202 143 203 144
rect 201 143 202 144
rect 200 143 201 144
rect 199 143 200 144
rect 198 143 199 144
rect 197 143 198 144
rect 196 143 197 144
rect 195 143 196 144
rect 194 143 195 144
rect 193 143 194 144
rect 192 143 193 144
rect 191 143 192 144
rect 190 143 191 144
rect 189 143 190 144
rect 188 143 189 144
rect 187 143 188 144
rect 186 143 187 144
rect 185 143 186 144
rect 184 143 185 144
rect 183 143 184 144
rect 182 143 183 144
rect 181 143 182 144
rect 180 143 181 144
rect 179 143 180 144
rect 178 143 179 144
rect 177 143 178 144
rect 176 143 177 144
rect 175 143 176 144
rect 174 143 175 144
rect 173 143 174 144
rect 172 143 173 144
rect 171 143 172 144
rect 170 143 171 144
rect 169 143 170 144
rect 168 143 169 144
rect 167 143 168 144
rect 166 143 167 144
rect 165 143 166 144
rect 164 143 165 144
rect 163 143 164 144
rect 162 143 163 144
rect 161 143 162 144
rect 141 143 142 144
rect 140 143 141 144
rect 139 143 140 144
rect 138 143 139 144
rect 137 143 138 144
rect 136 143 137 144
rect 135 143 136 144
rect 134 143 135 144
rect 133 143 134 144
rect 132 143 133 144
rect 131 143 132 144
rect 130 143 131 144
rect 129 143 130 144
rect 128 143 129 144
rect 127 143 128 144
rect 126 143 127 144
rect 125 143 126 144
rect 124 143 125 144
rect 123 143 124 144
rect 122 143 123 144
rect 121 143 122 144
rect 120 143 121 144
rect 119 143 120 144
rect 118 143 119 144
rect 117 143 118 144
rect 116 143 117 144
rect 115 143 116 144
rect 114 143 115 144
rect 113 143 114 144
rect 112 143 113 144
rect 111 143 112 144
rect 110 143 111 144
rect 109 143 110 144
rect 108 143 109 144
rect 107 143 108 144
rect 106 143 107 144
rect 105 143 106 144
rect 104 143 105 144
rect 103 143 104 144
rect 102 143 103 144
rect 101 143 102 144
rect 100 143 101 144
rect 99 143 100 144
rect 98 143 99 144
rect 97 143 98 144
rect 96 143 97 144
rect 95 143 96 144
rect 94 143 95 144
rect 93 143 94 144
rect 92 143 93 144
rect 91 143 92 144
rect 90 143 91 144
rect 89 143 90 144
rect 88 143 89 144
rect 87 143 88 144
rect 86 143 87 144
rect 85 143 86 144
rect 84 143 85 144
rect 83 143 84 144
rect 82 143 83 144
rect 81 143 82 144
rect 80 143 81 144
rect 79 143 80 144
rect 78 143 79 144
rect 77 143 78 144
rect 76 143 77 144
rect 75 143 76 144
rect 74 143 75 144
rect 73 143 74 144
rect 72 143 73 144
rect 71 143 72 144
rect 70 143 71 144
rect 69 143 70 144
rect 68 143 69 144
rect 67 143 68 144
rect 66 143 67 144
rect 65 143 66 144
rect 64 143 65 144
rect 63 143 64 144
rect 62 143 63 144
rect 61 143 62 144
rect 60 143 61 144
rect 59 143 60 144
rect 58 143 59 144
rect 57 143 58 144
rect 56 143 57 144
rect 55 143 56 144
rect 54 143 55 144
rect 53 143 54 144
rect 52 143 53 144
rect 51 143 52 144
rect 50 143 51 144
rect 49 143 50 144
rect 48 143 49 144
rect 47 143 48 144
rect 46 143 47 144
rect 45 143 46 144
rect 44 143 45 144
rect 43 143 44 144
rect 42 143 43 144
rect 41 143 42 144
rect 482 144 483 145
rect 462 144 463 145
rect 433 144 434 145
rect 432 144 433 145
rect 431 144 432 145
rect 430 144 431 145
rect 429 144 430 145
rect 428 144 429 145
rect 427 144 428 145
rect 426 144 427 145
rect 425 144 426 145
rect 424 144 425 145
rect 423 144 424 145
rect 422 144 423 145
rect 421 144 422 145
rect 420 144 421 145
rect 419 144 420 145
rect 418 144 419 145
rect 417 144 418 145
rect 416 144 417 145
rect 415 144 416 145
rect 414 144 415 145
rect 413 144 414 145
rect 412 144 413 145
rect 411 144 412 145
rect 410 144 411 145
rect 409 144 410 145
rect 408 144 409 145
rect 407 144 408 145
rect 406 144 407 145
rect 405 144 406 145
rect 404 144 405 145
rect 403 144 404 145
rect 402 144 403 145
rect 401 144 402 145
rect 400 144 401 145
rect 399 144 400 145
rect 398 144 399 145
rect 397 144 398 145
rect 316 144 317 145
rect 315 144 316 145
rect 314 144 315 145
rect 313 144 314 145
rect 312 144 313 145
rect 311 144 312 145
rect 310 144 311 145
rect 309 144 310 145
rect 308 144 309 145
rect 307 144 308 145
rect 306 144 307 145
rect 305 144 306 145
rect 304 144 305 145
rect 303 144 304 145
rect 302 144 303 145
rect 301 144 302 145
rect 300 144 301 145
rect 299 144 300 145
rect 298 144 299 145
rect 297 144 298 145
rect 296 144 297 145
rect 295 144 296 145
rect 294 144 295 145
rect 293 144 294 145
rect 292 144 293 145
rect 291 144 292 145
rect 290 144 291 145
rect 289 144 290 145
rect 288 144 289 145
rect 287 144 288 145
rect 286 144 287 145
rect 285 144 286 145
rect 284 144 285 145
rect 283 144 284 145
rect 282 144 283 145
rect 281 144 282 145
rect 280 144 281 145
rect 279 144 280 145
rect 278 144 279 145
rect 277 144 278 145
rect 276 144 277 145
rect 275 144 276 145
rect 274 144 275 145
rect 273 144 274 145
rect 272 144 273 145
rect 271 144 272 145
rect 270 144 271 145
rect 269 144 270 145
rect 268 144 269 145
rect 267 144 268 145
rect 266 144 267 145
rect 265 144 266 145
rect 264 144 265 145
rect 263 144 264 145
rect 262 144 263 145
rect 261 144 262 145
rect 260 144 261 145
rect 259 144 260 145
rect 258 144 259 145
rect 257 144 258 145
rect 256 144 257 145
rect 255 144 256 145
rect 254 144 255 145
rect 253 144 254 145
rect 252 144 253 145
rect 251 144 252 145
rect 250 144 251 145
rect 249 144 250 145
rect 248 144 249 145
rect 247 144 248 145
rect 224 144 225 145
rect 223 144 224 145
rect 222 144 223 145
rect 221 144 222 145
rect 220 144 221 145
rect 219 144 220 145
rect 218 144 219 145
rect 217 144 218 145
rect 216 144 217 145
rect 215 144 216 145
rect 214 144 215 145
rect 213 144 214 145
rect 212 144 213 145
rect 211 144 212 145
rect 210 144 211 145
rect 209 144 210 145
rect 208 144 209 145
rect 207 144 208 145
rect 206 144 207 145
rect 205 144 206 145
rect 204 144 205 145
rect 203 144 204 145
rect 202 144 203 145
rect 201 144 202 145
rect 200 144 201 145
rect 199 144 200 145
rect 198 144 199 145
rect 197 144 198 145
rect 196 144 197 145
rect 195 144 196 145
rect 194 144 195 145
rect 193 144 194 145
rect 192 144 193 145
rect 191 144 192 145
rect 190 144 191 145
rect 189 144 190 145
rect 188 144 189 145
rect 187 144 188 145
rect 186 144 187 145
rect 185 144 186 145
rect 184 144 185 145
rect 183 144 184 145
rect 182 144 183 145
rect 181 144 182 145
rect 180 144 181 145
rect 179 144 180 145
rect 178 144 179 145
rect 177 144 178 145
rect 176 144 177 145
rect 175 144 176 145
rect 174 144 175 145
rect 173 144 174 145
rect 172 144 173 145
rect 171 144 172 145
rect 170 144 171 145
rect 169 144 170 145
rect 168 144 169 145
rect 167 144 168 145
rect 166 144 167 145
rect 165 144 166 145
rect 164 144 165 145
rect 163 144 164 145
rect 162 144 163 145
rect 161 144 162 145
rect 140 144 141 145
rect 139 144 140 145
rect 138 144 139 145
rect 137 144 138 145
rect 136 144 137 145
rect 135 144 136 145
rect 134 144 135 145
rect 133 144 134 145
rect 132 144 133 145
rect 131 144 132 145
rect 130 144 131 145
rect 129 144 130 145
rect 128 144 129 145
rect 127 144 128 145
rect 126 144 127 145
rect 125 144 126 145
rect 124 144 125 145
rect 123 144 124 145
rect 122 144 123 145
rect 121 144 122 145
rect 120 144 121 145
rect 119 144 120 145
rect 118 144 119 145
rect 117 144 118 145
rect 116 144 117 145
rect 115 144 116 145
rect 114 144 115 145
rect 113 144 114 145
rect 112 144 113 145
rect 111 144 112 145
rect 110 144 111 145
rect 109 144 110 145
rect 108 144 109 145
rect 107 144 108 145
rect 106 144 107 145
rect 105 144 106 145
rect 104 144 105 145
rect 103 144 104 145
rect 102 144 103 145
rect 101 144 102 145
rect 100 144 101 145
rect 99 144 100 145
rect 98 144 99 145
rect 97 144 98 145
rect 96 144 97 145
rect 95 144 96 145
rect 94 144 95 145
rect 93 144 94 145
rect 92 144 93 145
rect 91 144 92 145
rect 90 144 91 145
rect 89 144 90 145
rect 88 144 89 145
rect 87 144 88 145
rect 86 144 87 145
rect 85 144 86 145
rect 84 144 85 145
rect 83 144 84 145
rect 82 144 83 145
rect 81 144 82 145
rect 80 144 81 145
rect 79 144 80 145
rect 78 144 79 145
rect 77 144 78 145
rect 76 144 77 145
rect 75 144 76 145
rect 74 144 75 145
rect 73 144 74 145
rect 72 144 73 145
rect 71 144 72 145
rect 70 144 71 145
rect 69 144 70 145
rect 68 144 69 145
rect 67 144 68 145
rect 66 144 67 145
rect 65 144 66 145
rect 64 144 65 145
rect 63 144 64 145
rect 62 144 63 145
rect 61 144 62 145
rect 60 144 61 145
rect 59 144 60 145
rect 58 144 59 145
rect 57 144 58 145
rect 56 144 57 145
rect 55 144 56 145
rect 54 144 55 145
rect 53 144 54 145
rect 52 144 53 145
rect 51 144 52 145
rect 50 144 51 145
rect 49 144 50 145
rect 48 144 49 145
rect 47 144 48 145
rect 46 144 47 145
rect 45 144 46 145
rect 44 144 45 145
rect 43 144 44 145
rect 42 144 43 145
rect 41 144 42 145
rect 26 144 27 145
rect 25 144 26 145
rect 24 144 25 145
rect 23 144 24 145
rect 22 144 23 145
rect 482 145 483 146
rect 462 145 463 146
rect 429 145 430 146
rect 428 145 429 146
rect 427 145 428 146
rect 426 145 427 146
rect 425 145 426 146
rect 424 145 425 146
rect 423 145 424 146
rect 422 145 423 146
rect 421 145 422 146
rect 420 145 421 146
rect 419 145 420 146
rect 418 145 419 146
rect 417 145 418 146
rect 416 145 417 146
rect 415 145 416 146
rect 414 145 415 146
rect 413 145 414 146
rect 412 145 413 146
rect 411 145 412 146
rect 410 145 411 146
rect 409 145 410 146
rect 408 145 409 146
rect 407 145 408 146
rect 406 145 407 146
rect 405 145 406 146
rect 404 145 405 146
rect 403 145 404 146
rect 402 145 403 146
rect 401 145 402 146
rect 400 145 401 146
rect 399 145 400 146
rect 398 145 399 146
rect 397 145 398 146
rect 317 145 318 146
rect 316 145 317 146
rect 315 145 316 146
rect 314 145 315 146
rect 313 145 314 146
rect 312 145 313 146
rect 311 145 312 146
rect 310 145 311 146
rect 309 145 310 146
rect 308 145 309 146
rect 307 145 308 146
rect 306 145 307 146
rect 305 145 306 146
rect 304 145 305 146
rect 303 145 304 146
rect 302 145 303 146
rect 301 145 302 146
rect 300 145 301 146
rect 299 145 300 146
rect 298 145 299 146
rect 297 145 298 146
rect 296 145 297 146
rect 295 145 296 146
rect 294 145 295 146
rect 293 145 294 146
rect 292 145 293 146
rect 291 145 292 146
rect 290 145 291 146
rect 289 145 290 146
rect 288 145 289 146
rect 287 145 288 146
rect 286 145 287 146
rect 285 145 286 146
rect 284 145 285 146
rect 283 145 284 146
rect 282 145 283 146
rect 281 145 282 146
rect 280 145 281 146
rect 279 145 280 146
rect 278 145 279 146
rect 277 145 278 146
rect 276 145 277 146
rect 275 145 276 146
rect 274 145 275 146
rect 273 145 274 146
rect 272 145 273 146
rect 271 145 272 146
rect 270 145 271 146
rect 269 145 270 146
rect 268 145 269 146
rect 267 145 268 146
rect 266 145 267 146
rect 265 145 266 146
rect 264 145 265 146
rect 263 145 264 146
rect 262 145 263 146
rect 261 145 262 146
rect 260 145 261 146
rect 259 145 260 146
rect 258 145 259 146
rect 257 145 258 146
rect 256 145 257 146
rect 255 145 256 146
rect 254 145 255 146
rect 253 145 254 146
rect 252 145 253 146
rect 251 145 252 146
rect 250 145 251 146
rect 249 145 250 146
rect 248 145 249 146
rect 247 145 248 146
rect 246 145 247 146
rect 223 145 224 146
rect 222 145 223 146
rect 221 145 222 146
rect 220 145 221 146
rect 219 145 220 146
rect 218 145 219 146
rect 217 145 218 146
rect 216 145 217 146
rect 215 145 216 146
rect 214 145 215 146
rect 213 145 214 146
rect 212 145 213 146
rect 211 145 212 146
rect 210 145 211 146
rect 209 145 210 146
rect 208 145 209 146
rect 207 145 208 146
rect 206 145 207 146
rect 205 145 206 146
rect 204 145 205 146
rect 203 145 204 146
rect 202 145 203 146
rect 201 145 202 146
rect 200 145 201 146
rect 199 145 200 146
rect 198 145 199 146
rect 197 145 198 146
rect 196 145 197 146
rect 195 145 196 146
rect 194 145 195 146
rect 193 145 194 146
rect 192 145 193 146
rect 191 145 192 146
rect 190 145 191 146
rect 189 145 190 146
rect 188 145 189 146
rect 187 145 188 146
rect 186 145 187 146
rect 185 145 186 146
rect 184 145 185 146
rect 183 145 184 146
rect 182 145 183 146
rect 181 145 182 146
rect 180 145 181 146
rect 179 145 180 146
rect 178 145 179 146
rect 177 145 178 146
rect 176 145 177 146
rect 175 145 176 146
rect 174 145 175 146
rect 173 145 174 146
rect 172 145 173 146
rect 171 145 172 146
rect 170 145 171 146
rect 169 145 170 146
rect 168 145 169 146
rect 167 145 168 146
rect 166 145 167 146
rect 165 145 166 146
rect 164 145 165 146
rect 163 145 164 146
rect 162 145 163 146
rect 161 145 162 146
rect 160 145 161 146
rect 139 145 140 146
rect 138 145 139 146
rect 137 145 138 146
rect 136 145 137 146
rect 135 145 136 146
rect 134 145 135 146
rect 133 145 134 146
rect 132 145 133 146
rect 131 145 132 146
rect 130 145 131 146
rect 129 145 130 146
rect 128 145 129 146
rect 127 145 128 146
rect 126 145 127 146
rect 125 145 126 146
rect 124 145 125 146
rect 123 145 124 146
rect 122 145 123 146
rect 121 145 122 146
rect 120 145 121 146
rect 119 145 120 146
rect 118 145 119 146
rect 117 145 118 146
rect 116 145 117 146
rect 115 145 116 146
rect 114 145 115 146
rect 113 145 114 146
rect 112 145 113 146
rect 111 145 112 146
rect 110 145 111 146
rect 109 145 110 146
rect 108 145 109 146
rect 107 145 108 146
rect 106 145 107 146
rect 105 145 106 146
rect 104 145 105 146
rect 103 145 104 146
rect 102 145 103 146
rect 101 145 102 146
rect 100 145 101 146
rect 99 145 100 146
rect 98 145 99 146
rect 97 145 98 146
rect 96 145 97 146
rect 95 145 96 146
rect 94 145 95 146
rect 93 145 94 146
rect 92 145 93 146
rect 91 145 92 146
rect 90 145 91 146
rect 89 145 90 146
rect 88 145 89 146
rect 87 145 88 146
rect 86 145 87 146
rect 85 145 86 146
rect 84 145 85 146
rect 83 145 84 146
rect 82 145 83 146
rect 81 145 82 146
rect 80 145 81 146
rect 79 145 80 146
rect 78 145 79 146
rect 77 145 78 146
rect 76 145 77 146
rect 75 145 76 146
rect 74 145 75 146
rect 73 145 74 146
rect 72 145 73 146
rect 71 145 72 146
rect 70 145 71 146
rect 69 145 70 146
rect 68 145 69 146
rect 67 145 68 146
rect 66 145 67 146
rect 65 145 66 146
rect 64 145 65 146
rect 63 145 64 146
rect 62 145 63 146
rect 61 145 62 146
rect 60 145 61 146
rect 59 145 60 146
rect 58 145 59 146
rect 57 145 58 146
rect 56 145 57 146
rect 55 145 56 146
rect 54 145 55 146
rect 53 145 54 146
rect 52 145 53 146
rect 51 145 52 146
rect 50 145 51 146
rect 49 145 50 146
rect 48 145 49 146
rect 47 145 48 146
rect 46 145 47 146
rect 45 145 46 146
rect 44 145 45 146
rect 43 145 44 146
rect 42 145 43 146
rect 28 145 29 146
rect 27 145 28 146
rect 26 145 27 146
rect 25 145 26 146
rect 24 145 25 146
rect 23 145 24 146
rect 22 145 23 146
rect 21 145 22 146
rect 20 145 21 146
rect 19 145 20 146
rect 482 146 483 147
rect 481 146 482 147
rect 463 146 464 147
rect 462 146 463 147
rect 406 146 407 147
rect 405 146 406 147
rect 404 146 405 147
rect 403 146 404 147
rect 402 146 403 147
rect 401 146 402 147
rect 400 146 401 147
rect 399 146 400 147
rect 398 146 399 147
rect 397 146 398 147
rect 318 146 319 147
rect 317 146 318 147
rect 316 146 317 147
rect 315 146 316 147
rect 314 146 315 147
rect 313 146 314 147
rect 312 146 313 147
rect 311 146 312 147
rect 310 146 311 147
rect 309 146 310 147
rect 308 146 309 147
rect 307 146 308 147
rect 306 146 307 147
rect 305 146 306 147
rect 304 146 305 147
rect 303 146 304 147
rect 302 146 303 147
rect 301 146 302 147
rect 300 146 301 147
rect 299 146 300 147
rect 298 146 299 147
rect 297 146 298 147
rect 296 146 297 147
rect 295 146 296 147
rect 294 146 295 147
rect 293 146 294 147
rect 292 146 293 147
rect 291 146 292 147
rect 290 146 291 147
rect 289 146 290 147
rect 288 146 289 147
rect 287 146 288 147
rect 286 146 287 147
rect 285 146 286 147
rect 284 146 285 147
rect 283 146 284 147
rect 282 146 283 147
rect 281 146 282 147
rect 280 146 281 147
rect 279 146 280 147
rect 278 146 279 147
rect 277 146 278 147
rect 276 146 277 147
rect 275 146 276 147
rect 274 146 275 147
rect 273 146 274 147
rect 272 146 273 147
rect 271 146 272 147
rect 270 146 271 147
rect 269 146 270 147
rect 268 146 269 147
rect 267 146 268 147
rect 266 146 267 147
rect 265 146 266 147
rect 264 146 265 147
rect 263 146 264 147
rect 262 146 263 147
rect 261 146 262 147
rect 260 146 261 147
rect 259 146 260 147
rect 258 146 259 147
rect 257 146 258 147
rect 256 146 257 147
rect 255 146 256 147
rect 254 146 255 147
rect 253 146 254 147
rect 252 146 253 147
rect 251 146 252 147
rect 250 146 251 147
rect 249 146 250 147
rect 248 146 249 147
rect 247 146 248 147
rect 246 146 247 147
rect 245 146 246 147
rect 223 146 224 147
rect 222 146 223 147
rect 221 146 222 147
rect 220 146 221 147
rect 219 146 220 147
rect 218 146 219 147
rect 217 146 218 147
rect 216 146 217 147
rect 215 146 216 147
rect 214 146 215 147
rect 213 146 214 147
rect 212 146 213 147
rect 211 146 212 147
rect 210 146 211 147
rect 209 146 210 147
rect 208 146 209 147
rect 207 146 208 147
rect 206 146 207 147
rect 205 146 206 147
rect 204 146 205 147
rect 203 146 204 147
rect 202 146 203 147
rect 201 146 202 147
rect 200 146 201 147
rect 199 146 200 147
rect 198 146 199 147
rect 197 146 198 147
rect 196 146 197 147
rect 195 146 196 147
rect 194 146 195 147
rect 193 146 194 147
rect 192 146 193 147
rect 191 146 192 147
rect 190 146 191 147
rect 189 146 190 147
rect 188 146 189 147
rect 187 146 188 147
rect 186 146 187 147
rect 185 146 186 147
rect 184 146 185 147
rect 183 146 184 147
rect 182 146 183 147
rect 181 146 182 147
rect 180 146 181 147
rect 179 146 180 147
rect 178 146 179 147
rect 177 146 178 147
rect 176 146 177 147
rect 175 146 176 147
rect 174 146 175 147
rect 173 146 174 147
rect 172 146 173 147
rect 171 146 172 147
rect 170 146 171 147
rect 169 146 170 147
rect 168 146 169 147
rect 167 146 168 147
rect 166 146 167 147
rect 165 146 166 147
rect 164 146 165 147
rect 163 146 164 147
rect 162 146 163 147
rect 161 146 162 147
rect 160 146 161 147
rect 138 146 139 147
rect 137 146 138 147
rect 136 146 137 147
rect 135 146 136 147
rect 134 146 135 147
rect 133 146 134 147
rect 132 146 133 147
rect 131 146 132 147
rect 130 146 131 147
rect 129 146 130 147
rect 128 146 129 147
rect 127 146 128 147
rect 126 146 127 147
rect 125 146 126 147
rect 124 146 125 147
rect 123 146 124 147
rect 122 146 123 147
rect 121 146 122 147
rect 120 146 121 147
rect 119 146 120 147
rect 118 146 119 147
rect 117 146 118 147
rect 116 146 117 147
rect 115 146 116 147
rect 114 146 115 147
rect 113 146 114 147
rect 112 146 113 147
rect 111 146 112 147
rect 110 146 111 147
rect 109 146 110 147
rect 108 146 109 147
rect 107 146 108 147
rect 106 146 107 147
rect 105 146 106 147
rect 104 146 105 147
rect 103 146 104 147
rect 102 146 103 147
rect 101 146 102 147
rect 100 146 101 147
rect 99 146 100 147
rect 98 146 99 147
rect 97 146 98 147
rect 96 146 97 147
rect 95 146 96 147
rect 94 146 95 147
rect 93 146 94 147
rect 92 146 93 147
rect 91 146 92 147
rect 90 146 91 147
rect 89 146 90 147
rect 88 146 89 147
rect 87 146 88 147
rect 86 146 87 147
rect 85 146 86 147
rect 84 146 85 147
rect 83 146 84 147
rect 82 146 83 147
rect 81 146 82 147
rect 80 146 81 147
rect 79 146 80 147
rect 78 146 79 147
rect 77 146 78 147
rect 76 146 77 147
rect 75 146 76 147
rect 74 146 75 147
rect 73 146 74 147
rect 72 146 73 147
rect 71 146 72 147
rect 70 146 71 147
rect 69 146 70 147
rect 68 146 69 147
rect 67 146 68 147
rect 66 146 67 147
rect 65 146 66 147
rect 64 146 65 147
rect 63 146 64 147
rect 62 146 63 147
rect 61 146 62 147
rect 60 146 61 147
rect 59 146 60 147
rect 58 146 59 147
rect 57 146 58 147
rect 56 146 57 147
rect 55 146 56 147
rect 54 146 55 147
rect 53 146 54 147
rect 52 146 53 147
rect 51 146 52 147
rect 50 146 51 147
rect 49 146 50 147
rect 48 146 49 147
rect 47 146 48 147
rect 46 146 47 147
rect 45 146 46 147
rect 44 146 45 147
rect 43 146 44 147
rect 42 146 43 147
rect 29 146 30 147
rect 28 146 29 147
rect 27 146 28 147
rect 26 146 27 147
rect 25 146 26 147
rect 24 146 25 147
rect 23 146 24 147
rect 22 146 23 147
rect 21 146 22 147
rect 20 146 21 147
rect 19 146 20 147
rect 18 146 19 147
rect 482 147 483 148
rect 481 147 482 148
rect 480 147 481 148
rect 479 147 480 148
rect 478 147 479 148
rect 477 147 478 148
rect 476 147 477 148
rect 475 147 476 148
rect 474 147 475 148
rect 473 147 474 148
rect 472 147 473 148
rect 471 147 472 148
rect 470 147 471 148
rect 469 147 470 148
rect 468 147 469 148
rect 467 147 468 148
rect 466 147 467 148
rect 465 147 466 148
rect 464 147 465 148
rect 463 147 464 148
rect 462 147 463 148
rect 401 147 402 148
rect 400 147 401 148
rect 399 147 400 148
rect 398 147 399 148
rect 397 147 398 148
rect 318 147 319 148
rect 317 147 318 148
rect 316 147 317 148
rect 315 147 316 148
rect 314 147 315 148
rect 313 147 314 148
rect 312 147 313 148
rect 311 147 312 148
rect 310 147 311 148
rect 309 147 310 148
rect 308 147 309 148
rect 307 147 308 148
rect 306 147 307 148
rect 305 147 306 148
rect 304 147 305 148
rect 303 147 304 148
rect 302 147 303 148
rect 301 147 302 148
rect 300 147 301 148
rect 299 147 300 148
rect 298 147 299 148
rect 297 147 298 148
rect 296 147 297 148
rect 295 147 296 148
rect 294 147 295 148
rect 293 147 294 148
rect 292 147 293 148
rect 291 147 292 148
rect 290 147 291 148
rect 289 147 290 148
rect 288 147 289 148
rect 287 147 288 148
rect 286 147 287 148
rect 285 147 286 148
rect 284 147 285 148
rect 283 147 284 148
rect 282 147 283 148
rect 281 147 282 148
rect 280 147 281 148
rect 279 147 280 148
rect 278 147 279 148
rect 277 147 278 148
rect 276 147 277 148
rect 275 147 276 148
rect 274 147 275 148
rect 273 147 274 148
rect 272 147 273 148
rect 271 147 272 148
rect 270 147 271 148
rect 269 147 270 148
rect 268 147 269 148
rect 267 147 268 148
rect 266 147 267 148
rect 265 147 266 148
rect 264 147 265 148
rect 263 147 264 148
rect 262 147 263 148
rect 261 147 262 148
rect 260 147 261 148
rect 259 147 260 148
rect 258 147 259 148
rect 257 147 258 148
rect 256 147 257 148
rect 255 147 256 148
rect 254 147 255 148
rect 253 147 254 148
rect 252 147 253 148
rect 251 147 252 148
rect 250 147 251 148
rect 249 147 250 148
rect 248 147 249 148
rect 247 147 248 148
rect 246 147 247 148
rect 245 147 246 148
rect 223 147 224 148
rect 222 147 223 148
rect 221 147 222 148
rect 220 147 221 148
rect 219 147 220 148
rect 218 147 219 148
rect 217 147 218 148
rect 216 147 217 148
rect 215 147 216 148
rect 214 147 215 148
rect 213 147 214 148
rect 212 147 213 148
rect 211 147 212 148
rect 210 147 211 148
rect 209 147 210 148
rect 208 147 209 148
rect 207 147 208 148
rect 206 147 207 148
rect 205 147 206 148
rect 204 147 205 148
rect 203 147 204 148
rect 202 147 203 148
rect 201 147 202 148
rect 200 147 201 148
rect 199 147 200 148
rect 198 147 199 148
rect 197 147 198 148
rect 196 147 197 148
rect 195 147 196 148
rect 194 147 195 148
rect 193 147 194 148
rect 192 147 193 148
rect 191 147 192 148
rect 190 147 191 148
rect 189 147 190 148
rect 188 147 189 148
rect 187 147 188 148
rect 186 147 187 148
rect 185 147 186 148
rect 184 147 185 148
rect 183 147 184 148
rect 182 147 183 148
rect 181 147 182 148
rect 180 147 181 148
rect 179 147 180 148
rect 178 147 179 148
rect 177 147 178 148
rect 176 147 177 148
rect 175 147 176 148
rect 174 147 175 148
rect 173 147 174 148
rect 172 147 173 148
rect 171 147 172 148
rect 170 147 171 148
rect 169 147 170 148
rect 168 147 169 148
rect 167 147 168 148
rect 166 147 167 148
rect 165 147 166 148
rect 164 147 165 148
rect 163 147 164 148
rect 162 147 163 148
rect 161 147 162 148
rect 160 147 161 148
rect 159 147 160 148
rect 137 147 138 148
rect 136 147 137 148
rect 135 147 136 148
rect 134 147 135 148
rect 133 147 134 148
rect 132 147 133 148
rect 131 147 132 148
rect 130 147 131 148
rect 129 147 130 148
rect 128 147 129 148
rect 127 147 128 148
rect 126 147 127 148
rect 125 147 126 148
rect 124 147 125 148
rect 123 147 124 148
rect 122 147 123 148
rect 121 147 122 148
rect 120 147 121 148
rect 119 147 120 148
rect 118 147 119 148
rect 117 147 118 148
rect 116 147 117 148
rect 115 147 116 148
rect 114 147 115 148
rect 113 147 114 148
rect 112 147 113 148
rect 111 147 112 148
rect 110 147 111 148
rect 109 147 110 148
rect 108 147 109 148
rect 107 147 108 148
rect 106 147 107 148
rect 105 147 106 148
rect 104 147 105 148
rect 103 147 104 148
rect 102 147 103 148
rect 101 147 102 148
rect 100 147 101 148
rect 99 147 100 148
rect 98 147 99 148
rect 97 147 98 148
rect 96 147 97 148
rect 95 147 96 148
rect 94 147 95 148
rect 93 147 94 148
rect 92 147 93 148
rect 91 147 92 148
rect 90 147 91 148
rect 89 147 90 148
rect 88 147 89 148
rect 87 147 88 148
rect 86 147 87 148
rect 85 147 86 148
rect 84 147 85 148
rect 83 147 84 148
rect 82 147 83 148
rect 81 147 82 148
rect 80 147 81 148
rect 79 147 80 148
rect 78 147 79 148
rect 77 147 78 148
rect 76 147 77 148
rect 75 147 76 148
rect 74 147 75 148
rect 73 147 74 148
rect 72 147 73 148
rect 71 147 72 148
rect 70 147 71 148
rect 69 147 70 148
rect 68 147 69 148
rect 67 147 68 148
rect 66 147 67 148
rect 65 147 66 148
rect 64 147 65 148
rect 63 147 64 148
rect 62 147 63 148
rect 61 147 62 148
rect 60 147 61 148
rect 59 147 60 148
rect 58 147 59 148
rect 57 147 58 148
rect 56 147 57 148
rect 55 147 56 148
rect 54 147 55 148
rect 53 147 54 148
rect 52 147 53 148
rect 51 147 52 148
rect 50 147 51 148
rect 49 147 50 148
rect 48 147 49 148
rect 47 147 48 148
rect 46 147 47 148
rect 45 147 46 148
rect 44 147 45 148
rect 43 147 44 148
rect 42 147 43 148
rect 30 147 31 148
rect 29 147 30 148
rect 28 147 29 148
rect 27 147 28 148
rect 26 147 27 148
rect 25 147 26 148
rect 24 147 25 148
rect 23 147 24 148
rect 22 147 23 148
rect 21 147 22 148
rect 20 147 21 148
rect 19 147 20 148
rect 18 147 19 148
rect 17 147 18 148
rect 16 147 17 148
rect 482 148 483 149
rect 481 148 482 149
rect 480 148 481 149
rect 479 148 480 149
rect 478 148 479 149
rect 477 148 478 149
rect 476 148 477 149
rect 475 148 476 149
rect 474 148 475 149
rect 473 148 474 149
rect 472 148 473 149
rect 471 148 472 149
rect 470 148 471 149
rect 469 148 470 149
rect 468 148 469 149
rect 467 148 468 149
rect 466 148 467 149
rect 465 148 466 149
rect 464 148 465 149
rect 463 148 464 149
rect 462 148 463 149
rect 400 148 401 149
rect 399 148 400 149
rect 398 148 399 149
rect 397 148 398 149
rect 319 148 320 149
rect 318 148 319 149
rect 317 148 318 149
rect 316 148 317 149
rect 315 148 316 149
rect 314 148 315 149
rect 313 148 314 149
rect 312 148 313 149
rect 311 148 312 149
rect 310 148 311 149
rect 309 148 310 149
rect 308 148 309 149
rect 307 148 308 149
rect 306 148 307 149
rect 305 148 306 149
rect 304 148 305 149
rect 303 148 304 149
rect 302 148 303 149
rect 301 148 302 149
rect 300 148 301 149
rect 299 148 300 149
rect 298 148 299 149
rect 297 148 298 149
rect 296 148 297 149
rect 295 148 296 149
rect 294 148 295 149
rect 293 148 294 149
rect 292 148 293 149
rect 291 148 292 149
rect 290 148 291 149
rect 289 148 290 149
rect 288 148 289 149
rect 287 148 288 149
rect 286 148 287 149
rect 285 148 286 149
rect 284 148 285 149
rect 283 148 284 149
rect 282 148 283 149
rect 281 148 282 149
rect 280 148 281 149
rect 279 148 280 149
rect 278 148 279 149
rect 277 148 278 149
rect 276 148 277 149
rect 275 148 276 149
rect 274 148 275 149
rect 273 148 274 149
rect 272 148 273 149
rect 271 148 272 149
rect 270 148 271 149
rect 269 148 270 149
rect 268 148 269 149
rect 267 148 268 149
rect 266 148 267 149
rect 265 148 266 149
rect 264 148 265 149
rect 263 148 264 149
rect 262 148 263 149
rect 261 148 262 149
rect 260 148 261 149
rect 259 148 260 149
rect 258 148 259 149
rect 257 148 258 149
rect 256 148 257 149
rect 255 148 256 149
rect 254 148 255 149
rect 253 148 254 149
rect 252 148 253 149
rect 251 148 252 149
rect 250 148 251 149
rect 249 148 250 149
rect 248 148 249 149
rect 247 148 248 149
rect 246 148 247 149
rect 245 148 246 149
rect 244 148 245 149
rect 222 148 223 149
rect 221 148 222 149
rect 220 148 221 149
rect 219 148 220 149
rect 218 148 219 149
rect 217 148 218 149
rect 216 148 217 149
rect 215 148 216 149
rect 214 148 215 149
rect 213 148 214 149
rect 212 148 213 149
rect 211 148 212 149
rect 210 148 211 149
rect 209 148 210 149
rect 208 148 209 149
rect 207 148 208 149
rect 206 148 207 149
rect 205 148 206 149
rect 204 148 205 149
rect 203 148 204 149
rect 202 148 203 149
rect 201 148 202 149
rect 200 148 201 149
rect 199 148 200 149
rect 198 148 199 149
rect 197 148 198 149
rect 196 148 197 149
rect 195 148 196 149
rect 194 148 195 149
rect 193 148 194 149
rect 192 148 193 149
rect 191 148 192 149
rect 190 148 191 149
rect 189 148 190 149
rect 188 148 189 149
rect 187 148 188 149
rect 186 148 187 149
rect 185 148 186 149
rect 184 148 185 149
rect 183 148 184 149
rect 182 148 183 149
rect 181 148 182 149
rect 180 148 181 149
rect 179 148 180 149
rect 178 148 179 149
rect 177 148 178 149
rect 176 148 177 149
rect 175 148 176 149
rect 174 148 175 149
rect 173 148 174 149
rect 172 148 173 149
rect 171 148 172 149
rect 170 148 171 149
rect 169 148 170 149
rect 168 148 169 149
rect 167 148 168 149
rect 166 148 167 149
rect 165 148 166 149
rect 164 148 165 149
rect 163 148 164 149
rect 162 148 163 149
rect 161 148 162 149
rect 160 148 161 149
rect 159 148 160 149
rect 158 148 159 149
rect 136 148 137 149
rect 135 148 136 149
rect 134 148 135 149
rect 133 148 134 149
rect 132 148 133 149
rect 131 148 132 149
rect 130 148 131 149
rect 129 148 130 149
rect 128 148 129 149
rect 127 148 128 149
rect 126 148 127 149
rect 125 148 126 149
rect 124 148 125 149
rect 123 148 124 149
rect 122 148 123 149
rect 121 148 122 149
rect 120 148 121 149
rect 119 148 120 149
rect 118 148 119 149
rect 117 148 118 149
rect 116 148 117 149
rect 115 148 116 149
rect 114 148 115 149
rect 113 148 114 149
rect 112 148 113 149
rect 111 148 112 149
rect 110 148 111 149
rect 109 148 110 149
rect 108 148 109 149
rect 107 148 108 149
rect 106 148 107 149
rect 105 148 106 149
rect 104 148 105 149
rect 103 148 104 149
rect 102 148 103 149
rect 101 148 102 149
rect 100 148 101 149
rect 99 148 100 149
rect 98 148 99 149
rect 97 148 98 149
rect 96 148 97 149
rect 95 148 96 149
rect 94 148 95 149
rect 93 148 94 149
rect 92 148 93 149
rect 91 148 92 149
rect 90 148 91 149
rect 89 148 90 149
rect 88 148 89 149
rect 87 148 88 149
rect 86 148 87 149
rect 85 148 86 149
rect 84 148 85 149
rect 83 148 84 149
rect 82 148 83 149
rect 81 148 82 149
rect 80 148 81 149
rect 79 148 80 149
rect 78 148 79 149
rect 77 148 78 149
rect 76 148 77 149
rect 75 148 76 149
rect 74 148 75 149
rect 73 148 74 149
rect 72 148 73 149
rect 71 148 72 149
rect 70 148 71 149
rect 69 148 70 149
rect 68 148 69 149
rect 67 148 68 149
rect 66 148 67 149
rect 65 148 66 149
rect 64 148 65 149
rect 63 148 64 149
rect 62 148 63 149
rect 61 148 62 149
rect 60 148 61 149
rect 59 148 60 149
rect 58 148 59 149
rect 57 148 58 149
rect 56 148 57 149
rect 55 148 56 149
rect 54 148 55 149
rect 53 148 54 149
rect 52 148 53 149
rect 51 148 52 149
rect 50 148 51 149
rect 49 148 50 149
rect 48 148 49 149
rect 47 148 48 149
rect 46 148 47 149
rect 45 148 46 149
rect 44 148 45 149
rect 43 148 44 149
rect 42 148 43 149
rect 30 148 31 149
rect 29 148 30 149
rect 28 148 29 149
rect 27 148 28 149
rect 26 148 27 149
rect 25 148 26 149
rect 24 148 25 149
rect 23 148 24 149
rect 22 148 23 149
rect 21 148 22 149
rect 20 148 21 149
rect 19 148 20 149
rect 18 148 19 149
rect 17 148 18 149
rect 16 148 17 149
rect 15 148 16 149
rect 482 149 483 150
rect 481 149 482 150
rect 480 149 481 150
rect 479 149 480 150
rect 478 149 479 150
rect 477 149 478 150
rect 476 149 477 150
rect 475 149 476 150
rect 474 149 475 150
rect 473 149 474 150
rect 472 149 473 150
rect 471 149 472 150
rect 470 149 471 150
rect 469 149 470 150
rect 468 149 469 150
rect 467 149 468 150
rect 466 149 467 150
rect 465 149 466 150
rect 464 149 465 150
rect 463 149 464 150
rect 462 149 463 150
rect 399 149 400 150
rect 398 149 399 150
rect 397 149 398 150
rect 320 149 321 150
rect 319 149 320 150
rect 318 149 319 150
rect 317 149 318 150
rect 316 149 317 150
rect 315 149 316 150
rect 314 149 315 150
rect 313 149 314 150
rect 312 149 313 150
rect 311 149 312 150
rect 310 149 311 150
rect 309 149 310 150
rect 308 149 309 150
rect 307 149 308 150
rect 306 149 307 150
rect 305 149 306 150
rect 304 149 305 150
rect 303 149 304 150
rect 302 149 303 150
rect 301 149 302 150
rect 300 149 301 150
rect 299 149 300 150
rect 298 149 299 150
rect 297 149 298 150
rect 296 149 297 150
rect 295 149 296 150
rect 294 149 295 150
rect 293 149 294 150
rect 292 149 293 150
rect 291 149 292 150
rect 290 149 291 150
rect 289 149 290 150
rect 288 149 289 150
rect 287 149 288 150
rect 286 149 287 150
rect 285 149 286 150
rect 284 149 285 150
rect 283 149 284 150
rect 282 149 283 150
rect 281 149 282 150
rect 280 149 281 150
rect 279 149 280 150
rect 278 149 279 150
rect 277 149 278 150
rect 276 149 277 150
rect 275 149 276 150
rect 274 149 275 150
rect 273 149 274 150
rect 272 149 273 150
rect 271 149 272 150
rect 270 149 271 150
rect 269 149 270 150
rect 268 149 269 150
rect 267 149 268 150
rect 266 149 267 150
rect 265 149 266 150
rect 264 149 265 150
rect 263 149 264 150
rect 262 149 263 150
rect 261 149 262 150
rect 260 149 261 150
rect 259 149 260 150
rect 258 149 259 150
rect 257 149 258 150
rect 256 149 257 150
rect 255 149 256 150
rect 254 149 255 150
rect 253 149 254 150
rect 252 149 253 150
rect 251 149 252 150
rect 250 149 251 150
rect 249 149 250 150
rect 248 149 249 150
rect 247 149 248 150
rect 246 149 247 150
rect 245 149 246 150
rect 244 149 245 150
rect 243 149 244 150
rect 222 149 223 150
rect 221 149 222 150
rect 220 149 221 150
rect 219 149 220 150
rect 218 149 219 150
rect 217 149 218 150
rect 216 149 217 150
rect 215 149 216 150
rect 214 149 215 150
rect 213 149 214 150
rect 212 149 213 150
rect 211 149 212 150
rect 210 149 211 150
rect 209 149 210 150
rect 208 149 209 150
rect 207 149 208 150
rect 206 149 207 150
rect 205 149 206 150
rect 204 149 205 150
rect 203 149 204 150
rect 202 149 203 150
rect 201 149 202 150
rect 200 149 201 150
rect 199 149 200 150
rect 198 149 199 150
rect 197 149 198 150
rect 196 149 197 150
rect 195 149 196 150
rect 194 149 195 150
rect 193 149 194 150
rect 192 149 193 150
rect 191 149 192 150
rect 190 149 191 150
rect 189 149 190 150
rect 188 149 189 150
rect 187 149 188 150
rect 186 149 187 150
rect 185 149 186 150
rect 184 149 185 150
rect 183 149 184 150
rect 182 149 183 150
rect 181 149 182 150
rect 180 149 181 150
rect 179 149 180 150
rect 178 149 179 150
rect 177 149 178 150
rect 176 149 177 150
rect 175 149 176 150
rect 174 149 175 150
rect 173 149 174 150
rect 172 149 173 150
rect 171 149 172 150
rect 170 149 171 150
rect 169 149 170 150
rect 168 149 169 150
rect 167 149 168 150
rect 166 149 167 150
rect 165 149 166 150
rect 164 149 165 150
rect 163 149 164 150
rect 162 149 163 150
rect 161 149 162 150
rect 160 149 161 150
rect 159 149 160 150
rect 158 149 159 150
rect 134 149 135 150
rect 133 149 134 150
rect 132 149 133 150
rect 131 149 132 150
rect 130 149 131 150
rect 129 149 130 150
rect 128 149 129 150
rect 127 149 128 150
rect 126 149 127 150
rect 125 149 126 150
rect 124 149 125 150
rect 123 149 124 150
rect 122 149 123 150
rect 121 149 122 150
rect 120 149 121 150
rect 119 149 120 150
rect 118 149 119 150
rect 117 149 118 150
rect 116 149 117 150
rect 115 149 116 150
rect 114 149 115 150
rect 113 149 114 150
rect 112 149 113 150
rect 111 149 112 150
rect 110 149 111 150
rect 109 149 110 150
rect 108 149 109 150
rect 107 149 108 150
rect 106 149 107 150
rect 105 149 106 150
rect 104 149 105 150
rect 103 149 104 150
rect 102 149 103 150
rect 101 149 102 150
rect 100 149 101 150
rect 99 149 100 150
rect 98 149 99 150
rect 97 149 98 150
rect 96 149 97 150
rect 95 149 96 150
rect 94 149 95 150
rect 93 149 94 150
rect 92 149 93 150
rect 91 149 92 150
rect 90 149 91 150
rect 89 149 90 150
rect 88 149 89 150
rect 87 149 88 150
rect 86 149 87 150
rect 85 149 86 150
rect 84 149 85 150
rect 83 149 84 150
rect 82 149 83 150
rect 81 149 82 150
rect 80 149 81 150
rect 79 149 80 150
rect 78 149 79 150
rect 77 149 78 150
rect 76 149 77 150
rect 75 149 76 150
rect 74 149 75 150
rect 73 149 74 150
rect 72 149 73 150
rect 71 149 72 150
rect 70 149 71 150
rect 69 149 70 150
rect 68 149 69 150
rect 67 149 68 150
rect 66 149 67 150
rect 65 149 66 150
rect 64 149 65 150
rect 63 149 64 150
rect 62 149 63 150
rect 61 149 62 150
rect 60 149 61 150
rect 59 149 60 150
rect 58 149 59 150
rect 57 149 58 150
rect 56 149 57 150
rect 55 149 56 150
rect 54 149 55 150
rect 53 149 54 150
rect 52 149 53 150
rect 51 149 52 150
rect 50 149 51 150
rect 49 149 50 150
rect 48 149 49 150
rect 47 149 48 150
rect 46 149 47 150
rect 45 149 46 150
rect 44 149 45 150
rect 43 149 44 150
rect 42 149 43 150
rect 31 149 32 150
rect 30 149 31 150
rect 29 149 30 150
rect 28 149 29 150
rect 27 149 28 150
rect 26 149 27 150
rect 25 149 26 150
rect 24 149 25 150
rect 23 149 24 150
rect 22 149 23 150
rect 21 149 22 150
rect 20 149 21 150
rect 19 149 20 150
rect 18 149 19 150
rect 17 149 18 150
rect 16 149 17 150
rect 15 149 16 150
rect 14 149 15 150
rect 482 150 483 151
rect 481 150 482 151
rect 480 150 481 151
rect 479 150 480 151
rect 478 150 479 151
rect 477 150 478 151
rect 476 150 477 151
rect 475 150 476 151
rect 474 150 475 151
rect 473 150 474 151
rect 472 150 473 151
rect 471 150 472 151
rect 470 150 471 151
rect 469 150 470 151
rect 468 150 469 151
rect 467 150 468 151
rect 466 150 467 151
rect 465 150 466 151
rect 464 150 465 151
rect 463 150 464 151
rect 462 150 463 151
rect 399 150 400 151
rect 398 150 399 151
rect 397 150 398 151
rect 321 150 322 151
rect 320 150 321 151
rect 319 150 320 151
rect 318 150 319 151
rect 317 150 318 151
rect 316 150 317 151
rect 315 150 316 151
rect 314 150 315 151
rect 313 150 314 151
rect 312 150 313 151
rect 311 150 312 151
rect 310 150 311 151
rect 309 150 310 151
rect 308 150 309 151
rect 307 150 308 151
rect 306 150 307 151
rect 305 150 306 151
rect 304 150 305 151
rect 303 150 304 151
rect 302 150 303 151
rect 301 150 302 151
rect 300 150 301 151
rect 299 150 300 151
rect 298 150 299 151
rect 297 150 298 151
rect 296 150 297 151
rect 295 150 296 151
rect 294 150 295 151
rect 293 150 294 151
rect 292 150 293 151
rect 291 150 292 151
rect 290 150 291 151
rect 289 150 290 151
rect 288 150 289 151
rect 287 150 288 151
rect 286 150 287 151
rect 285 150 286 151
rect 284 150 285 151
rect 283 150 284 151
rect 282 150 283 151
rect 281 150 282 151
rect 280 150 281 151
rect 279 150 280 151
rect 278 150 279 151
rect 277 150 278 151
rect 276 150 277 151
rect 275 150 276 151
rect 274 150 275 151
rect 273 150 274 151
rect 272 150 273 151
rect 271 150 272 151
rect 270 150 271 151
rect 269 150 270 151
rect 268 150 269 151
rect 267 150 268 151
rect 266 150 267 151
rect 265 150 266 151
rect 264 150 265 151
rect 263 150 264 151
rect 262 150 263 151
rect 261 150 262 151
rect 260 150 261 151
rect 259 150 260 151
rect 258 150 259 151
rect 257 150 258 151
rect 256 150 257 151
rect 255 150 256 151
rect 254 150 255 151
rect 253 150 254 151
rect 252 150 253 151
rect 251 150 252 151
rect 250 150 251 151
rect 249 150 250 151
rect 248 150 249 151
rect 247 150 248 151
rect 246 150 247 151
rect 245 150 246 151
rect 244 150 245 151
rect 243 150 244 151
rect 242 150 243 151
rect 221 150 222 151
rect 220 150 221 151
rect 219 150 220 151
rect 218 150 219 151
rect 217 150 218 151
rect 216 150 217 151
rect 215 150 216 151
rect 214 150 215 151
rect 213 150 214 151
rect 212 150 213 151
rect 211 150 212 151
rect 210 150 211 151
rect 209 150 210 151
rect 208 150 209 151
rect 207 150 208 151
rect 206 150 207 151
rect 205 150 206 151
rect 204 150 205 151
rect 203 150 204 151
rect 202 150 203 151
rect 201 150 202 151
rect 200 150 201 151
rect 199 150 200 151
rect 198 150 199 151
rect 197 150 198 151
rect 196 150 197 151
rect 195 150 196 151
rect 194 150 195 151
rect 193 150 194 151
rect 192 150 193 151
rect 191 150 192 151
rect 190 150 191 151
rect 189 150 190 151
rect 188 150 189 151
rect 187 150 188 151
rect 186 150 187 151
rect 185 150 186 151
rect 184 150 185 151
rect 183 150 184 151
rect 182 150 183 151
rect 181 150 182 151
rect 180 150 181 151
rect 179 150 180 151
rect 178 150 179 151
rect 177 150 178 151
rect 176 150 177 151
rect 175 150 176 151
rect 174 150 175 151
rect 173 150 174 151
rect 172 150 173 151
rect 171 150 172 151
rect 170 150 171 151
rect 169 150 170 151
rect 168 150 169 151
rect 167 150 168 151
rect 166 150 167 151
rect 165 150 166 151
rect 164 150 165 151
rect 163 150 164 151
rect 162 150 163 151
rect 161 150 162 151
rect 160 150 161 151
rect 159 150 160 151
rect 158 150 159 151
rect 157 150 158 151
rect 133 150 134 151
rect 132 150 133 151
rect 131 150 132 151
rect 130 150 131 151
rect 129 150 130 151
rect 128 150 129 151
rect 127 150 128 151
rect 126 150 127 151
rect 125 150 126 151
rect 124 150 125 151
rect 123 150 124 151
rect 122 150 123 151
rect 121 150 122 151
rect 120 150 121 151
rect 119 150 120 151
rect 118 150 119 151
rect 117 150 118 151
rect 116 150 117 151
rect 115 150 116 151
rect 114 150 115 151
rect 113 150 114 151
rect 112 150 113 151
rect 111 150 112 151
rect 110 150 111 151
rect 109 150 110 151
rect 108 150 109 151
rect 107 150 108 151
rect 106 150 107 151
rect 105 150 106 151
rect 104 150 105 151
rect 103 150 104 151
rect 102 150 103 151
rect 101 150 102 151
rect 100 150 101 151
rect 99 150 100 151
rect 98 150 99 151
rect 97 150 98 151
rect 96 150 97 151
rect 95 150 96 151
rect 94 150 95 151
rect 93 150 94 151
rect 92 150 93 151
rect 91 150 92 151
rect 90 150 91 151
rect 89 150 90 151
rect 88 150 89 151
rect 87 150 88 151
rect 86 150 87 151
rect 85 150 86 151
rect 84 150 85 151
rect 83 150 84 151
rect 82 150 83 151
rect 81 150 82 151
rect 80 150 81 151
rect 79 150 80 151
rect 78 150 79 151
rect 77 150 78 151
rect 76 150 77 151
rect 75 150 76 151
rect 74 150 75 151
rect 73 150 74 151
rect 72 150 73 151
rect 71 150 72 151
rect 70 150 71 151
rect 69 150 70 151
rect 68 150 69 151
rect 67 150 68 151
rect 66 150 67 151
rect 65 150 66 151
rect 64 150 65 151
rect 63 150 64 151
rect 62 150 63 151
rect 61 150 62 151
rect 60 150 61 151
rect 59 150 60 151
rect 58 150 59 151
rect 57 150 58 151
rect 56 150 57 151
rect 55 150 56 151
rect 54 150 55 151
rect 53 150 54 151
rect 52 150 53 151
rect 51 150 52 151
rect 50 150 51 151
rect 49 150 50 151
rect 48 150 49 151
rect 47 150 48 151
rect 46 150 47 151
rect 45 150 46 151
rect 44 150 45 151
rect 43 150 44 151
rect 42 150 43 151
rect 31 150 32 151
rect 30 150 31 151
rect 29 150 30 151
rect 28 150 29 151
rect 27 150 28 151
rect 26 150 27 151
rect 25 150 26 151
rect 24 150 25 151
rect 23 150 24 151
rect 22 150 23 151
rect 21 150 22 151
rect 20 150 21 151
rect 19 150 20 151
rect 18 150 19 151
rect 17 150 18 151
rect 16 150 17 151
rect 15 150 16 151
rect 14 150 15 151
rect 13 150 14 151
rect 482 151 483 152
rect 481 151 482 152
rect 480 151 481 152
rect 479 151 480 152
rect 478 151 479 152
rect 477 151 478 152
rect 476 151 477 152
rect 475 151 476 152
rect 474 151 475 152
rect 473 151 474 152
rect 472 151 473 152
rect 471 151 472 152
rect 470 151 471 152
rect 469 151 470 152
rect 468 151 469 152
rect 467 151 468 152
rect 466 151 467 152
rect 465 151 466 152
rect 464 151 465 152
rect 463 151 464 152
rect 462 151 463 152
rect 399 151 400 152
rect 398 151 399 152
rect 397 151 398 152
rect 321 151 322 152
rect 320 151 321 152
rect 319 151 320 152
rect 318 151 319 152
rect 317 151 318 152
rect 316 151 317 152
rect 315 151 316 152
rect 314 151 315 152
rect 313 151 314 152
rect 312 151 313 152
rect 311 151 312 152
rect 310 151 311 152
rect 309 151 310 152
rect 308 151 309 152
rect 307 151 308 152
rect 306 151 307 152
rect 305 151 306 152
rect 304 151 305 152
rect 303 151 304 152
rect 302 151 303 152
rect 301 151 302 152
rect 300 151 301 152
rect 299 151 300 152
rect 298 151 299 152
rect 297 151 298 152
rect 296 151 297 152
rect 295 151 296 152
rect 294 151 295 152
rect 293 151 294 152
rect 292 151 293 152
rect 291 151 292 152
rect 290 151 291 152
rect 289 151 290 152
rect 288 151 289 152
rect 287 151 288 152
rect 286 151 287 152
rect 285 151 286 152
rect 284 151 285 152
rect 283 151 284 152
rect 282 151 283 152
rect 281 151 282 152
rect 280 151 281 152
rect 279 151 280 152
rect 278 151 279 152
rect 277 151 278 152
rect 276 151 277 152
rect 275 151 276 152
rect 274 151 275 152
rect 273 151 274 152
rect 272 151 273 152
rect 271 151 272 152
rect 270 151 271 152
rect 269 151 270 152
rect 268 151 269 152
rect 267 151 268 152
rect 266 151 267 152
rect 265 151 266 152
rect 264 151 265 152
rect 263 151 264 152
rect 262 151 263 152
rect 261 151 262 152
rect 260 151 261 152
rect 259 151 260 152
rect 258 151 259 152
rect 257 151 258 152
rect 256 151 257 152
rect 255 151 256 152
rect 254 151 255 152
rect 253 151 254 152
rect 252 151 253 152
rect 251 151 252 152
rect 250 151 251 152
rect 249 151 250 152
rect 248 151 249 152
rect 247 151 248 152
rect 246 151 247 152
rect 245 151 246 152
rect 244 151 245 152
rect 243 151 244 152
rect 242 151 243 152
rect 221 151 222 152
rect 220 151 221 152
rect 219 151 220 152
rect 218 151 219 152
rect 217 151 218 152
rect 216 151 217 152
rect 215 151 216 152
rect 214 151 215 152
rect 213 151 214 152
rect 212 151 213 152
rect 211 151 212 152
rect 210 151 211 152
rect 209 151 210 152
rect 208 151 209 152
rect 207 151 208 152
rect 206 151 207 152
rect 205 151 206 152
rect 204 151 205 152
rect 203 151 204 152
rect 202 151 203 152
rect 201 151 202 152
rect 200 151 201 152
rect 199 151 200 152
rect 198 151 199 152
rect 197 151 198 152
rect 196 151 197 152
rect 195 151 196 152
rect 194 151 195 152
rect 193 151 194 152
rect 192 151 193 152
rect 191 151 192 152
rect 190 151 191 152
rect 189 151 190 152
rect 188 151 189 152
rect 187 151 188 152
rect 186 151 187 152
rect 185 151 186 152
rect 184 151 185 152
rect 183 151 184 152
rect 182 151 183 152
rect 181 151 182 152
rect 180 151 181 152
rect 179 151 180 152
rect 178 151 179 152
rect 177 151 178 152
rect 176 151 177 152
rect 175 151 176 152
rect 174 151 175 152
rect 173 151 174 152
rect 172 151 173 152
rect 171 151 172 152
rect 170 151 171 152
rect 169 151 170 152
rect 168 151 169 152
rect 167 151 168 152
rect 166 151 167 152
rect 165 151 166 152
rect 164 151 165 152
rect 163 151 164 152
rect 162 151 163 152
rect 161 151 162 152
rect 160 151 161 152
rect 159 151 160 152
rect 158 151 159 152
rect 157 151 158 152
rect 131 151 132 152
rect 130 151 131 152
rect 129 151 130 152
rect 128 151 129 152
rect 127 151 128 152
rect 126 151 127 152
rect 125 151 126 152
rect 124 151 125 152
rect 123 151 124 152
rect 122 151 123 152
rect 121 151 122 152
rect 120 151 121 152
rect 119 151 120 152
rect 118 151 119 152
rect 117 151 118 152
rect 116 151 117 152
rect 115 151 116 152
rect 114 151 115 152
rect 113 151 114 152
rect 112 151 113 152
rect 111 151 112 152
rect 110 151 111 152
rect 109 151 110 152
rect 108 151 109 152
rect 107 151 108 152
rect 106 151 107 152
rect 105 151 106 152
rect 104 151 105 152
rect 103 151 104 152
rect 102 151 103 152
rect 101 151 102 152
rect 100 151 101 152
rect 99 151 100 152
rect 98 151 99 152
rect 97 151 98 152
rect 96 151 97 152
rect 95 151 96 152
rect 94 151 95 152
rect 93 151 94 152
rect 92 151 93 152
rect 91 151 92 152
rect 90 151 91 152
rect 89 151 90 152
rect 88 151 89 152
rect 87 151 88 152
rect 86 151 87 152
rect 85 151 86 152
rect 84 151 85 152
rect 83 151 84 152
rect 82 151 83 152
rect 81 151 82 152
rect 80 151 81 152
rect 79 151 80 152
rect 78 151 79 152
rect 77 151 78 152
rect 76 151 77 152
rect 75 151 76 152
rect 74 151 75 152
rect 73 151 74 152
rect 72 151 73 152
rect 71 151 72 152
rect 70 151 71 152
rect 69 151 70 152
rect 68 151 69 152
rect 67 151 68 152
rect 66 151 67 152
rect 65 151 66 152
rect 64 151 65 152
rect 63 151 64 152
rect 62 151 63 152
rect 61 151 62 152
rect 60 151 61 152
rect 59 151 60 152
rect 58 151 59 152
rect 57 151 58 152
rect 56 151 57 152
rect 55 151 56 152
rect 54 151 55 152
rect 53 151 54 152
rect 52 151 53 152
rect 51 151 52 152
rect 50 151 51 152
rect 49 151 50 152
rect 48 151 49 152
rect 47 151 48 152
rect 46 151 47 152
rect 45 151 46 152
rect 44 151 45 152
rect 43 151 44 152
rect 42 151 43 152
rect 41 151 42 152
rect 31 151 32 152
rect 30 151 31 152
rect 29 151 30 152
rect 28 151 29 152
rect 27 151 28 152
rect 26 151 27 152
rect 25 151 26 152
rect 24 151 25 152
rect 23 151 24 152
rect 22 151 23 152
rect 21 151 22 152
rect 20 151 21 152
rect 19 151 20 152
rect 18 151 19 152
rect 17 151 18 152
rect 16 151 17 152
rect 15 151 16 152
rect 14 151 15 152
rect 13 151 14 152
rect 482 152 483 153
rect 462 152 463 153
rect 322 152 323 153
rect 321 152 322 153
rect 320 152 321 153
rect 319 152 320 153
rect 318 152 319 153
rect 317 152 318 153
rect 316 152 317 153
rect 315 152 316 153
rect 314 152 315 153
rect 313 152 314 153
rect 312 152 313 153
rect 311 152 312 153
rect 310 152 311 153
rect 309 152 310 153
rect 308 152 309 153
rect 307 152 308 153
rect 306 152 307 153
rect 305 152 306 153
rect 304 152 305 153
rect 303 152 304 153
rect 302 152 303 153
rect 301 152 302 153
rect 300 152 301 153
rect 299 152 300 153
rect 298 152 299 153
rect 297 152 298 153
rect 296 152 297 153
rect 295 152 296 153
rect 294 152 295 153
rect 293 152 294 153
rect 292 152 293 153
rect 291 152 292 153
rect 290 152 291 153
rect 289 152 290 153
rect 288 152 289 153
rect 287 152 288 153
rect 286 152 287 153
rect 285 152 286 153
rect 284 152 285 153
rect 283 152 284 153
rect 282 152 283 153
rect 281 152 282 153
rect 280 152 281 153
rect 279 152 280 153
rect 278 152 279 153
rect 277 152 278 153
rect 276 152 277 153
rect 275 152 276 153
rect 274 152 275 153
rect 273 152 274 153
rect 272 152 273 153
rect 271 152 272 153
rect 270 152 271 153
rect 269 152 270 153
rect 268 152 269 153
rect 267 152 268 153
rect 266 152 267 153
rect 265 152 266 153
rect 264 152 265 153
rect 263 152 264 153
rect 262 152 263 153
rect 261 152 262 153
rect 260 152 261 153
rect 259 152 260 153
rect 258 152 259 153
rect 257 152 258 153
rect 256 152 257 153
rect 255 152 256 153
rect 254 152 255 153
rect 253 152 254 153
rect 252 152 253 153
rect 251 152 252 153
rect 250 152 251 153
rect 249 152 250 153
rect 248 152 249 153
rect 247 152 248 153
rect 246 152 247 153
rect 245 152 246 153
rect 244 152 245 153
rect 243 152 244 153
rect 242 152 243 153
rect 241 152 242 153
rect 220 152 221 153
rect 219 152 220 153
rect 218 152 219 153
rect 217 152 218 153
rect 216 152 217 153
rect 215 152 216 153
rect 214 152 215 153
rect 213 152 214 153
rect 212 152 213 153
rect 211 152 212 153
rect 210 152 211 153
rect 209 152 210 153
rect 208 152 209 153
rect 207 152 208 153
rect 206 152 207 153
rect 205 152 206 153
rect 204 152 205 153
rect 203 152 204 153
rect 202 152 203 153
rect 201 152 202 153
rect 200 152 201 153
rect 199 152 200 153
rect 198 152 199 153
rect 197 152 198 153
rect 196 152 197 153
rect 195 152 196 153
rect 194 152 195 153
rect 193 152 194 153
rect 192 152 193 153
rect 191 152 192 153
rect 190 152 191 153
rect 189 152 190 153
rect 188 152 189 153
rect 187 152 188 153
rect 186 152 187 153
rect 185 152 186 153
rect 184 152 185 153
rect 183 152 184 153
rect 182 152 183 153
rect 181 152 182 153
rect 180 152 181 153
rect 179 152 180 153
rect 178 152 179 153
rect 177 152 178 153
rect 176 152 177 153
rect 175 152 176 153
rect 174 152 175 153
rect 173 152 174 153
rect 172 152 173 153
rect 171 152 172 153
rect 170 152 171 153
rect 169 152 170 153
rect 168 152 169 153
rect 167 152 168 153
rect 166 152 167 153
rect 165 152 166 153
rect 164 152 165 153
rect 163 152 164 153
rect 162 152 163 153
rect 161 152 162 153
rect 160 152 161 153
rect 159 152 160 153
rect 158 152 159 153
rect 157 152 158 153
rect 156 152 157 153
rect 130 152 131 153
rect 129 152 130 153
rect 128 152 129 153
rect 127 152 128 153
rect 126 152 127 153
rect 125 152 126 153
rect 124 152 125 153
rect 123 152 124 153
rect 122 152 123 153
rect 121 152 122 153
rect 120 152 121 153
rect 119 152 120 153
rect 118 152 119 153
rect 117 152 118 153
rect 116 152 117 153
rect 115 152 116 153
rect 114 152 115 153
rect 113 152 114 153
rect 112 152 113 153
rect 111 152 112 153
rect 110 152 111 153
rect 109 152 110 153
rect 108 152 109 153
rect 107 152 108 153
rect 106 152 107 153
rect 105 152 106 153
rect 104 152 105 153
rect 103 152 104 153
rect 102 152 103 153
rect 101 152 102 153
rect 100 152 101 153
rect 99 152 100 153
rect 98 152 99 153
rect 97 152 98 153
rect 96 152 97 153
rect 95 152 96 153
rect 94 152 95 153
rect 93 152 94 153
rect 92 152 93 153
rect 91 152 92 153
rect 90 152 91 153
rect 89 152 90 153
rect 88 152 89 153
rect 87 152 88 153
rect 86 152 87 153
rect 85 152 86 153
rect 84 152 85 153
rect 83 152 84 153
rect 82 152 83 153
rect 81 152 82 153
rect 80 152 81 153
rect 79 152 80 153
rect 78 152 79 153
rect 77 152 78 153
rect 76 152 77 153
rect 75 152 76 153
rect 74 152 75 153
rect 73 152 74 153
rect 72 152 73 153
rect 71 152 72 153
rect 70 152 71 153
rect 69 152 70 153
rect 68 152 69 153
rect 67 152 68 153
rect 66 152 67 153
rect 65 152 66 153
rect 64 152 65 153
rect 63 152 64 153
rect 62 152 63 153
rect 61 152 62 153
rect 60 152 61 153
rect 59 152 60 153
rect 58 152 59 153
rect 57 152 58 153
rect 56 152 57 153
rect 55 152 56 153
rect 54 152 55 153
rect 53 152 54 153
rect 52 152 53 153
rect 51 152 52 153
rect 50 152 51 153
rect 49 152 50 153
rect 48 152 49 153
rect 47 152 48 153
rect 46 152 47 153
rect 45 152 46 153
rect 44 152 45 153
rect 43 152 44 153
rect 42 152 43 153
rect 41 152 42 153
rect 31 152 32 153
rect 30 152 31 153
rect 29 152 30 153
rect 28 152 29 153
rect 27 152 28 153
rect 26 152 27 153
rect 25 152 26 153
rect 24 152 25 153
rect 23 152 24 153
rect 22 152 23 153
rect 21 152 22 153
rect 20 152 21 153
rect 19 152 20 153
rect 18 152 19 153
rect 17 152 18 153
rect 16 152 17 153
rect 15 152 16 153
rect 14 152 15 153
rect 13 152 14 153
rect 12 152 13 153
rect 482 153 483 154
rect 462 153 463 154
rect 323 153 324 154
rect 322 153 323 154
rect 321 153 322 154
rect 320 153 321 154
rect 319 153 320 154
rect 318 153 319 154
rect 317 153 318 154
rect 316 153 317 154
rect 315 153 316 154
rect 314 153 315 154
rect 313 153 314 154
rect 312 153 313 154
rect 311 153 312 154
rect 310 153 311 154
rect 309 153 310 154
rect 308 153 309 154
rect 307 153 308 154
rect 306 153 307 154
rect 305 153 306 154
rect 304 153 305 154
rect 303 153 304 154
rect 302 153 303 154
rect 301 153 302 154
rect 300 153 301 154
rect 299 153 300 154
rect 298 153 299 154
rect 297 153 298 154
rect 296 153 297 154
rect 295 153 296 154
rect 294 153 295 154
rect 293 153 294 154
rect 292 153 293 154
rect 291 153 292 154
rect 290 153 291 154
rect 289 153 290 154
rect 288 153 289 154
rect 287 153 288 154
rect 286 153 287 154
rect 285 153 286 154
rect 284 153 285 154
rect 283 153 284 154
rect 282 153 283 154
rect 281 153 282 154
rect 280 153 281 154
rect 279 153 280 154
rect 278 153 279 154
rect 277 153 278 154
rect 276 153 277 154
rect 275 153 276 154
rect 274 153 275 154
rect 273 153 274 154
rect 272 153 273 154
rect 271 153 272 154
rect 270 153 271 154
rect 269 153 270 154
rect 268 153 269 154
rect 267 153 268 154
rect 266 153 267 154
rect 265 153 266 154
rect 264 153 265 154
rect 263 153 264 154
rect 262 153 263 154
rect 261 153 262 154
rect 260 153 261 154
rect 259 153 260 154
rect 258 153 259 154
rect 257 153 258 154
rect 256 153 257 154
rect 255 153 256 154
rect 254 153 255 154
rect 253 153 254 154
rect 252 153 253 154
rect 251 153 252 154
rect 250 153 251 154
rect 249 153 250 154
rect 248 153 249 154
rect 247 153 248 154
rect 246 153 247 154
rect 245 153 246 154
rect 244 153 245 154
rect 243 153 244 154
rect 242 153 243 154
rect 241 153 242 154
rect 240 153 241 154
rect 220 153 221 154
rect 219 153 220 154
rect 218 153 219 154
rect 217 153 218 154
rect 216 153 217 154
rect 215 153 216 154
rect 214 153 215 154
rect 213 153 214 154
rect 212 153 213 154
rect 211 153 212 154
rect 210 153 211 154
rect 209 153 210 154
rect 208 153 209 154
rect 207 153 208 154
rect 206 153 207 154
rect 205 153 206 154
rect 204 153 205 154
rect 203 153 204 154
rect 202 153 203 154
rect 201 153 202 154
rect 200 153 201 154
rect 199 153 200 154
rect 198 153 199 154
rect 197 153 198 154
rect 196 153 197 154
rect 195 153 196 154
rect 194 153 195 154
rect 193 153 194 154
rect 192 153 193 154
rect 191 153 192 154
rect 190 153 191 154
rect 189 153 190 154
rect 188 153 189 154
rect 187 153 188 154
rect 186 153 187 154
rect 185 153 186 154
rect 184 153 185 154
rect 183 153 184 154
rect 182 153 183 154
rect 181 153 182 154
rect 180 153 181 154
rect 179 153 180 154
rect 178 153 179 154
rect 177 153 178 154
rect 176 153 177 154
rect 175 153 176 154
rect 174 153 175 154
rect 173 153 174 154
rect 172 153 173 154
rect 171 153 172 154
rect 170 153 171 154
rect 169 153 170 154
rect 168 153 169 154
rect 167 153 168 154
rect 166 153 167 154
rect 165 153 166 154
rect 164 153 165 154
rect 163 153 164 154
rect 162 153 163 154
rect 161 153 162 154
rect 160 153 161 154
rect 159 153 160 154
rect 158 153 159 154
rect 157 153 158 154
rect 156 153 157 154
rect 155 153 156 154
rect 128 153 129 154
rect 127 153 128 154
rect 126 153 127 154
rect 125 153 126 154
rect 124 153 125 154
rect 123 153 124 154
rect 122 153 123 154
rect 121 153 122 154
rect 120 153 121 154
rect 119 153 120 154
rect 118 153 119 154
rect 117 153 118 154
rect 116 153 117 154
rect 115 153 116 154
rect 114 153 115 154
rect 113 153 114 154
rect 112 153 113 154
rect 111 153 112 154
rect 110 153 111 154
rect 109 153 110 154
rect 108 153 109 154
rect 107 153 108 154
rect 106 153 107 154
rect 105 153 106 154
rect 104 153 105 154
rect 103 153 104 154
rect 102 153 103 154
rect 101 153 102 154
rect 100 153 101 154
rect 99 153 100 154
rect 98 153 99 154
rect 97 153 98 154
rect 96 153 97 154
rect 95 153 96 154
rect 94 153 95 154
rect 93 153 94 154
rect 92 153 93 154
rect 91 153 92 154
rect 90 153 91 154
rect 89 153 90 154
rect 88 153 89 154
rect 87 153 88 154
rect 86 153 87 154
rect 85 153 86 154
rect 84 153 85 154
rect 83 153 84 154
rect 82 153 83 154
rect 81 153 82 154
rect 80 153 81 154
rect 79 153 80 154
rect 78 153 79 154
rect 77 153 78 154
rect 76 153 77 154
rect 75 153 76 154
rect 74 153 75 154
rect 73 153 74 154
rect 72 153 73 154
rect 71 153 72 154
rect 70 153 71 154
rect 69 153 70 154
rect 68 153 69 154
rect 67 153 68 154
rect 66 153 67 154
rect 65 153 66 154
rect 64 153 65 154
rect 63 153 64 154
rect 62 153 63 154
rect 61 153 62 154
rect 60 153 61 154
rect 59 153 60 154
rect 58 153 59 154
rect 57 153 58 154
rect 56 153 57 154
rect 55 153 56 154
rect 54 153 55 154
rect 53 153 54 154
rect 52 153 53 154
rect 51 153 52 154
rect 50 153 51 154
rect 49 153 50 154
rect 48 153 49 154
rect 47 153 48 154
rect 46 153 47 154
rect 45 153 46 154
rect 44 153 45 154
rect 43 153 44 154
rect 42 153 43 154
rect 41 153 42 154
rect 40 153 41 154
rect 31 153 32 154
rect 30 153 31 154
rect 29 153 30 154
rect 28 153 29 154
rect 27 153 28 154
rect 26 153 27 154
rect 25 153 26 154
rect 24 153 25 154
rect 23 153 24 154
rect 22 153 23 154
rect 21 153 22 154
rect 20 153 21 154
rect 19 153 20 154
rect 18 153 19 154
rect 17 153 18 154
rect 16 153 17 154
rect 15 153 16 154
rect 14 153 15 154
rect 13 153 14 154
rect 12 153 13 154
rect 11 153 12 154
rect 324 154 325 155
rect 323 154 324 155
rect 322 154 323 155
rect 321 154 322 155
rect 320 154 321 155
rect 319 154 320 155
rect 318 154 319 155
rect 317 154 318 155
rect 316 154 317 155
rect 315 154 316 155
rect 314 154 315 155
rect 313 154 314 155
rect 312 154 313 155
rect 311 154 312 155
rect 310 154 311 155
rect 309 154 310 155
rect 308 154 309 155
rect 307 154 308 155
rect 306 154 307 155
rect 305 154 306 155
rect 304 154 305 155
rect 303 154 304 155
rect 302 154 303 155
rect 301 154 302 155
rect 300 154 301 155
rect 299 154 300 155
rect 298 154 299 155
rect 297 154 298 155
rect 296 154 297 155
rect 295 154 296 155
rect 294 154 295 155
rect 293 154 294 155
rect 292 154 293 155
rect 291 154 292 155
rect 290 154 291 155
rect 289 154 290 155
rect 288 154 289 155
rect 287 154 288 155
rect 286 154 287 155
rect 285 154 286 155
rect 284 154 285 155
rect 283 154 284 155
rect 282 154 283 155
rect 281 154 282 155
rect 280 154 281 155
rect 279 154 280 155
rect 278 154 279 155
rect 277 154 278 155
rect 276 154 277 155
rect 275 154 276 155
rect 274 154 275 155
rect 273 154 274 155
rect 272 154 273 155
rect 271 154 272 155
rect 270 154 271 155
rect 269 154 270 155
rect 268 154 269 155
rect 267 154 268 155
rect 266 154 267 155
rect 265 154 266 155
rect 264 154 265 155
rect 263 154 264 155
rect 262 154 263 155
rect 261 154 262 155
rect 260 154 261 155
rect 259 154 260 155
rect 258 154 259 155
rect 257 154 258 155
rect 256 154 257 155
rect 255 154 256 155
rect 254 154 255 155
rect 253 154 254 155
rect 252 154 253 155
rect 251 154 252 155
rect 250 154 251 155
rect 249 154 250 155
rect 248 154 249 155
rect 247 154 248 155
rect 246 154 247 155
rect 245 154 246 155
rect 244 154 245 155
rect 243 154 244 155
rect 242 154 243 155
rect 241 154 242 155
rect 240 154 241 155
rect 220 154 221 155
rect 219 154 220 155
rect 218 154 219 155
rect 217 154 218 155
rect 216 154 217 155
rect 215 154 216 155
rect 214 154 215 155
rect 213 154 214 155
rect 212 154 213 155
rect 211 154 212 155
rect 210 154 211 155
rect 209 154 210 155
rect 208 154 209 155
rect 207 154 208 155
rect 206 154 207 155
rect 205 154 206 155
rect 204 154 205 155
rect 203 154 204 155
rect 202 154 203 155
rect 201 154 202 155
rect 200 154 201 155
rect 199 154 200 155
rect 198 154 199 155
rect 197 154 198 155
rect 196 154 197 155
rect 195 154 196 155
rect 194 154 195 155
rect 193 154 194 155
rect 192 154 193 155
rect 191 154 192 155
rect 190 154 191 155
rect 189 154 190 155
rect 188 154 189 155
rect 187 154 188 155
rect 186 154 187 155
rect 185 154 186 155
rect 184 154 185 155
rect 183 154 184 155
rect 182 154 183 155
rect 181 154 182 155
rect 180 154 181 155
rect 179 154 180 155
rect 178 154 179 155
rect 177 154 178 155
rect 176 154 177 155
rect 175 154 176 155
rect 174 154 175 155
rect 173 154 174 155
rect 172 154 173 155
rect 171 154 172 155
rect 170 154 171 155
rect 169 154 170 155
rect 168 154 169 155
rect 167 154 168 155
rect 166 154 167 155
rect 165 154 166 155
rect 164 154 165 155
rect 163 154 164 155
rect 162 154 163 155
rect 161 154 162 155
rect 160 154 161 155
rect 159 154 160 155
rect 158 154 159 155
rect 157 154 158 155
rect 156 154 157 155
rect 155 154 156 155
rect 154 154 155 155
rect 126 154 127 155
rect 125 154 126 155
rect 124 154 125 155
rect 123 154 124 155
rect 122 154 123 155
rect 121 154 122 155
rect 120 154 121 155
rect 119 154 120 155
rect 118 154 119 155
rect 117 154 118 155
rect 116 154 117 155
rect 115 154 116 155
rect 114 154 115 155
rect 113 154 114 155
rect 112 154 113 155
rect 111 154 112 155
rect 110 154 111 155
rect 109 154 110 155
rect 108 154 109 155
rect 107 154 108 155
rect 106 154 107 155
rect 105 154 106 155
rect 104 154 105 155
rect 103 154 104 155
rect 102 154 103 155
rect 101 154 102 155
rect 100 154 101 155
rect 99 154 100 155
rect 98 154 99 155
rect 97 154 98 155
rect 96 154 97 155
rect 95 154 96 155
rect 94 154 95 155
rect 93 154 94 155
rect 92 154 93 155
rect 91 154 92 155
rect 90 154 91 155
rect 89 154 90 155
rect 88 154 89 155
rect 87 154 88 155
rect 86 154 87 155
rect 85 154 86 155
rect 84 154 85 155
rect 83 154 84 155
rect 82 154 83 155
rect 81 154 82 155
rect 80 154 81 155
rect 79 154 80 155
rect 78 154 79 155
rect 77 154 78 155
rect 76 154 77 155
rect 75 154 76 155
rect 74 154 75 155
rect 73 154 74 155
rect 72 154 73 155
rect 71 154 72 155
rect 70 154 71 155
rect 69 154 70 155
rect 68 154 69 155
rect 67 154 68 155
rect 66 154 67 155
rect 65 154 66 155
rect 64 154 65 155
rect 63 154 64 155
rect 62 154 63 155
rect 61 154 62 155
rect 60 154 61 155
rect 59 154 60 155
rect 58 154 59 155
rect 57 154 58 155
rect 56 154 57 155
rect 55 154 56 155
rect 54 154 55 155
rect 53 154 54 155
rect 52 154 53 155
rect 51 154 52 155
rect 50 154 51 155
rect 49 154 50 155
rect 48 154 49 155
rect 47 154 48 155
rect 46 154 47 155
rect 45 154 46 155
rect 44 154 45 155
rect 43 154 44 155
rect 42 154 43 155
rect 41 154 42 155
rect 40 154 41 155
rect 30 154 31 155
rect 29 154 30 155
rect 28 154 29 155
rect 27 154 28 155
rect 26 154 27 155
rect 25 154 26 155
rect 24 154 25 155
rect 23 154 24 155
rect 22 154 23 155
rect 21 154 22 155
rect 20 154 21 155
rect 19 154 20 155
rect 18 154 19 155
rect 17 154 18 155
rect 16 154 17 155
rect 15 154 16 155
rect 14 154 15 155
rect 13 154 14 155
rect 12 154 13 155
rect 11 154 12 155
rect 325 155 326 156
rect 324 155 325 156
rect 323 155 324 156
rect 322 155 323 156
rect 321 155 322 156
rect 320 155 321 156
rect 319 155 320 156
rect 318 155 319 156
rect 317 155 318 156
rect 316 155 317 156
rect 315 155 316 156
rect 314 155 315 156
rect 313 155 314 156
rect 312 155 313 156
rect 311 155 312 156
rect 310 155 311 156
rect 309 155 310 156
rect 308 155 309 156
rect 307 155 308 156
rect 306 155 307 156
rect 305 155 306 156
rect 304 155 305 156
rect 303 155 304 156
rect 302 155 303 156
rect 301 155 302 156
rect 300 155 301 156
rect 299 155 300 156
rect 298 155 299 156
rect 297 155 298 156
rect 296 155 297 156
rect 295 155 296 156
rect 294 155 295 156
rect 293 155 294 156
rect 292 155 293 156
rect 291 155 292 156
rect 290 155 291 156
rect 289 155 290 156
rect 288 155 289 156
rect 287 155 288 156
rect 286 155 287 156
rect 285 155 286 156
rect 284 155 285 156
rect 283 155 284 156
rect 282 155 283 156
rect 281 155 282 156
rect 280 155 281 156
rect 279 155 280 156
rect 278 155 279 156
rect 277 155 278 156
rect 276 155 277 156
rect 275 155 276 156
rect 274 155 275 156
rect 273 155 274 156
rect 272 155 273 156
rect 271 155 272 156
rect 270 155 271 156
rect 269 155 270 156
rect 268 155 269 156
rect 267 155 268 156
rect 266 155 267 156
rect 265 155 266 156
rect 264 155 265 156
rect 263 155 264 156
rect 262 155 263 156
rect 261 155 262 156
rect 260 155 261 156
rect 259 155 260 156
rect 258 155 259 156
rect 257 155 258 156
rect 256 155 257 156
rect 255 155 256 156
rect 254 155 255 156
rect 253 155 254 156
rect 252 155 253 156
rect 251 155 252 156
rect 250 155 251 156
rect 249 155 250 156
rect 248 155 249 156
rect 247 155 248 156
rect 246 155 247 156
rect 245 155 246 156
rect 244 155 245 156
rect 243 155 244 156
rect 242 155 243 156
rect 241 155 242 156
rect 240 155 241 156
rect 239 155 240 156
rect 219 155 220 156
rect 218 155 219 156
rect 217 155 218 156
rect 216 155 217 156
rect 215 155 216 156
rect 214 155 215 156
rect 213 155 214 156
rect 212 155 213 156
rect 211 155 212 156
rect 210 155 211 156
rect 209 155 210 156
rect 208 155 209 156
rect 207 155 208 156
rect 206 155 207 156
rect 205 155 206 156
rect 204 155 205 156
rect 203 155 204 156
rect 202 155 203 156
rect 201 155 202 156
rect 200 155 201 156
rect 199 155 200 156
rect 198 155 199 156
rect 197 155 198 156
rect 196 155 197 156
rect 195 155 196 156
rect 194 155 195 156
rect 193 155 194 156
rect 192 155 193 156
rect 191 155 192 156
rect 190 155 191 156
rect 189 155 190 156
rect 188 155 189 156
rect 187 155 188 156
rect 186 155 187 156
rect 185 155 186 156
rect 184 155 185 156
rect 183 155 184 156
rect 182 155 183 156
rect 181 155 182 156
rect 180 155 181 156
rect 179 155 180 156
rect 178 155 179 156
rect 177 155 178 156
rect 176 155 177 156
rect 175 155 176 156
rect 174 155 175 156
rect 173 155 174 156
rect 172 155 173 156
rect 171 155 172 156
rect 170 155 171 156
rect 169 155 170 156
rect 168 155 169 156
rect 167 155 168 156
rect 166 155 167 156
rect 165 155 166 156
rect 164 155 165 156
rect 163 155 164 156
rect 162 155 163 156
rect 161 155 162 156
rect 160 155 161 156
rect 159 155 160 156
rect 158 155 159 156
rect 157 155 158 156
rect 156 155 157 156
rect 155 155 156 156
rect 154 155 155 156
rect 125 155 126 156
rect 124 155 125 156
rect 123 155 124 156
rect 122 155 123 156
rect 121 155 122 156
rect 120 155 121 156
rect 119 155 120 156
rect 118 155 119 156
rect 117 155 118 156
rect 116 155 117 156
rect 115 155 116 156
rect 114 155 115 156
rect 113 155 114 156
rect 112 155 113 156
rect 111 155 112 156
rect 110 155 111 156
rect 109 155 110 156
rect 108 155 109 156
rect 107 155 108 156
rect 106 155 107 156
rect 105 155 106 156
rect 104 155 105 156
rect 103 155 104 156
rect 102 155 103 156
rect 101 155 102 156
rect 100 155 101 156
rect 99 155 100 156
rect 98 155 99 156
rect 97 155 98 156
rect 96 155 97 156
rect 95 155 96 156
rect 94 155 95 156
rect 93 155 94 156
rect 92 155 93 156
rect 91 155 92 156
rect 90 155 91 156
rect 89 155 90 156
rect 88 155 89 156
rect 87 155 88 156
rect 86 155 87 156
rect 85 155 86 156
rect 84 155 85 156
rect 83 155 84 156
rect 82 155 83 156
rect 81 155 82 156
rect 80 155 81 156
rect 79 155 80 156
rect 78 155 79 156
rect 77 155 78 156
rect 76 155 77 156
rect 75 155 76 156
rect 74 155 75 156
rect 73 155 74 156
rect 72 155 73 156
rect 71 155 72 156
rect 70 155 71 156
rect 69 155 70 156
rect 68 155 69 156
rect 67 155 68 156
rect 66 155 67 156
rect 65 155 66 156
rect 64 155 65 156
rect 63 155 64 156
rect 62 155 63 156
rect 61 155 62 156
rect 60 155 61 156
rect 59 155 60 156
rect 58 155 59 156
rect 57 155 58 156
rect 56 155 57 156
rect 55 155 56 156
rect 54 155 55 156
rect 53 155 54 156
rect 52 155 53 156
rect 51 155 52 156
rect 50 155 51 156
rect 49 155 50 156
rect 48 155 49 156
rect 47 155 48 156
rect 46 155 47 156
rect 45 155 46 156
rect 44 155 45 156
rect 43 155 44 156
rect 42 155 43 156
rect 41 155 42 156
rect 40 155 41 156
rect 39 155 40 156
rect 30 155 31 156
rect 29 155 30 156
rect 28 155 29 156
rect 27 155 28 156
rect 26 155 27 156
rect 25 155 26 156
rect 24 155 25 156
rect 23 155 24 156
rect 22 155 23 156
rect 21 155 22 156
rect 20 155 21 156
rect 19 155 20 156
rect 18 155 19 156
rect 17 155 18 156
rect 16 155 17 156
rect 15 155 16 156
rect 14 155 15 156
rect 13 155 14 156
rect 12 155 13 156
rect 11 155 12 156
rect 10 155 11 156
rect 398 156 399 157
rect 397 156 398 157
rect 325 156 326 157
rect 324 156 325 157
rect 323 156 324 157
rect 322 156 323 157
rect 321 156 322 157
rect 320 156 321 157
rect 319 156 320 157
rect 318 156 319 157
rect 317 156 318 157
rect 316 156 317 157
rect 315 156 316 157
rect 314 156 315 157
rect 313 156 314 157
rect 312 156 313 157
rect 311 156 312 157
rect 310 156 311 157
rect 309 156 310 157
rect 308 156 309 157
rect 307 156 308 157
rect 306 156 307 157
rect 305 156 306 157
rect 304 156 305 157
rect 303 156 304 157
rect 302 156 303 157
rect 301 156 302 157
rect 300 156 301 157
rect 299 156 300 157
rect 298 156 299 157
rect 297 156 298 157
rect 296 156 297 157
rect 295 156 296 157
rect 294 156 295 157
rect 293 156 294 157
rect 292 156 293 157
rect 291 156 292 157
rect 290 156 291 157
rect 289 156 290 157
rect 288 156 289 157
rect 287 156 288 157
rect 286 156 287 157
rect 285 156 286 157
rect 284 156 285 157
rect 283 156 284 157
rect 282 156 283 157
rect 281 156 282 157
rect 280 156 281 157
rect 279 156 280 157
rect 278 156 279 157
rect 277 156 278 157
rect 276 156 277 157
rect 275 156 276 157
rect 274 156 275 157
rect 273 156 274 157
rect 272 156 273 157
rect 271 156 272 157
rect 270 156 271 157
rect 269 156 270 157
rect 268 156 269 157
rect 267 156 268 157
rect 266 156 267 157
rect 265 156 266 157
rect 264 156 265 157
rect 263 156 264 157
rect 262 156 263 157
rect 261 156 262 157
rect 260 156 261 157
rect 259 156 260 157
rect 258 156 259 157
rect 257 156 258 157
rect 256 156 257 157
rect 255 156 256 157
rect 254 156 255 157
rect 253 156 254 157
rect 252 156 253 157
rect 251 156 252 157
rect 250 156 251 157
rect 249 156 250 157
rect 248 156 249 157
rect 247 156 248 157
rect 246 156 247 157
rect 245 156 246 157
rect 244 156 245 157
rect 243 156 244 157
rect 242 156 243 157
rect 241 156 242 157
rect 240 156 241 157
rect 239 156 240 157
rect 238 156 239 157
rect 219 156 220 157
rect 218 156 219 157
rect 217 156 218 157
rect 216 156 217 157
rect 215 156 216 157
rect 214 156 215 157
rect 213 156 214 157
rect 212 156 213 157
rect 211 156 212 157
rect 210 156 211 157
rect 209 156 210 157
rect 208 156 209 157
rect 207 156 208 157
rect 206 156 207 157
rect 205 156 206 157
rect 204 156 205 157
rect 203 156 204 157
rect 202 156 203 157
rect 201 156 202 157
rect 200 156 201 157
rect 199 156 200 157
rect 198 156 199 157
rect 197 156 198 157
rect 196 156 197 157
rect 195 156 196 157
rect 194 156 195 157
rect 193 156 194 157
rect 192 156 193 157
rect 191 156 192 157
rect 190 156 191 157
rect 189 156 190 157
rect 188 156 189 157
rect 187 156 188 157
rect 186 156 187 157
rect 185 156 186 157
rect 184 156 185 157
rect 183 156 184 157
rect 182 156 183 157
rect 181 156 182 157
rect 180 156 181 157
rect 179 156 180 157
rect 178 156 179 157
rect 177 156 178 157
rect 176 156 177 157
rect 175 156 176 157
rect 174 156 175 157
rect 173 156 174 157
rect 172 156 173 157
rect 171 156 172 157
rect 170 156 171 157
rect 169 156 170 157
rect 168 156 169 157
rect 167 156 168 157
rect 166 156 167 157
rect 165 156 166 157
rect 164 156 165 157
rect 163 156 164 157
rect 162 156 163 157
rect 161 156 162 157
rect 160 156 161 157
rect 159 156 160 157
rect 158 156 159 157
rect 157 156 158 157
rect 156 156 157 157
rect 155 156 156 157
rect 154 156 155 157
rect 153 156 154 157
rect 123 156 124 157
rect 122 156 123 157
rect 121 156 122 157
rect 120 156 121 157
rect 119 156 120 157
rect 118 156 119 157
rect 117 156 118 157
rect 116 156 117 157
rect 115 156 116 157
rect 114 156 115 157
rect 113 156 114 157
rect 112 156 113 157
rect 111 156 112 157
rect 110 156 111 157
rect 109 156 110 157
rect 108 156 109 157
rect 107 156 108 157
rect 106 156 107 157
rect 105 156 106 157
rect 104 156 105 157
rect 103 156 104 157
rect 102 156 103 157
rect 101 156 102 157
rect 100 156 101 157
rect 99 156 100 157
rect 98 156 99 157
rect 97 156 98 157
rect 96 156 97 157
rect 95 156 96 157
rect 94 156 95 157
rect 93 156 94 157
rect 92 156 93 157
rect 91 156 92 157
rect 90 156 91 157
rect 89 156 90 157
rect 88 156 89 157
rect 87 156 88 157
rect 86 156 87 157
rect 85 156 86 157
rect 84 156 85 157
rect 83 156 84 157
rect 82 156 83 157
rect 81 156 82 157
rect 80 156 81 157
rect 79 156 80 157
rect 78 156 79 157
rect 77 156 78 157
rect 76 156 77 157
rect 75 156 76 157
rect 74 156 75 157
rect 73 156 74 157
rect 72 156 73 157
rect 71 156 72 157
rect 70 156 71 157
rect 69 156 70 157
rect 68 156 69 157
rect 67 156 68 157
rect 66 156 67 157
rect 65 156 66 157
rect 64 156 65 157
rect 63 156 64 157
rect 62 156 63 157
rect 61 156 62 157
rect 60 156 61 157
rect 59 156 60 157
rect 58 156 59 157
rect 57 156 58 157
rect 56 156 57 157
rect 55 156 56 157
rect 54 156 55 157
rect 53 156 54 157
rect 52 156 53 157
rect 51 156 52 157
rect 50 156 51 157
rect 49 156 50 157
rect 48 156 49 157
rect 47 156 48 157
rect 46 156 47 157
rect 45 156 46 157
rect 44 156 45 157
rect 43 156 44 157
rect 42 156 43 157
rect 41 156 42 157
rect 40 156 41 157
rect 39 156 40 157
rect 30 156 31 157
rect 29 156 30 157
rect 28 156 29 157
rect 27 156 28 157
rect 26 156 27 157
rect 25 156 26 157
rect 24 156 25 157
rect 23 156 24 157
rect 22 156 23 157
rect 21 156 22 157
rect 20 156 21 157
rect 19 156 20 157
rect 18 156 19 157
rect 17 156 18 157
rect 16 156 17 157
rect 15 156 16 157
rect 14 156 15 157
rect 13 156 14 157
rect 12 156 13 157
rect 11 156 12 157
rect 10 156 11 157
rect 441 157 442 158
rect 440 157 441 158
rect 399 157 400 158
rect 398 157 399 158
rect 397 157 398 158
rect 326 157 327 158
rect 325 157 326 158
rect 324 157 325 158
rect 323 157 324 158
rect 322 157 323 158
rect 321 157 322 158
rect 320 157 321 158
rect 319 157 320 158
rect 318 157 319 158
rect 317 157 318 158
rect 316 157 317 158
rect 315 157 316 158
rect 314 157 315 158
rect 313 157 314 158
rect 312 157 313 158
rect 311 157 312 158
rect 310 157 311 158
rect 309 157 310 158
rect 308 157 309 158
rect 307 157 308 158
rect 306 157 307 158
rect 305 157 306 158
rect 304 157 305 158
rect 303 157 304 158
rect 302 157 303 158
rect 301 157 302 158
rect 300 157 301 158
rect 299 157 300 158
rect 298 157 299 158
rect 297 157 298 158
rect 296 157 297 158
rect 295 157 296 158
rect 294 157 295 158
rect 293 157 294 158
rect 292 157 293 158
rect 291 157 292 158
rect 290 157 291 158
rect 289 157 290 158
rect 288 157 289 158
rect 287 157 288 158
rect 286 157 287 158
rect 285 157 286 158
rect 284 157 285 158
rect 283 157 284 158
rect 282 157 283 158
rect 281 157 282 158
rect 280 157 281 158
rect 279 157 280 158
rect 278 157 279 158
rect 277 157 278 158
rect 276 157 277 158
rect 275 157 276 158
rect 274 157 275 158
rect 273 157 274 158
rect 272 157 273 158
rect 271 157 272 158
rect 270 157 271 158
rect 269 157 270 158
rect 268 157 269 158
rect 267 157 268 158
rect 266 157 267 158
rect 265 157 266 158
rect 264 157 265 158
rect 263 157 264 158
rect 262 157 263 158
rect 261 157 262 158
rect 260 157 261 158
rect 259 157 260 158
rect 258 157 259 158
rect 257 157 258 158
rect 256 157 257 158
rect 255 157 256 158
rect 254 157 255 158
rect 253 157 254 158
rect 252 157 253 158
rect 251 157 252 158
rect 250 157 251 158
rect 249 157 250 158
rect 248 157 249 158
rect 247 157 248 158
rect 246 157 247 158
rect 245 157 246 158
rect 244 157 245 158
rect 243 157 244 158
rect 242 157 243 158
rect 241 157 242 158
rect 240 157 241 158
rect 239 157 240 158
rect 238 157 239 158
rect 218 157 219 158
rect 217 157 218 158
rect 216 157 217 158
rect 215 157 216 158
rect 214 157 215 158
rect 213 157 214 158
rect 212 157 213 158
rect 211 157 212 158
rect 210 157 211 158
rect 209 157 210 158
rect 208 157 209 158
rect 207 157 208 158
rect 206 157 207 158
rect 205 157 206 158
rect 204 157 205 158
rect 203 157 204 158
rect 202 157 203 158
rect 201 157 202 158
rect 200 157 201 158
rect 199 157 200 158
rect 198 157 199 158
rect 197 157 198 158
rect 196 157 197 158
rect 195 157 196 158
rect 194 157 195 158
rect 193 157 194 158
rect 192 157 193 158
rect 191 157 192 158
rect 190 157 191 158
rect 189 157 190 158
rect 188 157 189 158
rect 187 157 188 158
rect 186 157 187 158
rect 185 157 186 158
rect 184 157 185 158
rect 183 157 184 158
rect 182 157 183 158
rect 181 157 182 158
rect 180 157 181 158
rect 179 157 180 158
rect 178 157 179 158
rect 177 157 178 158
rect 176 157 177 158
rect 175 157 176 158
rect 174 157 175 158
rect 173 157 174 158
rect 172 157 173 158
rect 171 157 172 158
rect 170 157 171 158
rect 169 157 170 158
rect 168 157 169 158
rect 167 157 168 158
rect 166 157 167 158
rect 165 157 166 158
rect 164 157 165 158
rect 163 157 164 158
rect 162 157 163 158
rect 161 157 162 158
rect 160 157 161 158
rect 159 157 160 158
rect 158 157 159 158
rect 157 157 158 158
rect 156 157 157 158
rect 155 157 156 158
rect 154 157 155 158
rect 153 157 154 158
rect 152 157 153 158
rect 121 157 122 158
rect 120 157 121 158
rect 119 157 120 158
rect 118 157 119 158
rect 117 157 118 158
rect 116 157 117 158
rect 115 157 116 158
rect 114 157 115 158
rect 113 157 114 158
rect 112 157 113 158
rect 111 157 112 158
rect 110 157 111 158
rect 109 157 110 158
rect 108 157 109 158
rect 107 157 108 158
rect 106 157 107 158
rect 105 157 106 158
rect 104 157 105 158
rect 103 157 104 158
rect 102 157 103 158
rect 101 157 102 158
rect 100 157 101 158
rect 99 157 100 158
rect 98 157 99 158
rect 97 157 98 158
rect 96 157 97 158
rect 95 157 96 158
rect 94 157 95 158
rect 93 157 94 158
rect 92 157 93 158
rect 91 157 92 158
rect 90 157 91 158
rect 89 157 90 158
rect 88 157 89 158
rect 87 157 88 158
rect 86 157 87 158
rect 85 157 86 158
rect 84 157 85 158
rect 83 157 84 158
rect 82 157 83 158
rect 81 157 82 158
rect 80 157 81 158
rect 79 157 80 158
rect 78 157 79 158
rect 77 157 78 158
rect 76 157 77 158
rect 75 157 76 158
rect 74 157 75 158
rect 73 157 74 158
rect 72 157 73 158
rect 71 157 72 158
rect 70 157 71 158
rect 69 157 70 158
rect 68 157 69 158
rect 67 157 68 158
rect 66 157 67 158
rect 65 157 66 158
rect 64 157 65 158
rect 63 157 64 158
rect 62 157 63 158
rect 61 157 62 158
rect 60 157 61 158
rect 59 157 60 158
rect 58 157 59 158
rect 57 157 58 158
rect 56 157 57 158
rect 55 157 56 158
rect 54 157 55 158
rect 53 157 54 158
rect 52 157 53 158
rect 51 157 52 158
rect 50 157 51 158
rect 49 157 50 158
rect 48 157 49 158
rect 47 157 48 158
rect 46 157 47 158
rect 45 157 46 158
rect 44 157 45 158
rect 43 157 44 158
rect 42 157 43 158
rect 41 157 42 158
rect 40 157 41 158
rect 39 157 40 158
rect 38 157 39 158
rect 30 157 31 158
rect 29 157 30 158
rect 28 157 29 158
rect 27 157 28 158
rect 26 157 27 158
rect 25 157 26 158
rect 24 157 25 158
rect 23 157 24 158
rect 22 157 23 158
rect 21 157 22 158
rect 20 157 21 158
rect 19 157 20 158
rect 18 157 19 158
rect 17 157 18 158
rect 16 157 17 158
rect 15 157 16 158
rect 14 157 15 158
rect 13 157 14 158
rect 12 157 13 158
rect 11 157 12 158
rect 10 157 11 158
rect 441 158 442 159
rect 440 158 441 159
rect 439 158 440 159
rect 399 158 400 159
rect 398 158 399 159
rect 397 158 398 159
rect 327 158 328 159
rect 326 158 327 159
rect 325 158 326 159
rect 324 158 325 159
rect 323 158 324 159
rect 322 158 323 159
rect 321 158 322 159
rect 320 158 321 159
rect 319 158 320 159
rect 318 158 319 159
rect 317 158 318 159
rect 316 158 317 159
rect 315 158 316 159
rect 314 158 315 159
rect 313 158 314 159
rect 312 158 313 159
rect 311 158 312 159
rect 310 158 311 159
rect 309 158 310 159
rect 308 158 309 159
rect 307 158 308 159
rect 306 158 307 159
rect 305 158 306 159
rect 304 158 305 159
rect 303 158 304 159
rect 302 158 303 159
rect 301 158 302 159
rect 300 158 301 159
rect 299 158 300 159
rect 298 158 299 159
rect 297 158 298 159
rect 296 158 297 159
rect 295 158 296 159
rect 294 158 295 159
rect 293 158 294 159
rect 292 158 293 159
rect 291 158 292 159
rect 290 158 291 159
rect 289 158 290 159
rect 288 158 289 159
rect 287 158 288 159
rect 286 158 287 159
rect 285 158 286 159
rect 284 158 285 159
rect 283 158 284 159
rect 282 158 283 159
rect 281 158 282 159
rect 280 158 281 159
rect 279 158 280 159
rect 278 158 279 159
rect 277 158 278 159
rect 276 158 277 159
rect 275 158 276 159
rect 274 158 275 159
rect 273 158 274 159
rect 272 158 273 159
rect 271 158 272 159
rect 270 158 271 159
rect 269 158 270 159
rect 268 158 269 159
rect 267 158 268 159
rect 266 158 267 159
rect 265 158 266 159
rect 264 158 265 159
rect 263 158 264 159
rect 262 158 263 159
rect 261 158 262 159
rect 260 158 261 159
rect 259 158 260 159
rect 258 158 259 159
rect 257 158 258 159
rect 256 158 257 159
rect 255 158 256 159
rect 254 158 255 159
rect 253 158 254 159
rect 252 158 253 159
rect 251 158 252 159
rect 250 158 251 159
rect 249 158 250 159
rect 248 158 249 159
rect 247 158 248 159
rect 246 158 247 159
rect 245 158 246 159
rect 244 158 245 159
rect 243 158 244 159
rect 242 158 243 159
rect 241 158 242 159
rect 240 158 241 159
rect 239 158 240 159
rect 238 158 239 159
rect 237 158 238 159
rect 218 158 219 159
rect 217 158 218 159
rect 216 158 217 159
rect 215 158 216 159
rect 214 158 215 159
rect 213 158 214 159
rect 212 158 213 159
rect 211 158 212 159
rect 210 158 211 159
rect 209 158 210 159
rect 208 158 209 159
rect 207 158 208 159
rect 206 158 207 159
rect 205 158 206 159
rect 204 158 205 159
rect 203 158 204 159
rect 202 158 203 159
rect 201 158 202 159
rect 200 158 201 159
rect 199 158 200 159
rect 198 158 199 159
rect 197 158 198 159
rect 196 158 197 159
rect 195 158 196 159
rect 194 158 195 159
rect 193 158 194 159
rect 192 158 193 159
rect 191 158 192 159
rect 190 158 191 159
rect 189 158 190 159
rect 188 158 189 159
rect 187 158 188 159
rect 186 158 187 159
rect 185 158 186 159
rect 184 158 185 159
rect 183 158 184 159
rect 182 158 183 159
rect 181 158 182 159
rect 180 158 181 159
rect 179 158 180 159
rect 178 158 179 159
rect 177 158 178 159
rect 176 158 177 159
rect 175 158 176 159
rect 174 158 175 159
rect 173 158 174 159
rect 172 158 173 159
rect 171 158 172 159
rect 170 158 171 159
rect 169 158 170 159
rect 168 158 169 159
rect 167 158 168 159
rect 166 158 167 159
rect 165 158 166 159
rect 164 158 165 159
rect 163 158 164 159
rect 162 158 163 159
rect 161 158 162 159
rect 160 158 161 159
rect 159 158 160 159
rect 158 158 159 159
rect 157 158 158 159
rect 156 158 157 159
rect 155 158 156 159
rect 154 158 155 159
rect 153 158 154 159
rect 152 158 153 159
rect 151 158 152 159
rect 120 158 121 159
rect 119 158 120 159
rect 118 158 119 159
rect 117 158 118 159
rect 116 158 117 159
rect 115 158 116 159
rect 114 158 115 159
rect 113 158 114 159
rect 112 158 113 159
rect 111 158 112 159
rect 110 158 111 159
rect 109 158 110 159
rect 108 158 109 159
rect 107 158 108 159
rect 106 158 107 159
rect 105 158 106 159
rect 104 158 105 159
rect 103 158 104 159
rect 102 158 103 159
rect 101 158 102 159
rect 100 158 101 159
rect 99 158 100 159
rect 98 158 99 159
rect 97 158 98 159
rect 96 158 97 159
rect 95 158 96 159
rect 94 158 95 159
rect 93 158 94 159
rect 92 158 93 159
rect 91 158 92 159
rect 90 158 91 159
rect 89 158 90 159
rect 88 158 89 159
rect 87 158 88 159
rect 86 158 87 159
rect 85 158 86 159
rect 84 158 85 159
rect 83 158 84 159
rect 82 158 83 159
rect 81 158 82 159
rect 80 158 81 159
rect 79 158 80 159
rect 78 158 79 159
rect 77 158 78 159
rect 76 158 77 159
rect 75 158 76 159
rect 74 158 75 159
rect 73 158 74 159
rect 72 158 73 159
rect 71 158 72 159
rect 70 158 71 159
rect 69 158 70 159
rect 68 158 69 159
rect 67 158 68 159
rect 66 158 67 159
rect 65 158 66 159
rect 64 158 65 159
rect 63 158 64 159
rect 62 158 63 159
rect 61 158 62 159
rect 60 158 61 159
rect 59 158 60 159
rect 58 158 59 159
rect 57 158 58 159
rect 56 158 57 159
rect 55 158 56 159
rect 54 158 55 159
rect 53 158 54 159
rect 52 158 53 159
rect 51 158 52 159
rect 50 158 51 159
rect 49 158 50 159
rect 48 158 49 159
rect 47 158 48 159
rect 46 158 47 159
rect 45 158 46 159
rect 44 158 45 159
rect 43 158 44 159
rect 42 158 43 159
rect 41 158 42 159
rect 40 158 41 159
rect 39 158 40 159
rect 38 158 39 159
rect 29 158 30 159
rect 28 158 29 159
rect 27 158 28 159
rect 26 158 27 159
rect 25 158 26 159
rect 24 158 25 159
rect 23 158 24 159
rect 22 158 23 159
rect 21 158 22 159
rect 20 158 21 159
rect 19 158 20 159
rect 18 158 19 159
rect 17 158 18 159
rect 16 158 17 159
rect 15 158 16 159
rect 14 158 15 159
rect 13 158 14 159
rect 12 158 13 159
rect 11 158 12 159
rect 10 158 11 159
rect 441 159 442 160
rect 440 159 441 160
rect 439 159 440 160
rect 399 159 400 160
rect 398 159 399 160
rect 397 159 398 160
rect 328 159 329 160
rect 327 159 328 160
rect 326 159 327 160
rect 325 159 326 160
rect 324 159 325 160
rect 323 159 324 160
rect 322 159 323 160
rect 321 159 322 160
rect 320 159 321 160
rect 319 159 320 160
rect 318 159 319 160
rect 317 159 318 160
rect 316 159 317 160
rect 315 159 316 160
rect 314 159 315 160
rect 313 159 314 160
rect 312 159 313 160
rect 311 159 312 160
rect 310 159 311 160
rect 309 159 310 160
rect 308 159 309 160
rect 307 159 308 160
rect 306 159 307 160
rect 305 159 306 160
rect 304 159 305 160
rect 303 159 304 160
rect 302 159 303 160
rect 301 159 302 160
rect 300 159 301 160
rect 299 159 300 160
rect 298 159 299 160
rect 297 159 298 160
rect 296 159 297 160
rect 295 159 296 160
rect 294 159 295 160
rect 293 159 294 160
rect 292 159 293 160
rect 291 159 292 160
rect 290 159 291 160
rect 289 159 290 160
rect 288 159 289 160
rect 287 159 288 160
rect 286 159 287 160
rect 285 159 286 160
rect 284 159 285 160
rect 283 159 284 160
rect 282 159 283 160
rect 281 159 282 160
rect 280 159 281 160
rect 279 159 280 160
rect 278 159 279 160
rect 277 159 278 160
rect 276 159 277 160
rect 275 159 276 160
rect 274 159 275 160
rect 273 159 274 160
rect 272 159 273 160
rect 271 159 272 160
rect 270 159 271 160
rect 269 159 270 160
rect 268 159 269 160
rect 267 159 268 160
rect 266 159 267 160
rect 265 159 266 160
rect 264 159 265 160
rect 263 159 264 160
rect 262 159 263 160
rect 261 159 262 160
rect 260 159 261 160
rect 259 159 260 160
rect 258 159 259 160
rect 257 159 258 160
rect 256 159 257 160
rect 255 159 256 160
rect 254 159 255 160
rect 253 159 254 160
rect 252 159 253 160
rect 251 159 252 160
rect 250 159 251 160
rect 249 159 250 160
rect 248 159 249 160
rect 247 159 248 160
rect 246 159 247 160
rect 245 159 246 160
rect 244 159 245 160
rect 243 159 244 160
rect 242 159 243 160
rect 241 159 242 160
rect 240 159 241 160
rect 239 159 240 160
rect 238 159 239 160
rect 237 159 238 160
rect 217 159 218 160
rect 216 159 217 160
rect 215 159 216 160
rect 214 159 215 160
rect 213 159 214 160
rect 212 159 213 160
rect 211 159 212 160
rect 210 159 211 160
rect 209 159 210 160
rect 208 159 209 160
rect 207 159 208 160
rect 206 159 207 160
rect 205 159 206 160
rect 204 159 205 160
rect 203 159 204 160
rect 202 159 203 160
rect 201 159 202 160
rect 200 159 201 160
rect 199 159 200 160
rect 198 159 199 160
rect 197 159 198 160
rect 196 159 197 160
rect 195 159 196 160
rect 194 159 195 160
rect 193 159 194 160
rect 192 159 193 160
rect 191 159 192 160
rect 190 159 191 160
rect 189 159 190 160
rect 188 159 189 160
rect 187 159 188 160
rect 186 159 187 160
rect 185 159 186 160
rect 184 159 185 160
rect 183 159 184 160
rect 182 159 183 160
rect 181 159 182 160
rect 180 159 181 160
rect 179 159 180 160
rect 178 159 179 160
rect 177 159 178 160
rect 176 159 177 160
rect 175 159 176 160
rect 174 159 175 160
rect 173 159 174 160
rect 172 159 173 160
rect 171 159 172 160
rect 170 159 171 160
rect 169 159 170 160
rect 168 159 169 160
rect 167 159 168 160
rect 166 159 167 160
rect 165 159 166 160
rect 164 159 165 160
rect 163 159 164 160
rect 162 159 163 160
rect 161 159 162 160
rect 160 159 161 160
rect 159 159 160 160
rect 158 159 159 160
rect 157 159 158 160
rect 156 159 157 160
rect 155 159 156 160
rect 154 159 155 160
rect 153 159 154 160
rect 152 159 153 160
rect 151 159 152 160
rect 150 159 151 160
rect 119 159 120 160
rect 118 159 119 160
rect 117 159 118 160
rect 116 159 117 160
rect 115 159 116 160
rect 114 159 115 160
rect 113 159 114 160
rect 112 159 113 160
rect 111 159 112 160
rect 110 159 111 160
rect 109 159 110 160
rect 108 159 109 160
rect 107 159 108 160
rect 106 159 107 160
rect 105 159 106 160
rect 104 159 105 160
rect 103 159 104 160
rect 102 159 103 160
rect 101 159 102 160
rect 100 159 101 160
rect 99 159 100 160
rect 98 159 99 160
rect 97 159 98 160
rect 96 159 97 160
rect 95 159 96 160
rect 94 159 95 160
rect 93 159 94 160
rect 92 159 93 160
rect 91 159 92 160
rect 90 159 91 160
rect 89 159 90 160
rect 88 159 89 160
rect 87 159 88 160
rect 86 159 87 160
rect 85 159 86 160
rect 84 159 85 160
rect 83 159 84 160
rect 82 159 83 160
rect 81 159 82 160
rect 80 159 81 160
rect 79 159 80 160
rect 78 159 79 160
rect 77 159 78 160
rect 76 159 77 160
rect 75 159 76 160
rect 74 159 75 160
rect 73 159 74 160
rect 72 159 73 160
rect 71 159 72 160
rect 70 159 71 160
rect 69 159 70 160
rect 68 159 69 160
rect 67 159 68 160
rect 66 159 67 160
rect 65 159 66 160
rect 64 159 65 160
rect 63 159 64 160
rect 62 159 63 160
rect 61 159 62 160
rect 60 159 61 160
rect 59 159 60 160
rect 58 159 59 160
rect 57 159 58 160
rect 56 159 57 160
rect 55 159 56 160
rect 54 159 55 160
rect 53 159 54 160
rect 52 159 53 160
rect 51 159 52 160
rect 50 159 51 160
rect 49 159 50 160
rect 48 159 49 160
rect 47 159 48 160
rect 46 159 47 160
rect 45 159 46 160
rect 44 159 45 160
rect 43 159 44 160
rect 42 159 43 160
rect 41 159 42 160
rect 40 159 41 160
rect 39 159 40 160
rect 38 159 39 160
rect 37 159 38 160
rect 29 159 30 160
rect 28 159 29 160
rect 27 159 28 160
rect 26 159 27 160
rect 25 159 26 160
rect 24 159 25 160
rect 23 159 24 160
rect 22 159 23 160
rect 21 159 22 160
rect 20 159 21 160
rect 19 159 20 160
rect 18 159 19 160
rect 17 159 18 160
rect 16 159 17 160
rect 15 159 16 160
rect 14 159 15 160
rect 13 159 14 160
rect 12 159 13 160
rect 11 159 12 160
rect 10 159 11 160
rect 9 159 10 160
rect 441 160 442 161
rect 440 160 441 161
rect 439 160 440 161
rect 400 160 401 161
rect 399 160 400 161
rect 398 160 399 161
rect 397 160 398 161
rect 328 160 329 161
rect 327 160 328 161
rect 326 160 327 161
rect 325 160 326 161
rect 324 160 325 161
rect 323 160 324 161
rect 322 160 323 161
rect 321 160 322 161
rect 320 160 321 161
rect 319 160 320 161
rect 318 160 319 161
rect 317 160 318 161
rect 298 160 299 161
rect 297 160 298 161
rect 296 160 297 161
rect 295 160 296 161
rect 294 160 295 161
rect 293 160 294 161
rect 292 160 293 161
rect 291 160 292 161
rect 290 160 291 161
rect 289 160 290 161
rect 288 160 289 161
rect 287 160 288 161
rect 286 160 287 161
rect 285 160 286 161
rect 284 160 285 161
rect 283 160 284 161
rect 282 160 283 161
rect 281 160 282 161
rect 280 160 281 161
rect 279 160 280 161
rect 278 160 279 161
rect 277 160 278 161
rect 276 160 277 161
rect 275 160 276 161
rect 274 160 275 161
rect 273 160 274 161
rect 272 160 273 161
rect 271 160 272 161
rect 270 160 271 161
rect 269 160 270 161
rect 268 160 269 161
rect 267 160 268 161
rect 266 160 267 161
rect 265 160 266 161
rect 264 160 265 161
rect 263 160 264 161
rect 262 160 263 161
rect 261 160 262 161
rect 260 160 261 161
rect 259 160 260 161
rect 258 160 259 161
rect 257 160 258 161
rect 256 160 257 161
rect 255 160 256 161
rect 254 160 255 161
rect 253 160 254 161
rect 252 160 253 161
rect 251 160 252 161
rect 250 160 251 161
rect 249 160 250 161
rect 248 160 249 161
rect 247 160 248 161
rect 246 160 247 161
rect 245 160 246 161
rect 244 160 245 161
rect 243 160 244 161
rect 242 160 243 161
rect 241 160 242 161
rect 240 160 241 161
rect 239 160 240 161
rect 238 160 239 161
rect 237 160 238 161
rect 236 160 237 161
rect 217 160 218 161
rect 216 160 217 161
rect 215 160 216 161
rect 214 160 215 161
rect 213 160 214 161
rect 212 160 213 161
rect 211 160 212 161
rect 210 160 211 161
rect 209 160 210 161
rect 208 160 209 161
rect 207 160 208 161
rect 206 160 207 161
rect 205 160 206 161
rect 204 160 205 161
rect 203 160 204 161
rect 202 160 203 161
rect 201 160 202 161
rect 200 160 201 161
rect 199 160 200 161
rect 198 160 199 161
rect 197 160 198 161
rect 196 160 197 161
rect 195 160 196 161
rect 194 160 195 161
rect 193 160 194 161
rect 192 160 193 161
rect 191 160 192 161
rect 190 160 191 161
rect 189 160 190 161
rect 188 160 189 161
rect 187 160 188 161
rect 186 160 187 161
rect 185 160 186 161
rect 184 160 185 161
rect 183 160 184 161
rect 182 160 183 161
rect 181 160 182 161
rect 180 160 181 161
rect 179 160 180 161
rect 178 160 179 161
rect 177 160 178 161
rect 176 160 177 161
rect 175 160 176 161
rect 174 160 175 161
rect 173 160 174 161
rect 172 160 173 161
rect 171 160 172 161
rect 170 160 171 161
rect 169 160 170 161
rect 168 160 169 161
rect 167 160 168 161
rect 166 160 167 161
rect 165 160 166 161
rect 164 160 165 161
rect 163 160 164 161
rect 162 160 163 161
rect 161 160 162 161
rect 160 160 161 161
rect 159 160 160 161
rect 158 160 159 161
rect 157 160 158 161
rect 156 160 157 161
rect 155 160 156 161
rect 154 160 155 161
rect 153 160 154 161
rect 152 160 153 161
rect 151 160 152 161
rect 150 160 151 161
rect 149 160 150 161
rect 117 160 118 161
rect 116 160 117 161
rect 115 160 116 161
rect 114 160 115 161
rect 113 160 114 161
rect 112 160 113 161
rect 111 160 112 161
rect 110 160 111 161
rect 109 160 110 161
rect 108 160 109 161
rect 107 160 108 161
rect 106 160 107 161
rect 105 160 106 161
rect 104 160 105 161
rect 103 160 104 161
rect 102 160 103 161
rect 101 160 102 161
rect 100 160 101 161
rect 99 160 100 161
rect 98 160 99 161
rect 97 160 98 161
rect 96 160 97 161
rect 95 160 96 161
rect 94 160 95 161
rect 93 160 94 161
rect 92 160 93 161
rect 91 160 92 161
rect 90 160 91 161
rect 89 160 90 161
rect 88 160 89 161
rect 87 160 88 161
rect 86 160 87 161
rect 85 160 86 161
rect 84 160 85 161
rect 83 160 84 161
rect 82 160 83 161
rect 81 160 82 161
rect 80 160 81 161
rect 79 160 80 161
rect 78 160 79 161
rect 77 160 78 161
rect 76 160 77 161
rect 75 160 76 161
rect 74 160 75 161
rect 73 160 74 161
rect 72 160 73 161
rect 71 160 72 161
rect 70 160 71 161
rect 69 160 70 161
rect 68 160 69 161
rect 67 160 68 161
rect 66 160 67 161
rect 65 160 66 161
rect 64 160 65 161
rect 63 160 64 161
rect 62 160 63 161
rect 61 160 62 161
rect 60 160 61 161
rect 59 160 60 161
rect 58 160 59 161
rect 57 160 58 161
rect 56 160 57 161
rect 55 160 56 161
rect 54 160 55 161
rect 53 160 54 161
rect 52 160 53 161
rect 51 160 52 161
rect 50 160 51 161
rect 49 160 50 161
rect 48 160 49 161
rect 47 160 48 161
rect 46 160 47 161
rect 45 160 46 161
rect 44 160 45 161
rect 43 160 44 161
rect 42 160 43 161
rect 41 160 42 161
rect 40 160 41 161
rect 39 160 40 161
rect 38 160 39 161
rect 37 160 38 161
rect 28 160 29 161
rect 27 160 28 161
rect 26 160 27 161
rect 25 160 26 161
rect 24 160 25 161
rect 23 160 24 161
rect 22 160 23 161
rect 21 160 22 161
rect 20 160 21 161
rect 19 160 20 161
rect 18 160 19 161
rect 17 160 18 161
rect 16 160 17 161
rect 15 160 16 161
rect 14 160 15 161
rect 13 160 14 161
rect 12 160 13 161
rect 11 160 12 161
rect 10 160 11 161
rect 9 160 10 161
rect 441 161 442 162
rect 440 161 441 162
rect 439 161 440 162
rect 438 161 439 162
rect 400 161 401 162
rect 399 161 400 162
rect 398 161 399 162
rect 397 161 398 162
rect 329 161 330 162
rect 328 161 329 162
rect 327 161 328 162
rect 326 161 327 162
rect 325 161 326 162
rect 324 161 325 162
rect 323 161 324 162
rect 294 161 295 162
rect 293 161 294 162
rect 292 161 293 162
rect 291 161 292 162
rect 290 161 291 162
rect 289 161 290 162
rect 288 161 289 162
rect 287 161 288 162
rect 286 161 287 162
rect 285 161 286 162
rect 284 161 285 162
rect 283 161 284 162
rect 282 161 283 162
rect 281 161 282 162
rect 280 161 281 162
rect 279 161 280 162
rect 278 161 279 162
rect 277 161 278 162
rect 276 161 277 162
rect 275 161 276 162
rect 274 161 275 162
rect 273 161 274 162
rect 272 161 273 162
rect 271 161 272 162
rect 270 161 271 162
rect 269 161 270 162
rect 268 161 269 162
rect 267 161 268 162
rect 266 161 267 162
rect 265 161 266 162
rect 264 161 265 162
rect 263 161 264 162
rect 262 161 263 162
rect 261 161 262 162
rect 260 161 261 162
rect 259 161 260 162
rect 258 161 259 162
rect 257 161 258 162
rect 256 161 257 162
rect 255 161 256 162
rect 254 161 255 162
rect 253 161 254 162
rect 252 161 253 162
rect 251 161 252 162
rect 250 161 251 162
rect 249 161 250 162
rect 248 161 249 162
rect 247 161 248 162
rect 246 161 247 162
rect 245 161 246 162
rect 244 161 245 162
rect 243 161 244 162
rect 242 161 243 162
rect 241 161 242 162
rect 240 161 241 162
rect 239 161 240 162
rect 238 161 239 162
rect 237 161 238 162
rect 236 161 237 162
rect 235 161 236 162
rect 216 161 217 162
rect 215 161 216 162
rect 214 161 215 162
rect 213 161 214 162
rect 212 161 213 162
rect 211 161 212 162
rect 210 161 211 162
rect 209 161 210 162
rect 208 161 209 162
rect 207 161 208 162
rect 206 161 207 162
rect 205 161 206 162
rect 204 161 205 162
rect 203 161 204 162
rect 202 161 203 162
rect 201 161 202 162
rect 200 161 201 162
rect 199 161 200 162
rect 198 161 199 162
rect 197 161 198 162
rect 196 161 197 162
rect 195 161 196 162
rect 194 161 195 162
rect 193 161 194 162
rect 192 161 193 162
rect 191 161 192 162
rect 190 161 191 162
rect 189 161 190 162
rect 188 161 189 162
rect 187 161 188 162
rect 186 161 187 162
rect 185 161 186 162
rect 184 161 185 162
rect 183 161 184 162
rect 182 161 183 162
rect 181 161 182 162
rect 180 161 181 162
rect 179 161 180 162
rect 178 161 179 162
rect 177 161 178 162
rect 176 161 177 162
rect 175 161 176 162
rect 174 161 175 162
rect 173 161 174 162
rect 172 161 173 162
rect 171 161 172 162
rect 170 161 171 162
rect 169 161 170 162
rect 168 161 169 162
rect 167 161 168 162
rect 166 161 167 162
rect 165 161 166 162
rect 164 161 165 162
rect 163 161 164 162
rect 162 161 163 162
rect 161 161 162 162
rect 160 161 161 162
rect 159 161 160 162
rect 158 161 159 162
rect 157 161 158 162
rect 156 161 157 162
rect 155 161 156 162
rect 154 161 155 162
rect 153 161 154 162
rect 152 161 153 162
rect 151 161 152 162
rect 150 161 151 162
rect 149 161 150 162
rect 116 161 117 162
rect 115 161 116 162
rect 114 161 115 162
rect 113 161 114 162
rect 112 161 113 162
rect 111 161 112 162
rect 110 161 111 162
rect 109 161 110 162
rect 108 161 109 162
rect 107 161 108 162
rect 106 161 107 162
rect 105 161 106 162
rect 104 161 105 162
rect 103 161 104 162
rect 102 161 103 162
rect 101 161 102 162
rect 100 161 101 162
rect 99 161 100 162
rect 98 161 99 162
rect 97 161 98 162
rect 96 161 97 162
rect 95 161 96 162
rect 94 161 95 162
rect 93 161 94 162
rect 92 161 93 162
rect 91 161 92 162
rect 90 161 91 162
rect 89 161 90 162
rect 88 161 89 162
rect 87 161 88 162
rect 86 161 87 162
rect 85 161 86 162
rect 84 161 85 162
rect 83 161 84 162
rect 82 161 83 162
rect 81 161 82 162
rect 80 161 81 162
rect 79 161 80 162
rect 78 161 79 162
rect 77 161 78 162
rect 76 161 77 162
rect 75 161 76 162
rect 74 161 75 162
rect 73 161 74 162
rect 72 161 73 162
rect 71 161 72 162
rect 70 161 71 162
rect 69 161 70 162
rect 68 161 69 162
rect 67 161 68 162
rect 66 161 67 162
rect 65 161 66 162
rect 64 161 65 162
rect 63 161 64 162
rect 62 161 63 162
rect 61 161 62 162
rect 60 161 61 162
rect 59 161 60 162
rect 58 161 59 162
rect 57 161 58 162
rect 56 161 57 162
rect 55 161 56 162
rect 54 161 55 162
rect 53 161 54 162
rect 52 161 53 162
rect 51 161 52 162
rect 50 161 51 162
rect 49 161 50 162
rect 48 161 49 162
rect 47 161 48 162
rect 46 161 47 162
rect 45 161 46 162
rect 44 161 45 162
rect 43 161 44 162
rect 42 161 43 162
rect 41 161 42 162
rect 40 161 41 162
rect 39 161 40 162
rect 38 161 39 162
rect 37 161 38 162
rect 36 161 37 162
rect 27 161 28 162
rect 26 161 27 162
rect 25 161 26 162
rect 24 161 25 162
rect 23 161 24 162
rect 22 161 23 162
rect 21 161 22 162
rect 20 161 21 162
rect 19 161 20 162
rect 18 161 19 162
rect 17 161 18 162
rect 16 161 17 162
rect 15 161 16 162
rect 14 161 15 162
rect 13 161 14 162
rect 12 161 13 162
rect 11 161 12 162
rect 10 161 11 162
rect 9 161 10 162
rect 462 162 463 163
rect 441 162 442 163
rect 440 162 441 163
rect 439 162 440 163
rect 438 162 439 163
rect 437 162 438 163
rect 436 162 437 163
rect 402 162 403 163
rect 401 162 402 163
rect 400 162 401 163
rect 399 162 400 163
rect 398 162 399 163
rect 397 162 398 163
rect 330 162 331 163
rect 329 162 330 163
rect 328 162 329 163
rect 327 162 328 163
rect 291 162 292 163
rect 290 162 291 163
rect 289 162 290 163
rect 288 162 289 163
rect 287 162 288 163
rect 286 162 287 163
rect 285 162 286 163
rect 284 162 285 163
rect 283 162 284 163
rect 282 162 283 163
rect 281 162 282 163
rect 280 162 281 163
rect 279 162 280 163
rect 278 162 279 163
rect 277 162 278 163
rect 276 162 277 163
rect 275 162 276 163
rect 274 162 275 163
rect 273 162 274 163
rect 272 162 273 163
rect 271 162 272 163
rect 270 162 271 163
rect 269 162 270 163
rect 268 162 269 163
rect 267 162 268 163
rect 266 162 267 163
rect 265 162 266 163
rect 264 162 265 163
rect 263 162 264 163
rect 262 162 263 163
rect 261 162 262 163
rect 260 162 261 163
rect 259 162 260 163
rect 258 162 259 163
rect 257 162 258 163
rect 256 162 257 163
rect 255 162 256 163
rect 254 162 255 163
rect 253 162 254 163
rect 252 162 253 163
rect 251 162 252 163
rect 250 162 251 163
rect 249 162 250 163
rect 248 162 249 163
rect 247 162 248 163
rect 246 162 247 163
rect 245 162 246 163
rect 244 162 245 163
rect 243 162 244 163
rect 242 162 243 163
rect 241 162 242 163
rect 240 162 241 163
rect 239 162 240 163
rect 238 162 239 163
rect 237 162 238 163
rect 236 162 237 163
rect 235 162 236 163
rect 216 162 217 163
rect 215 162 216 163
rect 214 162 215 163
rect 213 162 214 163
rect 212 162 213 163
rect 211 162 212 163
rect 210 162 211 163
rect 209 162 210 163
rect 208 162 209 163
rect 207 162 208 163
rect 206 162 207 163
rect 205 162 206 163
rect 204 162 205 163
rect 203 162 204 163
rect 202 162 203 163
rect 201 162 202 163
rect 200 162 201 163
rect 199 162 200 163
rect 198 162 199 163
rect 197 162 198 163
rect 196 162 197 163
rect 195 162 196 163
rect 194 162 195 163
rect 193 162 194 163
rect 192 162 193 163
rect 191 162 192 163
rect 190 162 191 163
rect 189 162 190 163
rect 188 162 189 163
rect 187 162 188 163
rect 186 162 187 163
rect 185 162 186 163
rect 184 162 185 163
rect 183 162 184 163
rect 182 162 183 163
rect 181 162 182 163
rect 180 162 181 163
rect 179 162 180 163
rect 178 162 179 163
rect 177 162 178 163
rect 176 162 177 163
rect 175 162 176 163
rect 174 162 175 163
rect 173 162 174 163
rect 172 162 173 163
rect 171 162 172 163
rect 170 162 171 163
rect 169 162 170 163
rect 168 162 169 163
rect 167 162 168 163
rect 166 162 167 163
rect 165 162 166 163
rect 164 162 165 163
rect 163 162 164 163
rect 162 162 163 163
rect 161 162 162 163
rect 160 162 161 163
rect 159 162 160 163
rect 158 162 159 163
rect 157 162 158 163
rect 156 162 157 163
rect 155 162 156 163
rect 154 162 155 163
rect 153 162 154 163
rect 152 162 153 163
rect 151 162 152 163
rect 150 162 151 163
rect 149 162 150 163
rect 148 162 149 163
rect 114 162 115 163
rect 113 162 114 163
rect 112 162 113 163
rect 111 162 112 163
rect 110 162 111 163
rect 109 162 110 163
rect 108 162 109 163
rect 107 162 108 163
rect 106 162 107 163
rect 105 162 106 163
rect 104 162 105 163
rect 103 162 104 163
rect 102 162 103 163
rect 101 162 102 163
rect 100 162 101 163
rect 99 162 100 163
rect 98 162 99 163
rect 97 162 98 163
rect 96 162 97 163
rect 95 162 96 163
rect 94 162 95 163
rect 93 162 94 163
rect 92 162 93 163
rect 91 162 92 163
rect 90 162 91 163
rect 89 162 90 163
rect 88 162 89 163
rect 87 162 88 163
rect 86 162 87 163
rect 85 162 86 163
rect 84 162 85 163
rect 83 162 84 163
rect 82 162 83 163
rect 81 162 82 163
rect 80 162 81 163
rect 79 162 80 163
rect 78 162 79 163
rect 77 162 78 163
rect 76 162 77 163
rect 75 162 76 163
rect 74 162 75 163
rect 73 162 74 163
rect 72 162 73 163
rect 71 162 72 163
rect 70 162 71 163
rect 69 162 70 163
rect 68 162 69 163
rect 67 162 68 163
rect 66 162 67 163
rect 65 162 66 163
rect 64 162 65 163
rect 63 162 64 163
rect 62 162 63 163
rect 61 162 62 163
rect 60 162 61 163
rect 59 162 60 163
rect 58 162 59 163
rect 57 162 58 163
rect 56 162 57 163
rect 55 162 56 163
rect 54 162 55 163
rect 53 162 54 163
rect 52 162 53 163
rect 51 162 52 163
rect 50 162 51 163
rect 49 162 50 163
rect 48 162 49 163
rect 47 162 48 163
rect 46 162 47 163
rect 45 162 46 163
rect 44 162 45 163
rect 43 162 44 163
rect 42 162 43 163
rect 41 162 42 163
rect 40 162 41 163
rect 39 162 40 163
rect 38 162 39 163
rect 37 162 38 163
rect 36 162 37 163
rect 27 162 28 163
rect 26 162 27 163
rect 25 162 26 163
rect 24 162 25 163
rect 23 162 24 163
rect 22 162 23 163
rect 21 162 22 163
rect 20 162 21 163
rect 19 162 20 163
rect 18 162 19 163
rect 17 162 18 163
rect 16 162 17 163
rect 15 162 16 163
rect 14 162 15 163
rect 13 162 14 163
rect 12 162 13 163
rect 11 162 12 163
rect 10 162 11 163
rect 9 162 10 163
rect 462 163 463 164
rect 441 163 442 164
rect 440 163 441 164
rect 439 163 440 164
rect 438 163 439 164
rect 437 163 438 164
rect 436 163 437 164
rect 435 163 436 164
rect 434 163 435 164
rect 433 163 434 164
rect 432 163 433 164
rect 431 163 432 164
rect 430 163 431 164
rect 429 163 430 164
rect 428 163 429 164
rect 427 163 428 164
rect 426 163 427 164
rect 425 163 426 164
rect 424 163 425 164
rect 423 163 424 164
rect 422 163 423 164
rect 421 163 422 164
rect 420 163 421 164
rect 419 163 420 164
rect 418 163 419 164
rect 417 163 418 164
rect 416 163 417 164
rect 415 163 416 164
rect 414 163 415 164
rect 413 163 414 164
rect 412 163 413 164
rect 411 163 412 164
rect 410 163 411 164
rect 409 163 410 164
rect 408 163 409 164
rect 407 163 408 164
rect 406 163 407 164
rect 405 163 406 164
rect 404 163 405 164
rect 403 163 404 164
rect 402 163 403 164
rect 401 163 402 164
rect 400 163 401 164
rect 399 163 400 164
rect 398 163 399 164
rect 397 163 398 164
rect 288 163 289 164
rect 287 163 288 164
rect 286 163 287 164
rect 285 163 286 164
rect 284 163 285 164
rect 283 163 284 164
rect 282 163 283 164
rect 281 163 282 164
rect 280 163 281 164
rect 279 163 280 164
rect 278 163 279 164
rect 277 163 278 164
rect 276 163 277 164
rect 275 163 276 164
rect 274 163 275 164
rect 273 163 274 164
rect 272 163 273 164
rect 271 163 272 164
rect 270 163 271 164
rect 269 163 270 164
rect 268 163 269 164
rect 267 163 268 164
rect 266 163 267 164
rect 265 163 266 164
rect 264 163 265 164
rect 263 163 264 164
rect 262 163 263 164
rect 261 163 262 164
rect 260 163 261 164
rect 259 163 260 164
rect 258 163 259 164
rect 257 163 258 164
rect 256 163 257 164
rect 255 163 256 164
rect 254 163 255 164
rect 253 163 254 164
rect 252 163 253 164
rect 251 163 252 164
rect 250 163 251 164
rect 249 163 250 164
rect 248 163 249 164
rect 247 163 248 164
rect 246 163 247 164
rect 245 163 246 164
rect 244 163 245 164
rect 243 163 244 164
rect 242 163 243 164
rect 241 163 242 164
rect 240 163 241 164
rect 239 163 240 164
rect 238 163 239 164
rect 237 163 238 164
rect 236 163 237 164
rect 235 163 236 164
rect 234 163 235 164
rect 215 163 216 164
rect 214 163 215 164
rect 213 163 214 164
rect 212 163 213 164
rect 211 163 212 164
rect 210 163 211 164
rect 209 163 210 164
rect 208 163 209 164
rect 207 163 208 164
rect 206 163 207 164
rect 205 163 206 164
rect 204 163 205 164
rect 203 163 204 164
rect 202 163 203 164
rect 201 163 202 164
rect 200 163 201 164
rect 199 163 200 164
rect 198 163 199 164
rect 197 163 198 164
rect 196 163 197 164
rect 195 163 196 164
rect 194 163 195 164
rect 193 163 194 164
rect 192 163 193 164
rect 191 163 192 164
rect 190 163 191 164
rect 189 163 190 164
rect 188 163 189 164
rect 187 163 188 164
rect 186 163 187 164
rect 185 163 186 164
rect 184 163 185 164
rect 183 163 184 164
rect 182 163 183 164
rect 181 163 182 164
rect 180 163 181 164
rect 179 163 180 164
rect 178 163 179 164
rect 177 163 178 164
rect 176 163 177 164
rect 175 163 176 164
rect 174 163 175 164
rect 173 163 174 164
rect 172 163 173 164
rect 171 163 172 164
rect 170 163 171 164
rect 169 163 170 164
rect 168 163 169 164
rect 167 163 168 164
rect 166 163 167 164
rect 165 163 166 164
rect 164 163 165 164
rect 163 163 164 164
rect 162 163 163 164
rect 161 163 162 164
rect 160 163 161 164
rect 159 163 160 164
rect 158 163 159 164
rect 157 163 158 164
rect 156 163 157 164
rect 155 163 156 164
rect 154 163 155 164
rect 153 163 154 164
rect 152 163 153 164
rect 151 163 152 164
rect 150 163 151 164
rect 149 163 150 164
rect 148 163 149 164
rect 147 163 148 164
rect 113 163 114 164
rect 112 163 113 164
rect 111 163 112 164
rect 110 163 111 164
rect 109 163 110 164
rect 108 163 109 164
rect 107 163 108 164
rect 106 163 107 164
rect 105 163 106 164
rect 104 163 105 164
rect 103 163 104 164
rect 102 163 103 164
rect 101 163 102 164
rect 100 163 101 164
rect 99 163 100 164
rect 98 163 99 164
rect 97 163 98 164
rect 96 163 97 164
rect 95 163 96 164
rect 94 163 95 164
rect 93 163 94 164
rect 92 163 93 164
rect 91 163 92 164
rect 90 163 91 164
rect 89 163 90 164
rect 88 163 89 164
rect 87 163 88 164
rect 86 163 87 164
rect 85 163 86 164
rect 84 163 85 164
rect 83 163 84 164
rect 82 163 83 164
rect 81 163 82 164
rect 80 163 81 164
rect 79 163 80 164
rect 78 163 79 164
rect 77 163 78 164
rect 76 163 77 164
rect 75 163 76 164
rect 74 163 75 164
rect 73 163 74 164
rect 72 163 73 164
rect 71 163 72 164
rect 70 163 71 164
rect 69 163 70 164
rect 68 163 69 164
rect 67 163 68 164
rect 66 163 67 164
rect 65 163 66 164
rect 64 163 65 164
rect 63 163 64 164
rect 62 163 63 164
rect 61 163 62 164
rect 60 163 61 164
rect 59 163 60 164
rect 58 163 59 164
rect 57 163 58 164
rect 56 163 57 164
rect 55 163 56 164
rect 54 163 55 164
rect 53 163 54 164
rect 52 163 53 164
rect 51 163 52 164
rect 50 163 51 164
rect 49 163 50 164
rect 48 163 49 164
rect 47 163 48 164
rect 46 163 47 164
rect 45 163 46 164
rect 44 163 45 164
rect 43 163 44 164
rect 42 163 43 164
rect 41 163 42 164
rect 40 163 41 164
rect 39 163 40 164
rect 38 163 39 164
rect 37 163 38 164
rect 36 163 37 164
rect 26 163 27 164
rect 25 163 26 164
rect 24 163 25 164
rect 23 163 24 164
rect 22 163 23 164
rect 21 163 22 164
rect 20 163 21 164
rect 19 163 20 164
rect 18 163 19 164
rect 17 163 18 164
rect 16 163 17 164
rect 15 163 16 164
rect 14 163 15 164
rect 13 163 14 164
rect 12 163 13 164
rect 11 163 12 164
rect 10 163 11 164
rect 463 164 464 165
rect 462 164 463 165
rect 441 164 442 165
rect 440 164 441 165
rect 439 164 440 165
rect 438 164 439 165
rect 437 164 438 165
rect 436 164 437 165
rect 435 164 436 165
rect 434 164 435 165
rect 433 164 434 165
rect 432 164 433 165
rect 431 164 432 165
rect 430 164 431 165
rect 429 164 430 165
rect 428 164 429 165
rect 427 164 428 165
rect 426 164 427 165
rect 425 164 426 165
rect 424 164 425 165
rect 423 164 424 165
rect 422 164 423 165
rect 421 164 422 165
rect 420 164 421 165
rect 419 164 420 165
rect 418 164 419 165
rect 417 164 418 165
rect 416 164 417 165
rect 415 164 416 165
rect 414 164 415 165
rect 413 164 414 165
rect 412 164 413 165
rect 411 164 412 165
rect 410 164 411 165
rect 409 164 410 165
rect 408 164 409 165
rect 407 164 408 165
rect 406 164 407 165
rect 405 164 406 165
rect 404 164 405 165
rect 403 164 404 165
rect 402 164 403 165
rect 401 164 402 165
rect 400 164 401 165
rect 399 164 400 165
rect 398 164 399 165
rect 397 164 398 165
rect 286 164 287 165
rect 285 164 286 165
rect 284 164 285 165
rect 283 164 284 165
rect 282 164 283 165
rect 281 164 282 165
rect 280 164 281 165
rect 279 164 280 165
rect 278 164 279 165
rect 277 164 278 165
rect 276 164 277 165
rect 275 164 276 165
rect 274 164 275 165
rect 273 164 274 165
rect 272 164 273 165
rect 271 164 272 165
rect 270 164 271 165
rect 269 164 270 165
rect 268 164 269 165
rect 267 164 268 165
rect 266 164 267 165
rect 265 164 266 165
rect 264 164 265 165
rect 263 164 264 165
rect 262 164 263 165
rect 261 164 262 165
rect 260 164 261 165
rect 259 164 260 165
rect 258 164 259 165
rect 257 164 258 165
rect 256 164 257 165
rect 255 164 256 165
rect 254 164 255 165
rect 253 164 254 165
rect 252 164 253 165
rect 251 164 252 165
rect 250 164 251 165
rect 249 164 250 165
rect 248 164 249 165
rect 247 164 248 165
rect 246 164 247 165
rect 245 164 246 165
rect 244 164 245 165
rect 243 164 244 165
rect 242 164 243 165
rect 241 164 242 165
rect 240 164 241 165
rect 239 164 240 165
rect 238 164 239 165
rect 237 164 238 165
rect 236 164 237 165
rect 235 164 236 165
rect 234 164 235 165
rect 215 164 216 165
rect 214 164 215 165
rect 213 164 214 165
rect 212 164 213 165
rect 211 164 212 165
rect 210 164 211 165
rect 209 164 210 165
rect 208 164 209 165
rect 207 164 208 165
rect 206 164 207 165
rect 205 164 206 165
rect 204 164 205 165
rect 203 164 204 165
rect 202 164 203 165
rect 201 164 202 165
rect 200 164 201 165
rect 199 164 200 165
rect 198 164 199 165
rect 197 164 198 165
rect 196 164 197 165
rect 195 164 196 165
rect 194 164 195 165
rect 193 164 194 165
rect 192 164 193 165
rect 191 164 192 165
rect 190 164 191 165
rect 189 164 190 165
rect 188 164 189 165
rect 187 164 188 165
rect 186 164 187 165
rect 185 164 186 165
rect 184 164 185 165
rect 183 164 184 165
rect 182 164 183 165
rect 181 164 182 165
rect 180 164 181 165
rect 179 164 180 165
rect 178 164 179 165
rect 177 164 178 165
rect 176 164 177 165
rect 175 164 176 165
rect 174 164 175 165
rect 173 164 174 165
rect 172 164 173 165
rect 171 164 172 165
rect 170 164 171 165
rect 169 164 170 165
rect 168 164 169 165
rect 167 164 168 165
rect 166 164 167 165
rect 165 164 166 165
rect 164 164 165 165
rect 163 164 164 165
rect 162 164 163 165
rect 161 164 162 165
rect 160 164 161 165
rect 159 164 160 165
rect 158 164 159 165
rect 157 164 158 165
rect 156 164 157 165
rect 155 164 156 165
rect 154 164 155 165
rect 153 164 154 165
rect 152 164 153 165
rect 151 164 152 165
rect 150 164 151 165
rect 149 164 150 165
rect 148 164 149 165
rect 147 164 148 165
rect 146 164 147 165
rect 145 164 146 165
rect 111 164 112 165
rect 110 164 111 165
rect 109 164 110 165
rect 108 164 109 165
rect 107 164 108 165
rect 106 164 107 165
rect 105 164 106 165
rect 104 164 105 165
rect 103 164 104 165
rect 102 164 103 165
rect 101 164 102 165
rect 100 164 101 165
rect 99 164 100 165
rect 98 164 99 165
rect 97 164 98 165
rect 96 164 97 165
rect 95 164 96 165
rect 94 164 95 165
rect 93 164 94 165
rect 92 164 93 165
rect 91 164 92 165
rect 90 164 91 165
rect 89 164 90 165
rect 88 164 89 165
rect 87 164 88 165
rect 86 164 87 165
rect 85 164 86 165
rect 84 164 85 165
rect 83 164 84 165
rect 82 164 83 165
rect 81 164 82 165
rect 80 164 81 165
rect 79 164 80 165
rect 78 164 79 165
rect 77 164 78 165
rect 76 164 77 165
rect 75 164 76 165
rect 74 164 75 165
rect 73 164 74 165
rect 72 164 73 165
rect 71 164 72 165
rect 70 164 71 165
rect 69 164 70 165
rect 68 164 69 165
rect 67 164 68 165
rect 66 164 67 165
rect 65 164 66 165
rect 64 164 65 165
rect 63 164 64 165
rect 62 164 63 165
rect 61 164 62 165
rect 60 164 61 165
rect 59 164 60 165
rect 58 164 59 165
rect 57 164 58 165
rect 56 164 57 165
rect 55 164 56 165
rect 54 164 55 165
rect 53 164 54 165
rect 52 164 53 165
rect 51 164 52 165
rect 50 164 51 165
rect 49 164 50 165
rect 48 164 49 165
rect 47 164 48 165
rect 46 164 47 165
rect 45 164 46 165
rect 44 164 45 165
rect 43 164 44 165
rect 42 164 43 165
rect 41 164 42 165
rect 40 164 41 165
rect 39 164 40 165
rect 38 164 39 165
rect 37 164 38 165
rect 36 164 37 165
rect 26 164 27 165
rect 25 164 26 165
rect 24 164 25 165
rect 23 164 24 165
rect 22 164 23 165
rect 21 164 22 165
rect 20 164 21 165
rect 19 164 20 165
rect 18 164 19 165
rect 17 164 18 165
rect 16 164 17 165
rect 15 164 16 165
rect 14 164 15 165
rect 13 164 14 165
rect 12 164 13 165
rect 11 164 12 165
rect 10 164 11 165
rect 465 165 466 166
rect 464 165 465 166
rect 463 165 464 166
rect 462 165 463 166
rect 441 165 442 166
rect 440 165 441 166
rect 439 165 440 166
rect 438 165 439 166
rect 437 165 438 166
rect 436 165 437 166
rect 435 165 436 166
rect 434 165 435 166
rect 433 165 434 166
rect 432 165 433 166
rect 431 165 432 166
rect 430 165 431 166
rect 429 165 430 166
rect 428 165 429 166
rect 427 165 428 166
rect 426 165 427 166
rect 425 165 426 166
rect 424 165 425 166
rect 423 165 424 166
rect 422 165 423 166
rect 421 165 422 166
rect 420 165 421 166
rect 419 165 420 166
rect 418 165 419 166
rect 417 165 418 166
rect 416 165 417 166
rect 415 165 416 166
rect 414 165 415 166
rect 413 165 414 166
rect 412 165 413 166
rect 411 165 412 166
rect 410 165 411 166
rect 409 165 410 166
rect 408 165 409 166
rect 407 165 408 166
rect 406 165 407 166
rect 405 165 406 166
rect 404 165 405 166
rect 403 165 404 166
rect 402 165 403 166
rect 401 165 402 166
rect 400 165 401 166
rect 399 165 400 166
rect 398 165 399 166
rect 397 165 398 166
rect 284 165 285 166
rect 283 165 284 166
rect 282 165 283 166
rect 281 165 282 166
rect 280 165 281 166
rect 279 165 280 166
rect 278 165 279 166
rect 277 165 278 166
rect 276 165 277 166
rect 275 165 276 166
rect 274 165 275 166
rect 273 165 274 166
rect 272 165 273 166
rect 271 165 272 166
rect 270 165 271 166
rect 269 165 270 166
rect 268 165 269 166
rect 267 165 268 166
rect 266 165 267 166
rect 265 165 266 166
rect 264 165 265 166
rect 263 165 264 166
rect 262 165 263 166
rect 261 165 262 166
rect 260 165 261 166
rect 259 165 260 166
rect 258 165 259 166
rect 257 165 258 166
rect 256 165 257 166
rect 255 165 256 166
rect 254 165 255 166
rect 253 165 254 166
rect 252 165 253 166
rect 251 165 252 166
rect 250 165 251 166
rect 249 165 250 166
rect 248 165 249 166
rect 247 165 248 166
rect 246 165 247 166
rect 245 165 246 166
rect 244 165 245 166
rect 243 165 244 166
rect 242 165 243 166
rect 241 165 242 166
rect 240 165 241 166
rect 239 165 240 166
rect 238 165 239 166
rect 237 165 238 166
rect 236 165 237 166
rect 235 165 236 166
rect 234 165 235 166
rect 233 165 234 166
rect 215 165 216 166
rect 214 165 215 166
rect 213 165 214 166
rect 212 165 213 166
rect 211 165 212 166
rect 210 165 211 166
rect 209 165 210 166
rect 208 165 209 166
rect 207 165 208 166
rect 206 165 207 166
rect 205 165 206 166
rect 204 165 205 166
rect 203 165 204 166
rect 202 165 203 166
rect 201 165 202 166
rect 200 165 201 166
rect 199 165 200 166
rect 198 165 199 166
rect 197 165 198 166
rect 196 165 197 166
rect 195 165 196 166
rect 194 165 195 166
rect 193 165 194 166
rect 192 165 193 166
rect 191 165 192 166
rect 190 165 191 166
rect 189 165 190 166
rect 188 165 189 166
rect 187 165 188 166
rect 186 165 187 166
rect 185 165 186 166
rect 184 165 185 166
rect 183 165 184 166
rect 182 165 183 166
rect 181 165 182 166
rect 180 165 181 166
rect 179 165 180 166
rect 178 165 179 166
rect 177 165 178 166
rect 176 165 177 166
rect 175 165 176 166
rect 174 165 175 166
rect 173 165 174 166
rect 172 165 173 166
rect 171 165 172 166
rect 170 165 171 166
rect 169 165 170 166
rect 168 165 169 166
rect 167 165 168 166
rect 166 165 167 166
rect 165 165 166 166
rect 164 165 165 166
rect 163 165 164 166
rect 162 165 163 166
rect 161 165 162 166
rect 160 165 161 166
rect 159 165 160 166
rect 158 165 159 166
rect 157 165 158 166
rect 156 165 157 166
rect 155 165 156 166
rect 154 165 155 166
rect 153 165 154 166
rect 152 165 153 166
rect 151 165 152 166
rect 150 165 151 166
rect 149 165 150 166
rect 148 165 149 166
rect 147 165 148 166
rect 146 165 147 166
rect 145 165 146 166
rect 144 165 145 166
rect 110 165 111 166
rect 109 165 110 166
rect 108 165 109 166
rect 107 165 108 166
rect 106 165 107 166
rect 105 165 106 166
rect 104 165 105 166
rect 103 165 104 166
rect 102 165 103 166
rect 101 165 102 166
rect 100 165 101 166
rect 99 165 100 166
rect 98 165 99 166
rect 97 165 98 166
rect 96 165 97 166
rect 95 165 96 166
rect 94 165 95 166
rect 93 165 94 166
rect 92 165 93 166
rect 91 165 92 166
rect 90 165 91 166
rect 89 165 90 166
rect 88 165 89 166
rect 87 165 88 166
rect 86 165 87 166
rect 85 165 86 166
rect 84 165 85 166
rect 83 165 84 166
rect 82 165 83 166
rect 81 165 82 166
rect 80 165 81 166
rect 79 165 80 166
rect 78 165 79 166
rect 77 165 78 166
rect 76 165 77 166
rect 75 165 76 166
rect 74 165 75 166
rect 73 165 74 166
rect 72 165 73 166
rect 71 165 72 166
rect 70 165 71 166
rect 69 165 70 166
rect 68 165 69 166
rect 67 165 68 166
rect 66 165 67 166
rect 65 165 66 166
rect 64 165 65 166
rect 63 165 64 166
rect 62 165 63 166
rect 61 165 62 166
rect 60 165 61 166
rect 59 165 60 166
rect 58 165 59 166
rect 57 165 58 166
rect 56 165 57 166
rect 55 165 56 166
rect 54 165 55 166
rect 53 165 54 166
rect 52 165 53 166
rect 51 165 52 166
rect 50 165 51 166
rect 49 165 50 166
rect 48 165 49 166
rect 47 165 48 166
rect 46 165 47 166
rect 45 165 46 166
rect 44 165 45 166
rect 43 165 44 166
rect 42 165 43 166
rect 41 165 42 166
rect 40 165 41 166
rect 39 165 40 166
rect 38 165 39 166
rect 37 165 38 166
rect 36 165 37 166
rect 35 165 36 166
rect 26 165 27 166
rect 25 165 26 166
rect 24 165 25 166
rect 23 165 24 166
rect 22 165 23 166
rect 21 165 22 166
rect 20 165 21 166
rect 19 165 20 166
rect 18 165 19 166
rect 17 165 18 166
rect 16 165 17 166
rect 15 165 16 166
rect 14 165 15 166
rect 13 165 14 166
rect 12 165 13 166
rect 11 165 12 166
rect 10 165 11 166
rect 467 166 468 167
rect 466 166 467 167
rect 465 166 466 167
rect 464 166 465 167
rect 463 166 464 167
rect 462 166 463 167
rect 441 166 442 167
rect 440 166 441 167
rect 439 166 440 167
rect 438 166 439 167
rect 437 166 438 167
rect 436 166 437 167
rect 435 166 436 167
rect 434 166 435 167
rect 433 166 434 167
rect 432 166 433 167
rect 431 166 432 167
rect 430 166 431 167
rect 429 166 430 167
rect 428 166 429 167
rect 427 166 428 167
rect 426 166 427 167
rect 425 166 426 167
rect 424 166 425 167
rect 423 166 424 167
rect 422 166 423 167
rect 421 166 422 167
rect 420 166 421 167
rect 419 166 420 167
rect 418 166 419 167
rect 417 166 418 167
rect 416 166 417 167
rect 415 166 416 167
rect 414 166 415 167
rect 413 166 414 167
rect 412 166 413 167
rect 411 166 412 167
rect 410 166 411 167
rect 409 166 410 167
rect 408 166 409 167
rect 407 166 408 167
rect 406 166 407 167
rect 405 166 406 167
rect 404 166 405 167
rect 403 166 404 167
rect 402 166 403 167
rect 401 166 402 167
rect 400 166 401 167
rect 399 166 400 167
rect 398 166 399 167
rect 397 166 398 167
rect 282 166 283 167
rect 281 166 282 167
rect 280 166 281 167
rect 279 166 280 167
rect 278 166 279 167
rect 277 166 278 167
rect 276 166 277 167
rect 275 166 276 167
rect 274 166 275 167
rect 273 166 274 167
rect 272 166 273 167
rect 271 166 272 167
rect 270 166 271 167
rect 269 166 270 167
rect 268 166 269 167
rect 267 166 268 167
rect 266 166 267 167
rect 265 166 266 167
rect 264 166 265 167
rect 263 166 264 167
rect 262 166 263 167
rect 261 166 262 167
rect 260 166 261 167
rect 259 166 260 167
rect 258 166 259 167
rect 257 166 258 167
rect 256 166 257 167
rect 255 166 256 167
rect 254 166 255 167
rect 253 166 254 167
rect 252 166 253 167
rect 251 166 252 167
rect 250 166 251 167
rect 249 166 250 167
rect 248 166 249 167
rect 247 166 248 167
rect 246 166 247 167
rect 245 166 246 167
rect 244 166 245 167
rect 243 166 244 167
rect 242 166 243 167
rect 241 166 242 167
rect 240 166 241 167
rect 239 166 240 167
rect 238 166 239 167
rect 237 166 238 167
rect 236 166 237 167
rect 235 166 236 167
rect 234 166 235 167
rect 233 166 234 167
rect 214 166 215 167
rect 213 166 214 167
rect 212 166 213 167
rect 211 166 212 167
rect 210 166 211 167
rect 209 166 210 167
rect 208 166 209 167
rect 207 166 208 167
rect 206 166 207 167
rect 205 166 206 167
rect 204 166 205 167
rect 203 166 204 167
rect 202 166 203 167
rect 201 166 202 167
rect 200 166 201 167
rect 199 166 200 167
rect 198 166 199 167
rect 197 166 198 167
rect 196 166 197 167
rect 195 166 196 167
rect 194 166 195 167
rect 193 166 194 167
rect 192 166 193 167
rect 191 166 192 167
rect 190 166 191 167
rect 189 166 190 167
rect 188 166 189 167
rect 187 166 188 167
rect 186 166 187 167
rect 185 166 186 167
rect 184 166 185 167
rect 183 166 184 167
rect 182 166 183 167
rect 181 166 182 167
rect 180 166 181 167
rect 179 166 180 167
rect 178 166 179 167
rect 177 166 178 167
rect 176 166 177 167
rect 175 166 176 167
rect 174 166 175 167
rect 173 166 174 167
rect 172 166 173 167
rect 171 166 172 167
rect 170 166 171 167
rect 169 166 170 167
rect 168 166 169 167
rect 167 166 168 167
rect 166 166 167 167
rect 165 166 166 167
rect 164 166 165 167
rect 163 166 164 167
rect 162 166 163 167
rect 161 166 162 167
rect 160 166 161 167
rect 159 166 160 167
rect 158 166 159 167
rect 157 166 158 167
rect 156 166 157 167
rect 155 166 156 167
rect 154 166 155 167
rect 153 166 154 167
rect 152 166 153 167
rect 151 166 152 167
rect 150 166 151 167
rect 149 166 150 167
rect 148 166 149 167
rect 147 166 148 167
rect 146 166 147 167
rect 145 166 146 167
rect 144 166 145 167
rect 143 166 144 167
rect 108 166 109 167
rect 107 166 108 167
rect 106 166 107 167
rect 105 166 106 167
rect 104 166 105 167
rect 103 166 104 167
rect 102 166 103 167
rect 101 166 102 167
rect 100 166 101 167
rect 99 166 100 167
rect 98 166 99 167
rect 97 166 98 167
rect 96 166 97 167
rect 95 166 96 167
rect 94 166 95 167
rect 93 166 94 167
rect 92 166 93 167
rect 91 166 92 167
rect 90 166 91 167
rect 89 166 90 167
rect 88 166 89 167
rect 87 166 88 167
rect 86 166 87 167
rect 85 166 86 167
rect 84 166 85 167
rect 83 166 84 167
rect 82 166 83 167
rect 81 166 82 167
rect 80 166 81 167
rect 79 166 80 167
rect 78 166 79 167
rect 77 166 78 167
rect 76 166 77 167
rect 75 166 76 167
rect 70 166 71 167
rect 69 166 70 167
rect 68 166 69 167
rect 67 166 68 167
rect 66 166 67 167
rect 65 166 66 167
rect 64 166 65 167
rect 63 166 64 167
rect 62 166 63 167
rect 61 166 62 167
rect 60 166 61 167
rect 59 166 60 167
rect 58 166 59 167
rect 57 166 58 167
rect 56 166 57 167
rect 55 166 56 167
rect 54 166 55 167
rect 53 166 54 167
rect 52 166 53 167
rect 51 166 52 167
rect 50 166 51 167
rect 49 166 50 167
rect 48 166 49 167
rect 47 166 48 167
rect 46 166 47 167
rect 45 166 46 167
rect 44 166 45 167
rect 43 166 44 167
rect 42 166 43 167
rect 41 166 42 167
rect 40 166 41 167
rect 39 166 40 167
rect 38 166 39 167
rect 37 166 38 167
rect 36 166 37 167
rect 35 166 36 167
rect 25 166 26 167
rect 24 166 25 167
rect 23 166 24 167
rect 22 166 23 167
rect 21 166 22 167
rect 20 166 21 167
rect 19 166 20 167
rect 18 166 19 167
rect 17 166 18 167
rect 16 166 17 167
rect 15 166 16 167
rect 14 166 15 167
rect 13 166 14 167
rect 12 166 13 167
rect 11 166 12 167
rect 10 166 11 167
rect 470 167 471 168
rect 469 167 470 168
rect 468 167 469 168
rect 467 167 468 168
rect 466 167 467 168
rect 465 167 466 168
rect 464 167 465 168
rect 463 167 464 168
rect 462 167 463 168
rect 441 167 442 168
rect 440 167 441 168
rect 439 167 440 168
rect 438 167 439 168
rect 437 167 438 168
rect 436 167 437 168
rect 435 167 436 168
rect 408 167 409 168
rect 407 167 408 168
rect 406 167 407 168
rect 405 167 406 168
rect 404 167 405 168
rect 403 167 404 168
rect 402 167 403 168
rect 401 167 402 168
rect 400 167 401 168
rect 399 167 400 168
rect 398 167 399 168
rect 397 167 398 168
rect 281 167 282 168
rect 280 167 281 168
rect 279 167 280 168
rect 278 167 279 168
rect 277 167 278 168
rect 276 167 277 168
rect 275 167 276 168
rect 274 167 275 168
rect 273 167 274 168
rect 272 167 273 168
rect 271 167 272 168
rect 270 167 271 168
rect 269 167 270 168
rect 268 167 269 168
rect 267 167 268 168
rect 266 167 267 168
rect 265 167 266 168
rect 264 167 265 168
rect 263 167 264 168
rect 262 167 263 168
rect 261 167 262 168
rect 260 167 261 168
rect 259 167 260 168
rect 258 167 259 168
rect 257 167 258 168
rect 256 167 257 168
rect 255 167 256 168
rect 254 167 255 168
rect 253 167 254 168
rect 252 167 253 168
rect 251 167 252 168
rect 250 167 251 168
rect 249 167 250 168
rect 248 167 249 168
rect 247 167 248 168
rect 246 167 247 168
rect 245 167 246 168
rect 244 167 245 168
rect 243 167 244 168
rect 242 167 243 168
rect 241 167 242 168
rect 240 167 241 168
rect 239 167 240 168
rect 238 167 239 168
rect 237 167 238 168
rect 236 167 237 168
rect 235 167 236 168
rect 234 167 235 168
rect 233 167 234 168
rect 232 167 233 168
rect 213 167 214 168
rect 212 167 213 168
rect 211 167 212 168
rect 210 167 211 168
rect 209 167 210 168
rect 208 167 209 168
rect 207 167 208 168
rect 206 167 207 168
rect 205 167 206 168
rect 204 167 205 168
rect 203 167 204 168
rect 202 167 203 168
rect 201 167 202 168
rect 200 167 201 168
rect 199 167 200 168
rect 198 167 199 168
rect 197 167 198 168
rect 196 167 197 168
rect 195 167 196 168
rect 194 167 195 168
rect 193 167 194 168
rect 192 167 193 168
rect 191 167 192 168
rect 190 167 191 168
rect 189 167 190 168
rect 188 167 189 168
rect 187 167 188 168
rect 186 167 187 168
rect 185 167 186 168
rect 184 167 185 168
rect 183 167 184 168
rect 182 167 183 168
rect 181 167 182 168
rect 180 167 181 168
rect 179 167 180 168
rect 178 167 179 168
rect 177 167 178 168
rect 176 167 177 168
rect 175 167 176 168
rect 174 167 175 168
rect 173 167 174 168
rect 172 167 173 168
rect 171 167 172 168
rect 170 167 171 168
rect 169 167 170 168
rect 168 167 169 168
rect 167 167 168 168
rect 166 167 167 168
rect 165 167 166 168
rect 164 167 165 168
rect 163 167 164 168
rect 162 167 163 168
rect 161 167 162 168
rect 160 167 161 168
rect 159 167 160 168
rect 158 167 159 168
rect 157 167 158 168
rect 156 167 157 168
rect 155 167 156 168
rect 154 167 155 168
rect 153 167 154 168
rect 152 167 153 168
rect 151 167 152 168
rect 150 167 151 168
rect 149 167 150 168
rect 148 167 149 168
rect 147 167 148 168
rect 146 167 147 168
rect 145 167 146 168
rect 144 167 145 168
rect 143 167 144 168
rect 142 167 143 168
rect 106 167 107 168
rect 105 167 106 168
rect 104 167 105 168
rect 103 167 104 168
rect 102 167 103 168
rect 101 167 102 168
rect 100 167 101 168
rect 99 167 100 168
rect 98 167 99 168
rect 97 167 98 168
rect 96 167 97 168
rect 95 167 96 168
rect 94 167 95 168
rect 93 167 94 168
rect 92 167 93 168
rect 91 167 92 168
rect 90 167 91 168
rect 89 167 90 168
rect 88 167 89 168
rect 87 167 88 168
rect 86 167 87 168
rect 85 167 86 168
rect 84 167 85 168
rect 83 167 84 168
rect 82 167 83 168
rect 81 167 82 168
rect 80 167 81 168
rect 68 167 69 168
rect 67 167 68 168
rect 66 167 67 168
rect 65 167 66 168
rect 64 167 65 168
rect 63 167 64 168
rect 62 167 63 168
rect 61 167 62 168
rect 60 167 61 168
rect 59 167 60 168
rect 58 167 59 168
rect 57 167 58 168
rect 56 167 57 168
rect 55 167 56 168
rect 54 167 55 168
rect 53 167 54 168
rect 52 167 53 168
rect 51 167 52 168
rect 50 167 51 168
rect 49 167 50 168
rect 48 167 49 168
rect 47 167 48 168
rect 46 167 47 168
rect 45 167 46 168
rect 44 167 45 168
rect 43 167 44 168
rect 42 167 43 168
rect 41 167 42 168
rect 40 167 41 168
rect 39 167 40 168
rect 38 167 39 168
rect 37 167 38 168
rect 36 167 37 168
rect 35 167 36 168
rect 25 167 26 168
rect 24 167 25 168
rect 23 167 24 168
rect 22 167 23 168
rect 21 167 22 168
rect 20 167 21 168
rect 19 167 20 168
rect 18 167 19 168
rect 17 167 18 168
rect 16 167 17 168
rect 15 167 16 168
rect 14 167 15 168
rect 13 167 14 168
rect 12 167 13 168
rect 11 167 12 168
rect 10 167 11 168
rect 472 168 473 169
rect 471 168 472 169
rect 470 168 471 169
rect 469 168 470 169
rect 468 168 469 169
rect 467 168 468 169
rect 466 168 467 169
rect 465 168 466 169
rect 464 168 465 169
rect 463 168 464 169
rect 462 168 463 169
rect 441 168 442 169
rect 440 168 441 169
rect 439 168 440 169
rect 438 168 439 169
rect 409 168 410 169
rect 408 168 409 169
rect 407 168 408 169
rect 406 168 407 169
rect 405 168 406 169
rect 404 168 405 169
rect 403 168 404 169
rect 402 168 403 169
rect 401 168 402 169
rect 400 168 401 169
rect 399 168 400 169
rect 398 168 399 169
rect 397 168 398 169
rect 279 168 280 169
rect 278 168 279 169
rect 277 168 278 169
rect 276 168 277 169
rect 275 168 276 169
rect 274 168 275 169
rect 273 168 274 169
rect 272 168 273 169
rect 271 168 272 169
rect 270 168 271 169
rect 269 168 270 169
rect 268 168 269 169
rect 267 168 268 169
rect 266 168 267 169
rect 265 168 266 169
rect 264 168 265 169
rect 263 168 264 169
rect 262 168 263 169
rect 261 168 262 169
rect 260 168 261 169
rect 259 168 260 169
rect 258 168 259 169
rect 257 168 258 169
rect 256 168 257 169
rect 255 168 256 169
rect 254 168 255 169
rect 253 168 254 169
rect 252 168 253 169
rect 251 168 252 169
rect 250 168 251 169
rect 249 168 250 169
rect 248 168 249 169
rect 247 168 248 169
rect 246 168 247 169
rect 245 168 246 169
rect 244 168 245 169
rect 243 168 244 169
rect 242 168 243 169
rect 241 168 242 169
rect 240 168 241 169
rect 239 168 240 169
rect 238 168 239 169
rect 237 168 238 169
rect 236 168 237 169
rect 235 168 236 169
rect 234 168 235 169
rect 233 168 234 169
rect 232 168 233 169
rect 213 168 214 169
rect 212 168 213 169
rect 211 168 212 169
rect 210 168 211 169
rect 209 168 210 169
rect 208 168 209 169
rect 207 168 208 169
rect 206 168 207 169
rect 205 168 206 169
rect 204 168 205 169
rect 203 168 204 169
rect 202 168 203 169
rect 201 168 202 169
rect 200 168 201 169
rect 199 168 200 169
rect 198 168 199 169
rect 197 168 198 169
rect 196 168 197 169
rect 195 168 196 169
rect 194 168 195 169
rect 193 168 194 169
rect 192 168 193 169
rect 191 168 192 169
rect 190 168 191 169
rect 189 168 190 169
rect 188 168 189 169
rect 187 168 188 169
rect 186 168 187 169
rect 185 168 186 169
rect 184 168 185 169
rect 183 168 184 169
rect 182 168 183 169
rect 181 168 182 169
rect 180 168 181 169
rect 179 168 180 169
rect 178 168 179 169
rect 177 168 178 169
rect 176 168 177 169
rect 175 168 176 169
rect 174 168 175 169
rect 173 168 174 169
rect 172 168 173 169
rect 171 168 172 169
rect 170 168 171 169
rect 169 168 170 169
rect 168 168 169 169
rect 167 168 168 169
rect 166 168 167 169
rect 165 168 166 169
rect 164 168 165 169
rect 163 168 164 169
rect 162 168 163 169
rect 161 168 162 169
rect 160 168 161 169
rect 159 168 160 169
rect 158 168 159 169
rect 157 168 158 169
rect 156 168 157 169
rect 155 168 156 169
rect 154 168 155 169
rect 153 168 154 169
rect 152 168 153 169
rect 151 168 152 169
rect 150 168 151 169
rect 149 168 150 169
rect 148 168 149 169
rect 147 168 148 169
rect 146 168 147 169
rect 145 168 146 169
rect 144 168 145 169
rect 143 168 144 169
rect 142 168 143 169
rect 141 168 142 169
rect 103 168 104 169
rect 102 168 103 169
rect 101 168 102 169
rect 100 168 101 169
rect 99 168 100 169
rect 98 168 99 169
rect 97 168 98 169
rect 96 168 97 169
rect 95 168 96 169
rect 94 168 95 169
rect 93 168 94 169
rect 92 168 93 169
rect 91 168 92 169
rect 90 168 91 169
rect 89 168 90 169
rect 88 168 89 169
rect 87 168 88 169
rect 86 168 87 169
rect 85 168 86 169
rect 84 168 85 169
rect 66 168 67 169
rect 65 168 66 169
rect 64 168 65 169
rect 63 168 64 169
rect 62 168 63 169
rect 61 168 62 169
rect 60 168 61 169
rect 59 168 60 169
rect 58 168 59 169
rect 57 168 58 169
rect 56 168 57 169
rect 55 168 56 169
rect 54 168 55 169
rect 53 168 54 169
rect 52 168 53 169
rect 51 168 52 169
rect 50 168 51 169
rect 49 168 50 169
rect 48 168 49 169
rect 47 168 48 169
rect 46 168 47 169
rect 45 168 46 169
rect 44 168 45 169
rect 43 168 44 169
rect 42 168 43 169
rect 41 168 42 169
rect 40 168 41 169
rect 39 168 40 169
rect 38 168 39 169
rect 37 168 38 169
rect 36 168 37 169
rect 35 168 36 169
rect 25 168 26 169
rect 24 168 25 169
rect 23 168 24 169
rect 22 168 23 169
rect 21 168 22 169
rect 20 168 21 169
rect 19 168 20 169
rect 18 168 19 169
rect 17 168 18 169
rect 16 168 17 169
rect 15 168 16 169
rect 14 168 15 169
rect 13 168 14 169
rect 12 168 13 169
rect 11 168 12 169
rect 10 168 11 169
rect 475 169 476 170
rect 474 169 475 170
rect 473 169 474 170
rect 472 169 473 170
rect 471 169 472 170
rect 470 169 471 170
rect 469 169 470 170
rect 468 169 469 170
rect 467 169 468 170
rect 466 169 467 170
rect 465 169 466 170
rect 464 169 465 170
rect 463 169 464 170
rect 462 169 463 170
rect 441 169 442 170
rect 440 169 441 170
rect 439 169 440 170
rect 411 169 412 170
rect 410 169 411 170
rect 409 169 410 170
rect 408 169 409 170
rect 407 169 408 170
rect 406 169 407 170
rect 405 169 406 170
rect 404 169 405 170
rect 403 169 404 170
rect 402 169 403 170
rect 401 169 402 170
rect 400 169 401 170
rect 399 169 400 170
rect 398 169 399 170
rect 397 169 398 170
rect 278 169 279 170
rect 277 169 278 170
rect 276 169 277 170
rect 275 169 276 170
rect 274 169 275 170
rect 273 169 274 170
rect 272 169 273 170
rect 271 169 272 170
rect 270 169 271 170
rect 269 169 270 170
rect 268 169 269 170
rect 267 169 268 170
rect 266 169 267 170
rect 265 169 266 170
rect 264 169 265 170
rect 263 169 264 170
rect 262 169 263 170
rect 261 169 262 170
rect 260 169 261 170
rect 259 169 260 170
rect 258 169 259 170
rect 257 169 258 170
rect 256 169 257 170
rect 255 169 256 170
rect 254 169 255 170
rect 253 169 254 170
rect 252 169 253 170
rect 251 169 252 170
rect 250 169 251 170
rect 249 169 250 170
rect 248 169 249 170
rect 247 169 248 170
rect 246 169 247 170
rect 245 169 246 170
rect 244 169 245 170
rect 243 169 244 170
rect 242 169 243 170
rect 241 169 242 170
rect 240 169 241 170
rect 239 169 240 170
rect 238 169 239 170
rect 237 169 238 170
rect 236 169 237 170
rect 235 169 236 170
rect 234 169 235 170
rect 233 169 234 170
rect 232 169 233 170
rect 231 169 232 170
rect 212 169 213 170
rect 211 169 212 170
rect 210 169 211 170
rect 209 169 210 170
rect 208 169 209 170
rect 207 169 208 170
rect 206 169 207 170
rect 205 169 206 170
rect 204 169 205 170
rect 203 169 204 170
rect 202 169 203 170
rect 201 169 202 170
rect 200 169 201 170
rect 199 169 200 170
rect 198 169 199 170
rect 197 169 198 170
rect 196 169 197 170
rect 195 169 196 170
rect 194 169 195 170
rect 193 169 194 170
rect 192 169 193 170
rect 191 169 192 170
rect 190 169 191 170
rect 189 169 190 170
rect 188 169 189 170
rect 187 169 188 170
rect 186 169 187 170
rect 185 169 186 170
rect 184 169 185 170
rect 183 169 184 170
rect 182 169 183 170
rect 181 169 182 170
rect 180 169 181 170
rect 179 169 180 170
rect 178 169 179 170
rect 177 169 178 170
rect 176 169 177 170
rect 175 169 176 170
rect 174 169 175 170
rect 173 169 174 170
rect 172 169 173 170
rect 171 169 172 170
rect 170 169 171 170
rect 169 169 170 170
rect 168 169 169 170
rect 167 169 168 170
rect 166 169 167 170
rect 165 169 166 170
rect 164 169 165 170
rect 163 169 164 170
rect 162 169 163 170
rect 161 169 162 170
rect 160 169 161 170
rect 159 169 160 170
rect 158 169 159 170
rect 157 169 158 170
rect 156 169 157 170
rect 155 169 156 170
rect 154 169 155 170
rect 153 169 154 170
rect 152 169 153 170
rect 151 169 152 170
rect 150 169 151 170
rect 149 169 150 170
rect 148 169 149 170
rect 147 169 148 170
rect 146 169 147 170
rect 145 169 146 170
rect 144 169 145 170
rect 143 169 144 170
rect 142 169 143 170
rect 141 169 142 170
rect 140 169 141 170
rect 139 169 140 170
rect 99 169 100 170
rect 98 169 99 170
rect 97 169 98 170
rect 96 169 97 170
rect 95 169 96 170
rect 94 169 95 170
rect 93 169 94 170
rect 92 169 93 170
rect 91 169 92 170
rect 90 169 91 170
rect 65 169 66 170
rect 64 169 65 170
rect 63 169 64 170
rect 62 169 63 170
rect 61 169 62 170
rect 60 169 61 170
rect 59 169 60 170
rect 58 169 59 170
rect 57 169 58 170
rect 56 169 57 170
rect 55 169 56 170
rect 54 169 55 170
rect 53 169 54 170
rect 52 169 53 170
rect 51 169 52 170
rect 50 169 51 170
rect 49 169 50 170
rect 48 169 49 170
rect 47 169 48 170
rect 46 169 47 170
rect 45 169 46 170
rect 44 169 45 170
rect 43 169 44 170
rect 42 169 43 170
rect 41 169 42 170
rect 40 169 41 170
rect 39 169 40 170
rect 38 169 39 170
rect 37 169 38 170
rect 36 169 37 170
rect 35 169 36 170
rect 25 169 26 170
rect 24 169 25 170
rect 23 169 24 170
rect 22 169 23 170
rect 21 169 22 170
rect 20 169 21 170
rect 19 169 20 170
rect 18 169 19 170
rect 17 169 18 170
rect 16 169 17 170
rect 15 169 16 170
rect 14 169 15 170
rect 13 169 14 170
rect 12 169 13 170
rect 11 169 12 170
rect 477 170 478 171
rect 476 170 477 171
rect 475 170 476 171
rect 474 170 475 171
rect 473 170 474 171
rect 472 170 473 171
rect 471 170 472 171
rect 470 170 471 171
rect 469 170 470 171
rect 468 170 469 171
rect 467 170 468 171
rect 466 170 467 171
rect 465 170 466 171
rect 463 170 464 171
rect 462 170 463 171
rect 441 170 442 171
rect 440 170 441 171
rect 439 170 440 171
rect 412 170 413 171
rect 411 170 412 171
rect 410 170 411 171
rect 409 170 410 171
rect 408 170 409 171
rect 407 170 408 171
rect 406 170 407 171
rect 405 170 406 171
rect 404 170 405 171
rect 403 170 404 171
rect 402 170 403 171
rect 401 170 402 171
rect 400 170 401 171
rect 399 170 400 171
rect 398 170 399 171
rect 277 170 278 171
rect 276 170 277 171
rect 275 170 276 171
rect 274 170 275 171
rect 273 170 274 171
rect 272 170 273 171
rect 271 170 272 171
rect 270 170 271 171
rect 269 170 270 171
rect 268 170 269 171
rect 267 170 268 171
rect 266 170 267 171
rect 265 170 266 171
rect 264 170 265 171
rect 263 170 264 171
rect 262 170 263 171
rect 261 170 262 171
rect 260 170 261 171
rect 259 170 260 171
rect 258 170 259 171
rect 257 170 258 171
rect 256 170 257 171
rect 255 170 256 171
rect 254 170 255 171
rect 253 170 254 171
rect 252 170 253 171
rect 251 170 252 171
rect 250 170 251 171
rect 249 170 250 171
rect 248 170 249 171
rect 247 170 248 171
rect 246 170 247 171
rect 245 170 246 171
rect 244 170 245 171
rect 243 170 244 171
rect 242 170 243 171
rect 241 170 242 171
rect 240 170 241 171
rect 239 170 240 171
rect 238 170 239 171
rect 237 170 238 171
rect 236 170 237 171
rect 235 170 236 171
rect 234 170 235 171
rect 233 170 234 171
rect 232 170 233 171
rect 231 170 232 171
rect 212 170 213 171
rect 211 170 212 171
rect 210 170 211 171
rect 209 170 210 171
rect 208 170 209 171
rect 207 170 208 171
rect 206 170 207 171
rect 205 170 206 171
rect 204 170 205 171
rect 203 170 204 171
rect 202 170 203 171
rect 201 170 202 171
rect 200 170 201 171
rect 199 170 200 171
rect 198 170 199 171
rect 197 170 198 171
rect 196 170 197 171
rect 195 170 196 171
rect 194 170 195 171
rect 193 170 194 171
rect 192 170 193 171
rect 191 170 192 171
rect 190 170 191 171
rect 189 170 190 171
rect 188 170 189 171
rect 187 170 188 171
rect 186 170 187 171
rect 185 170 186 171
rect 184 170 185 171
rect 183 170 184 171
rect 182 170 183 171
rect 181 170 182 171
rect 180 170 181 171
rect 179 170 180 171
rect 178 170 179 171
rect 177 170 178 171
rect 176 170 177 171
rect 175 170 176 171
rect 174 170 175 171
rect 173 170 174 171
rect 172 170 173 171
rect 171 170 172 171
rect 170 170 171 171
rect 169 170 170 171
rect 168 170 169 171
rect 167 170 168 171
rect 166 170 167 171
rect 165 170 166 171
rect 164 170 165 171
rect 163 170 164 171
rect 162 170 163 171
rect 161 170 162 171
rect 160 170 161 171
rect 159 170 160 171
rect 158 170 159 171
rect 157 170 158 171
rect 156 170 157 171
rect 155 170 156 171
rect 154 170 155 171
rect 153 170 154 171
rect 152 170 153 171
rect 151 170 152 171
rect 150 170 151 171
rect 149 170 150 171
rect 148 170 149 171
rect 147 170 148 171
rect 146 170 147 171
rect 145 170 146 171
rect 144 170 145 171
rect 143 170 144 171
rect 142 170 143 171
rect 141 170 142 171
rect 140 170 141 171
rect 139 170 140 171
rect 138 170 139 171
rect 64 170 65 171
rect 63 170 64 171
rect 62 170 63 171
rect 61 170 62 171
rect 60 170 61 171
rect 59 170 60 171
rect 58 170 59 171
rect 57 170 58 171
rect 56 170 57 171
rect 55 170 56 171
rect 54 170 55 171
rect 53 170 54 171
rect 52 170 53 171
rect 51 170 52 171
rect 50 170 51 171
rect 49 170 50 171
rect 48 170 49 171
rect 47 170 48 171
rect 46 170 47 171
rect 45 170 46 171
rect 44 170 45 171
rect 43 170 44 171
rect 42 170 43 171
rect 41 170 42 171
rect 40 170 41 171
rect 39 170 40 171
rect 38 170 39 171
rect 37 170 38 171
rect 36 170 37 171
rect 35 170 36 171
rect 25 170 26 171
rect 24 170 25 171
rect 23 170 24 171
rect 22 170 23 171
rect 21 170 22 171
rect 20 170 21 171
rect 19 170 20 171
rect 18 170 19 171
rect 17 170 18 171
rect 16 170 17 171
rect 15 170 16 171
rect 14 170 15 171
rect 13 170 14 171
rect 12 170 13 171
rect 11 170 12 171
rect 480 171 481 172
rect 479 171 480 172
rect 478 171 479 172
rect 477 171 478 172
rect 476 171 477 172
rect 475 171 476 172
rect 474 171 475 172
rect 473 171 474 172
rect 472 171 473 172
rect 471 171 472 172
rect 470 171 471 172
rect 469 171 470 172
rect 468 171 469 172
rect 462 171 463 172
rect 441 171 442 172
rect 440 171 441 172
rect 439 171 440 172
rect 413 171 414 172
rect 412 171 413 172
rect 411 171 412 172
rect 410 171 411 172
rect 409 171 410 172
rect 408 171 409 172
rect 407 171 408 172
rect 406 171 407 172
rect 405 171 406 172
rect 404 171 405 172
rect 403 171 404 172
rect 402 171 403 172
rect 401 171 402 172
rect 400 171 401 172
rect 276 171 277 172
rect 275 171 276 172
rect 274 171 275 172
rect 273 171 274 172
rect 272 171 273 172
rect 271 171 272 172
rect 270 171 271 172
rect 269 171 270 172
rect 268 171 269 172
rect 267 171 268 172
rect 266 171 267 172
rect 265 171 266 172
rect 264 171 265 172
rect 263 171 264 172
rect 262 171 263 172
rect 261 171 262 172
rect 260 171 261 172
rect 259 171 260 172
rect 258 171 259 172
rect 257 171 258 172
rect 256 171 257 172
rect 255 171 256 172
rect 254 171 255 172
rect 253 171 254 172
rect 252 171 253 172
rect 251 171 252 172
rect 250 171 251 172
rect 249 171 250 172
rect 248 171 249 172
rect 247 171 248 172
rect 246 171 247 172
rect 245 171 246 172
rect 244 171 245 172
rect 243 171 244 172
rect 242 171 243 172
rect 241 171 242 172
rect 240 171 241 172
rect 239 171 240 172
rect 238 171 239 172
rect 237 171 238 172
rect 236 171 237 172
rect 235 171 236 172
rect 234 171 235 172
rect 233 171 234 172
rect 232 171 233 172
rect 231 171 232 172
rect 230 171 231 172
rect 211 171 212 172
rect 210 171 211 172
rect 209 171 210 172
rect 208 171 209 172
rect 207 171 208 172
rect 206 171 207 172
rect 205 171 206 172
rect 204 171 205 172
rect 203 171 204 172
rect 202 171 203 172
rect 201 171 202 172
rect 200 171 201 172
rect 199 171 200 172
rect 198 171 199 172
rect 197 171 198 172
rect 196 171 197 172
rect 195 171 196 172
rect 194 171 195 172
rect 193 171 194 172
rect 192 171 193 172
rect 191 171 192 172
rect 190 171 191 172
rect 189 171 190 172
rect 188 171 189 172
rect 187 171 188 172
rect 186 171 187 172
rect 185 171 186 172
rect 184 171 185 172
rect 183 171 184 172
rect 182 171 183 172
rect 181 171 182 172
rect 180 171 181 172
rect 179 171 180 172
rect 178 171 179 172
rect 177 171 178 172
rect 176 171 177 172
rect 175 171 176 172
rect 174 171 175 172
rect 173 171 174 172
rect 172 171 173 172
rect 171 171 172 172
rect 170 171 171 172
rect 169 171 170 172
rect 168 171 169 172
rect 167 171 168 172
rect 166 171 167 172
rect 165 171 166 172
rect 164 171 165 172
rect 163 171 164 172
rect 162 171 163 172
rect 161 171 162 172
rect 160 171 161 172
rect 159 171 160 172
rect 158 171 159 172
rect 157 171 158 172
rect 156 171 157 172
rect 155 171 156 172
rect 154 171 155 172
rect 153 171 154 172
rect 152 171 153 172
rect 151 171 152 172
rect 150 171 151 172
rect 149 171 150 172
rect 148 171 149 172
rect 147 171 148 172
rect 146 171 147 172
rect 145 171 146 172
rect 144 171 145 172
rect 143 171 144 172
rect 142 171 143 172
rect 141 171 142 172
rect 140 171 141 172
rect 139 171 140 172
rect 138 171 139 172
rect 137 171 138 172
rect 63 171 64 172
rect 62 171 63 172
rect 61 171 62 172
rect 60 171 61 172
rect 59 171 60 172
rect 58 171 59 172
rect 57 171 58 172
rect 56 171 57 172
rect 55 171 56 172
rect 54 171 55 172
rect 53 171 54 172
rect 52 171 53 172
rect 51 171 52 172
rect 50 171 51 172
rect 49 171 50 172
rect 48 171 49 172
rect 47 171 48 172
rect 46 171 47 172
rect 45 171 46 172
rect 44 171 45 172
rect 43 171 44 172
rect 42 171 43 172
rect 41 171 42 172
rect 40 171 41 172
rect 39 171 40 172
rect 38 171 39 172
rect 37 171 38 172
rect 36 171 37 172
rect 35 171 36 172
rect 25 171 26 172
rect 24 171 25 172
rect 23 171 24 172
rect 22 171 23 172
rect 21 171 22 172
rect 20 171 21 172
rect 19 171 20 172
rect 18 171 19 172
rect 17 171 18 172
rect 16 171 17 172
rect 15 171 16 172
rect 14 171 15 172
rect 13 171 14 172
rect 12 171 13 172
rect 11 171 12 172
rect 483 172 484 173
rect 482 172 483 173
rect 481 172 482 173
rect 480 172 481 173
rect 479 172 480 173
rect 478 172 479 173
rect 477 172 478 173
rect 476 172 477 173
rect 475 172 476 173
rect 474 172 475 173
rect 473 172 474 173
rect 472 172 473 173
rect 471 172 472 173
rect 441 172 442 173
rect 440 172 441 173
rect 439 172 440 173
rect 414 172 415 173
rect 413 172 414 173
rect 412 172 413 173
rect 411 172 412 173
rect 410 172 411 173
rect 409 172 410 173
rect 408 172 409 173
rect 407 172 408 173
rect 406 172 407 173
rect 405 172 406 173
rect 404 172 405 173
rect 403 172 404 173
rect 402 172 403 173
rect 401 172 402 173
rect 274 172 275 173
rect 273 172 274 173
rect 272 172 273 173
rect 271 172 272 173
rect 270 172 271 173
rect 269 172 270 173
rect 268 172 269 173
rect 267 172 268 173
rect 266 172 267 173
rect 265 172 266 173
rect 264 172 265 173
rect 263 172 264 173
rect 262 172 263 173
rect 261 172 262 173
rect 260 172 261 173
rect 259 172 260 173
rect 258 172 259 173
rect 257 172 258 173
rect 256 172 257 173
rect 255 172 256 173
rect 254 172 255 173
rect 253 172 254 173
rect 252 172 253 173
rect 251 172 252 173
rect 250 172 251 173
rect 249 172 250 173
rect 248 172 249 173
rect 247 172 248 173
rect 246 172 247 173
rect 245 172 246 173
rect 244 172 245 173
rect 243 172 244 173
rect 242 172 243 173
rect 241 172 242 173
rect 240 172 241 173
rect 239 172 240 173
rect 238 172 239 173
rect 237 172 238 173
rect 236 172 237 173
rect 235 172 236 173
rect 234 172 235 173
rect 233 172 234 173
rect 232 172 233 173
rect 231 172 232 173
rect 230 172 231 173
rect 211 172 212 173
rect 210 172 211 173
rect 209 172 210 173
rect 208 172 209 173
rect 207 172 208 173
rect 206 172 207 173
rect 205 172 206 173
rect 204 172 205 173
rect 203 172 204 173
rect 202 172 203 173
rect 201 172 202 173
rect 200 172 201 173
rect 199 172 200 173
rect 198 172 199 173
rect 197 172 198 173
rect 196 172 197 173
rect 195 172 196 173
rect 194 172 195 173
rect 193 172 194 173
rect 192 172 193 173
rect 191 172 192 173
rect 190 172 191 173
rect 189 172 190 173
rect 188 172 189 173
rect 187 172 188 173
rect 186 172 187 173
rect 185 172 186 173
rect 184 172 185 173
rect 183 172 184 173
rect 182 172 183 173
rect 181 172 182 173
rect 180 172 181 173
rect 179 172 180 173
rect 178 172 179 173
rect 177 172 178 173
rect 176 172 177 173
rect 175 172 176 173
rect 174 172 175 173
rect 173 172 174 173
rect 172 172 173 173
rect 171 172 172 173
rect 170 172 171 173
rect 169 172 170 173
rect 168 172 169 173
rect 167 172 168 173
rect 166 172 167 173
rect 165 172 166 173
rect 164 172 165 173
rect 163 172 164 173
rect 162 172 163 173
rect 161 172 162 173
rect 160 172 161 173
rect 159 172 160 173
rect 158 172 159 173
rect 157 172 158 173
rect 156 172 157 173
rect 155 172 156 173
rect 154 172 155 173
rect 153 172 154 173
rect 152 172 153 173
rect 151 172 152 173
rect 150 172 151 173
rect 149 172 150 173
rect 148 172 149 173
rect 147 172 148 173
rect 146 172 147 173
rect 145 172 146 173
rect 144 172 145 173
rect 143 172 144 173
rect 142 172 143 173
rect 141 172 142 173
rect 140 172 141 173
rect 139 172 140 173
rect 138 172 139 173
rect 137 172 138 173
rect 136 172 137 173
rect 135 172 136 173
rect 62 172 63 173
rect 61 172 62 173
rect 60 172 61 173
rect 59 172 60 173
rect 58 172 59 173
rect 57 172 58 173
rect 56 172 57 173
rect 55 172 56 173
rect 54 172 55 173
rect 53 172 54 173
rect 52 172 53 173
rect 51 172 52 173
rect 50 172 51 173
rect 49 172 50 173
rect 48 172 49 173
rect 47 172 48 173
rect 46 172 47 173
rect 45 172 46 173
rect 44 172 45 173
rect 43 172 44 173
rect 42 172 43 173
rect 41 172 42 173
rect 40 172 41 173
rect 39 172 40 173
rect 38 172 39 173
rect 37 172 38 173
rect 36 172 37 173
rect 35 172 36 173
rect 25 172 26 173
rect 24 172 25 173
rect 23 172 24 173
rect 22 172 23 173
rect 21 172 22 173
rect 20 172 21 173
rect 19 172 20 173
rect 18 172 19 173
rect 17 172 18 173
rect 16 172 17 173
rect 15 172 16 173
rect 14 172 15 173
rect 13 172 14 173
rect 12 172 13 173
rect 11 172 12 173
rect 483 173 484 174
rect 482 173 483 174
rect 481 173 482 174
rect 480 173 481 174
rect 479 173 480 174
rect 478 173 479 174
rect 477 173 478 174
rect 476 173 477 174
rect 475 173 476 174
rect 474 173 475 174
rect 473 173 474 174
rect 441 173 442 174
rect 440 173 441 174
rect 415 173 416 174
rect 414 173 415 174
rect 413 173 414 174
rect 412 173 413 174
rect 411 173 412 174
rect 410 173 411 174
rect 409 173 410 174
rect 408 173 409 174
rect 407 173 408 174
rect 406 173 407 174
rect 405 173 406 174
rect 404 173 405 174
rect 403 173 404 174
rect 402 173 403 174
rect 273 173 274 174
rect 272 173 273 174
rect 271 173 272 174
rect 270 173 271 174
rect 269 173 270 174
rect 268 173 269 174
rect 267 173 268 174
rect 266 173 267 174
rect 265 173 266 174
rect 264 173 265 174
rect 263 173 264 174
rect 262 173 263 174
rect 261 173 262 174
rect 260 173 261 174
rect 259 173 260 174
rect 258 173 259 174
rect 257 173 258 174
rect 256 173 257 174
rect 255 173 256 174
rect 254 173 255 174
rect 253 173 254 174
rect 252 173 253 174
rect 251 173 252 174
rect 250 173 251 174
rect 249 173 250 174
rect 248 173 249 174
rect 247 173 248 174
rect 246 173 247 174
rect 245 173 246 174
rect 244 173 245 174
rect 243 173 244 174
rect 242 173 243 174
rect 241 173 242 174
rect 240 173 241 174
rect 239 173 240 174
rect 238 173 239 174
rect 237 173 238 174
rect 236 173 237 174
rect 235 173 236 174
rect 234 173 235 174
rect 233 173 234 174
rect 232 173 233 174
rect 231 173 232 174
rect 230 173 231 174
rect 229 173 230 174
rect 210 173 211 174
rect 209 173 210 174
rect 208 173 209 174
rect 207 173 208 174
rect 206 173 207 174
rect 205 173 206 174
rect 204 173 205 174
rect 203 173 204 174
rect 202 173 203 174
rect 201 173 202 174
rect 200 173 201 174
rect 199 173 200 174
rect 198 173 199 174
rect 197 173 198 174
rect 196 173 197 174
rect 195 173 196 174
rect 194 173 195 174
rect 193 173 194 174
rect 192 173 193 174
rect 191 173 192 174
rect 190 173 191 174
rect 189 173 190 174
rect 188 173 189 174
rect 187 173 188 174
rect 186 173 187 174
rect 185 173 186 174
rect 184 173 185 174
rect 183 173 184 174
rect 182 173 183 174
rect 181 173 182 174
rect 180 173 181 174
rect 179 173 180 174
rect 178 173 179 174
rect 177 173 178 174
rect 176 173 177 174
rect 175 173 176 174
rect 174 173 175 174
rect 173 173 174 174
rect 172 173 173 174
rect 171 173 172 174
rect 170 173 171 174
rect 169 173 170 174
rect 168 173 169 174
rect 167 173 168 174
rect 166 173 167 174
rect 165 173 166 174
rect 164 173 165 174
rect 163 173 164 174
rect 162 173 163 174
rect 161 173 162 174
rect 160 173 161 174
rect 159 173 160 174
rect 158 173 159 174
rect 157 173 158 174
rect 156 173 157 174
rect 155 173 156 174
rect 154 173 155 174
rect 153 173 154 174
rect 152 173 153 174
rect 151 173 152 174
rect 150 173 151 174
rect 149 173 150 174
rect 148 173 149 174
rect 147 173 148 174
rect 146 173 147 174
rect 145 173 146 174
rect 144 173 145 174
rect 143 173 144 174
rect 142 173 143 174
rect 141 173 142 174
rect 140 173 141 174
rect 139 173 140 174
rect 138 173 139 174
rect 137 173 138 174
rect 136 173 137 174
rect 135 173 136 174
rect 134 173 135 174
rect 61 173 62 174
rect 60 173 61 174
rect 59 173 60 174
rect 58 173 59 174
rect 57 173 58 174
rect 56 173 57 174
rect 55 173 56 174
rect 54 173 55 174
rect 53 173 54 174
rect 52 173 53 174
rect 51 173 52 174
rect 50 173 51 174
rect 49 173 50 174
rect 48 173 49 174
rect 47 173 48 174
rect 46 173 47 174
rect 45 173 46 174
rect 44 173 45 174
rect 43 173 44 174
rect 42 173 43 174
rect 41 173 42 174
rect 40 173 41 174
rect 39 173 40 174
rect 38 173 39 174
rect 37 173 38 174
rect 36 173 37 174
rect 24 173 25 174
rect 23 173 24 174
rect 22 173 23 174
rect 21 173 22 174
rect 20 173 21 174
rect 19 173 20 174
rect 18 173 19 174
rect 17 173 18 174
rect 16 173 17 174
rect 15 173 16 174
rect 14 173 15 174
rect 13 173 14 174
rect 12 173 13 174
rect 482 174 483 175
rect 481 174 482 175
rect 480 174 481 175
rect 479 174 480 175
rect 478 174 479 175
rect 477 174 478 175
rect 476 174 477 175
rect 416 174 417 175
rect 415 174 416 175
rect 414 174 415 175
rect 413 174 414 175
rect 412 174 413 175
rect 411 174 412 175
rect 410 174 411 175
rect 409 174 410 175
rect 408 174 409 175
rect 407 174 408 175
rect 406 174 407 175
rect 405 174 406 175
rect 404 174 405 175
rect 403 174 404 175
rect 272 174 273 175
rect 271 174 272 175
rect 270 174 271 175
rect 269 174 270 175
rect 268 174 269 175
rect 267 174 268 175
rect 266 174 267 175
rect 265 174 266 175
rect 264 174 265 175
rect 263 174 264 175
rect 262 174 263 175
rect 261 174 262 175
rect 260 174 261 175
rect 259 174 260 175
rect 258 174 259 175
rect 257 174 258 175
rect 256 174 257 175
rect 255 174 256 175
rect 254 174 255 175
rect 253 174 254 175
rect 252 174 253 175
rect 251 174 252 175
rect 250 174 251 175
rect 249 174 250 175
rect 248 174 249 175
rect 247 174 248 175
rect 246 174 247 175
rect 245 174 246 175
rect 244 174 245 175
rect 243 174 244 175
rect 242 174 243 175
rect 241 174 242 175
rect 240 174 241 175
rect 239 174 240 175
rect 238 174 239 175
rect 237 174 238 175
rect 236 174 237 175
rect 235 174 236 175
rect 234 174 235 175
rect 233 174 234 175
rect 232 174 233 175
rect 231 174 232 175
rect 230 174 231 175
rect 229 174 230 175
rect 228 174 229 175
rect 210 174 211 175
rect 209 174 210 175
rect 208 174 209 175
rect 207 174 208 175
rect 206 174 207 175
rect 205 174 206 175
rect 204 174 205 175
rect 203 174 204 175
rect 202 174 203 175
rect 201 174 202 175
rect 200 174 201 175
rect 199 174 200 175
rect 198 174 199 175
rect 197 174 198 175
rect 196 174 197 175
rect 195 174 196 175
rect 194 174 195 175
rect 193 174 194 175
rect 192 174 193 175
rect 191 174 192 175
rect 190 174 191 175
rect 189 174 190 175
rect 188 174 189 175
rect 187 174 188 175
rect 186 174 187 175
rect 185 174 186 175
rect 184 174 185 175
rect 183 174 184 175
rect 182 174 183 175
rect 181 174 182 175
rect 180 174 181 175
rect 179 174 180 175
rect 178 174 179 175
rect 177 174 178 175
rect 176 174 177 175
rect 175 174 176 175
rect 174 174 175 175
rect 173 174 174 175
rect 172 174 173 175
rect 171 174 172 175
rect 170 174 171 175
rect 169 174 170 175
rect 168 174 169 175
rect 167 174 168 175
rect 166 174 167 175
rect 165 174 166 175
rect 164 174 165 175
rect 163 174 164 175
rect 162 174 163 175
rect 161 174 162 175
rect 160 174 161 175
rect 159 174 160 175
rect 158 174 159 175
rect 157 174 158 175
rect 156 174 157 175
rect 155 174 156 175
rect 154 174 155 175
rect 153 174 154 175
rect 152 174 153 175
rect 151 174 152 175
rect 150 174 151 175
rect 149 174 150 175
rect 148 174 149 175
rect 147 174 148 175
rect 146 174 147 175
rect 145 174 146 175
rect 144 174 145 175
rect 143 174 144 175
rect 142 174 143 175
rect 141 174 142 175
rect 140 174 141 175
rect 139 174 140 175
rect 138 174 139 175
rect 137 174 138 175
rect 136 174 137 175
rect 135 174 136 175
rect 134 174 135 175
rect 133 174 134 175
rect 132 174 133 175
rect 60 174 61 175
rect 59 174 60 175
rect 58 174 59 175
rect 57 174 58 175
rect 56 174 57 175
rect 55 174 56 175
rect 54 174 55 175
rect 53 174 54 175
rect 52 174 53 175
rect 51 174 52 175
rect 50 174 51 175
rect 49 174 50 175
rect 48 174 49 175
rect 47 174 48 175
rect 46 174 47 175
rect 45 174 46 175
rect 44 174 45 175
rect 43 174 44 175
rect 42 174 43 175
rect 41 174 42 175
rect 40 174 41 175
rect 39 174 40 175
rect 38 174 39 175
rect 37 174 38 175
rect 36 174 37 175
rect 24 174 25 175
rect 23 174 24 175
rect 22 174 23 175
rect 21 174 22 175
rect 20 174 21 175
rect 19 174 20 175
rect 18 174 19 175
rect 17 174 18 175
rect 16 174 17 175
rect 15 174 16 175
rect 14 174 15 175
rect 13 174 14 175
rect 12 174 13 175
rect 480 175 481 176
rect 479 175 480 176
rect 478 175 479 176
rect 477 175 478 176
rect 476 175 477 176
rect 418 175 419 176
rect 417 175 418 176
rect 416 175 417 176
rect 415 175 416 176
rect 414 175 415 176
rect 413 175 414 176
rect 412 175 413 176
rect 411 175 412 176
rect 410 175 411 176
rect 409 175 410 176
rect 408 175 409 176
rect 407 175 408 176
rect 406 175 407 176
rect 405 175 406 176
rect 404 175 405 176
rect 271 175 272 176
rect 270 175 271 176
rect 269 175 270 176
rect 268 175 269 176
rect 267 175 268 176
rect 266 175 267 176
rect 265 175 266 176
rect 264 175 265 176
rect 263 175 264 176
rect 262 175 263 176
rect 261 175 262 176
rect 260 175 261 176
rect 259 175 260 176
rect 258 175 259 176
rect 257 175 258 176
rect 256 175 257 176
rect 255 175 256 176
rect 254 175 255 176
rect 253 175 254 176
rect 252 175 253 176
rect 251 175 252 176
rect 250 175 251 176
rect 249 175 250 176
rect 248 175 249 176
rect 247 175 248 176
rect 246 175 247 176
rect 245 175 246 176
rect 244 175 245 176
rect 243 175 244 176
rect 242 175 243 176
rect 241 175 242 176
rect 240 175 241 176
rect 239 175 240 176
rect 238 175 239 176
rect 237 175 238 176
rect 236 175 237 176
rect 235 175 236 176
rect 234 175 235 176
rect 233 175 234 176
rect 232 175 233 176
rect 231 175 232 176
rect 230 175 231 176
rect 229 175 230 176
rect 228 175 229 176
rect 209 175 210 176
rect 208 175 209 176
rect 207 175 208 176
rect 206 175 207 176
rect 205 175 206 176
rect 204 175 205 176
rect 203 175 204 176
rect 202 175 203 176
rect 201 175 202 176
rect 200 175 201 176
rect 199 175 200 176
rect 198 175 199 176
rect 197 175 198 176
rect 196 175 197 176
rect 195 175 196 176
rect 194 175 195 176
rect 193 175 194 176
rect 192 175 193 176
rect 191 175 192 176
rect 190 175 191 176
rect 189 175 190 176
rect 188 175 189 176
rect 187 175 188 176
rect 186 175 187 176
rect 185 175 186 176
rect 184 175 185 176
rect 183 175 184 176
rect 182 175 183 176
rect 181 175 182 176
rect 180 175 181 176
rect 179 175 180 176
rect 178 175 179 176
rect 177 175 178 176
rect 176 175 177 176
rect 175 175 176 176
rect 174 175 175 176
rect 173 175 174 176
rect 172 175 173 176
rect 171 175 172 176
rect 170 175 171 176
rect 169 175 170 176
rect 168 175 169 176
rect 167 175 168 176
rect 166 175 167 176
rect 165 175 166 176
rect 164 175 165 176
rect 163 175 164 176
rect 162 175 163 176
rect 161 175 162 176
rect 160 175 161 176
rect 159 175 160 176
rect 158 175 159 176
rect 157 175 158 176
rect 156 175 157 176
rect 155 175 156 176
rect 154 175 155 176
rect 153 175 154 176
rect 152 175 153 176
rect 151 175 152 176
rect 150 175 151 176
rect 149 175 150 176
rect 148 175 149 176
rect 147 175 148 176
rect 146 175 147 176
rect 145 175 146 176
rect 144 175 145 176
rect 143 175 144 176
rect 142 175 143 176
rect 141 175 142 176
rect 140 175 141 176
rect 139 175 140 176
rect 138 175 139 176
rect 137 175 138 176
rect 136 175 137 176
rect 135 175 136 176
rect 134 175 135 176
rect 133 175 134 176
rect 132 175 133 176
rect 131 175 132 176
rect 130 175 131 176
rect 59 175 60 176
rect 58 175 59 176
rect 57 175 58 176
rect 56 175 57 176
rect 55 175 56 176
rect 54 175 55 176
rect 53 175 54 176
rect 52 175 53 176
rect 51 175 52 176
rect 50 175 51 176
rect 49 175 50 176
rect 48 175 49 176
rect 47 175 48 176
rect 46 175 47 176
rect 45 175 46 176
rect 44 175 45 176
rect 43 175 44 176
rect 42 175 43 176
rect 41 175 42 176
rect 40 175 41 176
rect 39 175 40 176
rect 38 175 39 176
rect 37 175 38 176
rect 36 175 37 176
rect 24 175 25 176
rect 23 175 24 176
rect 22 175 23 176
rect 21 175 22 176
rect 20 175 21 176
rect 19 175 20 176
rect 18 175 19 176
rect 17 175 18 176
rect 16 175 17 176
rect 15 175 16 176
rect 14 175 15 176
rect 13 175 14 176
rect 12 175 13 176
rect 477 176 478 177
rect 476 176 477 177
rect 475 176 476 177
rect 474 176 475 177
rect 473 176 474 177
rect 419 176 420 177
rect 418 176 419 177
rect 417 176 418 177
rect 416 176 417 177
rect 415 176 416 177
rect 414 176 415 177
rect 413 176 414 177
rect 412 176 413 177
rect 411 176 412 177
rect 410 176 411 177
rect 409 176 410 177
rect 408 176 409 177
rect 407 176 408 177
rect 406 176 407 177
rect 405 176 406 177
rect 270 176 271 177
rect 269 176 270 177
rect 268 176 269 177
rect 267 176 268 177
rect 266 176 267 177
rect 265 176 266 177
rect 264 176 265 177
rect 263 176 264 177
rect 262 176 263 177
rect 261 176 262 177
rect 260 176 261 177
rect 259 176 260 177
rect 258 176 259 177
rect 257 176 258 177
rect 256 176 257 177
rect 255 176 256 177
rect 254 176 255 177
rect 253 176 254 177
rect 252 176 253 177
rect 251 176 252 177
rect 250 176 251 177
rect 249 176 250 177
rect 248 176 249 177
rect 247 176 248 177
rect 246 176 247 177
rect 245 176 246 177
rect 244 176 245 177
rect 243 176 244 177
rect 242 176 243 177
rect 241 176 242 177
rect 240 176 241 177
rect 239 176 240 177
rect 238 176 239 177
rect 237 176 238 177
rect 236 176 237 177
rect 235 176 236 177
rect 234 176 235 177
rect 233 176 234 177
rect 232 176 233 177
rect 231 176 232 177
rect 230 176 231 177
rect 229 176 230 177
rect 228 176 229 177
rect 227 176 228 177
rect 208 176 209 177
rect 207 176 208 177
rect 206 176 207 177
rect 205 176 206 177
rect 204 176 205 177
rect 203 176 204 177
rect 202 176 203 177
rect 201 176 202 177
rect 200 176 201 177
rect 199 176 200 177
rect 198 176 199 177
rect 197 176 198 177
rect 196 176 197 177
rect 195 176 196 177
rect 194 176 195 177
rect 193 176 194 177
rect 192 176 193 177
rect 191 176 192 177
rect 190 176 191 177
rect 189 176 190 177
rect 188 176 189 177
rect 187 176 188 177
rect 186 176 187 177
rect 185 176 186 177
rect 184 176 185 177
rect 183 176 184 177
rect 182 176 183 177
rect 181 176 182 177
rect 180 176 181 177
rect 179 176 180 177
rect 178 176 179 177
rect 177 176 178 177
rect 176 176 177 177
rect 175 176 176 177
rect 174 176 175 177
rect 173 176 174 177
rect 172 176 173 177
rect 171 176 172 177
rect 170 176 171 177
rect 169 176 170 177
rect 168 176 169 177
rect 167 176 168 177
rect 166 176 167 177
rect 165 176 166 177
rect 164 176 165 177
rect 163 176 164 177
rect 162 176 163 177
rect 161 176 162 177
rect 160 176 161 177
rect 159 176 160 177
rect 158 176 159 177
rect 157 176 158 177
rect 156 176 157 177
rect 155 176 156 177
rect 154 176 155 177
rect 153 176 154 177
rect 152 176 153 177
rect 151 176 152 177
rect 150 176 151 177
rect 149 176 150 177
rect 148 176 149 177
rect 147 176 148 177
rect 146 176 147 177
rect 145 176 146 177
rect 144 176 145 177
rect 143 176 144 177
rect 142 176 143 177
rect 141 176 142 177
rect 140 176 141 177
rect 139 176 140 177
rect 138 176 139 177
rect 137 176 138 177
rect 136 176 137 177
rect 135 176 136 177
rect 134 176 135 177
rect 133 176 134 177
rect 132 176 133 177
rect 131 176 132 177
rect 130 176 131 177
rect 129 176 130 177
rect 59 176 60 177
rect 58 176 59 177
rect 57 176 58 177
rect 56 176 57 177
rect 55 176 56 177
rect 54 176 55 177
rect 53 176 54 177
rect 52 176 53 177
rect 51 176 52 177
rect 50 176 51 177
rect 49 176 50 177
rect 48 176 49 177
rect 47 176 48 177
rect 46 176 47 177
rect 45 176 46 177
rect 44 176 45 177
rect 43 176 44 177
rect 42 176 43 177
rect 41 176 42 177
rect 40 176 41 177
rect 39 176 40 177
rect 38 176 39 177
rect 37 176 38 177
rect 24 176 25 177
rect 23 176 24 177
rect 22 176 23 177
rect 21 176 22 177
rect 20 176 21 177
rect 19 176 20 177
rect 18 176 19 177
rect 17 176 18 177
rect 16 176 17 177
rect 15 176 16 177
rect 14 176 15 177
rect 13 176 14 177
rect 475 177 476 178
rect 474 177 475 178
rect 473 177 474 178
rect 472 177 473 178
rect 471 177 472 178
rect 462 177 463 178
rect 420 177 421 178
rect 419 177 420 178
rect 418 177 419 178
rect 417 177 418 178
rect 416 177 417 178
rect 415 177 416 178
rect 414 177 415 178
rect 413 177 414 178
rect 412 177 413 178
rect 411 177 412 178
rect 410 177 411 178
rect 409 177 410 178
rect 408 177 409 178
rect 407 177 408 178
rect 269 177 270 178
rect 268 177 269 178
rect 267 177 268 178
rect 266 177 267 178
rect 265 177 266 178
rect 264 177 265 178
rect 263 177 264 178
rect 262 177 263 178
rect 261 177 262 178
rect 260 177 261 178
rect 259 177 260 178
rect 258 177 259 178
rect 257 177 258 178
rect 256 177 257 178
rect 255 177 256 178
rect 254 177 255 178
rect 253 177 254 178
rect 252 177 253 178
rect 251 177 252 178
rect 250 177 251 178
rect 249 177 250 178
rect 248 177 249 178
rect 247 177 248 178
rect 246 177 247 178
rect 245 177 246 178
rect 244 177 245 178
rect 243 177 244 178
rect 242 177 243 178
rect 241 177 242 178
rect 240 177 241 178
rect 239 177 240 178
rect 238 177 239 178
rect 237 177 238 178
rect 236 177 237 178
rect 235 177 236 178
rect 234 177 235 178
rect 233 177 234 178
rect 232 177 233 178
rect 231 177 232 178
rect 230 177 231 178
rect 229 177 230 178
rect 228 177 229 178
rect 227 177 228 178
rect 208 177 209 178
rect 207 177 208 178
rect 206 177 207 178
rect 205 177 206 178
rect 204 177 205 178
rect 203 177 204 178
rect 202 177 203 178
rect 201 177 202 178
rect 200 177 201 178
rect 199 177 200 178
rect 198 177 199 178
rect 197 177 198 178
rect 196 177 197 178
rect 195 177 196 178
rect 194 177 195 178
rect 193 177 194 178
rect 192 177 193 178
rect 191 177 192 178
rect 190 177 191 178
rect 189 177 190 178
rect 188 177 189 178
rect 187 177 188 178
rect 186 177 187 178
rect 185 177 186 178
rect 184 177 185 178
rect 183 177 184 178
rect 182 177 183 178
rect 181 177 182 178
rect 180 177 181 178
rect 179 177 180 178
rect 178 177 179 178
rect 177 177 178 178
rect 176 177 177 178
rect 175 177 176 178
rect 174 177 175 178
rect 173 177 174 178
rect 172 177 173 178
rect 171 177 172 178
rect 170 177 171 178
rect 169 177 170 178
rect 168 177 169 178
rect 167 177 168 178
rect 166 177 167 178
rect 165 177 166 178
rect 164 177 165 178
rect 163 177 164 178
rect 162 177 163 178
rect 161 177 162 178
rect 160 177 161 178
rect 159 177 160 178
rect 158 177 159 178
rect 157 177 158 178
rect 156 177 157 178
rect 155 177 156 178
rect 154 177 155 178
rect 153 177 154 178
rect 152 177 153 178
rect 151 177 152 178
rect 150 177 151 178
rect 149 177 150 178
rect 148 177 149 178
rect 147 177 148 178
rect 146 177 147 178
rect 145 177 146 178
rect 144 177 145 178
rect 143 177 144 178
rect 142 177 143 178
rect 141 177 142 178
rect 140 177 141 178
rect 139 177 140 178
rect 138 177 139 178
rect 137 177 138 178
rect 136 177 137 178
rect 135 177 136 178
rect 134 177 135 178
rect 133 177 134 178
rect 132 177 133 178
rect 131 177 132 178
rect 130 177 131 178
rect 129 177 130 178
rect 128 177 129 178
rect 127 177 128 178
rect 58 177 59 178
rect 57 177 58 178
rect 56 177 57 178
rect 55 177 56 178
rect 54 177 55 178
rect 53 177 54 178
rect 52 177 53 178
rect 51 177 52 178
rect 50 177 51 178
rect 49 177 50 178
rect 48 177 49 178
rect 47 177 48 178
rect 46 177 47 178
rect 45 177 46 178
rect 44 177 45 178
rect 43 177 44 178
rect 42 177 43 178
rect 41 177 42 178
rect 40 177 41 178
rect 39 177 40 178
rect 38 177 39 178
rect 37 177 38 178
rect 25 177 26 178
rect 24 177 25 178
rect 23 177 24 178
rect 22 177 23 178
rect 21 177 22 178
rect 20 177 21 178
rect 19 177 20 178
rect 18 177 19 178
rect 17 177 18 178
rect 16 177 17 178
rect 15 177 16 178
rect 14 177 15 178
rect 13 177 14 178
rect 472 178 473 179
rect 471 178 472 179
rect 470 178 471 179
rect 469 178 470 179
rect 468 178 469 179
rect 462 178 463 179
rect 421 178 422 179
rect 420 178 421 179
rect 419 178 420 179
rect 418 178 419 179
rect 417 178 418 179
rect 416 178 417 179
rect 415 178 416 179
rect 414 178 415 179
rect 413 178 414 179
rect 412 178 413 179
rect 411 178 412 179
rect 410 178 411 179
rect 409 178 410 179
rect 408 178 409 179
rect 268 178 269 179
rect 267 178 268 179
rect 266 178 267 179
rect 265 178 266 179
rect 264 178 265 179
rect 263 178 264 179
rect 262 178 263 179
rect 261 178 262 179
rect 260 178 261 179
rect 259 178 260 179
rect 258 178 259 179
rect 257 178 258 179
rect 256 178 257 179
rect 255 178 256 179
rect 254 178 255 179
rect 253 178 254 179
rect 252 178 253 179
rect 251 178 252 179
rect 250 178 251 179
rect 249 178 250 179
rect 248 178 249 179
rect 247 178 248 179
rect 246 178 247 179
rect 245 178 246 179
rect 244 178 245 179
rect 243 178 244 179
rect 242 178 243 179
rect 241 178 242 179
rect 240 178 241 179
rect 239 178 240 179
rect 238 178 239 179
rect 237 178 238 179
rect 236 178 237 179
rect 235 178 236 179
rect 234 178 235 179
rect 233 178 234 179
rect 232 178 233 179
rect 231 178 232 179
rect 230 178 231 179
rect 229 178 230 179
rect 228 178 229 179
rect 227 178 228 179
rect 226 178 227 179
rect 207 178 208 179
rect 206 178 207 179
rect 205 178 206 179
rect 204 178 205 179
rect 203 178 204 179
rect 202 178 203 179
rect 201 178 202 179
rect 200 178 201 179
rect 199 178 200 179
rect 198 178 199 179
rect 197 178 198 179
rect 196 178 197 179
rect 195 178 196 179
rect 194 178 195 179
rect 193 178 194 179
rect 192 178 193 179
rect 191 178 192 179
rect 190 178 191 179
rect 189 178 190 179
rect 188 178 189 179
rect 187 178 188 179
rect 186 178 187 179
rect 185 178 186 179
rect 184 178 185 179
rect 183 178 184 179
rect 182 178 183 179
rect 181 178 182 179
rect 180 178 181 179
rect 179 178 180 179
rect 178 178 179 179
rect 177 178 178 179
rect 176 178 177 179
rect 175 178 176 179
rect 174 178 175 179
rect 173 178 174 179
rect 172 178 173 179
rect 171 178 172 179
rect 170 178 171 179
rect 169 178 170 179
rect 168 178 169 179
rect 167 178 168 179
rect 166 178 167 179
rect 165 178 166 179
rect 164 178 165 179
rect 163 178 164 179
rect 162 178 163 179
rect 161 178 162 179
rect 160 178 161 179
rect 159 178 160 179
rect 158 178 159 179
rect 157 178 158 179
rect 156 178 157 179
rect 155 178 156 179
rect 154 178 155 179
rect 153 178 154 179
rect 152 178 153 179
rect 151 178 152 179
rect 150 178 151 179
rect 149 178 150 179
rect 148 178 149 179
rect 147 178 148 179
rect 146 178 147 179
rect 145 178 146 179
rect 144 178 145 179
rect 143 178 144 179
rect 142 178 143 179
rect 141 178 142 179
rect 140 178 141 179
rect 139 178 140 179
rect 138 178 139 179
rect 137 178 138 179
rect 136 178 137 179
rect 135 178 136 179
rect 134 178 135 179
rect 133 178 134 179
rect 132 178 133 179
rect 131 178 132 179
rect 130 178 131 179
rect 129 178 130 179
rect 128 178 129 179
rect 127 178 128 179
rect 126 178 127 179
rect 125 178 126 179
rect 57 178 58 179
rect 56 178 57 179
rect 55 178 56 179
rect 54 178 55 179
rect 53 178 54 179
rect 52 178 53 179
rect 51 178 52 179
rect 50 178 51 179
rect 49 178 50 179
rect 48 178 49 179
rect 47 178 48 179
rect 46 178 47 179
rect 45 178 46 179
rect 44 178 45 179
rect 43 178 44 179
rect 42 178 43 179
rect 41 178 42 179
rect 40 178 41 179
rect 39 178 40 179
rect 38 178 39 179
rect 25 178 26 179
rect 24 178 25 179
rect 23 178 24 179
rect 22 178 23 179
rect 21 178 22 179
rect 20 178 21 179
rect 19 178 20 179
rect 18 178 19 179
rect 17 178 18 179
rect 16 178 17 179
rect 15 178 16 179
rect 14 178 15 179
rect 13 178 14 179
rect 469 179 470 180
rect 468 179 469 180
rect 467 179 468 180
rect 466 179 467 180
rect 465 179 466 180
rect 464 179 465 180
rect 463 179 464 180
rect 462 179 463 180
rect 422 179 423 180
rect 421 179 422 180
rect 420 179 421 180
rect 419 179 420 180
rect 418 179 419 180
rect 417 179 418 180
rect 416 179 417 180
rect 415 179 416 180
rect 414 179 415 180
rect 413 179 414 180
rect 412 179 413 180
rect 411 179 412 180
rect 410 179 411 180
rect 409 179 410 180
rect 267 179 268 180
rect 266 179 267 180
rect 265 179 266 180
rect 264 179 265 180
rect 263 179 264 180
rect 262 179 263 180
rect 261 179 262 180
rect 260 179 261 180
rect 259 179 260 180
rect 258 179 259 180
rect 257 179 258 180
rect 256 179 257 180
rect 255 179 256 180
rect 254 179 255 180
rect 253 179 254 180
rect 252 179 253 180
rect 251 179 252 180
rect 250 179 251 180
rect 249 179 250 180
rect 248 179 249 180
rect 247 179 248 180
rect 246 179 247 180
rect 245 179 246 180
rect 244 179 245 180
rect 243 179 244 180
rect 242 179 243 180
rect 241 179 242 180
rect 240 179 241 180
rect 239 179 240 180
rect 238 179 239 180
rect 237 179 238 180
rect 236 179 237 180
rect 235 179 236 180
rect 234 179 235 180
rect 233 179 234 180
rect 232 179 233 180
rect 231 179 232 180
rect 230 179 231 180
rect 229 179 230 180
rect 228 179 229 180
rect 227 179 228 180
rect 226 179 227 180
rect 206 179 207 180
rect 205 179 206 180
rect 204 179 205 180
rect 203 179 204 180
rect 202 179 203 180
rect 201 179 202 180
rect 200 179 201 180
rect 199 179 200 180
rect 198 179 199 180
rect 197 179 198 180
rect 196 179 197 180
rect 195 179 196 180
rect 194 179 195 180
rect 193 179 194 180
rect 192 179 193 180
rect 191 179 192 180
rect 190 179 191 180
rect 189 179 190 180
rect 188 179 189 180
rect 187 179 188 180
rect 186 179 187 180
rect 185 179 186 180
rect 184 179 185 180
rect 183 179 184 180
rect 182 179 183 180
rect 181 179 182 180
rect 180 179 181 180
rect 179 179 180 180
rect 178 179 179 180
rect 177 179 178 180
rect 176 179 177 180
rect 175 179 176 180
rect 174 179 175 180
rect 173 179 174 180
rect 172 179 173 180
rect 171 179 172 180
rect 170 179 171 180
rect 169 179 170 180
rect 168 179 169 180
rect 167 179 168 180
rect 166 179 167 180
rect 165 179 166 180
rect 164 179 165 180
rect 163 179 164 180
rect 162 179 163 180
rect 161 179 162 180
rect 160 179 161 180
rect 159 179 160 180
rect 158 179 159 180
rect 157 179 158 180
rect 156 179 157 180
rect 155 179 156 180
rect 154 179 155 180
rect 153 179 154 180
rect 152 179 153 180
rect 151 179 152 180
rect 150 179 151 180
rect 149 179 150 180
rect 148 179 149 180
rect 147 179 148 180
rect 146 179 147 180
rect 145 179 146 180
rect 144 179 145 180
rect 143 179 144 180
rect 142 179 143 180
rect 141 179 142 180
rect 140 179 141 180
rect 139 179 140 180
rect 138 179 139 180
rect 137 179 138 180
rect 136 179 137 180
rect 135 179 136 180
rect 134 179 135 180
rect 133 179 134 180
rect 132 179 133 180
rect 131 179 132 180
rect 130 179 131 180
rect 129 179 130 180
rect 128 179 129 180
rect 127 179 128 180
rect 126 179 127 180
rect 125 179 126 180
rect 124 179 125 180
rect 123 179 124 180
rect 56 179 57 180
rect 55 179 56 180
rect 54 179 55 180
rect 53 179 54 180
rect 52 179 53 180
rect 51 179 52 180
rect 50 179 51 180
rect 49 179 50 180
rect 48 179 49 180
rect 47 179 48 180
rect 46 179 47 180
rect 45 179 46 180
rect 44 179 45 180
rect 43 179 44 180
rect 42 179 43 180
rect 41 179 42 180
rect 40 179 41 180
rect 39 179 40 180
rect 38 179 39 180
rect 25 179 26 180
rect 24 179 25 180
rect 23 179 24 180
rect 22 179 23 180
rect 21 179 22 180
rect 20 179 21 180
rect 19 179 20 180
rect 18 179 19 180
rect 17 179 18 180
rect 16 179 17 180
rect 15 179 16 180
rect 14 179 15 180
rect 13 179 14 180
rect 467 180 468 181
rect 466 180 467 181
rect 465 180 466 181
rect 464 180 465 181
rect 463 180 464 181
rect 462 180 463 181
rect 424 180 425 181
rect 423 180 424 181
rect 422 180 423 181
rect 421 180 422 181
rect 420 180 421 181
rect 419 180 420 181
rect 418 180 419 181
rect 417 180 418 181
rect 416 180 417 181
rect 415 180 416 181
rect 414 180 415 181
rect 413 180 414 181
rect 412 180 413 181
rect 411 180 412 181
rect 410 180 411 181
rect 267 180 268 181
rect 266 180 267 181
rect 265 180 266 181
rect 264 180 265 181
rect 263 180 264 181
rect 262 180 263 181
rect 261 180 262 181
rect 260 180 261 181
rect 259 180 260 181
rect 258 180 259 181
rect 257 180 258 181
rect 256 180 257 181
rect 255 180 256 181
rect 254 180 255 181
rect 253 180 254 181
rect 252 180 253 181
rect 251 180 252 181
rect 250 180 251 181
rect 249 180 250 181
rect 248 180 249 181
rect 247 180 248 181
rect 246 180 247 181
rect 245 180 246 181
rect 244 180 245 181
rect 243 180 244 181
rect 242 180 243 181
rect 241 180 242 181
rect 240 180 241 181
rect 239 180 240 181
rect 238 180 239 181
rect 237 180 238 181
rect 236 180 237 181
rect 235 180 236 181
rect 234 180 235 181
rect 233 180 234 181
rect 232 180 233 181
rect 231 180 232 181
rect 230 180 231 181
rect 229 180 230 181
rect 228 180 229 181
rect 227 180 228 181
rect 226 180 227 181
rect 225 180 226 181
rect 206 180 207 181
rect 205 180 206 181
rect 204 180 205 181
rect 203 180 204 181
rect 202 180 203 181
rect 201 180 202 181
rect 200 180 201 181
rect 199 180 200 181
rect 198 180 199 181
rect 197 180 198 181
rect 196 180 197 181
rect 195 180 196 181
rect 194 180 195 181
rect 193 180 194 181
rect 192 180 193 181
rect 191 180 192 181
rect 190 180 191 181
rect 189 180 190 181
rect 188 180 189 181
rect 187 180 188 181
rect 186 180 187 181
rect 185 180 186 181
rect 184 180 185 181
rect 183 180 184 181
rect 182 180 183 181
rect 181 180 182 181
rect 180 180 181 181
rect 179 180 180 181
rect 178 180 179 181
rect 177 180 178 181
rect 176 180 177 181
rect 175 180 176 181
rect 174 180 175 181
rect 173 180 174 181
rect 172 180 173 181
rect 171 180 172 181
rect 170 180 171 181
rect 169 180 170 181
rect 168 180 169 181
rect 167 180 168 181
rect 166 180 167 181
rect 165 180 166 181
rect 164 180 165 181
rect 163 180 164 181
rect 162 180 163 181
rect 161 180 162 181
rect 160 180 161 181
rect 159 180 160 181
rect 158 180 159 181
rect 157 180 158 181
rect 156 180 157 181
rect 155 180 156 181
rect 154 180 155 181
rect 153 180 154 181
rect 152 180 153 181
rect 151 180 152 181
rect 150 180 151 181
rect 149 180 150 181
rect 148 180 149 181
rect 147 180 148 181
rect 146 180 147 181
rect 145 180 146 181
rect 144 180 145 181
rect 143 180 144 181
rect 142 180 143 181
rect 141 180 142 181
rect 140 180 141 181
rect 139 180 140 181
rect 138 180 139 181
rect 137 180 138 181
rect 136 180 137 181
rect 135 180 136 181
rect 134 180 135 181
rect 133 180 134 181
rect 132 180 133 181
rect 131 180 132 181
rect 130 180 131 181
rect 129 180 130 181
rect 128 180 129 181
rect 127 180 128 181
rect 126 180 127 181
rect 125 180 126 181
rect 124 180 125 181
rect 123 180 124 181
rect 122 180 123 181
rect 121 180 122 181
rect 120 180 121 181
rect 55 180 56 181
rect 54 180 55 181
rect 53 180 54 181
rect 52 180 53 181
rect 51 180 52 181
rect 50 180 51 181
rect 49 180 50 181
rect 48 180 49 181
rect 47 180 48 181
rect 46 180 47 181
rect 45 180 46 181
rect 44 180 45 181
rect 43 180 44 181
rect 42 180 43 181
rect 41 180 42 181
rect 40 180 41 181
rect 39 180 40 181
rect 25 180 26 181
rect 24 180 25 181
rect 23 180 24 181
rect 22 180 23 181
rect 21 180 22 181
rect 20 180 21 181
rect 19 180 20 181
rect 18 180 19 181
rect 17 180 18 181
rect 16 180 17 181
rect 15 180 16 181
rect 14 180 15 181
rect 13 180 14 181
rect 465 181 466 182
rect 464 181 465 182
rect 463 181 464 182
rect 462 181 463 182
rect 425 181 426 182
rect 424 181 425 182
rect 423 181 424 182
rect 422 181 423 182
rect 421 181 422 182
rect 420 181 421 182
rect 419 181 420 182
rect 418 181 419 182
rect 417 181 418 182
rect 416 181 417 182
rect 415 181 416 182
rect 414 181 415 182
rect 413 181 414 182
rect 412 181 413 182
rect 411 181 412 182
rect 266 181 267 182
rect 265 181 266 182
rect 264 181 265 182
rect 263 181 264 182
rect 262 181 263 182
rect 261 181 262 182
rect 260 181 261 182
rect 259 181 260 182
rect 258 181 259 182
rect 257 181 258 182
rect 256 181 257 182
rect 255 181 256 182
rect 254 181 255 182
rect 253 181 254 182
rect 252 181 253 182
rect 251 181 252 182
rect 250 181 251 182
rect 249 181 250 182
rect 248 181 249 182
rect 247 181 248 182
rect 246 181 247 182
rect 245 181 246 182
rect 244 181 245 182
rect 243 181 244 182
rect 242 181 243 182
rect 241 181 242 182
rect 240 181 241 182
rect 239 181 240 182
rect 238 181 239 182
rect 237 181 238 182
rect 236 181 237 182
rect 235 181 236 182
rect 234 181 235 182
rect 233 181 234 182
rect 232 181 233 182
rect 231 181 232 182
rect 230 181 231 182
rect 229 181 230 182
rect 228 181 229 182
rect 227 181 228 182
rect 226 181 227 182
rect 225 181 226 182
rect 205 181 206 182
rect 204 181 205 182
rect 203 181 204 182
rect 202 181 203 182
rect 201 181 202 182
rect 200 181 201 182
rect 199 181 200 182
rect 198 181 199 182
rect 197 181 198 182
rect 196 181 197 182
rect 195 181 196 182
rect 194 181 195 182
rect 193 181 194 182
rect 192 181 193 182
rect 191 181 192 182
rect 190 181 191 182
rect 189 181 190 182
rect 188 181 189 182
rect 187 181 188 182
rect 186 181 187 182
rect 185 181 186 182
rect 184 181 185 182
rect 183 181 184 182
rect 182 181 183 182
rect 181 181 182 182
rect 180 181 181 182
rect 179 181 180 182
rect 178 181 179 182
rect 177 181 178 182
rect 176 181 177 182
rect 175 181 176 182
rect 174 181 175 182
rect 173 181 174 182
rect 172 181 173 182
rect 171 181 172 182
rect 170 181 171 182
rect 169 181 170 182
rect 168 181 169 182
rect 167 181 168 182
rect 166 181 167 182
rect 165 181 166 182
rect 164 181 165 182
rect 163 181 164 182
rect 162 181 163 182
rect 161 181 162 182
rect 160 181 161 182
rect 159 181 160 182
rect 158 181 159 182
rect 157 181 158 182
rect 156 181 157 182
rect 155 181 156 182
rect 154 181 155 182
rect 153 181 154 182
rect 152 181 153 182
rect 151 181 152 182
rect 150 181 151 182
rect 149 181 150 182
rect 148 181 149 182
rect 147 181 148 182
rect 146 181 147 182
rect 145 181 146 182
rect 144 181 145 182
rect 143 181 144 182
rect 142 181 143 182
rect 141 181 142 182
rect 140 181 141 182
rect 139 181 140 182
rect 138 181 139 182
rect 137 181 138 182
rect 136 181 137 182
rect 135 181 136 182
rect 134 181 135 182
rect 133 181 134 182
rect 132 181 133 182
rect 131 181 132 182
rect 130 181 131 182
rect 129 181 130 182
rect 128 181 129 182
rect 127 181 128 182
rect 126 181 127 182
rect 125 181 126 182
rect 124 181 125 182
rect 123 181 124 182
rect 122 181 123 182
rect 121 181 122 182
rect 120 181 121 182
rect 119 181 120 182
rect 118 181 119 182
rect 54 181 55 182
rect 53 181 54 182
rect 52 181 53 182
rect 51 181 52 182
rect 50 181 51 182
rect 49 181 50 182
rect 48 181 49 182
rect 47 181 48 182
rect 46 181 47 182
rect 45 181 46 182
rect 44 181 45 182
rect 43 181 44 182
rect 42 181 43 182
rect 41 181 42 182
rect 40 181 41 182
rect 25 181 26 182
rect 24 181 25 182
rect 23 181 24 182
rect 22 181 23 182
rect 21 181 22 182
rect 20 181 21 182
rect 19 181 20 182
rect 18 181 19 182
rect 17 181 18 182
rect 16 181 17 182
rect 15 181 16 182
rect 14 181 15 182
rect 463 182 464 183
rect 462 182 463 183
rect 426 182 427 183
rect 425 182 426 183
rect 424 182 425 183
rect 423 182 424 183
rect 422 182 423 183
rect 421 182 422 183
rect 420 182 421 183
rect 419 182 420 183
rect 418 182 419 183
rect 417 182 418 183
rect 416 182 417 183
rect 415 182 416 183
rect 414 182 415 183
rect 413 182 414 183
rect 412 182 413 183
rect 319 182 320 183
rect 318 182 319 183
rect 317 182 318 183
rect 316 182 317 183
rect 315 182 316 183
rect 314 182 315 183
rect 313 182 314 183
rect 312 182 313 183
rect 311 182 312 183
rect 310 182 311 183
rect 309 182 310 183
rect 308 182 309 183
rect 307 182 308 183
rect 306 182 307 183
rect 305 182 306 183
rect 304 182 305 183
rect 303 182 304 183
rect 265 182 266 183
rect 264 182 265 183
rect 263 182 264 183
rect 262 182 263 183
rect 261 182 262 183
rect 260 182 261 183
rect 259 182 260 183
rect 258 182 259 183
rect 257 182 258 183
rect 256 182 257 183
rect 255 182 256 183
rect 254 182 255 183
rect 253 182 254 183
rect 252 182 253 183
rect 251 182 252 183
rect 250 182 251 183
rect 249 182 250 183
rect 248 182 249 183
rect 247 182 248 183
rect 246 182 247 183
rect 245 182 246 183
rect 244 182 245 183
rect 243 182 244 183
rect 242 182 243 183
rect 241 182 242 183
rect 240 182 241 183
rect 239 182 240 183
rect 238 182 239 183
rect 237 182 238 183
rect 236 182 237 183
rect 235 182 236 183
rect 234 182 235 183
rect 233 182 234 183
rect 232 182 233 183
rect 231 182 232 183
rect 230 182 231 183
rect 229 182 230 183
rect 228 182 229 183
rect 227 182 228 183
rect 226 182 227 183
rect 225 182 226 183
rect 224 182 225 183
rect 204 182 205 183
rect 203 182 204 183
rect 202 182 203 183
rect 201 182 202 183
rect 200 182 201 183
rect 199 182 200 183
rect 198 182 199 183
rect 197 182 198 183
rect 196 182 197 183
rect 195 182 196 183
rect 194 182 195 183
rect 193 182 194 183
rect 192 182 193 183
rect 191 182 192 183
rect 190 182 191 183
rect 189 182 190 183
rect 188 182 189 183
rect 187 182 188 183
rect 186 182 187 183
rect 185 182 186 183
rect 184 182 185 183
rect 183 182 184 183
rect 182 182 183 183
rect 181 182 182 183
rect 180 182 181 183
rect 179 182 180 183
rect 178 182 179 183
rect 177 182 178 183
rect 176 182 177 183
rect 175 182 176 183
rect 174 182 175 183
rect 173 182 174 183
rect 172 182 173 183
rect 171 182 172 183
rect 170 182 171 183
rect 169 182 170 183
rect 168 182 169 183
rect 167 182 168 183
rect 166 182 167 183
rect 165 182 166 183
rect 164 182 165 183
rect 163 182 164 183
rect 162 182 163 183
rect 161 182 162 183
rect 160 182 161 183
rect 159 182 160 183
rect 158 182 159 183
rect 157 182 158 183
rect 156 182 157 183
rect 155 182 156 183
rect 154 182 155 183
rect 153 182 154 183
rect 152 182 153 183
rect 151 182 152 183
rect 150 182 151 183
rect 149 182 150 183
rect 148 182 149 183
rect 147 182 148 183
rect 146 182 147 183
rect 145 182 146 183
rect 144 182 145 183
rect 143 182 144 183
rect 142 182 143 183
rect 141 182 142 183
rect 140 182 141 183
rect 139 182 140 183
rect 138 182 139 183
rect 137 182 138 183
rect 136 182 137 183
rect 135 182 136 183
rect 134 182 135 183
rect 133 182 134 183
rect 132 182 133 183
rect 131 182 132 183
rect 130 182 131 183
rect 129 182 130 183
rect 128 182 129 183
rect 127 182 128 183
rect 126 182 127 183
rect 125 182 126 183
rect 124 182 125 183
rect 123 182 124 183
rect 122 182 123 183
rect 121 182 122 183
rect 120 182 121 183
rect 119 182 120 183
rect 118 182 119 183
rect 117 182 118 183
rect 116 182 117 183
rect 115 182 116 183
rect 72 182 73 183
rect 71 182 72 183
rect 52 182 53 183
rect 51 182 52 183
rect 50 182 51 183
rect 49 182 50 183
rect 48 182 49 183
rect 47 182 48 183
rect 46 182 47 183
rect 45 182 46 183
rect 44 182 45 183
rect 43 182 44 183
rect 42 182 43 183
rect 41 182 42 183
rect 25 182 26 183
rect 24 182 25 183
rect 23 182 24 183
rect 22 182 23 183
rect 21 182 22 183
rect 20 182 21 183
rect 19 182 20 183
rect 18 182 19 183
rect 17 182 18 183
rect 16 182 17 183
rect 15 182 16 183
rect 14 182 15 183
rect 462 183 463 184
rect 427 183 428 184
rect 426 183 427 184
rect 425 183 426 184
rect 424 183 425 184
rect 423 183 424 184
rect 422 183 423 184
rect 421 183 422 184
rect 420 183 421 184
rect 419 183 420 184
rect 418 183 419 184
rect 417 183 418 184
rect 416 183 417 184
rect 415 183 416 184
rect 414 183 415 184
rect 413 183 414 184
rect 324 183 325 184
rect 323 183 324 184
rect 322 183 323 184
rect 321 183 322 184
rect 320 183 321 184
rect 319 183 320 184
rect 318 183 319 184
rect 317 183 318 184
rect 316 183 317 184
rect 315 183 316 184
rect 314 183 315 184
rect 313 183 314 184
rect 312 183 313 184
rect 311 183 312 184
rect 310 183 311 184
rect 309 183 310 184
rect 308 183 309 184
rect 307 183 308 184
rect 306 183 307 184
rect 305 183 306 184
rect 304 183 305 184
rect 303 183 304 184
rect 302 183 303 184
rect 301 183 302 184
rect 300 183 301 184
rect 299 183 300 184
rect 298 183 299 184
rect 264 183 265 184
rect 263 183 264 184
rect 262 183 263 184
rect 261 183 262 184
rect 260 183 261 184
rect 259 183 260 184
rect 258 183 259 184
rect 257 183 258 184
rect 256 183 257 184
rect 255 183 256 184
rect 254 183 255 184
rect 253 183 254 184
rect 252 183 253 184
rect 251 183 252 184
rect 250 183 251 184
rect 249 183 250 184
rect 248 183 249 184
rect 247 183 248 184
rect 246 183 247 184
rect 245 183 246 184
rect 244 183 245 184
rect 243 183 244 184
rect 242 183 243 184
rect 241 183 242 184
rect 240 183 241 184
rect 239 183 240 184
rect 238 183 239 184
rect 237 183 238 184
rect 236 183 237 184
rect 235 183 236 184
rect 234 183 235 184
rect 233 183 234 184
rect 232 183 233 184
rect 231 183 232 184
rect 230 183 231 184
rect 229 183 230 184
rect 228 183 229 184
rect 227 183 228 184
rect 226 183 227 184
rect 225 183 226 184
rect 224 183 225 184
rect 203 183 204 184
rect 202 183 203 184
rect 201 183 202 184
rect 200 183 201 184
rect 199 183 200 184
rect 198 183 199 184
rect 197 183 198 184
rect 196 183 197 184
rect 195 183 196 184
rect 194 183 195 184
rect 193 183 194 184
rect 192 183 193 184
rect 191 183 192 184
rect 190 183 191 184
rect 189 183 190 184
rect 188 183 189 184
rect 187 183 188 184
rect 186 183 187 184
rect 185 183 186 184
rect 184 183 185 184
rect 183 183 184 184
rect 182 183 183 184
rect 181 183 182 184
rect 180 183 181 184
rect 179 183 180 184
rect 178 183 179 184
rect 177 183 178 184
rect 176 183 177 184
rect 175 183 176 184
rect 174 183 175 184
rect 173 183 174 184
rect 172 183 173 184
rect 171 183 172 184
rect 170 183 171 184
rect 169 183 170 184
rect 168 183 169 184
rect 167 183 168 184
rect 166 183 167 184
rect 165 183 166 184
rect 164 183 165 184
rect 163 183 164 184
rect 162 183 163 184
rect 161 183 162 184
rect 160 183 161 184
rect 159 183 160 184
rect 158 183 159 184
rect 157 183 158 184
rect 156 183 157 184
rect 155 183 156 184
rect 154 183 155 184
rect 153 183 154 184
rect 152 183 153 184
rect 151 183 152 184
rect 150 183 151 184
rect 149 183 150 184
rect 148 183 149 184
rect 147 183 148 184
rect 146 183 147 184
rect 145 183 146 184
rect 144 183 145 184
rect 143 183 144 184
rect 142 183 143 184
rect 141 183 142 184
rect 140 183 141 184
rect 139 183 140 184
rect 138 183 139 184
rect 137 183 138 184
rect 136 183 137 184
rect 135 183 136 184
rect 134 183 135 184
rect 133 183 134 184
rect 132 183 133 184
rect 131 183 132 184
rect 130 183 131 184
rect 129 183 130 184
rect 128 183 129 184
rect 127 183 128 184
rect 126 183 127 184
rect 125 183 126 184
rect 124 183 125 184
rect 123 183 124 184
rect 122 183 123 184
rect 121 183 122 184
rect 120 183 121 184
rect 119 183 120 184
rect 118 183 119 184
rect 117 183 118 184
rect 116 183 117 184
rect 115 183 116 184
rect 114 183 115 184
rect 113 183 114 184
rect 74 183 75 184
rect 73 183 74 184
rect 72 183 73 184
rect 71 183 72 184
rect 50 183 51 184
rect 49 183 50 184
rect 48 183 49 184
rect 47 183 48 184
rect 46 183 47 184
rect 45 183 46 184
rect 44 183 45 184
rect 43 183 44 184
rect 25 183 26 184
rect 24 183 25 184
rect 23 183 24 184
rect 22 183 23 184
rect 21 183 22 184
rect 20 183 21 184
rect 19 183 20 184
rect 18 183 19 184
rect 17 183 18 184
rect 16 183 17 184
rect 15 183 16 184
rect 14 183 15 184
rect 462 184 463 185
rect 428 184 429 185
rect 427 184 428 185
rect 426 184 427 185
rect 425 184 426 185
rect 424 184 425 185
rect 423 184 424 185
rect 422 184 423 185
rect 421 184 422 185
rect 420 184 421 185
rect 419 184 420 185
rect 418 184 419 185
rect 417 184 418 185
rect 416 184 417 185
rect 415 184 416 185
rect 327 184 328 185
rect 326 184 327 185
rect 325 184 326 185
rect 324 184 325 185
rect 323 184 324 185
rect 322 184 323 185
rect 321 184 322 185
rect 320 184 321 185
rect 319 184 320 185
rect 318 184 319 185
rect 317 184 318 185
rect 316 184 317 185
rect 315 184 316 185
rect 314 184 315 185
rect 313 184 314 185
rect 312 184 313 185
rect 311 184 312 185
rect 310 184 311 185
rect 309 184 310 185
rect 308 184 309 185
rect 307 184 308 185
rect 306 184 307 185
rect 305 184 306 185
rect 304 184 305 185
rect 303 184 304 185
rect 302 184 303 185
rect 301 184 302 185
rect 300 184 301 185
rect 299 184 300 185
rect 298 184 299 185
rect 297 184 298 185
rect 296 184 297 185
rect 295 184 296 185
rect 294 184 295 185
rect 263 184 264 185
rect 262 184 263 185
rect 261 184 262 185
rect 260 184 261 185
rect 259 184 260 185
rect 258 184 259 185
rect 257 184 258 185
rect 256 184 257 185
rect 255 184 256 185
rect 254 184 255 185
rect 253 184 254 185
rect 252 184 253 185
rect 251 184 252 185
rect 250 184 251 185
rect 249 184 250 185
rect 248 184 249 185
rect 247 184 248 185
rect 246 184 247 185
rect 245 184 246 185
rect 244 184 245 185
rect 243 184 244 185
rect 242 184 243 185
rect 241 184 242 185
rect 240 184 241 185
rect 239 184 240 185
rect 238 184 239 185
rect 237 184 238 185
rect 236 184 237 185
rect 235 184 236 185
rect 234 184 235 185
rect 233 184 234 185
rect 232 184 233 185
rect 231 184 232 185
rect 230 184 231 185
rect 229 184 230 185
rect 228 184 229 185
rect 227 184 228 185
rect 226 184 227 185
rect 225 184 226 185
rect 224 184 225 185
rect 223 184 224 185
rect 203 184 204 185
rect 202 184 203 185
rect 201 184 202 185
rect 200 184 201 185
rect 199 184 200 185
rect 198 184 199 185
rect 197 184 198 185
rect 196 184 197 185
rect 195 184 196 185
rect 194 184 195 185
rect 193 184 194 185
rect 192 184 193 185
rect 191 184 192 185
rect 190 184 191 185
rect 189 184 190 185
rect 188 184 189 185
rect 187 184 188 185
rect 186 184 187 185
rect 185 184 186 185
rect 184 184 185 185
rect 183 184 184 185
rect 182 184 183 185
rect 181 184 182 185
rect 180 184 181 185
rect 179 184 180 185
rect 178 184 179 185
rect 177 184 178 185
rect 176 184 177 185
rect 175 184 176 185
rect 174 184 175 185
rect 173 184 174 185
rect 172 184 173 185
rect 171 184 172 185
rect 170 184 171 185
rect 169 184 170 185
rect 168 184 169 185
rect 167 184 168 185
rect 166 184 167 185
rect 165 184 166 185
rect 164 184 165 185
rect 163 184 164 185
rect 162 184 163 185
rect 161 184 162 185
rect 160 184 161 185
rect 159 184 160 185
rect 158 184 159 185
rect 157 184 158 185
rect 156 184 157 185
rect 155 184 156 185
rect 154 184 155 185
rect 153 184 154 185
rect 152 184 153 185
rect 151 184 152 185
rect 150 184 151 185
rect 149 184 150 185
rect 148 184 149 185
rect 147 184 148 185
rect 146 184 147 185
rect 145 184 146 185
rect 144 184 145 185
rect 143 184 144 185
rect 142 184 143 185
rect 141 184 142 185
rect 140 184 141 185
rect 139 184 140 185
rect 138 184 139 185
rect 137 184 138 185
rect 136 184 137 185
rect 135 184 136 185
rect 134 184 135 185
rect 133 184 134 185
rect 132 184 133 185
rect 131 184 132 185
rect 130 184 131 185
rect 129 184 130 185
rect 128 184 129 185
rect 127 184 128 185
rect 126 184 127 185
rect 125 184 126 185
rect 124 184 125 185
rect 123 184 124 185
rect 122 184 123 185
rect 121 184 122 185
rect 120 184 121 185
rect 119 184 120 185
rect 118 184 119 185
rect 117 184 118 185
rect 116 184 117 185
rect 115 184 116 185
rect 114 184 115 185
rect 113 184 114 185
rect 112 184 113 185
rect 111 184 112 185
rect 110 184 111 185
rect 109 184 110 185
rect 77 184 78 185
rect 76 184 77 185
rect 75 184 76 185
rect 74 184 75 185
rect 73 184 74 185
rect 72 184 73 185
rect 71 184 72 185
rect 26 184 27 185
rect 25 184 26 185
rect 24 184 25 185
rect 23 184 24 185
rect 22 184 23 185
rect 21 184 22 185
rect 20 184 21 185
rect 19 184 20 185
rect 18 184 19 185
rect 17 184 18 185
rect 16 184 17 185
rect 15 184 16 185
rect 14 184 15 185
rect 430 185 431 186
rect 429 185 430 186
rect 428 185 429 186
rect 427 185 428 186
rect 426 185 427 186
rect 425 185 426 186
rect 424 185 425 186
rect 423 185 424 186
rect 422 185 423 186
rect 421 185 422 186
rect 420 185 421 186
rect 419 185 420 186
rect 418 185 419 186
rect 417 185 418 186
rect 416 185 417 186
rect 329 185 330 186
rect 328 185 329 186
rect 327 185 328 186
rect 326 185 327 186
rect 325 185 326 186
rect 324 185 325 186
rect 323 185 324 186
rect 322 185 323 186
rect 321 185 322 186
rect 320 185 321 186
rect 319 185 320 186
rect 318 185 319 186
rect 317 185 318 186
rect 316 185 317 186
rect 315 185 316 186
rect 314 185 315 186
rect 313 185 314 186
rect 312 185 313 186
rect 311 185 312 186
rect 310 185 311 186
rect 309 185 310 186
rect 308 185 309 186
rect 307 185 308 186
rect 306 185 307 186
rect 305 185 306 186
rect 304 185 305 186
rect 303 185 304 186
rect 302 185 303 186
rect 301 185 302 186
rect 300 185 301 186
rect 299 185 300 186
rect 298 185 299 186
rect 297 185 298 186
rect 296 185 297 186
rect 295 185 296 186
rect 294 185 295 186
rect 293 185 294 186
rect 292 185 293 186
rect 291 185 292 186
rect 263 185 264 186
rect 262 185 263 186
rect 261 185 262 186
rect 260 185 261 186
rect 259 185 260 186
rect 258 185 259 186
rect 257 185 258 186
rect 256 185 257 186
rect 255 185 256 186
rect 254 185 255 186
rect 253 185 254 186
rect 252 185 253 186
rect 251 185 252 186
rect 250 185 251 186
rect 249 185 250 186
rect 248 185 249 186
rect 247 185 248 186
rect 246 185 247 186
rect 245 185 246 186
rect 244 185 245 186
rect 243 185 244 186
rect 242 185 243 186
rect 241 185 242 186
rect 240 185 241 186
rect 239 185 240 186
rect 238 185 239 186
rect 237 185 238 186
rect 236 185 237 186
rect 235 185 236 186
rect 234 185 235 186
rect 233 185 234 186
rect 232 185 233 186
rect 231 185 232 186
rect 230 185 231 186
rect 229 185 230 186
rect 228 185 229 186
rect 227 185 228 186
rect 226 185 227 186
rect 225 185 226 186
rect 224 185 225 186
rect 223 185 224 186
rect 202 185 203 186
rect 201 185 202 186
rect 200 185 201 186
rect 199 185 200 186
rect 198 185 199 186
rect 197 185 198 186
rect 196 185 197 186
rect 195 185 196 186
rect 194 185 195 186
rect 193 185 194 186
rect 192 185 193 186
rect 191 185 192 186
rect 190 185 191 186
rect 189 185 190 186
rect 188 185 189 186
rect 187 185 188 186
rect 186 185 187 186
rect 185 185 186 186
rect 184 185 185 186
rect 183 185 184 186
rect 182 185 183 186
rect 181 185 182 186
rect 180 185 181 186
rect 179 185 180 186
rect 178 185 179 186
rect 177 185 178 186
rect 176 185 177 186
rect 175 185 176 186
rect 174 185 175 186
rect 173 185 174 186
rect 172 185 173 186
rect 171 185 172 186
rect 170 185 171 186
rect 169 185 170 186
rect 168 185 169 186
rect 167 185 168 186
rect 166 185 167 186
rect 165 185 166 186
rect 164 185 165 186
rect 163 185 164 186
rect 162 185 163 186
rect 161 185 162 186
rect 160 185 161 186
rect 159 185 160 186
rect 158 185 159 186
rect 157 185 158 186
rect 156 185 157 186
rect 155 185 156 186
rect 154 185 155 186
rect 153 185 154 186
rect 152 185 153 186
rect 151 185 152 186
rect 150 185 151 186
rect 149 185 150 186
rect 148 185 149 186
rect 147 185 148 186
rect 146 185 147 186
rect 145 185 146 186
rect 144 185 145 186
rect 143 185 144 186
rect 142 185 143 186
rect 141 185 142 186
rect 140 185 141 186
rect 139 185 140 186
rect 138 185 139 186
rect 137 185 138 186
rect 136 185 137 186
rect 135 185 136 186
rect 134 185 135 186
rect 133 185 134 186
rect 132 185 133 186
rect 131 185 132 186
rect 130 185 131 186
rect 129 185 130 186
rect 128 185 129 186
rect 127 185 128 186
rect 126 185 127 186
rect 125 185 126 186
rect 124 185 125 186
rect 123 185 124 186
rect 122 185 123 186
rect 121 185 122 186
rect 120 185 121 186
rect 119 185 120 186
rect 118 185 119 186
rect 117 185 118 186
rect 116 185 117 186
rect 115 185 116 186
rect 114 185 115 186
rect 113 185 114 186
rect 112 185 113 186
rect 111 185 112 186
rect 110 185 111 186
rect 109 185 110 186
rect 108 185 109 186
rect 107 185 108 186
rect 106 185 107 186
rect 79 185 80 186
rect 78 185 79 186
rect 77 185 78 186
rect 76 185 77 186
rect 75 185 76 186
rect 74 185 75 186
rect 73 185 74 186
rect 72 185 73 186
rect 26 185 27 186
rect 25 185 26 186
rect 24 185 25 186
rect 23 185 24 186
rect 22 185 23 186
rect 21 185 22 186
rect 20 185 21 186
rect 19 185 20 186
rect 18 185 19 186
rect 17 185 18 186
rect 16 185 17 186
rect 15 185 16 186
rect 14 185 15 186
rect 431 186 432 187
rect 430 186 431 187
rect 429 186 430 187
rect 428 186 429 187
rect 427 186 428 187
rect 426 186 427 187
rect 425 186 426 187
rect 424 186 425 187
rect 423 186 424 187
rect 422 186 423 187
rect 421 186 422 187
rect 420 186 421 187
rect 419 186 420 187
rect 418 186 419 187
rect 417 186 418 187
rect 331 186 332 187
rect 330 186 331 187
rect 329 186 330 187
rect 328 186 329 187
rect 327 186 328 187
rect 326 186 327 187
rect 325 186 326 187
rect 324 186 325 187
rect 323 186 324 187
rect 322 186 323 187
rect 321 186 322 187
rect 320 186 321 187
rect 319 186 320 187
rect 318 186 319 187
rect 317 186 318 187
rect 316 186 317 187
rect 315 186 316 187
rect 314 186 315 187
rect 313 186 314 187
rect 312 186 313 187
rect 311 186 312 187
rect 310 186 311 187
rect 309 186 310 187
rect 308 186 309 187
rect 307 186 308 187
rect 306 186 307 187
rect 305 186 306 187
rect 304 186 305 187
rect 303 186 304 187
rect 302 186 303 187
rect 301 186 302 187
rect 300 186 301 187
rect 299 186 300 187
rect 298 186 299 187
rect 297 186 298 187
rect 296 186 297 187
rect 295 186 296 187
rect 294 186 295 187
rect 293 186 294 187
rect 292 186 293 187
rect 291 186 292 187
rect 290 186 291 187
rect 289 186 290 187
rect 262 186 263 187
rect 261 186 262 187
rect 260 186 261 187
rect 259 186 260 187
rect 258 186 259 187
rect 257 186 258 187
rect 256 186 257 187
rect 255 186 256 187
rect 254 186 255 187
rect 253 186 254 187
rect 252 186 253 187
rect 251 186 252 187
rect 250 186 251 187
rect 249 186 250 187
rect 248 186 249 187
rect 247 186 248 187
rect 246 186 247 187
rect 245 186 246 187
rect 244 186 245 187
rect 243 186 244 187
rect 242 186 243 187
rect 241 186 242 187
rect 240 186 241 187
rect 239 186 240 187
rect 238 186 239 187
rect 237 186 238 187
rect 236 186 237 187
rect 235 186 236 187
rect 234 186 235 187
rect 233 186 234 187
rect 232 186 233 187
rect 231 186 232 187
rect 230 186 231 187
rect 229 186 230 187
rect 228 186 229 187
rect 227 186 228 187
rect 226 186 227 187
rect 225 186 226 187
rect 224 186 225 187
rect 223 186 224 187
rect 222 186 223 187
rect 201 186 202 187
rect 200 186 201 187
rect 199 186 200 187
rect 198 186 199 187
rect 197 186 198 187
rect 196 186 197 187
rect 195 186 196 187
rect 194 186 195 187
rect 193 186 194 187
rect 192 186 193 187
rect 191 186 192 187
rect 190 186 191 187
rect 189 186 190 187
rect 188 186 189 187
rect 187 186 188 187
rect 186 186 187 187
rect 185 186 186 187
rect 184 186 185 187
rect 183 186 184 187
rect 182 186 183 187
rect 181 186 182 187
rect 180 186 181 187
rect 179 186 180 187
rect 178 186 179 187
rect 177 186 178 187
rect 176 186 177 187
rect 175 186 176 187
rect 174 186 175 187
rect 173 186 174 187
rect 172 186 173 187
rect 171 186 172 187
rect 170 186 171 187
rect 169 186 170 187
rect 168 186 169 187
rect 167 186 168 187
rect 166 186 167 187
rect 165 186 166 187
rect 164 186 165 187
rect 163 186 164 187
rect 162 186 163 187
rect 161 186 162 187
rect 160 186 161 187
rect 159 186 160 187
rect 158 186 159 187
rect 157 186 158 187
rect 156 186 157 187
rect 155 186 156 187
rect 154 186 155 187
rect 153 186 154 187
rect 152 186 153 187
rect 151 186 152 187
rect 150 186 151 187
rect 149 186 150 187
rect 148 186 149 187
rect 147 186 148 187
rect 146 186 147 187
rect 145 186 146 187
rect 144 186 145 187
rect 143 186 144 187
rect 142 186 143 187
rect 141 186 142 187
rect 140 186 141 187
rect 139 186 140 187
rect 138 186 139 187
rect 137 186 138 187
rect 136 186 137 187
rect 135 186 136 187
rect 134 186 135 187
rect 133 186 134 187
rect 132 186 133 187
rect 131 186 132 187
rect 130 186 131 187
rect 129 186 130 187
rect 128 186 129 187
rect 127 186 128 187
rect 126 186 127 187
rect 125 186 126 187
rect 124 186 125 187
rect 123 186 124 187
rect 122 186 123 187
rect 121 186 122 187
rect 120 186 121 187
rect 119 186 120 187
rect 118 186 119 187
rect 117 186 118 187
rect 116 186 117 187
rect 115 186 116 187
rect 114 186 115 187
rect 113 186 114 187
rect 112 186 113 187
rect 111 186 112 187
rect 110 186 111 187
rect 109 186 110 187
rect 108 186 109 187
rect 107 186 108 187
rect 106 186 107 187
rect 105 186 106 187
rect 104 186 105 187
rect 103 186 104 187
rect 102 186 103 187
rect 101 186 102 187
rect 83 186 84 187
rect 82 186 83 187
rect 81 186 82 187
rect 80 186 81 187
rect 79 186 80 187
rect 78 186 79 187
rect 77 186 78 187
rect 76 186 77 187
rect 75 186 76 187
rect 74 186 75 187
rect 73 186 74 187
rect 72 186 73 187
rect 26 186 27 187
rect 25 186 26 187
rect 24 186 25 187
rect 23 186 24 187
rect 22 186 23 187
rect 21 186 22 187
rect 20 186 21 187
rect 19 186 20 187
rect 18 186 19 187
rect 17 186 18 187
rect 16 186 17 187
rect 15 186 16 187
rect 14 186 15 187
rect 432 187 433 188
rect 431 187 432 188
rect 430 187 431 188
rect 429 187 430 188
rect 428 187 429 188
rect 427 187 428 188
rect 426 187 427 188
rect 425 187 426 188
rect 424 187 425 188
rect 423 187 424 188
rect 422 187 423 188
rect 421 187 422 188
rect 420 187 421 188
rect 419 187 420 188
rect 418 187 419 188
rect 333 187 334 188
rect 332 187 333 188
rect 331 187 332 188
rect 330 187 331 188
rect 329 187 330 188
rect 328 187 329 188
rect 327 187 328 188
rect 326 187 327 188
rect 325 187 326 188
rect 324 187 325 188
rect 323 187 324 188
rect 322 187 323 188
rect 321 187 322 188
rect 320 187 321 188
rect 319 187 320 188
rect 318 187 319 188
rect 317 187 318 188
rect 316 187 317 188
rect 315 187 316 188
rect 314 187 315 188
rect 313 187 314 188
rect 312 187 313 188
rect 311 187 312 188
rect 310 187 311 188
rect 309 187 310 188
rect 308 187 309 188
rect 307 187 308 188
rect 306 187 307 188
rect 305 187 306 188
rect 304 187 305 188
rect 303 187 304 188
rect 302 187 303 188
rect 301 187 302 188
rect 300 187 301 188
rect 299 187 300 188
rect 298 187 299 188
rect 297 187 298 188
rect 296 187 297 188
rect 295 187 296 188
rect 294 187 295 188
rect 293 187 294 188
rect 292 187 293 188
rect 291 187 292 188
rect 290 187 291 188
rect 289 187 290 188
rect 288 187 289 188
rect 287 187 288 188
rect 286 187 287 188
rect 261 187 262 188
rect 260 187 261 188
rect 259 187 260 188
rect 258 187 259 188
rect 257 187 258 188
rect 256 187 257 188
rect 255 187 256 188
rect 254 187 255 188
rect 253 187 254 188
rect 252 187 253 188
rect 251 187 252 188
rect 250 187 251 188
rect 249 187 250 188
rect 248 187 249 188
rect 247 187 248 188
rect 246 187 247 188
rect 245 187 246 188
rect 244 187 245 188
rect 243 187 244 188
rect 242 187 243 188
rect 241 187 242 188
rect 240 187 241 188
rect 239 187 240 188
rect 238 187 239 188
rect 237 187 238 188
rect 236 187 237 188
rect 235 187 236 188
rect 234 187 235 188
rect 233 187 234 188
rect 232 187 233 188
rect 231 187 232 188
rect 230 187 231 188
rect 229 187 230 188
rect 228 187 229 188
rect 227 187 228 188
rect 226 187 227 188
rect 225 187 226 188
rect 224 187 225 188
rect 223 187 224 188
rect 222 187 223 188
rect 221 187 222 188
rect 200 187 201 188
rect 199 187 200 188
rect 198 187 199 188
rect 197 187 198 188
rect 196 187 197 188
rect 195 187 196 188
rect 194 187 195 188
rect 193 187 194 188
rect 192 187 193 188
rect 191 187 192 188
rect 190 187 191 188
rect 189 187 190 188
rect 188 187 189 188
rect 187 187 188 188
rect 186 187 187 188
rect 185 187 186 188
rect 184 187 185 188
rect 183 187 184 188
rect 182 187 183 188
rect 181 187 182 188
rect 180 187 181 188
rect 179 187 180 188
rect 178 187 179 188
rect 177 187 178 188
rect 176 187 177 188
rect 175 187 176 188
rect 174 187 175 188
rect 173 187 174 188
rect 172 187 173 188
rect 171 187 172 188
rect 170 187 171 188
rect 169 187 170 188
rect 168 187 169 188
rect 167 187 168 188
rect 166 187 167 188
rect 165 187 166 188
rect 164 187 165 188
rect 163 187 164 188
rect 162 187 163 188
rect 161 187 162 188
rect 160 187 161 188
rect 159 187 160 188
rect 158 187 159 188
rect 157 187 158 188
rect 156 187 157 188
rect 155 187 156 188
rect 154 187 155 188
rect 153 187 154 188
rect 152 187 153 188
rect 151 187 152 188
rect 150 187 151 188
rect 149 187 150 188
rect 148 187 149 188
rect 147 187 148 188
rect 146 187 147 188
rect 145 187 146 188
rect 144 187 145 188
rect 143 187 144 188
rect 142 187 143 188
rect 141 187 142 188
rect 140 187 141 188
rect 139 187 140 188
rect 138 187 139 188
rect 137 187 138 188
rect 136 187 137 188
rect 135 187 136 188
rect 134 187 135 188
rect 133 187 134 188
rect 132 187 133 188
rect 131 187 132 188
rect 130 187 131 188
rect 129 187 130 188
rect 128 187 129 188
rect 127 187 128 188
rect 126 187 127 188
rect 125 187 126 188
rect 124 187 125 188
rect 123 187 124 188
rect 122 187 123 188
rect 121 187 122 188
rect 120 187 121 188
rect 119 187 120 188
rect 118 187 119 188
rect 117 187 118 188
rect 116 187 117 188
rect 115 187 116 188
rect 114 187 115 188
rect 113 187 114 188
rect 112 187 113 188
rect 111 187 112 188
rect 110 187 111 188
rect 109 187 110 188
rect 108 187 109 188
rect 107 187 108 188
rect 106 187 107 188
rect 105 187 106 188
rect 104 187 105 188
rect 103 187 104 188
rect 102 187 103 188
rect 101 187 102 188
rect 100 187 101 188
rect 99 187 100 188
rect 98 187 99 188
rect 97 187 98 188
rect 96 187 97 188
rect 95 187 96 188
rect 94 187 95 188
rect 93 187 94 188
rect 92 187 93 188
rect 91 187 92 188
rect 90 187 91 188
rect 89 187 90 188
rect 88 187 89 188
rect 87 187 88 188
rect 86 187 87 188
rect 85 187 86 188
rect 84 187 85 188
rect 83 187 84 188
rect 82 187 83 188
rect 81 187 82 188
rect 80 187 81 188
rect 79 187 80 188
rect 78 187 79 188
rect 77 187 78 188
rect 76 187 77 188
rect 75 187 76 188
rect 74 187 75 188
rect 73 187 74 188
rect 72 187 73 188
rect 26 187 27 188
rect 25 187 26 188
rect 24 187 25 188
rect 23 187 24 188
rect 22 187 23 188
rect 21 187 22 188
rect 20 187 21 188
rect 19 187 20 188
rect 18 187 19 188
rect 17 187 18 188
rect 16 187 17 188
rect 15 187 16 188
rect 14 187 15 188
rect 433 188 434 189
rect 432 188 433 189
rect 431 188 432 189
rect 430 188 431 189
rect 429 188 430 189
rect 428 188 429 189
rect 427 188 428 189
rect 426 188 427 189
rect 425 188 426 189
rect 424 188 425 189
rect 423 188 424 189
rect 422 188 423 189
rect 421 188 422 189
rect 420 188 421 189
rect 419 188 420 189
rect 398 188 399 189
rect 397 188 398 189
rect 335 188 336 189
rect 334 188 335 189
rect 333 188 334 189
rect 332 188 333 189
rect 331 188 332 189
rect 330 188 331 189
rect 329 188 330 189
rect 328 188 329 189
rect 327 188 328 189
rect 326 188 327 189
rect 325 188 326 189
rect 324 188 325 189
rect 323 188 324 189
rect 322 188 323 189
rect 321 188 322 189
rect 320 188 321 189
rect 319 188 320 189
rect 318 188 319 189
rect 317 188 318 189
rect 316 188 317 189
rect 315 188 316 189
rect 314 188 315 189
rect 313 188 314 189
rect 312 188 313 189
rect 311 188 312 189
rect 310 188 311 189
rect 309 188 310 189
rect 308 188 309 189
rect 307 188 308 189
rect 306 188 307 189
rect 305 188 306 189
rect 304 188 305 189
rect 303 188 304 189
rect 302 188 303 189
rect 301 188 302 189
rect 300 188 301 189
rect 299 188 300 189
rect 298 188 299 189
rect 297 188 298 189
rect 296 188 297 189
rect 295 188 296 189
rect 294 188 295 189
rect 293 188 294 189
rect 292 188 293 189
rect 291 188 292 189
rect 290 188 291 189
rect 289 188 290 189
rect 288 188 289 189
rect 287 188 288 189
rect 286 188 287 189
rect 285 188 286 189
rect 284 188 285 189
rect 261 188 262 189
rect 260 188 261 189
rect 259 188 260 189
rect 258 188 259 189
rect 257 188 258 189
rect 256 188 257 189
rect 255 188 256 189
rect 254 188 255 189
rect 253 188 254 189
rect 252 188 253 189
rect 251 188 252 189
rect 250 188 251 189
rect 249 188 250 189
rect 248 188 249 189
rect 247 188 248 189
rect 246 188 247 189
rect 245 188 246 189
rect 244 188 245 189
rect 243 188 244 189
rect 242 188 243 189
rect 241 188 242 189
rect 240 188 241 189
rect 239 188 240 189
rect 238 188 239 189
rect 237 188 238 189
rect 236 188 237 189
rect 235 188 236 189
rect 234 188 235 189
rect 233 188 234 189
rect 232 188 233 189
rect 231 188 232 189
rect 230 188 231 189
rect 229 188 230 189
rect 228 188 229 189
rect 227 188 228 189
rect 226 188 227 189
rect 225 188 226 189
rect 224 188 225 189
rect 223 188 224 189
rect 222 188 223 189
rect 221 188 222 189
rect 199 188 200 189
rect 198 188 199 189
rect 197 188 198 189
rect 196 188 197 189
rect 195 188 196 189
rect 194 188 195 189
rect 193 188 194 189
rect 192 188 193 189
rect 191 188 192 189
rect 190 188 191 189
rect 189 188 190 189
rect 188 188 189 189
rect 187 188 188 189
rect 186 188 187 189
rect 185 188 186 189
rect 184 188 185 189
rect 183 188 184 189
rect 182 188 183 189
rect 181 188 182 189
rect 180 188 181 189
rect 179 188 180 189
rect 178 188 179 189
rect 177 188 178 189
rect 176 188 177 189
rect 175 188 176 189
rect 174 188 175 189
rect 173 188 174 189
rect 172 188 173 189
rect 171 188 172 189
rect 170 188 171 189
rect 169 188 170 189
rect 168 188 169 189
rect 167 188 168 189
rect 166 188 167 189
rect 165 188 166 189
rect 164 188 165 189
rect 163 188 164 189
rect 162 188 163 189
rect 161 188 162 189
rect 160 188 161 189
rect 159 188 160 189
rect 158 188 159 189
rect 157 188 158 189
rect 156 188 157 189
rect 155 188 156 189
rect 154 188 155 189
rect 153 188 154 189
rect 152 188 153 189
rect 151 188 152 189
rect 150 188 151 189
rect 149 188 150 189
rect 148 188 149 189
rect 147 188 148 189
rect 146 188 147 189
rect 145 188 146 189
rect 144 188 145 189
rect 143 188 144 189
rect 142 188 143 189
rect 141 188 142 189
rect 140 188 141 189
rect 139 188 140 189
rect 138 188 139 189
rect 137 188 138 189
rect 136 188 137 189
rect 135 188 136 189
rect 134 188 135 189
rect 133 188 134 189
rect 132 188 133 189
rect 131 188 132 189
rect 130 188 131 189
rect 129 188 130 189
rect 128 188 129 189
rect 127 188 128 189
rect 126 188 127 189
rect 125 188 126 189
rect 124 188 125 189
rect 123 188 124 189
rect 122 188 123 189
rect 121 188 122 189
rect 120 188 121 189
rect 119 188 120 189
rect 118 188 119 189
rect 117 188 118 189
rect 116 188 117 189
rect 115 188 116 189
rect 114 188 115 189
rect 113 188 114 189
rect 112 188 113 189
rect 111 188 112 189
rect 110 188 111 189
rect 109 188 110 189
rect 108 188 109 189
rect 107 188 108 189
rect 106 188 107 189
rect 105 188 106 189
rect 104 188 105 189
rect 103 188 104 189
rect 102 188 103 189
rect 101 188 102 189
rect 100 188 101 189
rect 99 188 100 189
rect 98 188 99 189
rect 97 188 98 189
rect 96 188 97 189
rect 95 188 96 189
rect 94 188 95 189
rect 93 188 94 189
rect 92 188 93 189
rect 91 188 92 189
rect 90 188 91 189
rect 89 188 90 189
rect 88 188 89 189
rect 87 188 88 189
rect 86 188 87 189
rect 85 188 86 189
rect 84 188 85 189
rect 83 188 84 189
rect 82 188 83 189
rect 81 188 82 189
rect 80 188 81 189
rect 79 188 80 189
rect 78 188 79 189
rect 77 188 78 189
rect 76 188 77 189
rect 75 188 76 189
rect 74 188 75 189
rect 73 188 74 189
rect 72 188 73 189
rect 27 188 28 189
rect 26 188 27 189
rect 25 188 26 189
rect 24 188 25 189
rect 23 188 24 189
rect 22 188 23 189
rect 21 188 22 189
rect 20 188 21 189
rect 19 188 20 189
rect 18 188 19 189
rect 17 188 18 189
rect 16 188 17 189
rect 15 188 16 189
rect 14 188 15 189
rect 434 189 435 190
rect 433 189 434 190
rect 432 189 433 190
rect 431 189 432 190
rect 430 189 431 190
rect 429 189 430 190
rect 428 189 429 190
rect 427 189 428 190
rect 426 189 427 190
rect 425 189 426 190
rect 424 189 425 190
rect 423 189 424 190
rect 422 189 423 190
rect 421 189 422 190
rect 420 189 421 190
rect 399 189 400 190
rect 398 189 399 190
rect 397 189 398 190
rect 337 189 338 190
rect 336 189 337 190
rect 335 189 336 190
rect 334 189 335 190
rect 333 189 334 190
rect 332 189 333 190
rect 331 189 332 190
rect 330 189 331 190
rect 329 189 330 190
rect 328 189 329 190
rect 327 189 328 190
rect 326 189 327 190
rect 325 189 326 190
rect 324 189 325 190
rect 323 189 324 190
rect 322 189 323 190
rect 321 189 322 190
rect 320 189 321 190
rect 319 189 320 190
rect 318 189 319 190
rect 317 189 318 190
rect 316 189 317 190
rect 315 189 316 190
rect 314 189 315 190
rect 313 189 314 190
rect 312 189 313 190
rect 311 189 312 190
rect 310 189 311 190
rect 309 189 310 190
rect 308 189 309 190
rect 307 189 308 190
rect 306 189 307 190
rect 305 189 306 190
rect 304 189 305 190
rect 303 189 304 190
rect 302 189 303 190
rect 301 189 302 190
rect 300 189 301 190
rect 299 189 300 190
rect 298 189 299 190
rect 297 189 298 190
rect 296 189 297 190
rect 295 189 296 190
rect 294 189 295 190
rect 293 189 294 190
rect 292 189 293 190
rect 291 189 292 190
rect 290 189 291 190
rect 289 189 290 190
rect 288 189 289 190
rect 287 189 288 190
rect 286 189 287 190
rect 285 189 286 190
rect 284 189 285 190
rect 283 189 284 190
rect 282 189 283 190
rect 260 189 261 190
rect 259 189 260 190
rect 258 189 259 190
rect 257 189 258 190
rect 256 189 257 190
rect 255 189 256 190
rect 254 189 255 190
rect 253 189 254 190
rect 252 189 253 190
rect 251 189 252 190
rect 250 189 251 190
rect 249 189 250 190
rect 248 189 249 190
rect 247 189 248 190
rect 246 189 247 190
rect 245 189 246 190
rect 244 189 245 190
rect 243 189 244 190
rect 242 189 243 190
rect 241 189 242 190
rect 240 189 241 190
rect 239 189 240 190
rect 238 189 239 190
rect 237 189 238 190
rect 236 189 237 190
rect 235 189 236 190
rect 234 189 235 190
rect 233 189 234 190
rect 232 189 233 190
rect 231 189 232 190
rect 230 189 231 190
rect 229 189 230 190
rect 228 189 229 190
rect 227 189 228 190
rect 226 189 227 190
rect 225 189 226 190
rect 224 189 225 190
rect 223 189 224 190
rect 222 189 223 190
rect 221 189 222 190
rect 220 189 221 190
rect 198 189 199 190
rect 197 189 198 190
rect 196 189 197 190
rect 195 189 196 190
rect 194 189 195 190
rect 193 189 194 190
rect 192 189 193 190
rect 191 189 192 190
rect 190 189 191 190
rect 189 189 190 190
rect 188 189 189 190
rect 187 189 188 190
rect 186 189 187 190
rect 185 189 186 190
rect 184 189 185 190
rect 183 189 184 190
rect 182 189 183 190
rect 181 189 182 190
rect 180 189 181 190
rect 179 189 180 190
rect 178 189 179 190
rect 177 189 178 190
rect 176 189 177 190
rect 175 189 176 190
rect 174 189 175 190
rect 173 189 174 190
rect 172 189 173 190
rect 171 189 172 190
rect 170 189 171 190
rect 169 189 170 190
rect 168 189 169 190
rect 167 189 168 190
rect 166 189 167 190
rect 165 189 166 190
rect 164 189 165 190
rect 163 189 164 190
rect 162 189 163 190
rect 161 189 162 190
rect 160 189 161 190
rect 159 189 160 190
rect 158 189 159 190
rect 157 189 158 190
rect 156 189 157 190
rect 155 189 156 190
rect 154 189 155 190
rect 153 189 154 190
rect 152 189 153 190
rect 151 189 152 190
rect 150 189 151 190
rect 149 189 150 190
rect 148 189 149 190
rect 147 189 148 190
rect 146 189 147 190
rect 145 189 146 190
rect 144 189 145 190
rect 143 189 144 190
rect 142 189 143 190
rect 141 189 142 190
rect 140 189 141 190
rect 139 189 140 190
rect 138 189 139 190
rect 137 189 138 190
rect 136 189 137 190
rect 135 189 136 190
rect 134 189 135 190
rect 133 189 134 190
rect 132 189 133 190
rect 131 189 132 190
rect 130 189 131 190
rect 129 189 130 190
rect 128 189 129 190
rect 127 189 128 190
rect 126 189 127 190
rect 125 189 126 190
rect 124 189 125 190
rect 123 189 124 190
rect 122 189 123 190
rect 121 189 122 190
rect 120 189 121 190
rect 119 189 120 190
rect 118 189 119 190
rect 117 189 118 190
rect 116 189 117 190
rect 115 189 116 190
rect 114 189 115 190
rect 113 189 114 190
rect 112 189 113 190
rect 111 189 112 190
rect 110 189 111 190
rect 109 189 110 190
rect 108 189 109 190
rect 107 189 108 190
rect 106 189 107 190
rect 105 189 106 190
rect 104 189 105 190
rect 103 189 104 190
rect 102 189 103 190
rect 101 189 102 190
rect 100 189 101 190
rect 99 189 100 190
rect 98 189 99 190
rect 97 189 98 190
rect 96 189 97 190
rect 95 189 96 190
rect 94 189 95 190
rect 93 189 94 190
rect 92 189 93 190
rect 91 189 92 190
rect 90 189 91 190
rect 89 189 90 190
rect 88 189 89 190
rect 87 189 88 190
rect 86 189 87 190
rect 85 189 86 190
rect 84 189 85 190
rect 83 189 84 190
rect 82 189 83 190
rect 81 189 82 190
rect 80 189 81 190
rect 79 189 80 190
rect 78 189 79 190
rect 77 189 78 190
rect 76 189 77 190
rect 75 189 76 190
rect 74 189 75 190
rect 73 189 74 190
rect 72 189 73 190
rect 27 189 28 190
rect 26 189 27 190
rect 25 189 26 190
rect 24 189 25 190
rect 23 189 24 190
rect 22 189 23 190
rect 21 189 22 190
rect 20 189 21 190
rect 19 189 20 190
rect 18 189 19 190
rect 17 189 18 190
rect 16 189 17 190
rect 15 189 16 190
rect 14 189 15 190
rect 436 190 437 191
rect 435 190 436 191
rect 434 190 435 191
rect 433 190 434 191
rect 432 190 433 191
rect 431 190 432 191
rect 430 190 431 191
rect 429 190 430 191
rect 428 190 429 191
rect 427 190 428 191
rect 426 190 427 191
rect 425 190 426 191
rect 424 190 425 191
rect 423 190 424 191
rect 422 190 423 191
rect 421 190 422 191
rect 399 190 400 191
rect 398 190 399 191
rect 397 190 398 191
rect 338 190 339 191
rect 337 190 338 191
rect 336 190 337 191
rect 335 190 336 191
rect 334 190 335 191
rect 333 190 334 191
rect 332 190 333 191
rect 331 190 332 191
rect 330 190 331 191
rect 329 190 330 191
rect 328 190 329 191
rect 327 190 328 191
rect 326 190 327 191
rect 325 190 326 191
rect 324 190 325 191
rect 323 190 324 191
rect 322 190 323 191
rect 321 190 322 191
rect 320 190 321 191
rect 319 190 320 191
rect 318 190 319 191
rect 317 190 318 191
rect 316 190 317 191
rect 315 190 316 191
rect 314 190 315 191
rect 313 190 314 191
rect 312 190 313 191
rect 311 190 312 191
rect 310 190 311 191
rect 309 190 310 191
rect 308 190 309 191
rect 307 190 308 191
rect 306 190 307 191
rect 305 190 306 191
rect 304 190 305 191
rect 303 190 304 191
rect 302 190 303 191
rect 301 190 302 191
rect 300 190 301 191
rect 299 190 300 191
rect 298 190 299 191
rect 297 190 298 191
rect 296 190 297 191
rect 295 190 296 191
rect 294 190 295 191
rect 293 190 294 191
rect 292 190 293 191
rect 291 190 292 191
rect 290 190 291 191
rect 289 190 290 191
rect 288 190 289 191
rect 287 190 288 191
rect 286 190 287 191
rect 285 190 286 191
rect 284 190 285 191
rect 283 190 284 191
rect 282 190 283 191
rect 281 190 282 191
rect 280 190 281 191
rect 259 190 260 191
rect 258 190 259 191
rect 257 190 258 191
rect 256 190 257 191
rect 255 190 256 191
rect 254 190 255 191
rect 253 190 254 191
rect 252 190 253 191
rect 251 190 252 191
rect 250 190 251 191
rect 249 190 250 191
rect 248 190 249 191
rect 247 190 248 191
rect 246 190 247 191
rect 245 190 246 191
rect 244 190 245 191
rect 243 190 244 191
rect 242 190 243 191
rect 241 190 242 191
rect 240 190 241 191
rect 239 190 240 191
rect 238 190 239 191
rect 237 190 238 191
rect 236 190 237 191
rect 235 190 236 191
rect 234 190 235 191
rect 233 190 234 191
rect 232 190 233 191
rect 231 190 232 191
rect 230 190 231 191
rect 229 190 230 191
rect 228 190 229 191
rect 227 190 228 191
rect 226 190 227 191
rect 225 190 226 191
rect 224 190 225 191
rect 223 190 224 191
rect 222 190 223 191
rect 221 190 222 191
rect 220 190 221 191
rect 197 190 198 191
rect 196 190 197 191
rect 195 190 196 191
rect 194 190 195 191
rect 193 190 194 191
rect 192 190 193 191
rect 191 190 192 191
rect 190 190 191 191
rect 189 190 190 191
rect 188 190 189 191
rect 187 190 188 191
rect 186 190 187 191
rect 185 190 186 191
rect 184 190 185 191
rect 183 190 184 191
rect 182 190 183 191
rect 181 190 182 191
rect 180 190 181 191
rect 179 190 180 191
rect 178 190 179 191
rect 177 190 178 191
rect 176 190 177 191
rect 175 190 176 191
rect 174 190 175 191
rect 173 190 174 191
rect 172 190 173 191
rect 171 190 172 191
rect 170 190 171 191
rect 169 190 170 191
rect 168 190 169 191
rect 167 190 168 191
rect 166 190 167 191
rect 165 190 166 191
rect 164 190 165 191
rect 163 190 164 191
rect 162 190 163 191
rect 161 190 162 191
rect 160 190 161 191
rect 159 190 160 191
rect 158 190 159 191
rect 157 190 158 191
rect 156 190 157 191
rect 155 190 156 191
rect 154 190 155 191
rect 153 190 154 191
rect 152 190 153 191
rect 151 190 152 191
rect 150 190 151 191
rect 149 190 150 191
rect 148 190 149 191
rect 147 190 148 191
rect 146 190 147 191
rect 145 190 146 191
rect 144 190 145 191
rect 143 190 144 191
rect 142 190 143 191
rect 141 190 142 191
rect 140 190 141 191
rect 139 190 140 191
rect 138 190 139 191
rect 137 190 138 191
rect 136 190 137 191
rect 135 190 136 191
rect 134 190 135 191
rect 133 190 134 191
rect 132 190 133 191
rect 131 190 132 191
rect 130 190 131 191
rect 129 190 130 191
rect 128 190 129 191
rect 127 190 128 191
rect 126 190 127 191
rect 125 190 126 191
rect 124 190 125 191
rect 123 190 124 191
rect 122 190 123 191
rect 121 190 122 191
rect 120 190 121 191
rect 119 190 120 191
rect 118 190 119 191
rect 117 190 118 191
rect 116 190 117 191
rect 115 190 116 191
rect 114 190 115 191
rect 113 190 114 191
rect 112 190 113 191
rect 111 190 112 191
rect 110 190 111 191
rect 109 190 110 191
rect 108 190 109 191
rect 107 190 108 191
rect 106 190 107 191
rect 105 190 106 191
rect 104 190 105 191
rect 103 190 104 191
rect 102 190 103 191
rect 101 190 102 191
rect 100 190 101 191
rect 99 190 100 191
rect 98 190 99 191
rect 97 190 98 191
rect 96 190 97 191
rect 95 190 96 191
rect 94 190 95 191
rect 93 190 94 191
rect 92 190 93 191
rect 91 190 92 191
rect 90 190 91 191
rect 89 190 90 191
rect 88 190 89 191
rect 87 190 88 191
rect 86 190 87 191
rect 85 190 86 191
rect 84 190 85 191
rect 83 190 84 191
rect 82 190 83 191
rect 81 190 82 191
rect 80 190 81 191
rect 79 190 80 191
rect 78 190 79 191
rect 77 190 78 191
rect 76 190 77 191
rect 75 190 76 191
rect 74 190 75 191
rect 73 190 74 191
rect 72 190 73 191
rect 28 190 29 191
rect 27 190 28 191
rect 26 190 27 191
rect 25 190 26 191
rect 24 190 25 191
rect 23 190 24 191
rect 22 190 23 191
rect 21 190 22 191
rect 20 190 21 191
rect 19 190 20 191
rect 18 190 19 191
rect 17 190 18 191
rect 16 190 17 191
rect 15 190 16 191
rect 14 190 15 191
rect 437 191 438 192
rect 436 191 437 192
rect 435 191 436 192
rect 434 191 435 192
rect 433 191 434 192
rect 432 191 433 192
rect 431 191 432 192
rect 430 191 431 192
rect 429 191 430 192
rect 428 191 429 192
rect 427 191 428 192
rect 426 191 427 192
rect 425 191 426 192
rect 424 191 425 192
rect 423 191 424 192
rect 399 191 400 192
rect 398 191 399 192
rect 397 191 398 192
rect 340 191 341 192
rect 339 191 340 192
rect 338 191 339 192
rect 337 191 338 192
rect 336 191 337 192
rect 335 191 336 192
rect 334 191 335 192
rect 333 191 334 192
rect 332 191 333 192
rect 331 191 332 192
rect 330 191 331 192
rect 329 191 330 192
rect 328 191 329 192
rect 327 191 328 192
rect 326 191 327 192
rect 325 191 326 192
rect 324 191 325 192
rect 323 191 324 192
rect 322 191 323 192
rect 321 191 322 192
rect 320 191 321 192
rect 319 191 320 192
rect 318 191 319 192
rect 317 191 318 192
rect 316 191 317 192
rect 315 191 316 192
rect 314 191 315 192
rect 313 191 314 192
rect 312 191 313 192
rect 311 191 312 192
rect 310 191 311 192
rect 309 191 310 192
rect 308 191 309 192
rect 307 191 308 192
rect 306 191 307 192
rect 305 191 306 192
rect 304 191 305 192
rect 303 191 304 192
rect 302 191 303 192
rect 301 191 302 192
rect 300 191 301 192
rect 299 191 300 192
rect 298 191 299 192
rect 297 191 298 192
rect 296 191 297 192
rect 295 191 296 192
rect 294 191 295 192
rect 293 191 294 192
rect 292 191 293 192
rect 291 191 292 192
rect 290 191 291 192
rect 289 191 290 192
rect 288 191 289 192
rect 287 191 288 192
rect 286 191 287 192
rect 285 191 286 192
rect 284 191 285 192
rect 283 191 284 192
rect 282 191 283 192
rect 281 191 282 192
rect 280 191 281 192
rect 279 191 280 192
rect 278 191 279 192
rect 259 191 260 192
rect 258 191 259 192
rect 257 191 258 192
rect 256 191 257 192
rect 255 191 256 192
rect 254 191 255 192
rect 253 191 254 192
rect 252 191 253 192
rect 251 191 252 192
rect 250 191 251 192
rect 249 191 250 192
rect 248 191 249 192
rect 247 191 248 192
rect 246 191 247 192
rect 245 191 246 192
rect 244 191 245 192
rect 243 191 244 192
rect 242 191 243 192
rect 241 191 242 192
rect 240 191 241 192
rect 239 191 240 192
rect 238 191 239 192
rect 237 191 238 192
rect 236 191 237 192
rect 235 191 236 192
rect 234 191 235 192
rect 233 191 234 192
rect 232 191 233 192
rect 231 191 232 192
rect 230 191 231 192
rect 229 191 230 192
rect 228 191 229 192
rect 227 191 228 192
rect 226 191 227 192
rect 225 191 226 192
rect 224 191 225 192
rect 223 191 224 192
rect 222 191 223 192
rect 221 191 222 192
rect 220 191 221 192
rect 219 191 220 192
rect 196 191 197 192
rect 195 191 196 192
rect 194 191 195 192
rect 193 191 194 192
rect 192 191 193 192
rect 191 191 192 192
rect 190 191 191 192
rect 189 191 190 192
rect 188 191 189 192
rect 187 191 188 192
rect 186 191 187 192
rect 185 191 186 192
rect 184 191 185 192
rect 183 191 184 192
rect 182 191 183 192
rect 181 191 182 192
rect 180 191 181 192
rect 179 191 180 192
rect 178 191 179 192
rect 177 191 178 192
rect 176 191 177 192
rect 175 191 176 192
rect 174 191 175 192
rect 173 191 174 192
rect 172 191 173 192
rect 171 191 172 192
rect 170 191 171 192
rect 169 191 170 192
rect 168 191 169 192
rect 167 191 168 192
rect 166 191 167 192
rect 165 191 166 192
rect 164 191 165 192
rect 163 191 164 192
rect 162 191 163 192
rect 161 191 162 192
rect 160 191 161 192
rect 159 191 160 192
rect 158 191 159 192
rect 157 191 158 192
rect 156 191 157 192
rect 155 191 156 192
rect 154 191 155 192
rect 153 191 154 192
rect 152 191 153 192
rect 151 191 152 192
rect 150 191 151 192
rect 149 191 150 192
rect 148 191 149 192
rect 147 191 148 192
rect 146 191 147 192
rect 145 191 146 192
rect 144 191 145 192
rect 143 191 144 192
rect 142 191 143 192
rect 141 191 142 192
rect 140 191 141 192
rect 139 191 140 192
rect 138 191 139 192
rect 137 191 138 192
rect 136 191 137 192
rect 135 191 136 192
rect 134 191 135 192
rect 133 191 134 192
rect 132 191 133 192
rect 131 191 132 192
rect 130 191 131 192
rect 129 191 130 192
rect 128 191 129 192
rect 127 191 128 192
rect 126 191 127 192
rect 125 191 126 192
rect 124 191 125 192
rect 123 191 124 192
rect 122 191 123 192
rect 121 191 122 192
rect 120 191 121 192
rect 119 191 120 192
rect 118 191 119 192
rect 117 191 118 192
rect 116 191 117 192
rect 115 191 116 192
rect 114 191 115 192
rect 113 191 114 192
rect 112 191 113 192
rect 111 191 112 192
rect 110 191 111 192
rect 109 191 110 192
rect 108 191 109 192
rect 107 191 108 192
rect 106 191 107 192
rect 105 191 106 192
rect 104 191 105 192
rect 103 191 104 192
rect 102 191 103 192
rect 101 191 102 192
rect 100 191 101 192
rect 99 191 100 192
rect 98 191 99 192
rect 97 191 98 192
rect 96 191 97 192
rect 95 191 96 192
rect 94 191 95 192
rect 93 191 94 192
rect 92 191 93 192
rect 91 191 92 192
rect 90 191 91 192
rect 89 191 90 192
rect 88 191 89 192
rect 87 191 88 192
rect 86 191 87 192
rect 85 191 86 192
rect 84 191 85 192
rect 83 191 84 192
rect 82 191 83 192
rect 81 191 82 192
rect 80 191 81 192
rect 79 191 80 192
rect 78 191 79 192
rect 77 191 78 192
rect 76 191 77 192
rect 75 191 76 192
rect 74 191 75 192
rect 73 191 74 192
rect 72 191 73 192
rect 28 191 29 192
rect 27 191 28 192
rect 26 191 27 192
rect 25 191 26 192
rect 24 191 25 192
rect 23 191 24 192
rect 22 191 23 192
rect 21 191 22 192
rect 20 191 21 192
rect 19 191 20 192
rect 18 191 19 192
rect 17 191 18 192
rect 16 191 17 192
rect 15 191 16 192
rect 14 191 15 192
rect 482 192 483 193
rect 438 192 439 193
rect 437 192 438 193
rect 436 192 437 193
rect 435 192 436 193
rect 434 192 435 193
rect 433 192 434 193
rect 432 192 433 193
rect 431 192 432 193
rect 430 192 431 193
rect 429 192 430 193
rect 428 192 429 193
rect 427 192 428 193
rect 426 192 427 193
rect 425 192 426 193
rect 424 192 425 193
rect 399 192 400 193
rect 398 192 399 193
rect 397 192 398 193
rect 341 192 342 193
rect 340 192 341 193
rect 339 192 340 193
rect 338 192 339 193
rect 337 192 338 193
rect 336 192 337 193
rect 335 192 336 193
rect 334 192 335 193
rect 333 192 334 193
rect 332 192 333 193
rect 331 192 332 193
rect 330 192 331 193
rect 329 192 330 193
rect 328 192 329 193
rect 327 192 328 193
rect 326 192 327 193
rect 325 192 326 193
rect 324 192 325 193
rect 323 192 324 193
rect 322 192 323 193
rect 321 192 322 193
rect 320 192 321 193
rect 319 192 320 193
rect 318 192 319 193
rect 317 192 318 193
rect 316 192 317 193
rect 315 192 316 193
rect 314 192 315 193
rect 313 192 314 193
rect 312 192 313 193
rect 311 192 312 193
rect 310 192 311 193
rect 309 192 310 193
rect 308 192 309 193
rect 307 192 308 193
rect 306 192 307 193
rect 305 192 306 193
rect 304 192 305 193
rect 303 192 304 193
rect 302 192 303 193
rect 301 192 302 193
rect 300 192 301 193
rect 299 192 300 193
rect 298 192 299 193
rect 297 192 298 193
rect 296 192 297 193
rect 295 192 296 193
rect 294 192 295 193
rect 293 192 294 193
rect 292 192 293 193
rect 291 192 292 193
rect 290 192 291 193
rect 289 192 290 193
rect 288 192 289 193
rect 287 192 288 193
rect 286 192 287 193
rect 285 192 286 193
rect 284 192 285 193
rect 283 192 284 193
rect 282 192 283 193
rect 281 192 282 193
rect 280 192 281 193
rect 279 192 280 193
rect 278 192 279 193
rect 277 192 278 193
rect 258 192 259 193
rect 257 192 258 193
rect 256 192 257 193
rect 255 192 256 193
rect 254 192 255 193
rect 253 192 254 193
rect 252 192 253 193
rect 251 192 252 193
rect 250 192 251 193
rect 249 192 250 193
rect 248 192 249 193
rect 247 192 248 193
rect 246 192 247 193
rect 245 192 246 193
rect 244 192 245 193
rect 243 192 244 193
rect 242 192 243 193
rect 241 192 242 193
rect 240 192 241 193
rect 239 192 240 193
rect 238 192 239 193
rect 237 192 238 193
rect 236 192 237 193
rect 235 192 236 193
rect 234 192 235 193
rect 233 192 234 193
rect 232 192 233 193
rect 231 192 232 193
rect 230 192 231 193
rect 229 192 230 193
rect 228 192 229 193
rect 227 192 228 193
rect 226 192 227 193
rect 225 192 226 193
rect 224 192 225 193
rect 223 192 224 193
rect 222 192 223 193
rect 221 192 222 193
rect 220 192 221 193
rect 219 192 220 193
rect 218 192 219 193
rect 195 192 196 193
rect 194 192 195 193
rect 193 192 194 193
rect 192 192 193 193
rect 191 192 192 193
rect 190 192 191 193
rect 189 192 190 193
rect 188 192 189 193
rect 187 192 188 193
rect 186 192 187 193
rect 185 192 186 193
rect 184 192 185 193
rect 183 192 184 193
rect 182 192 183 193
rect 181 192 182 193
rect 180 192 181 193
rect 179 192 180 193
rect 178 192 179 193
rect 177 192 178 193
rect 176 192 177 193
rect 175 192 176 193
rect 174 192 175 193
rect 173 192 174 193
rect 172 192 173 193
rect 171 192 172 193
rect 170 192 171 193
rect 169 192 170 193
rect 168 192 169 193
rect 167 192 168 193
rect 166 192 167 193
rect 165 192 166 193
rect 164 192 165 193
rect 163 192 164 193
rect 162 192 163 193
rect 161 192 162 193
rect 160 192 161 193
rect 159 192 160 193
rect 158 192 159 193
rect 157 192 158 193
rect 156 192 157 193
rect 155 192 156 193
rect 154 192 155 193
rect 153 192 154 193
rect 152 192 153 193
rect 151 192 152 193
rect 150 192 151 193
rect 149 192 150 193
rect 148 192 149 193
rect 147 192 148 193
rect 146 192 147 193
rect 145 192 146 193
rect 144 192 145 193
rect 143 192 144 193
rect 142 192 143 193
rect 141 192 142 193
rect 140 192 141 193
rect 139 192 140 193
rect 138 192 139 193
rect 137 192 138 193
rect 136 192 137 193
rect 135 192 136 193
rect 134 192 135 193
rect 133 192 134 193
rect 132 192 133 193
rect 131 192 132 193
rect 130 192 131 193
rect 129 192 130 193
rect 128 192 129 193
rect 127 192 128 193
rect 126 192 127 193
rect 125 192 126 193
rect 124 192 125 193
rect 123 192 124 193
rect 122 192 123 193
rect 121 192 122 193
rect 120 192 121 193
rect 119 192 120 193
rect 118 192 119 193
rect 117 192 118 193
rect 116 192 117 193
rect 115 192 116 193
rect 114 192 115 193
rect 113 192 114 193
rect 112 192 113 193
rect 111 192 112 193
rect 110 192 111 193
rect 109 192 110 193
rect 108 192 109 193
rect 107 192 108 193
rect 106 192 107 193
rect 105 192 106 193
rect 104 192 105 193
rect 103 192 104 193
rect 102 192 103 193
rect 101 192 102 193
rect 100 192 101 193
rect 99 192 100 193
rect 98 192 99 193
rect 97 192 98 193
rect 96 192 97 193
rect 95 192 96 193
rect 94 192 95 193
rect 93 192 94 193
rect 92 192 93 193
rect 91 192 92 193
rect 90 192 91 193
rect 89 192 90 193
rect 88 192 89 193
rect 87 192 88 193
rect 86 192 87 193
rect 85 192 86 193
rect 84 192 85 193
rect 83 192 84 193
rect 82 192 83 193
rect 81 192 82 193
rect 80 192 81 193
rect 79 192 80 193
rect 78 192 79 193
rect 77 192 78 193
rect 76 192 77 193
rect 75 192 76 193
rect 74 192 75 193
rect 73 192 74 193
rect 72 192 73 193
rect 71 192 72 193
rect 29 192 30 193
rect 28 192 29 193
rect 27 192 28 193
rect 26 192 27 193
rect 25 192 26 193
rect 24 192 25 193
rect 23 192 24 193
rect 22 192 23 193
rect 21 192 22 193
rect 20 192 21 193
rect 19 192 20 193
rect 18 192 19 193
rect 17 192 18 193
rect 16 192 17 193
rect 15 192 16 193
rect 14 192 15 193
rect 482 193 483 194
rect 462 193 463 194
rect 439 193 440 194
rect 438 193 439 194
rect 437 193 438 194
rect 436 193 437 194
rect 435 193 436 194
rect 434 193 435 194
rect 433 193 434 194
rect 432 193 433 194
rect 431 193 432 194
rect 430 193 431 194
rect 429 193 430 194
rect 428 193 429 194
rect 427 193 428 194
rect 426 193 427 194
rect 425 193 426 194
rect 400 193 401 194
rect 399 193 400 194
rect 398 193 399 194
rect 397 193 398 194
rect 342 193 343 194
rect 341 193 342 194
rect 340 193 341 194
rect 339 193 340 194
rect 338 193 339 194
rect 337 193 338 194
rect 336 193 337 194
rect 335 193 336 194
rect 334 193 335 194
rect 333 193 334 194
rect 332 193 333 194
rect 331 193 332 194
rect 330 193 331 194
rect 329 193 330 194
rect 328 193 329 194
rect 327 193 328 194
rect 326 193 327 194
rect 325 193 326 194
rect 324 193 325 194
rect 323 193 324 194
rect 322 193 323 194
rect 321 193 322 194
rect 320 193 321 194
rect 319 193 320 194
rect 318 193 319 194
rect 317 193 318 194
rect 316 193 317 194
rect 315 193 316 194
rect 314 193 315 194
rect 313 193 314 194
rect 312 193 313 194
rect 311 193 312 194
rect 310 193 311 194
rect 309 193 310 194
rect 308 193 309 194
rect 307 193 308 194
rect 306 193 307 194
rect 305 193 306 194
rect 304 193 305 194
rect 303 193 304 194
rect 302 193 303 194
rect 301 193 302 194
rect 300 193 301 194
rect 299 193 300 194
rect 298 193 299 194
rect 297 193 298 194
rect 296 193 297 194
rect 295 193 296 194
rect 294 193 295 194
rect 293 193 294 194
rect 292 193 293 194
rect 291 193 292 194
rect 290 193 291 194
rect 289 193 290 194
rect 288 193 289 194
rect 287 193 288 194
rect 286 193 287 194
rect 285 193 286 194
rect 284 193 285 194
rect 283 193 284 194
rect 282 193 283 194
rect 281 193 282 194
rect 280 193 281 194
rect 279 193 280 194
rect 278 193 279 194
rect 277 193 278 194
rect 276 193 277 194
rect 275 193 276 194
rect 257 193 258 194
rect 256 193 257 194
rect 255 193 256 194
rect 254 193 255 194
rect 253 193 254 194
rect 252 193 253 194
rect 251 193 252 194
rect 250 193 251 194
rect 249 193 250 194
rect 248 193 249 194
rect 247 193 248 194
rect 246 193 247 194
rect 245 193 246 194
rect 244 193 245 194
rect 243 193 244 194
rect 242 193 243 194
rect 241 193 242 194
rect 240 193 241 194
rect 239 193 240 194
rect 238 193 239 194
rect 237 193 238 194
rect 236 193 237 194
rect 235 193 236 194
rect 234 193 235 194
rect 233 193 234 194
rect 232 193 233 194
rect 231 193 232 194
rect 230 193 231 194
rect 229 193 230 194
rect 228 193 229 194
rect 227 193 228 194
rect 226 193 227 194
rect 225 193 226 194
rect 224 193 225 194
rect 223 193 224 194
rect 222 193 223 194
rect 221 193 222 194
rect 220 193 221 194
rect 219 193 220 194
rect 218 193 219 194
rect 194 193 195 194
rect 193 193 194 194
rect 192 193 193 194
rect 191 193 192 194
rect 190 193 191 194
rect 189 193 190 194
rect 188 193 189 194
rect 187 193 188 194
rect 186 193 187 194
rect 185 193 186 194
rect 184 193 185 194
rect 183 193 184 194
rect 182 193 183 194
rect 181 193 182 194
rect 180 193 181 194
rect 179 193 180 194
rect 178 193 179 194
rect 177 193 178 194
rect 176 193 177 194
rect 175 193 176 194
rect 174 193 175 194
rect 173 193 174 194
rect 172 193 173 194
rect 171 193 172 194
rect 170 193 171 194
rect 169 193 170 194
rect 168 193 169 194
rect 167 193 168 194
rect 166 193 167 194
rect 165 193 166 194
rect 164 193 165 194
rect 163 193 164 194
rect 162 193 163 194
rect 161 193 162 194
rect 160 193 161 194
rect 159 193 160 194
rect 158 193 159 194
rect 157 193 158 194
rect 156 193 157 194
rect 155 193 156 194
rect 154 193 155 194
rect 153 193 154 194
rect 152 193 153 194
rect 151 193 152 194
rect 150 193 151 194
rect 149 193 150 194
rect 148 193 149 194
rect 147 193 148 194
rect 146 193 147 194
rect 145 193 146 194
rect 144 193 145 194
rect 143 193 144 194
rect 142 193 143 194
rect 141 193 142 194
rect 140 193 141 194
rect 139 193 140 194
rect 138 193 139 194
rect 137 193 138 194
rect 136 193 137 194
rect 135 193 136 194
rect 134 193 135 194
rect 133 193 134 194
rect 132 193 133 194
rect 131 193 132 194
rect 130 193 131 194
rect 129 193 130 194
rect 128 193 129 194
rect 127 193 128 194
rect 126 193 127 194
rect 125 193 126 194
rect 124 193 125 194
rect 123 193 124 194
rect 122 193 123 194
rect 121 193 122 194
rect 120 193 121 194
rect 119 193 120 194
rect 118 193 119 194
rect 117 193 118 194
rect 116 193 117 194
rect 115 193 116 194
rect 114 193 115 194
rect 113 193 114 194
rect 112 193 113 194
rect 111 193 112 194
rect 110 193 111 194
rect 109 193 110 194
rect 108 193 109 194
rect 107 193 108 194
rect 106 193 107 194
rect 105 193 106 194
rect 104 193 105 194
rect 103 193 104 194
rect 102 193 103 194
rect 101 193 102 194
rect 100 193 101 194
rect 99 193 100 194
rect 98 193 99 194
rect 97 193 98 194
rect 96 193 97 194
rect 95 193 96 194
rect 94 193 95 194
rect 93 193 94 194
rect 92 193 93 194
rect 91 193 92 194
rect 90 193 91 194
rect 89 193 90 194
rect 88 193 89 194
rect 87 193 88 194
rect 86 193 87 194
rect 85 193 86 194
rect 84 193 85 194
rect 83 193 84 194
rect 82 193 83 194
rect 81 193 82 194
rect 80 193 81 194
rect 79 193 80 194
rect 78 193 79 194
rect 77 193 78 194
rect 76 193 77 194
rect 75 193 76 194
rect 74 193 75 194
rect 73 193 74 194
rect 72 193 73 194
rect 71 193 72 194
rect 30 193 31 194
rect 29 193 30 194
rect 28 193 29 194
rect 27 193 28 194
rect 26 193 27 194
rect 25 193 26 194
rect 24 193 25 194
rect 23 193 24 194
rect 22 193 23 194
rect 21 193 22 194
rect 20 193 21 194
rect 19 193 20 194
rect 18 193 19 194
rect 17 193 18 194
rect 16 193 17 194
rect 15 193 16 194
rect 14 193 15 194
rect 482 194 483 195
rect 481 194 482 195
rect 462 194 463 195
rect 440 194 441 195
rect 439 194 440 195
rect 438 194 439 195
rect 437 194 438 195
rect 436 194 437 195
rect 435 194 436 195
rect 434 194 435 195
rect 433 194 434 195
rect 432 194 433 195
rect 431 194 432 195
rect 430 194 431 195
rect 429 194 430 195
rect 428 194 429 195
rect 427 194 428 195
rect 426 194 427 195
rect 401 194 402 195
rect 400 194 401 195
rect 399 194 400 195
rect 398 194 399 195
rect 397 194 398 195
rect 343 194 344 195
rect 342 194 343 195
rect 341 194 342 195
rect 340 194 341 195
rect 339 194 340 195
rect 338 194 339 195
rect 337 194 338 195
rect 336 194 337 195
rect 335 194 336 195
rect 334 194 335 195
rect 333 194 334 195
rect 332 194 333 195
rect 331 194 332 195
rect 330 194 331 195
rect 329 194 330 195
rect 328 194 329 195
rect 327 194 328 195
rect 326 194 327 195
rect 325 194 326 195
rect 324 194 325 195
rect 323 194 324 195
rect 322 194 323 195
rect 321 194 322 195
rect 320 194 321 195
rect 319 194 320 195
rect 318 194 319 195
rect 317 194 318 195
rect 316 194 317 195
rect 315 194 316 195
rect 314 194 315 195
rect 313 194 314 195
rect 312 194 313 195
rect 311 194 312 195
rect 310 194 311 195
rect 309 194 310 195
rect 308 194 309 195
rect 307 194 308 195
rect 306 194 307 195
rect 305 194 306 195
rect 304 194 305 195
rect 303 194 304 195
rect 302 194 303 195
rect 301 194 302 195
rect 300 194 301 195
rect 299 194 300 195
rect 298 194 299 195
rect 297 194 298 195
rect 296 194 297 195
rect 295 194 296 195
rect 294 194 295 195
rect 293 194 294 195
rect 292 194 293 195
rect 291 194 292 195
rect 290 194 291 195
rect 289 194 290 195
rect 288 194 289 195
rect 287 194 288 195
rect 286 194 287 195
rect 285 194 286 195
rect 284 194 285 195
rect 283 194 284 195
rect 282 194 283 195
rect 281 194 282 195
rect 280 194 281 195
rect 279 194 280 195
rect 278 194 279 195
rect 277 194 278 195
rect 276 194 277 195
rect 275 194 276 195
rect 274 194 275 195
rect 257 194 258 195
rect 256 194 257 195
rect 255 194 256 195
rect 254 194 255 195
rect 253 194 254 195
rect 252 194 253 195
rect 251 194 252 195
rect 250 194 251 195
rect 249 194 250 195
rect 248 194 249 195
rect 247 194 248 195
rect 246 194 247 195
rect 245 194 246 195
rect 244 194 245 195
rect 243 194 244 195
rect 242 194 243 195
rect 241 194 242 195
rect 240 194 241 195
rect 239 194 240 195
rect 238 194 239 195
rect 237 194 238 195
rect 236 194 237 195
rect 235 194 236 195
rect 234 194 235 195
rect 233 194 234 195
rect 232 194 233 195
rect 231 194 232 195
rect 230 194 231 195
rect 229 194 230 195
rect 228 194 229 195
rect 227 194 228 195
rect 226 194 227 195
rect 225 194 226 195
rect 224 194 225 195
rect 223 194 224 195
rect 222 194 223 195
rect 221 194 222 195
rect 220 194 221 195
rect 219 194 220 195
rect 218 194 219 195
rect 217 194 218 195
rect 193 194 194 195
rect 192 194 193 195
rect 191 194 192 195
rect 190 194 191 195
rect 189 194 190 195
rect 188 194 189 195
rect 187 194 188 195
rect 186 194 187 195
rect 185 194 186 195
rect 184 194 185 195
rect 183 194 184 195
rect 182 194 183 195
rect 181 194 182 195
rect 180 194 181 195
rect 179 194 180 195
rect 178 194 179 195
rect 177 194 178 195
rect 176 194 177 195
rect 175 194 176 195
rect 174 194 175 195
rect 173 194 174 195
rect 172 194 173 195
rect 171 194 172 195
rect 170 194 171 195
rect 169 194 170 195
rect 168 194 169 195
rect 167 194 168 195
rect 166 194 167 195
rect 165 194 166 195
rect 164 194 165 195
rect 163 194 164 195
rect 162 194 163 195
rect 161 194 162 195
rect 160 194 161 195
rect 159 194 160 195
rect 158 194 159 195
rect 157 194 158 195
rect 156 194 157 195
rect 155 194 156 195
rect 154 194 155 195
rect 153 194 154 195
rect 152 194 153 195
rect 151 194 152 195
rect 150 194 151 195
rect 149 194 150 195
rect 148 194 149 195
rect 147 194 148 195
rect 146 194 147 195
rect 145 194 146 195
rect 144 194 145 195
rect 143 194 144 195
rect 142 194 143 195
rect 141 194 142 195
rect 140 194 141 195
rect 139 194 140 195
rect 138 194 139 195
rect 137 194 138 195
rect 136 194 137 195
rect 135 194 136 195
rect 134 194 135 195
rect 133 194 134 195
rect 132 194 133 195
rect 131 194 132 195
rect 130 194 131 195
rect 129 194 130 195
rect 128 194 129 195
rect 127 194 128 195
rect 126 194 127 195
rect 125 194 126 195
rect 124 194 125 195
rect 123 194 124 195
rect 122 194 123 195
rect 121 194 122 195
rect 120 194 121 195
rect 119 194 120 195
rect 118 194 119 195
rect 117 194 118 195
rect 116 194 117 195
rect 115 194 116 195
rect 114 194 115 195
rect 113 194 114 195
rect 112 194 113 195
rect 111 194 112 195
rect 110 194 111 195
rect 109 194 110 195
rect 108 194 109 195
rect 107 194 108 195
rect 106 194 107 195
rect 105 194 106 195
rect 104 194 105 195
rect 103 194 104 195
rect 102 194 103 195
rect 101 194 102 195
rect 100 194 101 195
rect 99 194 100 195
rect 98 194 99 195
rect 97 194 98 195
rect 96 194 97 195
rect 95 194 96 195
rect 94 194 95 195
rect 93 194 94 195
rect 92 194 93 195
rect 91 194 92 195
rect 90 194 91 195
rect 89 194 90 195
rect 88 194 89 195
rect 87 194 88 195
rect 86 194 87 195
rect 85 194 86 195
rect 84 194 85 195
rect 83 194 84 195
rect 82 194 83 195
rect 81 194 82 195
rect 80 194 81 195
rect 79 194 80 195
rect 78 194 79 195
rect 77 194 78 195
rect 76 194 77 195
rect 75 194 76 195
rect 74 194 75 195
rect 73 194 74 195
rect 72 194 73 195
rect 71 194 72 195
rect 30 194 31 195
rect 29 194 30 195
rect 28 194 29 195
rect 27 194 28 195
rect 26 194 27 195
rect 25 194 26 195
rect 24 194 25 195
rect 23 194 24 195
rect 22 194 23 195
rect 21 194 22 195
rect 20 194 21 195
rect 19 194 20 195
rect 18 194 19 195
rect 17 194 18 195
rect 16 194 17 195
rect 15 194 16 195
rect 14 194 15 195
rect 482 195 483 196
rect 481 195 482 196
rect 480 195 481 196
rect 479 195 480 196
rect 478 195 479 196
rect 477 195 478 196
rect 476 195 477 196
rect 475 195 476 196
rect 474 195 475 196
rect 473 195 474 196
rect 472 195 473 196
rect 471 195 472 196
rect 470 195 471 196
rect 469 195 470 196
rect 468 195 469 196
rect 467 195 468 196
rect 466 195 467 196
rect 465 195 466 196
rect 464 195 465 196
rect 463 195 464 196
rect 462 195 463 196
rect 442 195 443 196
rect 441 195 442 196
rect 440 195 441 196
rect 439 195 440 196
rect 438 195 439 196
rect 437 195 438 196
rect 436 195 437 196
rect 435 195 436 196
rect 434 195 435 196
rect 433 195 434 196
rect 432 195 433 196
rect 431 195 432 196
rect 430 195 431 196
rect 429 195 430 196
rect 428 195 429 196
rect 427 195 428 196
rect 407 195 408 196
rect 406 195 407 196
rect 405 195 406 196
rect 404 195 405 196
rect 403 195 404 196
rect 402 195 403 196
rect 401 195 402 196
rect 400 195 401 196
rect 399 195 400 196
rect 398 195 399 196
rect 397 195 398 196
rect 344 195 345 196
rect 343 195 344 196
rect 342 195 343 196
rect 341 195 342 196
rect 340 195 341 196
rect 339 195 340 196
rect 338 195 339 196
rect 337 195 338 196
rect 336 195 337 196
rect 335 195 336 196
rect 334 195 335 196
rect 333 195 334 196
rect 332 195 333 196
rect 331 195 332 196
rect 330 195 331 196
rect 329 195 330 196
rect 328 195 329 196
rect 327 195 328 196
rect 326 195 327 196
rect 325 195 326 196
rect 324 195 325 196
rect 323 195 324 196
rect 322 195 323 196
rect 321 195 322 196
rect 320 195 321 196
rect 319 195 320 196
rect 318 195 319 196
rect 317 195 318 196
rect 316 195 317 196
rect 315 195 316 196
rect 314 195 315 196
rect 313 195 314 196
rect 312 195 313 196
rect 311 195 312 196
rect 310 195 311 196
rect 309 195 310 196
rect 308 195 309 196
rect 307 195 308 196
rect 306 195 307 196
rect 305 195 306 196
rect 304 195 305 196
rect 303 195 304 196
rect 302 195 303 196
rect 301 195 302 196
rect 300 195 301 196
rect 299 195 300 196
rect 298 195 299 196
rect 297 195 298 196
rect 296 195 297 196
rect 295 195 296 196
rect 294 195 295 196
rect 293 195 294 196
rect 292 195 293 196
rect 291 195 292 196
rect 290 195 291 196
rect 289 195 290 196
rect 288 195 289 196
rect 287 195 288 196
rect 286 195 287 196
rect 285 195 286 196
rect 284 195 285 196
rect 283 195 284 196
rect 282 195 283 196
rect 281 195 282 196
rect 280 195 281 196
rect 279 195 280 196
rect 278 195 279 196
rect 277 195 278 196
rect 276 195 277 196
rect 275 195 276 196
rect 274 195 275 196
rect 273 195 274 196
rect 256 195 257 196
rect 255 195 256 196
rect 254 195 255 196
rect 253 195 254 196
rect 252 195 253 196
rect 251 195 252 196
rect 250 195 251 196
rect 249 195 250 196
rect 248 195 249 196
rect 247 195 248 196
rect 246 195 247 196
rect 245 195 246 196
rect 244 195 245 196
rect 243 195 244 196
rect 242 195 243 196
rect 241 195 242 196
rect 240 195 241 196
rect 239 195 240 196
rect 238 195 239 196
rect 237 195 238 196
rect 236 195 237 196
rect 235 195 236 196
rect 234 195 235 196
rect 233 195 234 196
rect 232 195 233 196
rect 231 195 232 196
rect 230 195 231 196
rect 229 195 230 196
rect 228 195 229 196
rect 227 195 228 196
rect 226 195 227 196
rect 225 195 226 196
rect 224 195 225 196
rect 223 195 224 196
rect 222 195 223 196
rect 221 195 222 196
rect 220 195 221 196
rect 219 195 220 196
rect 218 195 219 196
rect 217 195 218 196
rect 216 195 217 196
rect 192 195 193 196
rect 191 195 192 196
rect 190 195 191 196
rect 189 195 190 196
rect 188 195 189 196
rect 187 195 188 196
rect 186 195 187 196
rect 185 195 186 196
rect 184 195 185 196
rect 183 195 184 196
rect 182 195 183 196
rect 181 195 182 196
rect 180 195 181 196
rect 179 195 180 196
rect 178 195 179 196
rect 177 195 178 196
rect 176 195 177 196
rect 175 195 176 196
rect 174 195 175 196
rect 173 195 174 196
rect 172 195 173 196
rect 171 195 172 196
rect 170 195 171 196
rect 169 195 170 196
rect 168 195 169 196
rect 167 195 168 196
rect 166 195 167 196
rect 165 195 166 196
rect 164 195 165 196
rect 163 195 164 196
rect 162 195 163 196
rect 161 195 162 196
rect 160 195 161 196
rect 159 195 160 196
rect 158 195 159 196
rect 157 195 158 196
rect 156 195 157 196
rect 155 195 156 196
rect 154 195 155 196
rect 153 195 154 196
rect 152 195 153 196
rect 151 195 152 196
rect 150 195 151 196
rect 149 195 150 196
rect 148 195 149 196
rect 147 195 148 196
rect 146 195 147 196
rect 145 195 146 196
rect 144 195 145 196
rect 143 195 144 196
rect 142 195 143 196
rect 141 195 142 196
rect 140 195 141 196
rect 139 195 140 196
rect 138 195 139 196
rect 137 195 138 196
rect 136 195 137 196
rect 135 195 136 196
rect 134 195 135 196
rect 133 195 134 196
rect 132 195 133 196
rect 131 195 132 196
rect 130 195 131 196
rect 129 195 130 196
rect 128 195 129 196
rect 127 195 128 196
rect 126 195 127 196
rect 125 195 126 196
rect 124 195 125 196
rect 123 195 124 196
rect 122 195 123 196
rect 121 195 122 196
rect 120 195 121 196
rect 119 195 120 196
rect 118 195 119 196
rect 117 195 118 196
rect 116 195 117 196
rect 115 195 116 196
rect 114 195 115 196
rect 113 195 114 196
rect 112 195 113 196
rect 111 195 112 196
rect 110 195 111 196
rect 109 195 110 196
rect 108 195 109 196
rect 107 195 108 196
rect 106 195 107 196
rect 105 195 106 196
rect 104 195 105 196
rect 103 195 104 196
rect 102 195 103 196
rect 101 195 102 196
rect 100 195 101 196
rect 99 195 100 196
rect 98 195 99 196
rect 97 195 98 196
rect 96 195 97 196
rect 95 195 96 196
rect 94 195 95 196
rect 93 195 94 196
rect 92 195 93 196
rect 91 195 92 196
rect 90 195 91 196
rect 89 195 90 196
rect 88 195 89 196
rect 87 195 88 196
rect 86 195 87 196
rect 85 195 86 196
rect 84 195 85 196
rect 83 195 84 196
rect 82 195 83 196
rect 81 195 82 196
rect 80 195 81 196
rect 79 195 80 196
rect 78 195 79 196
rect 77 195 78 196
rect 76 195 77 196
rect 75 195 76 196
rect 74 195 75 196
rect 73 195 74 196
rect 72 195 73 196
rect 52 195 53 196
rect 51 195 52 196
rect 50 195 51 196
rect 31 195 32 196
rect 30 195 31 196
rect 29 195 30 196
rect 28 195 29 196
rect 27 195 28 196
rect 26 195 27 196
rect 25 195 26 196
rect 24 195 25 196
rect 23 195 24 196
rect 22 195 23 196
rect 21 195 22 196
rect 20 195 21 196
rect 19 195 20 196
rect 18 195 19 196
rect 17 195 18 196
rect 16 195 17 196
rect 15 195 16 196
rect 14 195 15 196
rect 482 196 483 197
rect 481 196 482 197
rect 480 196 481 197
rect 479 196 480 197
rect 478 196 479 197
rect 477 196 478 197
rect 476 196 477 197
rect 475 196 476 197
rect 474 196 475 197
rect 473 196 474 197
rect 472 196 473 197
rect 471 196 472 197
rect 470 196 471 197
rect 469 196 470 197
rect 468 196 469 197
rect 467 196 468 197
rect 466 196 467 197
rect 465 196 466 197
rect 464 196 465 197
rect 463 196 464 197
rect 462 196 463 197
rect 442 196 443 197
rect 441 196 442 197
rect 440 196 441 197
rect 439 196 440 197
rect 438 196 439 197
rect 437 196 438 197
rect 436 196 437 197
rect 435 196 436 197
rect 434 196 435 197
rect 433 196 434 197
rect 432 196 433 197
rect 431 196 432 197
rect 430 196 431 197
rect 429 196 430 197
rect 428 196 429 197
rect 427 196 428 197
rect 426 196 427 197
rect 425 196 426 197
rect 424 196 425 197
rect 423 196 424 197
rect 422 196 423 197
rect 421 196 422 197
rect 420 196 421 197
rect 419 196 420 197
rect 418 196 419 197
rect 417 196 418 197
rect 416 196 417 197
rect 415 196 416 197
rect 414 196 415 197
rect 413 196 414 197
rect 412 196 413 197
rect 411 196 412 197
rect 410 196 411 197
rect 409 196 410 197
rect 408 196 409 197
rect 407 196 408 197
rect 406 196 407 197
rect 405 196 406 197
rect 404 196 405 197
rect 403 196 404 197
rect 402 196 403 197
rect 401 196 402 197
rect 400 196 401 197
rect 399 196 400 197
rect 398 196 399 197
rect 397 196 398 197
rect 345 196 346 197
rect 344 196 345 197
rect 343 196 344 197
rect 342 196 343 197
rect 341 196 342 197
rect 340 196 341 197
rect 339 196 340 197
rect 338 196 339 197
rect 337 196 338 197
rect 336 196 337 197
rect 335 196 336 197
rect 334 196 335 197
rect 333 196 334 197
rect 332 196 333 197
rect 331 196 332 197
rect 330 196 331 197
rect 329 196 330 197
rect 328 196 329 197
rect 327 196 328 197
rect 326 196 327 197
rect 325 196 326 197
rect 324 196 325 197
rect 323 196 324 197
rect 322 196 323 197
rect 321 196 322 197
rect 320 196 321 197
rect 319 196 320 197
rect 318 196 319 197
rect 317 196 318 197
rect 316 196 317 197
rect 315 196 316 197
rect 314 196 315 197
rect 313 196 314 197
rect 312 196 313 197
rect 311 196 312 197
rect 310 196 311 197
rect 309 196 310 197
rect 308 196 309 197
rect 307 196 308 197
rect 306 196 307 197
rect 305 196 306 197
rect 304 196 305 197
rect 303 196 304 197
rect 302 196 303 197
rect 301 196 302 197
rect 300 196 301 197
rect 299 196 300 197
rect 298 196 299 197
rect 297 196 298 197
rect 296 196 297 197
rect 295 196 296 197
rect 294 196 295 197
rect 293 196 294 197
rect 292 196 293 197
rect 291 196 292 197
rect 290 196 291 197
rect 289 196 290 197
rect 288 196 289 197
rect 287 196 288 197
rect 286 196 287 197
rect 285 196 286 197
rect 284 196 285 197
rect 283 196 284 197
rect 282 196 283 197
rect 281 196 282 197
rect 280 196 281 197
rect 279 196 280 197
rect 278 196 279 197
rect 277 196 278 197
rect 276 196 277 197
rect 275 196 276 197
rect 274 196 275 197
rect 273 196 274 197
rect 272 196 273 197
rect 271 196 272 197
rect 256 196 257 197
rect 255 196 256 197
rect 254 196 255 197
rect 253 196 254 197
rect 252 196 253 197
rect 251 196 252 197
rect 250 196 251 197
rect 249 196 250 197
rect 248 196 249 197
rect 247 196 248 197
rect 246 196 247 197
rect 245 196 246 197
rect 244 196 245 197
rect 243 196 244 197
rect 242 196 243 197
rect 241 196 242 197
rect 240 196 241 197
rect 239 196 240 197
rect 238 196 239 197
rect 237 196 238 197
rect 236 196 237 197
rect 235 196 236 197
rect 234 196 235 197
rect 233 196 234 197
rect 232 196 233 197
rect 231 196 232 197
rect 230 196 231 197
rect 229 196 230 197
rect 228 196 229 197
rect 227 196 228 197
rect 226 196 227 197
rect 225 196 226 197
rect 224 196 225 197
rect 223 196 224 197
rect 222 196 223 197
rect 221 196 222 197
rect 220 196 221 197
rect 219 196 220 197
rect 218 196 219 197
rect 217 196 218 197
rect 216 196 217 197
rect 191 196 192 197
rect 190 196 191 197
rect 189 196 190 197
rect 188 196 189 197
rect 187 196 188 197
rect 186 196 187 197
rect 185 196 186 197
rect 184 196 185 197
rect 183 196 184 197
rect 182 196 183 197
rect 181 196 182 197
rect 180 196 181 197
rect 179 196 180 197
rect 178 196 179 197
rect 177 196 178 197
rect 176 196 177 197
rect 175 196 176 197
rect 174 196 175 197
rect 173 196 174 197
rect 172 196 173 197
rect 171 196 172 197
rect 170 196 171 197
rect 169 196 170 197
rect 168 196 169 197
rect 167 196 168 197
rect 166 196 167 197
rect 165 196 166 197
rect 164 196 165 197
rect 163 196 164 197
rect 162 196 163 197
rect 161 196 162 197
rect 160 196 161 197
rect 159 196 160 197
rect 158 196 159 197
rect 157 196 158 197
rect 156 196 157 197
rect 155 196 156 197
rect 154 196 155 197
rect 153 196 154 197
rect 152 196 153 197
rect 151 196 152 197
rect 150 196 151 197
rect 149 196 150 197
rect 148 196 149 197
rect 147 196 148 197
rect 146 196 147 197
rect 145 196 146 197
rect 144 196 145 197
rect 143 196 144 197
rect 142 196 143 197
rect 141 196 142 197
rect 140 196 141 197
rect 139 196 140 197
rect 138 196 139 197
rect 137 196 138 197
rect 136 196 137 197
rect 135 196 136 197
rect 134 196 135 197
rect 133 196 134 197
rect 132 196 133 197
rect 131 196 132 197
rect 130 196 131 197
rect 129 196 130 197
rect 128 196 129 197
rect 127 196 128 197
rect 126 196 127 197
rect 125 196 126 197
rect 124 196 125 197
rect 123 196 124 197
rect 122 196 123 197
rect 121 196 122 197
rect 120 196 121 197
rect 119 196 120 197
rect 118 196 119 197
rect 117 196 118 197
rect 116 196 117 197
rect 115 196 116 197
rect 114 196 115 197
rect 113 196 114 197
rect 112 196 113 197
rect 111 196 112 197
rect 110 196 111 197
rect 109 196 110 197
rect 108 196 109 197
rect 107 196 108 197
rect 106 196 107 197
rect 105 196 106 197
rect 104 196 105 197
rect 103 196 104 197
rect 102 196 103 197
rect 101 196 102 197
rect 100 196 101 197
rect 99 196 100 197
rect 98 196 99 197
rect 97 196 98 197
rect 96 196 97 197
rect 95 196 96 197
rect 94 196 95 197
rect 93 196 94 197
rect 92 196 93 197
rect 91 196 92 197
rect 90 196 91 197
rect 89 196 90 197
rect 88 196 89 197
rect 87 196 88 197
rect 86 196 87 197
rect 85 196 86 197
rect 84 196 85 197
rect 83 196 84 197
rect 82 196 83 197
rect 81 196 82 197
rect 80 196 81 197
rect 79 196 80 197
rect 78 196 79 197
rect 77 196 78 197
rect 76 196 77 197
rect 75 196 76 197
rect 74 196 75 197
rect 73 196 74 197
rect 72 196 73 197
rect 53 196 54 197
rect 52 196 53 197
rect 51 196 52 197
rect 50 196 51 197
rect 49 196 50 197
rect 48 196 49 197
rect 33 196 34 197
rect 32 196 33 197
rect 31 196 32 197
rect 30 196 31 197
rect 29 196 30 197
rect 28 196 29 197
rect 27 196 28 197
rect 26 196 27 197
rect 25 196 26 197
rect 24 196 25 197
rect 23 196 24 197
rect 22 196 23 197
rect 21 196 22 197
rect 20 196 21 197
rect 19 196 20 197
rect 18 196 19 197
rect 17 196 18 197
rect 16 196 17 197
rect 15 196 16 197
rect 14 196 15 197
rect 482 197 483 198
rect 481 197 482 198
rect 480 197 481 198
rect 479 197 480 198
rect 478 197 479 198
rect 477 197 478 198
rect 476 197 477 198
rect 475 197 476 198
rect 474 197 475 198
rect 473 197 474 198
rect 472 197 473 198
rect 471 197 472 198
rect 470 197 471 198
rect 469 197 470 198
rect 468 197 469 198
rect 467 197 468 198
rect 466 197 467 198
rect 465 197 466 198
rect 464 197 465 198
rect 463 197 464 198
rect 462 197 463 198
rect 442 197 443 198
rect 441 197 442 198
rect 440 197 441 198
rect 439 197 440 198
rect 438 197 439 198
rect 437 197 438 198
rect 436 197 437 198
rect 435 197 436 198
rect 434 197 435 198
rect 433 197 434 198
rect 432 197 433 198
rect 431 197 432 198
rect 430 197 431 198
rect 429 197 430 198
rect 428 197 429 198
rect 427 197 428 198
rect 426 197 427 198
rect 425 197 426 198
rect 424 197 425 198
rect 423 197 424 198
rect 422 197 423 198
rect 421 197 422 198
rect 420 197 421 198
rect 419 197 420 198
rect 418 197 419 198
rect 417 197 418 198
rect 416 197 417 198
rect 415 197 416 198
rect 414 197 415 198
rect 413 197 414 198
rect 412 197 413 198
rect 411 197 412 198
rect 410 197 411 198
rect 409 197 410 198
rect 408 197 409 198
rect 407 197 408 198
rect 406 197 407 198
rect 405 197 406 198
rect 404 197 405 198
rect 403 197 404 198
rect 402 197 403 198
rect 401 197 402 198
rect 400 197 401 198
rect 399 197 400 198
rect 398 197 399 198
rect 397 197 398 198
rect 346 197 347 198
rect 345 197 346 198
rect 344 197 345 198
rect 343 197 344 198
rect 342 197 343 198
rect 341 197 342 198
rect 340 197 341 198
rect 339 197 340 198
rect 338 197 339 198
rect 337 197 338 198
rect 336 197 337 198
rect 335 197 336 198
rect 334 197 335 198
rect 333 197 334 198
rect 332 197 333 198
rect 331 197 332 198
rect 330 197 331 198
rect 329 197 330 198
rect 328 197 329 198
rect 327 197 328 198
rect 326 197 327 198
rect 325 197 326 198
rect 324 197 325 198
rect 323 197 324 198
rect 322 197 323 198
rect 321 197 322 198
rect 320 197 321 198
rect 319 197 320 198
rect 318 197 319 198
rect 317 197 318 198
rect 316 197 317 198
rect 315 197 316 198
rect 314 197 315 198
rect 313 197 314 198
rect 312 197 313 198
rect 311 197 312 198
rect 310 197 311 198
rect 309 197 310 198
rect 308 197 309 198
rect 307 197 308 198
rect 306 197 307 198
rect 305 197 306 198
rect 304 197 305 198
rect 303 197 304 198
rect 302 197 303 198
rect 301 197 302 198
rect 300 197 301 198
rect 299 197 300 198
rect 298 197 299 198
rect 297 197 298 198
rect 296 197 297 198
rect 295 197 296 198
rect 294 197 295 198
rect 293 197 294 198
rect 292 197 293 198
rect 291 197 292 198
rect 290 197 291 198
rect 289 197 290 198
rect 288 197 289 198
rect 287 197 288 198
rect 286 197 287 198
rect 285 197 286 198
rect 284 197 285 198
rect 283 197 284 198
rect 282 197 283 198
rect 281 197 282 198
rect 280 197 281 198
rect 279 197 280 198
rect 278 197 279 198
rect 277 197 278 198
rect 276 197 277 198
rect 275 197 276 198
rect 274 197 275 198
rect 273 197 274 198
rect 272 197 273 198
rect 271 197 272 198
rect 270 197 271 198
rect 255 197 256 198
rect 254 197 255 198
rect 253 197 254 198
rect 252 197 253 198
rect 251 197 252 198
rect 250 197 251 198
rect 249 197 250 198
rect 248 197 249 198
rect 247 197 248 198
rect 246 197 247 198
rect 245 197 246 198
rect 244 197 245 198
rect 243 197 244 198
rect 242 197 243 198
rect 241 197 242 198
rect 240 197 241 198
rect 239 197 240 198
rect 238 197 239 198
rect 237 197 238 198
rect 236 197 237 198
rect 235 197 236 198
rect 234 197 235 198
rect 233 197 234 198
rect 232 197 233 198
rect 231 197 232 198
rect 230 197 231 198
rect 229 197 230 198
rect 228 197 229 198
rect 227 197 228 198
rect 226 197 227 198
rect 225 197 226 198
rect 224 197 225 198
rect 223 197 224 198
rect 222 197 223 198
rect 221 197 222 198
rect 220 197 221 198
rect 219 197 220 198
rect 218 197 219 198
rect 217 197 218 198
rect 216 197 217 198
rect 215 197 216 198
rect 190 197 191 198
rect 189 197 190 198
rect 188 197 189 198
rect 187 197 188 198
rect 186 197 187 198
rect 185 197 186 198
rect 184 197 185 198
rect 183 197 184 198
rect 182 197 183 198
rect 181 197 182 198
rect 180 197 181 198
rect 179 197 180 198
rect 178 197 179 198
rect 177 197 178 198
rect 176 197 177 198
rect 175 197 176 198
rect 174 197 175 198
rect 173 197 174 198
rect 172 197 173 198
rect 171 197 172 198
rect 170 197 171 198
rect 169 197 170 198
rect 168 197 169 198
rect 167 197 168 198
rect 166 197 167 198
rect 165 197 166 198
rect 164 197 165 198
rect 163 197 164 198
rect 162 197 163 198
rect 161 197 162 198
rect 160 197 161 198
rect 159 197 160 198
rect 158 197 159 198
rect 157 197 158 198
rect 156 197 157 198
rect 155 197 156 198
rect 154 197 155 198
rect 153 197 154 198
rect 152 197 153 198
rect 151 197 152 198
rect 150 197 151 198
rect 149 197 150 198
rect 148 197 149 198
rect 147 197 148 198
rect 146 197 147 198
rect 145 197 146 198
rect 144 197 145 198
rect 143 197 144 198
rect 142 197 143 198
rect 141 197 142 198
rect 140 197 141 198
rect 139 197 140 198
rect 138 197 139 198
rect 137 197 138 198
rect 136 197 137 198
rect 135 197 136 198
rect 134 197 135 198
rect 133 197 134 198
rect 132 197 133 198
rect 131 197 132 198
rect 130 197 131 198
rect 129 197 130 198
rect 128 197 129 198
rect 127 197 128 198
rect 126 197 127 198
rect 125 197 126 198
rect 124 197 125 198
rect 123 197 124 198
rect 122 197 123 198
rect 121 197 122 198
rect 120 197 121 198
rect 119 197 120 198
rect 118 197 119 198
rect 117 197 118 198
rect 116 197 117 198
rect 115 197 116 198
rect 114 197 115 198
rect 113 197 114 198
rect 112 197 113 198
rect 111 197 112 198
rect 110 197 111 198
rect 109 197 110 198
rect 108 197 109 198
rect 107 197 108 198
rect 106 197 107 198
rect 105 197 106 198
rect 104 197 105 198
rect 103 197 104 198
rect 102 197 103 198
rect 101 197 102 198
rect 100 197 101 198
rect 99 197 100 198
rect 98 197 99 198
rect 97 197 98 198
rect 96 197 97 198
rect 95 197 96 198
rect 94 197 95 198
rect 93 197 94 198
rect 92 197 93 198
rect 91 197 92 198
rect 90 197 91 198
rect 89 197 90 198
rect 88 197 89 198
rect 87 197 88 198
rect 86 197 87 198
rect 85 197 86 198
rect 84 197 85 198
rect 83 197 84 198
rect 82 197 83 198
rect 81 197 82 198
rect 80 197 81 198
rect 79 197 80 198
rect 78 197 79 198
rect 77 197 78 198
rect 76 197 77 198
rect 75 197 76 198
rect 74 197 75 198
rect 73 197 74 198
rect 72 197 73 198
rect 53 197 54 198
rect 52 197 53 198
rect 51 197 52 198
rect 50 197 51 198
rect 49 197 50 198
rect 48 197 49 198
rect 47 197 48 198
rect 46 197 47 198
rect 34 197 35 198
rect 33 197 34 198
rect 32 197 33 198
rect 31 197 32 198
rect 30 197 31 198
rect 29 197 30 198
rect 28 197 29 198
rect 27 197 28 198
rect 26 197 27 198
rect 25 197 26 198
rect 24 197 25 198
rect 23 197 24 198
rect 22 197 23 198
rect 21 197 22 198
rect 20 197 21 198
rect 19 197 20 198
rect 18 197 19 198
rect 17 197 18 198
rect 16 197 17 198
rect 15 197 16 198
rect 14 197 15 198
rect 482 198 483 199
rect 481 198 482 199
rect 480 198 481 199
rect 479 198 480 199
rect 478 198 479 199
rect 477 198 478 199
rect 476 198 477 199
rect 475 198 476 199
rect 474 198 475 199
rect 473 198 474 199
rect 472 198 473 199
rect 471 198 472 199
rect 470 198 471 199
rect 469 198 470 199
rect 468 198 469 199
rect 467 198 468 199
rect 466 198 467 199
rect 465 198 466 199
rect 464 198 465 199
rect 463 198 464 199
rect 462 198 463 199
rect 442 198 443 199
rect 441 198 442 199
rect 440 198 441 199
rect 439 198 440 199
rect 438 198 439 199
rect 437 198 438 199
rect 436 198 437 199
rect 435 198 436 199
rect 434 198 435 199
rect 433 198 434 199
rect 432 198 433 199
rect 431 198 432 199
rect 430 198 431 199
rect 429 198 430 199
rect 428 198 429 199
rect 427 198 428 199
rect 426 198 427 199
rect 425 198 426 199
rect 424 198 425 199
rect 423 198 424 199
rect 422 198 423 199
rect 421 198 422 199
rect 420 198 421 199
rect 419 198 420 199
rect 418 198 419 199
rect 417 198 418 199
rect 416 198 417 199
rect 415 198 416 199
rect 414 198 415 199
rect 413 198 414 199
rect 412 198 413 199
rect 411 198 412 199
rect 410 198 411 199
rect 409 198 410 199
rect 408 198 409 199
rect 407 198 408 199
rect 406 198 407 199
rect 405 198 406 199
rect 404 198 405 199
rect 403 198 404 199
rect 402 198 403 199
rect 401 198 402 199
rect 400 198 401 199
rect 399 198 400 199
rect 398 198 399 199
rect 397 198 398 199
rect 347 198 348 199
rect 346 198 347 199
rect 345 198 346 199
rect 344 198 345 199
rect 343 198 344 199
rect 342 198 343 199
rect 341 198 342 199
rect 340 198 341 199
rect 339 198 340 199
rect 338 198 339 199
rect 337 198 338 199
rect 336 198 337 199
rect 335 198 336 199
rect 334 198 335 199
rect 333 198 334 199
rect 332 198 333 199
rect 331 198 332 199
rect 330 198 331 199
rect 329 198 330 199
rect 328 198 329 199
rect 327 198 328 199
rect 326 198 327 199
rect 325 198 326 199
rect 324 198 325 199
rect 323 198 324 199
rect 322 198 323 199
rect 321 198 322 199
rect 320 198 321 199
rect 319 198 320 199
rect 318 198 319 199
rect 317 198 318 199
rect 316 198 317 199
rect 315 198 316 199
rect 314 198 315 199
rect 313 198 314 199
rect 312 198 313 199
rect 311 198 312 199
rect 310 198 311 199
rect 309 198 310 199
rect 308 198 309 199
rect 307 198 308 199
rect 306 198 307 199
rect 305 198 306 199
rect 304 198 305 199
rect 303 198 304 199
rect 302 198 303 199
rect 301 198 302 199
rect 300 198 301 199
rect 299 198 300 199
rect 298 198 299 199
rect 297 198 298 199
rect 296 198 297 199
rect 295 198 296 199
rect 294 198 295 199
rect 293 198 294 199
rect 292 198 293 199
rect 291 198 292 199
rect 290 198 291 199
rect 289 198 290 199
rect 288 198 289 199
rect 287 198 288 199
rect 286 198 287 199
rect 285 198 286 199
rect 284 198 285 199
rect 283 198 284 199
rect 282 198 283 199
rect 281 198 282 199
rect 280 198 281 199
rect 279 198 280 199
rect 278 198 279 199
rect 277 198 278 199
rect 276 198 277 199
rect 275 198 276 199
rect 274 198 275 199
rect 273 198 274 199
rect 272 198 273 199
rect 271 198 272 199
rect 270 198 271 199
rect 269 198 270 199
rect 254 198 255 199
rect 253 198 254 199
rect 252 198 253 199
rect 251 198 252 199
rect 250 198 251 199
rect 249 198 250 199
rect 248 198 249 199
rect 247 198 248 199
rect 246 198 247 199
rect 245 198 246 199
rect 244 198 245 199
rect 243 198 244 199
rect 242 198 243 199
rect 241 198 242 199
rect 240 198 241 199
rect 239 198 240 199
rect 238 198 239 199
rect 237 198 238 199
rect 236 198 237 199
rect 235 198 236 199
rect 234 198 235 199
rect 233 198 234 199
rect 232 198 233 199
rect 231 198 232 199
rect 230 198 231 199
rect 229 198 230 199
rect 228 198 229 199
rect 227 198 228 199
rect 226 198 227 199
rect 225 198 226 199
rect 224 198 225 199
rect 223 198 224 199
rect 222 198 223 199
rect 221 198 222 199
rect 220 198 221 199
rect 219 198 220 199
rect 218 198 219 199
rect 217 198 218 199
rect 216 198 217 199
rect 215 198 216 199
rect 214 198 215 199
rect 189 198 190 199
rect 188 198 189 199
rect 187 198 188 199
rect 186 198 187 199
rect 185 198 186 199
rect 184 198 185 199
rect 183 198 184 199
rect 182 198 183 199
rect 181 198 182 199
rect 180 198 181 199
rect 179 198 180 199
rect 178 198 179 199
rect 177 198 178 199
rect 176 198 177 199
rect 175 198 176 199
rect 174 198 175 199
rect 173 198 174 199
rect 172 198 173 199
rect 171 198 172 199
rect 170 198 171 199
rect 169 198 170 199
rect 168 198 169 199
rect 167 198 168 199
rect 166 198 167 199
rect 165 198 166 199
rect 164 198 165 199
rect 163 198 164 199
rect 162 198 163 199
rect 161 198 162 199
rect 160 198 161 199
rect 159 198 160 199
rect 158 198 159 199
rect 157 198 158 199
rect 156 198 157 199
rect 155 198 156 199
rect 154 198 155 199
rect 153 198 154 199
rect 152 198 153 199
rect 151 198 152 199
rect 150 198 151 199
rect 149 198 150 199
rect 148 198 149 199
rect 147 198 148 199
rect 146 198 147 199
rect 145 198 146 199
rect 144 198 145 199
rect 143 198 144 199
rect 142 198 143 199
rect 141 198 142 199
rect 140 198 141 199
rect 139 198 140 199
rect 138 198 139 199
rect 137 198 138 199
rect 136 198 137 199
rect 135 198 136 199
rect 134 198 135 199
rect 133 198 134 199
rect 132 198 133 199
rect 131 198 132 199
rect 130 198 131 199
rect 129 198 130 199
rect 128 198 129 199
rect 127 198 128 199
rect 126 198 127 199
rect 125 198 126 199
rect 124 198 125 199
rect 123 198 124 199
rect 122 198 123 199
rect 121 198 122 199
rect 120 198 121 199
rect 119 198 120 199
rect 118 198 119 199
rect 117 198 118 199
rect 116 198 117 199
rect 115 198 116 199
rect 114 198 115 199
rect 113 198 114 199
rect 112 198 113 199
rect 111 198 112 199
rect 110 198 111 199
rect 109 198 110 199
rect 108 198 109 199
rect 107 198 108 199
rect 106 198 107 199
rect 105 198 106 199
rect 104 198 105 199
rect 103 198 104 199
rect 102 198 103 199
rect 101 198 102 199
rect 100 198 101 199
rect 99 198 100 199
rect 98 198 99 199
rect 97 198 98 199
rect 96 198 97 199
rect 95 198 96 199
rect 94 198 95 199
rect 93 198 94 199
rect 92 198 93 199
rect 91 198 92 199
rect 90 198 91 199
rect 89 198 90 199
rect 88 198 89 199
rect 87 198 88 199
rect 86 198 87 199
rect 85 198 86 199
rect 84 198 85 199
rect 83 198 84 199
rect 82 198 83 199
rect 81 198 82 199
rect 80 198 81 199
rect 79 198 80 199
rect 78 198 79 199
rect 77 198 78 199
rect 76 198 77 199
rect 75 198 76 199
rect 74 198 75 199
rect 73 198 74 199
rect 72 198 73 199
rect 54 198 55 199
rect 53 198 54 199
rect 52 198 53 199
rect 51 198 52 199
rect 50 198 51 199
rect 49 198 50 199
rect 48 198 49 199
rect 47 198 48 199
rect 46 198 47 199
rect 45 198 46 199
rect 44 198 45 199
rect 43 198 44 199
rect 42 198 43 199
rect 37 198 38 199
rect 36 198 37 199
rect 35 198 36 199
rect 34 198 35 199
rect 33 198 34 199
rect 32 198 33 199
rect 31 198 32 199
rect 30 198 31 199
rect 29 198 30 199
rect 28 198 29 199
rect 27 198 28 199
rect 26 198 27 199
rect 25 198 26 199
rect 24 198 25 199
rect 23 198 24 199
rect 22 198 23 199
rect 21 198 22 199
rect 20 198 21 199
rect 19 198 20 199
rect 18 198 19 199
rect 17 198 18 199
rect 16 198 17 199
rect 15 198 16 199
rect 14 198 15 199
rect 482 199 483 200
rect 481 199 482 200
rect 480 199 481 200
rect 479 199 480 200
rect 478 199 479 200
rect 477 199 478 200
rect 476 199 477 200
rect 475 199 476 200
rect 474 199 475 200
rect 473 199 474 200
rect 472 199 473 200
rect 471 199 472 200
rect 470 199 471 200
rect 469 199 470 200
rect 468 199 469 200
rect 467 199 468 200
rect 466 199 467 200
rect 465 199 466 200
rect 464 199 465 200
rect 463 199 464 200
rect 462 199 463 200
rect 407 199 408 200
rect 406 199 407 200
rect 405 199 406 200
rect 404 199 405 200
rect 403 199 404 200
rect 402 199 403 200
rect 401 199 402 200
rect 400 199 401 200
rect 399 199 400 200
rect 398 199 399 200
rect 397 199 398 200
rect 348 199 349 200
rect 347 199 348 200
rect 346 199 347 200
rect 345 199 346 200
rect 344 199 345 200
rect 343 199 344 200
rect 342 199 343 200
rect 341 199 342 200
rect 340 199 341 200
rect 339 199 340 200
rect 338 199 339 200
rect 337 199 338 200
rect 336 199 337 200
rect 335 199 336 200
rect 334 199 335 200
rect 333 199 334 200
rect 332 199 333 200
rect 331 199 332 200
rect 330 199 331 200
rect 329 199 330 200
rect 328 199 329 200
rect 327 199 328 200
rect 326 199 327 200
rect 325 199 326 200
rect 324 199 325 200
rect 323 199 324 200
rect 322 199 323 200
rect 321 199 322 200
rect 320 199 321 200
rect 319 199 320 200
rect 318 199 319 200
rect 317 199 318 200
rect 316 199 317 200
rect 315 199 316 200
rect 314 199 315 200
rect 313 199 314 200
rect 312 199 313 200
rect 311 199 312 200
rect 310 199 311 200
rect 309 199 310 200
rect 308 199 309 200
rect 307 199 308 200
rect 306 199 307 200
rect 305 199 306 200
rect 304 199 305 200
rect 303 199 304 200
rect 302 199 303 200
rect 301 199 302 200
rect 300 199 301 200
rect 299 199 300 200
rect 298 199 299 200
rect 297 199 298 200
rect 296 199 297 200
rect 295 199 296 200
rect 294 199 295 200
rect 293 199 294 200
rect 292 199 293 200
rect 291 199 292 200
rect 290 199 291 200
rect 289 199 290 200
rect 288 199 289 200
rect 287 199 288 200
rect 286 199 287 200
rect 285 199 286 200
rect 284 199 285 200
rect 283 199 284 200
rect 282 199 283 200
rect 281 199 282 200
rect 280 199 281 200
rect 279 199 280 200
rect 278 199 279 200
rect 277 199 278 200
rect 276 199 277 200
rect 275 199 276 200
rect 274 199 275 200
rect 273 199 274 200
rect 272 199 273 200
rect 271 199 272 200
rect 270 199 271 200
rect 269 199 270 200
rect 268 199 269 200
rect 267 199 268 200
rect 254 199 255 200
rect 253 199 254 200
rect 252 199 253 200
rect 251 199 252 200
rect 250 199 251 200
rect 249 199 250 200
rect 248 199 249 200
rect 247 199 248 200
rect 246 199 247 200
rect 245 199 246 200
rect 244 199 245 200
rect 243 199 244 200
rect 242 199 243 200
rect 241 199 242 200
rect 240 199 241 200
rect 239 199 240 200
rect 238 199 239 200
rect 237 199 238 200
rect 236 199 237 200
rect 235 199 236 200
rect 234 199 235 200
rect 233 199 234 200
rect 232 199 233 200
rect 231 199 232 200
rect 230 199 231 200
rect 229 199 230 200
rect 228 199 229 200
rect 227 199 228 200
rect 226 199 227 200
rect 225 199 226 200
rect 224 199 225 200
rect 223 199 224 200
rect 222 199 223 200
rect 221 199 222 200
rect 220 199 221 200
rect 219 199 220 200
rect 218 199 219 200
rect 217 199 218 200
rect 216 199 217 200
rect 215 199 216 200
rect 214 199 215 200
rect 213 199 214 200
rect 187 199 188 200
rect 186 199 187 200
rect 185 199 186 200
rect 184 199 185 200
rect 183 199 184 200
rect 182 199 183 200
rect 181 199 182 200
rect 180 199 181 200
rect 179 199 180 200
rect 178 199 179 200
rect 177 199 178 200
rect 176 199 177 200
rect 175 199 176 200
rect 174 199 175 200
rect 173 199 174 200
rect 172 199 173 200
rect 171 199 172 200
rect 170 199 171 200
rect 169 199 170 200
rect 168 199 169 200
rect 167 199 168 200
rect 166 199 167 200
rect 165 199 166 200
rect 164 199 165 200
rect 163 199 164 200
rect 162 199 163 200
rect 161 199 162 200
rect 160 199 161 200
rect 159 199 160 200
rect 158 199 159 200
rect 157 199 158 200
rect 156 199 157 200
rect 155 199 156 200
rect 154 199 155 200
rect 153 199 154 200
rect 152 199 153 200
rect 151 199 152 200
rect 150 199 151 200
rect 149 199 150 200
rect 148 199 149 200
rect 147 199 148 200
rect 146 199 147 200
rect 145 199 146 200
rect 144 199 145 200
rect 143 199 144 200
rect 142 199 143 200
rect 141 199 142 200
rect 140 199 141 200
rect 139 199 140 200
rect 138 199 139 200
rect 137 199 138 200
rect 136 199 137 200
rect 135 199 136 200
rect 134 199 135 200
rect 133 199 134 200
rect 132 199 133 200
rect 131 199 132 200
rect 130 199 131 200
rect 129 199 130 200
rect 128 199 129 200
rect 127 199 128 200
rect 126 199 127 200
rect 125 199 126 200
rect 124 199 125 200
rect 123 199 124 200
rect 122 199 123 200
rect 121 199 122 200
rect 120 199 121 200
rect 119 199 120 200
rect 118 199 119 200
rect 117 199 118 200
rect 116 199 117 200
rect 115 199 116 200
rect 114 199 115 200
rect 113 199 114 200
rect 112 199 113 200
rect 111 199 112 200
rect 110 199 111 200
rect 109 199 110 200
rect 108 199 109 200
rect 107 199 108 200
rect 106 199 107 200
rect 105 199 106 200
rect 104 199 105 200
rect 103 199 104 200
rect 102 199 103 200
rect 101 199 102 200
rect 100 199 101 200
rect 99 199 100 200
rect 98 199 99 200
rect 97 199 98 200
rect 96 199 97 200
rect 95 199 96 200
rect 94 199 95 200
rect 93 199 94 200
rect 92 199 93 200
rect 91 199 92 200
rect 90 199 91 200
rect 89 199 90 200
rect 88 199 89 200
rect 87 199 88 200
rect 86 199 87 200
rect 85 199 86 200
rect 84 199 85 200
rect 83 199 84 200
rect 82 199 83 200
rect 81 199 82 200
rect 80 199 81 200
rect 79 199 80 200
rect 78 199 79 200
rect 77 199 78 200
rect 76 199 77 200
rect 75 199 76 200
rect 74 199 75 200
rect 73 199 74 200
rect 72 199 73 200
rect 54 199 55 200
rect 53 199 54 200
rect 52 199 53 200
rect 51 199 52 200
rect 50 199 51 200
rect 49 199 50 200
rect 48 199 49 200
rect 47 199 48 200
rect 46 199 47 200
rect 45 199 46 200
rect 44 199 45 200
rect 43 199 44 200
rect 42 199 43 200
rect 41 199 42 200
rect 40 199 41 200
rect 39 199 40 200
rect 38 199 39 200
rect 37 199 38 200
rect 36 199 37 200
rect 35 199 36 200
rect 34 199 35 200
rect 33 199 34 200
rect 32 199 33 200
rect 31 199 32 200
rect 30 199 31 200
rect 29 199 30 200
rect 28 199 29 200
rect 27 199 28 200
rect 26 199 27 200
rect 25 199 26 200
rect 24 199 25 200
rect 23 199 24 200
rect 22 199 23 200
rect 21 199 22 200
rect 20 199 21 200
rect 19 199 20 200
rect 18 199 19 200
rect 17 199 18 200
rect 16 199 17 200
rect 15 199 16 200
rect 14 199 15 200
rect 482 200 483 201
rect 481 200 482 201
rect 472 200 473 201
rect 471 200 472 201
rect 462 200 463 201
rect 401 200 402 201
rect 400 200 401 201
rect 399 200 400 201
rect 398 200 399 201
rect 397 200 398 201
rect 349 200 350 201
rect 348 200 349 201
rect 347 200 348 201
rect 346 200 347 201
rect 345 200 346 201
rect 344 200 345 201
rect 343 200 344 201
rect 342 200 343 201
rect 341 200 342 201
rect 340 200 341 201
rect 339 200 340 201
rect 338 200 339 201
rect 337 200 338 201
rect 336 200 337 201
rect 335 200 336 201
rect 334 200 335 201
rect 333 200 334 201
rect 332 200 333 201
rect 331 200 332 201
rect 330 200 331 201
rect 329 200 330 201
rect 328 200 329 201
rect 327 200 328 201
rect 326 200 327 201
rect 325 200 326 201
rect 324 200 325 201
rect 323 200 324 201
rect 322 200 323 201
rect 321 200 322 201
rect 320 200 321 201
rect 319 200 320 201
rect 318 200 319 201
rect 317 200 318 201
rect 316 200 317 201
rect 315 200 316 201
rect 314 200 315 201
rect 313 200 314 201
rect 312 200 313 201
rect 311 200 312 201
rect 310 200 311 201
rect 309 200 310 201
rect 308 200 309 201
rect 307 200 308 201
rect 306 200 307 201
rect 305 200 306 201
rect 304 200 305 201
rect 303 200 304 201
rect 302 200 303 201
rect 301 200 302 201
rect 300 200 301 201
rect 299 200 300 201
rect 298 200 299 201
rect 297 200 298 201
rect 296 200 297 201
rect 295 200 296 201
rect 294 200 295 201
rect 293 200 294 201
rect 292 200 293 201
rect 291 200 292 201
rect 290 200 291 201
rect 289 200 290 201
rect 288 200 289 201
rect 287 200 288 201
rect 286 200 287 201
rect 285 200 286 201
rect 284 200 285 201
rect 283 200 284 201
rect 282 200 283 201
rect 281 200 282 201
rect 280 200 281 201
rect 279 200 280 201
rect 278 200 279 201
rect 277 200 278 201
rect 276 200 277 201
rect 275 200 276 201
rect 274 200 275 201
rect 273 200 274 201
rect 272 200 273 201
rect 271 200 272 201
rect 270 200 271 201
rect 269 200 270 201
rect 268 200 269 201
rect 267 200 268 201
rect 266 200 267 201
rect 253 200 254 201
rect 252 200 253 201
rect 251 200 252 201
rect 250 200 251 201
rect 249 200 250 201
rect 248 200 249 201
rect 247 200 248 201
rect 246 200 247 201
rect 245 200 246 201
rect 244 200 245 201
rect 243 200 244 201
rect 242 200 243 201
rect 241 200 242 201
rect 240 200 241 201
rect 239 200 240 201
rect 238 200 239 201
rect 237 200 238 201
rect 236 200 237 201
rect 235 200 236 201
rect 234 200 235 201
rect 233 200 234 201
rect 232 200 233 201
rect 231 200 232 201
rect 230 200 231 201
rect 229 200 230 201
rect 228 200 229 201
rect 227 200 228 201
rect 226 200 227 201
rect 225 200 226 201
rect 224 200 225 201
rect 223 200 224 201
rect 222 200 223 201
rect 221 200 222 201
rect 220 200 221 201
rect 219 200 220 201
rect 218 200 219 201
rect 217 200 218 201
rect 216 200 217 201
rect 215 200 216 201
rect 214 200 215 201
rect 213 200 214 201
rect 212 200 213 201
rect 186 200 187 201
rect 185 200 186 201
rect 184 200 185 201
rect 183 200 184 201
rect 182 200 183 201
rect 181 200 182 201
rect 180 200 181 201
rect 179 200 180 201
rect 178 200 179 201
rect 177 200 178 201
rect 176 200 177 201
rect 175 200 176 201
rect 174 200 175 201
rect 173 200 174 201
rect 172 200 173 201
rect 171 200 172 201
rect 170 200 171 201
rect 169 200 170 201
rect 168 200 169 201
rect 167 200 168 201
rect 166 200 167 201
rect 165 200 166 201
rect 164 200 165 201
rect 163 200 164 201
rect 162 200 163 201
rect 161 200 162 201
rect 160 200 161 201
rect 159 200 160 201
rect 158 200 159 201
rect 157 200 158 201
rect 156 200 157 201
rect 155 200 156 201
rect 154 200 155 201
rect 153 200 154 201
rect 152 200 153 201
rect 151 200 152 201
rect 150 200 151 201
rect 149 200 150 201
rect 148 200 149 201
rect 147 200 148 201
rect 146 200 147 201
rect 145 200 146 201
rect 144 200 145 201
rect 143 200 144 201
rect 142 200 143 201
rect 141 200 142 201
rect 140 200 141 201
rect 139 200 140 201
rect 138 200 139 201
rect 137 200 138 201
rect 136 200 137 201
rect 135 200 136 201
rect 134 200 135 201
rect 133 200 134 201
rect 132 200 133 201
rect 131 200 132 201
rect 130 200 131 201
rect 129 200 130 201
rect 128 200 129 201
rect 127 200 128 201
rect 126 200 127 201
rect 125 200 126 201
rect 124 200 125 201
rect 123 200 124 201
rect 122 200 123 201
rect 121 200 122 201
rect 120 200 121 201
rect 119 200 120 201
rect 118 200 119 201
rect 117 200 118 201
rect 116 200 117 201
rect 115 200 116 201
rect 114 200 115 201
rect 113 200 114 201
rect 112 200 113 201
rect 111 200 112 201
rect 110 200 111 201
rect 109 200 110 201
rect 108 200 109 201
rect 107 200 108 201
rect 106 200 107 201
rect 105 200 106 201
rect 104 200 105 201
rect 103 200 104 201
rect 102 200 103 201
rect 101 200 102 201
rect 100 200 101 201
rect 99 200 100 201
rect 98 200 99 201
rect 97 200 98 201
rect 96 200 97 201
rect 95 200 96 201
rect 94 200 95 201
rect 93 200 94 201
rect 92 200 93 201
rect 91 200 92 201
rect 90 200 91 201
rect 89 200 90 201
rect 88 200 89 201
rect 87 200 88 201
rect 86 200 87 201
rect 85 200 86 201
rect 84 200 85 201
rect 83 200 84 201
rect 82 200 83 201
rect 81 200 82 201
rect 80 200 81 201
rect 79 200 80 201
rect 78 200 79 201
rect 77 200 78 201
rect 76 200 77 201
rect 75 200 76 201
rect 74 200 75 201
rect 73 200 74 201
rect 55 200 56 201
rect 54 200 55 201
rect 53 200 54 201
rect 52 200 53 201
rect 51 200 52 201
rect 50 200 51 201
rect 49 200 50 201
rect 48 200 49 201
rect 47 200 48 201
rect 46 200 47 201
rect 45 200 46 201
rect 44 200 45 201
rect 43 200 44 201
rect 42 200 43 201
rect 41 200 42 201
rect 40 200 41 201
rect 39 200 40 201
rect 38 200 39 201
rect 37 200 38 201
rect 36 200 37 201
rect 35 200 36 201
rect 34 200 35 201
rect 33 200 34 201
rect 32 200 33 201
rect 31 200 32 201
rect 30 200 31 201
rect 29 200 30 201
rect 28 200 29 201
rect 27 200 28 201
rect 26 200 27 201
rect 25 200 26 201
rect 24 200 25 201
rect 23 200 24 201
rect 22 200 23 201
rect 21 200 22 201
rect 20 200 21 201
rect 19 200 20 201
rect 18 200 19 201
rect 17 200 18 201
rect 16 200 17 201
rect 15 200 16 201
rect 14 200 15 201
rect 13 200 14 201
rect 482 201 483 202
rect 472 201 473 202
rect 471 201 472 202
rect 462 201 463 202
rect 400 201 401 202
rect 399 201 400 202
rect 398 201 399 202
rect 397 201 398 202
rect 350 201 351 202
rect 349 201 350 202
rect 348 201 349 202
rect 347 201 348 202
rect 346 201 347 202
rect 345 201 346 202
rect 344 201 345 202
rect 343 201 344 202
rect 342 201 343 202
rect 341 201 342 202
rect 340 201 341 202
rect 339 201 340 202
rect 338 201 339 202
rect 337 201 338 202
rect 336 201 337 202
rect 335 201 336 202
rect 334 201 335 202
rect 333 201 334 202
rect 332 201 333 202
rect 331 201 332 202
rect 330 201 331 202
rect 329 201 330 202
rect 328 201 329 202
rect 327 201 328 202
rect 326 201 327 202
rect 325 201 326 202
rect 324 201 325 202
rect 323 201 324 202
rect 322 201 323 202
rect 321 201 322 202
rect 320 201 321 202
rect 319 201 320 202
rect 318 201 319 202
rect 317 201 318 202
rect 316 201 317 202
rect 315 201 316 202
rect 314 201 315 202
rect 313 201 314 202
rect 312 201 313 202
rect 311 201 312 202
rect 310 201 311 202
rect 309 201 310 202
rect 308 201 309 202
rect 307 201 308 202
rect 306 201 307 202
rect 305 201 306 202
rect 304 201 305 202
rect 303 201 304 202
rect 302 201 303 202
rect 301 201 302 202
rect 300 201 301 202
rect 299 201 300 202
rect 298 201 299 202
rect 297 201 298 202
rect 296 201 297 202
rect 295 201 296 202
rect 294 201 295 202
rect 293 201 294 202
rect 292 201 293 202
rect 291 201 292 202
rect 290 201 291 202
rect 289 201 290 202
rect 288 201 289 202
rect 287 201 288 202
rect 286 201 287 202
rect 285 201 286 202
rect 284 201 285 202
rect 283 201 284 202
rect 282 201 283 202
rect 281 201 282 202
rect 280 201 281 202
rect 279 201 280 202
rect 278 201 279 202
rect 277 201 278 202
rect 276 201 277 202
rect 275 201 276 202
rect 274 201 275 202
rect 273 201 274 202
rect 272 201 273 202
rect 271 201 272 202
rect 270 201 271 202
rect 269 201 270 202
rect 268 201 269 202
rect 267 201 268 202
rect 266 201 267 202
rect 265 201 266 202
rect 252 201 253 202
rect 251 201 252 202
rect 250 201 251 202
rect 249 201 250 202
rect 248 201 249 202
rect 247 201 248 202
rect 246 201 247 202
rect 245 201 246 202
rect 244 201 245 202
rect 243 201 244 202
rect 242 201 243 202
rect 241 201 242 202
rect 240 201 241 202
rect 239 201 240 202
rect 238 201 239 202
rect 237 201 238 202
rect 236 201 237 202
rect 235 201 236 202
rect 234 201 235 202
rect 233 201 234 202
rect 232 201 233 202
rect 231 201 232 202
rect 230 201 231 202
rect 229 201 230 202
rect 228 201 229 202
rect 227 201 228 202
rect 226 201 227 202
rect 225 201 226 202
rect 224 201 225 202
rect 223 201 224 202
rect 222 201 223 202
rect 221 201 222 202
rect 220 201 221 202
rect 219 201 220 202
rect 218 201 219 202
rect 217 201 218 202
rect 216 201 217 202
rect 215 201 216 202
rect 214 201 215 202
rect 213 201 214 202
rect 212 201 213 202
rect 185 201 186 202
rect 184 201 185 202
rect 183 201 184 202
rect 182 201 183 202
rect 181 201 182 202
rect 180 201 181 202
rect 179 201 180 202
rect 178 201 179 202
rect 177 201 178 202
rect 176 201 177 202
rect 175 201 176 202
rect 174 201 175 202
rect 173 201 174 202
rect 172 201 173 202
rect 171 201 172 202
rect 170 201 171 202
rect 169 201 170 202
rect 168 201 169 202
rect 167 201 168 202
rect 166 201 167 202
rect 165 201 166 202
rect 164 201 165 202
rect 163 201 164 202
rect 162 201 163 202
rect 161 201 162 202
rect 160 201 161 202
rect 159 201 160 202
rect 158 201 159 202
rect 157 201 158 202
rect 156 201 157 202
rect 155 201 156 202
rect 154 201 155 202
rect 153 201 154 202
rect 152 201 153 202
rect 151 201 152 202
rect 150 201 151 202
rect 149 201 150 202
rect 148 201 149 202
rect 147 201 148 202
rect 146 201 147 202
rect 145 201 146 202
rect 144 201 145 202
rect 143 201 144 202
rect 142 201 143 202
rect 141 201 142 202
rect 140 201 141 202
rect 139 201 140 202
rect 138 201 139 202
rect 137 201 138 202
rect 136 201 137 202
rect 135 201 136 202
rect 134 201 135 202
rect 133 201 134 202
rect 132 201 133 202
rect 131 201 132 202
rect 130 201 131 202
rect 129 201 130 202
rect 128 201 129 202
rect 127 201 128 202
rect 126 201 127 202
rect 125 201 126 202
rect 124 201 125 202
rect 123 201 124 202
rect 122 201 123 202
rect 121 201 122 202
rect 120 201 121 202
rect 119 201 120 202
rect 118 201 119 202
rect 117 201 118 202
rect 116 201 117 202
rect 115 201 116 202
rect 114 201 115 202
rect 113 201 114 202
rect 112 201 113 202
rect 111 201 112 202
rect 110 201 111 202
rect 109 201 110 202
rect 108 201 109 202
rect 107 201 108 202
rect 106 201 107 202
rect 105 201 106 202
rect 104 201 105 202
rect 103 201 104 202
rect 102 201 103 202
rect 101 201 102 202
rect 100 201 101 202
rect 99 201 100 202
rect 98 201 99 202
rect 97 201 98 202
rect 96 201 97 202
rect 95 201 96 202
rect 94 201 95 202
rect 93 201 94 202
rect 92 201 93 202
rect 91 201 92 202
rect 90 201 91 202
rect 89 201 90 202
rect 88 201 89 202
rect 87 201 88 202
rect 86 201 87 202
rect 85 201 86 202
rect 84 201 85 202
rect 83 201 84 202
rect 82 201 83 202
rect 81 201 82 202
rect 80 201 81 202
rect 79 201 80 202
rect 78 201 79 202
rect 77 201 78 202
rect 76 201 77 202
rect 75 201 76 202
rect 74 201 75 202
rect 73 201 74 202
rect 56 201 57 202
rect 55 201 56 202
rect 54 201 55 202
rect 53 201 54 202
rect 52 201 53 202
rect 51 201 52 202
rect 50 201 51 202
rect 49 201 50 202
rect 48 201 49 202
rect 47 201 48 202
rect 46 201 47 202
rect 45 201 46 202
rect 44 201 45 202
rect 43 201 44 202
rect 42 201 43 202
rect 41 201 42 202
rect 40 201 41 202
rect 39 201 40 202
rect 38 201 39 202
rect 37 201 38 202
rect 36 201 37 202
rect 35 201 36 202
rect 34 201 35 202
rect 33 201 34 202
rect 32 201 33 202
rect 31 201 32 202
rect 30 201 31 202
rect 29 201 30 202
rect 28 201 29 202
rect 27 201 28 202
rect 26 201 27 202
rect 25 201 26 202
rect 24 201 25 202
rect 23 201 24 202
rect 22 201 23 202
rect 21 201 22 202
rect 20 201 21 202
rect 19 201 20 202
rect 18 201 19 202
rect 17 201 18 202
rect 16 201 17 202
rect 15 201 16 202
rect 14 201 15 202
rect 13 201 14 202
rect 482 202 483 203
rect 472 202 473 203
rect 471 202 472 203
rect 462 202 463 203
rect 399 202 400 203
rect 398 202 399 203
rect 397 202 398 203
rect 351 202 352 203
rect 350 202 351 203
rect 349 202 350 203
rect 348 202 349 203
rect 347 202 348 203
rect 346 202 347 203
rect 345 202 346 203
rect 344 202 345 203
rect 343 202 344 203
rect 342 202 343 203
rect 341 202 342 203
rect 340 202 341 203
rect 339 202 340 203
rect 338 202 339 203
rect 337 202 338 203
rect 336 202 337 203
rect 335 202 336 203
rect 334 202 335 203
rect 333 202 334 203
rect 332 202 333 203
rect 331 202 332 203
rect 330 202 331 203
rect 329 202 330 203
rect 328 202 329 203
rect 327 202 328 203
rect 326 202 327 203
rect 325 202 326 203
rect 324 202 325 203
rect 323 202 324 203
rect 322 202 323 203
rect 321 202 322 203
rect 320 202 321 203
rect 319 202 320 203
rect 318 202 319 203
rect 317 202 318 203
rect 316 202 317 203
rect 315 202 316 203
rect 314 202 315 203
rect 313 202 314 203
rect 312 202 313 203
rect 311 202 312 203
rect 310 202 311 203
rect 309 202 310 203
rect 308 202 309 203
rect 307 202 308 203
rect 306 202 307 203
rect 305 202 306 203
rect 304 202 305 203
rect 303 202 304 203
rect 302 202 303 203
rect 301 202 302 203
rect 300 202 301 203
rect 299 202 300 203
rect 298 202 299 203
rect 297 202 298 203
rect 296 202 297 203
rect 295 202 296 203
rect 294 202 295 203
rect 293 202 294 203
rect 292 202 293 203
rect 291 202 292 203
rect 290 202 291 203
rect 289 202 290 203
rect 288 202 289 203
rect 287 202 288 203
rect 286 202 287 203
rect 285 202 286 203
rect 284 202 285 203
rect 283 202 284 203
rect 282 202 283 203
rect 281 202 282 203
rect 280 202 281 203
rect 279 202 280 203
rect 278 202 279 203
rect 277 202 278 203
rect 276 202 277 203
rect 275 202 276 203
rect 274 202 275 203
rect 273 202 274 203
rect 272 202 273 203
rect 271 202 272 203
rect 270 202 271 203
rect 269 202 270 203
rect 268 202 269 203
rect 267 202 268 203
rect 266 202 267 203
rect 265 202 266 203
rect 264 202 265 203
rect 263 202 264 203
rect 252 202 253 203
rect 251 202 252 203
rect 250 202 251 203
rect 249 202 250 203
rect 248 202 249 203
rect 247 202 248 203
rect 246 202 247 203
rect 245 202 246 203
rect 244 202 245 203
rect 243 202 244 203
rect 242 202 243 203
rect 241 202 242 203
rect 240 202 241 203
rect 239 202 240 203
rect 238 202 239 203
rect 237 202 238 203
rect 236 202 237 203
rect 235 202 236 203
rect 234 202 235 203
rect 233 202 234 203
rect 232 202 233 203
rect 231 202 232 203
rect 230 202 231 203
rect 229 202 230 203
rect 228 202 229 203
rect 227 202 228 203
rect 226 202 227 203
rect 225 202 226 203
rect 224 202 225 203
rect 223 202 224 203
rect 222 202 223 203
rect 221 202 222 203
rect 220 202 221 203
rect 219 202 220 203
rect 218 202 219 203
rect 217 202 218 203
rect 216 202 217 203
rect 215 202 216 203
rect 214 202 215 203
rect 213 202 214 203
rect 212 202 213 203
rect 211 202 212 203
rect 184 202 185 203
rect 183 202 184 203
rect 182 202 183 203
rect 181 202 182 203
rect 180 202 181 203
rect 179 202 180 203
rect 178 202 179 203
rect 177 202 178 203
rect 176 202 177 203
rect 175 202 176 203
rect 174 202 175 203
rect 173 202 174 203
rect 172 202 173 203
rect 171 202 172 203
rect 170 202 171 203
rect 169 202 170 203
rect 168 202 169 203
rect 167 202 168 203
rect 166 202 167 203
rect 165 202 166 203
rect 164 202 165 203
rect 163 202 164 203
rect 162 202 163 203
rect 161 202 162 203
rect 160 202 161 203
rect 159 202 160 203
rect 158 202 159 203
rect 157 202 158 203
rect 156 202 157 203
rect 155 202 156 203
rect 154 202 155 203
rect 153 202 154 203
rect 152 202 153 203
rect 151 202 152 203
rect 150 202 151 203
rect 149 202 150 203
rect 148 202 149 203
rect 147 202 148 203
rect 146 202 147 203
rect 145 202 146 203
rect 144 202 145 203
rect 143 202 144 203
rect 142 202 143 203
rect 141 202 142 203
rect 140 202 141 203
rect 139 202 140 203
rect 138 202 139 203
rect 137 202 138 203
rect 136 202 137 203
rect 135 202 136 203
rect 134 202 135 203
rect 133 202 134 203
rect 132 202 133 203
rect 131 202 132 203
rect 130 202 131 203
rect 129 202 130 203
rect 128 202 129 203
rect 127 202 128 203
rect 126 202 127 203
rect 125 202 126 203
rect 124 202 125 203
rect 123 202 124 203
rect 122 202 123 203
rect 121 202 122 203
rect 120 202 121 203
rect 119 202 120 203
rect 118 202 119 203
rect 117 202 118 203
rect 116 202 117 203
rect 115 202 116 203
rect 114 202 115 203
rect 113 202 114 203
rect 112 202 113 203
rect 111 202 112 203
rect 110 202 111 203
rect 109 202 110 203
rect 108 202 109 203
rect 107 202 108 203
rect 106 202 107 203
rect 105 202 106 203
rect 104 202 105 203
rect 103 202 104 203
rect 102 202 103 203
rect 101 202 102 203
rect 100 202 101 203
rect 99 202 100 203
rect 98 202 99 203
rect 97 202 98 203
rect 96 202 97 203
rect 95 202 96 203
rect 94 202 95 203
rect 93 202 94 203
rect 92 202 93 203
rect 91 202 92 203
rect 90 202 91 203
rect 89 202 90 203
rect 88 202 89 203
rect 87 202 88 203
rect 86 202 87 203
rect 85 202 86 203
rect 84 202 85 203
rect 83 202 84 203
rect 82 202 83 203
rect 81 202 82 203
rect 80 202 81 203
rect 79 202 80 203
rect 78 202 79 203
rect 77 202 78 203
rect 76 202 77 203
rect 75 202 76 203
rect 74 202 75 203
rect 73 202 74 203
rect 56 202 57 203
rect 55 202 56 203
rect 54 202 55 203
rect 53 202 54 203
rect 52 202 53 203
rect 51 202 52 203
rect 50 202 51 203
rect 49 202 50 203
rect 48 202 49 203
rect 47 202 48 203
rect 46 202 47 203
rect 45 202 46 203
rect 44 202 45 203
rect 43 202 44 203
rect 42 202 43 203
rect 41 202 42 203
rect 40 202 41 203
rect 39 202 40 203
rect 38 202 39 203
rect 37 202 38 203
rect 36 202 37 203
rect 35 202 36 203
rect 34 202 35 203
rect 33 202 34 203
rect 32 202 33 203
rect 31 202 32 203
rect 30 202 31 203
rect 29 202 30 203
rect 28 202 29 203
rect 27 202 28 203
rect 26 202 27 203
rect 25 202 26 203
rect 24 202 25 203
rect 23 202 24 203
rect 22 202 23 203
rect 21 202 22 203
rect 20 202 21 203
rect 19 202 20 203
rect 18 202 19 203
rect 17 202 18 203
rect 16 202 17 203
rect 15 202 16 203
rect 14 202 15 203
rect 13 202 14 203
rect 482 203 483 204
rect 472 203 473 204
rect 471 203 472 204
rect 462 203 463 204
rect 399 203 400 204
rect 398 203 399 204
rect 397 203 398 204
rect 352 203 353 204
rect 351 203 352 204
rect 350 203 351 204
rect 349 203 350 204
rect 348 203 349 204
rect 347 203 348 204
rect 346 203 347 204
rect 345 203 346 204
rect 344 203 345 204
rect 343 203 344 204
rect 342 203 343 204
rect 341 203 342 204
rect 340 203 341 204
rect 339 203 340 204
rect 338 203 339 204
rect 337 203 338 204
rect 336 203 337 204
rect 335 203 336 204
rect 334 203 335 204
rect 333 203 334 204
rect 332 203 333 204
rect 331 203 332 204
rect 330 203 331 204
rect 329 203 330 204
rect 328 203 329 204
rect 327 203 328 204
rect 326 203 327 204
rect 325 203 326 204
rect 324 203 325 204
rect 323 203 324 204
rect 322 203 323 204
rect 321 203 322 204
rect 320 203 321 204
rect 319 203 320 204
rect 318 203 319 204
rect 317 203 318 204
rect 316 203 317 204
rect 315 203 316 204
rect 314 203 315 204
rect 313 203 314 204
rect 312 203 313 204
rect 311 203 312 204
rect 310 203 311 204
rect 309 203 310 204
rect 308 203 309 204
rect 307 203 308 204
rect 306 203 307 204
rect 305 203 306 204
rect 304 203 305 204
rect 303 203 304 204
rect 302 203 303 204
rect 301 203 302 204
rect 300 203 301 204
rect 299 203 300 204
rect 298 203 299 204
rect 297 203 298 204
rect 296 203 297 204
rect 295 203 296 204
rect 294 203 295 204
rect 293 203 294 204
rect 292 203 293 204
rect 291 203 292 204
rect 290 203 291 204
rect 289 203 290 204
rect 288 203 289 204
rect 287 203 288 204
rect 286 203 287 204
rect 285 203 286 204
rect 284 203 285 204
rect 283 203 284 204
rect 282 203 283 204
rect 281 203 282 204
rect 280 203 281 204
rect 279 203 280 204
rect 278 203 279 204
rect 277 203 278 204
rect 276 203 277 204
rect 275 203 276 204
rect 274 203 275 204
rect 273 203 274 204
rect 272 203 273 204
rect 271 203 272 204
rect 270 203 271 204
rect 269 203 270 204
rect 268 203 269 204
rect 267 203 268 204
rect 266 203 267 204
rect 265 203 266 204
rect 264 203 265 204
rect 263 203 264 204
rect 262 203 263 204
rect 251 203 252 204
rect 250 203 251 204
rect 249 203 250 204
rect 248 203 249 204
rect 247 203 248 204
rect 246 203 247 204
rect 245 203 246 204
rect 244 203 245 204
rect 243 203 244 204
rect 242 203 243 204
rect 241 203 242 204
rect 240 203 241 204
rect 239 203 240 204
rect 238 203 239 204
rect 237 203 238 204
rect 236 203 237 204
rect 235 203 236 204
rect 234 203 235 204
rect 233 203 234 204
rect 232 203 233 204
rect 231 203 232 204
rect 230 203 231 204
rect 229 203 230 204
rect 228 203 229 204
rect 227 203 228 204
rect 226 203 227 204
rect 225 203 226 204
rect 224 203 225 204
rect 223 203 224 204
rect 222 203 223 204
rect 221 203 222 204
rect 220 203 221 204
rect 219 203 220 204
rect 218 203 219 204
rect 217 203 218 204
rect 216 203 217 204
rect 215 203 216 204
rect 214 203 215 204
rect 213 203 214 204
rect 212 203 213 204
rect 211 203 212 204
rect 210 203 211 204
rect 182 203 183 204
rect 181 203 182 204
rect 180 203 181 204
rect 179 203 180 204
rect 178 203 179 204
rect 177 203 178 204
rect 176 203 177 204
rect 175 203 176 204
rect 174 203 175 204
rect 173 203 174 204
rect 172 203 173 204
rect 171 203 172 204
rect 170 203 171 204
rect 169 203 170 204
rect 168 203 169 204
rect 167 203 168 204
rect 166 203 167 204
rect 165 203 166 204
rect 164 203 165 204
rect 163 203 164 204
rect 162 203 163 204
rect 161 203 162 204
rect 160 203 161 204
rect 159 203 160 204
rect 158 203 159 204
rect 157 203 158 204
rect 156 203 157 204
rect 155 203 156 204
rect 154 203 155 204
rect 153 203 154 204
rect 152 203 153 204
rect 151 203 152 204
rect 150 203 151 204
rect 149 203 150 204
rect 148 203 149 204
rect 147 203 148 204
rect 146 203 147 204
rect 145 203 146 204
rect 144 203 145 204
rect 143 203 144 204
rect 142 203 143 204
rect 141 203 142 204
rect 140 203 141 204
rect 139 203 140 204
rect 138 203 139 204
rect 137 203 138 204
rect 136 203 137 204
rect 135 203 136 204
rect 134 203 135 204
rect 133 203 134 204
rect 132 203 133 204
rect 131 203 132 204
rect 130 203 131 204
rect 129 203 130 204
rect 128 203 129 204
rect 127 203 128 204
rect 126 203 127 204
rect 125 203 126 204
rect 124 203 125 204
rect 123 203 124 204
rect 122 203 123 204
rect 121 203 122 204
rect 120 203 121 204
rect 119 203 120 204
rect 118 203 119 204
rect 117 203 118 204
rect 116 203 117 204
rect 115 203 116 204
rect 114 203 115 204
rect 113 203 114 204
rect 112 203 113 204
rect 111 203 112 204
rect 110 203 111 204
rect 109 203 110 204
rect 108 203 109 204
rect 107 203 108 204
rect 106 203 107 204
rect 105 203 106 204
rect 104 203 105 204
rect 103 203 104 204
rect 102 203 103 204
rect 101 203 102 204
rect 100 203 101 204
rect 99 203 100 204
rect 98 203 99 204
rect 97 203 98 204
rect 96 203 97 204
rect 95 203 96 204
rect 94 203 95 204
rect 93 203 94 204
rect 92 203 93 204
rect 91 203 92 204
rect 90 203 91 204
rect 89 203 90 204
rect 88 203 89 204
rect 87 203 88 204
rect 86 203 87 204
rect 85 203 86 204
rect 84 203 85 204
rect 83 203 84 204
rect 82 203 83 204
rect 81 203 82 204
rect 80 203 81 204
rect 79 203 80 204
rect 78 203 79 204
rect 77 203 78 204
rect 76 203 77 204
rect 75 203 76 204
rect 74 203 75 204
rect 57 203 58 204
rect 56 203 57 204
rect 55 203 56 204
rect 54 203 55 204
rect 53 203 54 204
rect 52 203 53 204
rect 51 203 52 204
rect 50 203 51 204
rect 49 203 50 204
rect 48 203 49 204
rect 47 203 48 204
rect 46 203 47 204
rect 45 203 46 204
rect 44 203 45 204
rect 43 203 44 204
rect 42 203 43 204
rect 41 203 42 204
rect 40 203 41 204
rect 39 203 40 204
rect 38 203 39 204
rect 37 203 38 204
rect 36 203 37 204
rect 35 203 36 204
rect 34 203 35 204
rect 33 203 34 204
rect 32 203 33 204
rect 31 203 32 204
rect 30 203 31 204
rect 29 203 30 204
rect 28 203 29 204
rect 27 203 28 204
rect 26 203 27 204
rect 25 203 26 204
rect 24 203 25 204
rect 23 203 24 204
rect 22 203 23 204
rect 21 203 22 204
rect 20 203 21 204
rect 19 203 20 204
rect 18 203 19 204
rect 17 203 18 204
rect 16 203 17 204
rect 15 203 16 204
rect 14 203 15 204
rect 13 203 14 204
rect 482 204 483 205
rect 472 204 473 205
rect 471 204 472 205
rect 462 204 463 205
rect 399 204 400 205
rect 398 204 399 205
rect 397 204 398 205
rect 352 204 353 205
rect 351 204 352 205
rect 350 204 351 205
rect 349 204 350 205
rect 348 204 349 205
rect 347 204 348 205
rect 346 204 347 205
rect 345 204 346 205
rect 344 204 345 205
rect 343 204 344 205
rect 342 204 343 205
rect 341 204 342 205
rect 340 204 341 205
rect 339 204 340 205
rect 338 204 339 205
rect 337 204 338 205
rect 336 204 337 205
rect 335 204 336 205
rect 334 204 335 205
rect 333 204 334 205
rect 332 204 333 205
rect 331 204 332 205
rect 330 204 331 205
rect 329 204 330 205
rect 328 204 329 205
rect 327 204 328 205
rect 326 204 327 205
rect 325 204 326 205
rect 324 204 325 205
rect 323 204 324 205
rect 322 204 323 205
rect 321 204 322 205
rect 320 204 321 205
rect 319 204 320 205
rect 318 204 319 205
rect 317 204 318 205
rect 316 204 317 205
rect 315 204 316 205
rect 314 204 315 205
rect 313 204 314 205
rect 312 204 313 205
rect 311 204 312 205
rect 310 204 311 205
rect 309 204 310 205
rect 308 204 309 205
rect 307 204 308 205
rect 306 204 307 205
rect 305 204 306 205
rect 304 204 305 205
rect 303 204 304 205
rect 302 204 303 205
rect 301 204 302 205
rect 300 204 301 205
rect 299 204 300 205
rect 298 204 299 205
rect 297 204 298 205
rect 296 204 297 205
rect 295 204 296 205
rect 294 204 295 205
rect 293 204 294 205
rect 292 204 293 205
rect 291 204 292 205
rect 290 204 291 205
rect 289 204 290 205
rect 288 204 289 205
rect 287 204 288 205
rect 286 204 287 205
rect 285 204 286 205
rect 284 204 285 205
rect 283 204 284 205
rect 282 204 283 205
rect 281 204 282 205
rect 280 204 281 205
rect 279 204 280 205
rect 278 204 279 205
rect 277 204 278 205
rect 276 204 277 205
rect 275 204 276 205
rect 274 204 275 205
rect 273 204 274 205
rect 272 204 273 205
rect 271 204 272 205
rect 270 204 271 205
rect 269 204 270 205
rect 268 204 269 205
rect 267 204 268 205
rect 266 204 267 205
rect 265 204 266 205
rect 264 204 265 205
rect 263 204 264 205
rect 262 204 263 205
rect 261 204 262 205
rect 260 204 261 205
rect 251 204 252 205
rect 250 204 251 205
rect 249 204 250 205
rect 248 204 249 205
rect 247 204 248 205
rect 246 204 247 205
rect 245 204 246 205
rect 244 204 245 205
rect 243 204 244 205
rect 242 204 243 205
rect 241 204 242 205
rect 240 204 241 205
rect 239 204 240 205
rect 238 204 239 205
rect 237 204 238 205
rect 236 204 237 205
rect 235 204 236 205
rect 234 204 235 205
rect 233 204 234 205
rect 232 204 233 205
rect 231 204 232 205
rect 230 204 231 205
rect 229 204 230 205
rect 228 204 229 205
rect 227 204 228 205
rect 226 204 227 205
rect 225 204 226 205
rect 224 204 225 205
rect 223 204 224 205
rect 222 204 223 205
rect 221 204 222 205
rect 220 204 221 205
rect 219 204 220 205
rect 218 204 219 205
rect 217 204 218 205
rect 216 204 217 205
rect 215 204 216 205
rect 214 204 215 205
rect 213 204 214 205
rect 212 204 213 205
rect 211 204 212 205
rect 210 204 211 205
rect 209 204 210 205
rect 181 204 182 205
rect 180 204 181 205
rect 179 204 180 205
rect 178 204 179 205
rect 177 204 178 205
rect 176 204 177 205
rect 175 204 176 205
rect 174 204 175 205
rect 173 204 174 205
rect 172 204 173 205
rect 171 204 172 205
rect 170 204 171 205
rect 169 204 170 205
rect 168 204 169 205
rect 167 204 168 205
rect 166 204 167 205
rect 165 204 166 205
rect 164 204 165 205
rect 163 204 164 205
rect 162 204 163 205
rect 161 204 162 205
rect 160 204 161 205
rect 159 204 160 205
rect 158 204 159 205
rect 157 204 158 205
rect 156 204 157 205
rect 155 204 156 205
rect 154 204 155 205
rect 153 204 154 205
rect 152 204 153 205
rect 151 204 152 205
rect 150 204 151 205
rect 149 204 150 205
rect 148 204 149 205
rect 147 204 148 205
rect 146 204 147 205
rect 145 204 146 205
rect 144 204 145 205
rect 143 204 144 205
rect 142 204 143 205
rect 141 204 142 205
rect 140 204 141 205
rect 139 204 140 205
rect 138 204 139 205
rect 137 204 138 205
rect 136 204 137 205
rect 135 204 136 205
rect 134 204 135 205
rect 133 204 134 205
rect 132 204 133 205
rect 131 204 132 205
rect 130 204 131 205
rect 129 204 130 205
rect 128 204 129 205
rect 127 204 128 205
rect 126 204 127 205
rect 125 204 126 205
rect 124 204 125 205
rect 123 204 124 205
rect 122 204 123 205
rect 121 204 122 205
rect 120 204 121 205
rect 119 204 120 205
rect 118 204 119 205
rect 117 204 118 205
rect 116 204 117 205
rect 115 204 116 205
rect 114 204 115 205
rect 113 204 114 205
rect 112 204 113 205
rect 111 204 112 205
rect 110 204 111 205
rect 109 204 110 205
rect 108 204 109 205
rect 107 204 108 205
rect 106 204 107 205
rect 105 204 106 205
rect 104 204 105 205
rect 103 204 104 205
rect 102 204 103 205
rect 101 204 102 205
rect 100 204 101 205
rect 99 204 100 205
rect 98 204 99 205
rect 97 204 98 205
rect 96 204 97 205
rect 95 204 96 205
rect 94 204 95 205
rect 93 204 94 205
rect 92 204 93 205
rect 91 204 92 205
rect 90 204 91 205
rect 89 204 90 205
rect 88 204 89 205
rect 87 204 88 205
rect 86 204 87 205
rect 85 204 86 205
rect 84 204 85 205
rect 83 204 84 205
rect 82 204 83 205
rect 81 204 82 205
rect 80 204 81 205
rect 79 204 80 205
rect 78 204 79 205
rect 77 204 78 205
rect 76 204 77 205
rect 75 204 76 205
rect 58 204 59 205
rect 57 204 58 205
rect 56 204 57 205
rect 55 204 56 205
rect 54 204 55 205
rect 53 204 54 205
rect 52 204 53 205
rect 51 204 52 205
rect 50 204 51 205
rect 49 204 50 205
rect 48 204 49 205
rect 47 204 48 205
rect 46 204 47 205
rect 45 204 46 205
rect 44 204 45 205
rect 43 204 44 205
rect 42 204 43 205
rect 41 204 42 205
rect 40 204 41 205
rect 39 204 40 205
rect 38 204 39 205
rect 37 204 38 205
rect 36 204 37 205
rect 35 204 36 205
rect 34 204 35 205
rect 33 204 34 205
rect 32 204 33 205
rect 31 204 32 205
rect 30 204 31 205
rect 29 204 30 205
rect 28 204 29 205
rect 27 204 28 205
rect 26 204 27 205
rect 25 204 26 205
rect 24 204 25 205
rect 23 204 24 205
rect 22 204 23 205
rect 21 204 22 205
rect 20 204 21 205
rect 19 204 20 205
rect 18 204 19 205
rect 17 204 18 205
rect 16 204 17 205
rect 15 204 16 205
rect 14 204 15 205
rect 13 204 14 205
rect 482 205 483 206
rect 474 205 475 206
rect 473 205 474 206
rect 472 205 473 206
rect 471 205 472 206
rect 470 205 471 206
rect 469 205 470 206
rect 463 205 464 206
rect 462 205 463 206
rect 398 205 399 206
rect 353 205 354 206
rect 352 205 353 206
rect 351 205 352 206
rect 350 205 351 206
rect 349 205 350 206
rect 348 205 349 206
rect 347 205 348 206
rect 346 205 347 206
rect 345 205 346 206
rect 344 205 345 206
rect 343 205 344 206
rect 342 205 343 206
rect 341 205 342 206
rect 340 205 341 206
rect 339 205 340 206
rect 338 205 339 206
rect 337 205 338 206
rect 336 205 337 206
rect 335 205 336 206
rect 334 205 335 206
rect 333 205 334 206
rect 332 205 333 206
rect 331 205 332 206
rect 330 205 331 206
rect 329 205 330 206
rect 328 205 329 206
rect 327 205 328 206
rect 326 205 327 206
rect 325 205 326 206
rect 324 205 325 206
rect 323 205 324 206
rect 322 205 323 206
rect 321 205 322 206
rect 320 205 321 206
rect 319 205 320 206
rect 318 205 319 206
rect 317 205 318 206
rect 316 205 317 206
rect 315 205 316 206
rect 314 205 315 206
rect 313 205 314 206
rect 312 205 313 206
rect 311 205 312 206
rect 310 205 311 206
rect 309 205 310 206
rect 308 205 309 206
rect 307 205 308 206
rect 306 205 307 206
rect 305 205 306 206
rect 304 205 305 206
rect 303 205 304 206
rect 302 205 303 206
rect 301 205 302 206
rect 300 205 301 206
rect 299 205 300 206
rect 298 205 299 206
rect 297 205 298 206
rect 296 205 297 206
rect 295 205 296 206
rect 294 205 295 206
rect 293 205 294 206
rect 292 205 293 206
rect 291 205 292 206
rect 290 205 291 206
rect 289 205 290 206
rect 288 205 289 206
rect 287 205 288 206
rect 286 205 287 206
rect 285 205 286 206
rect 284 205 285 206
rect 283 205 284 206
rect 282 205 283 206
rect 281 205 282 206
rect 280 205 281 206
rect 279 205 280 206
rect 278 205 279 206
rect 277 205 278 206
rect 276 205 277 206
rect 275 205 276 206
rect 274 205 275 206
rect 273 205 274 206
rect 272 205 273 206
rect 271 205 272 206
rect 270 205 271 206
rect 269 205 270 206
rect 268 205 269 206
rect 267 205 268 206
rect 266 205 267 206
rect 265 205 266 206
rect 264 205 265 206
rect 263 205 264 206
rect 262 205 263 206
rect 261 205 262 206
rect 260 205 261 206
rect 259 205 260 206
rect 250 205 251 206
rect 249 205 250 206
rect 248 205 249 206
rect 247 205 248 206
rect 246 205 247 206
rect 245 205 246 206
rect 244 205 245 206
rect 243 205 244 206
rect 242 205 243 206
rect 241 205 242 206
rect 240 205 241 206
rect 239 205 240 206
rect 238 205 239 206
rect 237 205 238 206
rect 236 205 237 206
rect 235 205 236 206
rect 234 205 235 206
rect 233 205 234 206
rect 232 205 233 206
rect 231 205 232 206
rect 230 205 231 206
rect 229 205 230 206
rect 228 205 229 206
rect 227 205 228 206
rect 226 205 227 206
rect 225 205 226 206
rect 224 205 225 206
rect 223 205 224 206
rect 222 205 223 206
rect 221 205 222 206
rect 220 205 221 206
rect 219 205 220 206
rect 218 205 219 206
rect 217 205 218 206
rect 216 205 217 206
rect 215 205 216 206
rect 214 205 215 206
rect 213 205 214 206
rect 212 205 213 206
rect 211 205 212 206
rect 210 205 211 206
rect 209 205 210 206
rect 208 205 209 206
rect 179 205 180 206
rect 178 205 179 206
rect 177 205 178 206
rect 176 205 177 206
rect 175 205 176 206
rect 174 205 175 206
rect 173 205 174 206
rect 172 205 173 206
rect 171 205 172 206
rect 170 205 171 206
rect 169 205 170 206
rect 168 205 169 206
rect 167 205 168 206
rect 166 205 167 206
rect 165 205 166 206
rect 164 205 165 206
rect 163 205 164 206
rect 162 205 163 206
rect 161 205 162 206
rect 160 205 161 206
rect 159 205 160 206
rect 158 205 159 206
rect 157 205 158 206
rect 156 205 157 206
rect 155 205 156 206
rect 154 205 155 206
rect 153 205 154 206
rect 152 205 153 206
rect 151 205 152 206
rect 150 205 151 206
rect 149 205 150 206
rect 148 205 149 206
rect 147 205 148 206
rect 146 205 147 206
rect 145 205 146 206
rect 144 205 145 206
rect 143 205 144 206
rect 142 205 143 206
rect 141 205 142 206
rect 140 205 141 206
rect 139 205 140 206
rect 138 205 139 206
rect 137 205 138 206
rect 136 205 137 206
rect 135 205 136 206
rect 134 205 135 206
rect 133 205 134 206
rect 132 205 133 206
rect 131 205 132 206
rect 130 205 131 206
rect 129 205 130 206
rect 128 205 129 206
rect 127 205 128 206
rect 126 205 127 206
rect 125 205 126 206
rect 124 205 125 206
rect 123 205 124 206
rect 122 205 123 206
rect 121 205 122 206
rect 120 205 121 206
rect 119 205 120 206
rect 118 205 119 206
rect 117 205 118 206
rect 116 205 117 206
rect 115 205 116 206
rect 114 205 115 206
rect 113 205 114 206
rect 112 205 113 206
rect 111 205 112 206
rect 110 205 111 206
rect 109 205 110 206
rect 108 205 109 206
rect 107 205 108 206
rect 106 205 107 206
rect 105 205 106 206
rect 104 205 105 206
rect 103 205 104 206
rect 102 205 103 206
rect 101 205 102 206
rect 100 205 101 206
rect 99 205 100 206
rect 98 205 99 206
rect 97 205 98 206
rect 96 205 97 206
rect 95 205 96 206
rect 94 205 95 206
rect 93 205 94 206
rect 92 205 93 206
rect 91 205 92 206
rect 90 205 91 206
rect 89 205 90 206
rect 88 205 89 206
rect 87 205 88 206
rect 86 205 87 206
rect 85 205 86 206
rect 84 205 85 206
rect 83 205 84 206
rect 82 205 83 206
rect 81 205 82 206
rect 80 205 81 206
rect 79 205 80 206
rect 78 205 79 206
rect 77 205 78 206
rect 76 205 77 206
rect 75 205 76 206
rect 58 205 59 206
rect 57 205 58 206
rect 56 205 57 206
rect 55 205 56 206
rect 54 205 55 206
rect 53 205 54 206
rect 52 205 53 206
rect 51 205 52 206
rect 50 205 51 206
rect 49 205 50 206
rect 48 205 49 206
rect 47 205 48 206
rect 46 205 47 206
rect 45 205 46 206
rect 44 205 45 206
rect 43 205 44 206
rect 42 205 43 206
rect 41 205 42 206
rect 40 205 41 206
rect 39 205 40 206
rect 38 205 39 206
rect 37 205 38 206
rect 36 205 37 206
rect 35 205 36 206
rect 34 205 35 206
rect 33 205 34 206
rect 32 205 33 206
rect 31 205 32 206
rect 30 205 31 206
rect 29 205 30 206
rect 28 205 29 206
rect 27 205 28 206
rect 26 205 27 206
rect 25 205 26 206
rect 24 205 25 206
rect 23 205 24 206
rect 22 205 23 206
rect 21 205 22 206
rect 20 205 21 206
rect 19 205 20 206
rect 18 205 19 206
rect 17 205 18 206
rect 16 205 17 206
rect 15 205 16 206
rect 14 205 15 206
rect 13 205 14 206
rect 482 206 483 207
rect 481 206 482 207
rect 475 206 476 207
rect 474 206 475 207
rect 473 206 474 207
rect 472 206 473 207
rect 471 206 472 207
rect 470 206 471 207
rect 469 206 470 207
rect 464 206 465 207
rect 463 206 464 207
rect 462 206 463 207
rect 354 206 355 207
rect 353 206 354 207
rect 352 206 353 207
rect 351 206 352 207
rect 350 206 351 207
rect 349 206 350 207
rect 348 206 349 207
rect 347 206 348 207
rect 346 206 347 207
rect 345 206 346 207
rect 344 206 345 207
rect 343 206 344 207
rect 342 206 343 207
rect 341 206 342 207
rect 340 206 341 207
rect 339 206 340 207
rect 338 206 339 207
rect 337 206 338 207
rect 336 206 337 207
rect 335 206 336 207
rect 334 206 335 207
rect 333 206 334 207
rect 332 206 333 207
rect 331 206 332 207
rect 330 206 331 207
rect 329 206 330 207
rect 328 206 329 207
rect 327 206 328 207
rect 326 206 327 207
rect 325 206 326 207
rect 324 206 325 207
rect 323 206 324 207
rect 322 206 323 207
rect 321 206 322 207
rect 320 206 321 207
rect 319 206 320 207
rect 318 206 319 207
rect 317 206 318 207
rect 316 206 317 207
rect 315 206 316 207
rect 314 206 315 207
rect 313 206 314 207
rect 312 206 313 207
rect 311 206 312 207
rect 310 206 311 207
rect 309 206 310 207
rect 308 206 309 207
rect 307 206 308 207
rect 306 206 307 207
rect 305 206 306 207
rect 304 206 305 207
rect 303 206 304 207
rect 302 206 303 207
rect 301 206 302 207
rect 300 206 301 207
rect 299 206 300 207
rect 298 206 299 207
rect 297 206 298 207
rect 296 206 297 207
rect 295 206 296 207
rect 294 206 295 207
rect 293 206 294 207
rect 292 206 293 207
rect 291 206 292 207
rect 290 206 291 207
rect 289 206 290 207
rect 288 206 289 207
rect 287 206 288 207
rect 286 206 287 207
rect 285 206 286 207
rect 284 206 285 207
rect 283 206 284 207
rect 282 206 283 207
rect 281 206 282 207
rect 280 206 281 207
rect 279 206 280 207
rect 278 206 279 207
rect 277 206 278 207
rect 276 206 277 207
rect 275 206 276 207
rect 274 206 275 207
rect 273 206 274 207
rect 272 206 273 207
rect 271 206 272 207
rect 270 206 271 207
rect 269 206 270 207
rect 268 206 269 207
rect 267 206 268 207
rect 266 206 267 207
rect 265 206 266 207
rect 264 206 265 207
rect 263 206 264 207
rect 262 206 263 207
rect 261 206 262 207
rect 260 206 261 207
rect 259 206 260 207
rect 258 206 259 207
rect 257 206 258 207
rect 249 206 250 207
rect 248 206 249 207
rect 247 206 248 207
rect 246 206 247 207
rect 245 206 246 207
rect 244 206 245 207
rect 243 206 244 207
rect 242 206 243 207
rect 241 206 242 207
rect 240 206 241 207
rect 239 206 240 207
rect 238 206 239 207
rect 237 206 238 207
rect 236 206 237 207
rect 235 206 236 207
rect 234 206 235 207
rect 233 206 234 207
rect 232 206 233 207
rect 231 206 232 207
rect 230 206 231 207
rect 229 206 230 207
rect 228 206 229 207
rect 227 206 228 207
rect 226 206 227 207
rect 225 206 226 207
rect 224 206 225 207
rect 223 206 224 207
rect 222 206 223 207
rect 221 206 222 207
rect 220 206 221 207
rect 219 206 220 207
rect 218 206 219 207
rect 217 206 218 207
rect 216 206 217 207
rect 215 206 216 207
rect 214 206 215 207
rect 213 206 214 207
rect 212 206 213 207
rect 211 206 212 207
rect 210 206 211 207
rect 209 206 210 207
rect 208 206 209 207
rect 207 206 208 207
rect 177 206 178 207
rect 176 206 177 207
rect 175 206 176 207
rect 174 206 175 207
rect 173 206 174 207
rect 172 206 173 207
rect 171 206 172 207
rect 170 206 171 207
rect 169 206 170 207
rect 168 206 169 207
rect 167 206 168 207
rect 166 206 167 207
rect 165 206 166 207
rect 164 206 165 207
rect 163 206 164 207
rect 162 206 163 207
rect 161 206 162 207
rect 160 206 161 207
rect 159 206 160 207
rect 158 206 159 207
rect 157 206 158 207
rect 156 206 157 207
rect 155 206 156 207
rect 154 206 155 207
rect 153 206 154 207
rect 152 206 153 207
rect 151 206 152 207
rect 150 206 151 207
rect 149 206 150 207
rect 148 206 149 207
rect 147 206 148 207
rect 146 206 147 207
rect 145 206 146 207
rect 144 206 145 207
rect 143 206 144 207
rect 142 206 143 207
rect 141 206 142 207
rect 140 206 141 207
rect 139 206 140 207
rect 138 206 139 207
rect 137 206 138 207
rect 136 206 137 207
rect 135 206 136 207
rect 134 206 135 207
rect 133 206 134 207
rect 132 206 133 207
rect 131 206 132 207
rect 130 206 131 207
rect 129 206 130 207
rect 128 206 129 207
rect 127 206 128 207
rect 126 206 127 207
rect 125 206 126 207
rect 124 206 125 207
rect 123 206 124 207
rect 122 206 123 207
rect 121 206 122 207
rect 120 206 121 207
rect 119 206 120 207
rect 118 206 119 207
rect 117 206 118 207
rect 116 206 117 207
rect 115 206 116 207
rect 114 206 115 207
rect 113 206 114 207
rect 112 206 113 207
rect 111 206 112 207
rect 110 206 111 207
rect 109 206 110 207
rect 108 206 109 207
rect 107 206 108 207
rect 106 206 107 207
rect 105 206 106 207
rect 104 206 105 207
rect 103 206 104 207
rect 102 206 103 207
rect 101 206 102 207
rect 100 206 101 207
rect 99 206 100 207
rect 98 206 99 207
rect 97 206 98 207
rect 96 206 97 207
rect 95 206 96 207
rect 94 206 95 207
rect 93 206 94 207
rect 92 206 93 207
rect 91 206 92 207
rect 90 206 91 207
rect 89 206 90 207
rect 88 206 89 207
rect 87 206 88 207
rect 86 206 87 207
rect 85 206 86 207
rect 84 206 85 207
rect 83 206 84 207
rect 82 206 83 207
rect 81 206 82 207
rect 80 206 81 207
rect 79 206 80 207
rect 78 206 79 207
rect 77 206 78 207
rect 76 206 77 207
rect 59 206 60 207
rect 58 206 59 207
rect 57 206 58 207
rect 56 206 57 207
rect 55 206 56 207
rect 54 206 55 207
rect 53 206 54 207
rect 52 206 53 207
rect 51 206 52 207
rect 50 206 51 207
rect 49 206 50 207
rect 48 206 49 207
rect 47 206 48 207
rect 46 206 47 207
rect 45 206 46 207
rect 44 206 45 207
rect 43 206 44 207
rect 42 206 43 207
rect 41 206 42 207
rect 40 206 41 207
rect 39 206 40 207
rect 38 206 39 207
rect 37 206 38 207
rect 36 206 37 207
rect 35 206 36 207
rect 34 206 35 207
rect 33 206 34 207
rect 32 206 33 207
rect 31 206 32 207
rect 30 206 31 207
rect 29 206 30 207
rect 28 206 29 207
rect 27 206 28 207
rect 26 206 27 207
rect 25 206 26 207
rect 24 206 25 207
rect 23 206 24 207
rect 22 206 23 207
rect 21 206 22 207
rect 20 206 21 207
rect 19 206 20 207
rect 18 206 19 207
rect 17 206 18 207
rect 16 206 17 207
rect 15 206 16 207
rect 14 206 15 207
rect 13 206 14 207
rect 12 206 13 207
rect 482 207 483 208
rect 481 207 482 208
rect 480 207 481 208
rect 466 207 467 208
rect 465 207 466 208
rect 464 207 465 208
rect 463 207 464 208
rect 462 207 463 208
rect 355 207 356 208
rect 354 207 355 208
rect 353 207 354 208
rect 352 207 353 208
rect 351 207 352 208
rect 350 207 351 208
rect 349 207 350 208
rect 348 207 349 208
rect 347 207 348 208
rect 346 207 347 208
rect 345 207 346 208
rect 344 207 345 208
rect 343 207 344 208
rect 342 207 343 208
rect 341 207 342 208
rect 340 207 341 208
rect 339 207 340 208
rect 338 207 339 208
rect 337 207 338 208
rect 336 207 337 208
rect 335 207 336 208
rect 334 207 335 208
rect 333 207 334 208
rect 332 207 333 208
rect 331 207 332 208
rect 330 207 331 208
rect 329 207 330 208
rect 328 207 329 208
rect 327 207 328 208
rect 326 207 327 208
rect 325 207 326 208
rect 324 207 325 208
rect 323 207 324 208
rect 322 207 323 208
rect 321 207 322 208
rect 320 207 321 208
rect 319 207 320 208
rect 318 207 319 208
rect 317 207 318 208
rect 316 207 317 208
rect 315 207 316 208
rect 314 207 315 208
rect 313 207 314 208
rect 312 207 313 208
rect 311 207 312 208
rect 310 207 311 208
rect 309 207 310 208
rect 308 207 309 208
rect 307 207 308 208
rect 306 207 307 208
rect 305 207 306 208
rect 304 207 305 208
rect 303 207 304 208
rect 302 207 303 208
rect 301 207 302 208
rect 300 207 301 208
rect 299 207 300 208
rect 298 207 299 208
rect 297 207 298 208
rect 296 207 297 208
rect 295 207 296 208
rect 294 207 295 208
rect 293 207 294 208
rect 292 207 293 208
rect 291 207 292 208
rect 290 207 291 208
rect 289 207 290 208
rect 288 207 289 208
rect 287 207 288 208
rect 286 207 287 208
rect 285 207 286 208
rect 284 207 285 208
rect 283 207 284 208
rect 282 207 283 208
rect 281 207 282 208
rect 280 207 281 208
rect 279 207 280 208
rect 278 207 279 208
rect 277 207 278 208
rect 276 207 277 208
rect 275 207 276 208
rect 274 207 275 208
rect 273 207 274 208
rect 272 207 273 208
rect 271 207 272 208
rect 270 207 271 208
rect 269 207 270 208
rect 268 207 269 208
rect 267 207 268 208
rect 266 207 267 208
rect 265 207 266 208
rect 264 207 265 208
rect 263 207 264 208
rect 262 207 263 208
rect 261 207 262 208
rect 260 207 261 208
rect 259 207 260 208
rect 258 207 259 208
rect 257 207 258 208
rect 256 207 257 208
rect 255 207 256 208
rect 249 207 250 208
rect 248 207 249 208
rect 247 207 248 208
rect 246 207 247 208
rect 245 207 246 208
rect 244 207 245 208
rect 243 207 244 208
rect 242 207 243 208
rect 241 207 242 208
rect 240 207 241 208
rect 239 207 240 208
rect 238 207 239 208
rect 237 207 238 208
rect 236 207 237 208
rect 235 207 236 208
rect 234 207 235 208
rect 233 207 234 208
rect 232 207 233 208
rect 231 207 232 208
rect 230 207 231 208
rect 229 207 230 208
rect 228 207 229 208
rect 227 207 228 208
rect 226 207 227 208
rect 225 207 226 208
rect 224 207 225 208
rect 223 207 224 208
rect 222 207 223 208
rect 221 207 222 208
rect 220 207 221 208
rect 219 207 220 208
rect 218 207 219 208
rect 217 207 218 208
rect 216 207 217 208
rect 215 207 216 208
rect 214 207 215 208
rect 213 207 214 208
rect 212 207 213 208
rect 211 207 212 208
rect 210 207 211 208
rect 209 207 210 208
rect 208 207 209 208
rect 207 207 208 208
rect 206 207 207 208
rect 175 207 176 208
rect 174 207 175 208
rect 173 207 174 208
rect 172 207 173 208
rect 171 207 172 208
rect 170 207 171 208
rect 169 207 170 208
rect 168 207 169 208
rect 167 207 168 208
rect 166 207 167 208
rect 165 207 166 208
rect 164 207 165 208
rect 163 207 164 208
rect 162 207 163 208
rect 161 207 162 208
rect 160 207 161 208
rect 159 207 160 208
rect 158 207 159 208
rect 157 207 158 208
rect 156 207 157 208
rect 155 207 156 208
rect 154 207 155 208
rect 153 207 154 208
rect 152 207 153 208
rect 151 207 152 208
rect 150 207 151 208
rect 149 207 150 208
rect 148 207 149 208
rect 147 207 148 208
rect 146 207 147 208
rect 145 207 146 208
rect 144 207 145 208
rect 143 207 144 208
rect 142 207 143 208
rect 141 207 142 208
rect 140 207 141 208
rect 139 207 140 208
rect 138 207 139 208
rect 137 207 138 208
rect 136 207 137 208
rect 135 207 136 208
rect 134 207 135 208
rect 133 207 134 208
rect 132 207 133 208
rect 131 207 132 208
rect 130 207 131 208
rect 129 207 130 208
rect 128 207 129 208
rect 127 207 128 208
rect 126 207 127 208
rect 125 207 126 208
rect 124 207 125 208
rect 123 207 124 208
rect 122 207 123 208
rect 121 207 122 208
rect 120 207 121 208
rect 119 207 120 208
rect 118 207 119 208
rect 117 207 118 208
rect 116 207 117 208
rect 115 207 116 208
rect 114 207 115 208
rect 113 207 114 208
rect 112 207 113 208
rect 111 207 112 208
rect 110 207 111 208
rect 109 207 110 208
rect 108 207 109 208
rect 107 207 108 208
rect 106 207 107 208
rect 105 207 106 208
rect 104 207 105 208
rect 103 207 104 208
rect 102 207 103 208
rect 101 207 102 208
rect 100 207 101 208
rect 99 207 100 208
rect 98 207 99 208
rect 97 207 98 208
rect 96 207 97 208
rect 95 207 96 208
rect 94 207 95 208
rect 93 207 94 208
rect 92 207 93 208
rect 91 207 92 208
rect 90 207 91 208
rect 89 207 90 208
rect 88 207 89 208
rect 87 207 88 208
rect 86 207 87 208
rect 85 207 86 208
rect 84 207 85 208
rect 83 207 84 208
rect 82 207 83 208
rect 81 207 82 208
rect 80 207 81 208
rect 79 207 80 208
rect 78 207 79 208
rect 77 207 78 208
rect 60 207 61 208
rect 59 207 60 208
rect 58 207 59 208
rect 57 207 58 208
rect 56 207 57 208
rect 55 207 56 208
rect 54 207 55 208
rect 53 207 54 208
rect 52 207 53 208
rect 51 207 52 208
rect 50 207 51 208
rect 49 207 50 208
rect 48 207 49 208
rect 47 207 48 208
rect 46 207 47 208
rect 45 207 46 208
rect 44 207 45 208
rect 43 207 44 208
rect 42 207 43 208
rect 41 207 42 208
rect 40 207 41 208
rect 39 207 40 208
rect 38 207 39 208
rect 37 207 38 208
rect 36 207 37 208
rect 35 207 36 208
rect 34 207 35 208
rect 33 207 34 208
rect 32 207 33 208
rect 31 207 32 208
rect 30 207 31 208
rect 29 207 30 208
rect 28 207 29 208
rect 27 207 28 208
rect 26 207 27 208
rect 25 207 26 208
rect 24 207 25 208
rect 23 207 24 208
rect 22 207 23 208
rect 21 207 22 208
rect 20 207 21 208
rect 19 207 20 208
rect 18 207 19 208
rect 17 207 18 208
rect 16 207 17 208
rect 15 207 16 208
rect 14 207 15 208
rect 13 207 14 208
rect 12 207 13 208
rect 482 208 483 209
rect 481 208 482 209
rect 480 208 481 209
rect 479 208 480 209
rect 478 208 479 209
rect 466 208 467 209
rect 465 208 466 209
rect 464 208 465 209
rect 355 208 356 209
rect 354 208 355 209
rect 353 208 354 209
rect 352 208 353 209
rect 351 208 352 209
rect 350 208 351 209
rect 349 208 350 209
rect 348 208 349 209
rect 347 208 348 209
rect 346 208 347 209
rect 345 208 346 209
rect 344 208 345 209
rect 343 208 344 209
rect 342 208 343 209
rect 341 208 342 209
rect 340 208 341 209
rect 339 208 340 209
rect 338 208 339 209
rect 337 208 338 209
rect 336 208 337 209
rect 335 208 336 209
rect 334 208 335 209
rect 333 208 334 209
rect 332 208 333 209
rect 331 208 332 209
rect 330 208 331 209
rect 329 208 330 209
rect 328 208 329 209
rect 327 208 328 209
rect 326 208 327 209
rect 325 208 326 209
rect 324 208 325 209
rect 323 208 324 209
rect 322 208 323 209
rect 321 208 322 209
rect 320 208 321 209
rect 319 208 320 209
rect 318 208 319 209
rect 317 208 318 209
rect 316 208 317 209
rect 315 208 316 209
rect 314 208 315 209
rect 313 208 314 209
rect 312 208 313 209
rect 311 208 312 209
rect 310 208 311 209
rect 309 208 310 209
rect 308 208 309 209
rect 307 208 308 209
rect 306 208 307 209
rect 305 208 306 209
rect 304 208 305 209
rect 303 208 304 209
rect 302 208 303 209
rect 301 208 302 209
rect 300 208 301 209
rect 299 208 300 209
rect 298 208 299 209
rect 297 208 298 209
rect 296 208 297 209
rect 295 208 296 209
rect 294 208 295 209
rect 293 208 294 209
rect 292 208 293 209
rect 291 208 292 209
rect 290 208 291 209
rect 289 208 290 209
rect 288 208 289 209
rect 287 208 288 209
rect 286 208 287 209
rect 285 208 286 209
rect 284 208 285 209
rect 283 208 284 209
rect 282 208 283 209
rect 281 208 282 209
rect 280 208 281 209
rect 279 208 280 209
rect 278 208 279 209
rect 277 208 278 209
rect 276 208 277 209
rect 275 208 276 209
rect 274 208 275 209
rect 273 208 274 209
rect 272 208 273 209
rect 271 208 272 209
rect 270 208 271 209
rect 269 208 270 209
rect 268 208 269 209
rect 267 208 268 209
rect 266 208 267 209
rect 265 208 266 209
rect 264 208 265 209
rect 263 208 264 209
rect 262 208 263 209
rect 261 208 262 209
rect 260 208 261 209
rect 259 208 260 209
rect 258 208 259 209
rect 257 208 258 209
rect 256 208 257 209
rect 255 208 256 209
rect 254 208 255 209
rect 253 208 254 209
rect 248 208 249 209
rect 247 208 248 209
rect 246 208 247 209
rect 245 208 246 209
rect 244 208 245 209
rect 243 208 244 209
rect 242 208 243 209
rect 241 208 242 209
rect 240 208 241 209
rect 239 208 240 209
rect 238 208 239 209
rect 237 208 238 209
rect 236 208 237 209
rect 235 208 236 209
rect 234 208 235 209
rect 233 208 234 209
rect 232 208 233 209
rect 231 208 232 209
rect 230 208 231 209
rect 229 208 230 209
rect 228 208 229 209
rect 227 208 228 209
rect 226 208 227 209
rect 225 208 226 209
rect 224 208 225 209
rect 223 208 224 209
rect 222 208 223 209
rect 221 208 222 209
rect 220 208 221 209
rect 219 208 220 209
rect 218 208 219 209
rect 217 208 218 209
rect 216 208 217 209
rect 215 208 216 209
rect 214 208 215 209
rect 213 208 214 209
rect 212 208 213 209
rect 211 208 212 209
rect 210 208 211 209
rect 209 208 210 209
rect 208 208 209 209
rect 207 208 208 209
rect 206 208 207 209
rect 205 208 206 209
rect 173 208 174 209
rect 172 208 173 209
rect 171 208 172 209
rect 170 208 171 209
rect 169 208 170 209
rect 168 208 169 209
rect 167 208 168 209
rect 166 208 167 209
rect 165 208 166 209
rect 164 208 165 209
rect 163 208 164 209
rect 162 208 163 209
rect 161 208 162 209
rect 160 208 161 209
rect 159 208 160 209
rect 158 208 159 209
rect 157 208 158 209
rect 156 208 157 209
rect 155 208 156 209
rect 154 208 155 209
rect 153 208 154 209
rect 152 208 153 209
rect 151 208 152 209
rect 150 208 151 209
rect 149 208 150 209
rect 148 208 149 209
rect 147 208 148 209
rect 146 208 147 209
rect 145 208 146 209
rect 144 208 145 209
rect 143 208 144 209
rect 142 208 143 209
rect 141 208 142 209
rect 140 208 141 209
rect 139 208 140 209
rect 138 208 139 209
rect 137 208 138 209
rect 136 208 137 209
rect 135 208 136 209
rect 134 208 135 209
rect 133 208 134 209
rect 132 208 133 209
rect 131 208 132 209
rect 130 208 131 209
rect 129 208 130 209
rect 128 208 129 209
rect 127 208 128 209
rect 126 208 127 209
rect 125 208 126 209
rect 124 208 125 209
rect 123 208 124 209
rect 122 208 123 209
rect 121 208 122 209
rect 120 208 121 209
rect 119 208 120 209
rect 118 208 119 209
rect 117 208 118 209
rect 116 208 117 209
rect 115 208 116 209
rect 114 208 115 209
rect 113 208 114 209
rect 112 208 113 209
rect 111 208 112 209
rect 110 208 111 209
rect 109 208 110 209
rect 108 208 109 209
rect 107 208 108 209
rect 106 208 107 209
rect 105 208 106 209
rect 104 208 105 209
rect 103 208 104 209
rect 102 208 103 209
rect 101 208 102 209
rect 100 208 101 209
rect 99 208 100 209
rect 98 208 99 209
rect 97 208 98 209
rect 96 208 97 209
rect 95 208 96 209
rect 94 208 95 209
rect 93 208 94 209
rect 92 208 93 209
rect 91 208 92 209
rect 90 208 91 209
rect 89 208 90 209
rect 88 208 89 209
rect 87 208 88 209
rect 86 208 87 209
rect 85 208 86 209
rect 84 208 85 209
rect 83 208 84 209
rect 82 208 83 209
rect 81 208 82 209
rect 80 208 81 209
rect 79 208 80 209
rect 78 208 79 209
rect 60 208 61 209
rect 59 208 60 209
rect 58 208 59 209
rect 57 208 58 209
rect 56 208 57 209
rect 55 208 56 209
rect 54 208 55 209
rect 53 208 54 209
rect 52 208 53 209
rect 51 208 52 209
rect 50 208 51 209
rect 49 208 50 209
rect 48 208 49 209
rect 47 208 48 209
rect 46 208 47 209
rect 45 208 46 209
rect 44 208 45 209
rect 43 208 44 209
rect 42 208 43 209
rect 41 208 42 209
rect 40 208 41 209
rect 39 208 40 209
rect 38 208 39 209
rect 37 208 38 209
rect 36 208 37 209
rect 35 208 36 209
rect 34 208 35 209
rect 33 208 34 209
rect 32 208 33 209
rect 31 208 32 209
rect 30 208 31 209
rect 29 208 30 209
rect 28 208 29 209
rect 27 208 28 209
rect 26 208 27 209
rect 25 208 26 209
rect 24 208 25 209
rect 23 208 24 209
rect 22 208 23 209
rect 21 208 22 209
rect 20 208 21 209
rect 19 208 20 209
rect 18 208 19 209
rect 17 208 18 209
rect 16 208 17 209
rect 15 208 16 209
rect 14 208 15 209
rect 13 208 14 209
rect 12 208 13 209
rect 481 209 482 210
rect 480 209 481 210
rect 479 209 480 210
rect 478 209 479 210
rect 477 209 478 210
rect 424 209 425 210
rect 423 209 424 210
rect 422 209 423 210
rect 421 209 422 210
rect 420 209 421 210
rect 419 209 420 210
rect 418 209 419 210
rect 417 209 418 210
rect 416 209 417 210
rect 415 209 416 210
rect 356 209 357 210
rect 355 209 356 210
rect 354 209 355 210
rect 353 209 354 210
rect 352 209 353 210
rect 351 209 352 210
rect 350 209 351 210
rect 349 209 350 210
rect 348 209 349 210
rect 347 209 348 210
rect 346 209 347 210
rect 345 209 346 210
rect 344 209 345 210
rect 343 209 344 210
rect 342 209 343 210
rect 341 209 342 210
rect 340 209 341 210
rect 339 209 340 210
rect 338 209 339 210
rect 337 209 338 210
rect 336 209 337 210
rect 335 209 336 210
rect 334 209 335 210
rect 333 209 334 210
rect 332 209 333 210
rect 331 209 332 210
rect 330 209 331 210
rect 329 209 330 210
rect 328 209 329 210
rect 327 209 328 210
rect 326 209 327 210
rect 325 209 326 210
rect 324 209 325 210
rect 323 209 324 210
rect 322 209 323 210
rect 321 209 322 210
rect 320 209 321 210
rect 319 209 320 210
rect 318 209 319 210
rect 317 209 318 210
rect 316 209 317 210
rect 315 209 316 210
rect 314 209 315 210
rect 313 209 314 210
rect 312 209 313 210
rect 311 209 312 210
rect 310 209 311 210
rect 309 209 310 210
rect 308 209 309 210
rect 307 209 308 210
rect 306 209 307 210
rect 305 209 306 210
rect 304 209 305 210
rect 303 209 304 210
rect 302 209 303 210
rect 301 209 302 210
rect 300 209 301 210
rect 299 209 300 210
rect 298 209 299 210
rect 297 209 298 210
rect 296 209 297 210
rect 295 209 296 210
rect 294 209 295 210
rect 293 209 294 210
rect 292 209 293 210
rect 291 209 292 210
rect 290 209 291 210
rect 289 209 290 210
rect 288 209 289 210
rect 287 209 288 210
rect 286 209 287 210
rect 285 209 286 210
rect 284 209 285 210
rect 283 209 284 210
rect 282 209 283 210
rect 281 209 282 210
rect 280 209 281 210
rect 279 209 280 210
rect 278 209 279 210
rect 277 209 278 210
rect 276 209 277 210
rect 275 209 276 210
rect 274 209 275 210
rect 273 209 274 210
rect 272 209 273 210
rect 271 209 272 210
rect 270 209 271 210
rect 269 209 270 210
rect 268 209 269 210
rect 267 209 268 210
rect 266 209 267 210
rect 265 209 266 210
rect 264 209 265 210
rect 263 209 264 210
rect 262 209 263 210
rect 261 209 262 210
rect 260 209 261 210
rect 259 209 260 210
rect 258 209 259 210
rect 257 209 258 210
rect 256 209 257 210
rect 255 209 256 210
rect 254 209 255 210
rect 253 209 254 210
rect 252 209 253 210
rect 251 209 252 210
rect 250 209 251 210
rect 249 209 250 210
rect 248 209 249 210
rect 247 209 248 210
rect 246 209 247 210
rect 245 209 246 210
rect 244 209 245 210
rect 243 209 244 210
rect 242 209 243 210
rect 241 209 242 210
rect 240 209 241 210
rect 239 209 240 210
rect 238 209 239 210
rect 237 209 238 210
rect 236 209 237 210
rect 235 209 236 210
rect 234 209 235 210
rect 233 209 234 210
rect 232 209 233 210
rect 231 209 232 210
rect 230 209 231 210
rect 229 209 230 210
rect 228 209 229 210
rect 227 209 228 210
rect 226 209 227 210
rect 225 209 226 210
rect 224 209 225 210
rect 223 209 224 210
rect 222 209 223 210
rect 221 209 222 210
rect 220 209 221 210
rect 219 209 220 210
rect 218 209 219 210
rect 217 209 218 210
rect 216 209 217 210
rect 215 209 216 210
rect 214 209 215 210
rect 213 209 214 210
rect 212 209 213 210
rect 211 209 212 210
rect 210 209 211 210
rect 209 209 210 210
rect 208 209 209 210
rect 207 209 208 210
rect 206 209 207 210
rect 205 209 206 210
rect 204 209 205 210
rect 171 209 172 210
rect 170 209 171 210
rect 169 209 170 210
rect 168 209 169 210
rect 167 209 168 210
rect 166 209 167 210
rect 165 209 166 210
rect 164 209 165 210
rect 163 209 164 210
rect 162 209 163 210
rect 161 209 162 210
rect 160 209 161 210
rect 159 209 160 210
rect 158 209 159 210
rect 157 209 158 210
rect 156 209 157 210
rect 155 209 156 210
rect 154 209 155 210
rect 153 209 154 210
rect 152 209 153 210
rect 151 209 152 210
rect 150 209 151 210
rect 149 209 150 210
rect 148 209 149 210
rect 147 209 148 210
rect 146 209 147 210
rect 145 209 146 210
rect 144 209 145 210
rect 143 209 144 210
rect 142 209 143 210
rect 141 209 142 210
rect 140 209 141 210
rect 139 209 140 210
rect 138 209 139 210
rect 137 209 138 210
rect 136 209 137 210
rect 135 209 136 210
rect 134 209 135 210
rect 133 209 134 210
rect 132 209 133 210
rect 131 209 132 210
rect 130 209 131 210
rect 129 209 130 210
rect 128 209 129 210
rect 127 209 128 210
rect 126 209 127 210
rect 125 209 126 210
rect 124 209 125 210
rect 123 209 124 210
rect 122 209 123 210
rect 121 209 122 210
rect 120 209 121 210
rect 119 209 120 210
rect 118 209 119 210
rect 117 209 118 210
rect 116 209 117 210
rect 115 209 116 210
rect 114 209 115 210
rect 113 209 114 210
rect 112 209 113 210
rect 111 209 112 210
rect 110 209 111 210
rect 109 209 110 210
rect 108 209 109 210
rect 107 209 108 210
rect 106 209 107 210
rect 105 209 106 210
rect 104 209 105 210
rect 103 209 104 210
rect 102 209 103 210
rect 101 209 102 210
rect 100 209 101 210
rect 99 209 100 210
rect 98 209 99 210
rect 97 209 98 210
rect 96 209 97 210
rect 95 209 96 210
rect 94 209 95 210
rect 93 209 94 210
rect 92 209 93 210
rect 91 209 92 210
rect 90 209 91 210
rect 89 209 90 210
rect 88 209 89 210
rect 87 209 88 210
rect 86 209 87 210
rect 85 209 86 210
rect 84 209 85 210
rect 83 209 84 210
rect 82 209 83 210
rect 81 209 82 210
rect 80 209 81 210
rect 61 209 62 210
rect 60 209 61 210
rect 59 209 60 210
rect 58 209 59 210
rect 57 209 58 210
rect 56 209 57 210
rect 55 209 56 210
rect 54 209 55 210
rect 53 209 54 210
rect 52 209 53 210
rect 51 209 52 210
rect 50 209 51 210
rect 49 209 50 210
rect 48 209 49 210
rect 47 209 48 210
rect 46 209 47 210
rect 45 209 46 210
rect 44 209 45 210
rect 43 209 44 210
rect 42 209 43 210
rect 41 209 42 210
rect 40 209 41 210
rect 39 209 40 210
rect 38 209 39 210
rect 37 209 38 210
rect 36 209 37 210
rect 35 209 36 210
rect 34 209 35 210
rect 33 209 34 210
rect 32 209 33 210
rect 31 209 32 210
rect 30 209 31 210
rect 29 209 30 210
rect 28 209 29 210
rect 27 209 28 210
rect 26 209 27 210
rect 25 209 26 210
rect 24 209 25 210
rect 23 209 24 210
rect 22 209 23 210
rect 21 209 22 210
rect 20 209 21 210
rect 19 209 20 210
rect 18 209 19 210
rect 17 209 18 210
rect 16 209 17 210
rect 15 209 16 210
rect 14 209 15 210
rect 13 209 14 210
rect 12 209 13 210
rect 428 210 429 211
rect 427 210 428 211
rect 426 210 427 211
rect 425 210 426 211
rect 424 210 425 211
rect 423 210 424 211
rect 422 210 423 211
rect 421 210 422 211
rect 420 210 421 211
rect 419 210 420 211
rect 418 210 419 211
rect 417 210 418 211
rect 416 210 417 211
rect 415 210 416 211
rect 414 210 415 211
rect 413 210 414 211
rect 412 210 413 211
rect 357 210 358 211
rect 356 210 357 211
rect 355 210 356 211
rect 354 210 355 211
rect 353 210 354 211
rect 352 210 353 211
rect 351 210 352 211
rect 350 210 351 211
rect 349 210 350 211
rect 348 210 349 211
rect 347 210 348 211
rect 346 210 347 211
rect 345 210 346 211
rect 344 210 345 211
rect 343 210 344 211
rect 342 210 343 211
rect 341 210 342 211
rect 340 210 341 211
rect 339 210 340 211
rect 338 210 339 211
rect 337 210 338 211
rect 336 210 337 211
rect 335 210 336 211
rect 334 210 335 211
rect 333 210 334 211
rect 332 210 333 211
rect 331 210 332 211
rect 330 210 331 211
rect 329 210 330 211
rect 328 210 329 211
rect 327 210 328 211
rect 326 210 327 211
rect 325 210 326 211
rect 324 210 325 211
rect 323 210 324 211
rect 322 210 323 211
rect 321 210 322 211
rect 320 210 321 211
rect 319 210 320 211
rect 318 210 319 211
rect 317 210 318 211
rect 316 210 317 211
rect 315 210 316 211
rect 314 210 315 211
rect 313 210 314 211
rect 312 210 313 211
rect 311 210 312 211
rect 310 210 311 211
rect 309 210 310 211
rect 308 210 309 211
rect 307 210 308 211
rect 306 210 307 211
rect 305 210 306 211
rect 304 210 305 211
rect 303 210 304 211
rect 302 210 303 211
rect 301 210 302 211
rect 300 210 301 211
rect 299 210 300 211
rect 298 210 299 211
rect 297 210 298 211
rect 296 210 297 211
rect 295 210 296 211
rect 294 210 295 211
rect 293 210 294 211
rect 292 210 293 211
rect 291 210 292 211
rect 290 210 291 211
rect 289 210 290 211
rect 288 210 289 211
rect 287 210 288 211
rect 286 210 287 211
rect 285 210 286 211
rect 284 210 285 211
rect 283 210 284 211
rect 282 210 283 211
rect 281 210 282 211
rect 280 210 281 211
rect 279 210 280 211
rect 278 210 279 211
rect 277 210 278 211
rect 276 210 277 211
rect 275 210 276 211
rect 274 210 275 211
rect 273 210 274 211
rect 272 210 273 211
rect 271 210 272 211
rect 270 210 271 211
rect 269 210 270 211
rect 268 210 269 211
rect 267 210 268 211
rect 266 210 267 211
rect 265 210 266 211
rect 264 210 265 211
rect 263 210 264 211
rect 262 210 263 211
rect 261 210 262 211
rect 260 210 261 211
rect 259 210 260 211
rect 258 210 259 211
rect 257 210 258 211
rect 256 210 257 211
rect 255 210 256 211
rect 254 210 255 211
rect 253 210 254 211
rect 252 210 253 211
rect 251 210 252 211
rect 250 210 251 211
rect 249 210 250 211
rect 248 210 249 211
rect 247 210 248 211
rect 246 210 247 211
rect 245 210 246 211
rect 244 210 245 211
rect 243 210 244 211
rect 242 210 243 211
rect 241 210 242 211
rect 240 210 241 211
rect 239 210 240 211
rect 238 210 239 211
rect 237 210 238 211
rect 236 210 237 211
rect 235 210 236 211
rect 234 210 235 211
rect 233 210 234 211
rect 232 210 233 211
rect 231 210 232 211
rect 230 210 231 211
rect 229 210 230 211
rect 228 210 229 211
rect 227 210 228 211
rect 226 210 227 211
rect 225 210 226 211
rect 224 210 225 211
rect 223 210 224 211
rect 222 210 223 211
rect 221 210 222 211
rect 220 210 221 211
rect 219 210 220 211
rect 218 210 219 211
rect 217 210 218 211
rect 216 210 217 211
rect 215 210 216 211
rect 214 210 215 211
rect 213 210 214 211
rect 212 210 213 211
rect 211 210 212 211
rect 210 210 211 211
rect 209 210 210 211
rect 208 210 209 211
rect 207 210 208 211
rect 206 210 207 211
rect 205 210 206 211
rect 204 210 205 211
rect 203 210 204 211
rect 202 210 203 211
rect 169 210 170 211
rect 168 210 169 211
rect 167 210 168 211
rect 166 210 167 211
rect 165 210 166 211
rect 164 210 165 211
rect 163 210 164 211
rect 162 210 163 211
rect 161 210 162 211
rect 160 210 161 211
rect 159 210 160 211
rect 158 210 159 211
rect 157 210 158 211
rect 156 210 157 211
rect 155 210 156 211
rect 154 210 155 211
rect 153 210 154 211
rect 152 210 153 211
rect 151 210 152 211
rect 150 210 151 211
rect 149 210 150 211
rect 148 210 149 211
rect 147 210 148 211
rect 146 210 147 211
rect 145 210 146 211
rect 144 210 145 211
rect 143 210 144 211
rect 142 210 143 211
rect 141 210 142 211
rect 140 210 141 211
rect 139 210 140 211
rect 138 210 139 211
rect 137 210 138 211
rect 136 210 137 211
rect 135 210 136 211
rect 134 210 135 211
rect 133 210 134 211
rect 132 210 133 211
rect 131 210 132 211
rect 130 210 131 211
rect 129 210 130 211
rect 128 210 129 211
rect 127 210 128 211
rect 126 210 127 211
rect 125 210 126 211
rect 124 210 125 211
rect 123 210 124 211
rect 122 210 123 211
rect 121 210 122 211
rect 120 210 121 211
rect 119 210 120 211
rect 118 210 119 211
rect 117 210 118 211
rect 116 210 117 211
rect 115 210 116 211
rect 114 210 115 211
rect 113 210 114 211
rect 112 210 113 211
rect 111 210 112 211
rect 110 210 111 211
rect 109 210 110 211
rect 108 210 109 211
rect 107 210 108 211
rect 106 210 107 211
rect 105 210 106 211
rect 104 210 105 211
rect 103 210 104 211
rect 102 210 103 211
rect 101 210 102 211
rect 100 210 101 211
rect 99 210 100 211
rect 98 210 99 211
rect 97 210 98 211
rect 96 210 97 211
rect 95 210 96 211
rect 94 210 95 211
rect 93 210 94 211
rect 92 210 93 211
rect 91 210 92 211
rect 90 210 91 211
rect 89 210 90 211
rect 88 210 89 211
rect 87 210 88 211
rect 86 210 87 211
rect 85 210 86 211
rect 84 210 85 211
rect 83 210 84 211
rect 82 210 83 211
rect 81 210 82 211
rect 62 210 63 211
rect 61 210 62 211
rect 60 210 61 211
rect 59 210 60 211
rect 58 210 59 211
rect 57 210 58 211
rect 56 210 57 211
rect 55 210 56 211
rect 54 210 55 211
rect 53 210 54 211
rect 52 210 53 211
rect 51 210 52 211
rect 50 210 51 211
rect 49 210 50 211
rect 48 210 49 211
rect 47 210 48 211
rect 46 210 47 211
rect 45 210 46 211
rect 44 210 45 211
rect 43 210 44 211
rect 42 210 43 211
rect 41 210 42 211
rect 40 210 41 211
rect 39 210 40 211
rect 38 210 39 211
rect 37 210 38 211
rect 36 210 37 211
rect 35 210 36 211
rect 34 210 35 211
rect 33 210 34 211
rect 32 210 33 211
rect 31 210 32 211
rect 30 210 31 211
rect 29 210 30 211
rect 28 210 29 211
rect 27 210 28 211
rect 26 210 27 211
rect 25 210 26 211
rect 24 210 25 211
rect 23 210 24 211
rect 22 210 23 211
rect 21 210 22 211
rect 20 210 21 211
rect 19 210 20 211
rect 18 210 19 211
rect 17 210 18 211
rect 16 210 17 211
rect 15 210 16 211
rect 14 210 15 211
rect 13 210 14 211
rect 12 210 13 211
rect 430 211 431 212
rect 429 211 430 212
rect 428 211 429 212
rect 427 211 428 212
rect 426 211 427 212
rect 425 211 426 212
rect 424 211 425 212
rect 423 211 424 212
rect 422 211 423 212
rect 421 211 422 212
rect 420 211 421 212
rect 419 211 420 212
rect 418 211 419 212
rect 417 211 418 212
rect 416 211 417 212
rect 415 211 416 212
rect 414 211 415 212
rect 413 211 414 212
rect 412 211 413 212
rect 411 211 412 212
rect 410 211 411 212
rect 409 211 410 212
rect 357 211 358 212
rect 356 211 357 212
rect 355 211 356 212
rect 354 211 355 212
rect 353 211 354 212
rect 352 211 353 212
rect 351 211 352 212
rect 350 211 351 212
rect 349 211 350 212
rect 348 211 349 212
rect 347 211 348 212
rect 346 211 347 212
rect 345 211 346 212
rect 344 211 345 212
rect 343 211 344 212
rect 342 211 343 212
rect 341 211 342 212
rect 340 211 341 212
rect 339 211 340 212
rect 338 211 339 212
rect 337 211 338 212
rect 336 211 337 212
rect 335 211 336 212
rect 334 211 335 212
rect 333 211 334 212
rect 332 211 333 212
rect 331 211 332 212
rect 330 211 331 212
rect 329 211 330 212
rect 328 211 329 212
rect 327 211 328 212
rect 326 211 327 212
rect 325 211 326 212
rect 324 211 325 212
rect 323 211 324 212
rect 322 211 323 212
rect 321 211 322 212
rect 320 211 321 212
rect 319 211 320 212
rect 318 211 319 212
rect 317 211 318 212
rect 316 211 317 212
rect 315 211 316 212
rect 314 211 315 212
rect 313 211 314 212
rect 312 211 313 212
rect 311 211 312 212
rect 310 211 311 212
rect 309 211 310 212
rect 308 211 309 212
rect 307 211 308 212
rect 306 211 307 212
rect 305 211 306 212
rect 304 211 305 212
rect 303 211 304 212
rect 302 211 303 212
rect 301 211 302 212
rect 300 211 301 212
rect 299 211 300 212
rect 298 211 299 212
rect 297 211 298 212
rect 296 211 297 212
rect 295 211 296 212
rect 294 211 295 212
rect 293 211 294 212
rect 292 211 293 212
rect 291 211 292 212
rect 290 211 291 212
rect 289 211 290 212
rect 288 211 289 212
rect 287 211 288 212
rect 286 211 287 212
rect 285 211 286 212
rect 284 211 285 212
rect 283 211 284 212
rect 282 211 283 212
rect 281 211 282 212
rect 280 211 281 212
rect 279 211 280 212
rect 278 211 279 212
rect 277 211 278 212
rect 276 211 277 212
rect 275 211 276 212
rect 274 211 275 212
rect 273 211 274 212
rect 272 211 273 212
rect 271 211 272 212
rect 270 211 271 212
rect 269 211 270 212
rect 268 211 269 212
rect 267 211 268 212
rect 266 211 267 212
rect 265 211 266 212
rect 264 211 265 212
rect 263 211 264 212
rect 262 211 263 212
rect 261 211 262 212
rect 260 211 261 212
rect 259 211 260 212
rect 258 211 259 212
rect 257 211 258 212
rect 256 211 257 212
rect 255 211 256 212
rect 254 211 255 212
rect 253 211 254 212
rect 252 211 253 212
rect 251 211 252 212
rect 250 211 251 212
rect 249 211 250 212
rect 248 211 249 212
rect 247 211 248 212
rect 246 211 247 212
rect 245 211 246 212
rect 244 211 245 212
rect 243 211 244 212
rect 242 211 243 212
rect 241 211 242 212
rect 240 211 241 212
rect 239 211 240 212
rect 238 211 239 212
rect 237 211 238 212
rect 236 211 237 212
rect 235 211 236 212
rect 234 211 235 212
rect 233 211 234 212
rect 232 211 233 212
rect 231 211 232 212
rect 230 211 231 212
rect 229 211 230 212
rect 228 211 229 212
rect 227 211 228 212
rect 226 211 227 212
rect 225 211 226 212
rect 224 211 225 212
rect 223 211 224 212
rect 222 211 223 212
rect 221 211 222 212
rect 220 211 221 212
rect 219 211 220 212
rect 218 211 219 212
rect 217 211 218 212
rect 216 211 217 212
rect 215 211 216 212
rect 214 211 215 212
rect 213 211 214 212
rect 212 211 213 212
rect 211 211 212 212
rect 210 211 211 212
rect 209 211 210 212
rect 208 211 209 212
rect 207 211 208 212
rect 206 211 207 212
rect 205 211 206 212
rect 204 211 205 212
rect 203 211 204 212
rect 202 211 203 212
rect 201 211 202 212
rect 167 211 168 212
rect 166 211 167 212
rect 165 211 166 212
rect 164 211 165 212
rect 163 211 164 212
rect 162 211 163 212
rect 161 211 162 212
rect 160 211 161 212
rect 159 211 160 212
rect 158 211 159 212
rect 157 211 158 212
rect 156 211 157 212
rect 155 211 156 212
rect 154 211 155 212
rect 153 211 154 212
rect 152 211 153 212
rect 151 211 152 212
rect 150 211 151 212
rect 149 211 150 212
rect 148 211 149 212
rect 147 211 148 212
rect 146 211 147 212
rect 145 211 146 212
rect 144 211 145 212
rect 143 211 144 212
rect 142 211 143 212
rect 141 211 142 212
rect 140 211 141 212
rect 139 211 140 212
rect 138 211 139 212
rect 137 211 138 212
rect 136 211 137 212
rect 135 211 136 212
rect 134 211 135 212
rect 133 211 134 212
rect 132 211 133 212
rect 131 211 132 212
rect 130 211 131 212
rect 129 211 130 212
rect 128 211 129 212
rect 127 211 128 212
rect 126 211 127 212
rect 125 211 126 212
rect 124 211 125 212
rect 123 211 124 212
rect 122 211 123 212
rect 121 211 122 212
rect 120 211 121 212
rect 119 211 120 212
rect 118 211 119 212
rect 117 211 118 212
rect 116 211 117 212
rect 115 211 116 212
rect 114 211 115 212
rect 113 211 114 212
rect 112 211 113 212
rect 111 211 112 212
rect 110 211 111 212
rect 109 211 110 212
rect 108 211 109 212
rect 107 211 108 212
rect 106 211 107 212
rect 105 211 106 212
rect 104 211 105 212
rect 103 211 104 212
rect 102 211 103 212
rect 101 211 102 212
rect 100 211 101 212
rect 99 211 100 212
rect 98 211 99 212
rect 97 211 98 212
rect 96 211 97 212
rect 95 211 96 212
rect 94 211 95 212
rect 93 211 94 212
rect 92 211 93 212
rect 91 211 92 212
rect 90 211 91 212
rect 89 211 90 212
rect 88 211 89 212
rect 87 211 88 212
rect 86 211 87 212
rect 85 211 86 212
rect 84 211 85 212
rect 83 211 84 212
rect 63 211 64 212
rect 62 211 63 212
rect 61 211 62 212
rect 60 211 61 212
rect 59 211 60 212
rect 58 211 59 212
rect 57 211 58 212
rect 56 211 57 212
rect 55 211 56 212
rect 54 211 55 212
rect 53 211 54 212
rect 52 211 53 212
rect 51 211 52 212
rect 50 211 51 212
rect 49 211 50 212
rect 48 211 49 212
rect 47 211 48 212
rect 46 211 47 212
rect 45 211 46 212
rect 44 211 45 212
rect 43 211 44 212
rect 42 211 43 212
rect 41 211 42 212
rect 40 211 41 212
rect 39 211 40 212
rect 38 211 39 212
rect 37 211 38 212
rect 36 211 37 212
rect 35 211 36 212
rect 34 211 35 212
rect 33 211 34 212
rect 32 211 33 212
rect 31 211 32 212
rect 30 211 31 212
rect 29 211 30 212
rect 28 211 29 212
rect 27 211 28 212
rect 26 211 27 212
rect 25 211 26 212
rect 24 211 25 212
rect 23 211 24 212
rect 22 211 23 212
rect 21 211 22 212
rect 20 211 21 212
rect 19 211 20 212
rect 18 211 19 212
rect 17 211 18 212
rect 16 211 17 212
rect 15 211 16 212
rect 14 211 15 212
rect 13 211 14 212
rect 12 211 13 212
rect 11 211 12 212
rect 432 212 433 213
rect 431 212 432 213
rect 430 212 431 213
rect 429 212 430 213
rect 428 212 429 213
rect 427 212 428 213
rect 426 212 427 213
rect 425 212 426 213
rect 424 212 425 213
rect 423 212 424 213
rect 422 212 423 213
rect 421 212 422 213
rect 420 212 421 213
rect 419 212 420 213
rect 418 212 419 213
rect 417 212 418 213
rect 416 212 417 213
rect 415 212 416 213
rect 414 212 415 213
rect 413 212 414 213
rect 412 212 413 213
rect 411 212 412 213
rect 410 212 411 213
rect 409 212 410 213
rect 408 212 409 213
rect 407 212 408 213
rect 358 212 359 213
rect 357 212 358 213
rect 356 212 357 213
rect 355 212 356 213
rect 354 212 355 213
rect 353 212 354 213
rect 352 212 353 213
rect 351 212 352 213
rect 350 212 351 213
rect 349 212 350 213
rect 348 212 349 213
rect 347 212 348 213
rect 346 212 347 213
rect 345 212 346 213
rect 344 212 345 213
rect 343 212 344 213
rect 342 212 343 213
rect 341 212 342 213
rect 340 212 341 213
rect 339 212 340 213
rect 338 212 339 213
rect 337 212 338 213
rect 336 212 337 213
rect 335 212 336 213
rect 334 212 335 213
rect 333 212 334 213
rect 332 212 333 213
rect 331 212 332 213
rect 330 212 331 213
rect 329 212 330 213
rect 328 212 329 213
rect 327 212 328 213
rect 326 212 327 213
rect 325 212 326 213
rect 324 212 325 213
rect 323 212 324 213
rect 322 212 323 213
rect 321 212 322 213
rect 320 212 321 213
rect 319 212 320 213
rect 318 212 319 213
rect 317 212 318 213
rect 316 212 317 213
rect 315 212 316 213
rect 314 212 315 213
rect 313 212 314 213
rect 312 212 313 213
rect 311 212 312 213
rect 310 212 311 213
rect 309 212 310 213
rect 308 212 309 213
rect 307 212 308 213
rect 306 212 307 213
rect 305 212 306 213
rect 304 212 305 213
rect 303 212 304 213
rect 302 212 303 213
rect 301 212 302 213
rect 300 212 301 213
rect 299 212 300 213
rect 298 212 299 213
rect 297 212 298 213
rect 296 212 297 213
rect 295 212 296 213
rect 294 212 295 213
rect 293 212 294 213
rect 292 212 293 213
rect 291 212 292 213
rect 290 212 291 213
rect 289 212 290 213
rect 288 212 289 213
rect 287 212 288 213
rect 286 212 287 213
rect 285 212 286 213
rect 284 212 285 213
rect 283 212 284 213
rect 282 212 283 213
rect 281 212 282 213
rect 280 212 281 213
rect 279 212 280 213
rect 278 212 279 213
rect 277 212 278 213
rect 276 212 277 213
rect 275 212 276 213
rect 274 212 275 213
rect 273 212 274 213
rect 272 212 273 213
rect 271 212 272 213
rect 270 212 271 213
rect 269 212 270 213
rect 268 212 269 213
rect 267 212 268 213
rect 266 212 267 213
rect 265 212 266 213
rect 264 212 265 213
rect 263 212 264 213
rect 262 212 263 213
rect 261 212 262 213
rect 260 212 261 213
rect 259 212 260 213
rect 258 212 259 213
rect 257 212 258 213
rect 256 212 257 213
rect 255 212 256 213
rect 254 212 255 213
rect 253 212 254 213
rect 252 212 253 213
rect 251 212 252 213
rect 250 212 251 213
rect 249 212 250 213
rect 248 212 249 213
rect 247 212 248 213
rect 246 212 247 213
rect 245 212 246 213
rect 244 212 245 213
rect 243 212 244 213
rect 242 212 243 213
rect 241 212 242 213
rect 240 212 241 213
rect 239 212 240 213
rect 238 212 239 213
rect 237 212 238 213
rect 236 212 237 213
rect 235 212 236 213
rect 234 212 235 213
rect 233 212 234 213
rect 232 212 233 213
rect 231 212 232 213
rect 230 212 231 213
rect 229 212 230 213
rect 228 212 229 213
rect 227 212 228 213
rect 226 212 227 213
rect 225 212 226 213
rect 224 212 225 213
rect 223 212 224 213
rect 222 212 223 213
rect 221 212 222 213
rect 220 212 221 213
rect 219 212 220 213
rect 218 212 219 213
rect 217 212 218 213
rect 216 212 217 213
rect 215 212 216 213
rect 214 212 215 213
rect 213 212 214 213
rect 212 212 213 213
rect 211 212 212 213
rect 210 212 211 213
rect 209 212 210 213
rect 208 212 209 213
rect 207 212 208 213
rect 206 212 207 213
rect 205 212 206 213
rect 204 212 205 213
rect 203 212 204 213
rect 202 212 203 213
rect 201 212 202 213
rect 200 212 201 213
rect 164 212 165 213
rect 163 212 164 213
rect 162 212 163 213
rect 161 212 162 213
rect 160 212 161 213
rect 159 212 160 213
rect 158 212 159 213
rect 157 212 158 213
rect 156 212 157 213
rect 155 212 156 213
rect 154 212 155 213
rect 153 212 154 213
rect 152 212 153 213
rect 151 212 152 213
rect 150 212 151 213
rect 149 212 150 213
rect 148 212 149 213
rect 147 212 148 213
rect 146 212 147 213
rect 145 212 146 213
rect 144 212 145 213
rect 143 212 144 213
rect 142 212 143 213
rect 141 212 142 213
rect 140 212 141 213
rect 139 212 140 213
rect 138 212 139 213
rect 137 212 138 213
rect 136 212 137 213
rect 135 212 136 213
rect 134 212 135 213
rect 133 212 134 213
rect 132 212 133 213
rect 131 212 132 213
rect 130 212 131 213
rect 129 212 130 213
rect 128 212 129 213
rect 127 212 128 213
rect 126 212 127 213
rect 125 212 126 213
rect 124 212 125 213
rect 123 212 124 213
rect 122 212 123 213
rect 121 212 122 213
rect 120 212 121 213
rect 119 212 120 213
rect 118 212 119 213
rect 117 212 118 213
rect 116 212 117 213
rect 115 212 116 213
rect 114 212 115 213
rect 113 212 114 213
rect 112 212 113 213
rect 111 212 112 213
rect 110 212 111 213
rect 109 212 110 213
rect 108 212 109 213
rect 107 212 108 213
rect 106 212 107 213
rect 105 212 106 213
rect 104 212 105 213
rect 103 212 104 213
rect 102 212 103 213
rect 101 212 102 213
rect 100 212 101 213
rect 99 212 100 213
rect 98 212 99 213
rect 97 212 98 213
rect 96 212 97 213
rect 95 212 96 213
rect 94 212 95 213
rect 93 212 94 213
rect 92 212 93 213
rect 91 212 92 213
rect 90 212 91 213
rect 89 212 90 213
rect 88 212 89 213
rect 87 212 88 213
rect 86 212 87 213
rect 85 212 86 213
rect 84 212 85 213
rect 63 212 64 213
rect 62 212 63 213
rect 61 212 62 213
rect 60 212 61 213
rect 59 212 60 213
rect 58 212 59 213
rect 57 212 58 213
rect 56 212 57 213
rect 55 212 56 213
rect 54 212 55 213
rect 53 212 54 213
rect 52 212 53 213
rect 51 212 52 213
rect 50 212 51 213
rect 49 212 50 213
rect 48 212 49 213
rect 47 212 48 213
rect 46 212 47 213
rect 45 212 46 213
rect 44 212 45 213
rect 43 212 44 213
rect 42 212 43 213
rect 41 212 42 213
rect 40 212 41 213
rect 39 212 40 213
rect 38 212 39 213
rect 37 212 38 213
rect 36 212 37 213
rect 35 212 36 213
rect 34 212 35 213
rect 33 212 34 213
rect 32 212 33 213
rect 31 212 32 213
rect 30 212 31 213
rect 29 212 30 213
rect 28 212 29 213
rect 27 212 28 213
rect 26 212 27 213
rect 25 212 26 213
rect 24 212 25 213
rect 23 212 24 213
rect 22 212 23 213
rect 21 212 22 213
rect 20 212 21 213
rect 19 212 20 213
rect 18 212 19 213
rect 17 212 18 213
rect 16 212 17 213
rect 15 212 16 213
rect 14 212 15 213
rect 13 212 14 213
rect 12 212 13 213
rect 11 212 12 213
rect 433 213 434 214
rect 432 213 433 214
rect 431 213 432 214
rect 430 213 431 214
rect 429 213 430 214
rect 428 213 429 214
rect 427 213 428 214
rect 426 213 427 214
rect 425 213 426 214
rect 424 213 425 214
rect 423 213 424 214
rect 422 213 423 214
rect 421 213 422 214
rect 420 213 421 214
rect 419 213 420 214
rect 418 213 419 214
rect 417 213 418 214
rect 416 213 417 214
rect 415 213 416 214
rect 414 213 415 214
rect 413 213 414 214
rect 412 213 413 214
rect 411 213 412 214
rect 410 213 411 214
rect 409 213 410 214
rect 408 213 409 214
rect 407 213 408 214
rect 406 213 407 214
rect 358 213 359 214
rect 357 213 358 214
rect 356 213 357 214
rect 355 213 356 214
rect 354 213 355 214
rect 353 213 354 214
rect 352 213 353 214
rect 351 213 352 214
rect 350 213 351 214
rect 349 213 350 214
rect 348 213 349 214
rect 347 213 348 214
rect 346 213 347 214
rect 345 213 346 214
rect 344 213 345 214
rect 343 213 344 214
rect 342 213 343 214
rect 341 213 342 214
rect 340 213 341 214
rect 339 213 340 214
rect 338 213 339 214
rect 337 213 338 214
rect 336 213 337 214
rect 335 213 336 214
rect 334 213 335 214
rect 333 213 334 214
rect 332 213 333 214
rect 331 213 332 214
rect 330 213 331 214
rect 329 213 330 214
rect 328 213 329 214
rect 327 213 328 214
rect 326 213 327 214
rect 325 213 326 214
rect 324 213 325 214
rect 323 213 324 214
rect 322 213 323 214
rect 321 213 322 214
rect 320 213 321 214
rect 319 213 320 214
rect 318 213 319 214
rect 317 213 318 214
rect 316 213 317 214
rect 315 213 316 214
rect 314 213 315 214
rect 313 213 314 214
rect 312 213 313 214
rect 311 213 312 214
rect 310 213 311 214
rect 309 213 310 214
rect 308 213 309 214
rect 307 213 308 214
rect 306 213 307 214
rect 305 213 306 214
rect 304 213 305 214
rect 303 213 304 214
rect 302 213 303 214
rect 301 213 302 214
rect 300 213 301 214
rect 299 213 300 214
rect 298 213 299 214
rect 297 213 298 214
rect 296 213 297 214
rect 295 213 296 214
rect 294 213 295 214
rect 293 213 294 214
rect 292 213 293 214
rect 291 213 292 214
rect 290 213 291 214
rect 289 213 290 214
rect 288 213 289 214
rect 287 213 288 214
rect 286 213 287 214
rect 285 213 286 214
rect 284 213 285 214
rect 283 213 284 214
rect 282 213 283 214
rect 281 213 282 214
rect 280 213 281 214
rect 279 213 280 214
rect 278 213 279 214
rect 277 213 278 214
rect 276 213 277 214
rect 275 213 276 214
rect 274 213 275 214
rect 273 213 274 214
rect 272 213 273 214
rect 271 213 272 214
rect 270 213 271 214
rect 269 213 270 214
rect 268 213 269 214
rect 267 213 268 214
rect 266 213 267 214
rect 265 213 266 214
rect 264 213 265 214
rect 263 213 264 214
rect 262 213 263 214
rect 261 213 262 214
rect 260 213 261 214
rect 259 213 260 214
rect 258 213 259 214
rect 257 213 258 214
rect 256 213 257 214
rect 255 213 256 214
rect 254 213 255 214
rect 253 213 254 214
rect 252 213 253 214
rect 251 213 252 214
rect 250 213 251 214
rect 249 213 250 214
rect 248 213 249 214
rect 247 213 248 214
rect 246 213 247 214
rect 245 213 246 214
rect 244 213 245 214
rect 243 213 244 214
rect 242 213 243 214
rect 241 213 242 214
rect 240 213 241 214
rect 239 213 240 214
rect 238 213 239 214
rect 237 213 238 214
rect 236 213 237 214
rect 235 213 236 214
rect 234 213 235 214
rect 233 213 234 214
rect 232 213 233 214
rect 231 213 232 214
rect 230 213 231 214
rect 229 213 230 214
rect 228 213 229 214
rect 227 213 228 214
rect 226 213 227 214
rect 225 213 226 214
rect 224 213 225 214
rect 223 213 224 214
rect 222 213 223 214
rect 221 213 222 214
rect 220 213 221 214
rect 219 213 220 214
rect 218 213 219 214
rect 217 213 218 214
rect 216 213 217 214
rect 215 213 216 214
rect 214 213 215 214
rect 213 213 214 214
rect 212 213 213 214
rect 211 213 212 214
rect 210 213 211 214
rect 209 213 210 214
rect 208 213 209 214
rect 207 213 208 214
rect 206 213 207 214
rect 205 213 206 214
rect 204 213 205 214
rect 203 213 204 214
rect 202 213 203 214
rect 201 213 202 214
rect 200 213 201 214
rect 199 213 200 214
rect 198 213 199 214
rect 161 213 162 214
rect 160 213 161 214
rect 159 213 160 214
rect 158 213 159 214
rect 157 213 158 214
rect 156 213 157 214
rect 155 213 156 214
rect 154 213 155 214
rect 153 213 154 214
rect 152 213 153 214
rect 151 213 152 214
rect 150 213 151 214
rect 149 213 150 214
rect 148 213 149 214
rect 147 213 148 214
rect 146 213 147 214
rect 145 213 146 214
rect 144 213 145 214
rect 143 213 144 214
rect 142 213 143 214
rect 141 213 142 214
rect 140 213 141 214
rect 139 213 140 214
rect 138 213 139 214
rect 137 213 138 214
rect 136 213 137 214
rect 135 213 136 214
rect 134 213 135 214
rect 133 213 134 214
rect 132 213 133 214
rect 131 213 132 214
rect 130 213 131 214
rect 129 213 130 214
rect 128 213 129 214
rect 127 213 128 214
rect 126 213 127 214
rect 125 213 126 214
rect 124 213 125 214
rect 123 213 124 214
rect 122 213 123 214
rect 121 213 122 214
rect 120 213 121 214
rect 119 213 120 214
rect 118 213 119 214
rect 117 213 118 214
rect 116 213 117 214
rect 115 213 116 214
rect 114 213 115 214
rect 113 213 114 214
rect 112 213 113 214
rect 111 213 112 214
rect 110 213 111 214
rect 109 213 110 214
rect 108 213 109 214
rect 107 213 108 214
rect 106 213 107 214
rect 105 213 106 214
rect 104 213 105 214
rect 103 213 104 214
rect 102 213 103 214
rect 101 213 102 214
rect 100 213 101 214
rect 99 213 100 214
rect 98 213 99 214
rect 97 213 98 214
rect 96 213 97 214
rect 95 213 96 214
rect 94 213 95 214
rect 93 213 94 214
rect 92 213 93 214
rect 91 213 92 214
rect 90 213 91 214
rect 89 213 90 214
rect 88 213 89 214
rect 87 213 88 214
rect 86 213 87 214
rect 64 213 65 214
rect 63 213 64 214
rect 62 213 63 214
rect 61 213 62 214
rect 60 213 61 214
rect 59 213 60 214
rect 58 213 59 214
rect 57 213 58 214
rect 56 213 57 214
rect 55 213 56 214
rect 54 213 55 214
rect 53 213 54 214
rect 52 213 53 214
rect 51 213 52 214
rect 50 213 51 214
rect 49 213 50 214
rect 48 213 49 214
rect 47 213 48 214
rect 46 213 47 214
rect 45 213 46 214
rect 44 213 45 214
rect 43 213 44 214
rect 42 213 43 214
rect 41 213 42 214
rect 40 213 41 214
rect 39 213 40 214
rect 38 213 39 214
rect 37 213 38 214
rect 36 213 37 214
rect 35 213 36 214
rect 34 213 35 214
rect 33 213 34 214
rect 32 213 33 214
rect 31 213 32 214
rect 30 213 31 214
rect 29 213 30 214
rect 28 213 29 214
rect 27 213 28 214
rect 26 213 27 214
rect 25 213 26 214
rect 24 213 25 214
rect 23 213 24 214
rect 22 213 23 214
rect 21 213 22 214
rect 20 213 21 214
rect 19 213 20 214
rect 18 213 19 214
rect 17 213 18 214
rect 16 213 17 214
rect 15 213 16 214
rect 14 213 15 214
rect 13 213 14 214
rect 12 213 13 214
rect 11 213 12 214
rect 434 214 435 215
rect 433 214 434 215
rect 432 214 433 215
rect 431 214 432 215
rect 430 214 431 215
rect 429 214 430 215
rect 428 214 429 215
rect 427 214 428 215
rect 426 214 427 215
rect 425 214 426 215
rect 424 214 425 215
rect 423 214 424 215
rect 422 214 423 215
rect 421 214 422 215
rect 420 214 421 215
rect 419 214 420 215
rect 418 214 419 215
rect 417 214 418 215
rect 416 214 417 215
rect 415 214 416 215
rect 414 214 415 215
rect 413 214 414 215
rect 412 214 413 215
rect 411 214 412 215
rect 410 214 411 215
rect 409 214 410 215
rect 408 214 409 215
rect 407 214 408 215
rect 406 214 407 215
rect 405 214 406 215
rect 359 214 360 215
rect 358 214 359 215
rect 357 214 358 215
rect 356 214 357 215
rect 355 214 356 215
rect 354 214 355 215
rect 353 214 354 215
rect 352 214 353 215
rect 351 214 352 215
rect 350 214 351 215
rect 349 214 350 215
rect 348 214 349 215
rect 347 214 348 215
rect 346 214 347 215
rect 345 214 346 215
rect 344 214 345 215
rect 343 214 344 215
rect 342 214 343 215
rect 341 214 342 215
rect 340 214 341 215
rect 339 214 340 215
rect 338 214 339 215
rect 337 214 338 215
rect 336 214 337 215
rect 335 214 336 215
rect 334 214 335 215
rect 333 214 334 215
rect 332 214 333 215
rect 331 214 332 215
rect 330 214 331 215
rect 329 214 330 215
rect 328 214 329 215
rect 327 214 328 215
rect 326 214 327 215
rect 325 214 326 215
rect 324 214 325 215
rect 323 214 324 215
rect 322 214 323 215
rect 321 214 322 215
rect 320 214 321 215
rect 319 214 320 215
rect 318 214 319 215
rect 317 214 318 215
rect 316 214 317 215
rect 315 214 316 215
rect 314 214 315 215
rect 313 214 314 215
rect 312 214 313 215
rect 311 214 312 215
rect 310 214 311 215
rect 309 214 310 215
rect 308 214 309 215
rect 307 214 308 215
rect 306 214 307 215
rect 305 214 306 215
rect 304 214 305 215
rect 303 214 304 215
rect 302 214 303 215
rect 301 214 302 215
rect 300 214 301 215
rect 299 214 300 215
rect 298 214 299 215
rect 297 214 298 215
rect 296 214 297 215
rect 295 214 296 215
rect 294 214 295 215
rect 293 214 294 215
rect 292 214 293 215
rect 291 214 292 215
rect 290 214 291 215
rect 289 214 290 215
rect 288 214 289 215
rect 287 214 288 215
rect 286 214 287 215
rect 285 214 286 215
rect 284 214 285 215
rect 283 214 284 215
rect 282 214 283 215
rect 281 214 282 215
rect 280 214 281 215
rect 279 214 280 215
rect 278 214 279 215
rect 277 214 278 215
rect 276 214 277 215
rect 275 214 276 215
rect 274 214 275 215
rect 273 214 274 215
rect 272 214 273 215
rect 271 214 272 215
rect 270 214 271 215
rect 269 214 270 215
rect 268 214 269 215
rect 267 214 268 215
rect 266 214 267 215
rect 265 214 266 215
rect 264 214 265 215
rect 263 214 264 215
rect 262 214 263 215
rect 261 214 262 215
rect 260 214 261 215
rect 259 214 260 215
rect 258 214 259 215
rect 257 214 258 215
rect 256 214 257 215
rect 255 214 256 215
rect 254 214 255 215
rect 253 214 254 215
rect 252 214 253 215
rect 251 214 252 215
rect 250 214 251 215
rect 249 214 250 215
rect 248 214 249 215
rect 247 214 248 215
rect 246 214 247 215
rect 245 214 246 215
rect 244 214 245 215
rect 243 214 244 215
rect 242 214 243 215
rect 241 214 242 215
rect 240 214 241 215
rect 239 214 240 215
rect 238 214 239 215
rect 237 214 238 215
rect 236 214 237 215
rect 235 214 236 215
rect 234 214 235 215
rect 233 214 234 215
rect 232 214 233 215
rect 231 214 232 215
rect 230 214 231 215
rect 229 214 230 215
rect 228 214 229 215
rect 227 214 228 215
rect 226 214 227 215
rect 225 214 226 215
rect 224 214 225 215
rect 223 214 224 215
rect 222 214 223 215
rect 221 214 222 215
rect 220 214 221 215
rect 219 214 220 215
rect 218 214 219 215
rect 217 214 218 215
rect 216 214 217 215
rect 215 214 216 215
rect 214 214 215 215
rect 213 214 214 215
rect 212 214 213 215
rect 211 214 212 215
rect 210 214 211 215
rect 209 214 210 215
rect 208 214 209 215
rect 207 214 208 215
rect 206 214 207 215
rect 205 214 206 215
rect 204 214 205 215
rect 203 214 204 215
rect 202 214 203 215
rect 201 214 202 215
rect 200 214 201 215
rect 199 214 200 215
rect 198 214 199 215
rect 197 214 198 215
rect 158 214 159 215
rect 157 214 158 215
rect 156 214 157 215
rect 155 214 156 215
rect 154 214 155 215
rect 153 214 154 215
rect 152 214 153 215
rect 151 214 152 215
rect 150 214 151 215
rect 149 214 150 215
rect 148 214 149 215
rect 147 214 148 215
rect 146 214 147 215
rect 145 214 146 215
rect 144 214 145 215
rect 143 214 144 215
rect 142 214 143 215
rect 141 214 142 215
rect 140 214 141 215
rect 139 214 140 215
rect 138 214 139 215
rect 137 214 138 215
rect 136 214 137 215
rect 135 214 136 215
rect 134 214 135 215
rect 133 214 134 215
rect 132 214 133 215
rect 131 214 132 215
rect 130 214 131 215
rect 129 214 130 215
rect 128 214 129 215
rect 127 214 128 215
rect 126 214 127 215
rect 125 214 126 215
rect 124 214 125 215
rect 123 214 124 215
rect 122 214 123 215
rect 121 214 122 215
rect 120 214 121 215
rect 119 214 120 215
rect 118 214 119 215
rect 117 214 118 215
rect 116 214 117 215
rect 115 214 116 215
rect 114 214 115 215
rect 113 214 114 215
rect 112 214 113 215
rect 111 214 112 215
rect 110 214 111 215
rect 109 214 110 215
rect 108 214 109 215
rect 107 214 108 215
rect 106 214 107 215
rect 105 214 106 215
rect 104 214 105 215
rect 103 214 104 215
rect 102 214 103 215
rect 101 214 102 215
rect 100 214 101 215
rect 99 214 100 215
rect 98 214 99 215
rect 97 214 98 215
rect 96 214 97 215
rect 95 214 96 215
rect 94 214 95 215
rect 93 214 94 215
rect 92 214 93 215
rect 91 214 92 215
rect 90 214 91 215
rect 89 214 90 215
rect 88 214 89 215
rect 65 214 66 215
rect 64 214 65 215
rect 63 214 64 215
rect 62 214 63 215
rect 61 214 62 215
rect 60 214 61 215
rect 59 214 60 215
rect 58 214 59 215
rect 57 214 58 215
rect 56 214 57 215
rect 55 214 56 215
rect 54 214 55 215
rect 53 214 54 215
rect 52 214 53 215
rect 51 214 52 215
rect 50 214 51 215
rect 49 214 50 215
rect 48 214 49 215
rect 47 214 48 215
rect 46 214 47 215
rect 45 214 46 215
rect 44 214 45 215
rect 43 214 44 215
rect 42 214 43 215
rect 41 214 42 215
rect 40 214 41 215
rect 39 214 40 215
rect 38 214 39 215
rect 37 214 38 215
rect 36 214 37 215
rect 35 214 36 215
rect 34 214 35 215
rect 33 214 34 215
rect 32 214 33 215
rect 31 214 32 215
rect 30 214 31 215
rect 29 214 30 215
rect 28 214 29 215
rect 27 214 28 215
rect 26 214 27 215
rect 25 214 26 215
rect 24 214 25 215
rect 23 214 24 215
rect 22 214 23 215
rect 21 214 22 215
rect 20 214 21 215
rect 19 214 20 215
rect 18 214 19 215
rect 17 214 18 215
rect 16 214 17 215
rect 15 214 16 215
rect 14 214 15 215
rect 13 214 14 215
rect 12 214 13 215
rect 11 214 12 215
rect 435 215 436 216
rect 434 215 435 216
rect 433 215 434 216
rect 432 215 433 216
rect 431 215 432 216
rect 430 215 431 216
rect 429 215 430 216
rect 428 215 429 216
rect 427 215 428 216
rect 426 215 427 216
rect 425 215 426 216
rect 424 215 425 216
rect 423 215 424 216
rect 422 215 423 216
rect 421 215 422 216
rect 420 215 421 216
rect 419 215 420 216
rect 418 215 419 216
rect 417 215 418 216
rect 416 215 417 216
rect 415 215 416 216
rect 414 215 415 216
rect 413 215 414 216
rect 412 215 413 216
rect 411 215 412 216
rect 410 215 411 216
rect 409 215 410 216
rect 408 215 409 216
rect 407 215 408 216
rect 406 215 407 216
rect 405 215 406 216
rect 404 215 405 216
rect 360 215 361 216
rect 359 215 360 216
rect 358 215 359 216
rect 357 215 358 216
rect 356 215 357 216
rect 355 215 356 216
rect 354 215 355 216
rect 353 215 354 216
rect 352 215 353 216
rect 351 215 352 216
rect 350 215 351 216
rect 349 215 350 216
rect 348 215 349 216
rect 347 215 348 216
rect 346 215 347 216
rect 345 215 346 216
rect 344 215 345 216
rect 343 215 344 216
rect 342 215 343 216
rect 341 215 342 216
rect 340 215 341 216
rect 339 215 340 216
rect 338 215 339 216
rect 337 215 338 216
rect 336 215 337 216
rect 335 215 336 216
rect 334 215 335 216
rect 333 215 334 216
rect 332 215 333 216
rect 331 215 332 216
rect 330 215 331 216
rect 329 215 330 216
rect 328 215 329 216
rect 327 215 328 216
rect 326 215 327 216
rect 325 215 326 216
rect 324 215 325 216
rect 323 215 324 216
rect 322 215 323 216
rect 321 215 322 216
rect 320 215 321 216
rect 319 215 320 216
rect 318 215 319 216
rect 317 215 318 216
rect 316 215 317 216
rect 315 215 316 216
rect 314 215 315 216
rect 313 215 314 216
rect 312 215 313 216
rect 311 215 312 216
rect 310 215 311 216
rect 309 215 310 216
rect 308 215 309 216
rect 307 215 308 216
rect 306 215 307 216
rect 305 215 306 216
rect 304 215 305 216
rect 303 215 304 216
rect 302 215 303 216
rect 301 215 302 216
rect 300 215 301 216
rect 299 215 300 216
rect 298 215 299 216
rect 297 215 298 216
rect 296 215 297 216
rect 295 215 296 216
rect 294 215 295 216
rect 293 215 294 216
rect 292 215 293 216
rect 291 215 292 216
rect 290 215 291 216
rect 289 215 290 216
rect 288 215 289 216
rect 287 215 288 216
rect 286 215 287 216
rect 285 215 286 216
rect 284 215 285 216
rect 283 215 284 216
rect 282 215 283 216
rect 281 215 282 216
rect 280 215 281 216
rect 279 215 280 216
rect 278 215 279 216
rect 277 215 278 216
rect 276 215 277 216
rect 275 215 276 216
rect 274 215 275 216
rect 273 215 274 216
rect 272 215 273 216
rect 271 215 272 216
rect 270 215 271 216
rect 269 215 270 216
rect 268 215 269 216
rect 267 215 268 216
rect 266 215 267 216
rect 265 215 266 216
rect 264 215 265 216
rect 263 215 264 216
rect 262 215 263 216
rect 261 215 262 216
rect 260 215 261 216
rect 259 215 260 216
rect 258 215 259 216
rect 257 215 258 216
rect 256 215 257 216
rect 255 215 256 216
rect 254 215 255 216
rect 253 215 254 216
rect 252 215 253 216
rect 251 215 252 216
rect 250 215 251 216
rect 249 215 250 216
rect 248 215 249 216
rect 247 215 248 216
rect 246 215 247 216
rect 245 215 246 216
rect 244 215 245 216
rect 243 215 244 216
rect 242 215 243 216
rect 241 215 242 216
rect 240 215 241 216
rect 239 215 240 216
rect 238 215 239 216
rect 237 215 238 216
rect 236 215 237 216
rect 235 215 236 216
rect 234 215 235 216
rect 233 215 234 216
rect 232 215 233 216
rect 231 215 232 216
rect 230 215 231 216
rect 229 215 230 216
rect 228 215 229 216
rect 227 215 228 216
rect 226 215 227 216
rect 225 215 226 216
rect 224 215 225 216
rect 223 215 224 216
rect 222 215 223 216
rect 221 215 222 216
rect 220 215 221 216
rect 219 215 220 216
rect 218 215 219 216
rect 217 215 218 216
rect 216 215 217 216
rect 215 215 216 216
rect 214 215 215 216
rect 213 215 214 216
rect 212 215 213 216
rect 211 215 212 216
rect 210 215 211 216
rect 209 215 210 216
rect 208 215 209 216
rect 207 215 208 216
rect 206 215 207 216
rect 205 215 206 216
rect 204 215 205 216
rect 203 215 204 216
rect 202 215 203 216
rect 201 215 202 216
rect 200 215 201 216
rect 199 215 200 216
rect 198 215 199 216
rect 197 215 198 216
rect 196 215 197 216
rect 195 215 196 216
rect 155 215 156 216
rect 154 215 155 216
rect 153 215 154 216
rect 152 215 153 216
rect 151 215 152 216
rect 150 215 151 216
rect 149 215 150 216
rect 148 215 149 216
rect 147 215 148 216
rect 146 215 147 216
rect 145 215 146 216
rect 144 215 145 216
rect 143 215 144 216
rect 142 215 143 216
rect 141 215 142 216
rect 140 215 141 216
rect 139 215 140 216
rect 138 215 139 216
rect 137 215 138 216
rect 136 215 137 216
rect 135 215 136 216
rect 134 215 135 216
rect 133 215 134 216
rect 132 215 133 216
rect 131 215 132 216
rect 130 215 131 216
rect 129 215 130 216
rect 128 215 129 216
rect 127 215 128 216
rect 126 215 127 216
rect 125 215 126 216
rect 124 215 125 216
rect 123 215 124 216
rect 122 215 123 216
rect 121 215 122 216
rect 120 215 121 216
rect 119 215 120 216
rect 118 215 119 216
rect 117 215 118 216
rect 116 215 117 216
rect 115 215 116 216
rect 114 215 115 216
rect 113 215 114 216
rect 112 215 113 216
rect 111 215 112 216
rect 110 215 111 216
rect 109 215 110 216
rect 108 215 109 216
rect 107 215 108 216
rect 106 215 107 216
rect 105 215 106 216
rect 104 215 105 216
rect 103 215 104 216
rect 102 215 103 216
rect 101 215 102 216
rect 100 215 101 216
rect 99 215 100 216
rect 98 215 99 216
rect 97 215 98 216
rect 96 215 97 216
rect 95 215 96 216
rect 94 215 95 216
rect 93 215 94 216
rect 92 215 93 216
rect 91 215 92 216
rect 90 215 91 216
rect 66 215 67 216
rect 65 215 66 216
rect 64 215 65 216
rect 63 215 64 216
rect 62 215 63 216
rect 61 215 62 216
rect 60 215 61 216
rect 59 215 60 216
rect 58 215 59 216
rect 57 215 58 216
rect 56 215 57 216
rect 55 215 56 216
rect 54 215 55 216
rect 53 215 54 216
rect 52 215 53 216
rect 51 215 52 216
rect 50 215 51 216
rect 49 215 50 216
rect 48 215 49 216
rect 47 215 48 216
rect 46 215 47 216
rect 45 215 46 216
rect 44 215 45 216
rect 43 215 44 216
rect 42 215 43 216
rect 41 215 42 216
rect 40 215 41 216
rect 39 215 40 216
rect 38 215 39 216
rect 37 215 38 216
rect 36 215 37 216
rect 35 215 36 216
rect 34 215 35 216
rect 33 215 34 216
rect 32 215 33 216
rect 31 215 32 216
rect 30 215 31 216
rect 29 215 30 216
rect 28 215 29 216
rect 27 215 28 216
rect 26 215 27 216
rect 25 215 26 216
rect 24 215 25 216
rect 23 215 24 216
rect 22 215 23 216
rect 21 215 22 216
rect 20 215 21 216
rect 19 215 20 216
rect 18 215 19 216
rect 17 215 18 216
rect 16 215 17 216
rect 15 215 16 216
rect 14 215 15 216
rect 13 215 14 216
rect 12 215 13 216
rect 11 215 12 216
rect 10 215 11 216
rect 436 216 437 217
rect 435 216 436 217
rect 434 216 435 217
rect 433 216 434 217
rect 432 216 433 217
rect 431 216 432 217
rect 430 216 431 217
rect 429 216 430 217
rect 428 216 429 217
rect 427 216 428 217
rect 426 216 427 217
rect 425 216 426 217
rect 424 216 425 217
rect 423 216 424 217
rect 422 216 423 217
rect 421 216 422 217
rect 420 216 421 217
rect 419 216 420 217
rect 418 216 419 217
rect 417 216 418 217
rect 416 216 417 217
rect 415 216 416 217
rect 414 216 415 217
rect 413 216 414 217
rect 412 216 413 217
rect 411 216 412 217
rect 410 216 411 217
rect 409 216 410 217
rect 408 216 409 217
rect 407 216 408 217
rect 406 216 407 217
rect 405 216 406 217
rect 404 216 405 217
rect 403 216 404 217
rect 360 216 361 217
rect 359 216 360 217
rect 358 216 359 217
rect 357 216 358 217
rect 356 216 357 217
rect 355 216 356 217
rect 354 216 355 217
rect 353 216 354 217
rect 352 216 353 217
rect 351 216 352 217
rect 350 216 351 217
rect 349 216 350 217
rect 348 216 349 217
rect 347 216 348 217
rect 346 216 347 217
rect 345 216 346 217
rect 344 216 345 217
rect 343 216 344 217
rect 342 216 343 217
rect 341 216 342 217
rect 340 216 341 217
rect 339 216 340 217
rect 338 216 339 217
rect 337 216 338 217
rect 336 216 337 217
rect 335 216 336 217
rect 334 216 335 217
rect 333 216 334 217
rect 332 216 333 217
rect 331 216 332 217
rect 330 216 331 217
rect 329 216 330 217
rect 328 216 329 217
rect 327 216 328 217
rect 326 216 327 217
rect 325 216 326 217
rect 324 216 325 217
rect 323 216 324 217
rect 322 216 323 217
rect 321 216 322 217
rect 320 216 321 217
rect 319 216 320 217
rect 318 216 319 217
rect 317 216 318 217
rect 316 216 317 217
rect 315 216 316 217
rect 314 216 315 217
rect 313 216 314 217
rect 312 216 313 217
rect 311 216 312 217
rect 310 216 311 217
rect 309 216 310 217
rect 308 216 309 217
rect 307 216 308 217
rect 306 216 307 217
rect 305 216 306 217
rect 304 216 305 217
rect 303 216 304 217
rect 302 216 303 217
rect 301 216 302 217
rect 300 216 301 217
rect 299 216 300 217
rect 298 216 299 217
rect 297 216 298 217
rect 296 216 297 217
rect 295 216 296 217
rect 294 216 295 217
rect 293 216 294 217
rect 292 216 293 217
rect 291 216 292 217
rect 290 216 291 217
rect 289 216 290 217
rect 288 216 289 217
rect 287 216 288 217
rect 286 216 287 217
rect 285 216 286 217
rect 284 216 285 217
rect 283 216 284 217
rect 282 216 283 217
rect 281 216 282 217
rect 280 216 281 217
rect 279 216 280 217
rect 278 216 279 217
rect 277 216 278 217
rect 276 216 277 217
rect 275 216 276 217
rect 274 216 275 217
rect 273 216 274 217
rect 272 216 273 217
rect 271 216 272 217
rect 270 216 271 217
rect 269 216 270 217
rect 268 216 269 217
rect 267 216 268 217
rect 266 216 267 217
rect 265 216 266 217
rect 264 216 265 217
rect 263 216 264 217
rect 262 216 263 217
rect 261 216 262 217
rect 260 216 261 217
rect 259 216 260 217
rect 258 216 259 217
rect 257 216 258 217
rect 256 216 257 217
rect 255 216 256 217
rect 254 216 255 217
rect 253 216 254 217
rect 252 216 253 217
rect 251 216 252 217
rect 250 216 251 217
rect 249 216 250 217
rect 248 216 249 217
rect 247 216 248 217
rect 246 216 247 217
rect 245 216 246 217
rect 244 216 245 217
rect 243 216 244 217
rect 242 216 243 217
rect 241 216 242 217
rect 240 216 241 217
rect 239 216 240 217
rect 238 216 239 217
rect 237 216 238 217
rect 236 216 237 217
rect 235 216 236 217
rect 234 216 235 217
rect 233 216 234 217
rect 232 216 233 217
rect 231 216 232 217
rect 230 216 231 217
rect 229 216 230 217
rect 228 216 229 217
rect 227 216 228 217
rect 226 216 227 217
rect 225 216 226 217
rect 224 216 225 217
rect 223 216 224 217
rect 222 216 223 217
rect 221 216 222 217
rect 220 216 221 217
rect 219 216 220 217
rect 218 216 219 217
rect 217 216 218 217
rect 216 216 217 217
rect 215 216 216 217
rect 214 216 215 217
rect 213 216 214 217
rect 212 216 213 217
rect 211 216 212 217
rect 210 216 211 217
rect 209 216 210 217
rect 208 216 209 217
rect 207 216 208 217
rect 206 216 207 217
rect 205 216 206 217
rect 204 216 205 217
rect 203 216 204 217
rect 202 216 203 217
rect 201 216 202 217
rect 200 216 201 217
rect 199 216 200 217
rect 198 216 199 217
rect 197 216 198 217
rect 196 216 197 217
rect 195 216 196 217
rect 194 216 195 217
rect 153 216 154 217
rect 152 216 153 217
rect 151 216 152 217
rect 150 216 151 217
rect 149 216 150 217
rect 148 216 149 217
rect 147 216 148 217
rect 146 216 147 217
rect 145 216 146 217
rect 144 216 145 217
rect 143 216 144 217
rect 142 216 143 217
rect 141 216 142 217
rect 140 216 141 217
rect 139 216 140 217
rect 138 216 139 217
rect 137 216 138 217
rect 136 216 137 217
rect 135 216 136 217
rect 134 216 135 217
rect 133 216 134 217
rect 132 216 133 217
rect 131 216 132 217
rect 130 216 131 217
rect 129 216 130 217
rect 128 216 129 217
rect 127 216 128 217
rect 126 216 127 217
rect 125 216 126 217
rect 124 216 125 217
rect 123 216 124 217
rect 122 216 123 217
rect 121 216 122 217
rect 120 216 121 217
rect 119 216 120 217
rect 118 216 119 217
rect 117 216 118 217
rect 116 216 117 217
rect 115 216 116 217
rect 114 216 115 217
rect 113 216 114 217
rect 112 216 113 217
rect 111 216 112 217
rect 110 216 111 217
rect 109 216 110 217
rect 108 216 109 217
rect 107 216 108 217
rect 106 216 107 217
rect 105 216 106 217
rect 104 216 105 217
rect 103 216 104 217
rect 102 216 103 217
rect 101 216 102 217
rect 100 216 101 217
rect 99 216 100 217
rect 98 216 99 217
rect 97 216 98 217
rect 96 216 97 217
rect 95 216 96 217
rect 94 216 95 217
rect 93 216 94 217
rect 92 216 93 217
rect 67 216 68 217
rect 66 216 67 217
rect 65 216 66 217
rect 64 216 65 217
rect 63 216 64 217
rect 62 216 63 217
rect 61 216 62 217
rect 60 216 61 217
rect 59 216 60 217
rect 58 216 59 217
rect 57 216 58 217
rect 56 216 57 217
rect 55 216 56 217
rect 54 216 55 217
rect 53 216 54 217
rect 52 216 53 217
rect 51 216 52 217
rect 50 216 51 217
rect 49 216 50 217
rect 48 216 49 217
rect 47 216 48 217
rect 46 216 47 217
rect 45 216 46 217
rect 44 216 45 217
rect 43 216 44 217
rect 42 216 43 217
rect 41 216 42 217
rect 40 216 41 217
rect 39 216 40 217
rect 38 216 39 217
rect 37 216 38 217
rect 36 216 37 217
rect 35 216 36 217
rect 34 216 35 217
rect 33 216 34 217
rect 32 216 33 217
rect 31 216 32 217
rect 30 216 31 217
rect 29 216 30 217
rect 28 216 29 217
rect 27 216 28 217
rect 26 216 27 217
rect 25 216 26 217
rect 24 216 25 217
rect 23 216 24 217
rect 22 216 23 217
rect 21 216 22 217
rect 20 216 21 217
rect 19 216 20 217
rect 18 216 19 217
rect 17 216 18 217
rect 16 216 17 217
rect 15 216 16 217
rect 14 216 15 217
rect 13 216 14 217
rect 12 216 13 217
rect 11 216 12 217
rect 10 216 11 217
rect 437 217 438 218
rect 436 217 437 218
rect 435 217 436 218
rect 434 217 435 218
rect 433 217 434 218
rect 432 217 433 218
rect 431 217 432 218
rect 430 217 431 218
rect 429 217 430 218
rect 428 217 429 218
rect 427 217 428 218
rect 426 217 427 218
rect 425 217 426 218
rect 424 217 425 218
rect 423 217 424 218
rect 422 217 423 218
rect 421 217 422 218
rect 420 217 421 218
rect 419 217 420 218
rect 418 217 419 218
rect 417 217 418 218
rect 416 217 417 218
rect 415 217 416 218
rect 414 217 415 218
rect 413 217 414 218
rect 412 217 413 218
rect 411 217 412 218
rect 410 217 411 218
rect 409 217 410 218
rect 408 217 409 218
rect 407 217 408 218
rect 406 217 407 218
rect 405 217 406 218
rect 404 217 405 218
rect 403 217 404 218
rect 402 217 403 218
rect 361 217 362 218
rect 360 217 361 218
rect 359 217 360 218
rect 358 217 359 218
rect 357 217 358 218
rect 356 217 357 218
rect 355 217 356 218
rect 354 217 355 218
rect 353 217 354 218
rect 352 217 353 218
rect 351 217 352 218
rect 350 217 351 218
rect 349 217 350 218
rect 348 217 349 218
rect 347 217 348 218
rect 346 217 347 218
rect 345 217 346 218
rect 344 217 345 218
rect 343 217 344 218
rect 342 217 343 218
rect 341 217 342 218
rect 340 217 341 218
rect 339 217 340 218
rect 338 217 339 218
rect 337 217 338 218
rect 336 217 337 218
rect 335 217 336 218
rect 334 217 335 218
rect 333 217 334 218
rect 313 217 314 218
rect 312 217 313 218
rect 311 217 312 218
rect 310 217 311 218
rect 309 217 310 218
rect 308 217 309 218
rect 307 217 308 218
rect 306 217 307 218
rect 305 217 306 218
rect 304 217 305 218
rect 303 217 304 218
rect 302 217 303 218
rect 301 217 302 218
rect 300 217 301 218
rect 299 217 300 218
rect 298 217 299 218
rect 297 217 298 218
rect 296 217 297 218
rect 295 217 296 218
rect 294 217 295 218
rect 293 217 294 218
rect 292 217 293 218
rect 291 217 292 218
rect 290 217 291 218
rect 289 217 290 218
rect 288 217 289 218
rect 287 217 288 218
rect 286 217 287 218
rect 285 217 286 218
rect 284 217 285 218
rect 283 217 284 218
rect 282 217 283 218
rect 281 217 282 218
rect 280 217 281 218
rect 279 217 280 218
rect 278 217 279 218
rect 277 217 278 218
rect 276 217 277 218
rect 275 217 276 218
rect 274 217 275 218
rect 273 217 274 218
rect 272 217 273 218
rect 271 217 272 218
rect 270 217 271 218
rect 269 217 270 218
rect 268 217 269 218
rect 267 217 268 218
rect 266 217 267 218
rect 265 217 266 218
rect 264 217 265 218
rect 263 217 264 218
rect 262 217 263 218
rect 261 217 262 218
rect 260 217 261 218
rect 259 217 260 218
rect 258 217 259 218
rect 257 217 258 218
rect 256 217 257 218
rect 255 217 256 218
rect 254 217 255 218
rect 253 217 254 218
rect 252 217 253 218
rect 251 217 252 218
rect 250 217 251 218
rect 249 217 250 218
rect 248 217 249 218
rect 247 217 248 218
rect 246 217 247 218
rect 245 217 246 218
rect 244 217 245 218
rect 243 217 244 218
rect 242 217 243 218
rect 241 217 242 218
rect 240 217 241 218
rect 239 217 240 218
rect 238 217 239 218
rect 237 217 238 218
rect 236 217 237 218
rect 235 217 236 218
rect 234 217 235 218
rect 233 217 234 218
rect 232 217 233 218
rect 231 217 232 218
rect 230 217 231 218
rect 229 217 230 218
rect 228 217 229 218
rect 227 217 228 218
rect 226 217 227 218
rect 225 217 226 218
rect 224 217 225 218
rect 223 217 224 218
rect 222 217 223 218
rect 221 217 222 218
rect 220 217 221 218
rect 219 217 220 218
rect 218 217 219 218
rect 217 217 218 218
rect 216 217 217 218
rect 215 217 216 218
rect 214 217 215 218
rect 213 217 214 218
rect 212 217 213 218
rect 211 217 212 218
rect 210 217 211 218
rect 209 217 210 218
rect 208 217 209 218
rect 207 217 208 218
rect 206 217 207 218
rect 205 217 206 218
rect 204 217 205 218
rect 203 217 204 218
rect 202 217 203 218
rect 201 217 202 218
rect 200 217 201 218
rect 199 217 200 218
rect 198 217 199 218
rect 197 217 198 218
rect 196 217 197 218
rect 195 217 196 218
rect 194 217 195 218
rect 193 217 194 218
rect 192 217 193 218
rect 151 217 152 218
rect 150 217 151 218
rect 149 217 150 218
rect 148 217 149 218
rect 147 217 148 218
rect 146 217 147 218
rect 145 217 146 218
rect 144 217 145 218
rect 143 217 144 218
rect 142 217 143 218
rect 141 217 142 218
rect 140 217 141 218
rect 139 217 140 218
rect 138 217 139 218
rect 137 217 138 218
rect 136 217 137 218
rect 135 217 136 218
rect 134 217 135 218
rect 133 217 134 218
rect 132 217 133 218
rect 131 217 132 218
rect 130 217 131 218
rect 129 217 130 218
rect 128 217 129 218
rect 127 217 128 218
rect 126 217 127 218
rect 125 217 126 218
rect 124 217 125 218
rect 123 217 124 218
rect 122 217 123 218
rect 121 217 122 218
rect 120 217 121 218
rect 119 217 120 218
rect 118 217 119 218
rect 117 217 118 218
rect 116 217 117 218
rect 115 217 116 218
rect 114 217 115 218
rect 113 217 114 218
rect 112 217 113 218
rect 111 217 112 218
rect 110 217 111 218
rect 109 217 110 218
rect 108 217 109 218
rect 107 217 108 218
rect 106 217 107 218
rect 105 217 106 218
rect 104 217 105 218
rect 103 217 104 218
rect 102 217 103 218
rect 101 217 102 218
rect 100 217 101 218
rect 99 217 100 218
rect 98 217 99 218
rect 97 217 98 218
rect 96 217 97 218
rect 95 217 96 218
rect 68 217 69 218
rect 67 217 68 218
rect 66 217 67 218
rect 65 217 66 218
rect 64 217 65 218
rect 63 217 64 218
rect 62 217 63 218
rect 61 217 62 218
rect 60 217 61 218
rect 59 217 60 218
rect 58 217 59 218
rect 57 217 58 218
rect 56 217 57 218
rect 55 217 56 218
rect 54 217 55 218
rect 53 217 54 218
rect 52 217 53 218
rect 51 217 52 218
rect 50 217 51 218
rect 49 217 50 218
rect 48 217 49 218
rect 47 217 48 218
rect 46 217 47 218
rect 45 217 46 218
rect 44 217 45 218
rect 43 217 44 218
rect 42 217 43 218
rect 41 217 42 218
rect 40 217 41 218
rect 39 217 40 218
rect 38 217 39 218
rect 37 217 38 218
rect 36 217 37 218
rect 35 217 36 218
rect 34 217 35 218
rect 33 217 34 218
rect 32 217 33 218
rect 31 217 32 218
rect 30 217 31 218
rect 29 217 30 218
rect 28 217 29 218
rect 27 217 28 218
rect 26 217 27 218
rect 25 217 26 218
rect 24 217 25 218
rect 23 217 24 218
rect 22 217 23 218
rect 21 217 22 218
rect 20 217 21 218
rect 19 217 20 218
rect 18 217 19 218
rect 17 217 18 218
rect 16 217 17 218
rect 15 217 16 218
rect 14 217 15 218
rect 13 217 14 218
rect 12 217 13 218
rect 11 217 12 218
rect 10 217 11 218
rect 482 218 483 219
rect 462 218 463 219
rect 438 218 439 219
rect 437 218 438 219
rect 436 218 437 219
rect 435 218 436 219
rect 434 218 435 219
rect 433 218 434 219
rect 432 218 433 219
rect 431 218 432 219
rect 430 218 431 219
rect 429 218 430 219
rect 428 218 429 219
rect 427 218 428 219
rect 426 218 427 219
rect 425 218 426 219
rect 424 218 425 219
rect 423 218 424 219
rect 422 218 423 219
rect 421 218 422 219
rect 420 218 421 219
rect 419 218 420 219
rect 418 218 419 219
rect 417 218 418 219
rect 416 218 417 219
rect 415 218 416 219
rect 414 218 415 219
rect 413 218 414 219
rect 412 218 413 219
rect 411 218 412 219
rect 410 218 411 219
rect 409 218 410 219
rect 408 218 409 219
rect 407 218 408 219
rect 406 218 407 219
rect 405 218 406 219
rect 404 218 405 219
rect 403 218 404 219
rect 402 218 403 219
rect 401 218 402 219
rect 361 218 362 219
rect 360 218 361 219
rect 359 218 360 219
rect 358 218 359 219
rect 357 218 358 219
rect 356 218 357 219
rect 355 218 356 219
rect 354 218 355 219
rect 353 218 354 219
rect 352 218 353 219
rect 351 218 352 219
rect 350 218 351 219
rect 349 218 350 219
rect 348 218 349 219
rect 347 218 348 219
rect 346 218 347 219
rect 345 218 346 219
rect 344 218 345 219
rect 343 218 344 219
rect 342 218 343 219
rect 341 218 342 219
rect 340 218 341 219
rect 339 218 340 219
rect 307 218 308 219
rect 306 218 307 219
rect 305 218 306 219
rect 304 218 305 219
rect 303 218 304 219
rect 302 218 303 219
rect 301 218 302 219
rect 300 218 301 219
rect 299 218 300 219
rect 298 218 299 219
rect 297 218 298 219
rect 296 218 297 219
rect 295 218 296 219
rect 294 218 295 219
rect 293 218 294 219
rect 292 218 293 219
rect 291 218 292 219
rect 290 218 291 219
rect 289 218 290 219
rect 288 218 289 219
rect 287 218 288 219
rect 286 218 287 219
rect 285 218 286 219
rect 284 218 285 219
rect 283 218 284 219
rect 282 218 283 219
rect 281 218 282 219
rect 280 218 281 219
rect 279 218 280 219
rect 278 218 279 219
rect 277 218 278 219
rect 276 218 277 219
rect 275 218 276 219
rect 274 218 275 219
rect 273 218 274 219
rect 272 218 273 219
rect 271 218 272 219
rect 270 218 271 219
rect 269 218 270 219
rect 268 218 269 219
rect 267 218 268 219
rect 266 218 267 219
rect 265 218 266 219
rect 264 218 265 219
rect 263 218 264 219
rect 262 218 263 219
rect 261 218 262 219
rect 260 218 261 219
rect 259 218 260 219
rect 258 218 259 219
rect 257 218 258 219
rect 256 218 257 219
rect 255 218 256 219
rect 254 218 255 219
rect 253 218 254 219
rect 252 218 253 219
rect 251 218 252 219
rect 250 218 251 219
rect 249 218 250 219
rect 248 218 249 219
rect 247 218 248 219
rect 246 218 247 219
rect 245 218 246 219
rect 244 218 245 219
rect 243 218 244 219
rect 242 218 243 219
rect 241 218 242 219
rect 240 218 241 219
rect 239 218 240 219
rect 238 218 239 219
rect 237 218 238 219
rect 236 218 237 219
rect 235 218 236 219
rect 234 218 235 219
rect 233 218 234 219
rect 232 218 233 219
rect 231 218 232 219
rect 230 218 231 219
rect 229 218 230 219
rect 228 218 229 219
rect 227 218 228 219
rect 226 218 227 219
rect 225 218 226 219
rect 224 218 225 219
rect 223 218 224 219
rect 222 218 223 219
rect 221 218 222 219
rect 220 218 221 219
rect 219 218 220 219
rect 218 218 219 219
rect 217 218 218 219
rect 216 218 217 219
rect 215 218 216 219
rect 214 218 215 219
rect 213 218 214 219
rect 212 218 213 219
rect 211 218 212 219
rect 210 218 211 219
rect 209 218 210 219
rect 208 218 209 219
rect 207 218 208 219
rect 206 218 207 219
rect 205 218 206 219
rect 204 218 205 219
rect 203 218 204 219
rect 202 218 203 219
rect 201 218 202 219
rect 200 218 201 219
rect 199 218 200 219
rect 198 218 199 219
rect 197 218 198 219
rect 196 218 197 219
rect 195 218 196 219
rect 194 218 195 219
rect 193 218 194 219
rect 192 218 193 219
rect 191 218 192 219
rect 190 218 191 219
rect 150 218 151 219
rect 149 218 150 219
rect 148 218 149 219
rect 147 218 148 219
rect 146 218 147 219
rect 145 218 146 219
rect 144 218 145 219
rect 143 218 144 219
rect 142 218 143 219
rect 141 218 142 219
rect 140 218 141 219
rect 139 218 140 219
rect 138 218 139 219
rect 137 218 138 219
rect 136 218 137 219
rect 135 218 136 219
rect 134 218 135 219
rect 133 218 134 219
rect 132 218 133 219
rect 131 218 132 219
rect 130 218 131 219
rect 129 218 130 219
rect 128 218 129 219
rect 127 218 128 219
rect 126 218 127 219
rect 125 218 126 219
rect 124 218 125 219
rect 123 218 124 219
rect 122 218 123 219
rect 121 218 122 219
rect 120 218 121 219
rect 119 218 120 219
rect 118 218 119 219
rect 117 218 118 219
rect 116 218 117 219
rect 115 218 116 219
rect 114 218 115 219
rect 113 218 114 219
rect 112 218 113 219
rect 111 218 112 219
rect 110 218 111 219
rect 109 218 110 219
rect 108 218 109 219
rect 107 218 108 219
rect 106 218 107 219
rect 105 218 106 219
rect 104 218 105 219
rect 103 218 104 219
rect 102 218 103 219
rect 101 218 102 219
rect 100 218 101 219
rect 99 218 100 219
rect 98 218 99 219
rect 97 218 98 219
rect 69 218 70 219
rect 68 218 69 219
rect 67 218 68 219
rect 66 218 67 219
rect 65 218 66 219
rect 64 218 65 219
rect 63 218 64 219
rect 62 218 63 219
rect 61 218 62 219
rect 60 218 61 219
rect 59 218 60 219
rect 58 218 59 219
rect 57 218 58 219
rect 56 218 57 219
rect 55 218 56 219
rect 54 218 55 219
rect 53 218 54 219
rect 52 218 53 219
rect 51 218 52 219
rect 50 218 51 219
rect 49 218 50 219
rect 48 218 49 219
rect 47 218 48 219
rect 46 218 47 219
rect 45 218 46 219
rect 44 218 45 219
rect 43 218 44 219
rect 42 218 43 219
rect 41 218 42 219
rect 40 218 41 219
rect 39 218 40 219
rect 38 218 39 219
rect 37 218 38 219
rect 36 218 37 219
rect 35 218 36 219
rect 34 218 35 219
rect 33 218 34 219
rect 32 218 33 219
rect 31 218 32 219
rect 30 218 31 219
rect 29 218 30 219
rect 28 218 29 219
rect 27 218 28 219
rect 26 218 27 219
rect 25 218 26 219
rect 24 218 25 219
rect 23 218 24 219
rect 22 218 23 219
rect 21 218 22 219
rect 20 218 21 219
rect 19 218 20 219
rect 18 218 19 219
rect 17 218 18 219
rect 16 218 17 219
rect 15 218 16 219
rect 14 218 15 219
rect 13 218 14 219
rect 12 218 13 219
rect 11 218 12 219
rect 10 218 11 219
rect 482 219 483 220
rect 462 219 463 220
rect 438 219 439 220
rect 437 219 438 220
rect 436 219 437 220
rect 435 219 436 220
rect 434 219 435 220
rect 433 219 434 220
rect 432 219 433 220
rect 431 219 432 220
rect 430 219 431 220
rect 429 219 430 220
rect 428 219 429 220
rect 427 219 428 220
rect 426 219 427 220
rect 425 219 426 220
rect 424 219 425 220
rect 423 219 424 220
rect 422 219 423 220
rect 421 219 422 220
rect 420 219 421 220
rect 419 219 420 220
rect 418 219 419 220
rect 417 219 418 220
rect 416 219 417 220
rect 415 219 416 220
rect 414 219 415 220
rect 413 219 414 220
rect 412 219 413 220
rect 411 219 412 220
rect 410 219 411 220
rect 409 219 410 220
rect 408 219 409 220
rect 407 219 408 220
rect 406 219 407 220
rect 405 219 406 220
rect 404 219 405 220
rect 403 219 404 220
rect 402 219 403 220
rect 401 219 402 220
rect 362 219 363 220
rect 361 219 362 220
rect 360 219 361 220
rect 359 219 360 220
rect 358 219 359 220
rect 357 219 358 220
rect 356 219 357 220
rect 355 219 356 220
rect 354 219 355 220
rect 353 219 354 220
rect 352 219 353 220
rect 351 219 352 220
rect 350 219 351 220
rect 349 219 350 220
rect 348 219 349 220
rect 347 219 348 220
rect 346 219 347 220
rect 345 219 346 220
rect 344 219 345 220
rect 303 219 304 220
rect 302 219 303 220
rect 301 219 302 220
rect 300 219 301 220
rect 299 219 300 220
rect 298 219 299 220
rect 297 219 298 220
rect 296 219 297 220
rect 295 219 296 220
rect 294 219 295 220
rect 293 219 294 220
rect 292 219 293 220
rect 291 219 292 220
rect 290 219 291 220
rect 289 219 290 220
rect 288 219 289 220
rect 287 219 288 220
rect 286 219 287 220
rect 285 219 286 220
rect 284 219 285 220
rect 283 219 284 220
rect 282 219 283 220
rect 281 219 282 220
rect 280 219 281 220
rect 279 219 280 220
rect 278 219 279 220
rect 277 219 278 220
rect 276 219 277 220
rect 275 219 276 220
rect 274 219 275 220
rect 273 219 274 220
rect 272 219 273 220
rect 271 219 272 220
rect 270 219 271 220
rect 269 219 270 220
rect 268 219 269 220
rect 267 219 268 220
rect 266 219 267 220
rect 265 219 266 220
rect 264 219 265 220
rect 263 219 264 220
rect 262 219 263 220
rect 261 219 262 220
rect 260 219 261 220
rect 259 219 260 220
rect 258 219 259 220
rect 257 219 258 220
rect 256 219 257 220
rect 255 219 256 220
rect 254 219 255 220
rect 253 219 254 220
rect 252 219 253 220
rect 251 219 252 220
rect 250 219 251 220
rect 249 219 250 220
rect 248 219 249 220
rect 247 219 248 220
rect 246 219 247 220
rect 245 219 246 220
rect 244 219 245 220
rect 243 219 244 220
rect 242 219 243 220
rect 241 219 242 220
rect 240 219 241 220
rect 239 219 240 220
rect 238 219 239 220
rect 237 219 238 220
rect 236 219 237 220
rect 235 219 236 220
rect 234 219 235 220
rect 233 219 234 220
rect 232 219 233 220
rect 231 219 232 220
rect 230 219 231 220
rect 229 219 230 220
rect 228 219 229 220
rect 227 219 228 220
rect 226 219 227 220
rect 225 219 226 220
rect 224 219 225 220
rect 223 219 224 220
rect 222 219 223 220
rect 221 219 222 220
rect 220 219 221 220
rect 219 219 220 220
rect 218 219 219 220
rect 217 219 218 220
rect 216 219 217 220
rect 215 219 216 220
rect 214 219 215 220
rect 213 219 214 220
rect 212 219 213 220
rect 211 219 212 220
rect 210 219 211 220
rect 209 219 210 220
rect 208 219 209 220
rect 207 219 208 220
rect 206 219 207 220
rect 205 219 206 220
rect 204 219 205 220
rect 203 219 204 220
rect 202 219 203 220
rect 201 219 202 220
rect 200 219 201 220
rect 199 219 200 220
rect 198 219 199 220
rect 197 219 198 220
rect 196 219 197 220
rect 195 219 196 220
rect 194 219 195 220
rect 193 219 194 220
rect 192 219 193 220
rect 191 219 192 220
rect 190 219 191 220
rect 189 219 190 220
rect 188 219 189 220
rect 149 219 150 220
rect 148 219 149 220
rect 147 219 148 220
rect 146 219 147 220
rect 145 219 146 220
rect 144 219 145 220
rect 143 219 144 220
rect 142 219 143 220
rect 141 219 142 220
rect 140 219 141 220
rect 139 219 140 220
rect 138 219 139 220
rect 137 219 138 220
rect 136 219 137 220
rect 135 219 136 220
rect 134 219 135 220
rect 133 219 134 220
rect 132 219 133 220
rect 131 219 132 220
rect 130 219 131 220
rect 129 219 130 220
rect 128 219 129 220
rect 127 219 128 220
rect 126 219 127 220
rect 125 219 126 220
rect 124 219 125 220
rect 123 219 124 220
rect 122 219 123 220
rect 121 219 122 220
rect 120 219 121 220
rect 119 219 120 220
rect 118 219 119 220
rect 117 219 118 220
rect 116 219 117 220
rect 115 219 116 220
rect 114 219 115 220
rect 113 219 114 220
rect 112 219 113 220
rect 111 219 112 220
rect 110 219 111 220
rect 109 219 110 220
rect 108 219 109 220
rect 107 219 108 220
rect 106 219 107 220
rect 105 219 106 220
rect 104 219 105 220
rect 103 219 104 220
rect 102 219 103 220
rect 101 219 102 220
rect 100 219 101 220
rect 99 219 100 220
rect 70 219 71 220
rect 69 219 70 220
rect 68 219 69 220
rect 67 219 68 220
rect 66 219 67 220
rect 65 219 66 220
rect 64 219 65 220
rect 63 219 64 220
rect 62 219 63 220
rect 61 219 62 220
rect 60 219 61 220
rect 59 219 60 220
rect 58 219 59 220
rect 57 219 58 220
rect 56 219 57 220
rect 55 219 56 220
rect 54 219 55 220
rect 53 219 54 220
rect 52 219 53 220
rect 51 219 52 220
rect 50 219 51 220
rect 49 219 50 220
rect 48 219 49 220
rect 47 219 48 220
rect 46 219 47 220
rect 45 219 46 220
rect 44 219 45 220
rect 43 219 44 220
rect 42 219 43 220
rect 41 219 42 220
rect 40 219 41 220
rect 39 219 40 220
rect 38 219 39 220
rect 37 219 38 220
rect 36 219 37 220
rect 35 219 36 220
rect 34 219 35 220
rect 33 219 34 220
rect 32 219 33 220
rect 31 219 32 220
rect 30 219 31 220
rect 29 219 30 220
rect 28 219 29 220
rect 27 219 28 220
rect 26 219 27 220
rect 25 219 26 220
rect 24 219 25 220
rect 23 219 24 220
rect 22 219 23 220
rect 21 219 22 220
rect 20 219 21 220
rect 19 219 20 220
rect 18 219 19 220
rect 17 219 18 220
rect 16 219 17 220
rect 15 219 16 220
rect 14 219 15 220
rect 13 219 14 220
rect 12 219 13 220
rect 11 219 12 220
rect 10 219 11 220
rect 9 219 10 220
rect 482 220 483 221
rect 481 220 482 221
rect 480 220 481 221
rect 464 220 465 221
rect 463 220 464 221
rect 462 220 463 221
rect 439 220 440 221
rect 438 220 439 221
rect 437 220 438 221
rect 436 220 437 221
rect 435 220 436 221
rect 434 220 435 221
rect 433 220 434 221
rect 432 220 433 221
rect 431 220 432 221
rect 430 220 431 221
rect 429 220 430 221
rect 428 220 429 221
rect 427 220 428 221
rect 426 220 427 221
rect 425 220 426 221
rect 412 220 413 221
rect 411 220 412 221
rect 410 220 411 221
rect 409 220 410 221
rect 408 220 409 221
rect 407 220 408 221
rect 406 220 407 221
rect 405 220 406 221
rect 404 220 405 221
rect 403 220 404 221
rect 402 220 403 221
rect 401 220 402 221
rect 400 220 401 221
rect 362 220 363 221
rect 361 220 362 221
rect 360 220 361 221
rect 359 220 360 221
rect 358 220 359 221
rect 357 220 358 221
rect 356 220 357 221
rect 355 220 356 221
rect 354 220 355 221
rect 353 220 354 221
rect 352 220 353 221
rect 351 220 352 221
rect 350 220 351 221
rect 349 220 350 221
rect 348 220 349 221
rect 300 220 301 221
rect 299 220 300 221
rect 298 220 299 221
rect 297 220 298 221
rect 296 220 297 221
rect 295 220 296 221
rect 294 220 295 221
rect 293 220 294 221
rect 292 220 293 221
rect 291 220 292 221
rect 290 220 291 221
rect 289 220 290 221
rect 288 220 289 221
rect 287 220 288 221
rect 286 220 287 221
rect 285 220 286 221
rect 284 220 285 221
rect 283 220 284 221
rect 282 220 283 221
rect 281 220 282 221
rect 280 220 281 221
rect 279 220 280 221
rect 278 220 279 221
rect 277 220 278 221
rect 276 220 277 221
rect 275 220 276 221
rect 274 220 275 221
rect 273 220 274 221
rect 272 220 273 221
rect 271 220 272 221
rect 270 220 271 221
rect 269 220 270 221
rect 268 220 269 221
rect 267 220 268 221
rect 266 220 267 221
rect 265 220 266 221
rect 264 220 265 221
rect 263 220 264 221
rect 262 220 263 221
rect 261 220 262 221
rect 260 220 261 221
rect 259 220 260 221
rect 258 220 259 221
rect 257 220 258 221
rect 256 220 257 221
rect 255 220 256 221
rect 254 220 255 221
rect 253 220 254 221
rect 252 220 253 221
rect 251 220 252 221
rect 250 220 251 221
rect 249 220 250 221
rect 248 220 249 221
rect 247 220 248 221
rect 246 220 247 221
rect 245 220 246 221
rect 244 220 245 221
rect 243 220 244 221
rect 242 220 243 221
rect 241 220 242 221
rect 240 220 241 221
rect 239 220 240 221
rect 238 220 239 221
rect 237 220 238 221
rect 236 220 237 221
rect 235 220 236 221
rect 234 220 235 221
rect 233 220 234 221
rect 232 220 233 221
rect 231 220 232 221
rect 230 220 231 221
rect 229 220 230 221
rect 228 220 229 221
rect 227 220 228 221
rect 226 220 227 221
rect 225 220 226 221
rect 224 220 225 221
rect 223 220 224 221
rect 222 220 223 221
rect 221 220 222 221
rect 220 220 221 221
rect 219 220 220 221
rect 218 220 219 221
rect 217 220 218 221
rect 216 220 217 221
rect 215 220 216 221
rect 214 220 215 221
rect 213 220 214 221
rect 212 220 213 221
rect 211 220 212 221
rect 210 220 211 221
rect 209 220 210 221
rect 208 220 209 221
rect 207 220 208 221
rect 206 220 207 221
rect 205 220 206 221
rect 204 220 205 221
rect 203 220 204 221
rect 202 220 203 221
rect 201 220 202 221
rect 200 220 201 221
rect 199 220 200 221
rect 198 220 199 221
rect 197 220 198 221
rect 196 220 197 221
rect 195 220 196 221
rect 194 220 195 221
rect 193 220 194 221
rect 192 220 193 221
rect 191 220 192 221
rect 190 220 191 221
rect 189 220 190 221
rect 188 220 189 221
rect 187 220 188 221
rect 186 220 187 221
rect 185 220 186 221
rect 148 220 149 221
rect 147 220 148 221
rect 146 220 147 221
rect 145 220 146 221
rect 144 220 145 221
rect 143 220 144 221
rect 142 220 143 221
rect 141 220 142 221
rect 140 220 141 221
rect 139 220 140 221
rect 138 220 139 221
rect 137 220 138 221
rect 136 220 137 221
rect 135 220 136 221
rect 134 220 135 221
rect 133 220 134 221
rect 132 220 133 221
rect 131 220 132 221
rect 130 220 131 221
rect 129 220 130 221
rect 128 220 129 221
rect 127 220 128 221
rect 126 220 127 221
rect 125 220 126 221
rect 124 220 125 221
rect 123 220 124 221
rect 122 220 123 221
rect 121 220 122 221
rect 120 220 121 221
rect 119 220 120 221
rect 118 220 119 221
rect 117 220 118 221
rect 116 220 117 221
rect 115 220 116 221
rect 114 220 115 221
rect 113 220 114 221
rect 112 220 113 221
rect 111 220 112 221
rect 110 220 111 221
rect 109 220 110 221
rect 108 220 109 221
rect 107 220 108 221
rect 106 220 107 221
rect 105 220 106 221
rect 104 220 105 221
rect 103 220 104 221
rect 102 220 103 221
rect 101 220 102 221
rect 71 220 72 221
rect 70 220 71 221
rect 69 220 70 221
rect 68 220 69 221
rect 67 220 68 221
rect 66 220 67 221
rect 65 220 66 221
rect 64 220 65 221
rect 63 220 64 221
rect 62 220 63 221
rect 61 220 62 221
rect 60 220 61 221
rect 59 220 60 221
rect 58 220 59 221
rect 57 220 58 221
rect 56 220 57 221
rect 55 220 56 221
rect 54 220 55 221
rect 53 220 54 221
rect 52 220 53 221
rect 51 220 52 221
rect 50 220 51 221
rect 49 220 50 221
rect 48 220 49 221
rect 47 220 48 221
rect 46 220 47 221
rect 45 220 46 221
rect 44 220 45 221
rect 43 220 44 221
rect 42 220 43 221
rect 41 220 42 221
rect 40 220 41 221
rect 39 220 40 221
rect 38 220 39 221
rect 37 220 38 221
rect 36 220 37 221
rect 35 220 36 221
rect 34 220 35 221
rect 33 220 34 221
rect 32 220 33 221
rect 31 220 32 221
rect 30 220 31 221
rect 29 220 30 221
rect 28 220 29 221
rect 27 220 28 221
rect 26 220 27 221
rect 25 220 26 221
rect 24 220 25 221
rect 23 220 24 221
rect 22 220 23 221
rect 21 220 22 221
rect 20 220 21 221
rect 19 220 20 221
rect 18 220 19 221
rect 17 220 18 221
rect 16 220 17 221
rect 15 220 16 221
rect 14 220 15 221
rect 13 220 14 221
rect 12 220 13 221
rect 11 220 12 221
rect 10 220 11 221
rect 9 220 10 221
rect 482 221 483 222
rect 481 221 482 222
rect 480 221 481 222
rect 479 221 480 222
rect 478 221 479 222
rect 477 221 478 222
rect 476 221 477 222
rect 475 221 476 222
rect 474 221 475 222
rect 473 221 474 222
rect 472 221 473 222
rect 471 221 472 222
rect 470 221 471 222
rect 469 221 470 222
rect 468 221 469 222
rect 467 221 468 222
rect 466 221 467 222
rect 465 221 466 222
rect 464 221 465 222
rect 463 221 464 222
rect 462 221 463 222
rect 439 221 440 222
rect 438 221 439 222
rect 437 221 438 222
rect 436 221 437 222
rect 435 221 436 222
rect 434 221 435 222
rect 433 221 434 222
rect 432 221 433 222
rect 431 221 432 222
rect 430 221 431 222
rect 429 221 430 222
rect 408 221 409 222
rect 407 221 408 222
rect 406 221 407 222
rect 405 221 406 222
rect 404 221 405 222
rect 403 221 404 222
rect 402 221 403 222
rect 401 221 402 222
rect 400 221 401 222
rect 399 221 400 222
rect 363 221 364 222
rect 362 221 363 222
rect 361 221 362 222
rect 360 221 361 222
rect 359 221 360 222
rect 358 221 359 222
rect 357 221 358 222
rect 356 221 357 222
rect 355 221 356 222
rect 354 221 355 222
rect 353 221 354 222
rect 352 221 353 222
rect 351 221 352 222
rect 297 221 298 222
rect 296 221 297 222
rect 295 221 296 222
rect 294 221 295 222
rect 293 221 294 222
rect 292 221 293 222
rect 291 221 292 222
rect 290 221 291 222
rect 289 221 290 222
rect 288 221 289 222
rect 287 221 288 222
rect 286 221 287 222
rect 285 221 286 222
rect 284 221 285 222
rect 283 221 284 222
rect 282 221 283 222
rect 281 221 282 222
rect 280 221 281 222
rect 279 221 280 222
rect 278 221 279 222
rect 277 221 278 222
rect 276 221 277 222
rect 275 221 276 222
rect 274 221 275 222
rect 273 221 274 222
rect 272 221 273 222
rect 271 221 272 222
rect 270 221 271 222
rect 269 221 270 222
rect 268 221 269 222
rect 267 221 268 222
rect 266 221 267 222
rect 265 221 266 222
rect 264 221 265 222
rect 263 221 264 222
rect 262 221 263 222
rect 261 221 262 222
rect 260 221 261 222
rect 259 221 260 222
rect 258 221 259 222
rect 257 221 258 222
rect 256 221 257 222
rect 255 221 256 222
rect 254 221 255 222
rect 253 221 254 222
rect 252 221 253 222
rect 251 221 252 222
rect 250 221 251 222
rect 249 221 250 222
rect 248 221 249 222
rect 247 221 248 222
rect 246 221 247 222
rect 245 221 246 222
rect 244 221 245 222
rect 243 221 244 222
rect 242 221 243 222
rect 241 221 242 222
rect 240 221 241 222
rect 239 221 240 222
rect 238 221 239 222
rect 237 221 238 222
rect 236 221 237 222
rect 235 221 236 222
rect 234 221 235 222
rect 233 221 234 222
rect 232 221 233 222
rect 231 221 232 222
rect 230 221 231 222
rect 229 221 230 222
rect 228 221 229 222
rect 227 221 228 222
rect 226 221 227 222
rect 225 221 226 222
rect 224 221 225 222
rect 223 221 224 222
rect 222 221 223 222
rect 221 221 222 222
rect 220 221 221 222
rect 219 221 220 222
rect 218 221 219 222
rect 217 221 218 222
rect 216 221 217 222
rect 215 221 216 222
rect 214 221 215 222
rect 213 221 214 222
rect 212 221 213 222
rect 211 221 212 222
rect 210 221 211 222
rect 209 221 210 222
rect 208 221 209 222
rect 207 221 208 222
rect 206 221 207 222
rect 205 221 206 222
rect 204 221 205 222
rect 203 221 204 222
rect 202 221 203 222
rect 201 221 202 222
rect 200 221 201 222
rect 199 221 200 222
rect 198 221 199 222
rect 197 221 198 222
rect 196 221 197 222
rect 195 221 196 222
rect 194 221 195 222
rect 193 221 194 222
rect 192 221 193 222
rect 191 221 192 222
rect 190 221 191 222
rect 189 221 190 222
rect 188 221 189 222
rect 187 221 188 222
rect 186 221 187 222
rect 185 221 186 222
rect 184 221 185 222
rect 183 221 184 222
rect 147 221 148 222
rect 146 221 147 222
rect 145 221 146 222
rect 144 221 145 222
rect 143 221 144 222
rect 142 221 143 222
rect 141 221 142 222
rect 140 221 141 222
rect 139 221 140 222
rect 138 221 139 222
rect 137 221 138 222
rect 136 221 137 222
rect 135 221 136 222
rect 134 221 135 222
rect 133 221 134 222
rect 132 221 133 222
rect 131 221 132 222
rect 130 221 131 222
rect 129 221 130 222
rect 128 221 129 222
rect 127 221 128 222
rect 126 221 127 222
rect 125 221 126 222
rect 124 221 125 222
rect 123 221 124 222
rect 122 221 123 222
rect 121 221 122 222
rect 120 221 121 222
rect 119 221 120 222
rect 118 221 119 222
rect 117 221 118 222
rect 116 221 117 222
rect 115 221 116 222
rect 114 221 115 222
rect 113 221 114 222
rect 112 221 113 222
rect 111 221 112 222
rect 110 221 111 222
rect 109 221 110 222
rect 108 221 109 222
rect 107 221 108 222
rect 106 221 107 222
rect 105 221 106 222
rect 104 221 105 222
rect 103 221 104 222
rect 72 221 73 222
rect 71 221 72 222
rect 70 221 71 222
rect 69 221 70 222
rect 68 221 69 222
rect 67 221 68 222
rect 66 221 67 222
rect 65 221 66 222
rect 64 221 65 222
rect 63 221 64 222
rect 62 221 63 222
rect 61 221 62 222
rect 60 221 61 222
rect 59 221 60 222
rect 58 221 59 222
rect 57 221 58 222
rect 56 221 57 222
rect 55 221 56 222
rect 54 221 55 222
rect 53 221 54 222
rect 52 221 53 222
rect 51 221 52 222
rect 50 221 51 222
rect 49 221 50 222
rect 48 221 49 222
rect 47 221 48 222
rect 46 221 47 222
rect 45 221 46 222
rect 44 221 45 222
rect 43 221 44 222
rect 42 221 43 222
rect 41 221 42 222
rect 40 221 41 222
rect 39 221 40 222
rect 38 221 39 222
rect 37 221 38 222
rect 36 221 37 222
rect 35 221 36 222
rect 34 221 35 222
rect 33 221 34 222
rect 32 221 33 222
rect 31 221 32 222
rect 30 221 31 222
rect 29 221 30 222
rect 28 221 29 222
rect 27 221 28 222
rect 26 221 27 222
rect 25 221 26 222
rect 24 221 25 222
rect 23 221 24 222
rect 22 221 23 222
rect 21 221 22 222
rect 20 221 21 222
rect 19 221 20 222
rect 18 221 19 222
rect 17 221 18 222
rect 16 221 17 222
rect 15 221 16 222
rect 14 221 15 222
rect 13 221 14 222
rect 12 221 13 222
rect 11 221 12 222
rect 10 221 11 222
rect 9 221 10 222
rect 482 222 483 223
rect 481 222 482 223
rect 480 222 481 223
rect 479 222 480 223
rect 478 222 479 223
rect 477 222 478 223
rect 476 222 477 223
rect 475 222 476 223
rect 474 222 475 223
rect 473 222 474 223
rect 472 222 473 223
rect 471 222 472 223
rect 470 222 471 223
rect 469 222 470 223
rect 468 222 469 223
rect 467 222 468 223
rect 466 222 467 223
rect 465 222 466 223
rect 464 222 465 223
rect 463 222 464 223
rect 462 222 463 223
rect 440 222 441 223
rect 439 222 440 223
rect 438 222 439 223
rect 437 222 438 223
rect 436 222 437 223
rect 435 222 436 223
rect 434 222 435 223
rect 433 222 434 223
rect 432 222 433 223
rect 431 222 432 223
rect 406 222 407 223
rect 405 222 406 223
rect 404 222 405 223
rect 403 222 404 223
rect 402 222 403 223
rect 401 222 402 223
rect 400 222 401 223
rect 399 222 400 223
rect 363 222 364 223
rect 362 222 363 223
rect 361 222 362 223
rect 360 222 361 223
rect 359 222 360 223
rect 358 222 359 223
rect 357 222 358 223
rect 356 222 357 223
rect 355 222 356 223
rect 354 222 355 223
rect 295 222 296 223
rect 294 222 295 223
rect 293 222 294 223
rect 292 222 293 223
rect 291 222 292 223
rect 290 222 291 223
rect 289 222 290 223
rect 288 222 289 223
rect 287 222 288 223
rect 286 222 287 223
rect 285 222 286 223
rect 284 222 285 223
rect 283 222 284 223
rect 282 222 283 223
rect 281 222 282 223
rect 280 222 281 223
rect 279 222 280 223
rect 278 222 279 223
rect 277 222 278 223
rect 276 222 277 223
rect 275 222 276 223
rect 274 222 275 223
rect 273 222 274 223
rect 272 222 273 223
rect 271 222 272 223
rect 270 222 271 223
rect 269 222 270 223
rect 268 222 269 223
rect 267 222 268 223
rect 266 222 267 223
rect 265 222 266 223
rect 264 222 265 223
rect 263 222 264 223
rect 262 222 263 223
rect 261 222 262 223
rect 260 222 261 223
rect 259 222 260 223
rect 258 222 259 223
rect 257 222 258 223
rect 256 222 257 223
rect 255 222 256 223
rect 254 222 255 223
rect 253 222 254 223
rect 252 222 253 223
rect 251 222 252 223
rect 250 222 251 223
rect 249 222 250 223
rect 248 222 249 223
rect 247 222 248 223
rect 246 222 247 223
rect 245 222 246 223
rect 244 222 245 223
rect 243 222 244 223
rect 242 222 243 223
rect 241 222 242 223
rect 240 222 241 223
rect 239 222 240 223
rect 238 222 239 223
rect 237 222 238 223
rect 236 222 237 223
rect 235 222 236 223
rect 234 222 235 223
rect 233 222 234 223
rect 232 222 233 223
rect 231 222 232 223
rect 230 222 231 223
rect 229 222 230 223
rect 228 222 229 223
rect 227 222 228 223
rect 226 222 227 223
rect 225 222 226 223
rect 224 222 225 223
rect 223 222 224 223
rect 222 222 223 223
rect 221 222 222 223
rect 220 222 221 223
rect 219 222 220 223
rect 218 222 219 223
rect 217 222 218 223
rect 216 222 217 223
rect 215 222 216 223
rect 214 222 215 223
rect 213 222 214 223
rect 212 222 213 223
rect 211 222 212 223
rect 210 222 211 223
rect 209 222 210 223
rect 208 222 209 223
rect 207 222 208 223
rect 206 222 207 223
rect 205 222 206 223
rect 204 222 205 223
rect 203 222 204 223
rect 202 222 203 223
rect 201 222 202 223
rect 200 222 201 223
rect 199 222 200 223
rect 198 222 199 223
rect 197 222 198 223
rect 196 222 197 223
rect 195 222 196 223
rect 194 222 195 223
rect 193 222 194 223
rect 192 222 193 223
rect 191 222 192 223
rect 190 222 191 223
rect 189 222 190 223
rect 188 222 189 223
rect 187 222 188 223
rect 186 222 187 223
rect 185 222 186 223
rect 184 222 185 223
rect 183 222 184 223
rect 182 222 183 223
rect 181 222 182 223
rect 147 222 148 223
rect 146 222 147 223
rect 145 222 146 223
rect 144 222 145 223
rect 143 222 144 223
rect 142 222 143 223
rect 141 222 142 223
rect 140 222 141 223
rect 139 222 140 223
rect 138 222 139 223
rect 137 222 138 223
rect 136 222 137 223
rect 135 222 136 223
rect 134 222 135 223
rect 133 222 134 223
rect 132 222 133 223
rect 131 222 132 223
rect 130 222 131 223
rect 129 222 130 223
rect 128 222 129 223
rect 127 222 128 223
rect 126 222 127 223
rect 125 222 126 223
rect 124 222 125 223
rect 123 222 124 223
rect 122 222 123 223
rect 121 222 122 223
rect 120 222 121 223
rect 119 222 120 223
rect 118 222 119 223
rect 117 222 118 223
rect 116 222 117 223
rect 115 222 116 223
rect 114 222 115 223
rect 113 222 114 223
rect 112 222 113 223
rect 111 222 112 223
rect 110 222 111 223
rect 109 222 110 223
rect 108 222 109 223
rect 107 222 108 223
rect 106 222 107 223
rect 105 222 106 223
rect 73 222 74 223
rect 72 222 73 223
rect 71 222 72 223
rect 70 222 71 223
rect 69 222 70 223
rect 68 222 69 223
rect 67 222 68 223
rect 66 222 67 223
rect 65 222 66 223
rect 64 222 65 223
rect 63 222 64 223
rect 62 222 63 223
rect 61 222 62 223
rect 60 222 61 223
rect 59 222 60 223
rect 58 222 59 223
rect 57 222 58 223
rect 56 222 57 223
rect 55 222 56 223
rect 54 222 55 223
rect 53 222 54 223
rect 52 222 53 223
rect 51 222 52 223
rect 50 222 51 223
rect 49 222 50 223
rect 48 222 49 223
rect 47 222 48 223
rect 46 222 47 223
rect 45 222 46 223
rect 44 222 45 223
rect 43 222 44 223
rect 42 222 43 223
rect 41 222 42 223
rect 40 222 41 223
rect 39 222 40 223
rect 38 222 39 223
rect 37 222 38 223
rect 36 222 37 223
rect 35 222 36 223
rect 34 222 35 223
rect 33 222 34 223
rect 32 222 33 223
rect 31 222 32 223
rect 30 222 31 223
rect 29 222 30 223
rect 28 222 29 223
rect 27 222 28 223
rect 26 222 27 223
rect 25 222 26 223
rect 24 222 25 223
rect 23 222 24 223
rect 22 222 23 223
rect 21 222 22 223
rect 20 222 21 223
rect 19 222 20 223
rect 18 222 19 223
rect 17 222 18 223
rect 16 222 17 223
rect 15 222 16 223
rect 14 222 15 223
rect 13 222 14 223
rect 12 222 13 223
rect 11 222 12 223
rect 10 222 11 223
rect 9 222 10 223
rect 482 223 483 224
rect 481 223 482 224
rect 480 223 481 224
rect 479 223 480 224
rect 478 223 479 224
rect 477 223 478 224
rect 476 223 477 224
rect 475 223 476 224
rect 474 223 475 224
rect 473 223 474 224
rect 472 223 473 224
rect 471 223 472 224
rect 470 223 471 224
rect 469 223 470 224
rect 468 223 469 224
rect 467 223 468 224
rect 466 223 467 224
rect 465 223 466 224
rect 464 223 465 224
rect 463 223 464 224
rect 462 223 463 224
rect 440 223 441 224
rect 439 223 440 224
rect 438 223 439 224
rect 437 223 438 224
rect 436 223 437 224
rect 435 223 436 224
rect 434 223 435 224
rect 433 223 434 224
rect 405 223 406 224
rect 404 223 405 224
rect 403 223 404 224
rect 402 223 403 224
rect 401 223 402 224
rect 400 223 401 224
rect 399 223 400 224
rect 398 223 399 224
rect 363 223 364 224
rect 362 223 363 224
rect 361 223 362 224
rect 360 223 361 224
rect 359 223 360 224
rect 358 223 359 224
rect 357 223 358 224
rect 292 223 293 224
rect 291 223 292 224
rect 290 223 291 224
rect 289 223 290 224
rect 288 223 289 224
rect 287 223 288 224
rect 286 223 287 224
rect 285 223 286 224
rect 284 223 285 224
rect 283 223 284 224
rect 282 223 283 224
rect 281 223 282 224
rect 280 223 281 224
rect 279 223 280 224
rect 278 223 279 224
rect 277 223 278 224
rect 276 223 277 224
rect 275 223 276 224
rect 274 223 275 224
rect 273 223 274 224
rect 272 223 273 224
rect 271 223 272 224
rect 270 223 271 224
rect 269 223 270 224
rect 268 223 269 224
rect 267 223 268 224
rect 266 223 267 224
rect 265 223 266 224
rect 264 223 265 224
rect 263 223 264 224
rect 262 223 263 224
rect 261 223 262 224
rect 260 223 261 224
rect 259 223 260 224
rect 258 223 259 224
rect 257 223 258 224
rect 256 223 257 224
rect 255 223 256 224
rect 254 223 255 224
rect 253 223 254 224
rect 252 223 253 224
rect 251 223 252 224
rect 250 223 251 224
rect 249 223 250 224
rect 248 223 249 224
rect 247 223 248 224
rect 246 223 247 224
rect 245 223 246 224
rect 244 223 245 224
rect 243 223 244 224
rect 242 223 243 224
rect 241 223 242 224
rect 240 223 241 224
rect 239 223 240 224
rect 238 223 239 224
rect 237 223 238 224
rect 236 223 237 224
rect 235 223 236 224
rect 234 223 235 224
rect 233 223 234 224
rect 232 223 233 224
rect 231 223 232 224
rect 230 223 231 224
rect 229 223 230 224
rect 228 223 229 224
rect 227 223 228 224
rect 226 223 227 224
rect 225 223 226 224
rect 224 223 225 224
rect 223 223 224 224
rect 222 223 223 224
rect 221 223 222 224
rect 220 223 221 224
rect 219 223 220 224
rect 218 223 219 224
rect 217 223 218 224
rect 216 223 217 224
rect 215 223 216 224
rect 214 223 215 224
rect 213 223 214 224
rect 212 223 213 224
rect 211 223 212 224
rect 210 223 211 224
rect 209 223 210 224
rect 208 223 209 224
rect 207 223 208 224
rect 206 223 207 224
rect 205 223 206 224
rect 204 223 205 224
rect 203 223 204 224
rect 202 223 203 224
rect 201 223 202 224
rect 200 223 201 224
rect 199 223 200 224
rect 198 223 199 224
rect 197 223 198 224
rect 196 223 197 224
rect 195 223 196 224
rect 194 223 195 224
rect 193 223 194 224
rect 192 223 193 224
rect 191 223 192 224
rect 190 223 191 224
rect 189 223 190 224
rect 188 223 189 224
rect 187 223 188 224
rect 186 223 187 224
rect 185 223 186 224
rect 184 223 185 224
rect 183 223 184 224
rect 182 223 183 224
rect 181 223 182 224
rect 180 223 181 224
rect 179 223 180 224
rect 146 223 147 224
rect 145 223 146 224
rect 144 223 145 224
rect 143 223 144 224
rect 142 223 143 224
rect 141 223 142 224
rect 140 223 141 224
rect 139 223 140 224
rect 138 223 139 224
rect 137 223 138 224
rect 136 223 137 224
rect 135 223 136 224
rect 134 223 135 224
rect 133 223 134 224
rect 132 223 133 224
rect 131 223 132 224
rect 130 223 131 224
rect 129 223 130 224
rect 128 223 129 224
rect 127 223 128 224
rect 126 223 127 224
rect 125 223 126 224
rect 124 223 125 224
rect 123 223 124 224
rect 122 223 123 224
rect 121 223 122 224
rect 120 223 121 224
rect 119 223 120 224
rect 118 223 119 224
rect 117 223 118 224
rect 116 223 117 224
rect 115 223 116 224
rect 114 223 115 224
rect 113 223 114 224
rect 112 223 113 224
rect 111 223 112 224
rect 110 223 111 224
rect 109 223 110 224
rect 108 223 109 224
rect 107 223 108 224
rect 106 223 107 224
rect 74 223 75 224
rect 73 223 74 224
rect 72 223 73 224
rect 71 223 72 224
rect 70 223 71 224
rect 69 223 70 224
rect 68 223 69 224
rect 67 223 68 224
rect 66 223 67 224
rect 65 223 66 224
rect 64 223 65 224
rect 63 223 64 224
rect 62 223 63 224
rect 61 223 62 224
rect 60 223 61 224
rect 59 223 60 224
rect 58 223 59 224
rect 57 223 58 224
rect 56 223 57 224
rect 55 223 56 224
rect 54 223 55 224
rect 53 223 54 224
rect 52 223 53 224
rect 51 223 52 224
rect 50 223 51 224
rect 49 223 50 224
rect 48 223 49 224
rect 47 223 48 224
rect 46 223 47 224
rect 45 223 46 224
rect 44 223 45 224
rect 43 223 44 224
rect 42 223 43 224
rect 41 223 42 224
rect 40 223 41 224
rect 39 223 40 224
rect 38 223 39 224
rect 37 223 38 224
rect 36 223 37 224
rect 35 223 36 224
rect 34 223 35 224
rect 33 223 34 224
rect 32 223 33 224
rect 31 223 32 224
rect 30 223 31 224
rect 29 223 30 224
rect 28 223 29 224
rect 27 223 28 224
rect 26 223 27 224
rect 25 223 26 224
rect 24 223 25 224
rect 23 223 24 224
rect 22 223 23 224
rect 21 223 22 224
rect 20 223 21 224
rect 19 223 20 224
rect 18 223 19 224
rect 17 223 18 224
rect 16 223 17 224
rect 15 223 16 224
rect 14 223 15 224
rect 13 223 14 224
rect 12 223 13 224
rect 11 223 12 224
rect 10 223 11 224
rect 9 223 10 224
rect 482 224 483 225
rect 481 224 482 225
rect 480 224 481 225
rect 479 224 480 225
rect 478 224 479 225
rect 477 224 478 225
rect 476 224 477 225
rect 475 224 476 225
rect 474 224 475 225
rect 473 224 474 225
rect 472 224 473 225
rect 471 224 472 225
rect 470 224 471 225
rect 469 224 470 225
rect 468 224 469 225
rect 467 224 468 225
rect 466 224 467 225
rect 465 224 466 225
rect 464 224 465 225
rect 463 224 464 225
rect 462 224 463 225
rect 441 224 442 225
rect 440 224 441 225
rect 439 224 440 225
rect 438 224 439 225
rect 437 224 438 225
rect 436 224 437 225
rect 435 224 436 225
rect 434 224 435 225
rect 403 224 404 225
rect 402 224 403 225
rect 401 224 402 225
rect 400 224 401 225
rect 399 224 400 225
rect 398 224 399 225
rect 364 224 365 225
rect 363 224 364 225
rect 362 224 363 225
rect 361 224 362 225
rect 360 224 361 225
rect 291 224 292 225
rect 290 224 291 225
rect 289 224 290 225
rect 288 224 289 225
rect 287 224 288 225
rect 286 224 287 225
rect 285 224 286 225
rect 284 224 285 225
rect 283 224 284 225
rect 282 224 283 225
rect 281 224 282 225
rect 280 224 281 225
rect 279 224 280 225
rect 278 224 279 225
rect 277 224 278 225
rect 276 224 277 225
rect 275 224 276 225
rect 274 224 275 225
rect 273 224 274 225
rect 272 224 273 225
rect 271 224 272 225
rect 270 224 271 225
rect 269 224 270 225
rect 268 224 269 225
rect 267 224 268 225
rect 266 224 267 225
rect 265 224 266 225
rect 264 224 265 225
rect 263 224 264 225
rect 262 224 263 225
rect 261 224 262 225
rect 260 224 261 225
rect 259 224 260 225
rect 258 224 259 225
rect 257 224 258 225
rect 256 224 257 225
rect 255 224 256 225
rect 254 224 255 225
rect 253 224 254 225
rect 252 224 253 225
rect 251 224 252 225
rect 250 224 251 225
rect 249 224 250 225
rect 248 224 249 225
rect 247 224 248 225
rect 246 224 247 225
rect 245 224 246 225
rect 244 224 245 225
rect 243 224 244 225
rect 242 224 243 225
rect 241 224 242 225
rect 240 224 241 225
rect 239 224 240 225
rect 238 224 239 225
rect 237 224 238 225
rect 236 224 237 225
rect 235 224 236 225
rect 234 224 235 225
rect 233 224 234 225
rect 232 224 233 225
rect 231 224 232 225
rect 230 224 231 225
rect 229 224 230 225
rect 228 224 229 225
rect 227 224 228 225
rect 226 224 227 225
rect 225 224 226 225
rect 224 224 225 225
rect 223 224 224 225
rect 222 224 223 225
rect 221 224 222 225
rect 220 224 221 225
rect 219 224 220 225
rect 218 224 219 225
rect 217 224 218 225
rect 216 224 217 225
rect 215 224 216 225
rect 214 224 215 225
rect 213 224 214 225
rect 212 224 213 225
rect 211 224 212 225
rect 210 224 211 225
rect 209 224 210 225
rect 208 224 209 225
rect 207 224 208 225
rect 206 224 207 225
rect 205 224 206 225
rect 204 224 205 225
rect 203 224 204 225
rect 202 224 203 225
rect 201 224 202 225
rect 200 224 201 225
rect 199 224 200 225
rect 198 224 199 225
rect 197 224 198 225
rect 196 224 197 225
rect 195 224 196 225
rect 194 224 195 225
rect 193 224 194 225
rect 192 224 193 225
rect 191 224 192 225
rect 190 224 191 225
rect 189 224 190 225
rect 188 224 189 225
rect 187 224 188 225
rect 186 224 187 225
rect 185 224 186 225
rect 184 224 185 225
rect 183 224 184 225
rect 182 224 183 225
rect 181 224 182 225
rect 180 224 181 225
rect 179 224 180 225
rect 178 224 179 225
rect 177 224 178 225
rect 146 224 147 225
rect 145 224 146 225
rect 144 224 145 225
rect 143 224 144 225
rect 142 224 143 225
rect 141 224 142 225
rect 140 224 141 225
rect 139 224 140 225
rect 138 224 139 225
rect 137 224 138 225
rect 136 224 137 225
rect 135 224 136 225
rect 134 224 135 225
rect 133 224 134 225
rect 132 224 133 225
rect 131 224 132 225
rect 130 224 131 225
rect 129 224 130 225
rect 128 224 129 225
rect 127 224 128 225
rect 126 224 127 225
rect 125 224 126 225
rect 124 224 125 225
rect 123 224 124 225
rect 122 224 123 225
rect 121 224 122 225
rect 120 224 121 225
rect 119 224 120 225
rect 118 224 119 225
rect 117 224 118 225
rect 116 224 117 225
rect 115 224 116 225
rect 114 224 115 225
rect 113 224 114 225
rect 112 224 113 225
rect 111 224 112 225
rect 110 224 111 225
rect 109 224 110 225
rect 108 224 109 225
rect 75 224 76 225
rect 74 224 75 225
rect 73 224 74 225
rect 72 224 73 225
rect 71 224 72 225
rect 70 224 71 225
rect 69 224 70 225
rect 68 224 69 225
rect 67 224 68 225
rect 66 224 67 225
rect 65 224 66 225
rect 64 224 65 225
rect 63 224 64 225
rect 62 224 63 225
rect 61 224 62 225
rect 60 224 61 225
rect 59 224 60 225
rect 58 224 59 225
rect 57 224 58 225
rect 56 224 57 225
rect 55 224 56 225
rect 54 224 55 225
rect 53 224 54 225
rect 52 224 53 225
rect 51 224 52 225
rect 50 224 51 225
rect 49 224 50 225
rect 48 224 49 225
rect 47 224 48 225
rect 46 224 47 225
rect 45 224 46 225
rect 44 224 45 225
rect 43 224 44 225
rect 42 224 43 225
rect 41 224 42 225
rect 40 224 41 225
rect 39 224 40 225
rect 38 224 39 225
rect 37 224 38 225
rect 36 224 37 225
rect 35 224 36 225
rect 34 224 35 225
rect 33 224 34 225
rect 32 224 33 225
rect 31 224 32 225
rect 30 224 31 225
rect 29 224 30 225
rect 28 224 29 225
rect 27 224 28 225
rect 26 224 27 225
rect 25 224 26 225
rect 24 224 25 225
rect 23 224 24 225
rect 22 224 23 225
rect 21 224 22 225
rect 20 224 21 225
rect 19 224 20 225
rect 18 224 19 225
rect 17 224 18 225
rect 16 224 17 225
rect 15 224 16 225
rect 14 224 15 225
rect 13 224 14 225
rect 12 224 13 225
rect 11 224 12 225
rect 10 224 11 225
rect 9 224 10 225
rect 8 224 9 225
rect 482 225 483 226
rect 481 225 482 226
rect 473 225 474 226
rect 472 225 473 226
rect 463 225 464 226
rect 462 225 463 226
rect 441 225 442 226
rect 440 225 441 226
rect 439 225 440 226
rect 438 225 439 226
rect 437 225 438 226
rect 436 225 437 226
rect 402 225 403 226
rect 401 225 402 226
rect 400 225 401 226
rect 399 225 400 226
rect 398 225 399 226
rect 364 225 365 226
rect 363 225 364 226
rect 362 225 363 226
rect 289 225 290 226
rect 288 225 289 226
rect 287 225 288 226
rect 286 225 287 226
rect 285 225 286 226
rect 284 225 285 226
rect 283 225 284 226
rect 282 225 283 226
rect 281 225 282 226
rect 280 225 281 226
rect 279 225 280 226
rect 278 225 279 226
rect 277 225 278 226
rect 276 225 277 226
rect 275 225 276 226
rect 274 225 275 226
rect 273 225 274 226
rect 272 225 273 226
rect 271 225 272 226
rect 270 225 271 226
rect 269 225 270 226
rect 268 225 269 226
rect 267 225 268 226
rect 266 225 267 226
rect 265 225 266 226
rect 264 225 265 226
rect 263 225 264 226
rect 262 225 263 226
rect 261 225 262 226
rect 260 225 261 226
rect 259 225 260 226
rect 258 225 259 226
rect 257 225 258 226
rect 256 225 257 226
rect 255 225 256 226
rect 254 225 255 226
rect 253 225 254 226
rect 252 225 253 226
rect 251 225 252 226
rect 250 225 251 226
rect 249 225 250 226
rect 248 225 249 226
rect 247 225 248 226
rect 246 225 247 226
rect 245 225 246 226
rect 244 225 245 226
rect 243 225 244 226
rect 242 225 243 226
rect 241 225 242 226
rect 240 225 241 226
rect 239 225 240 226
rect 238 225 239 226
rect 237 225 238 226
rect 236 225 237 226
rect 235 225 236 226
rect 234 225 235 226
rect 233 225 234 226
rect 232 225 233 226
rect 231 225 232 226
rect 230 225 231 226
rect 229 225 230 226
rect 228 225 229 226
rect 227 225 228 226
rect 226 225 227 226
rect 225 225 226 226
rect 224 225 225 226
rect 223 225 224 226
rect 222 225 223 226
rect 221 225 222 226
rect 220 225 221 226
rect 219 225 220 226
rect 218 225 219 226
rect 217 225 218 226
rect 216 225 217 226
rect 215 225 216 226
rect 214 225 215 226
rect 213 225 214 226
rect 212 225 213 226
rect 211 225 212 226
rect 210 225 211 226
rect 209 225 210 226
rect 208 225 209 226
rect 207 225 208 226
rect 206 225 207 226
rect 205 225 206 226
rect 204 225 205 226
rect 203 225 204 226
rect 202 225 203 226
rect 201 225 202 226
rect 200 225 201 226
rect 199 225 200 226
rect 198 225 199 226
rect 197 225 198 226
rect 196 225 197 226
rect 195 225 196 226
rect 194 225 195 226
rect 193 225 194 226
rect 192 225 193 226
rect 191 225 192 226
rect 190 225 191 226
rect 189 225 190 226
rect 188 225 189 226
rect 187 225 188 226
rect 186 225 187 226
rect 185 225 186 226
rect 184 225 185 226
rect 183 225 184 226
rect 182 225 183 226
rect 181 225 182 226
rect 180 225 181 226
rect 179 225 180 226
rect 178 225 179 226
rect 177 225 178 226
rect 176 225 177 226
rect 175 225 176 226
rect 146 225 147 226
rect 145 225 146 226
rect 144 225 145 226
rect 143 225 144 226
rect 142 225 143 226
rect 141 225 142 226
rect 140 225 141 226
rect 139 225 140 226
rect 138 225 139 226
rect 137 225 138 226
rect 136 225 137 226
rect 135 225 136 226
rect 134 225 135 226
rect 133 225 134 226
rect 132 225 133 226
rect 131 225 132 226
rect 130 225 131 226
rect 129 225 130 226
rect 128 225 129 226
rect 127 225 128 226
rect 126 225 127 226
rect 125 225 126 226
rect 124 225 125 226
rect 123 225 124 226
rect 122 225 123 226
rect 121 225 122 226
rect 120 225 121 226
rect 119 225 120 226
rect 118 225 119 226
rect 117 225 118 226
rect 116 225 117 226
rect 115 225 116 226
rect 114 225 115 226
rect 113 225 114 226
rect 112 225 113 226
rect 111 225 112 226
rect 110 225 111 226
rect 109 225 110 226
rect 77 225 78 226
rect 76 225 77 226
rect 75 225 76 226
rect 74 225 75 226
rect 73 225 74 226
rect 72 225 73 226
rect 71 225 72 226
rect 70 225 71 226
rect 69 225 70 226
rect 68 225 69 226
rect 67 225 68 226
rect 66 225 67 226
rect 65 225 66 226
rect 64 225 65 226
rect 63 225 64 226
rect 62 225 63 226
rect 61 225 62 226
rect 60 225 61 226
rect 59 225 60 226
rect 58 225 59 226
rect 57 225 58 226
rect 56 225 57 226
rect 55 225 56 226
rect 54 225 55 226
rect 53 225 54 226
rect 52 225 53 226
rect 51 225 52 226
rect 50 225 51 226
rect 49 225 50 226
rect 48 225 49 226
rect 47 225 48 226
rect 46 225 47 226
rect 45 225 46 226
rect 44 225 45 226
rect 43 225 44 226
rect 42 225 43 226
rect 41 225 42 226
rect 40 225 41 226
rect 39 225 40 226
rect 38 225 39 226
rect 37 225 38 226
rect 36 225 37 226
rect 35 225 36 226
rect 34 225 35 226
rect 33 225 34 226
rect 32 225 33 226
rect 31 225 32 226
rect 30 225 31 226
rect 29 225 30 226
rect 28 225 29 226
rect 27 225 28 226
rect 26 225 27 226
rect 25 225 26 226
rect 24 225 25 226
rect 23 225 24 226
rect 22 225 23 226
rect 21 225 22 226
rect 20 225 21 226
rect 19 225 20 226
rect 18 225 19 226
rect 17 225 18 226
rect 16 225 17 226
rect 15 225 16 226
rect 14 225 15 226
rect 13 225 14 226
rect 12 225 13 226
rect 11 225 12 226
rect 10 225 11 226
rect 9 225 10 226
rect 8 225 9 226
rect 482 226 483 227
rect 473 226 474 227
rect 462 226 463 227
rect 441 226 442 227
rect 440 226 441 227
rect 439 226 440 227
rect 438 226 439 227
rect 437 226 438 227
rect 401 226 402 227
rect 400 226 401 227
rect 399 226 400 227
rect 398 226 399 227
rect 397 226 398 227
rect 364 226 365 227
rect 287 226 288 227
rect 286 226 287 227
rect 285 226 286 227
rect 284 226 285 227
rect 283 226 284 227
rect 282 226 283 227
rect 281 226 282 227
rect 280 226 281 227
rect 279 226 280 227
rect 278 226 279 227
rect 277 226 278 227
rect 276 226 277 227
rect 275 226 276 227
rect 274 226 275 227
rect 273 226 274 227
rect 272 226 273 227
rect 271 226 272 227
rect 270 226 271 227
rect 269 226 270 227
rect 268 226 269 227
rect 267 226 268 227
rect 266 226 267 227
rect 265 226 266 227
rect 264 226 265 227
rect 263 226 264 227
rect 262 226 263 227
rect 261 226 262 227
rect 260 226 261 227
rect 259 226 260 227
rect 258 226 259 227
rect 257 226 258 227
rect 256 226 257 227
rect 255 226 256 227
rect 254 226 255 227
rect 253 226 254 227
rect 252 226 253 227
rect 251 226 252 227
rect 250 226 251 227
rect 249 226 250 227
rect 248 226 249 227
rect 247 226 248 227
rect 246 226 247 227
rect 245 226 246 227
rect 244 226 245 227
rect 243 226 244 227
rect 242 226 243 227
rect 241 226 242 227
rect 240 226 241 227
rect 239 226 240 227
rect 238 226 239 227
rect 237 226 238 227
rect 236 226 237 227
rect 235 226 236 227
rect 234 226 235 227
rect 233 226 234 227
rect 232 226 233 227
rect 231 226 232 227
rect 230 226 231 227
rect 229 226 230 227
rect 228 226 229 227
rect 227 226 228 227
rect 226 226 227 227
rect 225 226 226 227
rect 224 226 225 227
rect 223 226 224 227
rect 222 226 223 227
rect 221 226 222 227
rect 220 226 221 227
rect 219 226 220 227
rect 218 226 219 227
rect 217 226 218 227
rect 216 226 217 227
rect 215 226 216 227
rect 214 226 215 227
rect 213 226 214 227
rect 212 226 213 227
rect 211 226 212 227
rect 210 226 211 227
rect 209 226 210 227
rect 208 226 209 227
rect 207 226 208 227
rect 206 226 207 227
rect 205 226 206 227
rect 204 226 205 227
rect 203 226 204 227
rect 202 226 203 227
rect 201 226 202 227
rect 200 226 201 227
rect 199 226 200 227
rect 198 226 199 227
rect 197 226 198 227
rect 196 226 197 227
rect 195 226 196 227
rect 194 226 195 227
rect 193 226 194 227
rect 192 226 193 227
rect 191 226 192 227
rect 190 226 191 227
rect 189 226 190 227
rect 188 226 189 227
rect 187 226 188 227
rect 186 226 187 227
rect 185 226 186 227
rect 184 226 185 227
rect 183 226 184 227
rect 182 226 183 227
rect 181 226 182 227
rect 180 226 181 227
rect 179 226 180 227
rect 178 226 179 227
rect 177 226 178 227
rect 176 226 177 227
rect 175 226 176 227
rect 174 226 175 227
rect 173 226 174 227
rect 146 226 147 227
rect 145 226 146 227
rect 144 226 145 227
rect 143 226 144 227
rect 142 226 143 227
rect 141 226 142 227
rect 140 226 141 227
rect 139 226 140 227
rect 138 226 139 227
rect 137 226 138 227
rect 136 226 137 227
rect 135 226 136 227
rect 134 226 135 227
rect 133 226 134 227
rect 132 226 133 227
rect 131 226 132 227
rect 130 226 131 227
rect 129 226 130 227
rect 128 226 129 227
rect 127 226 128 227
rect 126 226 127 227
rect 125 226 126 227
rect 124 226 125 227
rect 123 226 124 227
rect 122 226 123 227
rect 121 226 122 227
rect 120 226 121 227
rect 119 226 120 227
rect 118 226 119 227
rect 117 226 118 227
rect 116 226 117 227
rect 115 226 116 227
rect 114 226 115 227
rect 113 226 114 227
rect 112 226 113 227
rect 111 226 112 227
rect 78 226 79 227
rect 77 226 78 227
rect 76 226 77 227
rect 75 226 76 227
rect 74 226 75 227
rect 73 226 74 227
rect 72 226 73 227
rect 71 226 72 227
rect 70 226 71 227
rect 69 226 70 227
rect 68 226 69 227
rect 67 226 68 227
rect 66 226 67 227
rect 65 226 66 227
rect 64 226 65 227
rect 63 226 64 227
rect 62 226 63 227
rect 61 226 62 227
rect 60 226 61 227
rect 59 226 60 227
rect 58 226 59 227
rect 57 226 58 227
rect 56 226 57 227
rect 55 226 56 227
rect 54 226 55 227
rect 53 226 54 227
rect 52 226 53 227
rect 51 226 52 227
rect 50 226 51 227
rect 49 226 50 227
rect 48 226 49 227
rect 47 226 48 227
rect 46 226 47 227
rect 45 226 46 227
rect 44 226 45 227
rect 43 226 44 227
rect 42 226 43 227
rect 41 226 42 227
rect 40 226 41 227
rect 39 226 40 227
rect 38 226 39 227
rect 37 226 38 227
rect 36 226 37 227
rect 35 226 36 227
rect 34 226 35 227
rect 33 226 34 227
rect 32 226 33 227
rect 31 226 32 227
rect 30 226 31 227
rect 29 226 30 227
rect 28 226 29 227
rect 27 226 28 227
rect 26 226 27 227
rect 25 226 26 227
rect 24 226 25 227
rect 23 226 24 227
rect 22 226 23 227
rect 21 226 22 227
rect 20 226 21 227
rect 19 226 20 227
rect 18 226 19 227
rect 17 226 18 227
rect 16 226 17 227
rect 15 226 16 227
rect 14 226 15 227
rect 13 226 14 227
rect 12 226 13 227
rect 11 226 12 227
rect 10 226 11 227
rect 9 226 10 227
rect 8 226 9 227
rect 482 227 483 228
rect 474 227 475 228
rect 473 227 474 228
rect 472 227 473 228
rect 462 227 463 228
rect 441 227 442 228
rect 440 227 441 228
rect 439 227 440 228
rect 438 227 439 228
rect 437 227 438 228
rect 401 227 402 228
rect 400 227 401 228
rect 399 227 400 228
rect 398 227 399 228
rect 397 227 398 228
rect 286 227 287 228
rect 285 227 286 228
rect 284 227 285 228
rect 283 227 284 228
rect 282 227 283 228
rect 281 227 282 228
rect 280 227 281 228
rect 279 227 280 228
rect 278 227 279 228
rect 277 227 278 228
rect 276 227 277 228
rect 275 227 276 228
rect 274 227 275 228
rect 273 227 274 228
rect 272 227 273 228
rect 271 227 272 228
rect 270 227 271 228
rect 269 227 270 228
rect 268 227 269 228
rect 267 227 268 228
rect 266 227 267 228
rect 265 227 266 228
rect 264 227 265 228
rect 263 227 264 228
rect 262 227 263 228
rect 261 227 262 228
rect 260 227 261 228
rect 259 227 260 228
rect 258 227 259 228
rect 257 227 258 228
rect 256 227 257 228
rect 255 227 256 228
rect 254 227 255 228
rect 253 227 254 228
rect 252 227 253 228
rect 251 227 252 228
rect 250 227 251 228
rect 249 227 250 228
rect 248 227 249 228
rect 247 227 248 228
rect 246 227 247 228
rect 245 227 246 228
rect 244 227 245 228
rect 243 227 244 228
rect 242 227 243 228
rect 241 227 242 228
rect 240 227 241 228
rect 239 227 240 228
rect 238 227 239 228
rect 237 227 238 228
rect 236 227 237 228
rect 235 227 236 228
rect 234 227 235 228
rect 233 227 234 228
rect 232 227 233 228
rect 231 227 232 228
rect 230 227 231 228
rect 229 227 230 228
rect 228 227 229 228
rect 227 227 228 228
rect 226 227 227 228
rect 225 227 226 228
rect 224 227 225 228
rect 223 227 224 228
rect 222 227 223 228
rect 221 227 222 228
rect 220 227 221 228
rect 219 227 220 228
rect 218 227 219 228
rect 217 227 218 228
rect 216 227 217 228
rect 215 227 216 228
rect 214 227 215 228
rect 213 227 214 228
rect 212 227 213 228
rect 211 227 212 228
rect 210 227 211 228
rect 209 227 210 228
rect 208 227 209 228
rect 207 227 208 228
rect 206 227 207 228
rect 205 227 206 228
rect 204 227 205 228
rect 203 227 204 228
rect 202 227 203 228
rect 201 227 202 228
rect 200 227 201 228
rect 199 227 200 228
rect 198 227 199 228
rect 197 227 198 228
rect 196 227 197 228
rect 195 227 196 228
rect 194 227 195 228
rect 193 227 194 228
rect 192 227 193 228
rect 191 227 192 228
rect 190 227 191 228
rect 189 227 190 228
rect 188 227 189 228
rect 187 227 188 228
rect 186 227 187 228
rect 185 227 186 228
rect 184 227 185 228
rect 183 227 184 228
rect 182 227 183 228
rect 181 227 182 228
rect 180 227 181 228
rect 179 227 180 228
rect 178 227 179 228
rect 177 227 178 228
rect 176 227 177 228
rect 175 227 176 228
rect 174 227 175 228
rect 173 227 174 228
rect 172 227 173 228
rect 171 227 172 228
rect 146 227 147 228
rect 145 227 146 228
rect 144 227 145 228
rect 143 227 144 228
rect 142 227 143 228
rect 141 227 142 228
rect 140 227 141 228
rect 139 227 140 228
rect 138 227 139 228
rect 137 227 138 228
rect 136 227 137 228
rect 135 227 136 228
rect 134 227 135 228
rect 133 227 134 228
rect 132 227 133 228
rect 131 227 132 228
rect 130 227 131 228
rect 129 227 130 228
rect 128 227 129 228
rect 127 227 128 228
rect 126 227 127 228
rect 125 227 126 228
rect 124 227 125 228
rect 123 227 124 228
rect 122 227 123 228
rect 121 227 122 228
rect 120 227 121 228
rect 119 227 120 228
rect 118 227 119 228
rect 117 227 118 228
rect 116 227 117 228
rect 115 227 116 228
rect 114 227 115 228
rect 113 227 114 228
rect 112 227 113 228
rect 79 227 80 228
rect 78 227 79 228
rect 77 227 78 228
rect 76 227 77 228
rect 75 227 76 228
rect 74 227 75 228
rect 73 227 74 228
rect 72 227 73 228
rect 71 227 72 228
rect 70 227 71 228
rect 69 227 70 228
rect 68 227 69 228
rect 67 227 68 228
rect 66 227 67 228
rect 65 227 66 228
rect 64 227 65 228
rect 63 227 64 228
rect 62 227 63 228
rect 61 227 62 228
rect 60 227 61 228
rect 59 227 60 228
rect 58 227 59 228
rect 57 227 58 228
rect 56 227 57 228
rect 55 227 56 228
rect 54 227 55 228
rect 53 227 54 228
rect 52 227 53 228
rect 51 227 52 228
rect 50 227 51 228
rect 49 227 50 228
rect 48 227 49 228
rect 47 227 48 228
rect 46 227 47 228
rect 45 227 46 228
rect 44 227 45 228
rect 43 227 44 228
rect 42 227 43 228
rect 41 227 42 228
rect 40 227 41 228
rect 39 227 40 228
rect 38 227 39 228
rect 37 227 38 228
rect 36 227 37 228
rect 35 227 36 228
rect 34 227 35 228
rect 33 227 34 228
rect 32 227 33 228
rect 31 227 32 228
rect 30 227 31 228
rect 29 227 30 228
rect 28 227 29 228
rect 27 227 28 228
rect 26 227 27 228
rect 25 227 26 228
rect 24 227 25 228
rect 23 227 24 228
rect 22 227 23 228
rect 21 227 22 228
rect 20 227 21 228
rect 19 227 20 228
rect 18 227 19 228
rect 17 227 18 228
rect 16 227 17 228
rect 15 227 16 228
rect 14 227 15 228
rect 13 227 14 228
rect 12 227 13 228
rect 11 227 12 228
rect 10 227 11 228
rect 9 227 10 228
rect 8 227 9 228
rect 476 228 477 229
rect 475 228 476 229
rect 474 228 475 229
rect 473 228 474 229
rect 472 228 473 229
rect 463 228 464 229
rect 462 228 463 229
rect 442 228 443 229
rect 441 228 442 229
rect 440 228 441 229
rect 439 228 440 229
rect 438 228 439 229
rect 400 228 401 229
rect 399 228 400 229
rect 398 228 399 229
rect 397 228 398 229
rect 284 228 285 229
rect 283 228 284 229
rect 282 228 283 229
rect 281 228 282 229
rect 280 228 281 229
rect 279 228 280 229
rect 278 228 279 229
rect 277 228 278 229
rect 276 228 277 229
rect 275 228 276 229
rect 274 228 275 229
rect 273 228 274 229
rect 272 228 273 229
rect 271 228 272 229
rect 270 228 271 229
rect 269 228 270 229
rect 268 228 269 229
rect 267 228 268 229
rect 266 228 267 229
rect 265 228 266 229
rect 264 228 265 229
rect 263 228 264 229
rect 262 228 263 229
rect 261 228 262 229
rect 260 228 261 229
rect 259 228 260 229
rect 258 228 259 229
rect 257 228 258 229
rect 256 228 257 229
rect 255 228 256 229
rect 254 228 255 229
rect 253 228 254 229
rect 252 228 253 229
rect 251 228 252 229
rect 250 228 251 229
rect 249 228 250 229
rect 248 228 249 229
rect 247 228 248 229
rect 246 228 247 229
rect 245 228 246 229
rect 244 228 245 229
rect 243 228 244 229
rect 242 228 243 229
rect 241 228 242 229
rect 240 228 241 229
rect 239 228 240 229
rect 238 228 239 229
rect 237 228 238 229
rect 236 228 237 229
rect 235 228 236 229
rect 234 228 235 229
rect 233 228 234 229
rect 232 228 233 229
rect 231 228 232 229
rect 230 228 231 229
rect 229 228 230 229
rect 228 228 229 229
rect 227 228 228 229
rect 226 228 227 229
rect 225 228 226 229
rect 224 228 225 229
rect 223 228 224 229
rect 222 228 223 229
rect 221 228 222 229
rect 220 228 221 229
rect 219 228 220 229
rect 218 228 219 229
rect 217 228 218 229
rect 216 228 217 229
rect 215 228 216 229
rect 214 228 215 229
rect 213 228 214 229
rect 212 228 213 229
rect 211 228 212 229
rect 210 228 211 229
rect 209 228 210 229
rect 208 228 209 229
rect 207 228 208 229
rect 206 228 207 229
rect 205 228 206 229
rect 204 228 205 229
rect 203 228 204 229
rect 202 228 203 229
rect 201 228 202 229
rect 200 228 201 229
rect 199 228 200 229
rect 198 228 199 229
rect 197 228 198 229
rect 196 228 197 229
rect 195 228 196 229
rect 194 228 195 229
rect 193 228 194 229
rect 192 228 193 229
rect 191 228 192 229
rect 190 228 191 229
rect 189 228 190 229
rect 188 228 189 229
rect 187 228 188 229
rect 186 228 187 229
rect 185 228 186 229
rect 184 228 185 229
rect 183 228 184 229
rect 182 228 183 229
rect 181 228 182 229
rect 180 228 181 229
rect 179 228 180 229
rect 178 228 179 229
rect 177 228 178 229
rect 176 228 177 229
rect 175 228 176 229
rect 174 228 175 229
rect 173 228 174 229
rect 172 228 173 229
rect 171 228 172 229
rect 170 228 171 229
rect 169 228 170 229
rect 146 228 147 229
rect 145 228 146 229
rect 144 228 145 229
rect 143 228 144 229
rect 142 228 143 229
rect 141 228 142 229
rect 140 228 141 229
rect 139 228 140 229
rect 138 228 139 229
rect 137 228 138 229
rect 136 228 137 229
rect 135 228 136 229
rect 134 228 135 229
rect 133 228 134 229
rect 132 228 133 229
rect 131 228 132 229
rect 130 228 131 229
rect 129 228 130 229
rect 128 228 129 229
rect 127 228 128 229
rect 126 228 127 229
rect 125 228 126 229
rect 124 228 125 229
rect 123 228 124 229
rect 122 228 123 229
rect 121 228 122 229
rect 120 228 121 229
rect 119 228 120 229
rect 118 228 119 229
rect 117 228 118 229
rect 116 228 117 229
rect 115 228 116 229
rect 114 228 115 229
rect 113 228 114 229
rect 81 228 82 229
rect 80 228 81 229
rect 79 228 80 229
rect 78 228 79 229
rect 77 228 78 229
rect 76 228 77 229
rect 75 228 76 229
rect 74 228 75 229
rect 73 228 74 229
rect 72 228 73 229
rect 71 228 72 229
rect 70 228 71 229
rect 69 228 70 229
rect 68 228 69 229
rect 67 228 68 229
rect 66 228 67 229
rect 65 228 66 229
rect 64 228 65 229
rect 63 228 64 229
rect 62 228 63 229
rect 61 228 62 229
rect 60 228 61 229
rect 59 228 60 229
rect 58 228 59 229
rect 57 228 58 229
rect 56 228 57 229
rect 55 228 56 229
rect 54 228 55 229
rect 53 228 54 229
rect 52 228 53 229
rect 51 228 52 229
rect 50 228 51 229
rect 49 228 50 229
rect 48 228 49 229
rect 47 228 48 229
rect 46 228 47 229
rect 45 228 46 229
rect 44 228 45 229
rect 43 228 44 229
rect 42 228 43 229
rect 41 228 42 229
rect 40 228 41 229
rect 39 228 40 229
rect 38 228 39 229
rect 37 228 38 229
rect 36 228 37 229
rect 35 228 36 229
rect 34 228 35 229
rect 33 228 34 229
rect 32 228 33 229
rect 31 228 32 229
rect 30 228 31 229
rect 29 228 30 229
rect 28 228 29 229
rect 27 228 28 229
rect 26 228 27 229
rect 25 228 26 229
rect 24 228 25 229
rect 23 228 24 229
rect 22 228 23 229
rect 21 228 22 229
rect 20 228 21 229
rect 19 228 20 229
rect 18 228 19 229
rect 17 228 18 229
rect 16 228 17 229
rect 15 228 16 229
rect 14 228 15 229
rect 13 228 14 229
rect 12 228 13 229
rect 11 228 12 229
rect 10 228 11 229
rect 9 228 10 229
rect 8 228 9 229
rect 7 228 8 229
rect 478 229 479 230
rect 477 229 478 230
rect 476 229 477 230
rect 475 229 476 230
rect 474 229 475 230
rect 473 229 474 230
rect 472 229 473 230
rect 471 229 472 230
rect 463 229 464 230
rect 462 229 463 230
rect 442 229 443 230
rect 441 229 442 230
rect 440 229 441 230
rect 439 229 440 230
rect 399 229 400 230
rect 398 229 399 230
rect 397 229 398 230
rect 283 229 284 230
rect 282 229 283 230
rect 281 229 282 230
rect 280 229 281 230
rect 279 229 280 230
rect 278 229 279 230
rect 277 229 278 230
rect 276 229 277 230
rect 275 229 276 230
rect 274 229 275 230
rect 273 229 274 230
rect 272 229 273 230
rect 271 229 272 230
rect 270 229 271 230
rect 269 229 270 230
rect 268 229 269 230
rect 267 229 268 230
rect 266 229 267 230
rect 265 229 266 230
rect 264 229 265 230
rect 263 229 264 230
rect 262 229 263 230
rect 261 229 262 230
rect 260 229 261 230
rect 259 229 260 230
rect 258 229 259 230
rect 257 229 258 230
rect 256 229 257 230
rect 255 229 256 230
rect 254 229 255 230
rect 253 229 254 230
rect 252 229 253 230
rect 251 229 252 230
rect 250 229 251 230
rect 249 229 250 230
rect 248 229 249 230
rect 247 229 248 230
rect 246 229 247 230
rect 245 229 246 230
rect 244 229 245 230
rect 243 229 244 230
rect 242 229 243 230
rect 241 229 242 230
rect 240 229 241 230
rect 239 229 240 230
rect 238 229 239 230
rect 237 229 238 230
rect 236 229 237 230
rect 235 229 236 230
rect 234 229 235 230
rect 233 229 234 230
rect 232 229 233 230
rect 231 229 232 230
rect 230 229 231 230
rect 229 229 230 230
rect 228 229 229 230
rect 227 229 228 230
rect 226 229 227 230
rect 225 229 226 230
rect 224 229 225 230
rect 223 229 224 230
rect 222 229 223 230
rect 221 229 222 230
rect 220 229 221 230
rect 219 229 220 230
rect 218 229 219 230
rect 217 229 218 230
rect 216 229 217 230
rect 215 229 216 230
rect 214 229 215 230
rect 213 229 214 230
rect 212 229 213 230
rect 211 229 212 230
rect 210 229 211 230
rect 209 229 210 230
rect 208 229 209 230
rect 207 229 208 230
rect 206 229 207 230
rect 205 229 206 230
rect 204 229 205 230
rect 203 229 204 230
rect 202 229 203 230
rect 201 229 202 230
rect 200 229 201 230
rect 199 229 200 230
rect 198 229 199 230
rect 197 229 198 230
rect 196 229 197 230
rect 195 229 196 230
rect 194 229 195 230
rect 193 229 194 230
rect 192 229 193 230
rect 191 229 192 230
rect 190 229 191 230
rect 189 229 190 230
rect 188 229 189 230
rect 187 229 188 230
rect 186 229 187 230
rect 185 229 186 230
rect 184 229 185 230
rect 183 229 184 230
rect 182 229 183 230
rect 181 229 182 230
rect 180 229 181 230
rect 179 229 180 230
rect 178 229 179 230
rect 177 229 178 230
rect 176 229 177 230
rect 175 229 176 230
rect 174 229 175 230
rect 173 229 174 230
rect 172 229 173 230
rect 171 229 172 230
rect 170 229 171 230
rect 169 229 170 230
rect 168 229 169 230
rect 167 229 168 230
rect 166 229 167 230
rect 146 229 147 230
rect 145 229 146 230
rect 144 229 145 230
rect 143 229 144 230
rect 142 229 143 230
rect 141 229 142 230
rect 140 229 141 230
rect 139 229 140 230
rect 138 229 139 230
rect 137 229 138 230
rect 136 229 137 230
rect 135 229 136 230
rect 134 229 135 230
rect 133 229 134 230
rect 132 229 133 230
rect 131 229 132 230
rect 130 229 131 230
rect 129 229 130 230
rect 128 229 129 230
rect 127 229 128 230
rect 126 229 127 230
rect 125 229 126 230
rect 124 229 125 230
rect 123 229 124 230
rect 122 229 123 230
rect 121 229 122 230
rect 120 229 121 230
rect 119 229 120 230
rect 118 229 119 230
rect 117 229 118 230
rect 116 229 117 230
rect 115 229 116 230
rect 114 229 115 230
rect 82 229 83 230
rect 81 229 82 230
rect 80 229 81 230
rect 79 229 80 230
rect 78 229 79 230
rect 77 229 78 230
rect 76 229 77 230
rect 75 229 76 230
rect 74 229 75 230
rect 73 229 74 230
rect 72 229 73 230
rect 71 229 72 230
rect 70 229 71 230
rect 69 229 70 230
rect 68 229 69 230
rect 67 229 68 230
rect 66 229 67 230
rect 65 229 66 230
rect 64 229 65 230
rect 63 229 64 230
rect 62 229 63 230
rect 61 229 62 230
rect 60 229 61 230
rect 59 229 60 230
rect 58 229 59 230
rect 57 229 58 230
rect 56 229 57 230
rect 55 229 56 230
rect 54 229 55 230
rect 53 229 54 230
rect 52 229 53 230
rect 51 229 52 230
rect 50 229 51 230
rect 49 229 50 230
rect 48 229 49 230
rect 47 229 48 230
rect 46 229 47 230
rect 45 229 46 230
rect 44 229 45 230
rect 43 229 44 230
rect 42 229 43 230
rect 41 229 42 230
rect 40 229 41 230
rect 39 229 40 230
rect 38 229 39 230
rect 37 229 38 230
rect 36 229 37 230
rect 35 229 36 230
rect 34 229 35 230
rect 33 229 34 230
rect 32 229 33 230
rect 31 229 32 230
rect 30 229 31 230
rect 29 229 30 230
rect 28 229 29 230
rect 27 229 28 230
rect 26 229 27 230
rect 25 229 26 230
rect 24 229 25 230
rect 23 229 24 230
rect 22 229 23 230
rect 21 229 22 230
rect 20 229 21 230
rect 19 229 20 230
rect 18 229 19 230
rect 17 229 18 230
rect 16 229 17 230
rect 15 229 16 230
rect 14 229 15 230
rect 13 229 14 230
rect 12 229 13 230
rect 11 229 12 230
rect 10 229 11 230
rect 9 229 10 230
rect 8 229 9 230
rect 7 229 8 230
rect 480 230 481 231
rect 479 230 480 231
rect 478 230 479 231
rect 477 230 478 231
rect 476 230 477 231
rect 475 230 476 231
rect 474 230 475 231
rect 473 230 474 231
rect 472 230 473 231
rect 471 230 472 231
rect 470 230 471 231
rect 469 230 470 231
rect 466 230 467 231
rect 465 230 466 231
rect 464 230 465 231
rect 463 230 464 231
rect 462 230 463 231
rect 442 230 443 231
rect 441 230 442 231
rect 440 230 441 231
rect 439 230 440 231
rect 399 230 400 231
rect 398 230 399 231
rect 397 230 398 231
rect 396 230 397 231
rect 282 230 283 231
rect 281 230 282 231
rect 280 230 281 231
rect 279 230 280 231
rect 278 230 279 231
rect 277 230 278 231
rect 276 230 277 231
rect 275 230 276 231
rect 274 230 275 231
rect 273 230 274 231
rect 272 230 273 231
rect 271 230 272 231
rect 270 230 271 231
rect 269 230 270 231
rect 268 230 269 231
rect 267 230 268 231
rect 266 230 267 231
rect 265 230 266 231
rect 264 230 265 231
rect 263 230 264 231
rect 262 230 263 231
rect 261 230 262 231
rect 260 230 261 231
rect 259 230 260 231
rect 258 230 259 231
rect 257 230 258 231
rect 256 230 257 231
rect 255 230 256 231
rect 254 230 255 231
rect 253 230 254 231
rect 252 230 253 231
rect 251 230 252 231
rect 250 230 251 231
rect 249 230 250 231
rect 248 230 249 231
rect 247 230 248 231
rect 246 230 247 231
rect 245 230 246 231
rect 244 230 245 231
rect 243 230 244 231
rect 242 230 243 231
rect 241 230 242 231
rect 240 230 241 231
rect 239 230 240 231
rect 238 230 239 231
rect 237 230 238 231
rect 236 230 237 231
rect 235 230 236 231
rect 234 230 235 231
rect 233 230 234 231
rect 232 230 233 231
rect 231 230 232 231
rect 230 230 231 231
rect 229 230 230 231
rect 228 230 229 231
rect 227 230 228 231
rect 226 230 227 231
rect 225 230 226 231
rect 224 230 225 231
rect 223 230 224 231
rect 222 230 223 231
rect 221 230 222 231
rect 220 230 221 231
rect 219 230 220 231
rect 218 230 219 231
rect 217 230 218 231
rect 216 230 217 231
rect 215 230 216 231
rect 214 230 215 231
rect 213 230 214 231
rect 212 230 213 231
rect 211 230 212 231
rect 210 230 211 231
rect 209 230 210 231
rect 208 230 209 231
rect 207 230 208 231
rect 206 230 207 231
rect 205 230 206 231
rect 204 230 205 231
rect 203 230 204 231
rect 202 230 203 231
rect 201 230 202 231
rect 200 230 201 231
rect 199 230 200 231
rect 198 230 199 231
rect 197 230 198 231
rect 196 230 197 231
rect 195 230 196 231
rect 194 230 195 231
rect 193 230 194 231
rect 192 230 193 231
rect 191 230 192 231
rect 190 230 191 231
rect 189 230 190 231
rect 188 230 189 231
rect 187 230 188 231
rect 186 230 187 231
rect 185 230 186 231
rect 184 230 185 231
rect 183 230 184 231
rect 182 230 183 231
rect 181 230 182 231
rect 180 230 181 231
rect 179 230 180 231
rect 178 230 179 231
rect 177 230 178 231
rect 176 230 177 231
rect 175 230 176 231
rect 174 230 175 231
rect 173 230 174 231
rect 172 230 173 231
rect 171 230 172 231
rect 170 230 171 231
rect 169 230 170 231
rect 168 230 169 231
rect 167 230 168 231
rect 166 230 167 231
rect 165 230 166 231
rect 164 230 165 231
rect 146 230 147 231
rect 145 230 146 231
rect 144 230 145 231
rect 143 230 144 231
rect 142 230 143 231
rect 141 230 142 231
rect 140 230 141 231
rect 139 230 140 231
rect 138 230 139 231
rect 137 230 138 231
rect 136 230 137 231
rect 135 230 136 231
rect 134 230 135 231
rect 133 230 134 231
rect 132 230 133 231
rect 131 230 132 231
rect 130 230 131 231
rect 129 230 130 231
rect 128 230 129 231
rect 127 230 128 231
rect 126 230 127 231
rect 125 230 126 231
rect 124 230 125 231
rect 123 230 124 231
rect 122 230 123 231
rect 121 230 122 231
rect 120 230 121 231
rect 119 230 120 231
rect 118 230 119 231
rect 117 230 118 231
rect 116 230 117 231
rect 115 230 116 231
rect 114 230 115 231
rect 84 230 85 231
rect 83 230 84 231
rect 82 230 83 231
rect 81 230 82 231
rect 80 230 81 231
rect 79 230 80 231
rect 78 230 79 231
rect 77 230 78 231
rect 76 230 77 231
rect 75 230 76 231
rect 74 230 75 231
rect 73 230 74 231
rect 72 230 73 231
rect 71 230 72 231
rect 70 230 71 231
rect 69 230 70 231
rect 68 230 69 231
rect 67 230 68 231
rect 66 230 67 231
rect 65 230 66 231
rect 64 230 65 231
rect 63 230 64 231
rect 62 230 63 231
rect 61 230 62 231
rect 60 230 61 231
rect 59 230 60 231
rect 58 230 59 231
rect 57 230 58 231
rect 56 230 57 231
rect 55 230 56 231
rect 54 230 55 231
rect 53 230 54 231
rect 52 230 53 231
rect 51 230 52 231
rect 50 230 51 231
rect 49 230 50 231
rect 48 230 49 231
rect 47 230 48 231
rect 46 230 47 231
rect 45 230 46 231
rect 44 230 45 231
rect 43 230 44 231
rect 42 230 43 231
rect 41 230 42 231
rect 40 230 41 231
rect 39 230 40 231
rect 38 230 39 231
rect 37 230 38 231
rect 36 230 37 231
rect 35 230 36 231
rect 34 230 35 231
rect 33 230 34 231
rect 32 230 33 231
rect 31 230 32 231
rect 30 230 31 231
rect 29 230 30 231
rect 28 230 29 231
rect 27 230 28 231
rect 26 230 27 231
rect 25 230 26 231
rect 24 230 25 231
rect 23 230 24 231
rect 22 230 23 231
rect 21 230 22 231
rect 20 230 21 231
rect 19 230 20 231
rect 18 230 19 231
rect 17 230 18 231
rect 16 230 17 231
rect 15 230 16 231
rect 14 230 15 231
rect 13 230 14 231
rect 12 230 13 231
rect 11 230 12 231
rect 10 230 11 231
rect 9 230 10 231
rect 8 230 9 231
rect 7 230 8 231
rect 481 231 482 232
rect 480 231 481 232
rect 479 231 480 232
rect 478 231 479 232
rect 477 231 478 232
rect 476 231 477 232
rect 475 231 476 232
rect 474 231 475 232
rect 473 231 474 232
rect 472 231 473 232
rect 471 231 472 232
rect 470 231 471 232
rect 469 231 470 232
rect 468 231 469 232
rect 467 231 468 232
rect 466 231 467 232
rect 465 231 466 232
rect 464 231 465 232
rect 463 231 464 232
rect 462 231 463 232
rect 442 231 443 232
rect 441 231 442 232
rect 440 231 441 232
rect 439 231 440 232
rect 399 231 400 232
rect 398 231 399 232
rect 397 231 398 232
rect 396 231 397 232
rect 280 231 281 232
rect 279 231 280 232
rect 278 231 279 232
rect 277 231 278 232
rect 276 231 277 232
rect 275 231 276 232
rect 274 231 275 232
rect 273 231 274 232
rect 272 231 273 232
rect 271 231 272 232
rect 270 231 271 232
rect 269 231 270 232
rect 268 231 269 232
rect 267 231 268 232
rect 266 231 267 232
rect 265 231 266 232
rect 264 231 265 232
rect 263 231 264 232
rect 262 231 263 232
rect 261 231 262 232
rect 260 231 261 232
rect 259 231 260 232
rect 258 231 259 232
rect 257 231 258 232
rect 256 231 257 232
rect 255 231 256 232
rect 254 231 255 232
rect 253 231 254 232
rect 252 231 253 232
rect 251 231 252 232
rect 250 231 251 232
rect 249 231 250 232
rect 248 231 249 232
rect 247 231 248 232
rect 246 231 247 232
rect 245 231 246 232
rect 244 231 245 232
rect 243 231 244 232
rect 242 231 243 232
rect 241 231 242 232
rect 240 231 241 232
rect 239 231 240 232
rect 238 231 239 232
rect 237 231 238 232
rect 236 231 237 232
rect 235 231 236 232
rect 234 231 235 232
rect 233 231 234 232
rect 232 231 233 232
rect 231 231 232 232
rect 230 231 231 232
rect 229 231 230 232
rect 228 231 229 232
rect 227 231 228 232
rect 226 231 227 232
rect 225 231 226 232
rect 224 231 225 232
rect 223 231 224 232
rect 222 231 223 232
rect 221 231 222 232
rect 220 231 221 232
rect 219 231 220 232
rect 218 231 219 232
rect 217 231 218 232
rect 216 231 217 232
rect 215 231 216 232
rect 214 231 215 232
rect 213 231 214 232
rect 212 231 213 232
rect 211 231 212 232
rect 210 231 211 232
rect 209 231 210 232
rect 208 231 209 232
rect 207 231 208 232
rect 206 231 207 232
rect 205 231 206 232
rect 204 231 205 232
rect 203 231 204 232
rect 202 231 203 232
rect 201 231 202 232
rect 200 231 201 232
rect 199 231 200 232
rect 198 231 199 232
rect 197 231 198 232
rect 196 231 197 232
rect 195 231 196 232
rect 194 231 195 232
rect 193 231 194 232
rect 192 231 193 232
rect 191 231 192 232
rect 190 231 191 232
rect 189 231 190 232
rect 188 231 189 232
rect 187 231 188 232
rect 186 231 187 232
rect 185 231 186 232
rect 184 231 185 232
rect 183 231 184 232
rect 182 231 183 232
rect 181 231 182 232
rect 180 231 181 232
rect 179 231 180 232
rect 178 231 179 232
rect 177 231 178 232
rect 176 231 177 232
rect 175 231 176 232
rect 174 231 175 232
rect 173 231 174 232
rect 172 231 173 232
rect 171 231 172 232
rect 170 231 171 232
rect 169 231 170 232
rect 168 231 169 232
rect 167 231 168 232
rect 166 231 167 232
rect 165 231 166 232
rect 164 231 165 232
rect 146 231 147 232
rect 145 231 146 232
rect 144 231 145 232
rect 143 231 144 232
rect 142 231 143 232
rect 141 231 142 232
rect 140 231 141 232
rect 139 231 140 232
rect 138 231 139 232
rect 137 231 138 232
rect 136 231 137 232
rect 135 231 136 232
rect 134 231 135 232
rect 133 231 134 232
rect 132 231 133 232
rect 131 231 132 232
rect 130 231 131 232
rect 129 231 130 232
rect 128 231 129 232
rect 127 231 128 232
rect 126 231 127 232
rect 125 231 126 232
rect 124 231 125 232
rect 123 231 124 232
rect 122 231 123 232
rect 121 231 122 232
rect 120 231 121 232
rect 119 231 120 232
rect 118 231 119 232
rect 117 231 118 232
rect 116 231 117 232
rect 115 231 116 232
rect 85 231 86 232
rect 84 231 85 232
rect 83 231 84 232
rect 82 231 83 232
rect 81 231 82 232
rect 80 231 81 232
rect 79 231 80 232
rect 78 231 79 232
rect 77 231 78 232
rect 76 231 77 232
rect 75 231 76 232
rect 74 231 75 232
rect 73 231 74 232
rect 72 231 73 232
rect 71 231 72 232
rect 70 231 71 232
rect 69 231 70 232
rect 68 231 69 232
rect 67 231 68 232
rect 66 231 67 232
rect 65 231 66 232
rect 64 231 65 232
rect 63 231 64 232
rect 62 231 63 232
rect 61 231 62 232
rect 60 231 61 232
rect 59 231 60 232
rect 58 231 59 232
rect 57 231 58 232
rect 56 231 57 232
rect 55 231 56 232
rect 54 231 55 232
rect 53 231 54 232
rect 52 231 53 232
rect 51 231 52 232
rect 50 231 51 232
rect 49 231 50 232
rect 48 231 49 232
rect 47 231 48 232
rect 46 231 47 232
rect 45 231 46 232
rect 44 231 45 232
rect 43 231 44 232
rect 42 231 43 232
rect 41 231 42 232
rect 40 231 41 232
rect 39 231 40 232
rect 38 231 39 232
rect 37 231 38 232
rect 36 231 37 232
rect 35 231 36 232
rect 34 231 35 232
rect 33 231 34 232
rect 32 231 33 232
rect 31 231 32 232
rect 30 231 31 232
rect 29 231 30 232
rect 28 231 29 232
rect 27 231 28 232
rect 26 231 27 232
rect 25 231 26 232
rect 24 231 25 232
rect 23 231 24 232
rect 22 231 23 232
rect 21 231 22 232
rect 20 231 21 232
rect 19 231 20 232
rect 18 231 19 232
rect 17 231 18 232
rect 16 231 17 232
rect 15 231 16 232
rect 14 231 15 232
rect 13 231 14 232
rect 12 231 13 232
rect 11 231 12 232
rect 10 231 11 232
rect 9 231 10 232
rect 8 231 9 232
rect 7 231 8 232
rect 482 232 483 233
rect 481 232 482 233
rect 480 232 481 233
rect 479 232 480 233
rect 478 232 479 233
rect 477 232 478 233
rect 476 232 477 233
rect 475 232 476 233
rect 471 232 472 233
rect 470 232 471 233
rect 469 232 470 233
rect 468 232 469 233
rect 467 232 468 233
rect 466 232 467 233
rect 465 232 466 233
rect 464 232 465 233
rect 463 232 464 233
rect 462 232 463 233
rect 442 232 443 233
rect 441 232 442 233
rect 440 232 441 233
rect 398 232 399 233
rect 397 232 398 233
rect 396 232 397 233
rect 279 232 280 233
rect 278 232 279 233
rect 277 232 278 233
rect 276 232 277 233
rect 275 232 276 233
rect 274 232 275 233
rect 273 232 274 233
rect 272 232 273 233
rect 271 232 272 233
rect 270 232 271 233
rect 269 232 270 233
rect 268 232 269 233
rect 267 232 268 233
rect 266 232 267 233
rect 265 232 266 233
rect 264 232 265 233
rect 263 232 264 233
rect 262 232 263 233
rect 261 232 262 233
rect 260 232 261 233
rect 259 232 260 233
rect 258 232 259 233
rect 257 232 258 233
rect 256 232 257 233
rect 255 232 256 233
rect 254 232 255 233
rect 253 232 254 233
rect 252 232 253 233
rect 251 232 252 233
rect 250 232 251 233
rect 249 232 250 233
rect 248 232 249 233
rect 247 232 248 233
rect 246 232 247 233
rect 245 232 246 233
rect 244 232 245 233
rect 243 232 244 233
rect 242 232 243 233
rect 241 232 242 233
rect 240 232 241 233
rect 239 232 240 233
rect 238 232 239 233
rect 237 232 238 233
rect 236 232 237 233
rect 235 232 236 233
rect 234 232 235 233
rect 233 232 234 233
rect 232 232 233 233
rect 231 232 232 233
rect 230 232 231 233
rect 229 232 230 233
rect 228 232 229 233
rect 227 232 228 233
rect 226 232 227 233
rect 225 232 226 233
rect 224 232 225 233
rect 223 232 224 233
rect 222 232 223 233
rect 221 232 222 233
rect 220 232 221 233
rect 219 232 220 233
rect 218 232 219 233
rect 217 232 218 233
rect 216 232 217 233
rect 215 232 216 233
rect 214 232 215 233
rect 213 232 214 233
rect 212 232 213 233
rect 211 232 212 233
rect 210 232 211 233
rect 209 232 210 233
rect 208 232 209 233
rect 207 232 208 233
rect 206 232 207 233
rect 205 232 206 233
rect 204 232 205 233
rect 203 232 204 233
rect 202 232 203 233
rect 201 232 202 233
rect 200 232 201 233
rect 199 232 200 233
rect 198 232 199 233
rect 197 232 198 233
rect 196 232 197 233
rect 195 232 196 233
rect 194 232 195 233
rect 193 232 194 233
rect 192 232 193 233
rect 191 232 192 233
rect 190 232 191 233
rect 189 232 190 233
rect 188 232 189 233
rect 187 232 188 233
rect 186 232 187 233
rect 185 232 186 233
rect 184 232 185 233
rect 183 232 184 233
rect 182 232 183 233
rect 181 232 182 233
rect 180 232 181 233
rect 179 232 180 233
rect 178 232 179 233
rect 177 232 178 233
rect 176 232 177 233
rect 175 232 176 233
rect 174 232 175 233
rect 173 232 174 233
rect 172 232 173 233
rect 171 232 172 233
rect 170 232 171 233
rect 169 232 170 233
rect 168 232 169 233
rect 167 232 168 233
rect 166 232 167 233
rect 165 232 166 233
rect 147 232 148 233
rect 146 232 147 233
rect 145 232 146 233
rect 144 232 145 233
rect 143 232 144 233
rect 142 232 143 233
rect 141 232 142 233
rect 140 232 141 233
rect 139 232 140 233
rect 138 232 139 233
rect 137 232 138 233
rect 136 232 137 233
rect 135 232 136 233
rect 134 232 135 233
rect 133 232 134 233
rect 132 232 133 233
rect 131 232 132 233
rect 130 232 131 233
rect 129 232 130 233
rect 128 232 129 233
rect 127 232 128 233
rect 126 232 127 233
rect 125 232 126 233
rect 124 232 125 233
rect 123 232 124 233
rect 122 232 123 233
rect 121 232 122 233
rect 120 232 121 233
rect 119 232 120 233
rect 118 232 119 233
rect 117 232 118 233
rect 116 232 117 233
rect 87 232 88 233
rect 86 232 87 233
rect 85 232 86 233
rect 84 232 85 233
rect 83 232 84 233
rect 82 232 83 233
rect 81 232 82 233
rect 80 232 81 233
rect 79 232 80 233
rect 78 232 79 233
rect 77 232 78 233
rect 76 232 77 233
rect 75 232 76 233
rect 74 232 75 233
rect 73 232 74 233
rect 72 232 73 233
rect 71 232 72 233
rect 70 232 71 233
rect 69 232 70 233
rect 68 232 69 233
rect 67 232 68 233
rect 66 232 67 233
rect 65 232 66 233
rect 64 232 65 233
rect 63 232 64 233
rect 62 232 63 233
rect 61 232 62 233
rect 60 232 61 233
rect 59 232 60 233
rect 58 232 59 233
rect 57 232 58 233
rect 56 232 57 233
rect 55 232 56 233
rect 54 232 55 233
rect 53 232 54 233
rect 52 232 53 233
rect 51 232 52 233
rect 50 232 51 233
rect 49 232 50 233
rect 48 232 49 233
rect 47 232 48 233
rect 46 232 47 233
rect 45 232 46 233
rect 44 232 45 233
rect 43 232 44 233
rect 42 232 43 233
rect 41 232 42 233
rect 40 232 41 233
rect 39 232 40 233
rect 38 232 39 233
rect 37 232 38 233
rect 36 232 37 233
rect 35 232 36 233
rect 34 232 35 233
rect 33 232 34 233
rect 32 232 33 233
rect 31 232 32 233
rect 30 232 31 233
rect 29 232 30 233
rect 28 232 29 233
rect 27 232 28 233
rect 26 232 27 233
rect 25 232 26 233
rect 24 232 25 233
rect 23 232 24 233
rect 22 232 23 233
rect 21 232 22 233
rect 20 232 21 233
rect 19 232 20 233
rect 18 232 19 233
rect 17 232 18 233
rect 16 232 17 233
rect 15 232 16 233
rect 14 232 15 233
rect 13 232 14 233
rect 12 232 13 233
rect 11 232 12 233
rect 10 232 11 233
rect 9 232 10 233
rect 8 232 9 233
rect 7 232 8 233
rect 482 233 483 234
rect 481 233 482 234
rect 480 233 481 234
rect 479 233 480 234
rect 478 233 479 234
rect 477 233 478 234
rect 476 233 477 234
rect 471 233 472 234
rect 470 233 471 234
rect 469 233 470 234
rect 468 233 469 234
rect 467 233 468 234
rect 466 233 467 234
rect 465 233 466 234
rect 464 233 465 234
rect 463 233 464 234
rect 442 233 443 234
rect 441 233 442 234
rect 440 233 441 234
rect 398 233 399 234
rect 397 233 398 234
rect 396 233 397 234
rect 278 233 279 234
rect 277 233 278 234
rect 276 233 277 234
rect 275 233 276 234
rect 274 233 275 234
rect 273 233 274 234
rect 272 233 273 234
rect 271 233 272 234
rect 270 233 271 234
rect 269 233 270 234
rect 268 233 269 234
rect 267 233 268 234
rect 266 233 267 234
rect 265 233 266 234
rect 264 233 265 234
rect 263 233 264 234
rect 262 233 263 234
rect 261 233 262 234
rect 260 233 261 234
rect 259 233 260 234
rect 258 233 259 234
rect 257 233 258 234
rect 256 233 257 234
rect 255 233 256 234
rect 254 233 255 234
rect 253 233 254 234
rect 252 233 253 234
rect 251 233 252 234
rect 250 233 251 234
rect 249 233 250 234
rect 248 233 249 234
rect 247 233 248 234
rect 246 233 247 234
rect 245 233 246 234
rect 244 233 245 234
rect 243 233 244 234
rect 242 233 243 234
rect 241 233 242 234
rect 240 233 241 234
rect 239 233 240 234
rect 238 233 239 234
rect 237 233 238 234
rect 236 233 237 234
rect 235 233 236 234
rect 234 233 235 234
rect 233 233 234 234
rect 232 233 233 234
rect 231 233 232 234
rect 230 233 231 234
rect 229 233 230 234
rect 228 233 229 234
rect 227 233 228 234
rect 226 233 227 234
rect 225 233 226 234
rect 224 233 225 234
rect 223 233 224 234
rect 222 233 223 234
rect 221 233 222 234
rect 220 233 221 234
rect 219 233 220 234
rect 218 233 219 234
rect 217 233 218 234
rect 216 233 217 234
rect 215 233 216 234
rect 214 233 215 234
rect 213 233 214 234
rect 212 233 213 234
rect 211 233 212 234
rect 210 233 211 234
rect 209 233 210 234
rect 208 233 209 234
rect 207 233 208 234
rect 206 233 207 234
rect 205 233 206 234
rect 204 233 205 234
rect 203 233 204 234
rect 202 233 203 234
rect 201 233 202 234
rect 200 233 201 234
rect 199 233 200 234
rect 198 233 199 234
rect 197 233 198 234
rect 196 233 197 234
rect 195 233 196 234
rect 194 233 195 234
rect 193 233 194 234
rect 192 233 193 234
rect 191 233 192 234
rect 190 233 191 234
rect 189 233 190 234
rect 188 233 189 234
rect 187 233 188 234
rect 186 233 187 234
rect 185 233 186 234
rect 184 233 185 234
rect 183 233 184 234
rect 182 233 183 234
rect 181 233 182 234
rect 180 233 181 234
rect 179 233 180 234
rect 178 233 179 234
rect 177 233 178 234
rect 176 233 177 234
rect 175 233 176 234
rect 174 233 175 234
rect 173 233 174 234
rect 172 233 173 234
rect 171 233 172 234
rect 170 233 171 234
rect 169 233 170 234
rect 168 233 169 234
rect 167 233 168 234
rect 166 233 167 234
rect 147 233 148 234
rect 146 233 147 234
rect 145 233 146 234
rect 144 233 145 234
rect 143 233 144 234
rect 142 233 143 234
rect 141 233 142 234
rect 140 233 141 234
rect 139 233 140 234
rect 138 233 139 234
rect 137 233 138 234
rect 136 233 137 234
rect 135 233 136 234
rect 134 233 135 234
rect 133 233 134 234
rect 132 233 133 234
rect 131 233 132 234
rect 130 233 131 234
rect 129 233 130 234
rect 128 233 129 234
rect 127 233 128 234
rect 126 233 127 234
rect 125 233 126 234
rect 124 233 125 234
rect 123 233 124 234
rect 122 233 123 234
rect 121 233 122 234
rect 120 233 121 234
rect 119 233 120 234
rect 118 233 119 234
rect 117 233 118 234
rect 116 233 117 234
rect 89 233 90 234
rect 88 233 89 234
rect 87 233 88 234
rect 86 233 87 234
rect 85 233 86 234
rect 84 233 85 234
rect 83 233 84 234
rect 82 233 83 234
rect 81 233 82 234
rect 80 233 81 234
rect 79 233 80 234
rect 78 233 79 234
rect 77 233 78 234
rect 76 233 77 234
rect 75 233 76 234
rect 74 233 75 234
rect 73 233 74 234
rect 72 233 73 234
rect 71 233 72 234
rect 70 233 71 234
rect 69 233 70 234
rect 68 233 69 234
rect 67 233 68 234
rect 66 233 67 234
rect 65 233 66 234
rect 64 233 65 234
rect 63 233 64 234
rect 62 233 63 234
rect 61 233 62 234
rect 60 233 61 234
rect 59 233 60 234
rect 58 233 59 234
rect 57 233 58 234
rect 56 233 57 234
rect 55 233 56 234
rect 54 233 55 234
rect 53 233 54 234
rect 52 233 53 234
rect 51 233 52 234
rect 50 233 51 234
rect 49 233 50 234
rect 48 233 49 234
rect 47 233 48 234
rect 46 233 47 234
rect 45 233 46 234
rect 44 233 45 234
rect 43 233 44 234
rect 42 233 43 234
rect 41 233 42 234
rect 40 233 41 234
rect 39 233 40 234
rect 38 233 39 234
rect 37 233 38 234
rect 36 233 37 234
rect 35 233 36 234
rect 34 233 35 234
rect 33 233 34 234
rect 32 233 33 234
rect 31 233 32 234
rect 30 233 31 234
rect 29 233 30 234
rect 28 233 29 234
rect 27 233 28 234
rect 26 233 27 234
rect 25 233 26 234
rect 24 233 25 234
rect 23 233 24 234
rect 22 233 23 234
rect 21 233 22 234
rect 20 233 21 234
rect 19 233 20 234
rect 18 233 19 234
rect 17 233 18 234
rect 16 233 17 234
rect 15 233 16 234
rect 14 233 15 234
rect 13 233 14 234
rect 12 233 13 234
rect 11 233 12 234
rect 10 233 11 234
rect 9 233 10 234
rect 8 233 9 234
rect 7 233 8 234
rect 482 234 483 235
rect 481 234 482 235
rect 480 234 481 235
rect 479 234 480 235
rect 478 234 479 235
rect 470 234 471 235
rect 469 234 470 235
rect 468 234 469 235
rect 467 234 468 235
rect 466 234 467 235
rect 465 234 466 235
rect 464 234 465 235
rect 442 234 443 235
rect 441 234 442 235
rect 440 234 441 235
rect 422 234 423 235
rect 421 234 422 235
rect 420 234 421 235
rect 398 234 399 235
rect 397 234 398 235
rect 396 234 397 235
rect 277 234 278 235
rect 276 234 277 235
rect 275 234 276 235
rect 274 234 275 235
rect 273 234 274 235
rect 272 234 273 235
rect 271 234 272 235
rect 270 234 271 235
rect 269 234 270 235
rect 268 234 269 235
rect 267 234 268 235
rect 266 234 267 235
rect 265 234 266 235
rect 264 234 265 235
rect 263 234 264 235
rect 262 234 263 235
rect 261 234 262 235
rect 260 234 261 235
rect 259 234 260 235
rect 258 234 259 235
rect 257 234 258 235
rect 256 234 257 235
rect 255 234 256 235
rect 254 234 255 235
rect 253 234 254 235
rect 252 234 253 235
rect 251 234 252 235
rect 250 234 251 235
rect 249 234 250 235
rect 248 234 249 235
rect 247 234 248 235
rect 246 234 247 235
rect 245 234 246 235
rect 244 234 245 235
rect 243 234 244 235
rect 242 234 243 235
rect 241 234 242 235
rect 240 234 241 235
rect 239 234 240 235
rect 238 234 239 235
rect 237 234 238 235
rect 236 234 237 235
rect 235 234 236 235
rect 234 234 235 235
rect 233 234 234 235
rect 232 234 233 235
rect 231 234 232 235
rect 230 234 231 235
rect 229 234 230 235
rect 228 234 229 235
rect 227 234 228 235
rect 226 234 227 235
rect 225 234 226 235
rect 224 234 225 235
rect 223 234 224 235
rect 222 234 223 235
rect 221 234 222 235
rect 220 234 221 235
rect 219 234 220 235
rect 218 234 219 235
rect 217 234 218 235
rect 216 234 217 235
rect 215 234 216 235
rect 214 234 215 235
rect 213 234 214 235
rect 212 234 213 235
rect 211 234 212 235
rect 210 234 211 235
rect 209 234 210 235
rect 208 234 209 235
rect 207 234 208 235
rect 206 234 207 235
rect 205 234 206 235
rect 204 234 205 235
rect 203 234 204 235
rect 202 234 203 235
rect 201 234 202 235
rect 200 234 201 235
rect 199 234 200 235
rect 198 234 199 235
rect 197 234 198 235
rect 196 234 197 235
rect 195 234 196 235
rect 194 234 195 235
rect 193 234 194 235
rect 192 234 193 235
rect 191 234 192 235
rect 190 234 191 235
rect 189 234 190 235
rect 188 234 189 235
rect 187 234 188 235
rect 186 234 187 235
rect 185 234 186 235
rect 184 234 185 235
rect 183 234 184 235
rect 182 234 183 235
rect 181 234 182 235
rect 180 234 181 235
rect 179 234 180 235
rect 178 234 179 235
rect 177 234 178 235
rect 176 234 177 235
rect 175 234 176 235
rect 174 234 175 235
rect 173 234 174 235
rect 172 234 173 235
rect 171 234 172 235
rect 170 234 171 235
rect 169 234 170 235
rect 168 234 169 235
rect 167 234 168 235
rect 147 234 148 235
rect 146 234 147 235
rect 145 234 146 235
rect 144 234 145 235
rect 143 234 144 235
rect 142 234 143 235
rect 141 234 142 235
rect 140 234 141 235
rect 139 234 140 235
rect 138 234 139 235
rect 137 234 138 235
rect 136 234 137 235
rect 135 234 136 235
rect 134 234 135 235
rect 133 234 134 235
rect 132 234 133 235
rect 131 234 132 235
rect 130 234 131 235
rect 129 234 130 235
rect 128 234 129 235
rect 127 234 128 235
rect 126 234 127 235
rect 125 234 126 235
rect 124 234 125 235
rect 123 234 124 235
rect 122 234 123 235
rect 121 234 122 235
rect 120 234 121 235
rect 119 234 120 235
rect 118 234 119 235
rect 117 234 118 235
rect 91 234 92 235
rect 90 234 91 235
rect 89 234 90 235
rect 88 234 89 235
rect 87 234 88 235
rect 86 234 87 235
rect 85 234 86 235
rect 84 234 85 235
rect 83 234 84 235
rect 82 234 83 235
rect 81 234 82 235
rect 80 234 81 235
rect 79 234 80 235
rect 78 234 79 235
rect 77 234 78 235
rect 76 234 77 235
rect 75 234 76 235
rect 74 234 75 235
rect 73 234 74 235
rect 72 234 73 235
rect 71 234 72 235
rect 70 234 71 235
rect 69 234 70 235
rect 68 234 69 235
rect 67 234 68 235
rect 66 234 67 235
rect 65 234 66 235
rect 64 234 65 235
rect 63 234 64 235
rect 62 234 63 235
rect 61 234 62 235
rect 60 234 61 235
rect 59 234 60 235
rect 58 234 59 235
rect 57 234 58 235
rect 56 234 57 235
rect 55 234 56 235
rect 54 234 55 235
rect 53 234 54 235
rect 52 234 53 235
rect 51 234 52 235
rect 50 234 51 235
rect 49 234 50 235
rect 48 234 49 235
rect 47 234 48 235
rect 46 234 47 235
rect 45 234 46 235
rect 44 234 45 235
rect 43 234 44 235
rect 42 234 43 235
rect 41 234 42 235
rect 40 234 41 235
rect 39 234 40 235
rect 38 234 39 235
rect 37 234 38 235
rect 36 234 37 235
rect 35 234 36 235
rect 34 234 35 235
rect 33 234 34 235
rect 32 234 33 235
rect 31 234 32 235
rect 30 234 31 235
rect 29 234 30 235
rect 28 234 29 235
rect 25 234 26 235
rect 24 234 25 235
rect 23 234 24 235
rect 22 234 23 235
rect 21 234 22 235
rect 20 234 21 235
rect 19 234 20 235
rect 18 234 19 235
rect 17 234 18 235
rect 16 234 17 235
rect 15 234 16 235
rect 14 234 15 235
rect 13 234 14 235
rect 12 234 13 235
rect 11 234 12 235
rect 10 234 11 235
rect 9 234 10 235
rect 8 234 9 235
rect 7 234 8 235
rect 6 234 7 235
rect 483 235 484 236
rect 482 235 483 236
rect 481 235 482 236
rect 480 235 481 236
rect 442 235 443 236
rect 441 235 442 236
rect 440 235 441 236
rect 422 235 423 236
rect 421 235 422 236
rect 420 235 421 236
rect 398 235 399 236
rect 397 235 398 236
rect 396 235 397 236
rect 276 235 277 236
rect 275 235 276 236
rect 274 235 275 236
rect 273 235 274 236
rect 272 235 273 236
rect 271 235 272 236
rect 270 235 271 236
rect 269 235 270 236
rect 268 235 269 236
rect 267 235 268 236
rect 266 235 267 236
rect 265 235 266 236
rect 264 235 265 236
rect 263 235 264 236
rect 262 235 263 236
rect 261 235 262 236
rect 260 235 261 236
rect 259 235 260 236
rect 258 235 259 236
rect 257 235 258 236
rect 256 235 257 236
rect 255 235 256 236
rect 254 235 255 236
rect 253 235 254 236
rect 252 235 253 236
rect 251 235 252 236
rect 250 235 251 236
rect 249 235 250 236
rect 248 235 249 236
rect 247 235 248 236
rect 246 235 247 236
rect 245 235 246 236
rect 244 235 245 236
rect 243 235 244 236
rect 242 235 243 236
rect 241 235 242 236
rect 240 235 241 236
rect 239 235 240 236
rect 238 235 239 236
rect 237 235 238 236
rect 236 235 237 236
rect 235 235 236 236
rect 234 235 235 236
rect 233 235 234 236
rect 232 235 233 236
rect 231 235 232 236
rect 230 235 231 236
rect 229 235 230 236
rect 228 235 229 236
rect 227 235 228 236
rect 226 235 227 236
rect 225 235 226 236
rect 224 235 225 236
rect 223 235 224 236
rect 222 235 223 236
rect 221 235 222 236
rect 220 235 221 236
rect 219 235 220 236
rect 218 235 219 236
rect 217 235 218 236
rect 216 235 217 236
rect 215 235 216 236
rect 214 235 215 236
rect 213 235 214 236
rect 212 235 213 236
rect 211 235 212 236
rect 210 235 211 236
rect 209 235 210 236
rect 208 235 209 236
rect 207 235 208 236
rect 206 235 207 236
rect 205 235 206 236
rect 204 235 205 236
rect 203 235 204 236
rect 202 235 203 236
rect 201 235 202 236
rect 200 235 201 236
rect 199 235 200 236
rect 198 235 199 236
rect 197 235 198 236
rect 196 235 197 236
rect 195 235 196 236
rect 194 235 195 236
rect 193 235 194 236
rect 192 235 193 236
rect 191 235 192 236
rect 190 235 191 236
rect 189 235 190 236
rect 188 235 189 236
rect 187 235 188 236
rect 186 235 187 236
rect 185 235 186 236
rect 184 235 185 236
rect 183 235 184 236
rect 182 235 183 236
rect 181 235 182 236
rect 180 235 181 236
rect 179 235 180 236
rect 178 235 179 236
rect 177 235 178 236
rect 176 235 177 236
rect 175 235 176 236
rect 174 235 175 236
rect 173 235 174 236
rect 172 235 173 236
rect 171 235 172 236
rect 170 235 171 236
rect 169 235 170 236
rect 147 235 148 236
rect 146 235 147 236
rect 145 235 146 236
rect 144 235 145 236
rect 143 235 144 236
rect 142 235 143 236
rect 141 235 142 236
rect 140 235 141 236
rect 139 235 140 236
rect 138 235 139 236
rect 137 235 138 236
rect 136 235 137 236
rect 135 235 136 236
rect 134 235 135 236
rect 133 235 134 236
rect 132 235 133 236
rect 131 235 132 236
rect 130 235 131 236
rect 129 235 130 236
rect 128 235 129 236
rect 127 235 128 236
rect 126 235 127 236
rect 125 235 126 236
rect 124 235 125 236
rect 123 235 124 236
rect 122 235 123 236
rect 121 235 122 236
rect 120 235 121 236
rect 119 235 120 236
rect 118 235 119 236
rect 94 235 95 236
rect 93 235 94 236
rect 92 235 93 236
rect 91 235 92 236
rect 90 235 91 236
rect 89 235 90 236
rect 88 235 89 236
rect 87 235 88 236
rect 86 235 87 236
rect 85 235 86 236
rect 84 235 85 236
rect 83 235 84 236
rect 82 235 83 236
rect 81 235 82 236
rect 80 235 81 236
rect 79 235 80 236
rect 78 235 79 236
rect 77 235 78 236
rect 76 235 77 236
rect 75 235 76 236
rect 74 235 75 236
rect 73 235 74 236
rect 72 235 73 236
rect 71 235 72 236
rect 70 235 71 236
rect 69 235 70 236
rect 68 235 69 236
rect 67 235 68 236
rect 66 235 67 236
rect 65 235 66 236
rect 64 235 65 236
rect 63 235 64 236
rect 62 235 63 236
rect 61 235 62 236
rect 60 235 61 236
rect 59 235 60 236
rect 58 235 59 236
rect 57 235 58 236
rect 56 235 57 236
rect 55 235 56 236
rect 54 235 55 236
rect 53 235 54 236
rect 52 235 53 236
rect 51 235 52 236
rect 50 235 51 236
rect 49 235 50 236
rect 48 235 49 236
rect 47 235 48 236
rect 46 235 47 236
rect 45 235 46 236
rect 44 235 45 236
rect 43 235 44 236
rect 42 235 43 236
rect 41 235 42 236
rect 40 235 41 236
rect 39 235 40 236
rect 38 235 39 236
rect 37 235 38 236
rect 36 235 37 236
rect 35 235 36 236
rect 34 235 35 236
rect 33 235 34 236
rect 32 235 33 236
rect 31 235 32 236
rect 30 235 31 236
rect 29 235 30 236
rect 28 235 29 236
rect 24 235 25 236
rect 23 235 24 236
rect 22 235 23 236
rect 21 235 22 236
rect 20 235 21 236
rect 19 235 20 236
rect 18 235 19 236
rect 17 235 18 236
rect 16 235 17 236
rect 15 235 16 236
rect 14 235 15 236
rect 13 235 14 236
rect 12 235 13 236
rect 11 235 12 236
rect 10 235 11 236
rect 9 235 10 236
rect 8 235 9 236
rect 7 235 8 236
rect 6 235 7 236
rect 483 236 484 237
rect 482 236 483 237
rect 481 236 482 237
rect 442 236 443 237
rect 441 236 442 237
rect 440 236 441 237
rect 422 236 423 237
rect 421 236 422 237
rect 420 236 421 237
rect 398 236 399 237
rect 397 236 398 237
rect 396 236 397 237
rect 275 236 276 237
rect 274 236 275 237
rect 273 236 274 237
rect 272 236 273 237
rect 271 236 272 237
rect 270 236 271 237
rect 269 236 270 237
rect 268 236 269 237
rect 267 236 268 237
rect 266 236 267 237
rect 265 236 266 237
rect 264 236 265 237
rect 263 236 264 237
rect 262 236 263 237
rect 261 236 262 237
rect 260 236 261 237
rect 259 236 260 237
rect 258 236 259 237
rect 257 236 258 237
rect 256 236 257 237
rect 255 236 256 237
rect 254 236 255 237
rect 253 236 254 237
rect 252 236 253 237
rect 251 236 252 237
rect 250 236 251 237
rect 249 236 250 237
rect 248 236 249 237
rect 247 236 248 237
rect 246 236 247 237
rect 245 236 246 237
rect 244 236 245 237
rect 243 236 244 237
rect 242 236 243 237
rect 241 236 242 237
rect 240 236 241 237
rect 239 236 240 237
rect 238 236 239 237
rect 237 236 238 237
rect 236 236 237 237
rect 235 236 236 237
rect 234 236 235 237
rect 233 236 234 237
rect 232 236 233 237
rect 231 236 232 237
rect 230 236 231 237
rect 229 236 230 237
rect 228 236 229 237
rect 227 236 228 237
rect 226 236 227 237
rect 225 236 226 237
rect 224 236 225 237
rect 223 236 224 237
rect 222 236 223 237
rect 221 236 222 237
rect 220 236 221 237
rect 219 236 220 237
rect 218 236 219 237
rect 217 236 218 237
rect 216 236 217 237
rect 215 236 216 237
rect 214 236 215 237
rect 213 236 214 237
rect 212 236 213 237
rect 211 236 212 237
rect 210 236 211 237
rect 209 236 210 237
rect 208 236 209 237
rect 207 236 208 237
rect 206 236 207 237
rect 205 236 206 237
rect 204 236 205 237
rect 203 236 204 237
rect 202 236 203 237
rect 201 236 202 237
rect 200 236 201 237
rect 199 236 200 237
rect 198 236 199 237
rect 197 236 198 237
rect 196 236 197 237
rect 195 236 196 237
rect 194 236 195 237
rect 193 236 194 237
rect 192 236 193 237
rect 191 236 192 237
rect 190 236 191 237
rect 189 236 190 237
rect 188 236 189 237
rect 187 236 188 237
rect 186 236 187 237
rect 185 236 186 237
rect 184 236 185 237
rect 183 236 184 237
rect 182 236 183 237
rect 181 236 182 237
rect 180 236 181 237
rect 179 236 180 237
rect 178 236 179 237
rect 177 236 178 237
rect 176 236 177 237
rect 175 236 176 237
rect 174 236 175 237
rect 173 236 174 237
rect 172 236 173 237
rect 171 236 172 237
rect 170 236 171 237
rect 148 236 149 237
rect 147 236 148 237
rect 146 236 147 237
rect 145 236 146 237
rect 144 236 145 237
rect 143 236 144 237
rect 142 236 143 237
rect 141 236 142 237
rect 140 236 141 237
rect 139 236 140 237
rect 138 236 139 237
rect 137 236 138 237
rect 136 236 137 237
rect 135 236 136 237
rect 134 236 135 237
rect 133 236 134 237
rect 132 236 133 237
rect 131 236 132 237
rect 130 236 131 237
rect 129 236 130 237
rect 128 236 129 237
rect 127 236 128 237
rect 126 236 127 237
rect 125 236 126 237
rect 124 236 125 237
rect 123 236 124 237
rect 122 236 123 237
rect 121 236 122 237
rect 120 236 121 237
rect 119 236 120 237
rect 118 236 119 237
rect 96 236 97 237
rect 95 236 96 237
rect 94 236 95 237
rect 93 236 94 237
rect 92 236 93 237
rect 91 236 92 237
rect 90 236 91 237
rect 89 236 90 237
rect 88 236 89 237
rect 87 236 88 237
rect 86 236 87 237
rect 85 236 86 237
rect 84 236 85 237
rect 83 236 84 237
rect 82 236 83 237
rect 81 236 82 237
rect 80 236 81 237
rect 79 236 80 237
rect 78 236 79 237
rect 77 236 78 237
rect 76 236 77 237
rect 75 236 76 237
rect 74 236 75 237
rect 73 236 74 237
rect 72 236 73 237
rect 71 236 72 237
rect 70 236 71 237
rect 69 236 70 237
rect 68 236 69 237
rect 67 236 68 237
rect 66 236 67 237
rect 65 236 66 237
rect 64 236 65 237
rect 63 236 64 237
rect 62 236 63 237
rect 61 236 62 237
rect 60 236 61 237
rect 59 236 60 237
rect 58 236 59 237
rect 57 236 58 237
rect 56 236 57 237
rect 55 236 56 237
rect 54 236 55 237
rect 53 236 54 237
rect 52 236 53 237
rect 51 236 52 237
rect 50 236 51 237
rect 49 236 50 237
rect 48 236 49 237
rect 47 236 48 237
rect 46 236 47 237
rect 45 236 46 237
rect 44 236 45 237
rect 43 236 44 237
rect 42 236 43 237
rect 41 236 42 237
rect 40 236 41 237
rect 39 236 40 237
rect 38 236 39 237
rect 37 236 38 237
rect 36 236 37 237
rect 35 236 36 237
rect 34 236 35 237
rect 33 236 34 237
rect 32 236 33 237
rect 31 236 32 237
rect 30 236 31 237
rect 29 236 30 237
rect 24 236 25 237
rect 23 236 24 237
rect 22 236 23 237
rect 21 236 22 237
rect 20 236 21 237
rect 19 236 20 237
rect 18 236 19 237
rect 17 236 18 237
rect 16 236 17 237
rect 15 236 16 237
rect 14 236 15 237
rect 13 236 14 237
rect 12 236 13 237
rect 11 236 12 237
rect 10 236 11 237
rect 9 236 10 237
rect 8 236 9 237
rect 7 236 8 237
rect 6 236 7 237
rect 483 237 484 238
rect 482 237 483 238
rect 442 237 443 238
rect 441 237 442 238
rect 440 237 441 238
rect 423 237 424 238
rect 422 237 423 238
rect 421 237 422 238
rect 420 237 421 238
rect 398 237 399 238
rect 397 237 398 238
rect 396 237 397 238
rect 274 237 275 238
rect 273 237 274 238
rect 272 237 273 238
rect 271 237 272 238
rect 270 237 271 238
rect 269 237 270 238
rect 268 237 269 238
rect 267 237 268 238
rect 266 237 267 238
rect 265 237 266 238
rect 264 237 265 238
rect 263 237 264 238
rect 262 237 263 238
rect 261 237 262 238
rect 260 237 261 238
rect 259 237 260 238
rect 258 237 259 238
rect 257 237 258 238
rect 256 237 257 238
rect 255 237 256 238
rect 254 237 255 238
rect 253 237 254 238
rect 252 237 253 238
rect 251 237 252 238
rect 250 237 251 238
rect 249 237 250 238
rect 248 237 249 238
rect 247 237 248 238
rect 246 237 247 238
rect 245 237 246 238
rect 244 237 245 238
rect 243 237 244 238
rect 242 237 243 238
rect 241 237 242 238
rect 240 237 241 238
rect 239 237 240 238
rect 238 237 239 238
rect 237 237 238 238
rect 236 237 237 238
rect 235 237 236 238
rect 234 237 235 238
rect 233 237 234 238
rect 232 237 233 238
rect 231 237 232 238
rect 230 237 231 238
rect 229 237 230 238
rect 228 237 229 238
rect 227 237 228 238
rect 226 237 227 238
rect 225 237 226 238
rect 224 237 225 238
rect 223 237 224 238
rect 222 237 223 238
rect 221 237 222 238
rect 220 237 221 238
rect 219 237 220 238
rect 218 237 219 238
rect 217 237 218 238
rect 216 237 217 238
rect 215 237 216 238
rect 214 237 215 238
rect 213 237 214 238
rect 212 237 213 238
rect 211 237 212 238
rect 210 237 211 238
rect 209 237 210 238
rect 208 237 209 238
rect 207 237 208 238
rect 206 237 207 238
rect 205 237 206 238
rect 204 237 205 238
rect 203 237 204 238
rect 202 237 203 238
rect 201 237 202 238
rect 200 237 201 238
rect 199 237 200 238
rect 198 237 199 238
rect 197 237 198 238
rect 196 237 197 238
rect 195 237 196 238
rect 194 237 195 238
rect 193 237 194 238
rect 192 237 193 238
rect 191 237 192 238
rect 190 237 191 238
rect 189 237 190 238
rect 188 237 189 238
rect 187 237 188 238
rect 186 237 187 238
rect 185 237 186 238
rect 184 237 185 238
rect 183 237 184 238
rect 182 237 183 238
rect 181 237 182 238
rect 180 237 181 238
rect 179 237 180 238
rect 178 237 179 238
rect 177 237 178 238
rect 176 237 177 238
rect 175 237 176 238
rect 174 237 175 238
rect 173 237 174 238
rect 172 237 173 238
rect 148 237 149 238
rect 147 237 148 238
rect 146 237 147 238
rect 145 237 146 238
rect 144 237 145 238
rect 143 237 144 238
rect 142 237 143 238
rect 141 237 142 238
rect 140 237 141 238
rect 139 237 140 238
rect 138 237 139 238
rect 137 237 138 238
rect 136 237 137 238
rect 135 237 136 238
rect 134 237 135 238
rect 133 237 134 238
rect 132 237 133 238
rect 131 237 132 238
rect 130 237 131 238
rect 129 237 130 238
rect 128 237 129 238
rect 127 237 128 238
rect 126 237 127 238
rect 125 237 126 238
rect 124 237 125 238
rect 123 237 124 238
rect 122 237 123 238
rect 121 237 122 238
rect 120 237 121 238
rect 119 237 120 238
rect 98 237 99 238
rect 97 237 98 238
rect 96 237 97 238
rect 95 237 96 238
rect 94 237 95 238
rect 93 237 94 238
rect 92 237 93 238
rect 91 237 92 238
rect 90 237 91 238
rect 89 237 90 238
rect 88 237 89 238
rect 87 237 88 238
rect 86 237 87 238
rect 85 237 86 238
rect 84 237 85 238
rect 83 237 84 238
rect 82 237 83 238
rect 81 237 82 238
rect 80 237 81 238
rect 79 237 80 238
rect 78 237 79 238
rect 77 237 78 238
rect 76 237 77 238
rect 75 237 76 238
rect 74 237 75 238
rect 73 237 74 238
rect 72 237 73 238
rect 71 237 72 238
rect 70 237 71 238
rect 69 237 70 238
rect 68 237 69 238
rect 67 237 68 238
rect 66 237 67 238
rect 65 237 66 238
rect 64 237 65 238
rect 63 237 64 238
rect 62 237 63 238
rect 61 237 62 238
rect 60 237 61 238
rect 59 237 60 238
rect 58 237 59 238
rect 57 237 58 238
rect 56 237 57 238
rect 55 237 56 238
rect 54 237 55 238
rect 53 237 54 238
rect 52 237 53 238
rect 51 237 52 238
rect 50 237 51 238
rect 49 237 50 238
rect 48 237 49 238
rect 47 237 48 238
rect 46 237 47 238
rect 45 237 46 238
rect 44 237 45 238
rect 43 237 44 238
rect 42 237 43 238
rect 41 237 42 238
rect 40 237 41 238
rect 39 237 40 238
rect 38 237 39 238
rect 37 237 38 238
rect 36 237 37 238
rect 35 237 36 238
rect 34 237 35 238
rect 33 237 34 238
rect 32 237 33 238
rect 31 237 32 238
rect 30 237 31 238
rect 29 237 30 238
rect 24 237 25 238
rect 23 237 24 238
rect 22 237 23 238
rect 21 237 22 238
rect 20 237 21 238
rect 19 237 20 238
rect 18 237 19 238
rect 17 237 18 238
rect 16 237 17 238
rect 15 237 16 238
rect 14 237 15 238
rect 13 237 14 238
rect 12 237 13 238
rect 11 237 12 238
rect 10 237 11 238
rect 9 237 10 238
rect 8 237 9 238
rect 7 237 8 238
rect 6 237 7 238
rect 442 238 443 239
rect 441 238 442 239
rect 440 238 441 239
rect 423 238 424 239
rect 422 238 423 239
rect 421 238 422 239
rect 420 238 421 239
rect 398 238 399 239
rect 397 238 398 239
rect 396 238 397 239
rect 273 238 274 239
rect 272 238 273 239
rect 271 238 272 239
rect 270 238 271 239
rect 269 238 270 239
rect 268 238 269 239
rect 267 238 268 239
rect 266 238 267 239
rect 265 238 266 239
rect 264 238 265 239
rect 263 238 264 239
rect 262 238 263 239
rect 261 238 262 239
rect 260 238 261 239
rect 259 238 260 239
rect 258 238 259 239
rect 257 238 258 239
rect 256 238 257 239
rect 255 238 256 239
rect 254 238 255 239
rect 253 238 254 239
rect 252 238 253 239
rect 251 238 252 239
rect 250 238 251 239
rect 249 238 250 239
rect 248 238 249 239
rect 247 238 248 239
rect 246 238 247 239
rect 245 238 246 239
rect 244 238 245 239
rect 243 238 244 239
rect 242 238 243 239
rect 241 238 242 239
rect 240 238 241 239
rect 239 238 240 239
rect 238 238 239 239
rect 237 238 238 239
rect 236 238 237 239
rect 235 238 236 239
rect 234 238 235 239
rect 233 238 234 239
rect 232 238 233 239
rect 231 238 232 239
rect 230 238 231 239
rect 229 238 230 239
rect 228 238 229 239
rect 227 238 228 239
rect 226 238 227 239
rect 225 238 226 239
rect 224 238 225 239
rect 223 238 224 239
rect 222 238 223 239
rect 221 238 222 239
rect 220 238 221 239
rect 219 238 220 239
rect 218 238 219 239
rect 217 238 218 239
rect 216 238 217 239
rect 215 238 216 239
rect 214 238 215 239
rect 213 238 214 239
rect 212 238 213 239
rect 211 238 212 239
rect 210 238 211 239
rect 209 238 210 239
rect 208 238 209 239
rect 207 238 208 239
rect 206 238 207 239
rect 205 238 206 239
rect 204 238 205 239
rect 203 238 204 239
rect 202 238 203 239
rect 201 238 202 239
rect 200 238 201 239
rect 199 238 200 239
rect 198 238 199 239
rect 197 238 198 239
rect 196 238 197 239
rect 195 238 196 239
rect 194 238 195 239
rect 193 238 194 239
rect 192 238 193 239
rect 191 238 192 239
rect 190 238 191 239
rect 189 238 190 239
rect 188 238 189 239
rect 187 238 188 239
rect 186 238 187 239
rect 185 238 186 239
rect 184 238 185 239
rect 183 238 184 239
rect 182 238 183 239
rect 181 238 182 239
rect 180 238 181 239
rect 179 238 180 239
rect 178 238 179 239
rect 177 238 178 239
rect 176 238 177 239
rect 175 238 176 239
rect 174 238 175 239
rect 173 238 174 239
rect 149 238 150 239
rect 148 238 149 239
rect 147 238 148 239
rect 146 238 147 239
rect 145 238 146 239
rect 144 238 145 239
rect 143 238 144 239
rect 142 238 143 239
rect 141 238 142 239
rect 140 238 141 239
rect 139 238 140 239
rect 138 238 139 239
rect 137 238 138 239
rect 136 238 137 239
rect 135 238 136 239
rect 134 238 135 239
rect 133 238 134 239
rect 132 238 133 239
rect 131 238 132 239
rect 130 238 131 239
rect 129 238 130 239
rect 128 238 129 239
rect 127 238 128 239
rect 126 238 127 239
rect 125 238 126 239
rect 124 238 125 239
rect 123 238 124 239
rect 122 238 123 239
rect 121 238 122 239
rect 120 238 121 239
rect 119 238 120 239
rect 99 238 100 239
rect 98 238 99 239
rect 97 238 98 239
rect 96 238 97 239
rect 95 238 96 239
rect 94 238 95 239
rect 93 238 94 239
rect 92 238 93 239
rect 91 238 92 239
rect 90 238 91 239
rect 89 238 90 239
rect 88 238 89 239
rect 87 238 88 239
rect 86 238 87 239
rect 85 238 86 239
rect 84 238 85 239
rect 83 238 84 239
rect 82 238 83 239
rect 81 238 82 239
rect 80 238 81 239
rect 79 238 80 239
rect 78 238 79 239
rect 77 238 78 239
rect 76 238 77 239
rect 75 238 76 239
rect 74 238 75 239
rect 73 238 74 239
rect 72 238 73 239
rect 71 238 72 239
rect 70 238 71 239
rect 69 238 70 239
rect 68 238 69 239
rect 67 238 68 239
rect 66 238 67 239
rect 65 238 66 239
rect 64 238 65 239
rect 63 238 64 239
rect 62 238 63 239
rect 61 238 62 239
rect 60 238 61 239
rect 59 238 60 239
rect 58 238 59 239
rect 57 238 58 239
rect 56 238 57 239
rect 55 238 56 239
rect 54 238 55 239
rect 53 238 54 239
rect 52 238 53 239
rect 51 238 52 239
rect 50 238 51 239
rect 49 238 50 239
rect 48 238 49 239
rect 47 238 48 239
rect 46 238 47 239
rect 45 238 46 239
rect 44 238 45 239
rect 43 238 44 239
rect 42 238 43 239
rect 41 238 42 239
rect 40 238 41 239
rect 39 238 40 239
rect 38 238 39 239
rect 37 238 38 239
rect 36 238 37 239
rect 35 238 36 239
rect 34 238 35 239
rect 33 238 34 239
rect 32 238 33 239
rect 31 238 32 239
rect 30 238 31 239
rect 29 238 30 239
rect 23 238 24 239
rect 22 238 23 239
rect 21 238 22 239
rect 20 238 21 239
rect 19 238 20 239
rect 18 238 19 239
rect 17 238 18 239
rect 16 238 17 239
rect 15 238 16 239
rect 14 238 15 239
rect 13 238 14 239
rect 12 238 13 239
rect 11 238 12 239
rect 10 238 11 239
rect 9 238 10 239
rect 8 238 9 239
rect 7 238 8 239
rect 6 238 7 239
rect 442 239 443 240
rect 441 239 442 240
rect 440 239 441 240
rect 423 239 424 240
rect 422 239 423 240
rect 421 239 422 240
rect 420 239 421 240
rect 399 239 400 240
rect 398 239 399 240
rect 397 239 398 240
rect 396 239 397 240
rect 273 239 274 240
rect 272 239 273 240
rect 271 239 272 240
rect 270 239 271 240
rect 269 239 270 240
rect 268 239 269 240
rect 267 239 268 240
rect 266 239 267 240
rect 265 239 266 240
rect 264 239 265 240
rect 263 239 264 240
rect 262 239 263 240
rect 261 239 262 240
rect 260 239 261 240
rect 259 239 260 240
rect 258 239 259 240
rect 257 239 258 240
rect 256 239 257 240
rect 255 239 256 240
rect 254 239 255 240
rect 253 239 254 240
rect 252 239 253 240
rect 251 239 252 240
rect 250 239 251 240
rect 249 239 250 240
rect 248 239 249 240
rect 247 239 248 240
rect 246 239 247 240
rect 245 239 246 240
rect 244 239 245 240
rect 243 239 244 240
rect 242 239 243 240
rect 241 239 242 240
rect 240 239 241 240
rect 239 239 240 240
rect 238 239 239 240
rect 237 239 238 240
rect 236 239 237 240
rect 235 239 236 240
rect 234 239 235 240
rect 233 239 234 240
rect 232 239 233 240
rect 231 239 232 240
rect 230 239 231 240
rect 229 239 230 240
rect 228 239 229 240
rect 227 239 228 240
rect 226 239 227 240
rect 225 239 226 240
rect 224 239 225 240
rect 223 239 224 240
rect 222 239 223 240
rect 221 239 222 240
rect 220 239 221 240
rect 219 239 220 240
rect 218 239 219 240
rect 217 239 218 240
rect 216 239 217 240
rect 215 239 216 240
rect 214 239 215 240
rect 213 239 214 240
rect 212 239 213 240
rect 211 239 212 240
rect 210 239 211 240
rect 209 239 210 240
rect 208 239 209 240
rect 207 239 208 240
rect 206 239 207 240
rect 205 239 206 240
rect 204 239 205 240
rect 203 239 204 240
rect 202 239 203 240
rect 201 239 202 240
rect 200 239 201 240
rect 199 239 200 240
rect 198 239 199 240
rect 197 239 198 240
rect 196 239 197 240
rect 195 239 196 240
rect 194 239 195 240
rect 193 239 194 240
rect 192 239 193 240
rect 191 239 192 240
rect 190 239 191 240
rect 189 239 190 240
rect 188 239 189 240
rect 187 239 188 240
rect 186 239 187 240
rect 185 239 186 240
rect 184 239 185 240
rect 183 239 184 240
rect 182 239 183 240
rect 181 239 182 240
rect 180 239 181 240
rect 179 239 180 240
rect 178 239 179 240
rect 177 239 178 240
rect 176 239 177 240
rect 175 239 176 240
rect 149 239 150 240
rect 148 239 149 240
rect 147 239 148 240
rect 146 239 147 240
rect 145 239 146 240
rect 144 239 145 240
rect 143 239 144 240
rect 142 239 143 240
rect 141 239 142 240
rect 140 239 141 240
rect 139 239 140 240
rect 138 239 139 240
rect 137 239 138 240
rect 136 239 137 240
rect 135 239 136 240
rect 134 239 135 240
rect 133 239 134 240
rect 132 239 133 240
rect 131 239 132 240
rect 130 239 131 240
rect 129 239 130 240
rect 128 239 129 240
rect 127 239 128 240
rect 126 239 127 240
rect 125 239 126 240
rect 124 239 125 240
rect 123 239 124 240
rect 122 239 123 240
rect 121 239 122 240
rect 120 239 121 240
rect 119 239 120 240
rect 101 239 102 240
rect 100 239 101 240
rect 99 239 100 240
rect 98 239 99 240
rect 97 239 98 240
rect 96 239 97 240
rect 95 239 96 240
rect 94 239 95 240
rect 93 239 94 240
rect 92 239 93 240
rect 91 239 92 240
rect 90 239 91 240
rect 89 239 90 240
rect 88 239 89 240
rect 87 239 88 240
rect 86 239 87 240
rect 85 239 86 240
rect 84 239 85 240
rect 83 239 84 240
rect 82 239 83 240
rect 81 239 82 240
rect 80 239 81 240
rect 79 239 80 240
rect 78 239 79 240
rect 77 239 78 240
rect 76 239 77 240
rect 75 239 76 240
rect 74 239 75 240
rect 73 239 74 240
rect 72 239 73 240
rect 71 239 72 240
rect 70 239 71 240
rect 69 239 70 240
rect 68 239 69 240
rect 67 239 68 240
rect 66 239 67 240
rect 65 239 66 240
rect 64 239 65 240
rect 63 239 64 240
rect 62 239 63 240
rect 61 239 62 240
rect 60 239 61 240
rect 59 239 60 240
rect 58 239 59 240
rect 57 239 58 240
rect 56 239 57 240
rect 55 239 56 240
rect 54 239 55 240
rect 53 239 54 240
rect 52 239 53 240
rect 51 239 52 240
rect 50 239 51 240
rect 49 239 50 240
rect 48 239 49 240
rect 47 239 48 240
rect 46 239 47 240
rect 45 239 46 240
rect 44 239 45 240
rect 43 239 44 240
rect 42 239 43 240
rect 41 239 42 240
rect 40 239 41 240
rect 39 239 40 240
rect 38 239 39 240
rect 37 239 38 240
rect 36 239 37 240
rect 35 239 36 240
rect 34 239 35 240
rect 33 239 34 240
rect 32 239 33 240
rect 31 239 32 240
rect 30 239 31 240
rect 29 239 30 240
rect 23 239 24 240
rect 22 239 23 240
rect 21 239 22 240
rect 20 239 21 240
rect 19 239 20 240
rect 18 239 19 240
rect 17 239 18 240
rect 16 239 17 240
rect 15 239 16 240
rect 14 239 15 240
rect 13 239 14 240
rect 12 239 13 240
rect 11 239 12 240
rect 10 239 11 240
rect 9 239 10 240
rect 8 239 9 240
rect 7 239 8 240
rect 6 239 7 240
rect 442 240 443 241
rect 441 240 442 241
rect 440 240 441 241
rect 439 240 440 241
rect 424 240 425 241
rect 423 240 424 241
rect 422 240 423 241
rect 421 240 422 241
rect 420 240 421 241
rect 399 240 400 241
rect 398 240 399 241
rect 397 240 398 241
rect 396 240 397 241
rect 272 240 273 241
rect 271 240 272 241
rect 270 240 271 241
rect 269 240 270 241
rect 268 240 269 241
rect 267 240 268 241
rect 266 240 267 241
rect 265 240 266 241
rect 264 240 265 241
rect 263 240 264 241
rect 262 240 263 241
rect 261 240 262 241
rect 260 240 261 241
rect 259 240 260 241
rect 258 240 259 241
rect 257 240 258 241
rect 256 240 257 241
rect 255 240 256 241
rect 254 240 255 241
rect 253 240 254 241
rect 252 240 253 241
rect 251 240 252 241
rect 250 240 251 241
rect 249 240 250 241
rect 248 240 249 241
rect 247 240 248 241
rect 246 240 247 241
rect 245 240 246 241
rect 244 240 245 241
rect 243 240 244 241
rect 242 240 243 241
rect 241 240 242 241
rect 240 240 241 241
rect 239 240 240 241
rect 238 240 239 241
rect 237 240 238 241
rect 236 240 237 241
rect 235 240 236 241
rect 234 240 235 241
rect 233 240 234 241
rect 232 240 233 241
rect 231 240 232 241
rect 230 240 231 241
rect 229 240 230 241
rect 228 240 229 241
rect 227 240 228 241
rect 226 240 227 241
rect 225 240 226 241
rect 224 240 225 241
rect 223 240 224 241
rect 222 240 223 241
rect 221 240 222 241
rect 220 240 221 241
rect 219 240 220 241
rect 218 240 219 241
rect 217 240 218 241
rect 216 240 217 241
rect 215 240 216 241
rect 214 240 215 241
rect 213 240 214 241
rect 212 240 213 241
rect 211 240 212 241
rect 210 240 211 241
rect 209 240 210 241
rect 208 240 209 241
rect 207 240 208 241
rect 206 240 207 241
rect 205 240 206 241
rect 204 240 205 241
rect 203 240 204 241
rect 202 240 203 241
rect 201 240 202 241
rect 200 240 201 241
rect 199 240 200 241
rect 198 240 199 241
rect 197 240 198 241
rect 196 240 197 241
rect 195 240 196 241
rect 194 240 195 241
rect 193 240 194 241
rect 192 240 193 241
rect 191 240 192 241
rect 190 240 191 241
rect 189 240 190 241
rect 188 240 189 241
rect 187 240 188 241
rect 186 240 187 241
rect 185 240 186 241
rect 184 240 185 241
rect 183 240 184 241
rect 182 240 183 241
rect 181 240 182 241
rect 180 240 181 241
rect 179 240 180 241
rect 178 240 179 241
rect 177 240 178 241
rect 150 240 151 241
rect 149 240 150 241
rect 148 240 149 241
rect 147 240 148 241
rect 146 240 147 241
rect 145 240 146 241
rect 144 240 145 241
rect 143 240 144 241
rect 142 240 143 241
rect 141 240 142 241
rect 140 240 141 241
rect 139 240 140 241
rect 138 240 139 241
rect 137 240 138 241
rect 136 240 137 241
rect 135 240 136 241
rect 134 240 135 241
rect 133 240 134 241
rect 132 240 133 241
rect 131 240 132 241
rect 130 240 131 241
rect 129 240 130 241
rect 128 240 129 241
rect 127 240 128 241
rect 126 240 127 241
rect 125 240 126 241
rect 124 240 125 241
rect 123 240 124 241
rect 122 240 123 241
rect 121 240 122 241
rect 120 240 121 241
rect 102 240 103 241
rect 101 240 102 241
rect 100 240 101 241
rect 99 240 100 241
rect 98 240 99 241
rect 97 240 98 241
rect 96 240 97 241
rect 95 240 96 241
rect 94 240 95 241
rect 93 240 94 241
rect 92 240 93 241
rect 91 240 92 241
rect 90 240 91 241
rect 89 240 90 241
rect 88 240 89 241
rect 87 240 88 241
rect 86 240 87 241
rect 85 240 86 241
rect 84 240 85 241
rect 83 240 84 241
rect 82 240 83 241
rect 81 240 82 241
rect 80 240 81 241
rect 79 240 80 241
rect 78 240 79 241
rect 77 240 78 241
rect 76 240 77 241
rect 75 240 76 241
rect 74 240 75 241
rect 73 240 74 241
rect 72 240 73 241
rect 71 240 72 241
rect 70 240 71 241
rect 69 240 70 241
rect 68 240 69 241
rect 67 240 68 241
rect 66 240 67 241
rect 65 240 66 241
rect 64 240 65 241
rect 63 240 64 241
rect 62 240 63 241
rect 61 240 62 241
rect 60 240 61 241
rect 59 240 60 241
rect 58 240 59 241
rect 57 240 58 241
rect 56 240 57 241
rect 55 240 56 241
rect 54 240 55 241
rect 53 240 54 241
rect 52 240 53 241
rect 51 240 52 241
rect 50 240 51 241
rect 49 240 50 241
rect 48 240 49 241
rect 47 240 48 241
rect 46 240 47 241
rect 45 240 46 241
rect 44 240 45 241
rect 43 240 44 241
rect 42 240 43 241
rect 41 240 42 241
rect 40 240 41 241
rect 39 240 40 241
rect 38 240 39 241
rect 37 240 38 241
rect 36 240 37 241
rect 35 240 36 241
rect 34 240 35 241
rect 33 240 34 241
rect 32 240 33 241
rect 31 240 32 241
rect 30 240 31 241
rect 29 240 30 241
rect 23 240 24 241
rect 22 240 23 241
rect 21 240 22 241
rect 20 240 21 241
rect 19 240 20 241
rect 18 240 19 241
rect 17 240 18 241
rect 16 240 17 241
rect 15 240 16 241
rect 14 240 15 241
rect 13 240 14 241
rect 12 240 13 241
rect 11 240 12 241
rect 10 240 11 241
rect 9 240 10 241
rect 8 240 9 241
rect 7 240 8 241
rect 6 240 7 241
rect 442 241 443 242
rect 441 241 442 242
rect 440 241 441 242
rect 439 241 440 242
rect 438 241 439 242
rect 437 241 438 242
rect 436 241 437 242
rect 426 241 427 242
rect 425 241 426 242
rect 424 241 425 242
rect 423 241 424 242
rect 422 241 423 242
rect 421 241 422 242
rect 420 241 421 242
rect 399 241 400 242
rect 398 241 399 242
rect 397 241 398 242
rect 396 241 397 242
rect 310 241 311 242
rect 309 241 310 242
rect 308 241 309 242
rect 307 241 308 242
rect 306 241 307 242
rect 305 241 306 242
rect 304 241 305 242
rect 303 241 304 242
rect 302 241 303 242
rect 301 241 302 242
rect 300 241 301 242
rect 299 241 300 242
rect 298 241 299 242
rect 297 241 298 242
rect 296 241 297 242
rect 295 241 296 242
rect 294 241 295 242
rect 271 241 272 242
rect 270 241 271 242
rect 269 241 270 242
rect 268 241 269 242
rect 267 241 268 242
rect 266 241 267 242
rect 265 241 266 242
rect 264 241 265 242
rect 263 241 264 242
rect 262 241 263 242
rect 261 241 262 242
rect 260 241 261 242
rect 259 241 260 242
rect 258 241 259 242
rect 257 241 258 242
rect 256 241 257 242
rect 255 241 256 242
rect 254 241 255 242
rect 253 241 254 242
rect 252 241 253 242
rect 251 241 252 242
rect 250 241 251 242
rect 249 241 250 242
rect 248 241 249 242
rect 247 241 248 242
rect 246 241 247 242
rect 245 241 246 242
rect 244 241 245 242
rect 243 241 244 242
rect 242 241 243 242
rect 241 241 242 242
rect 240 241 241 242
rect 239 241 240 242
rect 238 241 239 242
rect 237 241 238 242
rect 236 241 237 242
rect 235 241 236 242
rect 234 241 235 242
rect 233 241 234 242
rect 232 241 233 242
rect 231 241 232 242
rect 230 241 231 242
rect 229 241 230 242
rect 228 241 229 242
rect 227 241 228 242
rect 226 241 227 242
rect 225 241 226 242
rect 224 241 225 242
rect 223 241 224 242
rect 222 241 223 242
rect 221 241 222 242
rect 220 241 221 242
rect 219 241 220 242
rect 218 241 219 242
rect 217 241 218 242
rect 216 241 217 242
rect 215 241 216 242
rect 214 241 215 242
rect 213 241 214 242
rect 212 241 213 242
rect 211 241 212 242
rect 210 241 211 242
rect 209 241 210 242
rect 208 241 209 242
rect 207 241 208 242
rect 206 241 207 242
rect 205 241 206 242
rect 204 241 205 242
rect 203 241 204 242
rect 202 241 203 242
rect 201 241 202 242
rect 200 241 201 242
rect 199 241 200 242
rect 198 241 199 242
rect 197 241 198 242
rect 196 241 197 242
rect 195 241 196 242
rect 194 241 195 242
rect 193 241 194 242
rect 192 241 193 242
rect 191 241 192 242
rect 190 241 191 242
rect 189 241 190 242
rect 188 241 189 242
rect 187 241 188 242
rect 186 241 187 242
rect 185 241 186 242
rect 184 241 185 242
rect 183 241 184 242
rect 182 241 183 242
rect 181 241 182 242
rect 180 241 181 242
rect 179 241 180 242
rect 178 241 179 242
rect 150 241 151 242
rect 149 241 150 242
rect 148 241 149 242
rect 147 241 148 242
rect 146 241 147 242
rect 145 241 146 242
rect 144 241 145 242
rect 143 241 144 242
rect 142 241 143 242
rect 141 241 142 242
rect 140 241 141 242
rect 139 241 140 242
rect 138 241 139 242
rect 137 241 138 242
rect 136 241 137 242
rect 135 241 136 242
rect 134 241 135 242
rect 133 241 134 242
rect 132 241 133 242
rect 131 241 132 242
rect 130 241 131 242
rect 129 241 130 242
rect 128 241 129 242
rect 127 241 128 242
rect 126 241 127 242
rect 125 241 126 242
rect 124 241 125 242
rect 123 241 124 242
rect 122 241 123 242
rect 121 241 122 242
rect 120 241 121 242
rect 103 241 104 242
rect 102 241 103 242
rect 101 241 102 242
rect 100 241 101 242
rect 99 241 100 242
rect 98 241 99 242
rect 97 241 98 242
rect 96 241 97 242
rect 95 241 96 242
rect 94 241 95 242
rect 93 241 94 242
rect 92 241 93 242
rect 91 241 92 242
rect 90 241 91 242
rect 89 241 90 242
rect 88 241 89 242
rect 87 241 88 242
rect 86 241 87 242
rect 85 241 86 242
rect 84 241 85 242
rect 83 241 84 242
rect 82 241 83 242
rect 81 241 82 242
rect 80 241 81 242
rect 79 241 80 242
rect 78 241 79 242
rect 77 241 78 242
rect 76 241 77 242
rect 75 241 76 242
rect 74 241 75 242
rect 73 241 74 242
rect 72 241 73 242
rect 71 241 72 242
rect 70 241 71 242
rect 69 241 70 242
rect 68 241 69 242
rect 67 241 68 242
rect 66 241 67 242
rect 65 241 66 242
rect 64 241 65 242
rect 63 241 64 242
rect 62 241 63 242
rect 61 241 62 242
rect 60 241 61 242
rect 59 241 60 242
rect 58 241 59 242
rect 57 241 58 242
rect 56 241 57 242
rect 55 241 56 242
rect 54 241 55 242
rect 53 241 54 242
rect 52 241 53 242
rect 51 241 52 242
rect 50 241 51 242
rect 49 241 50 242
rect 48 241 49 242
rect 47 241 48 242
rect 46 241 47 242
rect 45 241 46 242
rect 44 241 45 242
rect 43 241 44 242
rect 42 241 43 242
rect 41 241 42 242
rect 40 241 41 242
rect 39 241 40 242
rect 38 241 39 242
rect 37 241 38 242
rect 36 241 37 242
rect 35 241 36 242
rect 34 241 35 242
rect 33 241 34 242
rect 32 241 33 242
rect 31 241 32 242
rect 30 241 31 242
rect 23 241 24 242
rect 22 241 23 242
rect 21 241 22 242
rect 20 241 21 242
rect 19 241 20 242
rect 18 241 19 242
rect 17 241 18 242
rect 16 241 17 242
rect 15 241 16 242
rect 14 241 15 242
rect 13 241 14 242
rect 12 241 13 242
rect 11 241 12 242
rect 10 241 11 242
rect 9 241 10 242
rect 8 241 9 242
rect 7 241 8 242
rect 6 241 7 242
rect 442 242 443 243
rect 441 242 442 243
rect 440 242 441 243
rect 439 242 440 243
rect 438 242 439 243
rect 437 242 438 243
rect 436 242 437 243
rect 435 242 436 243
rect 434 242 435 243
rect 433 242 434 243
rect 432 242 433 243
rect 431 242 432 243
rect 430 242 431 243
rect 429 242 430 243
rect 428 242 429 243
rect 427 242 428 243
rect 426 242 427 243
rect 425 242 426 243
rect 424 242 425 243
rect 423 242 424 243
rect 422 242 423 243
rect 421 242 422 243
rect 420 242 421 243
rect 400 242 401 243
rect 399 242 400 243
rect 398 242 399 243
rect 397 242 398 243
rect 396 242 397 243
rect 318 242 319 243
rect 317 242 318 243
rect 316 242 317 243
rect 315 242 316 243
rect 314 242 315 243
rect 313 242 314 243
rect 312 242 313 243
rect 311 242 312 243
rect 310 242 311 243
rect 309 242 310 243
rect 308 242 309 243
rect 307 242 308 243
rect 306 242 307 243
rect 305 242 306 243
rect 304 242 305 243
rect 303 242 304 243
rect 302 242 303 243
rect 301 242 302 243
rect 300 242 301 243
rect 299 242 300 243
rect 298 242 299 243
rect 297 242 298 243
rect 296 242 297 243
rect 295 242 296 243
rect 294 242 295 243
rect 293 242 294 243
rect 292 242 293 243
rect 291 242 292 243
rect 290 242 291 243
rect 289 242 290 243
rect 288 242 289 243
rect 287 242 288 243
rect 270 242 271 243
rect 269 242 270 243
rect 268 242 269 243
rect 267 242 268 243
rect 266 242 267 243
rect 265 242 266 243
rect 264 242 265 243
rect 263 242 264 243
rect 262 242 263 243
rect 261 242 262 243
rect 260 242 261 243
rect 259 242 260 243
rect 258 242 259 243
rect 257 242 258 243
rect 256 242 257 243
rect 255 242 256 243
rect 254 242 255 243
rect 253 242 254 243
rect 252 242 253 243
rect 251 242 252 243
rect 250 242 251 243
rect 249 242 250 243
rect 248 242 249 243
rect 247 242 248 243
rect 246 242 247 243
rect 245 242 246 243
rect 244 242 245 243
rect 243 242 244 243
rect 242 242 243 243
rect 241 242 242 243
rect 240 242 241 243
rect 239 242 240 243
rect 238 242 239 243
rect 237 242 238 243
rect 236 242 237 243
rect 235 242 236 243
rect 234 242 235 243
rect 233 242 234 243
rect 232 242 233 243
rect 231 242 232 243
rect 230 242 231 243
rect 229 242 230 243
rect 228 242 229 243
rect 227 242 228 243
rect 226 242 227 243
rect 225 242 226 243
rect 224 242 225 243
rect 223 242 224 243
rect 222 242 223 243
rect 221 242 222 243
rect 220 242 221 243
rect 219 242 220 243
rect 218 242 219 243
rect 217 242 218 243
rect 216 242 217 243
rect 215 242 216 243
rect 214 242 215 243
rect 213 242 214 243
rect 212 242 213 243
rect 211 242 212 243
rect 210 242 211 243
rect 209 242 210 243
rect 208 242 209 243
rect 207 242 208 243
rect 206 242 207 243
rect 205 242 206 243
rect 204 242 205 243
rect 203 242 204 243
rect 202 242 203 243
rect 201 242 202 243
rect 200 242 201 243
rect 199 242 200 243
rect 198 242 199 243
rect 197 242 198 243
rect 196 242 197 243
rect 195 242 196 243
rect 194 242 195 243
rect 193 242 194 243
rect 192 242 193 243
rect 191 242 192 243
rect 190 242 191 243
rect 189 242 190 243
rect 188 242 189 243
rect 187 242 188 243
rect 186 242 187 243
rect 185 242 186 243
rect 184 242 185 243
rect 183 242 184 243
rect 182 242 183 243
rect 181 242 182 243
rect 151 242 152 243
rect 150 242 151 243
rect 149 242 150 243
rect 148 242 149 243
rect 147 242 148 243
rect 146 242 147 243
rect 145 242 146 243
rect 144 242 145 243
rect 143 242 144 243
rect 142 242 143 243
rect 141 242 142 243
rect 140 242 141 243
rect 139 242 140 243
rect 138 242 139 243
rect 137 242 138 243
rect 136 242 137 243
rect 135 242 136 243
rect 134 242 135 243
rect 133 242 134 243
rect 132 242 133 243
rect 131 242 132 243
rect 130 242 131 243
rect 129 242 130 243
rect 128 242 129 243
rect 127 242 128 243
rect 126 242 127 243
rect 125 242 126 243
rect 124 242 125 243
rect 123 242 124 243
rect 122 242 123 243
rect 121 242 122 243
rect 120 242 121 243
rect 104 242 105 243
rect 103 242 104 243
rect 102 242 103 243
rect 101 242 102 243
rect 100 242 101 243
rect 99 242 100 243
rect 98 242 99 243
rect 97 242 98 243
rect 96 242 97 243
rect 95 242 96 243
rect 94 242 95 243
rect 93 242 94 243
rect 92 242 93 243
rect 91 242 92 243
rect 90 242 91 243
rect 89 242 90 243
rect 88 242 89 243
rect 87 242 88 243
rect 86 242 87 243
rect 85 242 86 243
rect 84 242 85 243
rect 83 242 84 243
rect 82 242 83 243
rect 81 242 82 243
rect 80 242 81 243
rect 79 242 80 243
rect 78 242 79 243
rect 77 242 78 243
rect 76 242 77 243
rect 75 242 76 243
rect 74 242 75 243
rect 73 242 74 243
rect 72 242 73 243
rect 71 242 72 243
rect 70 242 71 243
rect 69 242 70 243
rect 68 242 69 243
rect 67 242 68 243
rect 66 242 67 243
rect 65 242 66 243
rect 64 242 65 243
rect 63 242 64 243
rect 62 242 63 243
rect 61 242 62 243
rect 60 242 61 243
rect 59 242 60 243
rect 58 242 59 243
rect 57 242 58 243
rect 56 242 57 243
rect 55 242 56 243
rect 54 242 55 243
rect 53 242 54 243
rect 52 242 53 243
rect 51 242 52 243
rect 50 242 51 243
rect 49 242 50 243
rect 48 242 49 243
rect 47 242 48 243
rect 46 242 47 243
rect 45 242 46 243
rect 44 242 45 243
rect 43 242 44 243
rect 42 242 43 243
rect 41 242 42 243
rect 40 242 41 243
rect 39 242 40 243
rect 38 242 39 243
rect 37 242 38 243
rect 36 242 37 243
rect 35 242 36 243
rect 34 242 35 243
rect 33 242 34 243
rect 32 242 33 243
rect 31 242 32 243
rect 30 242 31 243
rect 23 242 24 243
rect 22 242 23 243
rect 21 242 22 243
rect 20 242 21 243
rect 19 242 20 243
rect 18 242 19 243
rect 17 242 18 243
rect 16 242 17 243
rect 15 242 16 243
rect 14 242 15 243
rect 13 242 14 243
rect 12 242 13 243
rect 11 242 12 243
rect 10 242 11 243
rect 9 242 10 243
rect 8 242 9 243
rect 7 242 8 243
rect 6 242 7 243
rect 5 242 6 243
rect 441 243 442 244
rect 440 243 441 244
rect 439 243 440 244
rect 438 243 439 244
rect 437 243 438 244
rect 436 243 437 244
rect 435 243 436 244
rect 434 243 435 244
rect 433 243 434 244
rect 432 243 433 244
rect 431 243 432 244
rect 430 243 431 244
rect 429 243 430 244
rect 428 243 429 244
rect 427 243 428 244
rect 426 243 427 244
rect 425 243 426 244
rect 424 243 425 244
rect 423 243 424 244
rect 422 243 423 244
rect 421 243 422 244
rect 420 243 421 244
rect 401 243 402 244
rect 400 243 401 244
rect 399 243 400 244
rect 398 243 399 244
rect 397 243 398 244
rect 322 243 323 244
rect 321 243 322 244
rect 320 243 321 244
rect 319 243 320 244
rect 318 243 319 244
rect 317 243 318 244
rect 316 243 317 244
rect 315 243 316 244
rect 314 243 315 244
rect 313 243 314 244
rect 312 243 313 244
rect 311 243 312 244
rect 310 243 311 244
rect 309 243 310 244
rect 308 243 309 244
rect 307 243 308 244
rect 306 243 307 244
rect 305 243 306 244
rect 304 243 305 244
rect 303 243 304 244
rect 302 243 303 244
rect 301 243 302 244
rect 300 243 301 244
rect 299 243 300 244
rect 298 243 299 244
rect 297 243 298 244
rect 296 243 297 244
rect 295 243 296 244
rect 294 243 295 244
rect 293 243 294 244
rect 292 243 293 244
rect 291 243 292 244
rect 290 243 291 244
rect 289 243 290 244
rect 288 243 289 244
rect 287 243 288 244
rect 286 243 287 244
rect 285 243 286 244
rect 284 243 285 244
rect 283 243 284 244
rect 282 243 283 244
rect 269 243 270 244
rect 268 243 269 244
rect 267 243 268 244
rect 266 243 267 244
rect 265 243 266 244
rect 264 243 265 244
rect 263 243 264 244
rect 262 243 263 244
rect 261 243 262 244
rect 260 243 261 244
rect 259 243 260 244
rect 258 243 259 244
rect 257 243 258 244
rect 256 243 257 244
rect 255 243 256 244
rect 254 243 255 244
rect 253 243 254 244
rect 252 243 253 244
rect 251 243 252 244
rect 250 243 251 244
rect 249 243 250 244
rect 248 243 249 244
rect 247 243 248 244
rect 246 243 247 244
rect 245 243 246 244
rect 244 243 245 244
rect 243 243 244 244
rect 242 243 243 244
rect 241 243 242 244
rect 240 243 241 244
rect 239 243 240 244
rect 238 243 239 244
rect 237 243 238 244
rect 236 243 237 244
rect 235 243 236 244
rect 234 243 235 244
rect 233 243 234 244
rect 232 243 233 244
rect 231 243 232 244
rect 230 243 231 244
rect 229 243 230 244
rect 228 243 229 244
rect 227 243 228 244
rect 226 243 227 244
rect 225 243 226 244
rect 224 243 225 244
rect 223 243 224 244
rect 222 243 223 244
rect 221 243 222 244
rect 220 243 221 244
rect 219 243 220 244
rect 218 243 219 244
rect 217 243 218 244
rect 216 243 217 244
rect 215 243 216 244
rect 214 243 215 244
rect 213 243 214 244
rect 212 243 213 244
rect 211 243 212 244
rect 210 243 211 244
rect 209 243 210 244
rect 208 243 209 244
rect 207 243 208 244
rect 206 243 207 244
rect 205 243 206 244
rect 204 243 205 244
rect 203 243 204 244
rect 202 243 203 244
rect 201 243 202 244
rect 200 243 201 244
rect 199 243 200 244
rect 198 243 199 244
rect 197 243 198 244
rect 196 243 197 244
rect 195 243 196 244
rect 194 243 195 244
rect 193 243 194 244
rect 192 243 193 244
rect 191 243 192 244
rect 190 243 191 244
rect 189 243 190 244
rect 188 243 189 244
rect 187 243 188 244
rect 186 243 187 244
rect 185 243 186 244
rect 184 243 185 244
rect 183 243 184 244
rect 152 243 153 244
rect 151 243 152 244
rect 150 243 151 244
rect 149 243 150 244
rect 148 243 149 244
rect 147 243 148 244
rect 146 243 147 244
rect 145 243 146 244
rect 144 243 145 244
rect 143 243 144 244
rect 142 243 143 244
rect 141 243 142 244
rect 140 243 141 244
rect 139 243 140 244
rect 138 243 139 244
rect 137 243 138 244
rect 136 243 137 244
rect 135 243 136 244
rect 134 243 135 244
rect 133 243 134 244
rect 132 243 133 244
rect 131 243 132 244
rect 130 243 131 244
rect 129 243 130 244
rect 128 243 129 244
rect 127 243 128 244
rect 126 243 127 244
rect 125 243 126 244
rect 124 243 125 244
rect 123 243 124 244
rect 122 243 123 244
rect 121 243 122 244
rect 105 243 106 244
rect 104 243 105 244
rect 103 243 104 244
rect 102 243 103 244
rect 101 243 102 244
rect 100 243 101 244
rect 99 243 100 244
rect 98 243 99 244
rect 97 243 98 244
rect 96 243 97 244
rect 95 243 96 244
rect 94 243 95 244
rect 93 243 94 244
rect 92 243 93 244
rect 91 243 92 244
rect 90 243 91 244
rect 89 243 90 244
rect 88 243 89 244
rect 87 243 88 244
rect 86 243 87 244
rect 85 243 86 244
rect 84 243 85 244
rect 83 243 84 244
rect 82 243 83 244
rect 81 243 82 244
rect 80 243 81 244
rect 79 243 80 244
rect 78 243 79 244
rect 77 243 78 244
rect 76 243 77 244
rect 75 243 76 244
rect 74 243 75 244
rect 73 243 74 244
rect 72 243 73 244
rect 71 243 72 244
rect 70 243 71 244
rect 69 243 70 244
rect 68 243 69 244
rect 67 243 68 244
rect 66 243 67 244
rect 65 243 66 244
rect 64 243 65 244
rect 63 243 64 244
rect 62 243 63 244
rect 61 243 62 244
rect 60 243 61 244
rect 59 243 60 244
rect 58 243 59 244
rect 57 243 58 244
rect 56 243 57 244
rect 55 243 56 244
rect 54 243 55 244
rect 53 243 54 244
rect 52 243 53 244
rect 51 243 52 244
rect 50 243 51 244
rect 49 243 50 244
rect 48 243 49 244
rect 47 243 48 244
rect 46 243 47 244
rect 45 243 46 244
rect 44 243 45 244
rect 43 243 44 244
rect 42 243 43 244
rect 41 243 42 244
rect 40 243 41 244
rect 39 243 40 244
rect 38 243 39 244
rect 37 243 38 244
rect 36 243 37 244
rect 35 243 36 244
rect 34 243 35 244
rect 33 243 34 244
rect 32 243 33 244
rect 31 243 32 244
rect 30 243 31 244
rect 23 243 24 244
rect 22 243 23 244
rect 21 243 22 244
rect 20 243 21 244
rect 19 243 20 244
rect 18 243 19 244
rect 17 243 18 244
rect 16 243 17 244
rect 15 243 16 244
rect 14 243 15 244
rect 13 243 14 244
rect 12 243 13 244
rect 11 243 12 244
rect 10 243 11 244
rect 9 243 10 244
rect 8 243 9 244
rect 7 243 8 244
rect 6 243 7 244
rect 5 243 6 244
rect 441 244 442 245
rect 440 244 441 245
rect 439 244 440 245
rect 438 244 439 245
rect 437 244 438 245
rect 436 244 437 245
rect 435 244 436 245
rect 434 244 435 245
rect 433 244 434 245
rect 432 244 433 245
rect 431 244 432 245
rect 430 244 431 245
rect 429 244 430 245
rect 428 244 429 245
rect 427 244 428 245
rect 426 244 427 245
rect 425 244 426 245
rect 424 244 425 245
rect 423 244 424 245
rect 422 244 423 245
rect 421 244 422 245
rect 420 244 421 245
rect 402 244 403 245
rect 401 244 402 245
rect 400 244 401 245
rect 399 244 400 245
rect 398 244 399 245
rect 397 244 398 245
rect 326 244 327 245
rect 325 244 326 245
rect 324 244 325 245
rect 323 244 324 245
rect 322 244 323 245
rect 321 244 322 245
rect 320 244 321 245
rect 319 244 320 245
rect 318 244 319 245
rect 317 244 318 245
rect 316 244 317 245
rect 315 244 316 245
rect 314 244 315 245
rect 313 244 314 245
rect 312 244 313 245
rect 311 244 312 245
rect 310 244 311 245
rect 309 244 310 245
rect 308 244 309 245
rect 307 244 308 245
rect 306 244 307 245
rect 305 244 306 245
rect 304 244 305 245
rect 303 244 304 245
rect 302 244 303 245
rect 301 244 302 245
rect 300 244 301 245
rect 299 244 300 245
rect 298 244 299 245
rect 297 244 298 245
rect 296 244 297 245
rect 295 244 296 245
rect 294 244 295 245
rect 293 244 294 245
rect 292 244 293 245
rect 291 244 292 245
rect 290 244 291 245
rect 289 244 290 245
rect 288 244 289 245
rect 287 244 288 245
rect 286 244 287 245
rect 285 244 286 245
rect 284 244 285 245
rect 283 244 284 245
rect 282 244 283 245
rect 281 244 282 245
rect 280 244 281 245
rect 279 244 280 245
rect 278 244 279 245
rect 269 244 270 245
rect 268 244 269 245
rect 267 244 268 245
rect 266 244 267 245
rect 265 244 266 245
rect 264 244 265 245
rect 263 244 264 245
rect 262 244 263 245
rect 261 244 262 245
rect 260 244 261 245
rect 259 244 260 245
rect 258 244 259 245
rect 257 244 258 245
rect 256 244 257 245
rect 255 244 256 245
rect 254 244 255 245
rect 253 244 254 245
rect 252 244 253 245
rect 251 244 252 245
rect 250 244 251 245
rect 249 244 250 245
rect 248 244 249 245
rect 247 244 248 245
rect 246 244 247 245
rect 245 244 246 245
rect 244 244 245 245
rect 243 244 244 245
rect 242 244 243 245
rect 241 244 242 245
rect 240 244 241 245
rect 239 244 240 245
rect 238 244 239 245
rect 237 244 238 245
rect 236 244 237 245
rect 235 244 236 245
rect 234 244 235 245
rect 230 244 231 245
rect 229 244 230 245
rect 228 244 229 245
rect 227 244 228 245
rect 226 244 227 245
rect 225 244 226 245
rect 224 244 225 245
rect 223 244 224 245
rect 222 244 223 245
rect 221 244 222 245
rect 220 244 221 245
rect 219 244 220 245
rect 218 244 219 245
rect 217 244 218 245
rect 216 244 217 245
rect 215 244 216 245
rect 214 244 215 245
rect 213 244 214 245
rect 212 244 213 245
rect 211 244 212 245
rect 210 244 211 245
rect 209 244 210 245
rect 208 244 209 245
rect 207 244 208 245
rect 206 244 207 245
rect 205 244 206 245
rect 204 244 205 245
rect 203 244 204 245
rect 202 244 203 245
rect 201 244 202 245
rect 200 244 201 245
rect 199 244 200 245
rect 198 244 199 245
rect 197 244 198 245
rect 196 244 197 245
rect 195 244 196 245
rect 194 244 195 245
rect 193 244 194 245
rect 192 244 193 245
rect 191 244 192 245
rect 190 244 191 245
rect 189 244 190 245
rect 188 244 189 245
rect 187 244 188 245
rect 186 244 187 245
rect 152 244 153 245
rect 151 244 152 245
rect 150 244 151 245
rect 149 244 150 245
rect 148 244 149 245
rect 147 244 148 245
rect 146 244 147 245
rect 145 244 146 245
rect 144 244 145 245
rect 143 244 144 245
rect 142 244 143 245
rect 141 244 142 245
rect 140 244 141 245
rect 139 244 140 245
rect 138 244 139 245
rect 137 244 138 245
rect 136 244 137 245
rect 135 244 136 245
rect 134 244 135 245
rect 133 244 134 245
rect 132 244 133 245
rect 131 244 132 245
rect 130 244 131 245
rect 129 244 130 245
rect 128 244 129 245
rect 127 244 128 245
rect 126 244 127 245
rect 125 244 126 245
rect 124 244 125 245
rect 123 244 124 245
rect 122 244 123 245
rect 121 244 122 245
rect 106 244 107 245
rect 105 244 106 245
rect 104 244 105 245
rect 103 244 104 245
rect 102 244 103 245
rect 101 244 102 245
rect 100 244 101 245
rect 99 244 100 245
rect 98 244 99 245
rect 97 244 98 245
rect 96 244 97 245
rect 95 244 96 245
rect 94 244 95 245
rect 93 244 94 245
rect 92 244 93 245
rect 91 244 92 245
rect 90 244 91 245
rect 89 244 90 245
rect 88 244 89 245
rect 87 244 88 245
rect 86 244 87 245
rect 85 244 86 245
rect 84 244 85 245
rect 83 244 84 245
rect 82 244 83 245
rect 81 244 82 245
rect 80 244 81 245
rect 79 244 80 245
rect 78 244 79 245
rect 77 244 78 245
rect 76 244 77 245
rect 75 244 76 245
rect 74 244 75 245
rect 73 244 74 245
rect 72 244 73 245
rect 71 244 72 245
rect 70 244 71 245
rect 69 244 70 245
rect 68 244 69 245
rect 67 244 68 245
rect 66 244 67 245
rect 65 244 66 245
rect 64 244 65 245
rect 63 244 64 245
rect 62 244 63 245
rect 61 244 62 245
rect 60 244 61 245
rect 59 244 60 245
rect 58 244 59 245
rect 57 244 58 245
rect 56 244 57 245
rect 55 244 56 245
rect 54 244 55 245
rect 53 244 54 245
rect 52 244 53 245
rect 51 244 52 245
rect 50 244 51 245
rect 49 244 50 245
rect 48 244 49 245
rect 47 244 48 245
rect 46 244 47 245
rect 45 244 46 245
rect 44 244 45 245
rect 43 244 44 245
rect 42 244 43 245
rect 41 244 42 245
rect 40 244 41 245
rect 39 244 40 245
rect 38 244 39 245
rect 37 244 38 245
rect 36 244 37 245
rect 35 244 36 245
rect 34 244 35 245
rect 33 244 34 245
rect 32 244 33 245
rect 31 244 32 245
rect 23 244 24 245
rect 22 244 23 245
rect 21 244 22 245
rect 20 244 21 245
rect 19 244 20 245
rect 18 244 19 245
rect 17 244 18 245
rect 16 244 17 245
rect 15 244 16 245
rect 14 244 15 245
rect 13 244 14 245
rect 12 244 13 245
rect 11 244 12 245
rect 10 244 11 245
rect 9 244 10 245
rect 8 244 9 245
rect 7 244 8 245
rect 6 244 7 245
rect 5 244 6 245
rect 441 245 442 246
rect 440 245 441 246
rect 439 245 440 246
rect 438 245 439 246
rect 437 245 438 246
rect 436 245 437 246
rect 435 245 436 246
rect 434 245 435 246
rect 433 245 434 246
rect 432 245 433 246
rect 431 245 432 246
rect 430 245 431 246
rect 429 245 430 246
rect 428 245 429 246
rect 427 245 428 246
rect 426 245 427 246
rect 425 245 426 246
rect 424 245 425 246
rect 423 245 424 246
rect 422 245 423 246
rect 421 245 422 246
rect 420 245 421 246
rect 403 245 404 246
rect 402 245 403 246
rect 401 245 402 246
rect 400 245 401 246
rect 399 245 400 246
rect 398 245 399 246
rect 397 245 398 246
rect 329 245 330 246
rect 328 245 329 246
rect 327 245 328 246
rect 326 245 327 246
rect 325 245 326 246
rect 324 245 325 246
rect 323 245 324 246
rect 322 245 323 246
rect 321 245 322 246
rect 320 245 321 246
rect 319 245 320 246
rect 318 245 319 246
rect 317 245 318 246
rect 316 245 317 246
rect 315 245 316 246
rect 314 245 315 246
rect 313 245 314 246
rect 312 245 313 246
rect 311 245 312 246
rect 310 245 311 246
rect 309 245 310 246
rect 308 245 309 246
rect 307 245 308 246
rect 306 245 307 246
rect 305 245 306 246
rect 304 245 305 246
rect 303 245 304 246
rect 302 245 303 246
rect 301 245 302 246
rect 300 245 301 246
rect 299 245 300 246
rect 298 245 299 246
rect 297 245 298 246
rect 296 245 297 246
rect 295 245 296 246
rect 294 245 295 246
rect 293 245 294 246
rect 292 245 293 246
rect 291 245 292 246
rect 290 245 291 246
rect 289 245 290 246
rect 288 245 289 246
rect 287 245 288 246
rect 286 245 287 246
rect 285 245 286 246
rect 284 245 285 246
rect 283 245 284 246
rect 282 245 283 246
rect 281 245 282 246
rect 280 245 281 246
rect 279 245 280 246
rect 278 245 279 246
rect 277 245 278 246
rect 276 245 277 246
rect 275 245 276 246
rect 268 245 269 246
rect 267 245 268 246
rect 266 245 267 246
rect 265 245 266 246
rect 264 245 265 246
rect 263 245 264 246
rect 262 245 263 246
rect 261 245 262 246
rect 260 245 261 246
rect 259 245 260 246
rect 258 245 259 246
rect 257 245 258 246
rect 256 245 257 246
rect 255 245 256 246
rect 254 245 255 246
rect 253 245 254 246
rect 252 245 253 246
rect 251 245 252 246
rect 250 245 251 246
rect 249 245 250 246
rect 248 245 249 246
rect 247 245 248 246
rect 246 245 247 246
rect 245 245 246 246
rect 244 245 245 246
rect 243 245 244 246
rect 242 245 243 246
rect 241 245 242 246
rect 240 245 241 246
rect 239 245 240 246
rect 238 245 239 246
rect 237 245 238 246
rect 236 245 237 246
rect 235 245 236 246
rect 234 245 235 246
rect 226 245 227 246
rect 225 245 226 246
rect 224 245 225 246
rect 223 245 224 246
rect 222 245 223 246
rect 221 245 222 246
rect 220 245 221 246
rect 219 245 220 246
rect 218 245 219 246
rect 217 245 218 246
rect 216 245 217 246
rect 215 245 216 246
rect 214 245 215 246
rect 213 245 214 246
rect 212 245 213 246
rect 211 245 212 246
rect 210 245 211 246
rect 209 245 210 246
rect 208 245 209 246
rect 207 245 208 246
rect 206 245 207 246
rect 205 245 206 246
rect 204 245 205 246
rect 203 245 204 246
rect 202 245 203 246
rect 201 245 202 246
rect 200 245 201 246
rect 199 245 200 246
rect 198 245 199 246
rect 197 245 198 246
rect 196 245 197 246
rect 195 245 196 246
rect 194 245 195 246
rect 193 245 194 246
rect 192 245 193 246
rect 191 245 192 246
rect 190 245 191 246
rect 189 245 190 246
rect 153 245 154 246
rect 152 245 153 246
rect 151 245 152 246
rect 150 245 151 246
rect 149 245 150 246
rect 148 245 149 246
rect 147 245 148 246
rect 146 245 147 246
rect 145 245 146 246
rect 144 245 145 246
rect 143 245 144 246
rect 142 245 143 246
rect 141 245 142 246
rect 140 245 141 246
rect 139 245 140 246
rect 138 245 139 246
rect 137 245 138 246
rect 136 245 137 246
rect 135 245 136 246
rect 134 245 135 246
rect 133 245 134 246
rect 132 245 133 246
rect 131 245 132 246
rect 130 245 131 246
rect 129 245 130 246
rect 128 245 129 246
rect 127 245 128 246
rect 126 245 127 246
rect 125 245 126 246
rect 124 245 125 246
rect 123 245 124 246
rect 122 245 123 246
rect 121 245 122 246
rect 106 245 107 246
rect 105 245 106 246
rect 104 245 105 246
rect 103 245 104 246
rect 102 245 103 246
rect 101 245 102 246
rect 100 245 101 246
rect 99 245 100 246
rect 98 245 99 246
rect 97 245 98 246
rect 96 245 97 246
rect 95 245 96 246
rect 94 245 95 246
rect 93 245 94 246
rect 92 245 93 246
rect 91 245 92 246
rect 90 245 91 246
rect 89 245 90 246
rect 88 245 89 246
rect 87 245 88 246
rect 86 245 87 246
rect 85 245 86 246
rect 84 245 85 246
rect 83 245 84 246
rect 82 245 83 246
rect 81 245 82 246
rect 80 245 81 246
rect 79 245 80 246
rect 78 245 79 246
rect 77 245 78 246
rect 76 245 77 246
rect 75 245 76 246
rect 74 245 75 246
rect 73 245 74 246
rect 72 245 73 246
rect 71 245 72 246
rect 70 245 71 246
rect 69 245 70 246
rect 68 245 69 246
rect 67 245 68 246
rect 66 245 67 246
rect 65 245 66 246
rect 64 245 65 246
rect 63 245 64 246
rect 62 245 63 246
rect 61 245 62 246
rect 60 245 61 246
rect 59 245 60 246
rect 58 245 59 246
rect 57 245 58 246
rect 56 245 57 246
rect 55 245 56 246
rect 54 245 55 246
rect 53 245 54 246
rect 52 245 53 246
rect 51 245 52 246
rect 50 245 51 246
rect 49 245 50 246
rect 48 245 49 246
rect 47 245 48 246
rect 46 245 47 246
rect 45 245 46 246
rect 44 245 45 246
rect 43 245 44 246
rect 42 245 43 246
rect 41 245 42 246
rect 40 245 41 246
rect 39 245 40 246
rect 38 245 39 246
rect 37 245 38 246
rect 36 245 37 246
rect 35 245 36 246
rect 34 245 35 246
rect 33 245 34 246
rect 32 245 33 246
rect 31 245 32 246
rect 23 245 24 246
rect 22 245 23 246
rect 21 245 22 246
rect 20 245 21 246
rect 19 245 20 246
rect 18 245 19 246
rect 17 245 18 246
rect 16 245 17 246
rect 15 245 16 246
rect 14 245 15 246
rect 13 245 14 246
rect 12 245 13 246
rect 11 245 12 246
rect 10 245 11 246
rect 9 245 10 246
rect 8 245 9 246
rect 7 245 8 246
rect 6 245 7 246
rect 5 245 6 246
rect 481 246 482 247
rect 480 246 481 247
rect 479 246 480 247
rect 478 246 479 247
rect 477 246 478 247
rect 468 246 469 247
rect 467 246 468 247
rect 466 246 467 247
rect 441 246 442 247
rect 440 246 441 247
rect 439 246 440 247
rect 438 246 439 247
rect 437 246 438 247
rect 436 246 437 247
rect 435 246 436 247
rect 434 246 435 247
rect 433 246 434 247
rect 432 246 433 247
rect 431 246 432 247
rect 430 246 431 247
rect 429 246 430 247
rect 428 246 429 247
rect 427 246 428 247
rect 426 246 427 247
rect 425 246 426 247
rect 424 246 425 247
rect 423 246 424 247
rect 422 246 423 247
rect 421 246 422 247
rect 420 246 421 247
rect 404 246 405 247
rect 403 246 404 247
rect 402 246 403 247
rect 401 246 402 247
rect 400 246 401 247
rect 399 246 400 247
rect 398 246 399 247
rect 397 246 398 247
rect 329 246 330 247
rect 328 246 329 247
rect 327 246 328 247
rect 326 246 327 247
rect 325 246 326 247
rect 324 246 325 247
rect 323 246 324 247
rect 322 246 323 247
rect 321 246 322 247
rect 320 246 321 247
rect 319 246 320 247
rect 318 246 319 247
rect 317 246 318 247
rect 316 246 317 247
rect 315 246 316 247
rect 314 246 315 247
rect 313 246 314 247
rect 312 246 313 247
rect 311 246 312 247
rect 310 246 311 247
rect 309 246 310 247
rect 308 246 309 247
rect 307 246 308 247
rect 306 246 307 247
rect 305 246 306 247
rect 304 246 305 247
rect 303 246 304 247
rect 302 246 303 247
rect 301 246 302 247
rect 300 246 301 247
rect 299 246 300 247
rect 298 246 299 247
rect 297 246 298 247
rect 296 246 297 247
rect 295 246 296 247
rect 294 246 295 247
rect 293 246 294 247
rect 292 246 293 247
rect 291 246 292 247
rect 290 246 291 247
rect 289 246 290 247
rect 288 246 289 247
rect 287 246 288 247
rect 286 246 287 247
rect 285 246 286 247
rect 284 246 285 247
rect 283 246 284 247
rect 282 246 283 247
rect 281 246 282 247
rect 280 246 281 247
rect 279 246 280 247
rect 278 246 279 247
rect 277 246 278 247
rect 276 246 277 247
rect 275 246 276 247
rect 274 246 275 247
rect 273 246 274 247
rect 267 246 268 247
rect 266 246 267 247
rect 265 246 266 247
rect 264 246 265 247
rect 263 246 264 247
rect 262 246 263 247
rect 261 246 262 247
rect 260 246 261 247
rect 259 246 260 247
rect 258 246 259 247
rect 257 246 258 247
rect 256 246 257 247
rect 255 246 256 247
rect 254 246 255 247
rect 253 246 254 247
rect 252 246 253 247
rect 251 246 252 247
rect 250 246 251 247
rect 249 246 250 247
rect 248 246 249 247
rect 247 246 248 247
rect 246 246 247 247
rect 245 246 246 247
rect 244 246 245 247
rect 243 246 244 247
rect 242 246 243 247
rect 241 246 242 247
rect 240 246 241 247
rect 239 246 240 247
rect 238 246 239 247
rect 237 246 238 247
rect 236 246 237 247
rect 235 246 236 247
rect 234 246 235 247
rect 222 246 223 247
rect 221 246 222 247
rect 220 246 221 247
rect 219 246 220 247
rect 218 246 219 247
rect 217 246 218 247
rect 216 246 217 247
rect 215 246 216 247
rect 214 246 215 247
rect 213 246 214 247
rect 212 246 213 247
rect 211 246 212 247
rect 210 246 211 247
rect 209 246 210 247
rect 208 246 209 247
rect 207 246 208 247
rect 206 246 207 247
rect 205 246 206 247
rect 204 246 205 247
rect 203 246 204 247
rect 202 246 203 247
rect 201 246 202 247
rect 200 246 201 247
rect 199 246 200 247
rect 198 246 199 247
rect 197 246 198 247
rect 196 246 197 247
rect 195 246 196 247
rect 194 246 195 247
rect 193 246 194 247
rect 154 246 155 247
rect 153 246 154 247
rect 152 246 153 247
rect 151 246 152 247
rect 150 246 151 247
rect 149 246 150 247
rect 148 246 149 247
rect 147 246 148 247
rect 146 246 147 247
rect 145 246 146 247
rect 144 246 145 247
rect 143 246 144 247
rect 142 246 143 247
rect 141 246 142 247
rect 140 246 141 247
rect 139 246 140 247
rect 138 246 139 247
rect 137 246 138 247
rect 136 246 137 247
rect 135 246 136 247
rect 134 246 135 247
rect 133 246 134 247
rect 132 246 133 247
rect 131 246 132 247
rect 130 246 131 247
rect 129 246 130 247
rect 128 246 129 247
rect 127 246 128 247
rect 126 246 127 247
rect 125 246 126 247
rect 124 246 125 247
rect 123 246 124 247
rect 122 246 123 247
rect 121 246 122 247
rect 107 246 108 247
rect 106 246 107 247
rect 105 246 106 247
rect 104 246 105 247
rect 103 246 104 247
rect 102 246 103 247
rect 101 246 102 247
rect 100 246 101 247
rect 99 246 100 247
rect 98 246 99 247
rect 97 246 98 247
rect 96 246 97 247
rect 95 246 96 247
rect 94 246 95 247
rect 93 246 94 247
rect 92 246 93 247
rect 91 246 92 247
rect 90 246 91 247
rect 89 246 90 247
rect 88 246 89 247
rect 87 246 88 247
rect 86 246 87 247
rect 85 246 86 247
rect 84 246 85 247
rect 83 246 84 247
rect 82 246 83 247
rect 81 246 82 247
rect 80 246 81 247
rect 79 246 80 247
rect 78 246 79 247
rect 77 246 78 247
rect 76 246 77 247
rect 75 246 76 247
rect 74 246 75 247
rect 73 246 74 247
rect 72 246 73 247
rect 71 246 72 247
rect 70 246 71 247
rect 69 246 70 247
rect 68 246 69 247
rect 67 246 68 247
rect 66 246 67 247
rect 65 246 66 247
rect 64 246 65 247
rect 63 246 64 247
rect 62 246 63 247
rect 61 246 62 247
rect 60 246 61 247
rect 59 246 60 247
rect 58 246 59 247
rect 57 246 58 247
rect 56 246 57 247
rect 55 246 56 247
rect 54 246 55 247
rect 53 246 54 247
rect 52 246 53 247
rect 51 246 52 247
rect 50 246 51 247
rect 49 246 50 247
rect 48 246 49 247
rect 47 246 48 247
rect 46 246 47 247
rect 45 246 46 247
rect 44 246 45 247
rect 43 246 44 247
rect 42 246 43 247
rect 41 246 42 247
rect 40 246 41 247
rect 39 246 40 247
rect 38 246 39 247
rect 37 246 38 247
rect 36 246 37 247
rect 35 246 36 247
rect 34 246 35 247
rect 33 246 34 247
rect 32 246 33 247
rect 31 246 32 247
rect 23 246 24 247
rect 22 246 23 247
rect 21 246 22 247
rect 20 246 21 247
rect 19 246 20 247
rect 18 246 19 247
rect 17 246 18 247
rect 16 246 17 247
rect 15 246 16 247
rect 14 246 15 247
rect 13 246 14 247
rect 12 246 13 247
rect 11 246 12 247
rect 10 246 11 247
rect 9 246 10 247
rect 8 246 9 247
rect 7 246 8 247
rect 6 246 7 247
rect 5 246 6 247
rect 482 247 483 248
rect 481 247 482 248
rect 480 247 481 248
rect 479 247 480 248
rect 478 247 479 248
rect 470 247 471 248
rect 469 247 470 248
rect 468 247 469 248
rect 467 247 468 248
rect 466 247 467 248
rect 465 247 466 248
rect 464 247 465 248
rect 441 247 442 248
rect 440 247 441 248
rect 439 247 440 248
rect 438 247 439 248
rect 437 247 438 248
rect 436 247 437 248
rect 435 247 436 248
rect 434 247 435 248
rect 433 247 434 248
rect 432 247 433 248
rect 431 247 432 248
rect 430 247 431 248
rect 429 247 430 248
rect 428 247 429 248
rect 427 247 428 248
rect 426 247 427 248
rect 425 247 426 248
rect 424 247 425 248
rect 423 247 424 248
rect 422 247 423 248
rect 421 247 422 248
rect 420 247 421 248
rect 406 247 407 248
rect 405 247 406 248
rect 404 247 405 248
rect 403 247 404 248
rect 402 247 403 248
rect 401 247 402 248
rect 400 247 401 248
rect 399 247 400 248
rect 398 247 399 248
rect 397 247 398 248
rect 327 247 328 248
rect 326 247 327 248
rect 325 247 326 248
rect 324 247 325 248
rect 323 247 324 248
rect 322 247 323 248
rect 321 247 322 248
rect 320 247 321 248
rect 319 247 320 248
rect 318 247 319 248
rect 317 247 318 248
rect 316 247 317 248
rect 315 247 316 248
rect 314 247 315 248
rect 313 247 314 248
rect 312 247 313 248
rect 311 247 312 248
rect 310 247 311 248
rect 309 247 310 248
rect 308 247 309 248
rect 307 247 308 248
rect 306 247 307 248
rect 305 247 306 248
rect 304 247 305 248
rect 303 247 304 248
rect 302 247 303 248
rect 301 247 302 248
rect 300 247 301 248
rect 299 247 300 248
rect 298 247 299 248
rect 297 247 298 248
rect 296 247 297 248
rect 295 247 296 248
rect 294 247 295 248
rect 293 247 294 248
rect 292 247 293 248
rect 291 247 292 248
rect 290 247 291 248
rect 289 247 290 248
rect 288 247 289 248
rect 287 247 288 248
rect 286 247 287 248
rect 285 247 286 248
rect 284 247 285 248
rect 283 247 284 248
rect 282 247 283 248
rect 281 247 282 248
rect 280 247 281 248
rect 279 247 280 248
rect 278 247 279 248
rect 277 247 278 248
rect 276 247 277 248
rect 275 247 276 248
rect 274 247 275 248
rect 273 247 274 248
rect 272 247 273 248
rect 271 247 272 248
rect 267 247 268 248
rect 266 247 267 248
rect 265 247 266 248
rect 264 247 265 248
rect 263 247 264 248
rect 262 247 263 248
rect 261 247 262 248
rect 260 247 261 248
rect 259 247 260 248
rect 258 247 259 248
rect 257 247 258 248
rect 256 247 257 248
rect 255 247 256 248
rect 254 247 255 248
rect 253 247 254 248
rect 252 247 253 248
rect 251 247 252 248
rect 250 247 251 248
rect 249 247 250 248
rect 248 247 249 248
rect 247 247 248 248
rect 246 247 247 248
rect 245 247 246 248
rect 244 247 245 248
rect 243 247 244 248
rect 242 247 243 248
rect 241 247 242 248
rect 240 247 241 248
rect 239 247 240 248
rect 238 247 239 248
rect 237 247 238 248
rect 236 247 237 248
rect 235 247 236 248
rect 234 247 235 248
rect 216 247 217 248
rect 215 247 216 248
rect 214 247 215 248
rect 213 247 214 248
rect 212 247 213 248
rect 211 247 212 248
rect 210 247 211 248
rect 209 247 210 248
rect 208 247 209 248
rect 207 247 208 248
rect 206 247 207 248
rect 205 247 206 248
rect 204 247 205 248
rect 203 247 204 248
rect 202 247 203 248
rect 201 247 202 248
rect 200 247 201 248
rect 199 247 200 248
rect 198 247 199 248
rect 155 247 156 248
rect 154 247 155 248
rect 153 247 154 248
rect 152 247 153 248
rect 151 247 152 248
rect 150 247 151 248
rect 149 247 150 248
rect 148 247 149 248
rect 147 247 148 248
rect 146 247 147 248
rect 145 247 146 248
rect 144 247 145 248
rect 143 247 144 248
rect 142 247 143 248
rect 141 247 142 248
rect 140 247 141 248
rect 139 247 140 248
rect 138 247 139 248
rect 137 247 138 248
rect 136 247 137 248
rect 135 247 136 248
rect 134 247 135 248
rect 133 247 134 248
rect 132 247 133 248
rect 131 247 132 248
rect 130 247 131 248
rect 129 247 130 248
rect 128 247 129 248
rect 127 247 128 248
rect 126 247 127 248
rect 125 247 126 248
rect 124 247 125 248
rect 123 247 124 248
rect 122 247 123 248
rect 107 247 108 248
rect 106 247 107 248
rect 105 247 106 248
rect 104 247 105 248
rect 103 247 104 248
rect 102 247 103 248
rect 101 247 102 248
rect 100 247 101 248
rect 99 247 100 248
rect 98 247 99 248
rect 97 247 98 248
rect 96 247 97 248
rect 95 247 96 248
rect 94 247 95 248
rect 93 247 94 248
rect 92 247 93 248
rect 91 247 92 248
rect 90 247 91 248
rect 89 247 90 248
rect 88 247 89 248
rect 87 247 88 248
rect 86 247 87 248
rect 85 247 86 248
rect 84 247 85 248
rect 83 247 84 248
rect 82 247 83 248
rect 81 247 82 248
rect 80 247 81 248
rect 79 247 80 248
rect 78 247 79 248
rect 77 247 78 248
rect 76 247 77 248
rect 75 247 76 248
rect 74 247 75 248
rect 73 247 74 248
rect 72 247 73 248
rect 71 247 72 248
rect 70 247 71 248
rect 69 247 70 248
rect 68 247 69 248
rect 67 247 68 248
rect 66 247 67 248
rect 65 247 66 248
rect 64 247 65 248
rect 63 247 64 248
rect 62 247 63 248
rect 61 247 62 248
rect 60 247 61 248
rect 59 247 60 248
rect 58 247 59 248
rect 57 247 58 248
rect 56 247 57 248
rect 55 247 56 248
rect 54 247 55 248
rect 53 247 54 248
rect 52 247 53 248
rect 51 247 52 248
rect 50 247 51 248
rect 49 247 50 248
rect 48 247 49 248
rect 47 247 48 248
rect 46 247 47 248
rect 45 247 46 248
rect 44 247 45 248
rect 43 247 44 248
rect 42 247 43 248
rect 41 247 42 248
rect 40 247 41 248
rect 39 247 40 248
rect 38 247 39 248
rect 37 247 38 248
rect 36 247 37 248
rect 35 247 36 248
rect 34 247 35 248
rect 33 247 34 248
rect 32 247 33 248
rect 31 247 32 248
rect 23 247 24 248
rect 22 247 23 248
rect 21 247 22 248
rect 20 247 21 248
rect 19 247 20 248
rect 18 247 19 248
rect 17 247 18 248
rect 16 247 17 248
rect 15 247 16 248
rect 14 247 15 248
rect 13 247 14 248
rect 12 247 13 248
rect 11 247 12 248
rect 10 247 11 248
rect 9 247 10 248
rect 8 247 9 248
rect 7 247 8 248
rect 6 247 7 248
rect 5 247 6 248
rect 482 248 483 249
rect 481 248 482 249
rect 480 248 481 249
rect 479 248 480 249
rect 471 248 472 249
rect 470 248 471 249
rect 469 248 470 249
rect 468 248 469 249
rect 467 248 468 249
rect 466 248 467 249
rect 465 248 466 249
rect 464 248 465 249
rect 463 248 464 249
rect 440 248 441 249
rect 439 248 440 249
rect 438 248 439 249
rect 437 248 438 249
rect 436 248 437 249
rect 435 248 436 249
rect 434 248 435 249
rect 433 248 434 249
rect 432 248 433 249
rect 431 248 432 249
rect 430 248 431 249
rect 429 248 430 249
rect 428 248 429 249
rect 427 248 428 249
rect 426 248 427 249
rect 425 248 426 249
rect 424 248 425 249
rect 423 248 424 249
rect 422 248 423 249
rect 421 248 422 249
rect 420 248 421 249
rect 409 248 410 249
rect 408 248 409 249
rect 407 248 408 249
rect 406 248 407 249
rect 405 248 406 249
rect 404 248 405 249
rect 403 248 404 249
rect 402 248 403 249
rect 401 248 402 249
rect 400 248 401 249
rect 399 248 400 249
rect 398 248 399 249
rect 325 248 326 249
rect 324 248 325 249
rect 323 248 324 249
rect 322 248 323 249
rect 321 248 322 249
rect 320 248 321 249
rect 319 248 320 249
rect 318 248 319 249
rect 317 248 318 249
rect 316 248 317 249
rect 315 248 316 249
rect 314 248 315 249
rect 313 248 314 249
rect 312 248 313 249
rect 311 248 312 249
rect 310 248 311 249
rect 309 248 310 249
rect 308 248 309 249
rect 307 248 308 249
rect 306 248 307 249
rect 305 248 306 249
rect 304 248 305 249
rect 303 248 304 249
rect 302 248 303 249
rect 301 248 302 249
rect 300 248 301 249
rect 299 248 300 249
rect 298 248 299 249
rect 297 248 298 249
rect 296 248 297 249
rect 295 248 296 249
rect 294 248 295 249
rect 293 248 294 249
rect 292 248 293 249
rect 291 248 292 249
rect 290 248 291 249
rect 289 248 290 249
rect 288 248 289 249
rect 287 248 288 249
rect 286 248 287 249
rect 285 248 286 249
rect 284 248 285 249
rect 283 248 284 249
rect 282 248 283 249
rect 281 248 282 249
rect 280 248 281 249
rect 279 248 280 249
rect 278 248 279 249
rect 277 248 278 249
rect 276 248 277 249
rect 275 248 276 249
rect 274 248 275 249
rect 273 248 274 249
rect 272 248 273 249
rect 271 248 272 249
rect 270 248 271 249
rect 269 248 270 249
rect 266 248 267 249
rect 265 248 266 249
rect 264 248 265 249
rect 263 248 264 249
rect 262 248 263 249
rect 261 248 262 249
rect 260 248 261 249
rect 259 248 260 249
rect 258 248 259 249
rect 257 248 258 249
rect 256 248 257 249
rect 255 248 256 249
rect 254 248 255 249
rect 253 248 254 249
rect 252 248 253 249
rect 251 248 252 249
rect 250 248 251 249
rect 249 248 250 249
rect 248 248 249 249
rect 247 248 248 249
rect 246 248 247 249
rect 245 248 246 249
rect 244 248 245 249
rect 243 248 244 249
rect 242 248 243 249
rect 241 248 242 249
rect 240 248 241 249
rect 239 248 240 249
rect 238 248 239 249
rect 237 248 238 249
rect 236 248 237 249
rect 235 248 236 249
rect 234 248 235 249
rect 156 248 157 249
rect 155 248 156 249
rect 154 248 155 249
rect 153 248 154 249
rect 152 248 153 249
rect 151 248 152 249
rect 150 248 151 249
rect 149 248 150 249
rect 148 248 149 249
rect 147 248 148 249
rect 146 248 147 249
rect 145 248 146 249
rect 144 248 145 249
rect 143 248 144 249
rect 142 248 143 249
rect 141 248 142 249
rect 140 248 141 249
rect 139 248 140 249
rect 138 248 139 249
rect 137 248 138 249
rect 136 248 137 249
rect 135 248 136 249
rect 134 248 135 249
rect 133 248 134 249
rect 132 248 133 249
rect 131 248 132 249
rect 130 248 131 249
rect 129 248 130 249
rect 128 248 129 249
rect 127 248 128 249
rect 126 248 127 249
rect 125 248 126 249
rect 124 248 125 249
rect 123 248 124 249
rect 122 248 123 249
rect 108 248 109 249
rect 107 248 108 249
rect 106 248 107 249
rect 105 248 106 249
rect 104 248 105 249
rect 103 248 104 249
rect 102 248 103 249
rect 101 248 102 249
rect 100 248 101 249
rect 99 248 100 249
rect 98 248 99 249
rect 97 248 98 249
rect 96 248 97 249
rect 95 248 96 249
rect 94 248 95 249
rect 93 248 94 249
rect 92 248 93 249
rect 91 248 92 249
rect 90 248 91 249
rect 89 248 90 249
rect 88 248 89 249
rect 87 248 88 249
rect 86 248 87 249
rect 85 248 86 249
rect 84 248 85 249
rect 83 248 84 249
rect 82 248 83 249
rect 81 248 82 249
rect 80 248 81 249
rect 79 248 80 249
rect 78 248 79 249
rect 77 248 78 249
rect 76 248 77 249
rect 75 248 76 249
rect 74 248 75 249
rect 73 248 74 249
rect 72 248 73 249
rect 71 248 72 249
rect 70 248 71 249
rect 69 248 70 249
rect 68 248 69 249
rect 67 248 68 249
rect 66 248 67 249
rect 65 248 66 249
rect 64 248 65 249
rect 63 248 64 249
rect 62 248 63 249
rect 61 248 62 249
rect 60 248 61 249
rect 59 248 60 249
rect 58 248 59 249
rect 57 248 58 249
rect 56 248 57 249
rect 55 248 56 249
rect 54 248 55 249
rect 53 248 54 249
rect 52 248 53 249
rect 51 248 52 249
rect 50 248 51 249
rect 49 248 50 249
rect 48 248 49 249
rect 47 248 48 249
rect 46 248 47 249
rect 45 248 46 249
rect 44 248 45 249
rect 43 248 44 249
rect 42 248 43 249
rect 41 248 42 249
rect 40 248 41 249
rect 39 248 40 249
rect 38 248 39 249
rect 37 248 38 249
rect 36 248 37 249
rect 35 248 36 249
rect 34 248 35 249
rect 33 248 34 249
rect 32 248 33 249
rect 23 248 24 249
rect 22 248 23 249
rect 21 248 22 249
rect 20 248 21 249
rect 19 248 20 249
rect 18 248 19 249
rect 17 248 18 249
rect 16 248 17 249
rect 15 248 16 249
rect 14 248 15 249
rect 13 248 14 249
rect 12 248 13 249
rect 11 248 12 249
rect 10 248 11 249
rect 9 248 10 249
rect 8 248 9 249
rect 7 248 8 249
rect 6 248 7 249
rect 5 248 6 249
rect 483 249 484 250
rect 482 249 483 250
rect 481 249 482 250
rect 472 249 473 250
rect 471 249 472 250
rect 470 249 471 250
rect 469 249 470 250
rect 468 249 469 250
rect 467 249 468 250
rect 466 249 467 250
rect 465 249 466 250
rect 464 249 465 250
rect 463 249 464 250
rect 462 249 463 250
rect 440 249 441 250
rect 439 249 440 250
rect 438 249 439 250
rect 437 249 438 250
rect 436 249 437 250
rect 435 249 436 250
rect 434 249 435 250
rect 433 249 434 250
rect 432 249 433 250
rect 431 249 432 250
rect 430 249 431 250
rect 429 249 430 250
rect 428 249 429 250
rect 427 249 428 250
rect 426 249 427 250
rect 425 249 426 250
rect 424 249 425 250
rect 423 249 424 250
rect 422 249 423 250
rect 421 249 422 250
rect 420 249 421 250
rect 409 249 410 250
rect 408 249 409 250
rect 407 249 408 250
rect 406 249 407 250
rect 405 249 406 250
rect 404 249 405 250
rect 403 249 404 250
rect 402 249 403 250
rect 401 249 402 250
rect 400 249 401 250
rect 399 249 400 250
rect 398 249 399 250
rect 323 249 324 250
rect 322 249 323 250
rect 321 249 322 250
rect 320 249 321 250
rect 319 249 320 250
rect 318 249 319 250
rect 317 249 318 250
rect 316 249 317 250
rect 315 249 316 250
rect 314 249 315 250
rect 313 249 314 250
rect 312 249 313 250
rect 311 249 312 250
rect 310 249 311 250
rect 309 249 310 250
rect 308 249 309 250
rect 307 249 308 250
rect 306 249 307 250
rect 305 249 306 250
rect 304 249 305 250
rect 303 249 304 250
rect 302 249 303 250
rect 301 249 302 250
rect 300 249 301 250
rect 299 249 300 250
rect 298 249 299 250
rect 297 249 298 250
rect 296 249 297 250
rect 295 249 296 250
rect 294 249 295 250
rect 293 249 294 250
rect 292 249 293 250
rect 291 249 292 250
rect 290 249 291 250
rect 289 249 290 250
rect 288 249 289 250
rect 287 249 288 250
rect 286 249 287 250
rect 285 249 286 250
rect 284 249 285 250
rect 283 249 284 250
rect 282 249 283 250
rect 281 249 282 250
rect 280 249 281 250
rect 279 249 280 250
rect 278 249 279 250
rect 277 249 278 250
rect 276 249 277 250
rect 275 249 276 250
rect 274 249 275 250
rect 273 249 274 250
rect 272 249 273 250
rect 271 249 272 250
rect 270 249 271 250
rect 269 249 270 250
rect 268 249 269 250
rect 267 249 268 250
rect 265 249 266 250
rect 264 249 265 250
rect 263 249 264 250
rect 262 249 263 250
rect 261 249 262 250
rect 260 249 261 250
rect 259 249 260 250
rect 258 249 259 250
rect 257 249 258 250
rect 256 249 257 250
rect 255 249 256 250
rect 254 249 255 250
rect 253 249 254 250
rect 252 249 253 250
rect 251 249 252 250
rect 250 249 251 250
rect 249 249 250 250
rect 248 249 249 250
rect 247 249 248 250
rect 246 249 247 250
rect 245 249 246 250
rect 244 249 245 250
rect 243 249 244 250
rect 242 249 243 250
rect 241 249 242 250
rect 240 249 241 250
rect 239 249 240 250
rect 238 249 239 250
rect 237 249 238 250
rect 236 249 237 250
rect 235 249 236 250
rect 234 249 235 250
rect 157 249 158 250
rect 156 249 157 250
rect 155 249 156 250
rect 154 249 155 250
rect 153 249 154 250
rect 152 249 153 250
rect 151 249 152 250
rect 150 249 151 250
rect 149 249 150 250
rect 148 249 149 250
rect 147 249 148 250
rect 146 249 147 250
rect 145 249 146 250
rect 144 249 145 250
rect 143 249 144 250
rect 142 249 143 250
rect 141 249 142 250
rect 140 249 141 250
rect 139 249 140 250
rect 138 249 139 250
rect 137 249 138 250
rect 136 249 137 250
rect 135 249 136 250
rect 134 249 135 250
rect 133 249 134 250
rect 132 249 133 250
rect 131 249 132 250
rect 130 249 131 250
rect 129 249 130 250
rect 128 249 129 250
rect 127 249 128 250
rect 126 249 127 250
rect 125 249 126 250
rect 124 249 125 250
rect 123 249 124 250
rect 122 249 123 250
rect 108 249 109 250
rect 107 249 108 250
rect 106 249 107 250
rect 105 249 106 250
rect 104 249 105 250
rect 103 249 104 250
rect 102 249 103 250
rect 101 249 102 250
rect 100 249 101 250
rect 99 249 100 250
rect 98 249 99 250
rect 97 249 98 250
rect 96 249 97 250
rect 95 249 96 250
rect 94 249 95 250
rect 93 249 94 250
rect 92 249 93 250
rect 91 249 92 250
rect 90 249 91 250
rect 89 249 90 250
rect 88 249 89 250
rect 87 249 88 250
rect 86 249 87 250
rect 85 249 86 250
rect 84 249 85 250
rect 83 249 84 250
rect 82 249 83 250
rect 81 249 82 250
rect 80 249 81 250
rect 79 249 80 250
rect 78 249 79 250
rect 77 249 78 250
rect 76 249 77 250
rect 75 249 76 250
rect 74 249 75 250
rect 73 249 74 250
rect 72 249 73 250
rect 71 249 72 250
rect 70 249 71 250
rect 69 249 70 250
rect 68 249 69 250
rect 67 249 68 250
rect 66 249 67 250
rect 65 249 66 250
rect 64 249 65 250
rect 63 249 64 250
rect 62 249 63 250
rect 61 249 62 250
rect 60 249 61 250
rect 59 249 60 250
rect 58 249 59 250
rect 57 249 58 250
rect 56 249 57 250
rect 55 249 56 250
rect 54 249 55 250
rect 53 249 54 250
rect 52 249 53 250
rect 51 249 52 250
rect 50 249 51 250
rect 49 249 50 250
rect 48 249 49 250
rect 47 249 48 250
rect 46 249 47 250
rect 45 249 46 250
rect 44 249 45 250
rect 43 249 44 250
rect 42 249 43 250
rect 41 249 42 250
rect 40 249 41 250
rect 39 249 40 250
rect 38 249 39 250
rect 37 249 38 250
rect 36 249 37 250
rect 35 249 36 250
rect 34 249 35 250
rect 33 249 34 250
rect 32 249 33 250
rect 23 249 24 250
rect 22 249 23 250
rect 21 249 22 250
rect 20 249 21 250
rect 19 249 20 250
rect 18 249 19 250
rect 17 249 18 250
rect 16 249 17 250
rect 15 249 16 250
rect 14 249 15 250
rect 13 249 14 250
rect 12 249 13 250
rect 11 249 12 250
rect 10 249 11 250
rect 9 249 10 250
rect 8 249 9 250
rect 7 249 8 250
rect 6 249 7 250
rect 5 249 6 250
rect 483 250 484 251
rect 482 250 483 251
rect 473 250 474 251
rect 472 250 473 251
rect 471 250 472 251
rect 470 250 471 251
rect 469 250 470 251
rect 468 250 469 251
rect 467 250 468 251
rect 464 250 465 251
rect 463 250 464 251
rect 462 250 463 251
rect 440 250 441 251
rect 439 250 440 251
rect 438 250 439 251
rect 437 250 438 251
rect 436 250 437 251
rect 435 250 436 251
rect 434 250 435 251
rect 433 250 434 251
rect 432 250 433 251
rect 431 250 432 251
rect 430 250 431 251
rect 429 250 430 251
rect 428 250 429 251
rect 427 250 428 251
rect 426 250 427 251
rect 425 250 426 251
rect 424 250 425 251
rect 423 250 424 251
rect 422 250 423 251
rect 421 250 422 251
rect 420 250 421 251
rect 409 250 410 251
rect 408 250 409 251
rect 407 250 408 251
rect 406 250 407 251
rect 405 250 406 251
rect 404 250 405 251
rect 403 250 404 251
rect 402 250 403 251
rect 401 250 402 251
rect 321 250 322 251
rect 320 250 321 251
rect 319 250 320 251
rect 318 250 319 251
rect 317 250 318 251
rect 316 250 317 251
rect 315 250 316 251
rect 314 250 315 251
rect 313 250 314 251
rect 312 250 313 251
rect 311 250 312 251
rect 310 250 311 251
rect 309 250 310 251
rect 308 250 309 251
rect 307 250 308 251
rect 306 250 307 251
rect 305 250 306 251
rect 304 250 305 251
rect 303 250 304 251
rect 302 250 303 251
rect 301 250 302 251
rect 300 250 301 251
rect 299 250 300 251
rect 298 250 299 251
rect 297 250 298 251
rect 296 250 297 251
rect 295 250 296 251
rect 294 250 295 251
rect 293 250 294 251
rect 292 250 293 251
rect 291 250 292 251
rect 290 250 291 251
rect 289 250 290 251
rect 288 250 289 251
rect 287 250 288 251
rect 286 250 287 251
rect 285 250 286 251
rect 284 250 285 251
rect 283 250 284 251
rect 282 250 283 251
rect 281 250 282 251
rect 280 250 281 251
rect 279 250 280 251
rect 278 250 279 251
rect 277 250 278 251
rect 276 250 277 251
rect 275 250 276 251
rect 274 250 275 251
rect 273 250 274 251
rect 272 250 273 251
rect 271 250 272 251
rect 270 250 271 251
rect 269 250 270 251
rect 268 250 269 251
rect 267 250 268 251
rect 266 250 267 251
rect 265 250 266 251
rect 264 250 265 251
rect 263 250 264 251
rect 262 250 263 251
rect 261 250 262 251
rect 260 250 261 251
rect 259 250 260 251
rect 258 250 259 251
rect 257 250 258 251
rect 256 250 257 251
rect 255 250 256 251
rect 254 250 255 251
rect 253 250 254 251
rect 252 250 253 251
rect 251 250 252 251
rect 250 250 251 251
rect 249 250 250 251
rect 248 250 249 251
rect 247 250 248 251
rect 246 250 247 251
rect 245 250 246 251
rect 244 250 245 251
rect 243 250 244 251
rect 242 250 243 251
rect 241 250 242 251
rect 240 250 241 251
rect 239 250 240 251
rect 238 250 239 251
rect 237 250 238 251
rect 236 250 237 251
rect 235 250 236 251
rect 234 250 235 251
rect 158 250 159 251
rect 157 250 158 251
rect 156 250 157 251
rect 155 250 156 251
rect 154 250 155 251
rect 153 250 154 251
rect 152 250 153 251
rect 151 250 152 251
rect 150 250 151 251
rect 149 250 150 251
rect 148 250 149 251
rect 147 250 148 251
rect 146 250 147 251
rect 145 250 146 251
rect 144 250 145 251
rect 143 250 144 251
rect 142 250 143 251
rect 141 250 142 251
rect 140 250 141 251
rect 139 250 140 251
rect 138 250 139 251
rect 137 250 138 251
rect 136 250 137 251
rect 135 250 136 251
rect 134 250 135 251
rect 133 250 134 251
rect 132 250 133 251
rect 131 250 132 251
rect 130 250 131 251
rect 129 250 130 251
rect 128 250 129 251
rect 127 250 128 251
rect 126 250 127 251
rect 125 250 126 251
rect 124 250 125 251
rect 123 250 124 251
rect 122 250 123 251
rect 109 250 110 251
rect 108 250 109 251
rect 107 250 108 251
rect 106 250 107 251
rect 105 250 106 251
rect 104 250 105 251
rect 103 250 104 251
rect 102 250 103 251
rect 101 250 102 251
rect 100 250 101 251
rect 99 250 100 251
rect 98 250 99 251
rect 97 250 98 251
rect 96 250 97 251
rect 95 250 96 251
rect 94 250 95 251
rect 93 250 94 251
rect 92 250 93 251
rect 91 250 92 251
rect 90 250 91 251
rect 89 250 90 251
rect 88 250 89 251
rect 87 250 88 251
rect 86 250 87 251
rect 85 250 86 251
rect 84 250 85 251
rect 83 250 84 251
rect 82 250 83 251
rect 81 250 82 251
rect 80 250 81 251
rect 79 250 80 251
rect 78 250 79 251
rect 77 250 78 251
rect 76 250 77 251
rect 75 250 76 251
rect 74 250 75 251
rect 73 250 74 251
rect 72 250 73 251
rect 71 250 72 251
rect 70 250 71 251
rect 69 250 70 251
rect 68 250 69 251
rect 67 250 68 251
rect 66 250 67 251
rect 65 250 66 251
rect 64 250 65 251
rect 63 250 64 251
rect 62 250 63 251
rect 61 250 62 251
rect 60 250 61 251
rect 59 250 60 251
rect 58 250 59 251
rect 57 250 58 251
rect 56 250 57 251
rect 55 250 56 251
rect 54 250 55 251
rect 53 250 54 251
rect 52 250 53 251
rect 51 250 52 251
rect 50 250 51 251
rect 49 250 50 251
rect 48 250 49 251
rect 47 250 48 251
rect 46 250 47 251
rect 45 250 46 251
rect 44 250 45 251
rect 43 250 44 251
rect 42 250 43 251
rect 41 250 42 251
rect 40 250 41 251
rect 39 250 40 251
rect 38 250 39 251
rect 37 250 38 251
rect 36 250 37 251
rect 35 250 36 251
rect 34 250 35 251
rect 33 250 34 251
rect 32 250 33 251
rect 23 250 24 251
rect 22 250 23 251
rect 21 250 22 251
rect 20 250 21 251
rect 19 250 20 251
rect 18 250 19 251
rect 17 250 18 251
rect 16 250 17 251
rect 15 250 16 251
rect 14 250 15 251
rect 13 250 14 251
rect 12 250 13 251
rect 11 250 12 251
rect 10 250 11 251
rect 9 250 10 251
rect 8 250 9 251
rect 7 250 8 251
rect 6 250 7 251
rect 5 250 6 251
rect 483 251 484 252
rect 482 251 483 252
rect 473 251 474 252
rect 472 251 473 252
rect 471 251 472 252
rect 470 251 471 252
rect 469 251 470 252
rect 468 251 469 252
rect 462 251 463 252
rect 461 251 462 252
rect 424 251 425 252
rect 423 251 424 252
rect 422 251 423 252
rect 421 251 422 252
rect 420 251 421 252
rect 320 251 321 252
rect 319 251 320 252
rect 318 251 319 252
rect 317 251 318 252
rect 316 251 317 252
rect 315 251 316 252
rect 314 251 315 252
rect 313 251 314 252
rect 312 251 313 252
rect 311 251 312 252
rect 310 251 311 252
rect 309 251 310 252
rect 308 251 309 252
rect 307 251 308 252
rect 306 251 307 252
rect 305 251 306 252
rect 304 251 305 252
rect 303 251 304 252
rect 302 251 303 252
rect 301 251 302 252
rect 300 251 301 252
rect 299 251 300 252
rect 298 251 299 252
rect 297 251 298 252
rect 296 251 297 252
rect 295 251 296 252
rect 294 251 295 252
rect 293 251 294 252
rect 292 251 293 252
rect 291 251 292 252
rect 290 251 291 252
rect 289 251 290 252
rect 288 251 289 252
rect 287 251 288 252
rect 286 251 287 252
rect 285 251 286 252
rect 284 251 285 252
rect 283 251 284 252
rect 282 251 283 252
rect 281 251 282 252
rect 280 251 281 252
rect 279 251 280 252
rect 278 251 279 252
rect 277 251 278 252
rect 276 251 277 252
rect 275 251 276 252
rect 274 251 275 252
rect 273 251 274 252
rect 272 251 273 252
rect 271 251 272 252
rect 270 251 271 252
rect 269 251 270 252
rect 268 251 269 252
rect 267 251 268 252
rect 266 251 267 252
rect 265 251 266 252
rect 264 251 265 252
rect 263 251 264 252
rect 262 251 263 252
rect 261 251 262 252
rect 260 251 261 252
rect 259 251 260 252
rect 258 251 259 252
rect 257 251 258 252
rect 256 251 257 252
rect 255 251 256 252
rect 254 251 255 252
rect 253 251 254 252
rect 252 251 253 252
rect 251 251 252 252
rect 250 251 251 252
rect 249 251 250 252
rect 248 251 249 252
rect 247 251 248 252
rect 246 251 247 252
rect 245 251 246 252
rect 244 251 245 252
rect 243 251 244 252
rect 242 251 243 252
rect 241 251 242 252
rect 240 251 241 252
rect 239 251 240 252
rect 238 251 239 252
rect 237 251 238 252
rect 236 251 237 252
rect 235 251 236 252
rect 234 251 235 252
rect 233 251 234 252
rect 159 251 160 252
rect 158 251 159 252
rect 157 251 158 252
rect 156 251 157 252
rect 155 251 156 252
rect 154 251 155 252
rect 153 251 154 252
rect 152 251 153 252
rect 151 251 152 252
rect 150 251 151 252
rect 149 251 150 252
rect 148 251 149 252
rect 147 251 148 252
rect 146 251 147 252
rect 145 251 146 252
rect 144 251 145 252
rect 143 251 144 252
rect 142 251 143 252
rect 141 251 142 252
rect 140 251 141 252
rect 139 251 140 252
rect 138 251 139 252
rect 137 251 138 252
rect 136 251 137 252
rect 135 251 136 252
rect 134 251 135 252
rect 133 251 134 252
rect 132 251 133 252
rect 131 251 132 252
rect 130 251 131 252
rect 129 251 130 252
rect 128 251 129 252
rect 127 251 128 252
rect 126 251 127 252
rect 125 251 126 252
rect 124 251 125 252
rect 123 251 124 252
rect 122 251 123 252
rect 109 251 110 252
rect 108 251 109 252
rect 107 251 108 252
rect 106 251 107 252
rect 105 251 106 252
rect 104 251 105 252
rect 103 251 104 252
rect 102 251 103 252
rect 101 251 102 252
rect 100 251 101 252
rect 99 251 100 252
rect 98 251 99 252
rect 97 251 98 252
rect 96 251 97 252
rect 95 251 96 252
rect 94 251 95 252
rect 93 251 94 252
rect 92 251 93 252
rect 91 251 92 252
rect 90 251 91 252
rect 89 251 90 252
rect 88 251 89 252
rect 87 251 88 252
rect 86 251 87 252
rect 85 251 86 252
rect 84 251 85 252
rect 83 251 84 252
rect 82 251 83 252
rect 81 251 82 252
rect 80 251 81 252
rect 79 251 80 252
rect 78 251 79 252
rect 77 251 78 252
rect 76 251 77 252
rect 75 251 76 252
rect 74 251 75 252
rect 73 251 74 252
rect 72 251 73 252
rect 71 251 72 252
rect 70 251 71 252
rect 69 251 70 252
rect 68 251 69 252
rect 67 251 68 252
rect 66 251 67 252
rect 65 251 66 252
rect 64 251 65 252
rect 63 251 64 252
rect 62 251 63 252
rect 61 251 62 252
rect 60 251 61 252
rect 59 251 60 252
rect 58 251 59 252
rect 57 251 58 252
rect 56 251 57 252
rect 55 251 56 252
rect 54 251 55 252
rect 53 251 54 252
rect 52 251 53 252
rect 51 251 52 252
rect 50 251 51 252
rect 49 251 50 252
rect 48 251 49 252
rect 47 251 48 252
rect 46 251 47 252
rect 45 251 46 252
rect 44 251 45 252
rect 43 251 44 252
rect 42 251 43 252
rect 41 251 42 252
rect 40 251 41 252
rect 39 251 40 252
rect 38 251 39 252
rect 37 251 38 252
rect 36 251 37 252
rect 35 251 36 252
rect 34 251 35 252
rect 33 251 34 252
rect 23 251 24 252
rect 22 251 23 252
rect 21 251 22 252
rect 20 251 21 252
rect 19 251 20 252
rect 18 251 19 252
rect 17 251 18 252
rect 16 251 17 252
rect 15 251 16 252
rect 14 251 15 252
rect 13 251 14 252
rect 12 251 13 252
rect 11 251 12 252
rect 10 251 11 252
rect 9 251 10 252
rect 8 251 9 252
rect 7 251 8 252
rect 6 251 7 252
rect 5 251 6 252
rect 483 252 484 253
rect 482 252 483 253
rect 474 252 475 253
rect 473 252 474 253
rect 472 252 473 253
rect 471 252 472 253
rect 470 252 471 253
rect 469 252 470 253
rect 462 252 463 253
rect 461 252 462 253
rect 423 252 424 253
rect 422 252 423 253
rect 421 252 422 253
rect 420 252 421 253
rect 318 252 319 253
rect 317 252 318 253
rect 316 252 317 253
rect 315 252 316 253
rect 314 252 315 253
rect 313 252 314 253
rect 312 252 313 253
rect 311 252 312 253
rect 310 252 311 253
rect 309 252 310 253
rect 308 252 309 253
rect 307 252 308 253
rect 306 252 307 253
rect 305 252 306 253
rect 304 252 305 253
rect 303 252 304 253
rect 302 252 303 253
rect 301 252 302 253
rect 300 252 301 253
rect 299 252 300 253
rect 298 252 299 253
rect 297 252 298 253
rect 296 252 297 253
rect 295 252 296 253
rect 294 252 295 253
rect 293 252 294 253
rect 292 252 293 253
rect 291 252 292 253
rect 290 252 291 253
rect 289 252 290 253
rect 288 252 289 253
rect 287 252 288 253
rect 286 252 287 253
rect 285 252 286 253
rect 284 252 285 253
rect 283 252 284 253
rect 282 252 283 253
rect 281 252 282 253
rect 280 252 281 253
rect 279 252 280 253
rect 278 252 279 253
rect 277 252 278 253
rect 276 252 277 253
rect 275 252 276 253
rect 274 252 275 253
rect 273 252 274 253
rect 272 252 273 253
rect 271 252 272 253
rect 270 252 271 253
rect 269 252 270 253
rect 268 252 269 253
rect 267 252 268 253
rect 266 252 267 253
rect 265 252 266 253
rect 264 252 265 253
rect 263 252 264 253
rect 262 252 263 253
rect 261 252 262 253
rect 260 252 261 253
rect 259 252 260 253
rect 258 252 259 253
rect 257 252 258 253
rect 256 252 257 253
rect 255 252 256 253
rect 254 252 255 253
rect 253 252 254 253
rect 252 252 253 253
rect 251 252 252 253
rect 250 252 251 253
rect 249 252 250 253
rect 248 252 249 253
rect 247 252 248 253
rect 246 252 247 253
rect 245 252 246 253
rect 244 252 245 253
rect 243 252 244 253
rect 242 252 243 253
rect 241 252 242 253
rect 240 252 241 253
rect 239 252 240 253
rect 238 252 239 253
rect 237 252 238 253
rect 236 252 237 253
rect 235 252 236 253
rect 234 252 235 253
rect 233 252 234 253
rect 160 252 161 253
rect 159 252 160 253
rect 158 252 159 253
rect 157 252 158 253
rect 156 252 157 253
rect 155 252 156 253
rect 154 252 155 253
rect 153 252 154 253
rect 152 252 153 253
rect 151 252 152 253
rect 150 252 151 253
rect 149 252 150 253
rect 148 252 149 253
rect 147 252 148 253
rect 146 252 147 253
rect 145 252 146 253
rect 144 252 145 253
rect 143 252 144 253
rect 142 252 143 253
rect 141 252 142 253
rect 140 252 141 253
rect 139 252 140 253
rect 138 252 139 253
rect 137 252 138 253
rect 136 252 137 253
rect 135 252 136 253
rect 134 252 135 253
rect 133 252 134 253
rect 132 252 133 253
rect 131 252 132 253
rect 130 252 131 253
rect 129 252 130 253
rect 128 252 129 253
rect 127 252 128 253
rect 126 252 127 253
rect 125 252 126 253
rect 124 252 125 253
rect 123 252 124 253
rect 110 252 111 253
rect 109 252 110 253
rect 108 252 109 253
rect 107 252 108 253
rect 106 252 107 253
rect 105 252 106 253
rect 104 252 105 253
rect 103 252 104 253
rect 102 252 103 253
rect 101 252 102 253
rect 100 252 101 253
rect 99 252 100 253
rect 98 252 99 253
rect 97 252 98 253
rect 96 252 97 253
rect 95 252 96 253
rect 94 252 95 253
rect 93 252 94 253
rect 92 252 93 253
rect 91 252 92 253
rect 90 252 91 253
rect 89 252 90 253
rect 88 252 89 253
rect 87 252 88 253
rect 86 252 87 253
rect 85 252 86 253
rect 84 252 85 253
rect 83 252 84 253
rect 82 252 83 253
rect 81 252 82 253
rect 80 252 81 253
rect 79 252 80 253
rect 78 252 79 253
rect 77 252 78 253
rect 76 252 77 253
rect 75 252 76 253
rect 74 252 75 253
rect 73 252 74 253
rect 72 252 73 253
rect 71 252 72 253
rect 70 252 71 253
rect 69 252 70 253
rect 68 252 69 253
rect 67 252 68 253
rect 66 252 67 253
rect 65 252 66 253
rect 64 252 65 253
rect 63 252 64 253
rect 62 252 63 253
rect 61 252 62 253
rect 60 252 61 253
rect 59 252 60 253
rect 58 252 59 253
rect 57 252 58 253
rect 56 252 57 253
rect 55 252 56 253
rect 54 252 55 253
rect 53 252 54 253
rect 52 252 53 253
rect 51 252 52 253
rect 50 252 51 253
rect 49 252 50 253
rect 48 252 49 253
rect 47 252 48 253
rect 46 252 47 253
rect 45 252 46 253
rect 44 252 45 253
rect 43 252 44 253
rect 42 252 43 253
rect 41 252 42 253
rect 40 252 41 253
rect 39 252 40 253
rect 38 252 39 253
rect 37 252 38 253
rect 36 252 37 253
rect 35 252 36 253
rect 34 252 35 253
rect 33 252 34 253
rect 23 252 24 253
rect 22 252 23 253
rect 21 252 22 253
rect 20 252 21 253
rect 19 252 20 253
rect 18 252 19 253
rect 17 252 18 253
rect 16 252 17 253
rect 15 252 16 253
rect 14 252 15 253
rect 13 252 14 253
rect 12 252 13 253
rect 11 252 12 253
rect 10 252 11 253
rect 9 252 10 253
rect 8 252 9 253
rect 7 252 8 253
rect 6 252 7 253
rect 5 252 6 253
rect 483 253 484 254
rect 482 253 483 254
rect 474 253 475 254
rect 473 253 474 254
rect 472 253 473 254
rect 471 253 472 254
rect 470 253 471 254
rect 462 253 463 254
rect 461 253 462 254
rect 422 253 423 254
rect 421 253 422 254
rect 420 253 421 254
rect 317 253 318 254
rect 316 253 317 254
rect 315 253 316 254
rect 314 253 315 254
rect 313 253 314 254
rect 312 253 313 254
rect 311 253 312 254
rect 310 253 311 254
rect 309 253 310 254
rect 308 253 309 254
rect 307 253 308 254
rect 306 253 307 254
rect 305 253 306 254
rect 304 253 305 254
rect 303 253 304 254
rect 302 253 303 254
rect 301 253 302 254
rect 300 253 301 254
rect 299 253 300 254
rect 298 253 299 254
rect 297 253 298 254
rect 296 253 297 254
rect 295 253 296 254
rect 294 253 295 254
rect 293 253 294 254
rect 292 253 293 254
rect 291 253 292 254
rect 290 253 291 254
rect 289 253 290 254
rect 288 253 289 254
rect 287 253 288 254
rect 286 253 287 254
rect 285 253 286 254
rect 284 253 285 254
rect 283 253 284 254
rect 282 253 283 254
rect 281 253 282 254
rect 280 253 281 254
rect 279 253 280 254
rect 278 253 279 254
rect 277 253 278 254
rect 276 253 277 254
rect 275 253 276 254
rect 274 253 275 254
rect 273 253 274 254
rect 272 253 273 254
rect 271 253 272 254
rect 270 253 271 254
rect 269 253 270 254
rect 268 253 269 254
rect 267 253 268 254
rect 266 253 267 254
rect 265 253 266 254
rect 264 253 265 254
rect 263 253 264 254
rect 262 253 263 254
rect 261 253 262 254
rect 260 253 261 254
rect 259 253 260 254
rect 258 253 259 254
rect 257 253 258 254
rect 256 253 257 254
rect 255 253 256 254
rect 254 253 255 254
rect 253 253 254 254
rect 252 253 253 254
rect 251 253 252 254
rect 250 253 251 254
rect 249 253 250 254
rect 248 253 249 254
rect 247 253 248 254
rect 246 253 247 254
rect 245 253 246 254
rect 244 253 245 254
rect 243 253 244 254
rect 242 253 243 254
rect 241 253 242 254
rect 240 253 241 254
rect 239 253 240 254
rect 238 253 239 254
rect 237 253 238 254
rect 236 253 237 254
rect 235 253 236 254
rect 234 253 235 254
rect 233 253 234 254
rect 161 253 162 254
rect 160 253 161 254
rect 159 253 160 254
rect 158 253 159 254
rect 157 253 158 254
rect 156 253 157 254
rect 155 253 156 254
rect 154 253 155 254
rect 153 253 154 254
rect 152 253 153 254
rect 151 253 152 254
rect 150 253 151 254
rect 149 253 150 254
rect 148 253 149 254
rect 147 253 148 254
rect 146 253 147 254
rect 145 253 146 254
rect 144 253 145 254
rect 143 253 144 254
rect 142 253 143 254
rect 141 253 142 254
rect 140 253 141 254
rect 139 253 140 254
rect 138 253 139 254
rect 137 253 138 254
rect 136 253 137 254
rect 135 253 136 254
rect 134 253 135 254
rect 133 253 134 254
rect 132 253 133 254
rect 131 253 132 254
rect 130 253 131 254
rect 129 253 130 254
rect 128 253 129 254
rect 127 253 128 254
rect 126 253 127 254
rect 125 253 126 254
rect 124 253 125 254
rect 123 253 124 254
rect 110 253 111 254
rect 109 253 110 254
rect 108 253 109 254
rect 107 253 108 254
rect 106 253 107 254
rect 105 253 106 254
rect 104 253 105 254
rect 103 253 104 254
rect 102 253 103 254
rect 101 253 102 254
rect 100 253 101 254
rect 99 253 100 254
rect 98 253 99 254
rect 97 253 98 254
rect 96 253 97 254
rect 95 253 96 254
rect 94 253 95 254
rect 93 253 94 254
rect 92 253 93 254
rect 91 253 92 254
rect 90 253 91 254
rect 89 253 90 254
rect 88 253 89 254
rect 87 253 88 254
rect 86 253 87 254
rect 85 253 86 254
rect 84 253 85 254
rect 83 253 84 254
rect 82 253 83 254
rect 81 253 82 254
rect 80 253 81 254
rect 79 253 80 254
rect 78 253 79 254
rect 77 253 78 254
rect 76 253 77 254
rect 75 253 76 254
rect 74 253 75 254
rect 73 253 74 254
rect 72 253 73 254
rect 71 253 72 254
rect 70 253 71 254
rect 69 253 70 254
rect 68 253 69 254
rect 67 253 68 254
rect 66 253 67 254
rect 65 253 66 254
rect 64 253 65 254
rect 63 253 64 254
rect 62 253 63 254
rect 61 253 62 254
rect 60 253 61 254
rect 59 253 60 254
rect 58 253 59 254
rect 57 253 58 254
rect 56 253 57 254
rect 55 253 56 254
rect 54 253 55 254
rect 53 253 54 254
rect 52 253 53 254
rect 51 253 52 254
rect 50 253 51 254
rect 49 253 50 254
rect 48 253 49 254
rect 47 253 48 254
rect 46 253 47 254
rect 45 253 46 254
rect 44 253 45 254
rect 43 253 44 254
rect 42 253 43 254
rect 41 253 42 254
rect 40 253 41 254
rect 39 253 40 254
rect 38 253 39 254
rect 37 253 38 254
rect 36 253 37 254
rect 35 253 36 254
rect 34 253 35 254
rect 33 253 34 254
rect 23 253 24 254
rect 22 253 23 254
rect 21 253 22 254
rect 20 253 21 254
rect 19 253 20 254
rect 18 253 19 254
rect 17 253 18 254
rect 16 253 17 254
rect 15 253 16 254
rect 14 253 15 254
rect 13 253 14 254
rect 12 253 13 254
rect 11 253 12 254
rect 10 253 11 254
rect 9 253 10 254
rect 8 253 9 254
rect 7 253 8 254
rect 6 253 7 254
rect 5 253 6 254
rect 483 254 484 255
rect 482 254 483 255
rect 475 254 476 255
rect 474 254 475 255
rect 473 254 474 255
rect 472 254 473 255
rect 471 254 472 255
rect 470 254 471 255
rect 462 254 463 255
rect 461 254 462 255
rect 422 254 423 255
rect 421 254 422 255
rect 315 254 316 255
rect 314 254 315 255
rect 313 254 314 255
rect 312 254 313 255
rect 311 254 312 255
rect 310 254 311 255
rect 309 254 310 255
rect 308 254 309 255
rect 307 254 308 255
rect 306 254 307 255
rect 305 254 306 255
rect 304 254 305 255
rect 303 254 304 255
rect 302 254 303 255
rect 301 254 302 255
rect 300 254 301 255
rect 299 254 300 255
rect 298 254 299 255
rect 297 254 298 255
rect 296 254 297 255
rect 295 254 296 255
rect 294 254 295 255
rect 293 254 294 255
rect 292 254 293 255
rect 291 254 292 255
rect 290 254 291 255
rect 289 254 290 255
rect 288 254 289 255
rect 287 254 288 255
rect 286 254 287 255
rect 285 254 286 255
rect 284 254 285 255
rect 283 254 284 255
rect 282 254 283 255
rect 281 254 282 255
rect 280 254 281 255
rect 279 254 280 255
rect 278 254 279 255
rect 277 254 278 255
rect 276 254 277 255
rect 275 254 276 255
rect 274 254 275 255
rect 273 254 274 255
rect 272 254 273 255
rect 271 254 272 255
rect 270 254 271 255
rect 269 254 270 255
rect 268 254 269 255
rect 267 254 268 255
rect 266 254 267 255
rect 265 254 266 255
rect 264 254 265 255
rect 263 254 264 255
rect 262 254 263 255
rect 261 254 262 255
rect 260 254 261 255
rect 259 254 260 255
rect 258 254 259 255
rect 257 254 258 255
rect 256 254 257 255
rect 255 254 256 255
rect 254 254 255 255
rect 253 254 254 255
rect 252 254 253 255
rect 251 254 252 255
rect 250 254 251 255
rect 249 254 250 255
rect 248 254 249 255
rect 247 254 248 255
rect 246 254 247 255
rect 245 254 246 255
rect 244 254 245 255
rect 243 254 244 255
rect 242 254 243 255
rect 241 254 242 255
rect 240 254 241 255
rect 239 254 240 255
rect 238 254 239 255
rect 237 254 238 255
rect 236 254 237 255
rect 235 254 236 255
rect 234 254 235 255
rect 233 254 234 255
rect 162 254 163 255
rect 161 254 162 255
rect 160 254 161 255
rect 159 254 160 255
rect 158 254 159 255
rect 157 254 158 255
rect 156 254 157 255
rect 155 254 156 255
rect 154 254 155 255
rect 153 254 154 255
rect 152 254 153 255
rect 151 254 152 255
rect 150 254 151 255
rect 149 254 150 255
rect 148 254 149 255
rect 147 254 148 255
rect 146 254 147 255
rect 145 254 146 255
rect 144 254 145 255
rect 143 254 144 255
rect 142 254 143 255
rect 141 254 142 255
rect 140 254 141 255
rect 139 254 140 255
rect 138 254 139 255
rect 137 254 138 255
rect 136 254 137 255
rect 135 254 136 255
rect 134 254 135 255
rect 133 254 134 255
rect 132 254 133 255
rect 131 254 132 255
rect 130 254 131 255
rect 129 254 130 255
rect 128 254 129 255
rect 127 254 128 255
rect 126 254 127 255
rect 125 254 126 255
rect 124 254 125 255
rect 123 254 124 255
rect 110 254 111 255
rect 109 254 110 255
rect 108 254 109 255
rect 107 254 108 255
rect 106 254 107 255
rect 105 254 106 255
rect 104 254 105 255
rect 103 254 104 255
rect 102 254 103 255
rect 101 254 102 255
rect 100 254 101 255
rect 99 254 100 255
rect 98 254 99 255
rect 97 254 98 255
rect 96 254 97 255
rect 95 254 96 255
rect 94 254 95 255
rect 93 254 94 255
rect 92 254 93 255
rect 91 254 92 255
rect 90 254 91 255
rect 89 254 90 255
rect 88 254 89 255
rect 87 254 88 255
rect 86 254 87 255
rect 85 254 86 255
rect 84 254 85 255
rect 83 254 84 255
rect 82 254 83 255
rect 81 254 82 255
rect 80 254 81 255
rect 79 254 80 255
rect 78 254 79 255
rect 77 254 78 255
rect 76 254 77 255
rect 75 254 76 255
rect 74 254 75 255
rect 73 254 74 255
rect 72 254 73 255
rect 71 254 72 255
rect 70 254 71 255
rect 69 254 70 255
rect 68 254 69 255
rect 67 254 68 255
rect 66 254 67 255
rect 65 254 66 255
rect 64 254 65 255
rect 63 254 64 255
rect 62 254 63 255
rect 61 254 62 255
rect 60 254 61 255
rect 59 254 60 255
rect 58 254 59 255
rect 57 254 58 255
rect 56 254 57 255
rect 55 254 56 255
rect 54 254 55 255
rect 53 254 54 255
rect 52 254 53 255
rect 51 254 52 255
rect 50 254 51 255
rect 49 254 50 255
rect 48 254 49 255
rect 47 254 48 255
rect 46 254 47 255
rect 45 254 46 255
rect 44 254 45 255
rect 43 254 44 255
rect 42 254 43 255
rect 41 254 42 255
rect 40 254 41 255
rect 39 254 40 255
rect 38 254 39 255
rect 37 254 38 255
rect 36 254 37 255
rect 35 254 36 255
rect 34 254 35 255
rect 23 254 24 255
rect 22 254 23 255
rect 21 254 22 255
rect 20 254 21 255
rect 19 254 20 255
rect 18 254 19 255
rect 17 254 18 255
rect 16 254 17 255
rect 15 254 16 255
rect 14 254 15 255
rect 13 254 14 255
rect 12 254 13 255
rect 11 254 12 255
rect 10 254 11 255
rect 9 254 10 255
rect 8 254 9 255
rect 7 254 8 255
rect 6 254 7 255
rect 5 254 6 255
rect 482 255 483 256
rect 481 255 482 256
rect 476 255 477 256
rect 475 255 476 256
rect 474 255 475 256
rect 473 255 474 256
rect 472 255 473 256
rect 471 255 472 256
rect 462 255 463 256
rect 461 255 462 256
rect 314 255 315 256
rect 313 255 314 256
rect 312 255 313 256
rect 311 255 312 256
rect 310 255 311 256
rect 309 255 310 256
rect 308 255 309 256
rect 307 255 308 256
rect 306 255 307 256
rect 305 255 306 256
rect 304 255 305 256
rect 303 255 304 256
rect 302 255 303 256
rect 301 255 302 256
rect 300 255 301 256
rect 299 255 300 256
rect 298 255 299 256
rect 297 255 298 256
rect 296 255 297 256
rect 295 255 296 256
rect 294 255 295 256
rect 293 255 294 256
rect 292 255 293 256
rect 291 255 292 256
rect 290 255 291 256
rect 289 255 290 256
rect 288 255 289 256
rect 287 255 288 256
rect 286 255 287 256
rect 285 255 286 256
rect 284 255 285 256
rect 283 255 284 256
rect 282 255 283 256
rect 281 255 282 256
rect 280 255 281 256
rect 279 255 280 256
rect 278 255 279 256
rect 277 255 278 256
rect 276 255 277 256
rect 275 255 276 256
rect 274 255 275 256
rect 273 255 274 256
rect 272 255 273 256
rect 271 255 272 256
rect 270 255 271 256
rect 269 255 270 256
rect 268 255 269 256
rect 267 255 268 256
rect 266 255 267 256
rect 265 255 266 256
rect 264 255 265 256
rect 263 255 264 256
rect 262 255 263 256
rect 261 255 262 256
rect 260 255 261 256
rect 259 255 260 256
rect 258 255 259 256
rect 257 255 258 256
rect 256 255 257 256
rect 255 255 256 256
rect 254 255 255 256
rect 253 255 254 256
rect 252 255 253 256
rect 251 255 252 256
rect 250 255 251 256
rect 249 255 250 256
rect 248 255 249 256
rect 247 255 248 256
rect 246 255 247 256
rect 245 255 246 256
rect 244 255 245 256
rect 243 255 244 256
rect 242 255 243 256
rect 241 255 242 256
rect 240 255 241 256
rect 239 255 240 256
rect 238 255 239 256
rect 237 255 238 256
rect 236 255 237 256
rect 235 255 236 256
rect 234 255 235 256
rect 233 255 234 256
rect 232 255 233 256
rect 164 255 165 256
rect 163 255 164 256
rect 162 255 163 256
rect 161 255 162 256
rect 160 255 161 256
rect 159 255 160 256
rect 158 255 159 256
rect 157 255 158 256
rect 156 255 157 256
rect 155 255 156 256
rect 154 255 155 256
rect 153 255 154 256
rect 152 255 153 256
rect 151 255 152 256
rect 150 255 151 256
rect 149 255 150 256
rect 148 255 149 256
rect 147 255 148 256
rect 146 255 147 256
rect 145 255 146 256
rect 144 255 145 256
rect 143 255 144 256
rect 142 255 143 256
rect 141 255 142 256
rect 140 255 141 256
rect 139 255 140 256
rect 138 255 139 256
rect 137 255 138 256
rect 136 255 137 256
rect 135 255 136 256
rect 134 255 135 256
rect 133 255 134 256
rect 132 255 133 256
rect 131 255 132 256
rect 130 255 131 256
rect 129 255 130 256
rect 128 255 129 256
rect 127 255 128 256
rect 126 255 127 256
rect 125 255 126 256
rect 124 255 125 256
rect 123 255 124 256
rect 110 255 111 256
rect 109 255 110 256
rect 108 255 109 256
rect 107 255 108 256
rect 106 255 107 256
rect 105 255 106 256
rect 104 255 105 256
rect 103 255 104 256
rect 102 255 103 256
rect 101 255 102 256
rect 100 255 101 256
rect 99 255 100 256
rect 98 255 99 256
rect 97 255 98 256
rect 96 255 97 256
rect 95 255 96 256
rect 94 255 95 256
rect 93 255 94 256
rect 92 255 93 256
rect 91 255 92 256
rect 90 255 91 256
rect 89 255 90 256
rect 88 255 89 256
rect 87 255 88 256
rect 86 255 87 256
rect 85 255 86 256
rect 84 255 85 256
rect 83 255 84 256
rect 82 255 83 256
rect 81 255 82 256
rect 80 255 81 256
rect 79 255 80 256
rect 78 255 79 256
rect 77 255 78 256
rect 76 255 77 256
rect 75 255 76 256
rect 74 255 75 256
rect 73 255 74 256
rect 72 255 73 256
rect 71 255 72 256
rect 70 255 71 256
rect 69 255 70 256
rect 68 255 69 256
rect 67 255 68 256
rect 66 255 67 256
rect 65 255 66 256
rect 64 255 65 256
rect 63 255 64 256
rect 62 255 63 256
rect 61 255 62 256
rect 60 255 61 256
rect 59 255 60 256
rect 58 255 59 256
rect 57 255 58 256
rect 56 255 57 256
rect 55 255 56 256
rect 54 255 55 256
rect 53 255 54 256
rect 52 255 53 256
rect 51 255 52 256
rect 50 255 51 256
rect 49 255 50 256
rect 48 255 49 256
rect 47 255 48 256
rect 46 255 47 256
rect 45 255 46 256
rect 44 255 45 256
rect 43 255 44 256
rect 42 255 43 256
rect 41 255 42 256
rect 40 255 41 256
rect 39 255 40 256
rect 38 255 39 256
rect 37 255 38 256
rect 36 255 37 256
rect 35 255 36 256
rect 34 255 35 256
rect 23 255 24 256
rect 22 255 23 256
rect 21 255 22 256
rect 20 255 21 256
rect 19 255 20 256
rect 18 255 19 256
rect 17 255 18 256
rect 16 255 17 256
rect 15 255 16 256
rect 14 255 15 256
rect 13 255 14 256
rect 12 255 13 256
rect 11 255 12 256
rect 10 255 11 256
rect 9 255 10 256
rect 8 255 9 256
rect 7 255 8 256
rect 6 255 7 256
rect 5 255 6 256
rect 482 256 483 257
rect 481 256 482 257
rect 480 256 481 257
rect 479 256 480 257
rect 478 256 479 257
rect 477 256 478 257
rect 476 256 477 257
rect 475 256 476 257
rect 474 256 475 257
rect 473 256 474 257
rect 472 256 473 257
rect 471 256 472 257
rect 463 256 464 257
rect 462 256 463 257
rect 461 256 462 257
rect 313 256 314 257
rect 312 256 313 257
rect 311 256 312 257
rect 310 256 311 257
rect 309 256 310 257
rect 308 256 309 257
rect 307 256 308 257
rect 306 256 307 257
rect 305 256 306 257
rect 304 256 305 257
rect 303 256 304 257
rect 302 256 303 257
rect 301 256 302 257
rect 300 256 301 257
rect 299 256 300 257
rect 298 256 299 257
rect 297 256 298 257
rect 296 256 297 257
rect 295 256 296 257
rect 294 256 295 257
rect 293 256 294 257
rect 292 256 293 257
rect 291 256 292 257
rect 290 256 291 257
rect 289 256 290 257
rect 288 256 289 257
rect 287 256 288 257
rect 286 256 287 257
rect 285 256 286 257
rect 284 256 285 257
rect 283 256 284 257
rect 282 256 283 257
rect 281 256 282 257
rect 280 256 281 257
rect 279 256 280 257
rect 278 256 279 257
rect 277 256 278 257
rect 276 256 277 257
rect 275 256 276 257
rect 274 256 275 257
rect 273 256 274 257
rect 272 256 273 257
rect 271 256 272 257
rect 270 256 271 257
rect 269 256 270 257
rect 268 256 269 257
rect 267 256 268 257
rect 266 256 267 257
rect 265 256 266 257
rect 264 256 265 257
rect 263 256 264 257
rect 262 256 263 257
rect 261 256 262 257
rect 260 256 261 257
rect 259 256 260 257
rect 258 256 259 257
rect 257 256 258 257
rect 256 256 257 257
rect 255 256 256 257
rect 254 256 255 257
rect 253 256 254 257
rect 252 256 253 257
rect 251 256 252 257
rect 250 256 251 257
rect 249 256 250 257
rect 248 256 249 257
rect 247 256 248 257
rect 246 256 247 257
rect 245 256 246 257
rect 244 256 245 257
rect 243 256 244 257
rect 242 256 243 257
rect 241 256 242 257
rect 240 256 241 257
rect 239 256 240 257
rect 238 256 239 257
rect 237 256 238 257
rect 236 256 237 257
rect 235 256 236 257
rect 234 256 235 257
rect 233 256 234 257
rect 232 256 233 257
rect 166 256 167 257
rect 165 256 166 257
rect 164 256 165 257
rect 163 256 164 257
rect 162 256 163 257
rect 161 256 162 257
rect 160 256 161 257
rect 159 256 160 257
rect 158 256 159 257
rect 157 256 158 257
rect 156 256 157 257
rect 155 256 156 257
rect 154 256 155 257
rect 153 256 154 257
rect 152 256 153 257
rect 151 256 152 257
rect 150 256 151 257
rect 149 256 150 257
rect 148 256 149 257
rect 147 256 148 257
rect 146 256 147 257
rect 145 256 146 257
rect 144 256 145 257
rect 143 256 144 257
rect 142 256 143 257
rect 141 256 142 257
rect 140 256 141 257
rect 139 256 140 257
rect 138 256 139 257
rect 137 256 138 257
rect 136 256 137 257
rect 135 256 136 257
rect 134 256 135 257
rect 133 256 134 257
rect 132 256 133 257
rect 131 256 132 257
rect 130 256 131 257
rect 129 256 130 257
rect 128 256 129 257
rect 127 256 128 257
rect 126 256 127 257
rect 125 256 126 257
rect 124 256 125 257
rect 123 256 124 257
rect 111 256 112 257
rect 110 256 111 257
rect 109 256 110 257
rect 108 256 109 257
rect 107 256 108 257
rect 106 256 107 257
rect 105 256 106 257
rect 104 256 105 257
rect 103 256 104 257
rect 102 256 103 257
rect 101 256 102 257
rect 100 256 101 257
rect 99 256 100 257
rect 98 256 99 257
rect 97 256 98 257
rect 96 256 97 257
rect 95 256 96 257
rect 94 256 95 257
rect 93 256 94 257
rect 92 256 93 257
rect 91 256 92 257
rect 90 256 91 257
rect 89 256 90 257
rect 88 256 89 257
rect 87 256 88 257
rect 86 256 87 257
rect 85 256 86 257
rect 84 256 85 257
rect 83 256 84 257
rect 82 256 83 257
rect 81 256 82 257
rect 80 256 81 257
rect 79 256 80 257
rect 78 256 79 257
rect 77 256 78 257
rect 76 256 77 257
rect 75 256 76 257
rect 74 256 75 257
rect 73 256 74 257
rect 72 256 73 257
rect 71 256 72 257
rect 70 256 71 257
rect 69 256 70 257
rect 68 256 69 257
rect 67 256 68 257
rect 66 256 67 257
rect 65 256 66 257
rect 64 256 65 257
rect 63 256 64 257
rect 62 256 63 257
rect 61 256 62 257
rect 60 256 61 257
rect 56 256 57 257
rect 55 256 56 257
rect 54 256 55 257
rect 53 256 54 257
rect 52 256 53 257
rect 51 256 52 257
rect 50 256 51 257
rect 49 256 50 257
rect 48 256 49 257
rect 47 256 48 257
rect 46 256 47 257
rect 45 256 46 257
rect 44 256 45 257
rect 43 256 44 257
rect 42 256 43 257
rect 41 256 42 257
rect 40 256 41 257
rect 39 256 40 257
rect 38 256 39 257
rect 37 256 38 257
rect 36 256 37 257
rect 35 256 36 257
rect 34 256 35 257
rect 24 256 25 257
rect 23 256 24 257
rect 22 256 23 257
rect 21 256 22 257
rect 20 256 21 257
rect 19 256 20 257
rect 18 256 19 257
rect 17 256 18 257
rect 16 256 17 257
rect 15 256 16 257
rect 14 256 15 257
rect 13 256 14 257
rect 12 256 13 257
rect 11 256 12 257
rect 10 256 11 257
rect 9 256 10 257
rect 8 256 9 257
rect 7 256 8 257
rect 6 256 7 257
rect 5 256 6 257
rect 481 257 482 258
rect 480 257 481 258
rect 479 257 480 258
rect 478 257 479 258
rect 477 257 478 258
rect 476 257 477 258
rect 475 257 476 258
rect 474 257 475 258
rect 473 257 474 258
rect 472 257 473 258
rect 465 257 466 258
rect 464 257 465 258
rect 463 257 464 258
rect 462 257 463 258
rect 311 257 312 258
rect 310 257 311 258
rect 309 257 310 258
rect 308 257 309 258
rect 307 257 308 258
rect 306 257 307 258
rect 305 257 306 258
rect 304 257 305 258
rect 303 257 304 258
rect 302 257 303 258
rect 301 257 302 258
rect 300 257 301 258
rect 299 257 300 258
rect 298 257 299 258
rect 297 257 298 258
rect 296 257 297 258
rect 295 257 296 258
rect 294 257 295 258
rect 293 257 294 258
rect 292 257 293 258
rect 291 257 292 258
rect 290 257 291 258
rect 289 257 290 258
rect 288 257 289 258
rect 287 257 288 258
rect 286 257 287 258
rect 285 257 286 258
rect 284 257 285 258
rect 283 257 284 258
rect 282 257 283 258
rect 281 257 282 258
rect 280 257 281 258
rect 279 257 280 258
rect 278 257 279 258
rect 277 257 278 258
rect 276 257 277 258
rect 275 257 276 258
rect 274 257 275 258
rect 273 257 274 258
rect 272 257 273 258
rect 271 257 272 258
rect 270 257 271 258
rect 269 257 270 258
rect 268 257 269 258
rect 267 257 268 258
rect 266 257 267 258
rect 265 257 266 258
rect 264 257 265 258
rect 263 257 264 258
rect 262 257 263 258
rect 261 257 262 258
rect 260 257 261 258
rect 259 257 260 258
rect 258 257 259 258
rect 257 257 258 258
rect 256 257 257 258
rect 255 257 256 258
rect 254 257 255 258
rect 253 257 254 258
rect 252 257 253 258
rect 251 257 252 258
rect 250 257 251 258
rect 249 257 250 258
rect 248 257 249 258
rect 247 257 248 258
rect 246 257 247 258
rect 245 257 246 258
rect 244 257 245 258
rect 243 257 244 258
rect 242 257 243 258
rect 241 257 242 258
rect 240 257 241 258
rect 239 257 240 258
rect 238 257 239 258
rect 237 257 238 258
rect 236 257 237 258
rect 235 257 236 258
rect 234 257 235 258
rect 233 257 234 258
rect 232 257 233 258
rect 168 257 169 258
rect 167 257 168 258
rect 166 257 167 258
rect 165 257 166 258
rect 164 257 165 258
rect 163 257 164 258
rect 162 257 163 258
rect 161 257 162 258
rect 160 257 161 258
rect 159 257 160 258
rect 158 257 159 258
rect 157 257 158 258
rect 156 257 157 258
rect 155 257 156 258
rect 154 257 155 258
rect 153 257 154 258
rect 152 257 153 258
rect 151 257 152 258
rect 150 257 151 258
rect 149 257 150 258
rect 148 257 149 258
rect 147 257 148 258
rect 146 257 147 258
rect 145 257 146 258
rect 144 257 145 258
rect 143 257 144 258
rect 142 257 143 258
rect 141 257 142 258
rect 140 257 141 258
rect 139 257 140 258
rect 138 257 139 258
rect 137 257 138 258
rect 136 257 137 258
rect 135 257 136 258
rect 134 257 135 258
rect 133 257 134 258
rect 132 257 133 258
rect 131 257 132 258
rect 130 257 131 258
rect 129 257 130 258
rect 128 257 129 258
rect 127 257 128 258
rect 126 257 127 258
rect 125 257 126 258
rect 124 257 125 258
rect 111 257 112 258
rect 110 257 111 258
rect 109 257 110 258
rect 108 257 109 258
rect 107 257 108 258
rect 106 257 107 258
rect 105 257 106 258
rect 104 257 105 258
rect 103 257 104 258
rect 102 257 103 258
rect 101 257 102 258
rect 100 257 101 258
rect 99 257 100 258
rect 98 257 99 258
rect 97 257 98 258
rect 96 257 97 258
rect 95 257 96 258
rect 94 257 95 258
rect 93 257 94 258
rect 92 257 93 258
rect 91 257 92 258
rect 90 257 91 258
rect 89 257 90 258
rect 88 257 89 258
rect 87 257 88 258
rect 86 257 87 258
rect 85 257 86 258
rect 84 257 85 258
rect 83 257 84 258
rect 82 257 83 258
rect 81 257 82 258
rect 80 257 81 258
rect 79 257 80 258
rect 78 257 79 258
rect 77 257 78 258
rect 76 257 77 258
rect 75 257 76 258
rect 74 257 75 258
rect 73 257 74 258
rect 72 257 73 258
rect 71 257 72 258
rect 70 257 71 258
rect 69 257 70 258
rect 68 257 69 258
rect 67 257 68 258
rect 66 257 67 258
rect 65 257 66 258
rect 56 257 57 258
rect 55 257 56 258
rect 54 257 55 258
rect 53 257 54 258
rect 52 257 53 258
rect 51 257 52 258
rect 50 257 51 258
rect 49 257 50 258
rect 48 257 49 258
rect 47 257 48 258
rect 46 257 47 258
rect 45 257 46 258
rect 44 257 45 258
rect 43 257 44 258
rect 42 257 43 258
rect 41 257 42 258
rect 40 257 41 258
rect 39 257 40 258
rect 38 257 39 258
rect 37 257 38 258
rect 36 257 37 258
rect 35 257 36 258
rect 24 257 25 258
rect 23 257 24 258
rect 22 257 23 258
rect 21 257 22 258
rect 20 257 21 258
rect 19 257 20 258
rect 18 257 19 258
rect 17 257 18 258
rect 16 257 17 258
rect 15 257 16 258
rect 14 257 15 258
rect 13 257 14 258
rect 12 257 13 258
rect 11 257 12 258
rect 10 257 11 258
rect 9 257 10 258
rect 8 257 9 258
rect 7 257 8 258
rect 6 257 7 258
rect 5 257 6 258
rect 480 258 481 259
rect 479 258 480 259
rect 478 258 479 259
rect 477 258 478 259
rect 476 258 477 259
rect 475 258 476 259
rect 474 258 475 259
rect 473 258 474 259
rect 466 258 467 259
rect 465 258 466 259
rect 464 258 465 259
rect 463 258 464 259
rect 462 258 463 259
rect 310 258 311 259
rect 309 258 310 259
rect 308 258 309 259
rect 307 258 308 259
rect 306 258 307 259
rect 305 258 306 259
rect 304 258 305 259
rect 303 258 304 259
rect 302 258 303 259
rect 301 258 302 259
rect 300 258 301 259
rect 299 258 300 259
rect 298 258 299 259
rect 297 258 298 259
rect 296 258 297 259
rect 295 258 296 259
rect 294 258 295 259
rect 293 258 294 259
rect 292 258 293 259
rect 291 258 292 259
rect 290 258 291 259
rect 289 258 290 259
rect 288 258 289 259
rect 287 258 288 259
rect 286 258 287 259
rect 285 258 286 259
rect 284 258 285 259
rect 283 258 284 259
rect 282 258 283 259
rect 281 258 282 259
rect 280 258 281 259
rect 279 258 280 259
rect 278 258 279 259
rect 277 258 278 259
rect 276 258 277 259
rect 275 258 276 259
rect 274 258 275 259
rect 273 258 274 259
rect 272 258 273 259
rect 271 258 272 259
rect 270 258 271 259
rect 269 258 270 259
rect 268 258 269 259
rect 267 258 268 259
rect 266 258 267 259
rect 265 258 266 259
rect 264 258 265 259
rect 263 258 264 259
rect 262 258 263 259
rect 261 258 262 259
rect 260 258 261 259
rect 259 258 260 259
rect 258 258 259 259
rect 257 258 258 259
rect 256 258 257 259
rect 255 258 256 259
rect 254 258 255 259
rect 253 258 254 259
rect 252 258 253 259
rect 251 258 252 259
rect 250 258 251 259
rect 249 258 250 259
rect 248 258 249 259
rect 247 258 248 259
rect 246 258 247 259
rect 245 258 246 259
rect 244 258 245 259
rect 243 258 244 259
rect 242 258 243 259
rect 241 258 242 259
rect 240 258 241 259
rect 239 258 240 259
rect 238 258 239 259
rect 237 258 238 259
rect 236 258 237 259
rect 235 258 236 259
rect 234 258 235 259
rect 233 258 234 259
rect 232 258 233 259
rect 170 258 171 259
rect 169 258 170 259
rect 168 258 169 259
rect 167 258 168 259
rect 166 258 167 259
rect 165 258 166 259
rect 164 258 165 259
rect 163 258 164 259
rect 162 258 163 259
rect 161 258 162 259
rect 160 258 161 259
rect 159 258 160 259
rect 158 258 159 259
rect 157 258 158 259
rect 156 258 157 259
rect 155 258 156 259
rect 154 258 155 259
rect 153 258 154 259
rect 152 258 153 259
rect 151 258 152 259
rect 150 258 151 259
rect 149 258 150 259
rect 148 258 149 259
rect 147 258 148 259
rect 146 258 147 259
rect 145 258 146 259
rect 144 258 145 259
rect 143 258 144 259
rect 142 258 143 259
rect 141 258 142 259
rect 140 258 141 259
rect 139 258 140 259
rect 138 258 139 259
rect 137 258 138 259
rect 136 258 137 259
rect 135 258 136 259
rect 134 258 135 259
rect 133 258 134 259
rect 132 258 133 259
rect 131 258 132 259
rect 130 258 131 259
rect 129 258 130 259
rect 128 258 129 259
rect 127 258 128 259
rect 126 258 127 259
rect 125 258 126 259
rect 124 258 125 259
rect 111 258 112 259
rect 110 258 111 259
rect 109 258 110 259
rect 108 258 109 259
rect 107 258 108 259
rect 106 258 107 259
rect 105 258 106 259
rect 104 258 105 259
rect 103 258 104 259
rect 102 258 103 259
rect 101 258 102 259
rect 100 258 101 259
rect 99 258 100 259
rect 98 258 99 259
rect 97 258 98 259
rect 96 258 97 259
rect 95 258 96 259
rect 94 258 95 259
rect 93 258 94 259
rect 92 258 93 259
rect 91 258 92 259
rect 90 258 91 259
rect 89 258 90 259
rect 88 258 89 259
rect 87 258 88 259
rect 86 258 87 259
rect 85 258 86 259
rect 84 258 85 259
rect 83 258 84 259
rect 82 258 83 259
rect 81 258 82 259
rect 80 258 81 259
rect 79 258 80 259
rect 78 258 79 259
rect 77 258 78 259
rect 76 258 77 259
rect 75 258 76 259
rect 74 258 75 259
rect 73 258 74 259
rect 72 258 73 259
rect 71 258 72 259
rect 70 258 71 259
rect 69 258 70 259
rect 68 258 69 259
rect 67 258 68 259
rect 56 258 57 259
rect 55 258 56 259
rect 54 258 55 259
rect 53 258 54 259
rect 52 258 53 259
rect 51 258 52 259
rect 50 258 51 259
rect 49 258 50 259
rect 48 258 49 259
rect 47 258 48 259
rect 46 258 47 259
rect 45 258 46 259
rect 44 258 45 259
rect 43 258 44 259
rect 42 258 43 259
rect 41 258 42 259
rect 40 258 41 259
rect 39 258 40 259
rect 38 258 39 259
rect 37 258 38 259
rect 36 258 37 259
rect 35 258 36 259
rect 24 258 25 259
rect 23 258 24 259
rect 22 258 23 259
rect 21 258 22 259
rect 20 258 21 259
rect 19 258 20 259
rect 18 258 19 259
rect 17 258 18 259
rect 16 258 17 259
rect 15 258 16 259
rect 14 258 15 259
rect 13 258 14 259
rect 12 258 13 259
rect 11 258 12 259
rect 10 258 11 259
rect 9 258 10 259
rect 8 258 9 259
rect 7 258 8 259
rect 6 258 7 259
rect 5 258 6 259
rect 479 259 480 260
rect 478 259 479 260
rect 477 259 478 260
rect 476 259 477 260
rect 475 259 476 260
rect 474 259 475 260
rect 309 259 310 260
rect 308 259 309 260
rect 307 259 308 260
rect 306 259 307 260
rect 305 259 306 260
rect 304 259 305 260
rect 303 259 304 260
rect 302 259 303 260
rect 301 259 302 260
rect 300 259 301 260
rect 299 259 300 260
rect 298 259 299 260
rect 297 259 298 260
rect 296 259 297 260
rect 295 259 296 260
rect 294 259 295 260
rect 293 259 294 260
rect 292 259 293 260
rect 291 259 292 260
rect 290 259 291 260
rect 289 259 290 260
rect 288 259 289 260
rect 287 259 288 260
rect 286 259 287 260
rect 285 259 286 260
rect 284 259 285 260
rect 283 259 284 260
rect 282 259 283 260
rect 281 259 282 260
rect 280 259 281 260
rect 279 259 280 260
rect 278 259 279 260
rect 277 259 278 260
rect 276 259 277 260
rect 275 259 276 260
rect 274 259 275 260
rect 273 259 274 260
rect 272 259 273 260
rect 271 259 272 260
rect 270 259 271 260
rect 269 259 270 260
rect 268 259 269 260
rect 267 259 268 260
rect 266 259 267 260
rect 265 259 266 260
rect 264 259 265 260
rect 263 259 264 260
rect 262 259 263 260
rect 261 259 262 260
rect 260 259 261 260
rect 259 259 260 260
rect 258 259 259 260
rect 257 259 258 260
rect 256 259 257 260
rect 255 259 256 260
rect 254 259 255 260
rect 253 259 254 260
rect 252 259 253 260
rect 251 259 252 260
rect 250 259 251 260
rect 249 259 250 260
rect 248 259 249 260
rect 247 259 248 260
rect 246 259 247 260
rect 245 259 246 260
rect 244 259 245 260
rect 243 259 244 260
rect 242 259 243 260
rect 241 259 242 260
rect 240 259 241 260
rect 239 259 240 260
rect 238 259 239 260
rect 237 259 238 260
rect 236 259 237 260
rect 235 259 236 260
rect 234 259 235 260
rect 233 259 234 260
rect 232 259 233 260
rect 231 259 232 260
rect 172 259 173 260
rect 171 259 172 260
rect 170 259 171 260
rect 169 259 170 260
rect 168 259 169 260
rect 167 259 168 260
rect 166 259 167 260
rect 165 259 166 260
rect 164 259 165 260
rect 163 259 164 260
rect 162 259 163 260
rect 161 259 162 260
rect 160 259 161 260
rect 159 259 160 260
rect 158 259 159 260
rect 157 259 158 260
rect 156 259 157 260
rect 155 259 156 260
rect 154 259 155 260
rect 153 259 154 260
rect 152 259 153 260
rect 151 259 152 260
rect 150 259 151 260
rect 149 259 150 260
rect 148 259 149 260
rect 147 259 148 260
rect 146 259 147 260
rect 145 259 146 260
rect 144 259 145 260
rect 143 259 144 260
rect 142 259 143 260
rect 141 259 142 260
rect 140 259 141 260
rect 139 259 140 260
rect 138 259 139 260
rect 137 259 138 260
rect 136 259 137 260
rect 135 259 136 260
rect 134 259 135 260
rect 133 259 134 260
rect 132 259 133 260
rect 131 259 132 260
rect 130 259 131 260
rect 129 259 130 260
rect 128 259 129 260
rect 127 259 128 260
rect 126 259 127 260
rect 125 259 126 260
rect 124 259 125 260
rect 111 259 112 260
rect 110 259 111 260
rect 109 259 110 260
rect 108 259 109 260
rect 107 259 108 260
rect 106 259 107 260
rect 105 259 106 260
rect 104 259 105 260
rect 103 259 104 260
rect 102 259 103 260
rect 101 259 102 260
rect 100 259 101 260
rect 99 259 100 260
rect 98 259 99 260
rect 97 259 98 260
rect 96 259 97 260
rect 95 259 96 260
rect 94 259 95 260
rect 93 259 94 260
rect 92 259 93 260
rect 91 259 92 260
rect 90 259 91 260
rect 89 259 90 260
rect 88 259 89 260
rect 87 259 88 260
rect 86 259 87 260
rect 85 259 86 260
rect 84 259 85 260
rect 83 259 84 260
rect 82 259 83 260
rect 81 259 82 260
rect 80 259 81 260
rect 79 259 80 260
rect 78 259 79 260
rect 77 259 78 260
rect 76 259 77 260
rect 75 259 76 260
rect 74 259 75 260
rect 73 259 74 260
rect 72 259 73 260
rect 71 259 72 260
rect 70 259 71 260
rect 69 259 70 260
rect 57 259 58 260
rect 56 259 57 260
rect 55 259 56 260
rect 54 259 55 260
rect 53 259 54 260
rect 52 259 53 260
rect 51 259 52 260
rect 50 259 51 260
rect 49 259 50 260
rect 48 259 49 260
rect 47 259 48 260
rect 46 259 47 260
rect 45 259 46 260
rect 44 259 45 260
rect 43 259 44 260
rect 42 259 43 260
rect 41 259 42 260
rect 40 259 41 260
rect 39 259 40 260
rect 38 259 39 260
rect 37 259 38 260
rect 36 259 37 260
rect 35 259 36 260
rect 24 259 25 260
rect 23 259 24 260
rect 22 259 23 260
rect 21 259 22 260
rect 20 259 21 260
rect 19 259 20 260
rect 18 259 19 260
rect 17 259 18 260
rect 16 259 17 260
rect 15 259 16 260
rect 14 259 15 260
rect 13 259 14 260
rect 12 259 13 260
rect 11 259 12 260
rect 10 259 11 260
rect 9 259 10 260
rect 8 259 9 260
rect 7 259 8 260
rect 6 259 7 260
rect 5 259 6 260
rect 308 260 309 261
rect 307 260 308 261
rect 306 260 307 261
rect 305 260 306 261
rect 304 260 305 261
rect 303 260 304 261
rect 302 260 303 261
rect 301 260 302 261
rect 300 260 301 261
rect 299 260 300 261
rect 298 260 299 261
rect 297 260 298 261
rect 296 260 297 261
rect 295 260 296 261
rect 294 260 295 261
rect 293 260 294 261
rect 292 260 293 261
rect 291 260 292 261
rect 290 260 291 261
rect 289 260 290 261
rect 288 260 289 261
rect 287 260 288 261
rect 286 260 287 261
rect 285 260 286 261
rect 284 260 285 261
rect 283 260 284 261
rect 282 260 283 261
rect 281 260 282 261
rect 280 260 281 261
rect 279 260 280 261
rect 278 260 279 261
rect 277 260 278 261
rect 276 260 277 261
rect 275 260 276 261
rect 274 260 275 261
rect 273 260 274 261
rect 272 260 273 261
rect 271 260 272 261
rect 270 260 271 261
rect 269 260 270 261
rect 268 260 269 261
rect 267 260 268 261
rect 266 260 267 261
rect 265 260 266 261
rect 264 260 265 261
rect 263 260 264 261
rect 262 260 263 261
rect 261 260 262 261
rect 260 260 261 261
rect 259 260 260 261
rect 258 260 259 261
rect 257 260 258 261
rect 256 260 257 261
rect 255 260 256 261
rect 254 260 255 261
rect 253 260 254 261
rect 252 260 253 261
rect 251 260 252 261
rect 250 260 251 261
rect 249 260 250 261
rect 248 260 249 261
rect 247 260 248 261
rect 246 260 247 261
rect 245 260 246 261
rect 244 260 245 261
rect 243 260 244 261
rect 242 260 243 261
rect 241 260 242 261
rect 240 260 241 261
rect 239 260 240 261
rect 238 260 239 261
rect 237 260 238 261
rect 236 260 237 261
rect 235 260 236 261
rect 234 260 235 261
rect 233 260 234 261
rect 232 260 233 261
rect 231 260 232 261
rect 175 260 176 261
rect 174 260 175 261
rect 173 260 174 261
rect 172 260 173 261
rect 171 260 172 261
rect 170 260 171 261
rect 169 260 170 261
rect 168 260 169 261
rect 167 260 168 261
rect 166 260 167 261
rect 165 260 166 261
rect 164 260 165 261
rect 163 260 164 261
rect 162 260 163 261
rect 161 260 162 261
rect 160 260 161 261
rect 159 260 160 261
rect 158 260 159 261
rect 157 260 158 261
rect 156 260 157 261
rect 155 260 156 261
rect 154 260 155 261
rect 153 260 154 261
rect 152 260 153 261
rect 151 260 152 261
rect 150 260 151 261
rect 149 260 150 261
rect 148 260 149 261
rect 147 260 148 261
rect 146 260 147 261
rect 145 260 146 261
rect 144 260 145 261
rect 143 260 144 261
rect 142 260 143 261
rect 141 260 142 261
rect 140 260 141 261
rect 139 260 140 261
rect 138 260 139 261
rect 137 260 138 261
rect 136 260 137 261
rect 135 260 136 261
rect 134 260 135 261
rect 133 260 134 261
rect 132 260 133 261
rect 131 260 132 261
rect 130 260 131 261
rect 129 260 130 261
rect 128 260 129 261
rect 127 260 128 261
rect 126 260 127 261
rect 125 260 126 261
rect 124 260 125 261
rect 111 260 112 261
rect 110 260 111 261
rect 109 260 110 261
rect 108 260 109 261
rect 107 260 108 261
rect 106 260 107 261
rect 105 260 106 261
rect 104 260 105 261
rect 103 260 104 261
rect 102 260 103 261
rect 101 260 102 261
rect 100 260 101 261
rect 99 260 100 261
rect 98 260 99 261
rect 97 260 98 261
rect 96 260 97 261
rect 95 260 96 261
rect 94 260 95 261
rect 93 260 94 261
rect 92 260 93 261
rect 91 260 92 261
rect 90 260 91 261
rect 89 260 90 261
rect 88 260 89 261
rect 87 260 88 261
rect 86 260 87 261
rect 85 260 86 261
rect 84 260 85 261
rect 83 260 84 261
rect 82 260 83 261
rect 81 260 82 261
rect 80 260 81 261
rect 79 260 80 261
rect 78 260 79 261
rect 77 260 78 261
rect 76 260 77 261
rect 75 260 76 261
rect 74 260 75 261
rect 73 260 74 261
rect 72 260 73 261
rect 71 260 72 261
rect 70 260 71 261
rect 57 260 58 261
rect 56 260 57 261
rect 55 260 56 261
rect 54 260 55 261
rect 53 260 54 261
rect 52 260 53 261
rect 51 260 52 261
rect 50 260 51 261
rect 49 260 50 261
rect 48 260 49 261
rect 47 260 48 261
rect 46 260 47 261
rect 45 260 46 261
rect 44 260 45 261
rect 43 260 44 261
rect 42 260 43 261
rect 41 260 42 261
rect 40 260 41 261
rect 39 260 40 261
rect 38 260 39 261
rect 37 260 38 261
rect 36 260 37 261
rect 24 260 25 261
rect 23 260 24 261
rect 22 260 23 261
rect 21 260 22 261
rect 20 260 21 261
rect 19 260 20 261
rect 18 260 19 261
rect 17 260 18 261
rect 16 260 17 261
rect 15 260 16 261
rect 14 260 15 261
rect 13 260 14 261
rect 12 260 13 261
rect 11 260 12 261
rect 10 260 11 261
rect 9 260 10 261
rect 8 260 9 261
rect 7 260 8 261
rect 6 260 7 261
rect 5 260 6 261
rect 307 261 308 262
rect 306 261 307 262
rect 305 261 306 262
rect 304 261 305 262
rect 303 261 304 262
rect 302 261 303 262
rect 301 261 302 262
rect 300 261 301 262
rect 299 261 300 262
rect 298 261 299 262
rect 297 261 298 262
rect 296 261 297 262
rect 295 261 296 262
rect 294 261 295 262
rect 293 261 294 262
rect 292 261 293 262
rect 291 261 292 262
rect 290 261 291 262
rect 289 261 290 262
rect 288 261 289 262
rect 287 261 288 262
rect 286 261 287 262
rect 285 261 286 262
rect 284 261 285 262
rect 283 261 284 262
rect 282 261 283 262
rect 281 261 282 262
rect 280 261 281 262
rect 279 261 280 262
rect 278 261 279 262
rect 277 261 278 262
rect 276 261 277 262
rect 275 261 276 262
rect 274 261 275 262
rect 273 261 274 262
rect 272 261 273 262
rect 271 261 272 262
rect 270 261 271 262
rect 269 261 270 262
rect 268 261 269 262
rect 267 261 268 262
rect 266 261 267 262
rect 265 261 266 262
rect 264 261 265 262
rect 263 261 264 262
rect 262 261 263 262
rect 261 261 262 262
rect 260 261 261 262
rect 259 261 260 262
rect 258 261 259 262
rect 257 261 258 262
rect 256 261 257 262
rect 255 261 256 262
rect 254 261 255 262
rect 253 261 254 262
rect 252 261 253 262
rect 251 261 252 262
rect 250 261 251 262
rect 249 261 250 262
rect 248 261 249 262
rect 247 261 248 262
rect 246 261 247 262
rect 245 261 246 262
rect 244 261 245 262
rect 243 261 244 262
rect 242 261 243 262
rect 241 261 242 262
rect 240 261 241 262
rect 239 261 240 262
rect 238 261 239 262
rect 237 261 238 262
rect 236 261 237 262
rect 235 261 236 262
rect 234 261 235 262
rect 233 261 234 262
rect 232 261 233 262
rect 231 261 232 262
rect 179 261 180 262
rect 178 261 179 262
rect 177 261 178 262
rect 176 261 177 262
rect 175 261 176 262
rect 174 261 175 262
rect 173 261 174 262
rect 172 261 173 262
rect 171 261 172 262
rect 170 261 171 262
rect 169 261 170 262
rect 168 261 169 262
rect 167 261 168 262
rect 166 261 167 262
rect 165 261 166 262
rect 164 261 165 262
rect 163 261 164 262
rect 162 261 163 262
rect 161 261 162 262
rect 160 261 161 262
rect 159 261 160 262
rect 158 261 159 262
rect 157 261 158 262
rect 156 261 157 262
rect 155 261 156 262
rect 154 261 155 262
rect 153 261 154 262
rect 152 261 153 262
rect 151 261 152 262
rect 150 261 151 262
rect 149 261 150 262
rect 148 261 149 262
rect 147 261 148 262
rect 146 261 147 262
rect 145 261 146 262
rect 144 261 145 262
rect 143 261 144 262
rect 142 261 143 262
rect 141 261 142 262
rect 140 261 141 262
rect 139 261 140 262
rect 138 261 139 262
rect 137 261 138 262
rect 136 261 137 262
rect 135 261 136 262
rect 134 261 135 262
rect 133 261 134 262
rect 132 261 133 262
rect 131 261 132 262
rect 130 261 131 262
rect 129 261 130 262
rect 128 261 129 262
rect 127 261 128 262
rect 126 261 127 262
rect 125 261 126 262
rect 124 261 125 262
rect 112 261 113 262
rect 111 261 112 262
rect 110 261 111 262
rect 109 261 110 262
rect 108 261 109 262
rect 107 261 108 262
rect 106 261 107 262
rect 105 261 106 262
rect 104 261 105 262
rect 103 261 104 262
rect 102 261 103 262
rect 101 261 102 262
rect 100 261 101 262
rect 99 261 100 262
rect 98 261 99 262
rect 97 261 98 262
rect 96 261 97 262
rect 95 261 96 262
rect 94 261 95 262
rect 93 261 94 262
rect 92 261 93 262
rect 91 261 92 262
rect 90 261 91 262
rect 89 261 90 262
rect 88 261 89 262
rect 87 261 88 262
rect 86 261 87 262
rect 85 261 86 262
rect 84 261 85 262
rect 83 261 84 262
rect 82 261 83 262
rect 81 261 82 262
rect 80 261 81 262
rect 79 261 80 262
rect 78 261 79 262
rect 77 261 78 262
rect 76 261 77 262
rect 75 261 76 262
rect 74 261 75 262
rect 73 261 74 262
rect 72 261 73 262
rect 71 261 72 262
rect 57 261 58 262
rect 56 261 57 262
rect 55 261 56 262
rect 54 261 55 262
rect 53 261 54 262
rect 52 261 53 262
rect 51 261 52 262
rect 50 261 51 262
rect 49 261 50 262
rect 48 261 49 262
rect 47 261 48 262
rect 46 261 47 262
rect 45 261 46 262
rect 44 261 45 262
rect 43 261 44 262
rect 42 261 43 262
rect 41 261 42 262
rect 40 261 41 262
rect 39 261 40 262
rect 38 261 39 262
rect 37 261 38 262
rect 36 261 37 262
rect 25 261 26 262
rect 24 261 25 262
rect 23 261 24 262
rect 22 261 23 262
rect 21 261 22 262
rect 20 261 21 262
rect 19 261 20 262
rect 18 261 19 262
rect 17 261 18 262
rect 16 261 17 262
rect 15 261 16 262
rect 14 261 15 262
rect 13 261 14 262
rect 12 261 13 262
rect 11 261 12 262
rect 10 261 11 262
rect 9 261 10 262
rect 8 261 9 262
rect 7 261 8 262
rect 6 261 7 262
rect 5 261 6 262
rect 306 262 307 263
rect 305 262 306 263
rect 304 262 305 263
rect 303 262 304 263
rect 302 262 303 263
rect 301 262 302 263
rect 300 262 301 263
rect 299 262 300 263
rect 298 262 299 263
rect 297 262 298 263
rect 296 262 297 263
rect 295 262 296 263
rect 294 262 295 263
rect 293 262 294 263
rect 292 262 293 263
rect 291 262 292 263
rect 290 262 291 263
rect 289 262 290 263
rect 288 262 289 263
rect 287 262 288 263
rect 286 262 287 263
rect 285 262 286 263
rect 284 262 285 263
rect 283 262 284 263
rect 282 262 283 263
rect 281 262 282 263
rect 280 262 281 263
rect 279 262 280 263
rect 278 262 279 263
rect 277 262 278 263
rect 276 262 277 263
rect 275 262 276 263
rect 274 262 275 263
rect 273 262 274 263
rect 272 262 273 263
rect 271 262 272 263
rect 270 262 271 263
rect 269 262 270 263
rect 268 262 269 263
rect 267 262 268 263
rect 266 262 267 263
rect 265 262 266 263
rect 264 262 265 263
rect 263 262 264 263
rect 262 262 263 263
rect 261 262 262 263
rect 260 262 261 263
rect 259 262 260 263
rect 258 262 259 263
rect 257 262 258 263
rect 256 262 257 263
rect 255 262 256 263
rect 254 262 255 263
rect 253 262 254 263
rect 252 262 253 263
rect 251 262 252 263
rect 250 262 251 263
rect 249 262 250 263
rect 248 262 249 263
rect 247 262 248 263
rect 246 262 247 263
rect 245 262 246 263
rect 244 262 245 263
rect 243 262 244 263
rect 242 262 243 263
rect 241 262 242 263
rect 240 262 241 263
rect 239 262 240 263
rect 238 262 239 263
rect 237 262 238 263
rect 236 262 237 263
rect 235 262 236 263
rect 234 262 235 263
rect 233 262 234 263
rect 232 262 233 263
rect 231 262 232 263
rect 230 262 231 263
rect 183 262 184 263
rect 182 262 183 263
rect 181 262 182 263
rect 180 262 181 263
rect 179 262 180 263
rect 178 262 179 263
rect 177 262 178 263
rect 176 262 177 263
rect 175 262 176 263
rect 174 262 175 263
rect 173 262 174 263
rect 172 262 173 263
rect 171 262 172 263
rect 170 262 171 263
rect 169 262 170 263
rect 168 262 169 263
rect 167 262 168 263
rect 166 262 167 263
rect 165 262 166 263
rect 164 262 165 263
rect 163 262 164 263
rect 162 262 163 263
rect 161 262 162 263
rect 160 262 161 263
rect 159 262 160 263
rect 158 262 159 263
rect 157 262 158 263
rect 156 262 157 263
rect 155 262 156 263
rect 154 262 155 263
rect 153 262 154 263
rect 152 262 153 263
rect 151 262 152 263
rect 150 262 151 263
rect 149 262 150 263
rect 148 262 149 263
rect 147 262 148 263
rect 146 262 147 263
rect 145 262 146 263
rect 144 262 145 263
rect 143 262 144 263
rect 142 262 143 263
rect 141 262 142 263
rect 140 262 141 263
rect 139 262 140 263
rect 138 262 139 263
rect 137 262 138 263
rect 136 262 137 263
rect 135 262 136 263
rect 134 262 135 263
rect 133 262 134 263
rect 132 262 133 263
rect 131 262 132 263
rect 130 262 131 263
rect 129 262 130 263
rect 128 262 129 263
rect 127 262 128 263
rect 126 262 127 263
rect 125 262 126 263
rect 124 262 125 263
rect 112 262 113 263
rect 111 262 112 263
rect 110 262 111 263
rect 109 262 110 263
rect 108 262 109 263
rect 107 262 108 263
rect 106 262 107 263
rect 105 262 106 263
rect 104 262 105 263
rect 103 262 104 263
rect 102 262 103 263
rect 101 262 102 263
rect 100 262 101 263
rect 99 262 100 263
rect 98 262 99 263
rect 97 262 98 263
rect 96 262 97 263
rect 95 262 96 263
rect 94 262 95 263
rect 93 262 94 263
rect 92 262 93 263
rect 91 262 92 263
rect 90 262 91 263
rect 89 262 90 263
rect 88 262 89 263
rect 87 262 88 263
rect 86 262 87 263
rect 85 262 86 263
rect 84 262 85 263
rect 83 262 84 263
rect 82 262 83 263
rect 81 262 82 263
rect 80 262 81 263
rect 79 262 80 263
rect 78 262 79 263
rect 77 262 78 263
rect 76 262 77 263
rect 75 262 76 263
rect 74 262 75 263
rect 73 262 74 263
rect 72 262 73 263
rect 57 262 58 263
rect 56 262 57 263
rect 55 262 56 263
rect 54 262 55 263
rect 53 262 54 263
rect 52 262 53 263
rect 51 262 52 263
rect 50 262 51 263
rect 49 262 50 263
rect 48 262 49 263
rect 47 262 48 263
rect 46 262 47 263
rect 45 262 46 263
rect 44 262 45 263
rect 43 262 44 263
rect 42 262 43 263
rect 41 262 42 263
rect 40 262 41 263
rect 39 262 40 263
rect 38 262 39 263
rect 37 262 38 263
rect 36 262 37 263
rect 25 262 26 263
rect 24 262 25 263
rect 23 262 24 263
rect 22 262 23 263
rect 21 262 22 263
rect 20 262 21 263
rect 19 262 20 263
rect 18 262 19 263
rect 17 262 18 263
rect 16 262 17 263
rect 15 262 16 263
rect 14 262 15 263
rect 13 262 14 263
rect 12 262 13 263
rect 11 262 12 263
rect 10 262 11 263
rect 9 262 10 263
rect 8 262 9 263
rect 7 262 8 263
rect 6 262 7 263
rect 5 262 6 263
rect 305 263 306 264
rect 304 263 305 264
rect 303 263 304 264
rect 302 263 303 264
rect 301 263 302 264
rect 300 263 301 264
rect 299 263 300 264
rect 298 263 299 264
rect 297 263 298 264
rect 296 263 297 264
rect 295 263 296 264
rect 294 263 295 264
rect 293 263 294 264
rect 292 263 293 264
rect 291 263 292 264
rect 290 263 291 264
rect 289 263 290 264
rect 288 263 289 264
rect 287 263 288 264
rect 286 263 287 264
rect 285 263 286 264
rect 284 263 285 264
rect 283 263 284 264
rect 282 263 283 264
rect 281 263 282 264
rect 280 263 281 264
rect 279 263 280 264
rect 278 263 279 264
rect 277 263 278 264
rect 276 263 277 264
rect 275 263 276 264
rect 274 263 275 264
rect 273 263 274 264
rect 272 263 273 264
rect 271 263 272 264
rect 270 263 271 264
rect 269 263 270 264
rect 268 263 269 264
rect 267 263 268 264
rect 266 263 267 264
rect 265 263 266 264
rect 264 263 265 264
rect 263 263 264 264
rect 262 263 263 264
rect 261 263 262 264
rect 260 263 261 264
rect 259 263 260 264
rect 258 263 259 264
rect 257 263 258 264
rect 256 263 257 264
rect 255 263 256 264
rect 254 263 255 264
rect 253 263 254 264
rect 252 263 253 264
rect 251 263 252 264
rect 250 263 251 264
rect 249 263 250 264
rect 248 263 249 264
rect 247 263 248 264
rect 246 263 247 264
rect 245 263 246 264
rect 244 263 245 264
rect 243 263 244 264
rect 242 263 243 264
rect 241 263 242 264
rect 240 263 241 264
rect 239 263 240 264
rect 238 263 239 264
rect 237 263 238 264
rect 236 263 237 264
rect 235 263 236 264
rect 234 263 235 264
rect 233 263 234 264
rect 232 263 233 264
rect 231 263 232 264
rect 230 263 231 264
rect 187 263 188 264
rect 186 263 187 264
rect 185 263 186 264
rect 184 263 185 264
rect 183 263 184 264
rect 182 263 183 264
rect 181 263 182 264
rect 180 263 181 264
rect 179 263 180 264
rect 178 263 179 264
rect 177 263 178 264
rect 176 263 177 264
rect 175 263 176 264
rect 174 263 175 264
rect 173 263 174 264
rect 172 263 173 264
rect 171 263 172 264
rect 170 263 171 264
rect 169 263 170 264
rect 168 263 169 264
rect 167 263 168 264
rect 166 263 167 264
rect 165 263 166 264
rect 164 263 165 264
rect 163 263 164 264
rect 162 263 163 264
rect 161 263 162 264
rect 160 263 161 264
rect 159 263 160 264
rect 158 263 159 264
rect 157 263 158 264
rect 156 263 157 264
rect 155 263 156 264
rect 154 263 155 264
rect 153 263 154 264
rect 152 263 153 264
rect 151 263 152 264
rect 150 263 151 264
rect 149 263 150 264
rect 148 263 149 264
rect 147 263 148 264
rect 146 263 147 264
rect 145 263 146 264
rect 144 263 145 264
rect 143 263 144 264
rect 142 263 143 264
rect 141 263 142 264
rect 140 263 141 264
rect 139 263 140 264
rect 138 263 139 264
rect 137 263 138 264
rect 136 263 137 264
rect 135 263 136 264
rect 134 263 135 264
rect 133 263 134 264
rect 132 263 133 264
rect 131 263 132 264
rect 130 263 131 264
rect 129 263 130 264
rect 128 263 129 264
rect 127 263 128 264
rect 126 263 127 264
rect 125 263 126 264
rect 112 263 113 264
rect 111 263 112 264
rect 110 263 111 264
rect 109 263 110 264
rect 108 263 109 264
rect 107 263 108 264
rect 106 263 107 264
rect 105 263 106 264
rect 104 263 105 264
rect 103 263 104 264
rect 102 263 103 264
rect 101 263 102 264
rect 100 263 101 264
rect 99 263 100 264
rect 98 263 99 264
rect 97 263 98 264
rect 96 263 97 264
rect 95 263 96 264
rect 94 263 95 264
rect 93 263 94 264
rect 92 263 93 264
rect 91 263 92 264
rect 90 263 91 264
rect 89 263 90 264
rect 88 263 89 264
rect 87 263 88 264
rect 86 263 87 264
rect 85 263 86 264
rect 84 263 85 264
rect 83 263 84 264
rect 82 263 83 264
rect 81 263 82 264
rect 80 263 81 264
rect 79 263 80 264
rect 78 263 79 264
rect 77 263 78 264
rect 76 263 77 264
rect 75 263 76 264
rect 74 263 75 264
rect 73 263 74 264
rect 58 263 59 264
rect 57 263 58 264
rect 56 263 57 264
rect 55 263 56 264
rect 54 263 55 264
rect 53 263 54 264
rect 52 263 53 264
rect 51 263 52 264
rect 50 263 51 264
rect 49 263 50 264
rect 48 263 49 264
rect 47 263 48 264
rect 46 263 47 264
rect 45 263 46 264
rect 44 263 45 264
rect 43 263 44 264
rect 42 263 43 264
rect 41 263 42 264
rect 40 263 41 264
rect 39 263 40 264
rect 38 263 39 264
rect 37 263 38 264
rect 25 263 26 264
rect 24 263 25 264
rect 23 263 24 264
rect 22 263 23 264
rect 21 263 22 264
rect 20 263 21 264
rect 19 263 20 264
rect 18 263 19 264
rect 17 263 18 264
rect 16 263 17 264
rect 15 263 16 264
rect 14 263 15 264
rect 13 263 14 264
rect 12 263 13 264
rect 11 263 12 264
rect 10 263 11 264
rect 9 263 10 264
rect 8 263 9 264
rect 7 263 8 264
rect 6 263 7 264
rect 5 263 6 264
rect 304 264 305 265
rect 303 264 304 265
rect 302 264 303 265
rect 301 264 302 265
rect 300 264 301 265
rect 299 264 300 265
rect 298 264 299 265
rect 297 264 298 265
rect 296 264 297 265
rect 295 264 296 265
rect 294 264 295 265
rect 293 264 294 265
rect 292 264 293 265
rect 291 264 292 265
rect 290 264 291 265
rect 289 264 290 265
rect 288 264 289 265
rect 287 264 288 265
rect 286 264 287 265
rect 285 264 286 265
rect 284 264 285 265
rect 283 264 284 265
rect 282 264 283 265
rect 281 264 282 265
rect 280 264 281 265
rect 279 264 280 265
rect 278 264 279 265
rect 277 264 278 265
rect 276 264 277 265
rect 275 264 276 265
rect 274 264 275 265
rect 273 264 274 265
rect 272 264 273 265
rect 271 264 272 265
rect 270 264 271 265
rect 269 264 270 265
rect 268 264 269 265
rect 267 264 268 265
rect 266 264 267 265
rect 265 264 266 265
rect 264 264 265 265
rect 263 264 264 265
rect 262 264 263 265
rect 261 264 262 265
rect 260 264 261 265
rect 259 264 260 265
rect 258 264 259 265
rect 257 264 258 265
rect 256 264 257 265
rect 255 264 256 265
rect 254 264 255 265
rect 253 264 254 265
rect 252 264 253 265
rect 251 264 252 265
rect 250 264 251 265
rect 249 264 250 265
rect 248 264 249 265
rect 247 264 248 265
rect 246 264 247 265
rect 245 264 246 265
rect 244 264 245 265
rect 243 264 244 265
rect 242 264 243 265
rect 241 264 242 265
rect 240 264 241 265
rect 239 264 240 265
rect 238 264 239 265
rect 237 264 238 265
rect 236 264 237 265
rect 235 264 236 265
rect 234 264 235 265
rect 233 264 234 265
rect 232 264 233 265
rect 231 264 232 265
rect 230 264 231 265
rect 209 264 210 265
rect 208 264 209 265
rect 207 264 208 265
rect 206 264 207 265
rect 205 264 206 265
rect 204 264 205 265
rect 194 264 195 265
rect 193 264 194 265
rect 192 264 193 265
rect 191 264 192 265
rect 190 264 191 265
rect 189 264 190 265
rect 188 264 189 265
rect 187 264 188 265
rect 186 264 187 265
rect 185 264 186 265
rect 184 264 185 265
rect 183 264 184 265
rect 182 264 183 265
rect 181 264 182 265
rect 180 264 181 265
rect 179 264 180 265
rect 178 264 179 265
rect 177 264 178 265
rect 176 264 177 265
rect 175 264 176 265
rect 174 264 175 265
rect 173 264 174 265
rect 172 264 173 265
rect 171 264 172 265
rect 170 264 171 265
rect 169 264 170 265
rect 168 264 169 265
rect 167 264 168 265
rect 166 264 167 265
rect 165 264 166 265
rect 164 264 165 265
rect 163 264 164 265
rect 162 264 163 265
rect 161 264 162 265
rect 160 264 161 265
rect 159 264 160 265
rect 158 264 159 265
rect 157 264 158 265
rect 156 264 157 265
rect 155 264 156 265
rect 154 264 155 265
rect 153 264 154 265
rect 152 264 153 265
rect 151 264 152 265
rect 150 264 151 265
rect 149 264 150 265
rect 148 264 149 265
rect 147 264 148 265
rect 146 264 147 265
rect 145 264 146 265
rect 144 264 145 265
rect 143 264 144 265
rect 142 264 143 265
rect 141 264 142 265
rect 140 264 141 265
rect 139 264 140 265
rect 138 264 139 265
rect 137 264 138 265
rect 136 264 137 265
rect 135 264 136 265
rect 134 264 135 265
rect 133 264 134 265
rect 132 264 133 265
rect 131 264 132 265
rect 130 264 131 265
rect 129 264 130 265
rect 128 264 129 265
rect 127 264 128 265
rect 126 264 127 265
rect 125 264 126 265
rect 112 264 113 265
rect 111 264 112 265
rect 110 264 111 265
rect 109 264 110 265
rect 108 264 109 265
rect 107 264 108 265
rect 106 264 107 265
rect 105 264 106 265
rect 104 264 105 265
rect 103 264 104 265
rect 102 264 103 265
rect 101 264 102 265
rect 100 264 101 265
rect 99 264 100 265
rect 98 264 99 265
rect 97 264 98 265
rect 96 264 97 265
rect 95 264 96 265
rect 94 264 95 265
rect 93 264 94 265
rect 92 264 93 265
rect 91 264 92 265
rect 90 264 91 265
rect 89 264 90 265
rect 88 264 89 265
rect 87 264 88 265
rect 86 264 87 265
rect 85 264 86 265
rect 84 264 85 265
rect 83 264 84 265
rect 82 264 83 265
rect 81 264 82 265
rect 80 264 81 265
rect 79 264 80 265
rect 78 264 79 265
rect 77 264 78 265
rect 76 264 77 265
rect 75 264 76 265
rect 74 264 75 265
rect 58 264 59 265
rect 57 264 58 265
rect 56 264 57 265
rect 55 264 56 265
rect 54 264 55 265
rect 53 264 54 265
rect 52 264 53 265
rect 51 264 52 265
rect 50 264 51 265
rect 49 264 50 265
rect 48 264 49 265
rect 47 264 48 265
rect 46 264 47 265
rect 45 264 46 265
rect 44 264 45 265
rect 43 264 44 265
rect 42 264 43 265
rect 41 264 42 265
rect 40 264 41 265
rect 39 264 40 265
rect 38 264 39 265
rect 37 264 38 265
rect 26 264 27 265
rect 25 264 26 265
rect 24 264 25 265
rect 23 264 24 265
rect 22 264 23 265
rect 21 264 22 265
rect 20 264 21 265
rect 19 264 20 265
rect 18 264 19 265
rect 17 264 18 265
rect 16 264 17 265
rect 15 264 16 265
rect 14 264 15 265
rect 13 264 14 265
rect 12 264 13 265
rect 11 264 12 265
rect 10 264 11 265
rect 9 264 10 265
rect 8 264 9 265
rect 7 264 8 265
rect 6 264 7 265
rect 5 264 6 265
rect 304 265 305 266
rect 303 265 304 266
rect 302 265 303 266
rect 301 265 302 266
rect 300 265 301 266
rect 299 265 300 266
rect 298 265 299 266
rect 297 265 298 266
rect 296 265 297 266
rect 295 265 296 266
rect 294 265 295 266
rect 293 265 294 266
rect 292 265 293 266
rect 291 265 292 266
rect 290 265 291 266
rect 289 265 290 266
rect 288 265 289 266
rect 287 265 288 266
rect 286 265 287 266
rect 285 265 286 266
rect 284 265 285 266
rect 283 265 284 266
rect 282 265 283 266
rect 281 265 282 266
rect 280 265 281 266
rect 279 265 280 266
rect 278 265 279 266
rect 277 265 278 266
rect 276 265 277 266
rect 275 265 276 266
rect 274 265 275 266
rect 273 265 274 266
rect 272 265 273 266
rect 271 265 272 266
rect 270 265 271 266
rect 269 265 270 266
rect 268 265 269 266
rect 267 265 268 266
rect 266 265 267 266
rect 265 265 266 266
rect 264 265 265 266
rect 263 265 264 266
rect 262 265 263 266
rect 261 265 262 266
rect 260 265 261 266
rect 259 265 260 266
rect 258 265 259 266
rect 257 265 258 266
rect 256 265 257 266
rect 255 265 256 266
rect 254 265 255 266
rect 253 265 254 266
rect 252 265 253 266
rect 251 265 252 266
rect 250 265 251 266
rect 249 265 250 266
rect 248 265 249 266
rect 247 265 248 266
rect 246 265 247 266
rect 245 265 246 266
rect 244 265 245 266
rect 243 265 244 266
rect 242 265 243 266
rect 241 265 242 266
rect 240 265 241 266
rect 239 265 240 266
rect 238 265 239 266
rect 237 265 238 266
rect 236 265 237 266
rect 235 265 236 266
rect 234 265 235 266
rect 233 265 234 266
rect 232 265 233 266
rect 231 265 232 266
rect 230 265 231 266
rect 229 265 230 266
rect 208 265 209 266
rect 207 265 208 266
rect 206 265 207 266
rect 205 265 206 266
rect 204 265 205 266
rect 203 265 204 266
rect 202 265 203 266
rect 201 265 202 266
rect 200 265 201 266
rect 199 265 200 266
rect 198 265 199 266
rect 197 265 198 266
rect 196 265 197 266
rect 195 265 196 266
rect 194 265 195 266
rect 193 265 194 266
rect 192 265 193 266
rect 191 265 192 266
rect 190 265 191 266
rect 189 265 190 266
rect 188 265 189 266
rect 187 265 188 266
rect 186 265 187 266
rect 185 265 186 266
rect 184 265 185 266
rect 183 265 184 266
rect 182 265 183 266
rect 181 265 182 266
rect 180 265 181 266
rect 179 265 180 266
rect 178 265 179 266
rect 177 265 178 266
rect 176 265 177 266
rect 175 265 176 266
rect 174 265 175 266
rect 173 265 174 266
rect 172 265 173 266
rect 171 265 172 266
rect 170 265 171 266
rect 169 265 170 266
rect 168 265 169 266
rect 167 265 168 266
rect 166 265 167 266
rect 165 265 166 266
rect 164 265 165 266
rect 163 265 164 266
rect 162 265 163 266
rect 161 265 162 266
rect 160 265 161 266
rect 159 265 160 266
rect 158 265 159 266
rect 157 265 158 266
rect 156 265 157 266
rect 155 265 156 266
rect 154 265 155 266
rect 153 265 154 266
rect 152 265 153 266
rect 151 265 152 266
rect 150 265 151 266
rect 149 265 150 266
rect 148 265 149 266
rect 147 265 148 266
rect 146 265 147 266
rect 145 265 146 266
rect 144 265 145 266
rect 143 265 144 266
rect 142 265 143 266
rect 141 265 142 266
rect 140 265 141 266
rect 139 265 140 266
rect 138 265 139 266
rect 137 265 138 266
rect 136 265 137 266
rect 135 265 136 266
rect 134 265 135 266
rect 133 265 134 266
rect 132 265 133 266
rect 131 265 132 266
rect 130 265 131 266
rect 129 265 130 266
rect 128 265 129 266
rect 127 265 128 266
rect 126 265 127 266
rect 125 265 126 266
rect 112 265 113 266
rect 111 265 112 266
rect 110 265 111 266
rect 109 265 110 266
rect 108 265 109 266
rect 107 265 108 266
rect 106 265 107 266
rect 105 265 106 266
rect 104 265 105 266
rect 103 265 104 266
rect 102 265 103 266
rect 101 265 102 266
rect 100 265 101 266
rect 99 265 100 266
rect 98 265 99 266
rect 97 265 98 266
rect 96 265 97 266
rect 95 265 96 266
rect 94 265 95 266
rect 93 265 94 266
rect 92 265 93 266
rect 91 265 92 266
rect 90 265 91 266
rect 89 265 90 266
rect 88 265 89 266
rect 87 265 88 266
rect 86 265 87 266
rect 85 265 86 266
rect 84 265 85 266
rect 83 265 84 266
rect 82 265 83 266
rect 81 265 82 266
rect 80 265 81 266
rect 79 265 80 266
rect 78 265 79 266
rect 77 265 78 266
rect 76 265 77 266
rect 75 265 76 266
rect 74 265 75 266
rect 59 265 60 266
rect 58 265 59 266
rect 57 265 58 266
rect 56 265 57 266
rect 55 265 56 266
rect 54 265 55 266
rect 53 265 54 266
rect 52 265 53 266
rect 51 265 52 266
rect 50 265 51 266
rect 49 265 50 266
rect 48 265 49 266
rect 47 265 48 266
rect 46 265 47 266
rect 45 265 46 266
rect 44 265 45 266
rect 43 265 44 266
rect 42 265 43 266
rect 41 265 42 266
rect 40 265 41 266
rect 39 265 40 266
rect 38 265 39 266
rect 37 265 38 266
rect 26 265 27 266
rect 25 265 26 266
rect 24 265 25 266
rect 23 265 24 266
rect 22 265 23 266
rect 21 265 22 266
rect 20 265 21 266
rect 19 265 20 266
rect 18 265 19 266
rect 17 265 18 266
rect 16 265 17 266
rect 15 265 16 266
rect 14 265 15 266
rect 13 265 14 266
rect 12 265 13 266
rect 11 265 12 266
rect 10 265 11 266
rect 9 265 10 266
rect 8 265 9 266
rect 7 265 8 266
rect 6 265 7 266
rect 5 265 6 266
rect 303 266 304 267
rect 302 266 303 267
rect 301 266 302 267
rect 300 266 301 267
rect 299 266 300 267
rect 298 266 299 267
rect 297 266 298 267
rect 296 266 297 267
rect 295 266 296 267
rect 294 266 295 267
rect 293 266 294 267
rect 292 266 293 267
rect 291 266 292 267
rect 290 266 291 267
rect 289 266 290 267
rect 288 266 289 267
rect 287 266 288 267
rect 286 266 287 267
rect 285 266 286 267
rect 284 266 285 267
rect 283 266 284 267
rect 282 266 283 267
rect 281 266 282 267
rect 280 266 281 267
rect 279 266 280 267
rect 278 266 279 267
rect 277 266 278 267
rect 276 266 277 267
rect 275 266 276 267
rect 274 266 275 267
rect 273 266 274 267
rect 272 266 273 267
rect 271 266 272 267
rect 270 266 271 267
rect 269 266 270 267
rect 268 266 269 267
rect 267 266 268 267
rect 266 266 267 267
rect 265 266 266 267
rect 264 266 265 267
rect 263 266 264 267
rect 262 266 263 267
rect 261 266 262 267
rect 260 266 261 267
rect 259 266 260 267
rect 258 266 259 267
rect 257 266 258 267
rect 256 266 257 267
rect 255 266 256 267
rect 254 266 255 267
rect 253 266 254 267
rect 252 266 253 267
rect 251 266 252 267
rect 250 266 251 267
rect 249 266 250 267
rect 248 266 249 267
rect 247 266 248 267
rect 246 266 247 267
rect 245 266 246 267
rect 244 266 245 267
rect 243 266 244 267
rect 242 266 243 267
rect 241 266 242 267
rect 240 266 241 267
rect 239 266 240 267
rect 238 266 239 267
rect 237 266 238 267
rect 236 266 237 267
rect 235 266 236 267
rect 234 266 235 267
rect 233 266 234 267
rect 232 266 233 267
rect 231 266 232 267
rect 230 266 231 267
rect 229 266 230 267
rect 208 266 209 267
rect 207 266 208 267
rect 206 266 207 267
rect 205 266 206 267
rect 204 266 205 267
rect 203 266 204 267
rect 202 266 203 267
rect 201 266 202 267
rect 200 266 201 267
rect 199 266 200 267
rect 198 266 199 267
rect 197 266 198 267
rect 196 266 197 267
rect 195 266 196 267
rect 194 266 195 267
rect 193 266 194 267
rect 192 266 193 267
rect 191 266 192 267
rect 190 266 191 267
rect 189 266 190 267
rect 188 266 189 267
rect 187 266 188 267
rect 186 266 187 267
rect 185 266 186 267
rect 184 266 185 267
rect 183 266 184 267
rect 182 266 183 267
rect 181 266 182 267
rect 180 266 181 267
rect 179 266 180 267
rect 178 266 179 267
rect 177 266 178 267
rect 176 266 177 267
rect 175 266 176 267
rect 174 266 175 267
rect 173 266 174 267
rect 172 266 173 267
rect 171 266 172 267
rect 170 266 171 267
rect 169 266 170 267
rect 168 266 169 267
rect 167 266 168 267
rect 166 266 167 267
rect 165 266 166 267
rect 164 266 165 267
rect 163 266 164 267
rect 162 266 163 267
rect 161 266 162 267
rect 160 266 161 267
rect 159 266 160 267
rect 158 266 159 267
rect 157 266 158 267
rect 156 266 157 267
rect 155 266 156 267
rect 154 266 155 267
rect 153 266 154 267
rect 152 266 153 267
rect 151 266 152 267
rect 150 266 151 267
rect 149 266 150 267
rect 148 266 149 267
rect 147 266 148 267
rect 146 266 147 267
rect 145 266 146 267
rect 144 266 145 267
rect 143 266 144 267
rect 142 266 143 267
rect 141 266 142 267
rect 140 266 141 267
rect 139 266 140 267
rect 138 266 139 267
rect 137 266 138 267
rect 136 266 137 267
rect 135 266 136 267
rect 134 266 135 267
rect 133 266 134 267
rect 132 266 133 267
rect 131 266 132 267
rect 130 266 131 267
rect 129 266 130 267
rect 128 266 129 267
rect 127 266 128 267
rect 126 266 127 267
rect 125 266 126 267
rect 112 266 113 267
rect 111 266 112 267
rect 110 266 111 267
rect 109 266 110 267
rect 108 266 109 267
rect 107 266 108 267
rect 106 266 107 267
rect 105 266 106 267
rect 104 266 105 267
rect 103 266 104 267
rect 102 266 103 267
rect 101 266 102 267
rect 100 266 101 267
rect 99 266 100 267
rect 98 266 99 267
rect 97 266 98 267
rect 96 266 97 267
rect 95 266 96 267
rect 94 266 95 267
rect 93 266 94 267
rect 92 266 93 267
rect 91 266 92 267
rect 90 266 91 267
rect 89 266 90 267
rect 88 266 89 267
rect 87 266 88 267
rect 86 266 87 267
rect 85 266 86 267
rect 84 266 85 267
rect 83 266 84 267
rect 82 266 83 267
rect 81 266 82 267
rect 80 266 81 267
rect 79 266 80 267
rect 78 266 79 267
rect 77 266 78 267
rect 76 266 77 267
rect 75 266 76 267
rect 59 266 60 267
rect 58 266 59 267
rect 57 266 58 267
rect 56 266 57 267
rect 55 266 56 267
rect 54 266 55 267
rect 53 266 54 267
rect 52 266 53 267
rect 51 266 52 267
rect 50 266 51 267
rect 49 266 50 267
rect 48 266 49 267
rect 47 266 48 267
rect 46 266 47 267
rect 45 266 46 267
rect 44 266 45 267
rect 43 266 44 267
rect 42 266 43 267
rect 41 266 42 267
rect 40 266 41 267
rect 39 266 40 267
rect 38 266 39 267
rect 37 266 38 267
rect 26 266 27 267
rect 25 266 26 267
rect 24 266 25 267
rect 23 266 24 267
rect 22 266 23 267
rect 21 266 22 267
rect 20 266 21 267
rect 19 266 20 267
rect 18 266 19 267
rect 17 266 18 267
rect 16 266 17 267
rect 15 266 16 267
rect 14 266 15 267
rect 13 266 14 267
rect 12 266 13 267
rect 11 266 12 267
rect 10 266 11 267
rect 9 266 10 267
rect 8 266 9 267
rect 7 266 8 267
rect 6 266 7 267
rect 5 266 6 267
rect 302 267 303 268
rect 301 267 302 268
rect 300 267 301 268
rect 299 267 300 268
rect 298 267 299 268
rect 297 267 298 268
rect 296 267 297 268
rect 295 267 296 268
rect 294 267 295 268
rect 293 267 294 268
rect 292 267 293 268
rect 291 267 292 268
rect 290 267 291 268
rect 289 267 290 268
rect 288 267 289 268
rect 287 267 288 268
rect 286 267 287 268
rect 285 267 286 268
rect 284 267 285 268
rect 283 267 284 268
rect 282 267 283 268
rect 281 267 282 268
rect 280 267 281 268
rect 279 267 280 268
rect 278 267 279 268
rect 277 267 278 268
rect 276 267 277 268
rect 275 267 276 268
rect 274 267 275 268
rect 273 267 274 268
rect 272 267 273 268
rect 271 267 272 268
rect 270 267 271 268
rect 269 267 270 268
rect 268 267 269 268
rect 267 267 268 268
rect 266 267 267 268
rect 265 267 266 268
rect 264 267 265 268
rect 263 267 264 268
rect 262 267 263 268
rect 261 267 262 268
rect 260 267 261 268
rect 259 267 260 268
rect 258 267 259 268
rect 257 267 258 268
rect 256 267 257 268
rect 255 267 256 268
rect 254 267 255 268
rect 253 267 254 268
rect 252 267 253 268
rect 251 267 252 268
rect 250 267 251 268
rect 249 267 250 268
rect 248 267 249 268
rect 247 267 248 268
rect 246 267 247 268
rect 245 267 246 268
rect 244 267 245 268
rect 243 267 244 268
rect 242 267 243 268
rect 241 267 242 268
rect 240 267 241 268
rect 239 267 240 268
rect 238 267 239 268
rect 237 267 238 268
rect 236 267 237 268
rect 235 267 236 268
rect 234 267 235 268
rect 233 267 234 268
rect 232 267 233 268
rect 231 267 232 268
rect 230 267 231 268
rect 229 267 230 268
rect 208 267 209 268
rect 207 267 208 268
rect 206 267 207 268
rect 205 267 206 268
rect 204 267 205 268
rect 203 267 204 268
rect 202 267 203 268
rect 201 267 202 268
rect 200 267 201 268
rect 199 267 200 268
rect 198 267 199 268
rect 197 267 198 268
rect 196 267 197 268
rect 195 267 196 268
rect 194 267 195 268
rect 193 267 194 268
rect 192 267 193 268
rect 191 267 192 268
rect 190 267 191 268
rect 189 267 190 268
rect 188 267 189 268
rect 187 267 188 268
rect 186 267 187 268
rect 185 267 186 268
rect 184 267 185 268
rect 183 267 184 268
rect 182 267 183 268
rect 181 267 182 268
rect 180 267 181 268
rect 179 267 180 268
rect 178 267 179 268
rect 177 267 178 268
rect 176 267 177 268
rect 175 267 176 268
rect 174 267 175 268
rect 173 267 174 268
rect 172 267 173 268
rect 171 267 172 268
rect 170 267 171 268
rect 169 267 170 268
rect 168 267 169 268
rect 167 267 168 268
rect 166 267 167 268
rect 165 267 166 268
rect 164 267 165 268
rect 163 267 164 268
rect 162 267 163 268
rect 161 267 162 268
rect 160 267 161 268
rect 159 267 160 268
rect 158 267 159 268
rect 157 267 158 268
rect 156 267 157 268
rect 155 267 156 268
rect 154 267 155 268
rect 153 267 154 268
rect 152 267 153 268
rect 151 267 152 268
rect 150 267 151 268
rect 149 267 150 268
rect 148 267 149 268
rect 147 267 148 268
rect 146 267 147 268
rect 145 267 146 268
rect 144 267 145 268
rect 143 267 144 268
rect 142 267 143 268
rect 141 267 142 268
rect 140 267 141 268
rect 139 267 140 268
rect 138 267 139 268
rect 137 267 138 268
rect 136 267 137 268
rect 135 267 136 268
rect 134 267 135 268
rect 133 267 134 268
rect 132 267 133 268
rect 131 267 132 268
rect 130 267 131 268
rect 129 267 130 268
rect 128 267 129 268
rect 127 267 128 268
rect 126 267 127 268
rect 113 267 114 268
rect 112 267 113 268
rect 111 267 112 268
rect 110 267 111 268
rect 109 267 110 268
rect 108 267 109 268
rect 107 267 108 268
rect 106 267 107 268
rect 105 267 106 268
rect 104 267 105 268
rect 103 267 104 268
rect 102 267 103 268
rect 101 267 102 268
rect 100 267 101 268
rect 99 267 100 268
rect 98 267 99 268
rect 97 267 98 268
rect 96 267 97 268
rect 95 267 96 268
rect 94 267 95 268
rect 93 267 94 268
rect 92 267 93 268
rect 91 267 92 268
rect 90 267 91 268
rect 89 267 90 268
rect 88 267 89 268
rect 87 267 88 268
rect 86 267 87 268
rect 85 267 86 268
rect 84 267 85 268
rect 83 267 84 268
rect 82 267 83 268
rect 81 267 82 268
rect 80 267 81 268
rect 79 267 80 268
rect 78 267 79 268
rect 77 267 78 268
rect 76 267 77 268
rect 59 267 60 268
rect 58 267 59 268
rect 57 267 58 268
rect 56 267 57 268
rect 55 267 56 268
rect 54 267 55 268
rect 53 267 54 268
rect 52 267 53 268
rect 51 267 52 268
rect 50 267 51 268
rect 49 267 50 268
rect 48 267 49 268
rect 47 267 48 268
rect 46 267 47 268
rect 45 267 46 268
rect 44 267 45 268
rect 43 267 44 268
rect 42 267 43 268
rect 41 267 42 268
rect 40 267 41 268
rect 39 267 40 268
rect 38 267 39 268
rect 26 267 27 268
rect 25 267 26 268
rect 24 267 25 268
rect 23 267 24 268
rect 22 267 23 268
rect 21 267 22 268
rect 20 267 21 268
rect 19 267 20 268
rect 18 267 19 268
rect 17 267 18 268
rect 16 267 17 268
rect 15 267 16 268
rect 14 267 15 268
rect 13 267 14 268
rect 12 267 13 268
rect 11 267 12 268
rect 10 267 11 268
rect 9 267 10 268
rect 8 267 9 268
rect 7 267 8 268
rect 6 267 7 268
rect 5 267 6 268
rect 482 268 483 269
rect 462 268 463 269
rect 301 268 302 269
rect 300 268 301 269
rect 299 268 300 269
rect 298 268 299 269
rect 297 268 298 269
rect 296 268 297 269
rect 295 268 296 269
rect 294 268 295 269
rect 293 268 294 269
rect 292 268 293 269
rect 291 268 292 269
rect 290 268 291 269
rect 289 268 290 269
rect 288 268 289 269
rect 287 268 288 269
rect 286 268 287 269
rect 285 268 286 269
rect 284 268 285 269
rect 283 268 284 269
rect 282 268 283 269
rect 281 268 282 269
rect 280 268 281 269
rect 279 268 280 269
rect 278 268 279 269
rect 277 268 278 269
rect 276 268 277 269
rect 275 268 276 269
rect 274 268 275 269
rect 273 268 274 269
rect 272 268 273 269
rect 271 268 272 269
rect 270 268 271 269
rect 269 268 270 269
rect 268 268 269 269
rect 267 268 268 269
rect 266 268 267 269
rect 265 268 266 269
rect 264 268 265 269
rect 263 268 264 269
rect 262 268 263 269
rect 261 268 262 269
rect 260 268 261 269
rect 259 268 260 269
rect 258 268 259 269
rect 257 268 258 269
rect 256 268 257 269
rect 255 268 256 269
rect 254 268 255 269
rect 253 268 254 269
rect 252 268 253 269
rect 251 268 252 269
rect 250 268 251 269
rect 249 268 250 269
rect 248 268 249 269
rect 247 268 248 269
rect 246 268 247 269
rect 245 268 246 269
rect 244 268 245 269
rect 243 268 244 269
rect 242 268 243 269
rect 241 268 242 269
rect 240 268 241 269
rect 239 268 240 269
rect 238 268 239 269
rect 237 268 238 269
rect 236 268 237 269
rect 235 268 236 269
rect 234 268 235 269
rect 233 268 234 269
rect 232 268 233 269
rect 231 268 232 269
rect 230 268 231 269
rect 229 268 230 269
rect 228 268 229 269
rect 207 268 208 269
rect 206 268 207 269
rect 205 268 206 269
rect 204 268 205 269
rect 203 268 204 269
rect 202 268 203 269
rect 201 268 202 269
rect 200 268 201 269
rect 199 268 200 269
rect 198 268 199 269
rect 197 268 198 269
rect 196 268 197 269
rect 195 268 196 269
rect 194 268 195 269
rect 193 268 194 269
rect 192 268 193 269
rect 191 268 192 269
rect 190 268 191 269
rect 189 268 190 269
rect 188 268 189 269
rect 187 268 188 269
rect 186 268 187 269
rect 185 268 186 269
rect 184 268 185 269
rect 183 268 184 269
rect 182 268 183 269
rect 181 268 182 269
rect 180 268 181 269
rect 179 268 180 269
rect 178 268 179 269
rect 177 268 178 269
rect 176 268 177 269
rect 175 268 176 269
rect 174 268 175 269
rect 173 268 174 269
rect 172 268 173 269
rect 171 268 172 269
rect 170 268 171 269
rect 169 268 170 269
rect 168 268 169 269
rect 167 268 168 269
rect 166 268 167 269
rect 165 268 166 269
rect 164 268 165 269
rect 163 268 164 269
rect 162 268 163 269
rect 161 268 162 269
rect 160 268 161 269
rect 159 268 160 269
rect 158 268 159 269
rect 157 268 158 269
rect 156 268 157 269
rect 155 268 156 269
rect 154 268 155 269
rect 153 268 154 269
rect 152 268 153 269
rect 151 268 152 269
rect 150 268 151 269
rect 149 268 150 269
rect 148 268 149 269
rect 147 268 148 269
rect 146 268 147 269
rect 145 268 146 269
rect 144 268 145 269
rect 143 268 144 269
rect 142 268 143 269
rect 141 268 142 269
rect 140 268 141 269
rect 139 268 140 269
rect 138 268 139 269
rect 137 268 138 269
rect 136 268 137 269
rect 135 268 136 269
rect 134 268 135 269
rect 133 268 134 269
rect 132 268 133 269
rect 131 268 132 269
rect 130 268 131 269
rect 129 268 130 269
rect 128 268 129 269
rect 127 268 128 269
rect 126 268 127 269
rect 113 268 114 269
rect 112 268 113 269
rect 111 268 112 269
rect 110 268 111 269
rect 109 268 110 269
rect 108 268 109 269
rect 107 268 108 269
rect 106 268 107 269
rect 105 268 106 269
rect 104 268 105 269
rect 103 268 104 269
rect 102 268 103 269
rect 101 268 102 269
rect 100 268 101 269
rect 99 268 100 269
rect 98 268 99 269
rect 97 268 98 269
rect 96 268 97 269
rect 95 268 96 269
rect 94 268 95 269
rect 93 268 94 269
rect 92 268 93 269
rect 91 268 92 269
rect 90 268 91 269
rect 89 268 90 269
rect 88 268 89 269
rect 87 268 88 269
rect 86 268 87 269
rect 85 268 86 269
rect 84 268 85 269
rect 83 268 84 269
rect 82 268 83 269
rect 81 268 82 269
rect 80 268 81 269
rect 79 268 80 269
rect 78 268 79 269
rect 77 268 78 269
rect 76 268 77 269
rect 60 268 61 269
rect 59 268 60 269
rect 58 268 59 269
rect 57 268 58 269
rect 56 268 57 269
rect 55 268 56 269
rect 54 268 55 269
rect 53 268 54 269
rect 52 268 53 269
rect 51 268 52 269
rect 50 268 51 269
rect 49 268 50 269
rect 48 268 49 269
rect 47 268 48 269
rect 46 268 47 269
rect 45 268 46 269
rect 44 268 45 269
rect 43 268 44 269
rect 42 268 43 269
rect 41 268 42 269
rect 40 268 41 269
rect 39 268 40 269
rect 38 268 39 269
rect 27 268 28 269
rect 26 268 27 269
rect 25 268 26 269
rect 24 268 25 269
rect 23 268 24 269
rect 22 268 23 269
rect 21 268 22 269
rect 20 268 21 269
rect 19 268 20 269
rect 18 268 19 269
rect 17 268 18 269
rect 16 268 17 269
rect 15 268 16 269
rect 14 268 15 269
rect 13 268 14 269
rect 12 268 13 269
rect 11 268 12 269
rect 10 268 11 269
rect 9 268 10 269
rect 8 268 9 269
rect 7 268 8 269
rect 6 268 7 269
rect 5 268 6 269
rect 482 269 483 270
rect 462 269 463 270
rect 301 269 302 270
rect 300 269 301 270
rect 299 269 300 270
rect 298 269 299 270
rect 297 269 298 270
rect 296 269 297 270
rect 295 269 296 270
rect 294 269 295 270
rect 293 269 294 270
rect 292 269 293 270
rect 291 269 292 270
rect 290 269 291 270
rect 289 269 290 270
rect 288 269 289 270
rect 287 269 288 270
rect 286 269 287 270
rect 285 269 286 270
rect 284 269 285 270
rect 283 269 284 270
rect 282 269 283 270
rect 281 269 282 270
rect 280 269 281 270
rect 279 269 280 270
rect 278 269 279 270
rect 277 269 278 270
rect 276 269 277 270
rect 275 269 276 270
rect 274 269 275 270
rect 273 269 274 270
rect 272 269 273 270
rect 271 269 272 270
rect 270 269 271 270
rect 269 269 270 270
rect 268 269 269 270
rect 267 269 268 270
rect 266 269 267 270
rect 265 269 266 270
rect 264 269 265 270
rect 263 269 264 270
rect 262 269 263 270
rect 261 269 262 270
rect 260 269 261 270
rect 259 269 260 270
rect 258 269 259 270
rect 257 269 258 270
rect 256 269 257 270
rect 255 269 256 270
rect 254 269 255 270
rect 253 269 254 270
rect 252 269 253 270
rect 251 269 252 270
rect 250 269 251 270
rect 249 269 250 270
rect 248 269 249 270
rect 247 269 248 270
rect 246 269 247 270
rect 245 269 246 270
rect 244 269 245 270
rect 243 269 244 270
rect 242 269 243 270
rect 241 269 242 270
rect 240 269 241 270
rect 239 269 240 270
rect 238 269 239 270
rect 237 269 238 270
rect 236 269 237 270
rect 235 269 236 270
rect 234 269 235 270
rect 233 269 234 270
rect 232 269 233 270
rect 231 269 232 270
rect 230 269 231 270
rect 229 269 230 270
rect 228 269 229 270
rect 207 269 208 270
rect 206 269 207 270
rect 205 269 206 270
rect 204 269 205 270
rect 203 269 204 270
rect 202 269 203 270
rect 201 269 202 270
rect 200 269 201 270
rect 199 269 200 270
rect 198 269 199 270
rect 197 269 198 270
rect 196 269 197 270
rect 195 269 196 270
rect 194 269 195 270
rect 193 269 194 270
rect 192 269 193 270
rect 191 269 192 270
rect 190 269 191 270
rect 189 269 190 270
rect 188 269 189 270
rect 187 269 188 270
rect 186 269 187 270
rect 185 269 186 270
rect 184 269 185 270
rect 183 269 184 270
rect 182 269 183 270
rect 181 269 182 270
rect 180 269 181 270
rect 179 269 180 270
rect 178 269 179 270
rect 177 269 178 270
rect 176 269 177 270
rect 175 269 176 270
rect 174 269 175 270
rect 173 269 174 270
rect 172 269 173 270
rect 171 269 172 270
rect 170 269 171 270
rect 169 269 170 270
rect 168 269 169 270
rect 167 269 168 270
rect 166 269 167 270
rect 165 269 166 270
rect 164 269 165 270
rect 163 269 164 270
rect 162 269 163 270
rect 161 269 162 270
rect 160 269 161 270
rect 159 269 160 270
rect 158 269 159 270
rect 157 269 158 270
rect 156 269 157 270
rect 155 269 156 270
rect 154 269 155 270
rect 153 269 154 270
rect 152 269 153 270
rect 151 269 152 270
rect 150 269 151 270
rect 149 269 150 270
rect 148 269 149 270
rect 147 269 148 270
rect 146 269 147 270
rect 145 269 146 270
rect 144 269 145 270
rect 143 269 144 270
rect 142 269 143 270
rect 141 269 142 270
rect 140 269 141 270
rect 139 269 140 270
rect 138 269 139 270
rect 137 269 138 270
rect 136 269 137 270
rect 135 269 136 270
rect 134 269 135 270
rect 133 269 134 270
rect 132 269 133 270
rect 131 269 132 270
rect 130 269 131 270
rect 129 269 130 270
rect 128 269 129 270
rect 127 269 128 270
rect 126 269 127 270
rect 113 269 114 270
rect 112 269 113 270
rect 111 269 112 270
rect 110 269 111 270
rect 109 269 110 270
rect 108 269 109 270
rect 107 269 108 270
rect 106 269 107 270
rect 105 269 106 270
rect 104 269 105 270
rect 103 269 104 270
rect 102 269 103 270
rect 101 269 102 270
rect 100 269 101 270
rect 99 269 100 270
rect 98 269 99 270
rect 97 269 98 270
rect 96 269 97 270
rect 95 269 96 270
rect 94 269 95 270
rect 93 269 94 270
rect 92 269 93 270
rect 91 269 92 270
rect 90 269 91 270
rect 89 269 90 270
rect 88 269 89 270
rect 87 269 88 270
rect 86 269 87 270
rect 85 269 86 270
rect 84 269 85 270
rect 83 269 84 270
rect 82 269 83 270
rect 81 269 82 270
rect 80 269 81 270
rect 79 269 80 270
rect 78 269 79 270
rect 77 269 78 270
rect 60 269 61 270
rect 59 269 60 270
rect 58 269 59 270
rect 57 269 58 270
rect 56 269 57 270
rect 55 269 56 270
rect 54 269 55 270
rect 53 269 54 270
rect 52 269 53 270
rect 51 269 52 270
rect 50 269 51 270
rect 49 269 50 270
rect 48 269 49 270
rect 47 269 48 270
rect 46 269 47 270
rect 45 269 46 270
rect 44 269 45 270
rect 43 269 44 270
rect 42 269 43 270
rect 41 269 42 270
rect 40 269 41 270
rect 39 269 40 270
rect 38 269 39 270
rect 27 269 28 270
rect 26 269 27 270
rect 25 269 26 270
rect 24 269 25 270
rect 23 269 24 270
rect 22 269 23 270
rect 21 269 22 270
rect 20 269 21 270
rect 19 269 20 270
rect 18 269 19 270
rect 17 269 18 270
rect 16 269 17 270
rect 15 269 16 270
rect 14 269 15 270
rect 13 269 14 270
rect 12 269 13 270
rect 11 269 12 270
rect 10 269 11 270
rect 9 269 10 270
rect 8 269 9 270
rect 7 269 8 270
rect 6 269 7 270
rect 5 269 6 270
rect 482 270 483 271
rect 481 270 482 271
rect 463 270 464 271
rect 462 270 463 271
rect 300 270 301 271
rect 299 270 300 271
rect 298 270 299 271
rect 297 270 298 271
rect 296 270 297 271
rect 295 270 296 271
rect 294 270 295 271
rect 293 270 294 271
rect 292 270 293 271
rect 291 270 292 271
rect 290 270 291 271
rect 289 270 290 271
rect 288 270 289 271
rect 287 270 288 271
rect 286 270 287 271
rect 285 270 286 271
rect 284 270 285 271
rect 283 270 284 271
rect 282 270 283 271
rect 281 270 282 271
rect 280 270 281 271
rect 279 270 280 271
rect 278 270 279 271
rect 277 270 278 271
rect 276 270 277 271
rect 275 270 276 271
rect 274 270 275 271
rect 273 270 274 271
rect 272 270 273 271
rect 271 270 272 271
rect 270 270 271 271
rect 269 270 270 271
rect 268 270 269 271
rect 267 270 268 271
rect 266 270 267 271
rect 265 270 266 271
rect 264 270 265 271
rect 263 270 264 271
rect 262 270 263 271
rect 261 270 262 271
rect 260 270 261 271
rect 259 270 260 271
rect 258 270 259 271
rect 257 270 258 271
rect 256 270 257 271
rect 255 270 256 271
rect 254 270 255 271
rect 253 270 254 271
rect 252 270 253 271
rect 251 270 252 271
rect 250 270 251 271
rect 249 270 250 271
rect 248 270 249 271
rect 247 270 248 271
rect 246 270 247 271
rect 245 270 246 271
rect 244 270 245 271
rect 243 270 244 271
rect 242 270 243 271
rect 241 270 242 271
rect 240 270 241 271
rect 239 270 240 271
rect 238 270 239 271
rect 237 270 238 271
rect 236 270 237 271
rect 235 270 236 271
rect 234 270 235 271
rect 233 270 234 271
rect 232 270 233 271
rect 231 270 232 271
rect 230 270 231 271
rect 229 270 230 271
rect 228 270 229 271
rect 227 270 228 271
rect 206 270 207 271
rect 205 270 206 271
rect 204 270 205 271
rect 203 270 204 271
rect 202 270 203 271
rect 201 270 202 271
rect 200 270 201 271
rect 199 270 200 271
rect 198 270 199 271
rect 197 270 198 271
rect 196 270 197 271
rect 195 270 196 271
rect 194 270 195 271
rect 193 270 194 271
rect 192 270 193 271
rect 191 270 192 271
rect 190 270 191 271
rect 189 270 190 271
rect 188 270 189 271
rect 187 270 188 271
rect 186 270 187 271
rect 185 270 186 271
rect 184 270 185 271
rect 183 270 184 271
rect 182 270 183 271
rect 181 270 182 271
rect 180 270 181 271
rect 179 270 180 271
rect 178 270 179 271
rect 177 270 178 271
rect 176 270 177 271
rect 175 270 176 271
rect 174 270 175 271
rect 173 270 174 271
rect 172 270 173 271
rect 171 270 172 271
rect 170 270 171 271
rect 169 270 170 271
rect 168 270 169 271
rect 167 270 168 271
rect 166 270 167 271
rect 165 270 166 271
rect 164 270 165 271
rect 163 270 164 271
rect 162 270 163 271
rect 161 270 162 271
rect 160 270 161 271
rect 159 270 160 271
rect 158 270 159 271
rect 157 270 158 271
rect 156 270 157 271
rect 155 270 156 271
rect 154 270 155 271
rect 153 270 154 271
rect 152 270 153 271
rect 151 270 152 271
rect 150 270 151 271
rect 149 270 150 271
rect 148 270 149 271
rect 147 270 148 271
rect 146 270 147 271
rect 145 270 146 271
rect 144 270 145 271
rect 143 270 144 271
rect 142 270 143 271
rect 141 270 142 271
rect 140 270 141 271
rect 139 270 140 271
rect 138 270 139 271
rect 137 270 138 271
rect 136 270 137 271
rect 135 270 136 271
rect 134 270 135 271
rect 133 270 134 271
rect 132 270 133 271
rect 131 270 132 271
rect 130 270 131 271
rect 129 270 130 271
rect 128 270 129 271
rect 127 270 128 271
rect 126 270 127 271
rect 113 270 114 271
rect 112 270 113 271
rect 111 270 112 271
rect 110 270 111 271
rect 109 270 110 271
rect 108 270 109 271
rect 107 270 108 271
rect 106 270 107 271
rect 105 270 106 271
rect 104 270 105 271
rect 103 270 104 271
rect 102 270 103 271
rect 101 270 102 271
rect 100 270 101 271
rect 99 270 100 271
rect 98 270 99 271
rect 97 270 98 271
rect 96 270 97 271
rect 95 270 96 271
rect 94 270 95 271
rect 93 270 94 271
rect 92 270 93 271
rect 91 270 92 271
rect 90 270 91 271
rect 89 270 90 271
rect 88 270 89 271
rect 87 270 88 271
rect 86 270 87 271
rect 85 270 86 271
rect 84 270 85 271
rect 83 270 84 271
rect 82 270 83 271
rect 81 270 82 271
rect 80 270 81 271
rect 79 270 80 271
rect 78 270 79 271
rect 77 270 78 271
rect 61 270 62 271
rect 60 270 61 271
rect 59 270 60 271
rect 58 270 59 271
rect 57 270 58 271
rect 56 270 57 271
rect 55 270 56 271
rect 54 270 55 271
rect 53 270 54 271
rect 52 270 53 271
rect 51 270 52 271
rect 50 270 51 271
rect 49 270 50 271
rect 48 270 49 271
rect 47 270 48 271
rect 46 270 47 271
rect 45 270 46 271
rect 44 270 45 271
rect 43 270 44 271
rect 42 270 43 271
rect 41 270 42 271
rect 40 270 41 271
rect 39 270 40 271
rect 38 270 39 271
rect 27 270 28 271
rect 26 270 27 271
rect 25 270 26 271
rect 24 270 25 271
rect 23 270 24 271
rect 22 270 23 271
rect 21 270 22 271
rect 20 270 21 271
rect 19 270 20 271
rect 18 270 19 271
rect 17 270 18 271
rect 16 270 17 271
rect 15 270 16 271
rect 14 270 15 271
rect 13 270 14 271
rect 12 270 13 271
rect 11 270 12 271
rect 10 270 11 271
rect 9 270 10 271
rect 8 270 9 271
rect 7 270 8 271
rect 6 270 7 271
rect 5 270 6 271
rect 482 271 483 272
rect 481 271 482 272
rect 480 271 481 272
rect 479 271 480 272
rect 478 271 479 272
rect 477 271 478 272
rect 476 271 477 272
rect 475 271 476 272
rect 474 271 475 272
rect 473 271 474 272
rect 472 271 473 272
rect 471 271 472 272
rect 470 271 471 272
rect 469 271 470 272
rect 468 271 469 272
rect 467 271 468 272
rect 466 271 467 272
rect 465 271 466 272
rect 464 271 465 272
rect 463 271 464 272
rect 462 271 463 272
rect 299 271 300 272
rect 298 271 299 272
rect 297 271 298 272
rect 296 271 297 272
rect 295 271 296 272
rect 294 271 295 272
rect 293 271 294 272
rect 292 271 293 272
rect 291 271 292 272
rect 290 271 291 272
rect 289 271 290 272
rect 288 271 289 272
rect 287 271 288 272
rect 286 271 287 272
rect 285 271 286 272
rect 284 271 285 272
rect 283 271 284 272
rect 282 271 283 272
rect 281 271 282 272
rect 280 271 281 272
rect 279 271 280 272
rect 278 271 279 272
rect 277 271 278 272
rect 276 271 277 272
rect 275 271 276 272
rect 274 271 275 272
rect 273 271 274 272
rect 272 271 273 272
rect 271 271 272 272
rect 270 271 271 272
rect 269 271 270 272
rect 268 271 269 272
rect 267 271 268 272
rect 266 271 267 272
rect 265 271 266 272
rect 264 271 265 272
rect 263 271 264 272
rect 262 271 263 272
rect 261 271 262 272
rect 260 271 261 272
rect 259 271 260 272
rect 258 271 259 272
rect 257 271 258 272
rect 256 271 257 272
rect 255 271 256 272
rect 254 271 255 272
rect 253 271 254 272
rect 252 271 253 272
rect 251 271 252 272
rect 250 271 251 272
rect 249 271 250 272
rect 248 271 249 272
rect 247 271 248 272
rect 246 271 247 272
rect 245 271 246 272
rect 244 271 245 272
rect 243 271 244 272
rect 242 271 243 272
rect 241 271 242 272
rect 240 271 241 272
rect 239 271 240 272
rect 238 271 239 272
rect 237 271 238 272
rect 236 271 237 272
rect 235 271 236 272
rect 234 271 235 272
rect 233 271 234 272
rect 232 271 233 272
rect 231 271 232 272
rect 230 271 231 272
rect 229 271 230 272
rect 228 271 229 272
rect 227 271 228 272
rect 206 271 207 272
rect 205 271 206 272
rect 204 271 205 272
rect 203 271 204 272
rect 202 271 203 272
rect 201 271 202 272
rect 200 271 201 272
rect 199 271 200 272
rect 198 271 199 272
rect 197 271 198 272
rect 196 271 197 272
rect 195 271 196 272
rect 194 271 195 272
rect 193 271 194 272
rect 192 271 193 272
rect 191 271 192 272
rect 190 271 191 272
rect 189 271 190 272
rect 188 271 189 272
rect 187 271 188 272
rect 186 271 187 272
rect 185 271 186 272
rect 184 271 185 272
rect 183 271 184 272
rect 182 271 183 272
rect 181 271 182 272
rect 180 271 181 272
rect 179 271 180 272
rect 178 271 179 272
rect 177 271 178 272
rect 176 271 177 272
rect 175 271 176 272
rect 174 271 175 272
rect 173 271 174 272
rect 172 271 173 272
rect 171 271 172 272
rect 170 271 171 272
rect 169 271 170 272
rect 168 271 169 272
rect 167 271 168 272
rect 166 271 167 272
rect 165 271 166 272
rect 164 271 165 272
rect 163 271 164 272
rect 162 271 163 272
rect 161 271 162 272
rect 160 271 161 272
rect 159 271 160 272
rect 158 271 159 272
rect 157 271 158 272
rect 156 271 157 272
rect 155 271 156 272
rect 154 271 155 272
rect 153 271 154 272
rect 152 271 153 272
rect 151 271 152 272
rect 150 271 151 272
rect 149 271 150 272
rect 148 271 149 272
rect 147 271 148 272
rect 146 271 147 272
rect 145 271 146 272
rect 144 271 145 272
rect 143 271 144 272
rect 142 271 143 272
rect 141 271 142 272
rect 140 271 141 272
rect 139 271 140 272
rect 138 271 139 272
rect 137 271 138 272
rect 136 271 137 272
rect 135 271 136 272
rect 134 271 135 272
rect 133 271 134 272
rect 132 271 133 272
rect 131 271 132 272
rect 130 271 131 272
rect 129 271 130 272
rect 128 271 129 272
rect 127 271 128 272
rect 113 271 114 272
rect 112 271 113 272
rect 111 271 112 272
rect 110 271 111 272
rect 109 271 110 272
rect 108 271 109 272
rect 107 271 108 272
rect 106 271 107 272
rect 105 271 106 272
rect 104 271 105 272
rect 103 271 104 272
rect 102 271 103 272
rect 101 271 102 272
rect 100 271 101 272
rect 99 271 100 272
rect 98 271 99 272
rect 97 271 98 272
rect 96 271 97 272
rect 95 271 96 272
rect 94 271 95 272
rect 93 271 94 272
rect 92 271 93 272
rect 91 271 92 272
rect 90 271 91 272
rect 89 271 90 272
rect 88 271 89 272
rect 87 271 88 272
rect 86 271 87 272
rect 85 271 86 272
rect 84 271 85 272
rect 83 271 84 272
rect 82 271 83 272
rect 81 271 82 272
rect 80 271 81 272
rect 79 271 80 272
rect 78 271 79 272
rect 61 271 62 272
rect 60 271 61 272
rect 59 271 60 272
rect 58 271 59 272
rect 57 271 58 272
rect 56 271 57 272
rect 55 271 56 272
rect 54 271 55 272
rect 53 271 54 272
rect 52 271 53 272
rect 51 271 52 272
rect 50 271 51 272
rect 49 271 50 272
rect 48 271 49 272
rect 47 271 48 272
rect 46 271 47 272
rect 45 271 46 272
rect 44 271 45 272
rect 43 271 44 272
rect 42 271 43 272
rect 41 271 42 272
rect 40 271 41 272
rect 39 271 40 272
rect 27 271 28 272
rect 26 271 27 272
rect 25 271 26 272
rect 24 271 25 272
rect 23 271 24 272
rect 22 271 23 272
rect 21 271 22 272
rect 20 271 21 272
rect 19 271 20 272
rect 18 271 19 272
rect 17 271 18 272
rect 16 271 17 272
rect 15 271 16 272
rect 14 271 15 272
rect 13 271 14 272
rect 12 271 13 272
rect 11 271 12 272
rect 10 271 11 272
rect 9 271 10 272
rect 8 271 9 272
rect 7 271 8 272
rect 6 271 7 272
rect 5 271 6 272
rect 482 272 483 273
rect 481 272 482 273
rect 480 272 481 273
rect 479 272 480 273
rect 478 272 479 273
rect 477 272 478 273
rect 476 272 477 273
rect 475 272 476 273
rect 474 272 475 273
rect 473 272 474 273
rect 472 272 473 273
rect 471 272 472 273
rect 470 272 471 273
rect 469 272 470 273
rect 468 272 469 273
rect 467 272 468 273
rect 466 272 467 273
rect 465 272 466 273
rect 464 272 465 273
rect 463 272 464 273
rect 462 272 463 273
rect 299 272 300 273
rect 298 272 299 273
rect 297 272 298 273
rect 296 272 297 273
rect 295 272 296 273
rect 294 272 295 273
rect 293 272 294 273
rect 292 272 293 273
rect 291 272 292 273
rect 290 272 291 273
rect 289 272 290 273
rect 288 272 289 273
rect 287 272 288 273
rect 286 272 287 273
rect 285 272 286 273
rect 284 272 285 273
rect 283 272 284 273
rect 282 272 283 273
rect 281 272 282 273
rect 280 272 281 273
rect 279 272 280 273
rect 278 272 279 273
rect 277 272 278 273
rect 276 272 277 273
rect 275 272 276 273
rect 274 272 275 273
rect 273 272 274 273
rect 272 272 273 273
rect 271 272 272 273
rect 270 272 271 273
rect 269 272 270 273
rect 268 272 269 273
rect 267 272 268 273
rect 266 272 267 273
rect 265 272 266 273
rect 264 272 265 273
rect 263 272 264 273
rect 262 272 263 273
rect 261 272 262 273
rect 260 272 261 273
rect 259 272 260 273
rect 258 272 259 273
rect 257 272 258 273
rect 256 272 257 273
rect 255 272 256 273
rect 254 272 255 273
rect 253 272 254 273
rect 252 272 253 273
rect 251 272 252 273
rect 250 272 251 273
rect 249 272 250 273
rect 248 272 249 273
rect 247 272 248 273
rect 246 272 247 273
rect 245 272 246 273
rect 244 272 245 273
rect 243 272 244 273
rect 242 272 243 273
rect 241 272 242 273
rect 240 272 241 273
rect 239 272 240 273
rect 238 272 239 273
rect 237 272 238 273
rect 236 272 237 273
rect 235 272 236 273
rect 234 272 235 273
rect 233 272 234 273
rect 232 272 233 273
rect 231 272 232 273
rect 230 272 231 273
rect 229 272 230 273
rect 228 272 229 273
rect 227 272 228 273
rect 206 272 207 273
rect 205 272 206 273
rect 204 272 205 273
rect 203 272 204 273
rect 202 272 203 273
rect 201 272 202 273
rect 200 272 201 273
rect 199 272 200 273
rect 198 272 199 273
rect 197 272 198 273
rect 196 272 197 273
rect 195 272 196 273
rect 194 272 195 273
rect 193 272 194 273
rect 192 272 193 273
rect 191 272 192 273
rect 190 272 191 273
rect 189 272 190 273
rect 188 272 189 273
rect 187 272 188 273
rect 186 272 187 273
rect 185 272 186 273
rect 184 272 185 273
rect 183 272 184 273
rect 182 272 183 273
rect 181 272 182 273
rect 180 272 181 273
rect 179 272 180 273
rect 178 272 179 273
rect 177 272 178 273
rect 176 272 177 273
rect 175 272 176 273
rect 174 272 175 273
rect 173 272 174 273
rect 172 272 173 273
rect 171 272 172 273
rect 170 272 171 273
rect 169 272 170 273
rect 168 272 169 273
rect 167 272 168 273
rect 166 272 167 273
rect 165 272 166 273
rect 164 272 165 273
rect 163 272 164 273
rect 162 272 163 273
rect 161 272 162 273
rect 160 272 161 273
rect 159 272 160 273
rect 158 272 159 273
rect 157 272 158 273
rect 156 272 157 273
rect 155 272 156 273
rect 154 272 155 273
rect 153 272 154 273
rect 152 272 153 273
rect 151 272 152 273
rect 150 272 151 273
rect 149 272 150 273
rect 148 272 149 273
rect 147 272 148 273
rect 146 272 147 273
rect 145 272 146 273
rect 144 272 145 273
rect 143 272 144 273
rect 142 272 143 273
rect 141 272 142 273
rect 140 272 141 273
rect 139 272 140 273
rect 138 272 139 273
rect 137 272 138 273
rect 136 272 137 273
rect 135 272 136 273
rect 134 272 135 273
rect 133 272 134 273
rect 132 272 133 273
rect 131 272 132 273
rect 130 272 131 273
rect 129 272 130 273
rect 128 272 129 273
rect 127 272 128 273
rect 113 272 114 273
rect 112 272 113 273
rect 111 272 112 273
rect 110 272 111 273
rect 109 272 110 273
rect 108 272 109 273
rect 107 272 108 273
rect 106 272 107 273
rect 105 272 106 273
rect 104 272 105 273
rect 103 272 104 273
rect 102 272 103 273
rect 101 272 102 273
rect 100 272 101 273
rect 99 272 100 273
rect 98 272 99 273
rect 97 272 98 273
rect 96 272 97 273
rect 95 272 96 273
rect 94 272 95 273
rect 93 272 94 273
rect 92 272 93 273
rect 91 272 92 273
rect 90 272 91 273
rect 89 272 90 273
rect 88 272 89 273
rect 87 272 88 273
rect 86 272 87 273
rect 85 272 86 273
rect 84 272 85 273
rect 83 272 84 273
rect 82 272 83 273
rect 81 272 82 273
rect 80 272 81 273
rect 79 272 80 273
rect 78 272 79 273
rect 61 272 62 273
rect 60 272 61 273
rect 59 272 60 273
rect 58 272 59 273
rect 57 272 58 273
rect 56 272 57 273
rect 55 272 56 273
rect 54 272 55 273
rect 53 272 54 273
rect 52 272 53 273
rect 51 272 52 273
rect 50 272 51 273
rect 49 272 50 273
rect 48 272 49 273
rect 47 272 48 273
rect 46 272 47 273
rect 45 272 46 273
rect 44 272 45 273
rect 43 272 44 273
rect 42 272 43 273
rect 41 272 42 273
rect 40 272 41 273
rect 39 272 40 273
rect 27 272 28 273
rect 26 272 27 273
rect 25 272 26 273
rect 24 272 25 273
rect 23 272 24 273
rect 22 272 23 273
rect 21 272 22 273
rect 20 272 21 273
rect 19 272 20 273
rect 18 272 19 273
rect 17 272 18 273
rect 16 272 17 273
rect 15 272 16 273
rect 14 272 15 273
rect 13 272 14 273
rect 12 272 13 273
rect 11 272 12 273
rect 10 272 11 273
rect 9 272 10 273
rect 8 272 9 273
rect 7 272 8 273
rect 6 272 7 273
rect 5 272 6 273
rect 482 273 483 274
rect 481 273 482 274
rect 480 273 481 274
rect 479 273 480 274
rect 478 273 479 274
rect 477 273 478 274
rect 476 273 477 274
rect 475 273 476 274
rect 474 273 475 274
rect 473 273 474 274
rect 472 273 473 274
rect 471 273 472 274
rect 470 273 471 274
rect 469 273 470 274
rect 468 273 469 274
rect 467 273 468 274
rect 466 273 467 274
rect 465 273 466 274
rect 464 273 465 274
rect 463 273 464 274
rect 462 273 463 274
rect 298 273 299 274
rect 297 273 298 274
rect 296 273 297 274
rect 295 273 296 274
rect 294 273 295 274
rect 293 273 294 274
rect 292 273 293 274
rect 291 273 292 274
rect 290 273 291 274
rect 289 273 290 274
rect 288 273 289 274
rect 287 273 288 274
rect 286 273 287 274
rect 285 273 286 274
rect 284 273 285 274
rect 283 273 284 274
rect 282 273 283 274
rect 281 273 282 274
rect 280 273 281 274
rect 279 273 280 274
rect 278 273 279 274
rect 277 273 278 274
rect 276 273 277 274
rect 275 273 276 274
rect 274 273 275 274
rect 273 273 274 274
rect 272 273 273 274
rect 271 273 272 274
rect 270 273 271 274
rect 269 273 270 274
rect 268 273 269 274
rect 267 273 268 274
rect 266 273 267 274
rect 265 273 266 274
rect 264 273 265 274
rect 263 273 264 274
rect 262 273 263 274
rect 261 273 262 274
rect 260 273 261 274
rect 259 273 260 274
rect 258 273 259 274
rect 257 273 258 274
rect 256 273 257 274
rect 255 273 256 274
rect 254 273 255 274
rect 253 273 254 274
rect 252 273 253 274
rect 251 273 252 274
rect 250 273 251 274
rect 249 273 250 274
rect 248 273 249 274
rect 247 273 248 274
rect 246 273 247 274
rect 245 273 246 274
rect 244 273 245 274
rect 243 273 244 274
rect 242 273 243 274
rect 241 273 242 274
rect 240 273 241 274
rect 239 273 240 274
rect 238 273 239 274
rect 237 273 238 274
rect 236 273 237 274
rect 235 273 236 274
rect 234 273 235 274
rect 233 273 234 274
rect 232 273 233 274
rect 231 273 232 274
rect 230 273 231 274
rect 229 273 230 274
rect 228 273 229 274
rect 227 273 228 274
rect 226 273 227 274
rect 205 273 206 274
rect 204 273 205 274
rect 203 273 204 274
rect 202 273 203 274
rect 201 273 202 274
rect 200 273 201 274
rect 199 273 200 274
rect 198 273 199 274
rect 197 273 198 274
rect 196 273 197 274
rect 195 273 196 274
rect 194 273 195 274
rect 193 273 194 274
rect 192 273 193 274
rect 191 273 192 274
rect 190 273 191 274
rect 189 273 190 274
rect 188 273 189 274
rect 187 273 188 274
rect 186 273 187 274
rect 185 273 186 274
rect 184 273 185 274
rect 183 273 184 274
rect 182 273 183 274
rect 181 273 182 274
rect 180 273 181 274
rect 179 273 180 274
rect 178 273 179 274
rect 177 273 178 274
rect 176 273 177 274
rect 175 273 176 274
rect 174 273 175 274
rect 173 273 174 274
rect 172 273 173 274
rect 171 273 172 274
rect 170 273 171 274
rect 169 273 170 274
rect 168 273 169 274
rect 167 273 168 274
rect 166 273 167 274
rect 165 273 166 274
rect 164 273 165 274
rect 163 273 164 274
rect 162 273 163 274
rect 161 273 162 274
rect 160 273 161 274
rect 159 273 160 274
rect 158 273 159 274
rect 157 273 158 274
rect 156 273 157 274
rect 155 273 156 274
rect 154 273 155 274
rect 153 273 154 274
rect 152 273 153 274
rect 151 273 152 274
rect 150 273 151 274
rect 149 273 150 274
rect 148 273 149 274
rect 147 273 148 274
rect 146 273 147 274
rect 145 273 146 274
rect 144 273 145 274
rect 143 273 144 274
rect 142 273 143 274
rect 141 273 142 274
rect 140 273 141 274
rect 139 273 140 274
rect 138 273 139 274
rect 137 273 138 274
rect 136 273 137 274
rect 135 273 136 274
rect 134 273 135 274
rect 133 273 134 274
rect 132 273 133 274
rect 131 273 132 274
rect 130 273 131 274
rect 129 273 130 274
rect 128 273 129 274
rect 114 273 115 274
rect 113 273 114 274
rect 112 273 113 274
rect 111 273 112 274
rect 110 273 111 274
rect 109 273 110 274
rect 108 273 109 274
rect 107 273 108 274
rect 106 273 107 274
rect 105 273 106 274
rect 104 273 105 274
rect 103 273 104 274
rect 102 273 103 274
rect 101 273 102 274
rect 100 273 101 274
rect 99 273 100 274
rect 98 273 99 274
rect 97 273 98 274
rect 96 273 97 274
rect 95 273 96 274
rect 94 273 95 274
rect 93 273 94 274
rect 92 273 93 274
rect 91 273 92 274
rect 90 273 91 274
rect 89 273 90 274
rect 88 273 89 274
rect 87 273 88 274
rect 86 273 87 274
rect 85 273 86 274
rect 84 273 85 274
rect 83 273 84 274
rect 82 273 83 274
rect 81 273 82 274
rect 80 273 81 274
rect 79 273 80 274
rect 62 273 63 274
rect 61 273 62 274
rect 60 273 61 274
rect 59 273 60 274
rect 58 273 59 274
rect 57 273 58 274
rect 56 273 57 274
rect 55 273 56 274
rect 54 273 55 274
rect 53 273 54 274
rect 52 273 53 274
rect 51 273 52 274
rect 50 273 51 274
rect 49 273 50 274
rect 48 273 49 274
rect 47 273 48 274
rect 46 273 47 274
rect 45 273 46 274
rect 44 273 45 274
rect 43 273 44 274
rect 42 273 43 274
rect 41 273 42 274
rect 40 273 41 274
rect 39 273 40 274
rect 28 273 29 274
rect 27 273 28 274
rect 26 273 27 274
rect 25 273 26 274
rect 24 273 25 274
rect 23 273 24 274
rect 22 273 23 274
rect 21 273 22 274
rect 20 273 21 274
rect 19 273 20 274
rect 18 273 19 274
rect 17 273 18 274
rect 16 273 17 274
rect 15 273 16 274
rect 14 273 15 274
rect 13 273 14 274
rect 12 273 13 274
rect 11 273 12 274
rect 10 273 11 274
rect 9 273 10 274
rect 8 273 9 274
rect 7 273 8 274
rect 6 273 7 274
rect 5 273 6 274
rect 482 274 483 275
rect 481 274 482 275
rect 480 274 481 275
rect 479 274 480 275
rect 478 274 479 275
rect 477 274 478 275
rect 476 274 477 275
rect 475 274 476 275
rect 474 274 475 275
rect 473 274 474 275
rect 472 274 473 275
rect 471 274 472 275
rect 470 274 471 275
rect 469 274 470 275
rect 468 274 469 275
rect 467 274 468 275
rect 466 274 467 275
rect 465 274 466 275
rect 464 274 465 275
rect 463 274 464 275
rect 462 274 463 275
rect 297 274 298 275
rect 296 274 297 275
rect 295 274 296 275
rect 294 274 295 275
rect 293 274 294 275
rect 292 274 293 275
rect 291 274 292 275
rect 290 274 291 275
rect 289 274 290 275
rect 288 274 289 275
rect 287 274 288 275
rect 286 274 287 275
rect 285 274 286 275
rect 284 274 285 275
rect 283 274 284 275
rect 282 274 283 275
rect 281 274 282 275
rect 280 274 281 275
rect 279 274 280 275
rect 278 274 279 275
rect 277 274 278 275
rect 276 274 277 275
rect 275 274 276 275
rect 274 274 275 275
rect 273 274 274 275
rect 272 274 273 275
rect 271 274 272 275
rect 270 274 271 275
rect 269 274 270 275
rect 268 274 269 275
rect 267 274 268 275
rect 266 274 267 275
rect 265 274 266 275
rect 264 274 265 275
rect 263 274 264 275
rect 262 274 263 275
rect 261 274 262 275
rect 260 274 261 275
rect 259 274 260 275
rect 258 274 259 275
rect 257 274 258 275
rect 256 274 257 275
rect 255 274 256 275
rect 254 274 255 275
rect 253 274 254 275
rect 252 274 253 275
rect 251 274 252 275
rect 250 274 251 275
rect 249 274 250 275
rect 248 274 249 275
rect 247 274 248 275
rect 246 274 247 275
rect 245 274 246 275
rect 244 274 245 275
rect 243 274 244 275
rect 242 274 243 275
rect 241 274 242 275
rect 240 274 241 275
rect 239 274 240 275
rect 238 274 239 275
rect 237 274 238 275
rect 236 274 237 275
rect 235 274 236 275
rect 234 274 235 275
rect 233 274 234 275
rect 232 274 233 275
rect 231 274 232 275
rect 230 274 231 275
rect 229 274 230 275
rect 228 274 229 275
rect 227 274 228 275
rect 226 274 227 275
rect 205 274 206 275
rect 204 274 205 275
rect 203 274 204 275
rect 202 274 203 275
rect 201 274 202 275
rect 200 274 201 275
rect 199 274 200 275
rect 198 274 199 275
rect 197 274 198 275
rect 196 274 197 275
rect 195 274 196 275
rect 194 274 195 275
rect 193 274 194 275
rect 192 274 193 275
rect 191 274 192 275
rect 190 274 191 275
rect 189 274 190 275
rect 188 274 189 275
rect 187 274 188 275
rect 186 274 187 275
rect 185 274 186 275
rect 184 274 185 275
rect 183 274 184 275
rect 182 274 183 275
rect 181 274 182 275
rect 180 274 181 275
rect 179 274 180 275
rect 178 274 179 275
rect 177 274 178 275
rect 176 274 177 275
rect 175 274 176 275
rect 174 274 175 275
rect 173 274 174 275
rect 172 274 173 275
rect 171 274 172 275
rect 170 274 171 275
rect 169 274 170 275
rect 168 274 169 275
rect 167 274 168 275
rect 166 274 167 275
rect 165 274 166 275
rect 164 274 165 275
rect 163 274 164 275
rect 162 274 163 275
rect 161 274 162 275
rect 160 274 161 275
rect 159 274 160 275
rect 158 274 159 275
rect 157 274 158 275
rect 156 274 157 275
rect 155 274 156 275
rect 154 274 155 275
rect 153 274 154 275
rect 152 274 153 275
rect 151 274 152 275
rect 150 274 151 275
rect 149 274 150 275
rect 148 274 149 275
rect 147 274 148 275
rect 146 274 147 275
rect 145 274 146 275
rect 144 274 145 275
rect 143 274 144 275
rect 142 274 143 275
rect 141 274 142 275
rect 140 274 141 275
rect 139 274 140 275
rect 138 274 139 275
rect 137 274 138 275
rect 136 274 137 275
rect 135 274 136 275
rect 134 274 135 275
rect 133 274 134 275
rect 132 274 133 275
rect 131 274 132 275
rect 130 274 131 275
rect 129 274 130 275
rect 128 274 129 275
rect 114 274 115 275
rect 113 274 114 275
rect 112 274 113 275
rect 111 274 112 275
rect 110 274 111 275
rect 109 274 110 275
rect 108 274 109 275
rect 107 274 108 275
rect 106 274 107 275
rect 105 274 106 275
rect 104 274 105 275
rect 103 274 104 275
rect 102 274 103 275
rect 101 274 102 275
rect 100 274 101 275
rect 99 274 100 275
rect 98 274 99 275
rect 97 274 98 275
rect 96 274 97 275
rect 95 274 96 275
rect 94 274 95 275
rect 93 274 94 275
rect 92 274 93 275
rect 91 274 92 275
rect 90 274 91 275
rect 89 274 90 275
rect 88 274 89 275
rect 87 274 88 275
rect 86 274 87 275
rect 85 274 86 275
rect 84 274 85 275
rect 83 274 84 275
rect 82 274 83 275
rect 81 274 82 275
rect 80 274 81 275
rect 79 274 80 275
rect 62 274 63 275
rect 61 274 62 275
rect 60 274 61 275
rect 59 274 60 275
rect 58 274 59 275
rect 57 274 58 275
rect 56 274 57 275
rect 55 274 56 275
rect 54 274 55 275
rect 53 274 54 275
rect 52 274 53 275
rect 51 274 52 275
rect 50 274 51 275
rect 49 274 50 275
rect 48 274 49 275
rect 47 274 48 275
rect 46 274 47 275
rect 45 274 46 275
rect 44 274 45 275
rect 43 274 44 275
rect 42 274 43 275
rect 41 274 42 275
rect 40 274 41 275
rect 39 274 40 275
rect 28 274 29 275
rect 27 274 28 275
rect 26 274 27 275
rect 25 274 26 275
rect 24 274 25 275
rect 23 274 24 275
rect 22 274 23 275
rect 21 274 22 275
rect 20 274 21 275
rect 19 274 20 275
rect 18 274 19 275
rect 17 274 18 275
rect 16 274 17 275
rect 15 274 16 275
rect 14 274 15 275
rect 13 274 14 275
rect 12 274 13 275
rect 11 274 12 275
rect 10 274 11 275
rect 9 274 10 275
rect 8 274 9 275
rect 7 274 8 275
rect 6 274 7 275
rect 5 274 6 275
rect 482 275 483 276
rect 481 275 482 276
rect 480 275 481 276
rect 479 275 480 276
rect 478 275 479 276
rect 477 275 478 276
rect 476 275 477 276
rect 475 275 476 276
rect 474 275 475 276
rect 473 275 474 276
rect 472 275 473 276
rect 471 275 472 276
rect 470 275 471 276
rect 469 275 470 276
rect 468 275 469 276
rect 467 275 468 276
rect 466 275 467 276
rect 465 275 466 276
rect 464 275 465 276
rect 463 275 464 276
rect 462 275 463 276
rect 296 275 297 276
rect 295 275 296 276
rect 294 275 295 276
rect 293 275 294 276
rect 292 275 293 276
rect 291 275 292 276
rect 290 275 291 276
rect 289 275 290 276
rect 288 275 289 276
rect 287 275 288 276
rect 286 275 287 276
rect 285 275 286 276
rect 284 275 285 276
rect 283 275 284 276
rect 282 275 283 276
rect 281 275 282 276
rect 280 275 281 276
rect 279 275 280 276
rect 278 275 279 276
rect 277 275 278 276
rect 276 275 277 276
rect 275 275 276 276
rect 274 275 275 276
rect 273 275 274 276
rect 272 275 273 276
rect 271 275 272 276
rect 270 275 271 276
rect 269 275 270 276
rect 268 275 269 276
rect 267 275 268 276
rect 266 275 267 276
rect 265 275 266 276
rect 264 275 265 276
rect 263 275 264 276
rect 262 275 263 276
rect 261 275 262 276
rect 260 275 261 276
rect 259 275 260 276
rect 258 275 259 276
rect 257 275 258 276
rect 256 275 257 276
rect 255 275 256 276
rect 254 275 255 276
rect 253 275 254 276
rect 252 275 253 276
rect 251 275 252 276
rect 250 275 251 276
rect 249 275 250 276
rect 248 275 249 276
rect 247 275 248 276
rect 246 275 247 276
rect 245 275 246 276
rect 244 275 245 276
rect 243 275 244 276
rect 242 275 243 276
rect 241 275 242 276
rect 240 275 241 276
rect 239 275 240 276
rect 238 275 239 276
rect 237 275 238 276
rect 236 275 237 276
rect 235 275 236 276
rect 234 275 235 276
rect 233 275 234 276
rect 232 275 233 276
rect 231 275 232 276
rect 230 275 231 276
rect 229 275 230 276
rect 228 275 229 276
rect 227 275 228 276
rect 226 275 227 276
rect 225 275 226 276
rect 204 275 205 276
rect 203 275 204 276
rect 202 275 203 276
rect 201 275 202 276
rect 200 275 201 276
rect 199 275 200 276
rect 198 275 199 276
rect 197 275 198 276
rect 196 275 197 276
rect 195 275 196 276
rect 194 275 195 276
rect 193 275 194 276
rect 192 275 193 276
rect 191 275 192 276
rect 190 275 191 276
rect 189 275 190 276
rect 188 275 189 276
rect 187 275 188 276
rect 186 275 187 276
rect 185 275 186 276
rect 184 275 185 276
rect 183 275 184 276
rect 182 275 183 276
rect 181 275 182 276
rect 180 275 181 276
rect 179 275 180 276
rect 178 275 179 276
rect 177 275 178 276
rect 176 275 177 276
rect 175 275 176 276
rect 174 275 175 276
rect 173 275 174 276
rect 172 275 173 276
rect 171 275 172 276
rect 170 275 171 276
rect 169 275 170 276
rect 168 275 169 276
rect 167 275 168 276
rect 166 275 167 276
rect 165 275 166 276
rect 164 275 165 276
rect 163 275 164 276
rect 162 275 163 276
rect 161 275 162 276
rect 160 275 161 276
rect 159 275 160 276
rect 158 275 159 276
rect 157 275 158 276
rect 156 275 157 276
rect 155 275 156 276
rect 154 275 155 276
rect 153 275 154 276
rect 152 275 153 276
rect 151 275 152 276
rect 150 275 151 276
rect 149 275 150 276
rect 148 275 149 276
rect 147 275 148 276
rect 146 275 147 276
rect 145 275 146 276
rect 144 275 145 276
rect 143 275 144 276
rect 142 275 143 276
rect 141 275 142 276
rect 140 275 141 276
rect 139 275 140 276
rect 138 275 139 276
rect 137 275 138 276
rect 136 275 137 276
rect 135 275 136 276
rect 134 275 135 276
rect 133 275 134 276
rect 132 275 133 276
rect 131 275 132 276
rect 130 275 131 276
rect 129 275 130 276
rect 128 275 129 276
rect 114 275 115 276
rect 113 275 114 276
rect 112 275 113 276
rect 111 275 112 276
rect 110 275 111 276
rect 109 275 110 276
rect 108 275 109 276
rect 107 275 108 276
rect 106 275 107 276
rect 105 275 106 276
rect 104 275 105 276
rect 103 275 104 276
rect 102 275 103 276
rect 101 275 102 276
rect 100 275 101 276
rect 99 275 100 276
rect 98 275 99 276
rect 97 275 98 276
rect 96 275 97 276
rect 95 275 96 276
rect 94 275 95 276
rect 93 275 94 276
rect 92 275 93 276
rect 91 275 92 276
rect 90 275 91 276
rect 89 275 90 276
rect 88 275 89 276
rect 87 275 88 276
rect 86 275 87 276
rect 85 275 86 276
rect 84 275 85 276
rect 83 275 84 276
rect 82 275 83 276
rect 81 275 82 276
rect 80 275 81 276
rect 63 275 64 276
rect 62 275 63 276
rect 61 275 62 276
rect 60 275 61 276
rect 59 275 60 276
rect 58 275 59 276
rect 57 275 58 276
rect 56 275 57 276
rect 55 275 56 276
rect 54 275 55 276
rect 53 275 54 276
rect 52 275 53 276
rect 51 275 52 276
rect 50 275 51 276
rect 49 275 50 276
rect 48 275 49 276
rect 47 275 48 276
rect 46 275 47 276
rect 45 275 46 276
rect 44 275 45 276
rect 43 275 44 276
rect 42 275 43 276
rect 41 275 42 276
rect 40 275 41 276
rect 39 275 40 276
rect 28 275 29 276
rect 27 275 28 276
rect 26 275 27 276
rect 25 275 26 276
rect 24 275 25 276
rect 23 275 24 276
rect 22 275 23 276
rect 21 275 22 276
rect 20 275 21 276
rect 19 275 20 276
rect 18 275 19 276
rect 17 275 18 276
rect 16 275 17 276
rect 15 275 16 276
rect 14 275 15 276
rect 13 275 14 276
rect 12 275 13 276
rect 11 275 12 276
rect 10 275 11 276
rect 9 275 10 276
rect 8 275 9 276
rect 7 275 8 276
rect 6 275 7 276
rect 5 275 6 276
rect 482 276 483 277
rect 462 276 463 277
rect 441 276 442 277
rect 440 276 441 277
rect 399 276 400 277
rect 398 276 399 277
rect 397 276 398 277
rect 296 276 297 277
rect 295 276 296 277
rect 294 276 295 277
rect 293 276 294 277
rect 292 276 293 277
rect 291 276 292 277
rect 290 276 291 277
rect 289 276 290 277
rect 288 276 289 277
rect 287 276 288 277
rect 286 276 287 277
rect 285 276 286 277
rect 284 276 285 277
rect 283 276 284 277
rect 282 276 283 277
rect 281 276 282 277
rect 280 276 281 277
rect 279 276 280 277
rect 278 276 279 277
rect 277 276 278 277
rect 276 276 277 277
rect 275 276 276 277
rect 274 276 275 277
rect 273 276 274 277
rect 272 276 273 277
rect 271 276 272 277
rect 270 276 271 277
rect 269 276 270 277
rect 268 276 269 277
rect 267 276 268 277
rect 266 276 267 277
rect 265 276 266 277
rect 264 276 265 277
rect 263 276 264 277
rect 262 276 263 277
rect 261 276 262 277
rect 260 276 261 277
rect 259 276 260 277
rect 258 276 259 277
rect 257 276 258 277
rect 256 276 257 277
rect 255 276 256 277
rect 254 276 255 277
rect 253 276 254 277
rect 252 276 253 277
rect 251 276 252 277
rect 250 276 251 277
rect 249 276 250 277
rect 248 276 249 277
rect 247 276 248 277
rect 246 276 247 277
rect 245 276 246 277
rect 244 276 245 277
rect 243 276 244 277
rect 242 276 243 277
rect 241 276 242 277
rect 240 276 241 277
rect 239 276 240 277
rect 238 276 239 277
rect 237 276 238 277
rect 236 276 237 277
rect 235 276 236 277
rect 234 276 235 277
rect 233 276 234 277
rect 232 276 233 277
rect 231 276 232 277
rect 230 276 231 277
rect 229 276 230 277
rect 228 276 229 277
rect 227 276 228 277
rect 226 276 227 277
rect 225 276 226 277
rect 204 276 205 277
rect 203 276 204 277
rect 202 276 203 277
rect 201 276 202 277
rect 200 276 201 277
rect 199 276 200 277
rect 198 276 199 277
rect 197 276 198 277
rect 196 276 197 277
rect 195 276 196 277
rect 194 276 195 277
rect 193 276 194 277
rect 192 276 193 277
rect 191 276 192 277
rect 190 276 191 277
rect 189 276 190 277
rect 188 276 189 277
rect 187 276 188 277
rect 186 276 187 277
rect 185 276 186 277
rect 184 276 185 277
rect 183 276 184 277
rect 182 276 183 277
rect 181 276 182 277
rect 180 276 181 277
rect 179 276 180 277
rect 178 276 179 277
rect 177 276 178 277
rect 176 276 177 277
rect 175 276 176 277
rect 174 276 175 277
rect 173 276 174 277
rect 172 276 173 277
rect 171 276 172 277
rect 170 276 171 277
rect 169 276 170 277
rect 168 276 169 277
rect 167 276 168 277
rect 166 276 167 277
rect 165 276 166 277
rect 164 276 165 277
rect 163 276 164 277
rect 162 276 163 277
rect 161 276 162 277
rect 160 276 161 277
rect 159 276 160 277
rect 158 276 159 277
rect 157 276 158 277
rect 156 276 157 277
rect 155 276 156 277
rect 154 276 155 277
rect 153 276 154 277
rect 152 276 153 277
rect 151 276 152 277
rect 150 276 151 277
rect 149 276 150 277
rect 148 276 149 277
rect 147 276 148 277
rect 146 276 147 277
rect 145 276 146 277
rect 144 276 145 277
rect 143 276 144 277
rect 142 276 143 277
rect 141 276 142 277
rect 140 276 141 277
rect 139 276 140 277
rect 138 276 139 277
rect 137 276 138 277
rect 136 276 137 277
rect 135 276 136 277
rect 134 276 135 277
rect 133 276 134 277
rect 132 276 133 277
rect 131 276 132 277
rect 130 276 131 277
rect 129 276 130 277
rect 114 276 115 277
rect 113 276 114 277
rect 112 276 113 277
rect 111 276 112 277
rect 110 276 111 277
rect 109 276 110 277
rect 108 276 109 277
rect 107 276 108 277
rect 106 276 107 277
rect 105 276 106 277
rect 104 276 105 277
rect 103 276 104 277
rect 102 276 103 277
rect 101 276 102 277
rect 100 276 101 277
rect 99 276 100 277
rect 98 276 99 277
rect 97 276 98 277
rect 96 276 97 277
rect 95 276 96 277
rect 94 276 95 277
rect 93 276 94 277
rect 92 276 93 277
rect 91 276 92 277
rect 90 276 91 277
rect 89 276 90 277
rect 88 276 89 277
rect 87 276 88 277
rect 86 276 87 277
rect 85 276 86 277
rect 84 276 85 277
rect 83 276 84 277
rect 82 276 83 277
rect 81 276 82 277
rect 80 276 81 277
rect 63 276 64 277
rect 62 276 63 277
rect 61 276 62 277
rect 60 276 61 277
rect 59 276 60 277
rect 58 276 59 277
rect 57 276 58 277
rect 56 276 57 277
rect 55 276 56 277
rect 54 276 55 277
rect 53 276 54 277
rect 52 276 53 277
rect 51 276 52 277
rect 50 276 51 277
rect 49 276 50 277
rect 48 276 49 277
rect 47 276 48 277
rect 46 276 47 277
rect 45 276 46 277
rect 44 276 45 277
rect 43 276 44 277
rect 42 276 43 277
rect 41 276 42 277
rect 40 276 41 277
rect 39 276 40 277
rect 28 276 29 277
rect 27 276 28 277
rect 26 276 27 277
rect 25 276 26 277
rect 24 276 25 277
rect 23 276 24 277
rect 22 276 23 277
rect 21 276 22 277
rect 20 276 21 277
rect 19 276 20 277
rect 18 276 19 277
rect 17 276 18 277
rect 16 276 17 277
rect 15 276 16 277
rect 14 276 15 277
rect 13 276 14 277
rect 12 276 13 277
rect 11 276 12 277
rect 10 276 11 277
rect 9 276 10 277
rect 8 276 9 277
rect 7 276 8 277
rect 6 276 7 277
rect 5 276 6 277
rect 482 277 483 278
rect 462 277 463 278
rect 441 277 442 278
rect 440 277 441 278
rect 439 277 440 278
rect 399 277 400 278
rect 398 277 399 278
rect 397 277 398 278
rect 295 277 296 278
rect 294 277 295 278
rect 293 277 294 278
rect 292 277 293 278
rect 291 277 292 278
rect 290 277 291 278
rect 289 277 290 278
rect 288 277 289 278
rect 287 277 288 278
rect 286 277 287 278
rect 285 277 286 278
rect 284 277 285 278
rect 283 277 284 278
rect 282 277 283 278
rect 281 277 282 278
rect 280 277 281 278
rect 279 277 280 278
rect 278 277 279 278
rect 277 277 278 278
rect 276 277 277 278
rect 275 277 276 278
rect 274 277 275 278
rect 273 277 274 278
rect 272 277 273 278
rect 271 277 272 278
rect 270 277 271 278
rect 269 277 270 278
rect 268 277 269 278
rect 267 277 268 278
rect 266 277 267 278
rect 265 277 266 278
rect 264 277 265 278
rect 263 277 264 278
rect 262 277 263 278
rect 261 277 262 278
rect 260 277 261 278
rect 259 277 260 278
rect 258 277 259 278
rect 257 277 258 278
rect 256 277 257 278
rect 255 277 256 278
rect 254 277 255 278
rect 253 277 254 278
rect 252 277 253 278
rect 251 277 252 278
rect 250 277 251 278
rect 249 277 250 278
rect 248 277 249 278
rect 247 277 248 278
rect 246 277 247 278
rect 245 277 246 278
rect 244 277 245 278
rect 243 277 244 278
rect 242 277 243 278
rect 241 277 242 278
rect 240 277 241 278
rect 239 277 240 278
rect 238 277 239 278
rect 237 277 238 278
rect 236 277 237 278
rect 235 277 236 278
rect 234 277 235 278
rect 233 277 234 278
rect 232 277 233 278
rect 231 277 232 278
rect 230 277 231 278
rect 229 277 230 278
rect 228 277 229 278
rect 227 277 228 278
rect 226 277 227 278
rect 225 277 226 278
rect 224 277 225 278
rect 203 277 204 278
rect 202 277 203 278
rect 201 277 202 278
rect 200 277 201 278
rect 199 277 200 278
rect 198 277 199 278
rect 197 277 198 278
rect 196 277 197 278
rect 195 277 196 278
rect 194 277 195 278
rect 193 277 194 278
rect 192 277 193 278
rect 191 277 192 278
rect 190 277 191 278
rect 189 277 190 278
rect 188 277 189 278
rect 187 277 188 278
rect 186 277 187 278
rect 185 277 186 278
rect 184 277 185 278
rect 183 277 184 278
rect 182 277 183 278
rect 181 277 182 278
rect 180 277 181 278
rect 179 277 180 278
rect 178 277 179 278
rect 177 277 178 278
rect 176 277 177 278
rect 175 277 176 278
rect 174 277 175 278
rect 173 277 174 278
rect 172 277 173 278
rect 171 277 172 278
rect 170 277 171 278
rect 169 277 170 278
rect 168 277 169 278
rect 167 277 168 278
rect 166 277 167 278
rect 165 277 166 278
rect 164 277 165 278
rect 163 277 164 278
rect 162 277 163 278
rect 161 277 162 278
rect 160 277 161 278
rect 159 277 160 278
rect 158 277 159 278
rect 157 277 158 278
rect 156 277 157 278
rect 155 277 156 278
rect 154 277 155 278
rect 153 277 154 278
rect 152 277 153 278
rect 151 277 152 278
rect 150 277 151 278
rect 149 277 150 278
rect 148 277 149 278
rect 147 277 148 278
rect 146 277 147 278
rect 145 277 146 278
rect 144 277 145 278
rect 143 277 144 278
rect 142 277 143 278
rect 141 277 142 278
rect 140 277 141 278
rect 139 277 140 278
rect 138 277 139 278
rect 137 277 138 278
rect 136 277 137 278
rect 135 277 136 278
rect 134 277 135 278
rect 133 277 134 278
rect 132 277 133 278
rect 131 277 132 278
rect 130 277 131 278
rect 129 277 130 278
rect 114 277 115 278
rect 113 277 114 278
rect 112 277 113 278
rect 111 277 112 278
rect 110 277 111 278
rect 109 277 110 278
rect 108 277 109 278
rect 107 277 108 278
rect 106 277 107 278
rect 105 277 106 278
rect 104 277 105 278
rect 103 277 104 278
rect 102 277 103 278
rect 101 277 102 278
rect 100 277 101 278
rect 99 277 100 278
rect 98 277 99 278
rect 97 277 98 278
rect 96 277 97 278
rect 95 277 96 278
rect 94 277 95 278
rect 93 277 94 278
rect 92 277 93 278
rect 91 277 92 278
rect 90 277 91 278
rect 89 277 90 278
rect 88 277 89 278
rect 87 277 88 278
rect 86 277 87 278
rect 85 277 86 278
rect 84 277 85 278
rect 83 277 84 278
rect 82 277 83 278
rect 81 277 82 278
rect 64 277 65 278
rect 63 277 64 278
rect 62 277 63 278
rect 61 277 62 278
rect 60 277 61 278
rect 59 277 60 278
rect 58 277 59 278
rect 57 277 58 278
rect 56 277 57 278
rect 55 277 56 278
rect 54 277 55 278
rect 53 277 54 278
rect 52 277 53 278
rect 51 277 52 278
rect 50 277 51 278
rect 49 277 50 278
rect 48 277 49 278
rect 47 277 48 278
rect 46 277 47 278
rect 45 277 46 278
rect 44 277 45 278
rect 43 277 44 278
rect 42 277 43 278
rect 41 277 42 278
rect 40 277 41 278
rect 29 277 30 278
rect 28 277 29 278
rect 27 277 28 278
rect 26 277 27 278
rect 25 277 26 278
rect 24 277 25 278
rect 23 277 24 278
rect 22 277 23 278
rect 21 277 22 278
rect 20 277 21 278
rect 19 277 20 278
rect 18 277 19 278
rect 17 277 18 278
rect 16 277 17 278
rect 15 277 16 278
rect 14 277 15 278
rect 13 277 14 278
rect 12 277 13 278
rect 11 277 12 278
rect 10 277 11 278
rect 9 277 10 278
rect 8 277 9 278
rect 7 277 8 278
rect 6 277 7 278
rect 5 277 6 278
rect 441 278 442 279
rect 440 278 441 279
rect 439 278 440 279
rect 399 278 400 279
rect 398 278 399 279
rect 397 278 398 279
rect 294 278 295 279
rect 293 278 294 279
rect 292 278 293 279
rect 291 278 292 279
rect 290 278 291 279
rect 289 278 290 279
rect 288 278 289 279
rect 287 278 288 279
rect 286 278 287 279
rect 285 278 286 279
rect 284 278 285 279
rect 283 278 284 279
rect 282 278 283 279
rect 281 278 282 279
rect 280 278 281 279
rect 279 278 280 279
rect 278 278 279 279
rect 277 278 278 279
rect 276 278 277 279
rect 275 278 276 279
rect 274 278 275 279
rect 273 278 274 279
rect 272 278 273 279
rect 271 278 272 279
rect 270 278 271 279
rect 269 278 270 279
rect 268 278 269 279
rect 267 278 268 279
rect 266 278 267 279
rect 265 278 266 279
rect 264 278 265 279
rect 263 278 264 279
rect 262 278 263 279
rect 261 278 262 279
rect 260 278 261 279
rect 259 278 260 279
rect 258 278 259 279
rect 257 278 258 279
rect 256 278 257 279
rect 255 278 256 279
rect 254 278 255 279
rect 253 278 254 279
rect 252 278 253 279
rect 251 278 252 279
rect 250 278 251 279
rect 249 278 250 279
rect 248 278 249 279
rect 247 278 248 279
rect 246 278 247 279
rect 245 278 246 279
rect 244 278 245 279
rect 243 278 244 279
rect 242 278 243 279
rect 241 278 242 279
rect 240 278 241 279
rect 239 278 240 279
rect 238 278 239 279
rect 237 278 238 279
rect 236 278 237 279
rect 235 278 236 279
rect 234 278 235 279
rect 233 278 234 279
rect 232 278 233 279
rect 231 278 232 279
rect 230 278 231 279
rect 229 278 230 279
rect 228 278 229 279
rect 227 278 228 279
rect 226 278 227 279
rect 225 278 226 279
rect 224 278 225 279
rect 203 278 204 279
rect 202 278 203 279
rect 201 278 202 279
rect 200 278 201 279
rect 199 278 200 279
rect 198 278 199 279
rect 197 278 198 279
rect 196 278 197 279
rect 195 278 196 279
rect 194 278 195 279
rect 193 278 194 279
rect 192 278 193 279
rect 191 278 192 279
rect 190 278 191 279
rect 189 278 190 279
rect 188 278 189 279
rect 187 278 188 279
rect 186 278 187 279
rect 185 278 186 279
rect 184 278 185 279
rect 183 278 184 279
rect 182 278 183 279
rect 181 278 182 279
rect 180 278 181 279
rect 179 278 180 279
rect 178 278 179 279
rect 177 278 178 279
rect 176 278 177 279
rect 175 278 176 279
rect 174 278 175 279
rect 173 278 174 279
rect 172 278 173 279
rect 171 278 172 279
rect 170 278 171 279
rect 169 278 170 279
rect 168 278 169 279
rect 167 278 168 279
rect 166 278 167 279
rect 165 278 166 279
rect 164 278 165 279
rect 163 278 164 279
rect 162 278 163 279
rect 161 278 162 279
rect 160 278 161 279
rect 159 278 160 279
rect 158 278 159 279
rect 157 278 158 279
rect 156 278 157 279
rect 155 278 156 279
rect 154 278 155 279
rect 153 278 154 279
rect 152 278 153 279
rect 151 278 152 279
rect 150 278 151 279
rect 149 278 150 279
rect 148 278 149 279
rect 147 278 148 279
rect 146 278 147 279
rect 145 278 146 279
rect 144 278 145 279
rect 143 278 144 279
rect 142 278 143 279
rect 141 278 142 279
rect 140 278 141 279
rect 139 278 140 279
rect 138 278 139 279
rect 137 278 138 279
rect 136 278 137 279
rect 135 278 136 279
rect 134 278 135 279
rect 133 278 134 279
rect 132 278 133 279
rect 131 278 132 279
rect 130 278 131 279
rect 129 278 130 279
rect 115 278 116 279
rect 114 278 115 279
rect 113 278 114 279
rect 112 278 113 279
rect 111 278 112 279
rect 110 278 111 279
rect 109 278 110 279
rect 108 278 109 279
rect 107 278 108 279
rect 106 278 107 279
rect 105 278 106 279
rect 104 278 105 279
rect 103 278 104 279
rect 102 278 103 279
rect 101 278 102 279
rect 100 278 101 279
rect 99 278 100 279
rect 98 278 99 279
rect 97 278 98 279
rect 96 278 97 279
rect 95 278 96 279
rect 94 278 95 279
rect 93 278 94 279
rect 92 278 93 279
rect 91 278 92 279
rect 90 278 91 279
rect 89 278 90 279
rect 88 278 89 279
rect 87 278 88 279
rect 86 278 87 279
rect 85 278 86 279
rect 84 278 85 279
rect 83 278 84 279
rect 82 278 83 279
rect 81 278 82 279
rect 64 278 65 279
rect 63 278 64 279
rect 62 278 63 279
rect 61 278 62 279
rect 60 278 61 279
rect 59 278 60 279
rect 58 278 59 279
rect 57 278 58 279
rect 56 278 57 279
rect 55 278 56 279
rect 54 278 55 279
rect 53 278 54 279
rect 52 278 53 279
rect 51 278 52 279
rect 50 278 51 279
rect 49 278 50 279
rect 48 278 49 279
rect 47 278 48 279
rect 46 278 47 279
rect 45 278 46 279
rect 44 278 45 279
rect 43 278 44 279
rect 42 278 43 279
rect 41 278 42 279
rect 40 278 41 279
rect 29 278 30 279
rect 28 278 29 279
rect 27 278 28 279
rect 26 278 27 279
rect 25 278 26 279
rect 24 278 25 279
rect 23 278 24 279
rect 22 278 23 279
rect 21 278 22 279
rect 20 278 21 279
rect 19 278 20 279
rect 18 278 19 279
rect 17 278 18 279
rect 16 278 17 279
rect 15 278 16 279
rect 14 278 15 279
rect 13 278 14 279
rect 12 278 13 279
rect 11 278 12 279
rect 10 278 11 279
rect 9 278 10 279
rect 8 278 9 279
rect 7 278 8 279
rect 6 278 7 279
rect 5 278 6 279
rect 441 279 442 280
rect 440 279 441 280
rect 439 279 440 280
rect 399 279 400 280
rect 398 279 399 280
rect 397 279 398 280
rect 293 279 294 280
rect 292 279 293 280
rect 291 279 292 280
rect 290 279 291 280
rect 289 279 290 280
rect 288 279 289 280
rect 287 279 288 280
rect 286 279 287 280
rect 285 279 286 280
rect 284 279 285 280
rect 283 279 284 280
rect 282 279 283 280
rect 281 279 282 280
rect 280 279 281 280
rect 279 279 280 280
rect 278 279 279 280
rect 277 279 278 280
rect 276 279 277 280
rect 275 279 276 280
rect 274 279 275 280
rect 273 279 274 280
rect 272 279 273 280
rect 271 279 272 280
rect 270 279 271 280
rect 269 279 270 280
rect 268 279 269 280
rect 267 279 268 280
rect 266 279 267 280
rect 265 279 266 280
rect 264 279 265 280
rect 263 279 264 280
rect 262 279 263 280
rect 261 279 262 280
rect 260 279 261 280
rect 259 279 260 280
rect 258 279 259 280
rect 257 279 258 280
rect 256 279 257 280
rect 255 279 256 280
rect 254 279 255 280
rect 253 279 254 280
rect 252 279 253 280
rect 251 279 252 280
rect 250 279 251 280
rect 249 279 250 280
rect 248 279 249 280
rect 247 279 248 280
rect 246 279 247 280
rect 245 279 246 280
rect 244 279 245 280
rect 243 279 244 280
rect 242 279 243 280
rect 241 279 242 280
rect 240 279 241 280
rect 239 279 240 280
rect 238 279 239 280
rect 237 279 238 280
rect 236 279 237 280
rect 235 279 236 280
rect 234 279 235 280
rect 233 279 234 280
rect 232 279 233 280
rect 231 279 232 280
rect 230 279 231 280
rect 229 279 230 280
rect 228 279 229 280
rect 227 279 228 280
rect 226 279 227 280
rect 225 279 226 280
rect 224 279 225 280
rect 202 279 203 280
rect 201 279 202 280
rect 200 279 201 280
rect 199 279 200 280
rect 198 279 199 280
rect 197 279 198 280
rect 196 279 197 280
rect 195 279 196 280
rect 194 279 195 280
rect 193 279 194 280
rect 192 279 193 280
rect 191 279 192 280
rect 190 279 191 280
rect 189 279 190 280
rect 188 279 189 280
rect 187 279 188 280
rect 186 279 187 280
rect 185 279 186 280
rect 184 279 185 280
rect 183 279 184 280
rect 182 279 183 280
rect 181 279 182 280
rect 180 279 181 280
rect 179 279 180 280
rect 178 279 179 280
rect 177 279 178 280
rect 176 279 177 280
rect 175 279 176 280
rect 174 279 175 280
rect 173 279 174 280
rect 172 279 173 280
rect 171 279 172 280
rect 170 279 171 280
rect 169 279 170 280
rect 168 279 169 280
rect 167 279 168 280
rect 166 279 167 280
rect 165 279 166 280
rect 164 279 165 280
rect 163 279 164 280
rect 162 279 163 280
rect 161 279 162 280
rect 160 279 161 280
rect 159 279 160 280
rect 158 279 159 280
rect 157 279 158 280
rect 156 279 157 280
rect 155 279 156 280
rect 154 279 155 280
rect 153 279 154 280
rect 152 279 153 280
rect 151 279 152 280
rect 150 279 151 280
rect 149 279 150 280
rect 148 279 149 280
rect 147 279 148 280
rect 146 279 147 280
rect 145 279 146 280
rect 144 279 145 280
rect 143 279 144 280
rect 142 279 143 280
rect 141 279 142 280
rect 140 279 141 280
rect 139 279 140 280
rect 138 279 139 280
rect 137 279 138 280
rect 136 279 137 280
rect 135 279 136 280
rect 134 279 135 280
rect 133 279 134 280
rect 132 279 133 280
rect 131 279 132 280
rect 130 279 131 280
rect 115 279 116 280
rect 114 279 115 280
rect 113 279 114 280
rect 112 279 113 280
rect 111 279 112 280
rect 110 279 111 280
rect 109 279 110 280
rect 108 279 109 280
rect 107 279 108 280
rect 106 279 107 280
rect 105 279 106 280
rect 104 279 105 280
rect 103 279 104 280
rect 102 279 103 280
rect 101 279 102 280
rect 100 279 101 280
rect 99 279 100 280
rect 98 279 99 280
rect 97 279 98 280
rect 96 279 97 280
rect 95 279 96 280
rect 94 279 95 280
rect 93 279 94 280
rect 92 279 93 280
rect 91 279 92 280
rect 90 279 91 280
rect 89 279 90 280
rect 88 279 89 280
rect 87 279 88 280
rect 86 279 87 280
rect 85 279 86 280
rect 84 279 85 280
rect 83 279 84 280
rect 82 279 83 280
rect 81 279 82 280
rect 64 279 65 280
rect 63 279 64 280
rect 62 279 63 280
rect 61 279 62 280
rect 60 279 61 280
rect 59 279 60 280
rect 58 279 59 280
rect 57 279 58 280
rect 56 279 57 280
rect 55 279 56 280
rect 54 279 55 280
rect 53 279 54 280
rect 52 279 53 280
rect 51 279 52 280
rect 50 279 51 280
rect 49 279 50 280
rect 48 279 49 280
rect 47 279 48 280
rect 46 279 47 280
rect 45 279 46 280
rect 44 279 45 280
rect 43 279 44 280
rect 42 279 43 280
rect 41 279 42 280
rect 40 279 41 280
rect 29 279 30 280
rect 28 279 29 280
rect 27 279 28 280
rect 26 279 27 280
rect 25 279 26 280
rect 24 279 25 280
rect 23 279 24 280
rect 22 279 23 280
rect 21 279 22 280
rect 20 279 21 280
rect 19 279 20 280
rect 18 279 19 280
rect 17 279 18 280
rect 16 279 17 280
rect 15 279 16 280
rect 14 279 15 280
rect 13 279 14 280
rect 12 279 13 280
rect 11 279 12 280
rect 10 279 11 280
rect 9 279 10 280
rect 8 279 9 280
rect 7 279 8 280
rect 6 279 7 280
rect 5 279 6 280
rect 441 280 442 281
rect 440 280 441 281
rect 439 280 440 281
rect 400 280 401 281
rect 399 280 400 281
rect 398 280 399 281
rect 397 280 398 281
rect 292 280 293 281
rect 291 280 292 281
rect 290 280 291 281
rect 289 280 290 281
rect 288 280 289 281
rect 287 280 288 281
rect 286 280 287 281
rect 285 280 286 281
rect 284 280 285 281
rect 283 280 284 281
rect 282 280 283 281
rect 281 280 282 281
rect 280 280 281 281
rect 279 280 280 281
rect 278 280 279 281
rect 277 280 278 281
rect 276 280 277 281
rect 275 280 276 281
rect 274 280 275 281
rect 273 280 274 281
rect 272 280 273 281
rect 271 280 272 281
rect 270 280 271 281
rect 269 280 270 281
rect 268 280 269 281
rect 267 280 268 281
rect 266 280 267 281
rect 265 280 266 281
rect 264 280 265 281
rect 263 280 264 281
rect 262 280 263 281
rect 261 280 262 281
rect 260 280 261 281
rect 259 280 260 281
rect 258 280 259 281
rect 257 280 258 281
rect 256 280 257 281
rect 255 280 256 281
rect 254 280 255 281
rect 253 280 254 281
rect 252 280 253 281
rect 251 280 252 281
rect 250 280 251 281
rect 249 280 250 281
rect 248 280 249 281
rect 247 280 248 281
rect 246 280 247 281
rect 245 280 246 281
rect 244 280 245 281
rect 243 280 244 281
rect 242 280 243 281
rect 241 280 242 281
rect 240 280 241 281
rect 239 280 240 281
rect 238 280 239 281
rect 237 280 238 281
rect 236 280 237 281
rect 235 280 236 281
rect 234 280 235 281
rect 233 280 234 281
rect 232 280 233 281
rect 231 280 232 281
rect 230 280 231 281
rect 229 280 230 281
rect 228 280 229 281
rect 227 280 228 281
rect 226 280 227 281
rect 225 280 226 281
rect 224 280 225 281
rect 223 280 224 281
rect 201 280 202 281
rect 200 280 201 281
rect 199 280 200 281
rect 198 280 199 281
rect 197 280 198 281
rect 196 280 197 281
rect 195 280 196 281
rect 194 280 195 281
rect 193 280 194 281
rect 192 280 193 281
rect 191 280 192 281
rect 190 280 191 281
rect 189 280 190 281
rect 188 280 189 281
rect 187 280 188 281
rect 186 280 187 281
rect 185 280 186 281
rect 184 280 185 281
rect 183 280 184 281
rect 182 280 183 281
rect 181 280 182 281
rect 180 280 181 281
rect 179 280 180 281
rect 178 280 179 281
rect 177 280 178 281
rect 176 280 177 281
rect 175 280 176 281
rect 174 280 175 281
rect 173 280 174 281
rect 172 280 173 281
rect 171 280 172 281
rect 170 280 171 281
rect 169 280 170 281
rect 168 280 169 281
rect 167 280 168 281
rect 166 280 167 281
rect 165 280 166 281
rect 164 280 165 281
rect 163 280 164 281
rect 162 280 163 281
rect 161 280 162 281
rect 160 280 161 281
rect 159 280 160 281
rect 158 280 159 281
rect 157 280 158 281
rect 156 280 157 281
rect 155 280 156 281
rect 154 280 155 281
rect 153 280 154 281
rect 152 280 153 281
rect 151 280 152 281
rect 150 280 151 281
rect 149 280 150 281
rect 148 280 149 281
rect 147 280 148 281
rect 146 280 147 281
rect 145 280 146 281
rect 144 280 145 281
rect 143 280 144 281
rect 142 280 143 281
rect 141 280 142 281
rect 140 280 141 281
rect 139 280 140 281
rect 138 280 139 281
rect 137 280 138 281
rect 136 280 137 281
rect 135 280 136 281
rect 134 280 135 281
rect 133 280 134 281
rect 132 280 133 281
rect 131 280 132 281
rect 130 280 131 281
rect 115 280 116 281
rect 114 280 115 281
rect 113 280 114 281
rect 112 280 113 281
rect 111 280 112 281
rect 110 280 111 281
rect 109 280 110 281
rect 108 280 109 281
rect 107 280 108 281
rect 106 280 107 281
rect 105 280 106 281
rect 104 280 105 281
rect 103 280 104 281
rect 102 280 103 281
rect 101 280 102 281
rect 100 280 101 281
rect 99 280 100 281
rect 98 280 99 281
rect 97 280 98 281
rect 96 280 97 281
rect 95 280 96 281
rect 94 280 95 281
rect 93 280 94 281
rect 92 280 93 281
rect 91 280 92 281
rect 90 280 91 281
rect 89 280 90 281
rect 88 280 89 281
rect 87 280 88 281
rect 86 280 87 281
rect 85 280 86 281
rect 84 280 85 281
rect 83 280 84 281
rect 82 280 83 281
rect 65 280 66 281
rect 64 280 65 281
rect 63 280 64 281
rect 62 280 63 281
rect 61 280 62 281
rect 60 280 61 281
rect 59 280 60 281
rect 58 280 59 281
rect 57 280 58 281
rect 56 280 57 281
rect 55 280 56 281
rect 54 280 55 281
rect 53 280 54 281
rect 52 280 53 281
rect 51 280 52 281
rect 50 280 51 281
rect 49 280 50 281
rect 48 280 49 281
rect 47 280 48 281
rect 46 280 47 281
rect 45 280 46 281
rect 44 280 45 281
rect 43 280 44 281
rect 42 280 43 281
rect 41 280 42 281
rect 40 280 41 281
rect 29 280 30 281
rect 28 280 29 281
rect 27 280 28 281
rect 26 280 27 281
rect 25 280 26 281
rect 24 280 25 281
rect 23 280 24 281
rect 22 280 23 281
rect 21 280 22 281
rect 20 280 21 281
rect 19 280 20 281
rect 18 280 19 281
rect 17 280 18 281
rect 16 280 17 281
rect 15 280 16 281
rect 14 280 15 281
rect 13 280 14 281
rect 12 280 13 281
rect 11 280 12 281
rect 10 280 11 281
rect 9 280 10 281
rect 8 280 9 281
rect 7 280 8 281
rect 6 280 7 281
rect 5 280 6 281
rect 441 281 442 282
rect 440 281 441 282
rect 439 281 440 282
rect 438 281 439 282
rect 437 281 438 282
rect 401 281 402 282
rect 400 281 401 282
rect 399 281 400 282
rect 398 281 399 282
rect 397 281 398 282
rect 292 281 293 282
rect 291 281 292 282
rect 290 281 291 282
rect 289 281 290 282
rect 288 281 289 282
rect 287 281 288 282
rect 286 281 287 282
rect 285 281 286 282
rect 284 281 285 282
rect 283 281 284 282
rect 282 281 283 282
rect 281 281 282 282
rect 280 281 281 282
rect 279 281 280 282
rect 278 281 279 282
rect 277 281 278 282
rect 276 281 277 282
rect 275 281 276 282
rect 274 281 275 282
rect 273 281 274 282
rect 272 281 273 282
rect 271 281 272 282
rect 270 281 271 282
rect 269 281 270 282
rect 268 281 269 282
rect 267 281 268 282
rect 266 281 267 282
rect 265 281 266 282
rect 264 281 265 282
rect 263 281 264 282
rect 262 281 263 282
rect 261 281 262 282
rect 260 281 261 282
rect 259 281 260 282
rect 258 281 259 282
rect 257 281 258 282
rect 256 281 257 282
rect 255 281 256 282
rect 254 281 255 282
rect 253 281 254 282
rect 252 281 253 282
rect 251 281 252 282
rect 250 281 251 282
rect 249 281 250 282
rect 248 281 249 282
rect 247 281 248 282
rect 246 281 247 282
rect 245 281 246 282
rect 244 281 245 282
rect 243 281 244 282
rect 242 281 243 282
rect 241 281 242 282
rect 240 281 241 282
rect 239 281 240 282
rect 238 281 239 282
rect 237 281 238 282
rect 236 281 237 282
rect 235 281 236 282
rect 234 281 235 282
rect 233 281 234 282
rect 232 281 233 282
rect 231 281 232 282
rect 230 281 231 282
rect 229 281 230 282
rect 228 281 229 282
rect 227 281 228 282
rect 226 281 227 282
rect 225 281 226 282
rect 224 281 225 282
rect 223 281 224 282
rect 201 281 202 282
rect 200 281 201 282
rect 199 281 200 282
rect 198 281 199 282
rect 197 281 198 282
rect 196 281 197 282
rect 195 281 196 282
rect 194 281 195 282
rect 193 281 194 282
rect 192 281 193 282
rect 191 281 192 282
rect 190 281 191 282
rect 189 281 190 282
rect 188 281 189 282
rect 187 281 188 282
rect 186 281 187 282
rect 185 281 186 282
rect 184 281 185 282
rect 183 281 184 282
rect 182 281 183 282
rect 181 281 182 282
rect 180 281 181 282
rect 179 281 180 282
rect 178 281 179 282
rect 177 281 178 282
rect 176 281 177 282
rect 175 281 176 282
rect 174 281 175 282
rect 173 281 174 282
rect 172 281 173 282
rect 171 281 172 282
rect 170 281 171 282
rect 169 281 170 282
rect 168 281 169 282
rect 167 281 168 282
rect 166 281 167 282
rect 165 281 166 282
rect 164 281 165 282
rect 163 281 164 282
rect 162 281 163 282
rect 161 281 162 282
rect 160 281 161 282
rect 159 281 160 282
rect 158 281 159 282
rect 157 281 158 282
rect 156 281 157 282
rect 155 281 156 282
rect 154 281 155 282
rect 153 281 154 282
rect 152 281 153 282
rect 151 281 152 282
rect 150 281 151 282
rect 149 281 150 282
rect 148 281 149 282
rect 147 281 148 282
rect 146 281 147 282
rect 145 281 146 282
rect 144 281 145 282
rect 143 281 144 282
rect 142 281 143 282
rect 141 281 142 282
rect 140 281 141 282
rect 139 281 140 282
rect 138 281 139 282
rect 137 281 138 282
rect 136 281 137 282
rect 135 281 136 282
rect 134 281 135 282
rect 133 281 134 282
rect 132 281 133 282
rect 131 281 132 282
rect 116 281 117 282
rect 115 281 116 282
rect 114 281 115 282
rect 113 281 114 282
rect 112 281 113 282
rect 111 281 112 282
rect 110 281 111 282
rect 109 281 110 282
rect 108 281 109 282
rect 107 281 108 282
rect 106 281 107 282
rect 105 281 106 282
rect 104 281 105 282
rect 103 281 104 282
rect 102 281 103 282
rect 101 281 102 282
rect 100 281 101 282
rect 99 281 100 282
rect 98 281 99 282
rect 97 281 98 282
rect 96 281 97 282
rect 95 281 96 282
rect 94 281 95 282
rect 93 281 94 282
rect 92 281 93 282
rect 91 281 92 282
rect 90 281 91 282
rect 89 281 90 282
rect 88 281 89 282
rect 87 281 88 282
rect 86 281 87 282
rect 85 281 86 282
rect 84 281 85 282
rect 83 281 84 282
rect 82 281 83 282
rect 65 281 66 282
rect 64 281 65 282
rect 63 281 64 282
rect 62 281 63 282
rect 61 281 62 282
rect 60 281 61 282
rect 59 281 60 282
rect 58 281 59 282
rect 57 281 58 282
rect 56 281 57 282
rect 55 281 56 282
rect 54 281 55 282
rect 53 281 54 282
rect 52 281 53 282
rect 51 281 52 282
rect 50 281 51 282
rect 49 281 50 282
rect 48 281 49 282
rect 47 281 48 282
rect 46 281 47 282
rect 45 281 46 282
rect 44 281 45 282
rect 43 281 44 282
rect 42 281 43 282
rect 41 281 42 282
rect 40 281 41 282
rect 29 281 30 282
rect 28 281 29 282
rect 27 281 28 282
rect 26 281 27 282
rect 25 281 26 282
rect 24 281 25 282
rect 23 281 24 282
rect 22 281 23 282
rect 21 281 22 282
rect 20 281 21 282
rect 19 281 20 282
rect 18 281 19 282
rect 17 281 18 282
rect 16 281 17 282
rect 15 281 16 282
rect 14 281 15 282
rect 13 281 14 282
rect 12 281 13 282
rect 11 281 12 282
rect 10 281 11 282
rect 9 281 10 282
rect 8 281 9 282
rect 7 281 8 282
rect 6 281 7 282
rect 5 281 6 282
rect 441 282 442 283
rect 440 282 441 283
rect 439 282 440 283
rect 438 282 439 283
rect 437 282 438 283
rect 436 282 437 283
rect 435 282 436 283
rect 434 282 435 283
rect 433 282 434 283
rect 432 282 433 283
rect 431 282 432 283
rect 430 282 431 283
rect 429 282 430 283
rect 428 282 429 283
rect 427 282 428 283
rect 426 282 427 283
rect 425 282 426 283
rect 424 282 425 283
rect 423 282 424 283
rect 422 282 423 283
rect 421 282 422 283
rect 420 282 421 283
rect 419 282 420 283
rect 418 282 419 283
rect 417 282 418 283
rect 416 282 417 283
rect 415 282 416 283
rect 414 282 415 283
rect 413 282 414 283
rect 412 282 413 283
rect 411 282 412 283
rect 410 282 411 283
rect 409 282 410 283
rect 408 282 409 283
rect 407 282 408 283
rect 406 282 407 283
rect 405 282 406 283
rect 404 282 405 283
rect 403 282 404 283
rect 402 282 403 283
rect 401 282 402 283
rect 400 282 401 283
rect 399 282 400 283
rect 398 282 399 283
rect 397 282 398 283
rect 291 282 292 283
rect 290 282 291 283
rect 289 282 290 283
rect 288 282 289 283
rect 287 282 288 283
rect 286 282 287 283
rect 285 282 286 283
rect 284 282 285 283
rect 283 282 284 283
rect 282 282 283 283
rect 281 282 282 283
rect 280 282 281 283
rect 279 282 280 283
rect 278 282 279 283
rect 277 282 278 283
rect 276 282 277 283
rect 275 282 276 283
rect 274 282 275 283
rect 273 282 274 283
rect 272 282 273 283
rect 271 282 272 283
rect 270 282 271 283
rect 269 282 270 283
rect 268 282 269 283
rect 267 282 268 283
rect 266 282 267 283
rect 265 282 266 283
rect 264 282 265 283
rect 263 282 264 283
rect 262 282 263 283
rect 261 282 262 283
rect 260 282 261 283
rect 259 282 260 283
rect 258 282 259 283
rect 257 282 258 283
rect 256 282 257 283
rect 255 282 256 283
rect 254 282 255 283
rect 253 282 254 283
rect 252 282 253 283
rect 251 282 252 283
rect 250 282 251 283
rect 249 282 250 283
rect 248 282 249 283
rect 247 282 248 283
rect 246 282 247 283
rect 245 282 246 283
rect 244 282 245 283
rect 243 282 244 283
rect 242 282 243 283
rect 241 282 242 283
rect 240 282 241 283
rect 239 282 240 283
rect 238 282 239 283
rect 237 282 238 283
rect 236 282 237 283
rect 235 282 236 283
rect 234 282 235 283
rect 233 282 234 283
rect 232 282 233 283
rect 231 282 232 283
rect 230 282 231 283
rect 229 282 230 283
rect 228 282 229 283
rect 227 282 228 283
rect 226 282 227 283
rect 225 282 226 283
rect 224 282 225 283
rect 223 282 224 283
rect 222 282 223 283
rect 200 282 201 283
rect 199 282 200 283
rect 198 282 199 283
rect 197 282 198 283
rect 196 282 197 283
rect 195 282 196 283
rect 194 282 195 283
rect 193 282 194 283
rect 192 282 193 283
rect 191 282 192 283
rect 190 282 191 283
rect 189 282 190 283
rect 188 282 189 283
rect 187 282 188 283
rect 186 282 187 283
rect 185 282 186 283
rect 184 282 185 283
rect 183 282 184 283
rect 182 282 183 283
rect 181 282 182 283
rect 180 282 181 283
rect 179 282 180 283
rect 178 282 179 283
rect 177 282 178 283
rect 176 282 177 283
rect 175 282 176 283
rect 174 282 175 283
rect 173 282 174 283
rect 172 282 173 283
rect 171 282 172 283
rect 170 282 171 283
rect 169 282 170 283
rect 168 282 169 283
rect 167 282 168 283
rect 166 282 167 283
rect 165 282 166 283
rect 164 282 165 283
rect 163 282 164 283
rect 162 282 163 283
rect 161 282 162 283
rect 160 282 161 283
rect 159 282 160 283
rect 158 282 159 283
rect 157 282 158 283
rect 156 282 157 283
rect 155 282 156 283
rect 154 282 155 283
rect 153 282 154 283
rect 152 282 153 283
rect 151 282 152 283
rect 150 282 151 283
rect 149 282 150 283
rect 148 282 149 283
rect 147 282 148 283
rect 146 282 147 283
rect 145 282 146 283
rect 144 282 145 283
rect 143 282 144 283
rect 142 282 143 283
rect 141 282 142 283
rect 140 282 141 283
rect 139 282 140 283
rect 138 282 139 283
rect 137 282 138 283
rect 136 282 137 283
rect 135 282 136 283
rect 134 282 135 283
rect 133 282 134 283
rect 132 282 133 283
rect 131 282 132 283
rect 116 282 117 283
rect 115 282 116 283
rect 114 282 115 283
rect 113 282 114 283
rect 112 282 113 283
rect 111 282 112 283
rect 110 282 111 283
rect 109 282 110 283
rect 108 282 109 283
rect 107 282 108 283
rect 106 282 107 283
rect 105 282 106 283
rect 104 282 105 283
rect 103 282 104 283
rect 102 282 103 283
rect 101 282 102 283
rect 100 282 101 283
rect 99 282 100 283
rect 98 282 99 283
rect 97 282 98 283
rect 96 282 97 283
rect 95 282 96 283
rect 94 282 95 283
rect 93 282 94 283
rect 92 282 93 283
rect 91 282 92 283
rect 90 282 91 283
rect 89 282 90 283
rect 88 282 89 283
rect 87 282 88 283
rect 86 282 87 283
rect 85 282 86 283
rect 84 282 85 283
rect 83 282 84 283
rect 82 282 83 283
rect 66 282 67 283
rect 65 282 66 283
rect 64 282 65 283
rect 63 282 64 283
rect 62 282 63 283
rect 61 282 62 283
rect 60 282 61 283
rect 59 282 60 283
rect 58 282 59 283
rect 57 282 58 283
rect 56 282 57 283
rect 55 282 56 283
rect 54 282 55 283
rect 53 282 54 283
rect 52 282 53 283
rect 51 282 52 283
rect 50 282 51 283
rect 49 282 50 283
rect 48 282 49 283
rect 47 282 48 283
rect 46 282 47 283
rect 45 282 46 283
rect 44 282 45 283
rect 43 282 44 283
rect 42 282 43 283
rect 41 282 42 283
rect 40 282 41 283
rect 30 282 31 283
rect 29 282 30 283
rect 28 282 29 283
rect 27 282 28 283
rect 26 282 27 283
rect 25 282 26 283
rect 24 282 25 283
rect 23 282 24 283
rect 22 282 23 283
rect 21 282 22 283
rect 20 282 21 283
rect 19 282 20 283
rect 18 282 19 283
rect 17 282 18 283
rect 16 282 17 283
rect 15 282 16 283
rect 14 282 15 283
rect 13 282 14 283
rect 12 282 13 283
rect 11 282 12 283
rect 10 282 11 283
rect 9 282 10 283
rect 8 282 9 283
rect 7 282 8 283
rect 6 282 7 283
rect 5 282 6 283
rect 441 283 442 284
rect 440 283 441 284
rect 439 283 440 284
rect 438 283 439 284
rect 437 283 438 284
rect 436 283 437 284
rect 435 283 436 284
rect 434 283 435 284
rect 433 283 434 284
rect 432 283 433 284
rect 431 283 432 284
rect 430 283 431 284
rect 429 283 430 284
rect 428 283 429 284
rect 427 283 428 284
rect 426 283 427 284
rect 425 283 426 284
rect 424 283 425 284
rect 423 283 424 284
rect 422 283 423 284
rect 421 283 422 284
rect 420 283 421 284
rect 419 283 420 284
rect 418 283 419 284
rect 417 283 418 284
rect 416 283 417 284
rect 415 283 416 284
rect 414 283 415 284
rect 413 283 414 284
rect 412 283 413 284
rect 411 283 412 284
rect 410 283 411 284
rect 409 283 410 284
rect 408 283 409 284
rect 407 283 408 284
rect 406 283 407 284
rect 405 283 406 284
rect 404 283 405 284
rect 403 283 404 284
rect 402 283 403 284
rect 401 283 402 284
rect 400 283 401 284
rect 399 283 400 284
rect 398 283 399 284
rect 397 283 398 284
rect 290 283 291 284
rect 289 283 290 284
rect 288 283 289 284
rect 287 283 288 284
rect 286 283 287 284
rect 285 283 286 284
rect 284 283 285 284
rect 283 283 284 284
rect 282 283 283 284
rect 281 283 282 284
rect 280 283 281 284
rect 279 283 280 284
rect 278 283 279 284
rect 277 283 278 284
rect 276 283 277 284
rect 275 283 276 284
rect 274 283 275 284
rect 273 283 274 284
rect 272 283 273 284
rect 271 283 272 284
rect 270 283 271 284
rect 269 283 270 284
rect 268 283 269 284
rect 267 283 268 284
rect 266 283 267 284
rect 265 283 266 284
rect 264 283 265 284
rect 263 283 264 284
rect 262 283 263 284
rect 261 283 262 284
rect 260 283 261 284
rect 259 283 260 284
rect 258 283 259 284
rect 257 283 258 284
rect 256 283 257 284
rect 255 283 256 284
rect 254 283 255 284
rect 253 283 254 284
rect 252 283 253 284
rect 251 283 252 284
rect 250 283 251 284
rect 249 283 250 284
rect 248 283 249 284
rect 247 283 248 284
rect 246 283 247 284
rect 245 283 246 284
rect 244 283 245 284
rect 243 283 244 284
rect 242 283 243 284
rect 241 283 242 284
rect 240 283 241 284
rect 239 283 240 284
rect 238 283 239 284
rect 237 283 238 284
rect 236 283 237 284
rect 235 283 236 284
rect 234 283 235 284
rect 233 283 234 284
rect 232 283 233 284
rect 231 283 232 284
rect 230 283 231 284
rect 229 283 230 284
rect 228 283 229 284
rect 227 283 228 284
rect 226 283 227 284
rect 225 283 226 284
rect 224 283 225 284
rect 223 283 224 284
rect 222 283 223 284
rect 200 283 201 284
rect 199 283 200 284
rect 198 283 199 284
rect 197 283 198 284
rect 196 283 197 284
rect 195 283 196 284
rect 194 283 195 284
rect 193 283 194 284
rect 192 283 193 284
rect 191 283 192 284
rect 190 283 191 284
rect 189 283 190 284
rect 188 283 189 284
rect 187 283 188 284
rect 186 283 187 284
rect 185 283 186 284
rect 184 283 185 284
rect 183 283 184 284
rect 182 283 183 284
rect 181 283 182 284
rect 180 283 181 284
rect 179 283 180 284
rect 178 283 179 284
rect 177 283 178 284
rect 176 283 177 284
rect 175 283 176 284
rect 174 283 175 284
rect 173 283 174 284
rect 172 283 173 284
rect 171 283 172 284
rect 170 283 171 284
rect 169 283 170 284
rect 168 283 169 284
rect 167 283 168 284
rect 166 283 167 284
rect 165 283 166 284
rect 164 283 165 284
rect 163 283 164 284
rect 162 283 163 284
rect 161 283 162 284
rect 160 283 161 284
rect 159 283 160 284
rect 158 283 159 284
rect 157 283 158 284
rect 156 283 157 284
rect 155 283 156 284
rect 154 283 155 284
rect 153 283 154 284
rect 152 283 153 284
rect 151 283 152 284
rect 150 283 151 284
rect 149 283 150 284
rect 148 283 149 284
rect 147 283 148 284
rect 146 283 147 284
rect 145 283 146 284
rect 144 283 145 284
rect 143 283 144 284
rect 142 283 143 284
rect 141 283 142 284
rect 140 283 141 284
rect 139 283 140 284
rect 138 283 139 284
rect 137 283 138 284
rect 136 283 137 284
rect 135 283 136 284
rect 134 283 135 284
rect 133 283 134 284
rect 132 283 133 284
rect 116 283 117 284
rect 115 283 116 284
rect 114 283 115 284
rect 113 283 114 284
rect 112 283 113 284
rect 111 283 112 284
rect 110 283 111 284
rect 109 283 110 284
rect 108 283 109 284
rect 107 283 108 284
rect 106 283 107 284
rect 105 283 106 284
rect 104 283 105 284
rect 103 283 104 284
rect 102 283 103 284
rect 101 283 102 284
rect 100 283 101 284
rect 99 283 100 284
rect 98 283 99 284
rect 97 283 98 284
rect 96 283 97 284
rect 95 283 96 284
rect 94 283 95 284
rect 93 283 94 284
rect 92 283 93 284
rect 91 283 92 284
rect 90 283 91 284
rect 89 283 90 284
rect 88 283 89 284
rect 87 283 88 284
rect 86 283 87 284
rect 85 283 86 284
rect 84 283 85 284
rect 83 283 84 284
rect 82 283 83 284
rect 66 283 67 284
rect 65 283 66 284
rect 64 283 65 284
rect 63 283 64 284
rect 62 283 63 284
rect 61 283 62 284
rect 60 283 61 284
rect 59 283 60 284
rect 58 283 59 284
rect 57 283 58 284
rect 56 283 57 284
rect 55 283 56 284
rect 54 283 55 284
rect 53 283 54 284
rect 52 283 53 284
rect 51 283 52 284
rect 50 283 51 284
rect 49 283 50 284
rect 48 283 49 284
rect 47 283 48 284
rect 46 283 47 284
rect 45 283 46 284
rect 44 283 45 284
rect 43 283 44 284
rect 42 283 43 284
rect 41 283 42 284
rect 40 283 41 284
rect 30 283 31 284
rect 29 283 30 284
rect 28 283 29 284
rect 27 283 28 284
rect 26 283 27 284
rect 25 283 26 284
rect 24 283 25 284
rect 23 283 24 284
rect 22 283 23 284
rect 21 283 22 284
rect 20 283 21 284
rect 19 283 20 284
rect 18 283 19 284
rect 17 283 18 284
rect 16 283 17 284
rect 15 283 16 284
rect 14 283 15 284
rect 13 283 14 284
rect 12 283 13 284
rect 11 283 12 284
rect 10 283 11 284
rect 9 283 10 284
rect 8 283 9 284
rect 7 283 8 284
rect 6 283 7 284
rect 5 283 6 284
rect 441 284 442 285
rect 440 284 441 285
rect 439 284 440 285
rect 438 284 439 285
rect 437 284 438 285
rect 436 284 437 285
rect 435 284 436 285
rect 434 284 435 285
rect 433 284 434 285
rect 432 284 433 285
rect 431 284 432 285
rect 430 284 431 285
rect 429 284 430 285
rect 428 284 429 285
rect 427 284 428 285
rect 426 284 427 285
rect 425 284 426 285
rect 424 284 425 285
rect 423 284 424 285
rect 422 284 423 285
rect 421 284 422 285
rect 420 284 421 285
rect 419 284 420 285
rect 418 284 419 285
rect 417 284 418 285
rect 416 284 417 285
rect 415 284 416 285
rect 414 284 415 285
rect 413 284 414 285
rect 412 284 413 285
rect 411 284 412 285
rect 410 284 411 285
rect 409 284 410 285
rect 408 284 409 285
rect 407 284 408 285
rect 406 284 407 285
rect 405 284 406 285
rect 404 284 405 285
rect 403 284 404 285
rect 402 284 403 285
rect 401 284 402 285
rect 400 284 401 285
rect 399 284 400 285
rect 398 284 399 285
rect 397 284 398 285
rect 289 284 290 285
rect 288 284 289 285
rect 287 284 288 285
rect 286 284 287 285
rect 285 284 286 285
rect 284 284 285 285
rect 283 284 284 285
rect 282 284 283 285
rect 281 284 282 285
rect 280 284 281 285
rect 279 284 280 285
rect 278 284 279 285
rect 277 284 278 285
rect 276 284 277 285
rect 275 284 276 285
rect 274 284 275 285
rect 273 284 274 285
rect 272 284 273 285
rect 271 284 272 285
rect 270 284 271 285
rect 269 284 270 285
rect 268 284 269 285
rect 267 284 268 285
rect 266 284 267 285
rect 265 284 266 285
rect 264 284 265 285
rect 263 284 264 285
rect 262 284 263 285
rect 261 284 262 285
rect 260 284 261 285
rect 259 284 260 285
rect 258 284 259 285
rect 257 284 258 285
rect 256 284 257 285
rect 255 284 256 285
rect 254 284 255 285
rect 253 284 254 285
rect 252 284 253 285
rect 251 284 252 285
rect 250 284 251 285
rect 249 284 250 285
rect 248 284 249 285
rect 247 284 248 285
rect 246 284 247 285
rect 245 284 246 285
rect 244 284 245 285
rect 243 284 244 285
rect 242 284 243 285
rect 241 284 242 285
rect 240 284 241 285
rect 239 284 240 285
rect 238 284 239 285
rect 237 284 238 285
rect 236 284 237 285
rect 235 284 236 285
rect 234 284 235 285
rect 233 284 234 285
rect 232 284 233 285
rect 231 284 232 285
rect 230 284 231 285
rect 229 284 230 285
rect 228 284 229 285
rect 227 284 228 285
rect 226 284 227 285
rect 225 284 226 285
rect 224 284 225 285
rect 223 284 224 285
rect 222 284 223 285
rect 221 284 222 285
rect 199 284 200 285
rect 198 284 199 285
rect 197 284 198 285
rect 196 284 197 285
rect 195 284 196 285
rect 194 284 195 285
rect 193 284 194 285
rect 192 284 193 285
rect 191 284 192 285
rect 190 284 191 285
rect 189 284 190 285
rect 188 284 189 285
rect 187 284 188 285
rect 186 284 187 285
rect 185 284 186 285
rect 184 284 185 285
rect 183 284 184 285
rect 182 284 183 285
rect 181 284 182 285
rect 180 284 181 285
rect 179 284 180 285
rect 178 284 179 285
rect 177 284 178 285
rect 176 284 177 285
rect 175 284 176 285
rect 174 284 175 285
rect 173 284 174 285
rect 172 284 173 285
rect 171 284 172 285
rect 170 284 171 285
rect 169 284 170 285
rect 168 284 169 285
rect 167 284 168 285
rect 166 284 167 285
rect 165 284 166 285
rect 164 284 165 285
rect 163 284 164 285
rect 162 284 163 285
rect 161 284 162 285
rect 160 284 161 285
rect 159 284 160 285
rect 158 284 159 285
rect 157 284 158 285
rect 156 284 157 285
rect 155 284 156 285
rect 154 284 155 285
rect 153 284 154 285
rect 152 284 153 285
rect 151 284 152 285
rect 150 284 151 285
rect 149 284 150 285
rect 148 284 149 285
rect 147 284 148 285
rect 146 284 147 285
rect 145 284 146 285
rect 144 284 145 285
rect 143 284 144 285
rect 142 284 143 285
rect 141 284 142 285
rect 140 284 141 285
rect 139 284 140 285
rect 138 284 139 285
rect 137 284 138 285
rect 136 284 137 285
rect 135 284 136 285
rect 134 284 135 285
rect 133 284 134 285
rect 132 284 133 285
rect 117 284 118 285
rect 116 284 117 285
rect 115 284 116 285
rect 114 284 115 285
rect 113 284 114 285
rect 112 284 113 285
rect 111 284 112 285
rect 110 284 111 285
rect 109 284 110 285
rect 108 284 109 285
rect 107 284 108 285
rect 106 284 107 285
rect 105 284 106 285
rect 104 284 105 285
rect 103 284 104 285
rect 102 284 103 285
rect 101 284 102 285
rect 100 284 101 285
rect 99 284 100 285
rect 98 284 99 285
rect 97 284 98 285
rect 96 284 97 285
rect 95 284 96 285
rect 94 284 95 285
rect 93 284 94 285
rect 92 284 93 285
rect 91 284 92 285
rect 90 284 91 285
rect 89 284 90 285
rect 88 284 89 285
rect 87 284 88 285
rect 86 284 87 285
rect 85 284 86 285
rect 84 284 85 285
rect 83 284 84 285
rect 66 284 67 285
rect 65 284 66 285
rect 64 284 65 285
rect 63 284 64 285
rect 62 284 63 285
rect 61 284 62 285
rect 60 284 61 285
rect 59 284 60 285
rect 58 284 59 285
rect 57 284 58 285
rect 56 284 57 285
rect 55 284 56 285
rect 54 284 55 285
rect 53 284 54 285
rect 52 284 53 285
rect 51 284 52 285
rect 50 284 51 285
rect 49 284 50 285
rect 48 284 49 285
rect 47 284 48 285
rect 46 284 47 285
rect 45 284 46 285
rect 44 284 45 285
rect 43 284 44 285
rect 42 284 43 285
rect 41 284 42 285
rect 40 284 41 285
rect 30 284 31 285
rect 29 284 30 285
rect 28 284 29 285
rect 27 284 28 285
rect 26 284 27 285
rect 25 284 26 285
rect 24 284 25 285
rect 23 284 24 285
rect 22 284 23 285
rect 21 284 22 285
rect 20 284 21 285
rect 19 284 20 285
rect 18 284 19 285
rect 17 284 18 285
rect 16 284 17 285
rect 15 284 16 285
rect 14 284 15 285
rect 13 284 14 285
rect 12 284 13 285
rect 11 284 12 285
rect 10 284 11 285
rect 9 284 10 285
rect 8 284 9 285
rect 7 284 8 285
rect 6 284 7 285
rect 5 284 6 285
rect 441 285 442 286
rect 440 285 441 286
rect 439 285 440 286
rect 438 285 439 286
rect 437 285 438 286
rect 436 285 437 286
rect 435 285 436 286
rect 434 285 435 286
rect 433 285 434 286
rect 432 285 433 286
rect 431 285 432 286
rect 430 285 431 286
rect 429 285 430 286
rect 428 285 429 286
rect 427 285 428 286
rect 426 285 427 286
rect 425 285 426 286
rect 424 285 425 286
rect 423 285 424 286
rect 422 285 423 286
rect 421 285 422 286
rect 420 285 421 286
rect 419 285 420 286
rect 418 285 419 286
rect 417 285 418 286
rect 416 285 417 286
rect 415 285 416 286
rect 414 285 415 286
rect 413 285 414 286
rect 412 285 413 286
rect 411 285 412 286
rect 410 285 411 286
rect 409 285 410 286
rect 408 285 409 286
rect 407 285 408 286
rect 406 285 407 286
rect 405 285 406 286
rect 404 285 405 286
rect 403 285 404 286
rect 402 285 403 286
rect 401 285 402 286
rect 400 285 401 286
rect 399 285 400 286
rect 398 285 399 286
rect 397 285 398 286
rect 288 285 289 286
rect 287 285 288 286
rect 286 285 287 286
rect 285 285 286 286
rect 284 285 285 286
rect 283 285 284 286
rect 282 285 283 286
rect 281 285 282 286
rect 280 285 281 286
rect 279 285 280 286
rect 278 285 279 286
rect 277 285 278 286
rect 276 285 277 286
rect 275 285 276 286
rect 274 285 275 286
rect 273 285 274 286
rect 272 285 273 286
rect 271 285 272 286
rect 270 285 271 286
rect 269 285 270 286
rect 268 285 269 286
rect 267 285 268 286
rect 266 285 267 286
rect 265 285 266 286
rect 264 285 265 286
rect 263 285 264 286
rect 262 285 263 286
rect 261 285 262 286
rect 260 285 261 286
rect 259 285 260 286
rect 258 285 259 286
rect 257 285 258 286
rect 256 285 257 286
rect 255 285 256 286
rect 254 285 255 286
rect 253 285 254 286
rect 252 285 253 286
rect 251 285 252 286
rect 250 285 251 286
rect 249 285 250 286
rect 248 285 249 286
rect 247 285 248 286
rect 246 285 247 286
rect 245 285 246 286
rect 244 285 245 286
rect 243 285 244 286
rect 242 285 243 286
rect 241 285 242 286
rect 240 285 241 286
rect 239 285 240 286
rect 238 285 239 286
rect 237 285 238 286
rect 236 285 237 286
rect 235 285 236 286
rect 234 285 235 286
rect 233 285 234 286
rect 232 285 233 286
rect 231 285 232 286
rect 230 285 231 286
rect 229 285 230 286
rect 228 285 229 286
rect 227 285 228 286
rect 226 285 227 286
rect 225 285 226 286
rect 224 285 225 286
rect 223 285 224 286
rect 222 285 223 286
rect 221 285 222 286
rect 198 285 199 286
rect 197 285 198 286
rect 196 285 197 286
rect 195 285 196 286
rect 194 285 195 286
rect 193 285 194 286
rect 192 285 193 286
rect 191 285 192 286
rect 190 285 191 286
rect 189 285 190 286
rect 188 285 189 286
rect 187 285 188 286
rect 186 285 187 286
rect 185 285 186 286
rect 184 285 185 286
rect 183 285 184 286
rect 182 285 183 286
rect 181 285 182 286
rect 180 285 181 286
rect 179 285 180 286
rect 178 285 179 286
rect 177 285 178 286
rect 176 285 177 286
rect 175 285 176 286
rect 174 285 175 286
rect 173 285 174 286
rect 172 285 173 286
rect 171 285 172 286
rect 170 285 171 286
rect 169 285 170 286
rect 168 285 169 286
rect 167 285 168 286
rect 166 285 167 286
rect 165 285 166 286
rect 164 285 165 286
rect 163 285 164 286
rect 162 285 163 286
rect 161 285 162 286
rect 160 285 161 286
rect 159 285 160 286
rect 158 285 159 286
rect 157 285 158 286
rect 156 285 157 286
rect 155 285 156 286
rect 154 285 155 286
rect 153 285 154 286
rect 152 285 153 286
rect 151 285 152 286
rect 150 285 151 286
rect 149 285 150 286
rect 148 285 149 286
rect 147 285 148 286
rect 146 285 147 286
rect 145 285 146 286
rect 144 285 145 286
rect 143 285 144 286
rect 142 285 143 286
rect 141 285 142 286
rect 140 285 141 286
rect 139 285 140 286
rect 138 285 139 286
rect 137 285 138 286
rect 136 285 137 286
rect 135 285 136 286
rect 134 285 135 286
rect 133 285 134 286
rect 117 285 118 286
rect 116 285 117 286
rect 115 285 116 286
rect 114 285 115 286
rect 113 285 114 286
rect 112 285 113 286
rect 111 285 112 286
rect 110 285 111 286
rect 109 285 110 286
rect 108 285 109 286
rect 107 285 108 286
rect 106 285 107 286
rect 105 285 106 286
rect 104 285 105 286
rect 103 285 104 286
rect 102 285 103 286
rect 101 285 102 286
rect 100 285 101 286
rect 99 285 100 286
rect 98 285 99 286
rect 97 285 98 286
rect 96 285 97 286
rect 95 285 96 286
rect 94 285 95 286
rect 93 285 94 286
rect 92 285 93 286
rect 91 285 92 286
rect 90 285 91 286
rect 89 285 90 286
rect 88 285 89 286
rect 87 285 88 286
rect 86 285 87 286
rect 85 285 86 286
rect 84 285 85 286
rect 83 285 84 286
rect 67 285 68 286
rect 66 285 67 286
rect 65 285 66 286
rect 64 285 65 286
rect 63 285 64 286
rect 62 285 63 286
rect 61 285 62 286
rect 60 285 61 286
rect 59 285 60 286
rect 58 285 59 286
rect 57 285 58 286
rect 56 285 57 286
rect 55 285 56 286
rect 54 285 55 286
rect 53 285 54 286
rect 52 285 53 286
rect 51 285 52 286
rect 50 285 51 286
rect 49 285 50 286
rect 48 285 49 286
rect 47 285 48 286
rect 46 285 47 286
rect 45 285 46 286
rect 44 285 45 286
rect 43 285 44 286
rect 42 285 43 286
rect 41 285 42 286
rect 40 285 41 286
rect 30 285 31 286
rect 29 285 30 286
rect 28 285 29 286
rect 27 285 28 286
rect 26 285 27 286
rect 25 285 26 286
rect 24 285 25 286
rect 23 285 24 286
rect 22 285 23 286
rect 21 285 22 286
rect 20 285 21 286
rect 19 285 20 286
rect 18 285 19 286
rect 17 285 18 286
rect 16 285 17 286
rect 15 285 16 286
rect 14 285 15 286
rect 13 285 14 286
rect 12 285 13 286
rect 11 285 12 286
rect 10 285 11 286
rect 9 285 10 286
rect 8 285 9 286
rect 7 285 8 286
rect 6 285 7 286
rect 5 285 6 286
rect 466 286 467 287
rect 441 286 442 287
rect 440 286 441 287
rect 439 286 440 287
rect 438 286 439 287
rect 437 286 438 287
rect 436 286 437 287
rect 435 286 436 287
rect 434 286 435 287
rect 433 286 434 287
rect 432 286 433 287
rect 431 286 432 287
rect 430 286 431 287
rect 429 286 430 287
rect 428 286 429 287
rect 427 286 428 287
rect 426 286 427 287
rect 425 286 426 287
rect 424 286 425 287
rect 423 286 424 287
rect 422 286 423 287
rect 421 286 422 287
rect 420 286 421 287
rect 419 286 420 287
rect 418 286 419 287
rect 417 286 418 287
rect 416 286 417 287
rect 415 286 416 287
rect 414 286 415 287
rect 413 286 414 287
rect 412 286 413 287
rect 411 286 412 287
rect 410 286 411 287
rect 409 286 410 287
rect 408 286 409 287
rect 407 286 408 287
rect 406 286 407 287
rect 405 286 406 287
rect 404 286 405 287
rect 403 286 404 287
rect 402 286 403 287
rect 401 286 402 287
rect 400 286 401 287
rect 399 286 400 287
rect 398 286 399 287
rect 397 286 398 287
rect 287 286 288 287
rect 286 286 287 287
rect 285 286 286 287
rect 284 286 285 287
rect 283 286 284 287
rect 282 286 283 287
rect 281 286 282 287
rect 280 286 281 287
rect 279 286 280 287
rect 278 286 279 287
rect 277 286 278 287
rect 276 286 277 287
rect 275 286 276 287
rect 274 286 275 287
rect 273 286 274 287
rect 272 286 273 287
rect 271 286 272 287
rect 270 286 271 287
rect 269 286 270 287
rect 268 286 269 287
rect 267 286 268 287
rect 266 286 267 287
rect 265 286 266 287
rect 264 286 265 287
rect 263 286 264 287
rect 262 286 263 287
rect 261 286 262 287
rect 260 286 261 287
rect 259 286 260 287
rect 258 286 259 287
rect 257 286 258 287
rect 256 286 257 287
rect 255 286 256 287
rect 254 286 255 287
rect 253 286 254 287
rect 252 286 253 287
rect 251 286 252 287
rect 250 286 251 287
rect 249 286 250 287
rect 248 286 249 287
rect 247 286 248 287
rect 246 286 247 287
rect 245 286 246 287
rect 244 286 245 287
rect 243 286 244 287
rect 242 286 243 287
rect 241 286 242 287
rect 240 286 241 287
rect 239 286 240 287
rect 238 286 239 287
rect 237 286 238 287
rect 236 286 237 287
rect 235 286 236 287
rect 234 286 235 287
rect 233 286 234 287
rect 232 286 233 287
rect 231 286 232 287
rect 230 286 231 287
rect 229 286 230 287
rect 228 286 229 287
rect 227 286 228 287
rect 226 286 227 287
rect 225 286 226 287
rect 224 286 225 287
rect 223 286 224 287
rect 222 286 223 287
rect 221 286 222 287
rect 220 286 221 287
rect 198 286 199 287
rect 197 286 198 287
rect 196 286 197 287
rect 195 286 196 287
rect 194 286 195 287
rect 193 286 194 287
rect 192 286 193 287
rect 191 286 192 287
rect 190 286 191 287
rect 189 286 190 287
rect 188 286 189 287
rect 187 286 188 287
rect 186 286 187 287
rect 185 286 186 287
rect 184 286 185 287
rect 183 286 184 287
rect 182 286 183 287
rect 181 286 182 287
rect 180 286 181 287
rect 179 286 180 287
rect 178 286 179 287
rect 177 286 178 287
rect 176 286 177 287
rect 175 286 176 287
rect 174 286 175 287
rect 173 286 174 287
rect 172 286 173 287
rect 171 286 172 287
rect 170 286 171 287
rect 169 286 170 287
rect 168 286 169 287
rect 167 286 168 287
rect 166 286 167 287
rect 165 286 166 287
rect 164 286 165 287
rect 163 286 164 287
rect 162 286 163 287
rect 161 286 162 287
rect 160 286 161 287
rect 159 286 160 287
rect 158 286 159 287
rect 157 286 158 287
rect 156 286 157 287
rect 155 286 156 287
rect 154 286 155 287
rect 153 286 154 287
rect 152 286 153 287
rect 151 286 152 287
rect 150 286 151 287
rect 149 286 150 287
rect 148 286 149 287
rect 147 286 148 287
rect 146 286 147 287
rect 145 286 146 287
rect 144 286 145 287
rect 143 286 144 287
rect 142 286 143 287
rect 141 286 142 287
rect 140 286 141 287
rect 139 286 140 287
rect 138 286 139 287
rect 137 286 138 287
rect 136 286 137 287
rect 135 286 136 287
rect 134 286 135 287
rect 133 286 134 287
rect 117 286 118 287
rect 116 286 117 287
rect 115 286 116 287
rect 114 286 115 287
rect 113 286 114 287
rect 112 286 113 287
rect 111 286 112 287
rect 110 286 111 287
rect 109 286 110 287
rect 108 286 109 287
rect 107 286 108 287
rect 106 286 107 287
rect 105 286 106 287
rect 104 286 105 287
rect 103 286 104 287
rect 102 286 103 287
rect 101 286 102 287
rect 100 286 101 287
rect 99 286 100 287
rect 98 286 99 287
rect 97 286 98 287
rect 96 286 97 287
rect 95 286 96 287
rect 94 286 95 287
rect 93 286 94 287
rect 92 286 93 287
rect 91 286 92 287
rect 90 286 91 287
rect 89 286 90 287
rect 88 286 89 287
rect 87 286 88 287
rect 86 286 87 287
rect 85 286 86 287
rect 84 286 85 287
rect 83 286 84 287
rect 67 286 68 287
rect 66 286 67 287
rect 65 286 66 287
rect 64 286 65 287
rect 63 286 64 287
rect 62 286 63 287
rect 61 286 62 287
rect 60 286 61 287
rect 59 286 60 287
rect 58 286 59 287
rect 57 286 58 287
rect 56 286 57 287
rect 55 286 56 287
rect 54 286 55 287
rect 53 286 54 287
rect 52 286 53 287
rect 51 286 52 287
rect 50 286 51 287
rect 49 286 50 287
rect 48 286 49 287
rect 47 286 48 287
rect 46 286 47 287
rect 45 286 46 287
rect 44 286 45 287
rect 43 286 44 287
rect 42 286 43 287
rect 41 286 42 287
rect 40 286 41 287
rect 30 286 31 287
rect 29 286 30 287
rect 28 286 29 287
rect 27 286 28 287
rect 26 286 27 287
rect 25 286 26 287
rect 24 286 25 287
rect 23 286 24 287
rect 22 286 23 287
rect 21 286 22 287
rect 20 286 21 287
rect 19 286 20 287
rect 18 286 19 287
rect 17 286 18 287
rect 16 286 17 287
rect 15 286 16 287
rect 14 286 15 287
rect 13 286 14 287
rect 12 286 13 287
rect 11 286 12 287
rect 10 286 11 287
rect 9 286 10 287
rect 8 286 9 287
rect 7 286 8 287
rect 6 286 7 287
rect 5 286 6 287
rect 467 287 468 288
rect 466 287 467 288
rect 465 287 466 288
rect 464 287 465 288
rect 463 287 464 288
rect 462 287 463 288
rect 461 287 462 288
rect 441 287 442 288
rect 440 287 441 288
rect 439 287 440 288
rect 438 287 439 288
rect 437 287 438 288
rect 436 287 437 288
rect 435 287 436 288
rect 434 287 435 288
rect 433 287 434 288
rect 432 287 433 288
rect 431 287 432 288
rect 430 287 431 288
rect 429 287 430 288
rect 428 287 429 288
rect 427 287 428 288
rect 426 287 427 288
rect 425 287 426 288
rect 424 287 425 288
rect 423 287 424 288
rect 422 287 423 288
rect 421 287 422 288
rect 420 287 421 288
rect 419 287 420 288
rect 418 287 419 288
rect 417 287 418 288
rect 416 287 417 288
rect 415 287 416 288
rect 414 287 415 288
rect 413 287 414 288
rect 412 287 413 288
rect 411 287 412 288
rect 410 287 411 288
rect 409 287 410 288
rect 408 287 409 288
rect 407 287 408 288
rect 406 287 407 288
rect 405 287 406 288
rect 404 287 405 288
rect 403 287 404 288
rect 402 287 403 288
rect 401 287 402 288
rect 400 287 401 288
rect 399 287 400 288
rect 398 287 399 288
rect 397 287 398 288
rect 286 287 287 288
rect 285 287 286 288
rect 284 287 285 288
rect 283 287 284 288
rect 282 287 283 288
rect 281 287 282 288
rect 280 287 281 288
rect 279 287 280 288
rect 278 287 279 288
rect 277 287 278 288
rect 276 287 277 288
rect 275 287 276 288
rect 274 287 275 288
rect 273 287 274 288
rect 272 287 273 288
rect 271 287 272 288
rect 270 287 271 288
rect 269 287 270 288
rect 268 287 269 288
rect 267 287 268 288
rect 266 287 267 288
rect 265 287 266 288
rect 264 287 265 288
rect 263 287 264 288
rect 262 287 263 288
rect 261 287 262 288
rect 260 287 261 288
rect 259 287 260 288
rect 258 287 259 288
rect 257 287 258 288
rect 256 287 257 288
rect 255 287 256 288
rect 254 287 255 288
rect 253 287 254 288
rect 252 287 253 288
rect 251 287 252 288
rect 250 287 251 288
rect 249 287 250 288
rect 248 287 249 288
rect 247 287 248 288
rect 246 287 247 288
rect 245 287 246 288
rect 244 287 245 288
rect 243 287 244 288
rect 242 287 243 288
rect 241 287 242 288
rect 240 287 241 288
rect 239 287 240 288
rect 238 287 239 288
rect 237 287 238 288
rect 236 287 237 288
rect 235 287 236 288
rect 234 287 235 288
rect 233 287 234 288
rect 232 287 233 288
rect 231 287 232 288
rect 230 287 231 288
rect 229 287 230 288
rect 228 287 229 288
rect 227 287 228 288
rect 226 287 227 288
rect 225 287 226 288
rect 224 287 225 288
rect 223 287 224 288
rect 222 287 223 288
rect 221 287 222 288
rect 220 287 221 288
rect 219 287 220 288
rect 197 287 198 288
rect 196 287 197 288
rect 195 287 196 288
rect 194 287 195 288
rect 193 287 194 288
rect 192 287 193 288
rect 191 287 192 288
rect 190 287 191 288
rect 189 287 190 288
rect 188 287 189 288
rect 187 287 188 288
rect 186 287 187 288
rect 185 287 186 288
rect 184 287 185 288
rect 183 287 184 288
rect 182 287 183 288
rect 181 287 182 288
rect 180 287 181 288
rect 179 287 180 288
rect 178 287 179 288
rect 177 287 178 288
rect 176 287 177 288
rect 175 287 176 288
rect 174 287 175 288
rect 173 287 174 288
rect 172 287 173 288
rect 171 287 172 288
rect 170 287 171 288
rect 169 287 170 288
rect 168 287 169 288
rect 167 287 168 288
rect 166 287 167 288
rect 165 287 166 288
rect 164 287 165 288
rect 163 287 164 288
rect 162 287 163 288
rect 161 287 162 288
rect 160 287 161 288
rect 159 287 160 288
rect 158 287 159 288
rect 157 287 158 288
rect 156 287 157 288
rect 155 287 156 288
rect 154 287 155 288
rect 153 287 154 288
rect 152 287 153 288
rect 151 287 152 288
rect 150 287 151 288
rect 149 287 150 288
rect 148 287 149 288
rect 147 287 148 288
rect 146 287 147 288
rect 145 287 146 288
rect 144 287 145 288
rect 143 287 144 288
rect 142 287 143 288
rect 141 287 142 288
rect 140 287 141 288
rect 139 287 140 288
rect 138 287 139 288
rect 137 287 138 288
rect 136 287 137 288
rect 135 287 136 288
rect 134 287 135 288
rect 118 287 119 288
rect 117 287 118 288
rect 116 287 117 288
rect 115 287 116 288
rect 114 287 115 288
rect 113 287 114 288
rect 112 287 113 288
rect 111 287 112 288
rect 110 287 111 288
rect 109 287 110 288
rect 108 287 109 288
rect 107 287 108 288
rect 106 287 107 288
rect 105 287 106 288
rect 104 287 105 288
rect 103 287 104 288
rect 102 287 103 288
rect 101 287 102 288
rect 100 287 101 288
rect 99 287 100 288
rect 98 287 99 288
rect 97 287 98 288
rect 96 287 97 288
rect 95 287 96 288
rect 94 287 95 288
rect 93 287 94 288
rect 92 287 93 288
rect 91 287 92 288
rect 90 287 91 288
rect 89 287 90 288
rect 88 287 89 288
rect 87 287 88 288
rect 86 287 87 288
rect 85 287 86 288
rect 84 287 85 288
rect 68 287 69 288
rect 67 287 68 288
rect 66 287 67 288
rect 65 287 66 288
rect 64 287 65 288
rect 63 287 64 288
rect 62 287 63 288
rect 61 287 62 288
rect 60 287 61 288
rect 59 287 60 288
rect 58 287 59 288
rect 57 287 58 288
rect 56 287 57 288
rect 55 287 56 288
rect 54 287 55 288
rect 53 287 54 288
rect 52 287 53 288
rect 51 287 52 288
rect 50 287 51 288
rect 49 287 50 288
rect 48 287 49 288
rect 47 287 48 288
rect 46 287 47 288
rect 45 287 46 288
rect 44 287 45 288
rect 43 287 44 288
rect 42 287 43 288
rect 41 287 42 288
rect 40 287 41 288
rect 30 287 31 288
rect 29 287 30 288
rect 28 287 29 288
rect 27 287 28 288
rect 26 287 27 288
rect 25 287 26 288
rect 24 287 25 288
rect 23 287 24 288
rect 22 287 23 288
rect 21 287 22 288
rect 20 287 21 288
rect 19 287 20 288
rect 18 287 19 288
rect 17 287 18 288
rect 16 287 17 288
rect 15 287 16 288
rect 14 287 15 288
rect 13 287 14 288
rect 12 287 13 288
rect 11 287 12 288
rect 10 287 11 288
rect 9 287 10 288
rect 8 287 9 288
rect 7 287 8 288
rect 6 287 7 288
rect 5 287 6 288
rect 464 288 465 289
rect 463 288 464 289
rect 462 288 463 289
rect 461 288 462 289
rect 441 288 442 289
rect 440 288 441 289
rect 439 288 440 289
rect 438 288 439 289
rect 437 288 438 289
rect 436 288 437 289
rect 435 288 436 289
rect 434 288 435 289
rect 433 288 434 289
rect 432 288 433 289
rect 431 288 432 289
rect 430 288 431 289
rect 429 288 430 289
rect 428 288 429 289
rect 427 288 428 289
rect 426 288 427 289
rect 425 288 426 289
rect 424 288 425 289
rect 423 288 424 289
rect 422 288 423 289
rect 421 288 422 289
rect 420 288 421 289
rect 419 288 420 289
rect 418 288 419 289
rect 417 288 418 289
rect 416 288 417 289
rect 415 288 416 289
rect 414 288 415 289
rect 413 288 414 289
rect 412 288 413 289
rect 411 288 412 289
rect 410 288 411 289
rect 409 288 410 289
rect 408 288 409 289
rect 407 288 408 289
rect 406 288 407 289
rect 405 288 406 289
rect 404 288 405 289
rect 403 288 404 289
rect 402 288 403 289
rect 401 288 402 289
rect 400 288 401 289
rect 399 288 400 289
rect 398 288 399 289
rect 397 288 398 289
rect 286 288 287 289
rect 285 288 286 289
rect 284 288 285 289
rect 283 288 284 289
rect 282 288 283 289
rect 281 288 282 289
rect 280 288 281 289
rect 279 288 280 289
rect 278 288 279 289
rect 277 288 278 289
rect 276 288 277 289
rect 275 288 276 289
rect 274 288 275 289
rect 273 288 274 289
rect 272 288 273 289
rect 271 288 272 289
rect 270 288 271 289
rect 269 288 270 289
rect 268 288 269 289
rect 267 288 268 289
rect 266 288 267 289
rect 265 288 266 289
rect 264 288 265 289
rect 263 288 264 289
rect 262 288 263 289
rect 261 288 262 289
rect 260 288 261 289
rect 259 288 260 289
rect 258 288 259 289
rect 257 288 258 289
rect 256 288 257 289
rect 255 288 256 289
rect 254 288 255 289
rect 253 288 254 289
rect 252 288 253 289
rect 251 288 252 289
rect 250 288 251 289
rect 249 288 250 289
rect 248 288 249 289
rect 247 288 248 289
rect 246 288 247 289
rect 245 288 246 289
rect 244 288 245 289
rect 243 288 244 289
rect 242 288 243 289
rect 241 288 242 289
rect 240 288 241 289
rect 239 288 240 289
rect 238 288 239 289
rect 237 288 238 289
rect 236 288 237 289
rect 235 288 236 289
rect 234 288 235 289
rect 233 288 234 289
rect 232 288 233 289
rect 231 288 232 289
rect 230 288 231 289
rect 229 288 230 289
rect 228 288 229 289
rect 227 288 228 289
rect 226 288 227 289
rect 225 288 226 289
rect 224 288 225 289
rect 223 288 224 289
rect 222 288 223 289
rect 221 288 222 289
rect 220 288 221 289
rect 219 288 220 289
rect 196 288 197 289
rect 195 288 196 289
rect 194 288 195 289
rect 193 288 194 289
rect 192 288 193 289
rect 191 288 192 289
rect 190 288 191 289
rect 189 288 190 289
rect 188 288 189 289
rect 187 288 188 289
rect 186 288 187 289
rect 185 288 186 289
rect 184 288 185 289
rect 183 288 184 289
rect 182 288 183 289
rect 181 288 182 289
rect 180 288 181 289
rect 179 288 180 289
rect 178 288 179 289
rect 177 288 178 289
rect 176 288 177 289
rect 175 288 176 289
rect 174 288 175 289
rect 173 288 174 289
rect 172 288 173 289
rect 171 288 172 289
rect 170 288 171 289
rect 169 288 170 289
rect 168 288 169 289
rect 167 288 168 289
rect 166 288 167 289
rect 165 288 166 289
rect 164 288 165 289
rect 163 288 164 289
rect 162 288 163 289
rect 161 288 162 289
rect 160 288 161 289
rect 159 288 160 289
rect 158 288 159 289
rect 157 288 158 289
rect 156 288 157 289
rect 155 288 156 289
rect 154 288 155 289
rect 153 288 154 289
rect 152 288 153 289
rect 151 288 152 289
rect 150 288 151 289
rect 149 288 150 289
rect 148 288 149 289
rect 147 288 148 289
rect 146 288 147 289
rect 145 288 146 289
rect 144 288 145 289
rect 143 288 144 289
rect 142 288 143 289
rect 141 288 142 289
rect 140 288 141 289
rect 139 288 140 289
rect 138 288 139 289
rect 137 288 138 289
rect 136 288 137 289
rect 135 288 136 289
rect 134 288 135 289
rect 118 288 119 289
rect 117 288 118 289
rect 116 288 117 289
rect 115 288 116 289
rect 114 288 115 289
rect 113 288 114 289
rect 112 288 113 289
rect 111 288 112 289
rect 110 288 111 289
rect 109 288 110 289
rect 108 288 109 289
rect 107 288 108 289
rect 106 288 107 289
rect 105 288 106 289
rect 104 288 105 289
rect 103 288 104 289
rect 102 288 103 289
rect 101 288 102 289
rect 100 288 101 289
rect 99 288 100 289
rect 98 288 99 289
rect 97 288 98 289
rect 96 288 97 289
rect 95 288 96 289
rect 94 288 95 289
rect 93 288 94 289
rect 92 288 93 289
rect 91 288 92 289
rect 90 288 91 289
rect 89 288 90 289
rect 88 288 89 289
rect 87 288 88 289
rect 86 288 87 289
rect 85 288 86 289
rect 84 288 85 289
rect 68 288 69 289
rect 67 288 68 289
rect 66 288 67 289
rect 65 288 66 289
rect 64 288 65 289
rect 63 288 64 289
rect 62 288 63 289
rect 61 288 62 289
rect 60 288 61 289
rect 59 288 60 289
rect 58 288 59 289
rect 57 288 58 289
rect 56 288 57 289
rect 55 288 56 289
rect 54 288 55 289
rect 53 288 54 289
rect 52 288 53 289
rect 51 288 52 289
rect 50 288 51 289
rect 49 288 50 289
rect 48 288 49 289
rect 47 288 48 289
rect 46 288 47 289
rect 45 288 46 289
rect 44 288 45 289
rect 43 288 44 289
rect 42 288 43 289
rect 41 288 42 289
rect 40 288 41 289
rect 30 288 31 289
rect 29 288 30 289
rect 28 288 29 289
rect 27 288 28 289
rect 26 288 27 289
rect 25 288 26 289
rect 24 288 25 289
rect 23 288 24 289
rect 22 288 23 289
rect 21 288 22 289
rect 20 288 21 289
rect 19 288 20 289
rect 18 288 19 289
rect 17 288 18 289
rect 16 288 17 289
rect 15 288 16 289
rect 14 288 15 289
rect 13 288 14 289
rect 12 288 13 289
rect 11 288 12 289
rect 10 288 11 289
rect 9 288 10 289
rect 8 288 9 289
rect 7 288 8 289
rect 6 288 7 289
rect 5 288 6 289
rect 463 289 464 290
rect 462 289 463 290
rect 441 289 442 290
rect 440 289 441 290
rect 439 289 440 290
rect 438 289 439 290
rect 437 289 438 290
rect 436 289 437 290
rect 435 289 436 290
rect 434 289 435 290
rect 433 289 434 290
rect 432 289 433 290
rect 431 289 432 290
rect 430 289 431 290
rect 429 289 430 290
rect 428 289 429 290
rect 427 289 428 290
rect 426 289 427 290
rect 425 289 426 290
rect 424 289 425 290
rect 423 289 424 290
rect 422 289 423 290
rect 421 289 422 290
rect 420 289 421 290
rect 419 289 420 290
rect 418 289 419 290
rect 417 289 418 290
rect 416 289 417 290
rect 415 289 416 290
rect 414 289 415 290
rect 413 289 414 290
rect 412 289 413 290
rect 411 289 412 290
rect 410 289 411 290
rect 409 289 410 290
rect 408 289 409 290
rect 407 289 408 290
rect 406 289 407 290
rect 405 289 406 290
rect 404 289 405 290
rect 403 289 404 290
rect 402 289 403 290
rect 401 289 402 290
rect 400 289 401 290
rect 399 289 400 290
rect 398 289 399 290
rect 397 289 398 290
rect 285 289 286 290
rect 284 289 285 290
rect 283 289 284 290
rect 282 289 283 290
rect 281 289 282 290
rect 280 289 281 290
rect 279 289 280 290
rect 278 289 279 290
rect 277 289 278 290
rect 276 289 277 290
rect 275 289 276 290
rect 274 289 275 290
rect 273 289 274 290
rect 272 289 273 290
rect 271 289 272 290
rect 270 289 271 290
rect 269 289 270 290
rect 268 289 269 290
rect 267 289 268 290
rect 266 289 267 290
rect 265 289 266 290
rect 264 289 265 290
rect 263 289 264 290
rect 262 289 263 290
rect 261 289 262 290
rect 260 289 261 290
rect 259 289 260 290
rect 258 289 259 290
rect 257 289 258 290
rect 256 289 257 290
rect 255 289 256 290
rect 254 289 255 290
rect 253 289 254 290
rect 252 289 253 290
rect 251 289 252 290
rect 250 289 251 290
rect 249 289 250 290
rect 248 289 249 290
rect 247 289 248 290
rect 246 289 247 290
rect 245 289 246 290
rect 244 289 245 290
rect 243 289 244 290
rect 242 289 243 290
rect 241 289 242 290
rect 240 289 241 290
rect 239 289 240 290
rect 238 289 239 290
rect 237 289 238 290
rect 236 289 237 290
rect 235 289 236 290
rect 234 289 235 290
rect 233 289 234 290
rect 232 289 233 290
rect 231 289 232 290
rect 230 289 231 290
rect 229 289 230 290
rect 228 289 229 290
rect 227 289 228 290
rect 226 289 227 290
rect 225 289 226 290
rect 224 289 225 290
rect 223 289 224 290
rect 222 289 223 290
rect 221 289 222 290
rect 220 289 221 290
rect 219 289 220 290
rect 218 289 219 290
rect 196 289 197 290
rect 195 289 196 290
rect 194 289 195 290
rect 193 289 194 290
rect 192 289 193 290
rect 191 289 192 290
rect 190 289 191 290
rect 189 289 190 290
rect 188 289 189 290
rect 187 289 188 290
rect 186 289 187 290
rect 185 289 186 290
rect 184 289 185 290
rect 183 289 184 290
rect 182 289 183 290
rect 181 289 182 290
rect 180 289 181 290
rect 179 289 180 290
rect 178 289 179 290
rect 177 289 178 290
rect 176 289 177 290
rect 175 289 176 290
rect 174 289 175 290
rect 173 289 174 290
rect 172 289 173 290
rect 171 289 172 290
rect 170 289 171 290
rect 169 289 170 290
rect 168 289 169 290
rect 167 289 168 290
rect 166 289 167 290
rect 165 289 166 290
rect 164 289 165 290
rect 163 289 164 290
rect 162 289 163 290
rect 161 289 162 290
rect 160 289 161 290
rect 159 289 160 290
rect 158 289 159 290
rect 157 289 158 290
rect 156 289 157 290
rect 155 289 156 290
rect 154 289 155 290
rect 153 289 154 290
rect 152 289 153 290
rect 151 289 152 290
rect 150 289 151 290
rect 149 289 150 290
rect 148 289 149 290
rect 147 289 148 290
rect 146 289 147 290
rect 145 289 146 290
rect 144 289 145 290
rect 143 289 144 290
rect 142 289 143 290
rect 141 289 142 290
rect 140 289 141 290
rect 139 289 140 290
rect 138 289 139 290
rect 137 289 138 290
rect 136 289 137 290
rect 135 289 136 290
rect 118 289 119 290
rect 117 289 118 290
rect 116 289 117 290
rect 115 289 116 290
rect 114 289 115 290
rect 113 289 114 290
rect 112 289 113 290
rect 111 289 112 290
rect 110 289 111 290
rect 109 289 110 290
rect 108 289 109 290
rect 107 289 108 290
rect 106 289 107 290
rect 105 289 106 290
rect 104 289 105 290
rect 103 289 104 290
rect 102 289 103 290
rect 101 289 102 290
rect 100 289 101 290
rect 99 289 100 290
rect 98 289 99 290
rect 97 289 98 290
rect 96 289 97 290
rect 95 289 96 290
rect 94 289 95 290
rect 93 289 94 290
rect 92 289 93 290
rect 91 289 92 290
rect 90 289 91 290
rect 89 289 90 290
rect 88 289 89 290
rect 87 289 88 290
rect 86 289 87 290
rect 85 289 86 290
rect 84 289 85 290
rect 68 289 69 290
rect 67 289 68 290
rect 66 289 67 290
rect 65 289 66 290
rect 64 289 65 290
rect 63 289 64 290
rect 62 289 63 290
rect 61 289 62 290
rect 60 289 61 290
rect 59 289 60 290
rect 58 289 59 290
rect 57 289 58 290
rect 56 289 57 290
rect 55 289 56 290
rect 54 289 55 290
rect 53 289 54 290
rect 52 289 53 290
rect 51 289 52 290
rect 50 289 51 290
rect 49 289 50 290
rect 48 289 49 290
rect 47 289 48 290
rect 46 289 47 290
rect 45 289 46 290
rect 44 289 45 290
rect 43 289 44 290
rect 42 289 43 290
rect 41 289 42 290
rect 40 289 41 290
rect 31 289 32 290
rect 30 289 31 290
rect 29 289 30 290
rect 28 289 29 290
rect 27 289 28 290
rect 26 289 27 290
rect 25 289 26 290
rect 24 289 25 290
rect 23 289 24 290
rect 22 289 23 290
rect 21 289 22 290
rect 20 289 21 290
rect 19 289 20 290
rect 18 289 19 290
rect 17 289 18 290
rect 16 289 17 290
rect 15 289 16 290
rect 14 289 15 290
rect 13 289 14 290
rect 12 289 13 290
rect 11 289 12 290
rect 10 289 11 290
rect 9 289 10 290
rect 8 289 9 290
rect 7 289 8 290
rect 6 289 7 290
rect 5 289 6 290
rect 462 290 463 291
rect 441 290 442 291
rect 440 290 441 291
rect 439 290 440 291
rect 438 290 439 291
rect 437 290 438 291
rect 436 290 437 291
rect 435 290 436 291
rect 434 290 435 291
rect 433 290 434 291
rect 432 290 433 291
rect 431 290 432 291
rect 430 290 431 291
rect 429 290 430 291
rect 428 290 429 291
rect 427 290 428 291
rect 426 290 427 291
rect 425 290 426 291
rect 424 290 425 291
rect 423 290 424 291
rect 422 290 423 291
rect 421 290 422 291
rect 420 290 421 291
rect 419 290 420 291
rect 418 290 419 291
rect 417 290 418 291
rect 416 290 417 291
rect 415 290 416 291
rect 414 290 415 291
rect 413 290 414 291
rect 412 290 413 291
rect 411 290 412 291
rect 410 290 411 291
rect 409 290 410 291
rect 408 290 409 291
rect 407 290 408 291
rect 406 290 407 291
rect 405 290 406 291
rect 404 290 405 291
rect 403 290 404 291
rect 402 290 403 291
rect 401 290 402 291
rect 400 290 401 291
rect 399 290 400 291
rect 398 290 399 291
rect 397 290 398 291
rect 284 290 285 291
rect 283 290 284 291
rect 282 290 283 291
rect 281 290 282 291
rect 280 290 281 291
rect 279 290 280 291
rect 278 290 279 291
rect 277 290 278 291
rect 276 290 277 291
rect 275 290 276 291
rect 274 290 275 291
rect 273 290 274 291
rect 272 290 273 291
rect 271 290 272 291
rect 270 290 271 291
rect 269 290 270 291
rect 268 290 269 291
rect 267 290 268 291
rect 266 290 267 291
rect 265 290 266 291
rect 264 290 265 291
rect 263 290 264 291
rect 262 290 263 291
rect 261 290 262 291
rect 260 290 261 291
rect 259 290 260 291
rect 258 290 259 291
rect 257 290 258 291
rect 256 290 257 291
rect 255 290 256 291
rect 254 290 255 291
rect 253 290 254 291
rect 252 290 253 291
rect 251 290 252 291
rect 250 290 251 291
rect 249 290 250 291
rect 248 290 249 291
rect 247 290 248 291
rect 246 290 247 291
rect 245 290 246 291
rect 244 290 245 291
rect 243 290 244 291
rect 242 290 243 291
rect 241 290 242 291
rect 240 290 241 291
rect 239 290 240 291
rect 238 290 239 291
rect 237 290 238 291
rect 236 290 237 291
rect 235 290 236 291
rect 234 290 235 291
rect 233 290 234 291
rect 232 290 233 291
rect 231 290 232 291
rect 230 290 231 291
rect 229 290 230 291
rect 228 290 229 291
rect 227 290 228 291
rect 226 290 227 291
rect 225 290 226 291
rect 224 290 225 291
rect 223 290 224 291
rect 222 290 223 291
rect 221 290 222 291
rect 220 290 221 291
rect 219 290 220 291
rect 218 290 219 291
rect 195 290 196 291
rect 194 290 195 291
rect 193 290 194 291
rect 192 290 193 291
rect 191 290 192 291
rect 190 290 191 291
rect 189 290 190 291
rect 188 290 189 291
rect 187 290 188 291
rect 186 290 187 291
rect 185 290 186 291
rect 184 290 185 291
rect 183 290 184 291
rect 182 290 183 291
rect 181 290 182 291
rect 180 290 181 291
rect 179 290 180 291
rect 178 290 179 291
rect 177 290 178 291
rect 176 290 177 291
rect 175 290 176 291
rect 174 290 175 291
rect 173 290 174 291
rect 172 290 173 291
rect 171 290 172 291
rect 170 290 171 291
rect 169 290 170 291
rect 168 290 169 291
rect 167 290 168 291
rect 166 290 167 291
rect 165 290 166 291
rect 164 290 165 291
rect 163 290 164 291
rect 162 290 163 291
rect 161 290 162 291
rect 160 290 161 291
rect 159 290 160 291
rect 158 290 159 291
rect 157 290 158 291
rect 156 290 157 291
rect 155 290 156 291
rect 154 290 155 291
rect 153 290 154 291
rect 152 290 153 291
rect 151 290 152 291
rect 150 290 151 291
rect 149 290 150 291
rect 148 290 149 291
rect 147 290 148 291
rect 146 290 147 291
rect 145 290 146 291
rect 144 290 145 291
rect 143 290 144 291
rect 142 290 143 291
rect 141 290 142 291
rect 140 290 141 291
rect 139 290 140 291
rect 138 290 139 291
rect 137 290 138 291
rect 136 290 137 291
rect 135 290 136 291
rect 119 290 120 291
rect 118 290 119 291
rect 117 290 118 291
rect 116 290 117 291
rect 115 290 116 291
rect 114 290 115 291
rect 113 290 114 291
rect 112 290 113 291
rect 111 290 112 291
rect 110 290 111 291
rect 109 290 110 291
rect 108 290 109 291
rect 107 290 108 291
rect 106 290 107 291
rect 105 290 106 291
rect 104 290 105 291
rect 103 290 104 291
rect 102 290 103 291
rect 101 290 102 291
rect 100 290 101 291
rect 99 290 100 291
rect 98 290 99 291
rect 97 290 98 291
rect 96 290 97 291
rect 95 290 96 291
rect 94 290 95 291
rect 93 290 94 291
rect 92 290 93 291
rect 91 290 92 291
rect 90 290 91 291
rect 89 290 90 291
rect 88 290 89 291
rect 87 290 88 291
rect 86 290 87 291
rect 85 290 86 291
rect 84 290 85 291
rect 68 290 69 291
rect 67 290 68 291
rect 66 290 67 291
rect 65 290 66 291
rect 64 290 65 291
rect 63 290 64 291
rect 62 290 63 291
rect 61 290 62 291
rect 60 290 61 291
rect 59 290 60 291
rect 58 290 59 291
rect 57 290 58 291
rect 56 290 57 291
rect 55 290 56 291
rect 54 290 55 291
rect 53 290 54 291
rect 52 290 53 291
rect 51 290 52 291
rect 50 290 51 291
rect 49 290 50 291
rect 48 290 49 291
rect 47 290 48 291
rect 46 290 47 291
rect 45 290 46 291
rect 44 290 45 291
rect 43 290 44 291
rect 42 290 43 291
rect 41 290 42 291
rect 40 290 41 291
rect 31 290 32 291
rect 30 290 31 291
rect 29 290 30 291
rect 28 290 29 291
rect 27 290 28 291
rect 26 290 27 291
rect 25 290 26 291
rect 24 290 25 291
rect 23 290 24 291
rect 22 290 23 291
rect 21 290 22 291
rect 20 290 21 291
rect 19 290 20 291
rect 18 290 19 291
rect 17 290 18 291
rect 16 290 17 291
rect 15 290 16 291
rect 14 290 15 291
rect 13 290 14 291
rect 12 290 13 291
rect 11 290 12 291
rect 10 290 11 291
rect 9 290 10 291
rect 8 290 9 291
rect 7 290 8 291
rect 6 290 7 291
rect 5 290 6 291
rect 482 291 483 292
rect 462 291 463 292
rect 441 291 442 292
rect 440 291 441 292
rect 439 291 440 292
rect 438 291 439 292
rect 437 291 438 292
rect 436 291 437 292
rect 420 291 421 292
rect 419 291 420 292
rect 418 291 419 292
rect 417 291 418 292
rect 416 291 417 292
rect 403 291 404 292
rect 402 291 403 292
rect 401 291 402 292
rect 400 291 401 292
rect 399 291 400 292
rect 398 291 399 292
rect 397 291 398 292
rect 283 291 284 292
rect 282 291 283 292
rect 281 291 282 292
rect 280 291 281 292
rect 279 291 280 292
rect 278 291 279 292
rect 277 291 278 292
rect 276 291 277 292
rect 275 291 276 292
rect 274 291 275 292
rect 273 291 274 292
rect 272 291 273 292
rect 271 291 272 292
rect 270 291 271 292
rect 269 291 270 292
rect 268 291 269 292
rect 267 291 268 292
rect 266 291 267 292
rect 265 291 266 292
rect 264 291 265 292
rect 263 291 264 292
rect 262 291 263 292
rect 261 291 262 292
rect 260 291 261 292
rect 259 291 260 292
rect 258 291 259 292
rect 257 291 258 292
rect 256 291 257 292
rect 255 291 256 292
rect 254 291 255 292
rect 253 291 254 292
rect 252 291 253 292
rect 251 291 252 292
rect 250 291 251 292
rect 249 291 250 292
rect 248 291 249 292
rect 247 291 248 292
rect 246 291 247 292
rect 245 291 246 292
rect 244 291 245 292
rect 243 291 244 292
rect 242 291 243 292
rect 241 291 242 292
rect 240 291 241 292
rect 239 291 240 292
rect 238 291 239 292
rect 237 291 238 292
rect 236 291 237 292
rect 235 291 236 292
rect 234 291 235 292
rect 233 291 234 292
rect 232 291 233 292
rect 231 291 232 292
rect 230 291 231 292
rect 229 291 230 292
rect 228 291 229 292
rect 227 291 228 292
rect 226 291 227 292
rect 225 291 226 292
rect 224 291 225 292
rect 223 291 224 292
rect 222 291 223 292
rect 221 291 222 292
rect 220 291 221 292
rect 219 291 220 292
rect 218 291 219 292
rect 217 291 218 292
rect 194 291 195 292
rect 193 291 194 292
rect 192 291 193 292
rect 191 291 192 292
rect 190 291 191 292
rect 189 291 190 292
rect 188 291 189 292
rect 187 291 188 292
rect 186 291 187 292
rect 185 291 186 292
rect 184 291 185 292
rect 183 291 184 292
rect 182 291 183 292
rect 181 291 182 292
rect 180 291 181 292
rect 179 291 180 292
rect 178 291 179 292
rect 177 291 178 292
rect 176 291 177 292
rect 175 291 176 292
rect 174 291 175 292
rect 173 291 174 292
rect 172 291 173 292
rect 171 291 172 292
rect 170 291 171 292
rect 169 291 170 292
rect 168 291 169 292
rect 167 291 168 292
rect 166 291 167 292
rect 165 291 166 292
rect 164 291 165 292
rect 163 291 164 292
rect 162 291 163 292
rect 161 291 162 292
rect 160 291 161 292
rect 159 291 160 292
rect 158 291 159 292
rect 157 291 158 292
rect 156 291 157 292
rect 155 291 156 292
rect 154 291 155 292
rect 153 291 154 292
rect 152 291 153 292
rect 151 291 152 292
rect 150 291 151 292
rect 149 291 150 292
rect 148 291 149 292
rect 147 291 148 292
rect 146 291 147 292
rect 145 291 146 292
rect 144 291 145 292
rect 143 291 144 292
rect 142 291 143 292
rect 141 291 142 292
rect 140 291 141 292
rect 139 291 140 292
rect 138 291 139 292
rect 137 291 138 292
rect 136 291 137 292
rect 119 291 120 292
rect 118 291 119 292
rect 117 291 118 292
rect 116 291 117 292
rect 115 291 116 292
rect 114 291 115 292
rect 113 291 114 292
rect 112 291 113 292
rect 111 291 112 292
rect 110 291 111 292
rect 109 291 110 292
rect 108 291 109 292
rect 107 291 108 292
rect 106 291 107 292
rect 105 291 106 292
rect 104 291 105 292
rect 103 291 104 292
rect 102 291 103 292
rect 101 291 102 292
rect 100 291 101 292
rect 99 291 100 292
rect 98 291 99 292
rect 97 291 98 292
rect 96 291 97 292
rect 95 291 96 292
rect 94 291 95 292
rect 93 291 94 292
rect 92 291 93 292
rect 91 291 92 292
rect 90 291 91 292
rect 89 291 90 292
rect 88 291 89 292
rect 87 291 88 292
rect 86 291 87 292
rect 85 291 86 292
rect 69 291 70 292
rect 68 291 69 292
rect 67 291 68 292
rect 66 291 67 292
rect 65 291 66 292
rect 64 291 65 292
rect 63 291 64 292
rect 62 291 63 292
rect 61 291 62 292
rect 60 291 61 292
rect 59 291 60 292
rect 58 291 59 292
rect 57 291 58 292
rect 56 291 57 292
rect 55 291 56 292
rect 54 291 55 292
rect 53 291 54 292
rect 52 291 53 292
rect 51 291 52 292
rect 50 291 51 292
rect 49 291 50 292
rect 48 291 49 292
rect 47 291 48 292
rect 46 291 47 292
rect 45 291 46 292
rect 44 291 45 292
rect 43 291 44 292
rect 42 291 43 292
rect 41 291 42 292
rect 40 291 41 292
rect 31 291 32 292
rect 30 291 31 292
rect 29 291 30 292
rect 28 291 29 292
rect 27 291 28 292
rect 26 291 27 292
rect 25 291 26 292
rect 24 291 25 292
rect 23 291 24 292
rect 22 291 23 292
rect 21 291 22 292
rect 20 291 21 292
rect 19 291 20 292
rect 18 291 19 292
rect 17 291 18 292
rect 16 291 17 292
rect 15 291 16 292
rect 14 291 15 292
rect 13 291 14 292
rect 12 291 13 292
rect 11 291 12 292
rect 10 291 11 292
rect 9 291 10 292
rect 8 291 9 292
rect 7 291 8 292
rect 6 291 7 292
rect 5 291 6 292
rect 482 292 483 293
rect 462 292 463 293
rect 441 292 442 293
rect 440 292 441 293
rect 439 292 440 293
rect 438 292 439 293
rect 419 292 420 293
rect 418 292 419 293
rect 417 292 418 293
rect 416 292 417 293
rect 400 292 401 293
rect 399 292 400 293
rect 398 292 399 293
rect 397 292 398 293
rect 282 292 283 293
rect 281 292 282 293
rect 280 292 281 293
rect 279 292 280 293
rect 278 292 279 293
rect 277 292 278 293
rect 276 292 277 293
rect 275 292 276 293
rect 274 292 275 293
rect 273 292 274 293
rect 272 292 273 293
rect 271 292 272 293
rect 270 292 271 293
rect 269 292 270 293
rect 268 292 269 293
rect 267 292 268 293
rect 266 292 267 293
rect 265 292 266 293
rect 264 292 265 293
rect 263 292 264 293
rect 262 292 263 293
rect 261 292 262 293
rect 260 292 261 293
rect 259 292 260 293
rect 258 292 259 293
rect 257 292 258 293
rect 256 292 257 293
rect 255 292 256 293
rect 254 292 255 293
rect 253 292 254 293
rect 252 292 253 293
rect 251 292 252 293
rect 250 292 251 293
rect 249 292 250 293
rect 248 292 249 293
rect 247 292 248 293
rect 246 292 247 293
rect 245 292 246 293
rect 244 292 245 293
rect 243 292 244 293
rect 242 292 243 293
rect 241 292 242 293
rect 240 292 241 293
rect 239 292 240 293
rect 238 292 239 293
rect 237 292 238 293
rect 236 292 237 293
rect 235 292 236 293
rect 234 292 235 293
rect 233 292 234 293
rect 232 292 233 293
rect 231 292 232 293
rect 230 292 231 293
rect 229 292 230 293
rect 228 292 229 293
rect 227 292 228 293
rect 226 292 227 293
rect 225 292 226 293
rect 224 292 225 293
rect 223 292 224 293
rect 222 292 223 293
rect 221 292 222 293
rect 220 292 221 293
rect 219 292 220 293
rect 218 292 219 293
rect 217 292 218 293
rect 193 292 194 293
rect 192 292 193 293
rect 191 292 192 293
rect 190 292 191 293
rect 189 292 190 293
rect 188 292 189 293
rect 187 292 188 293
rect 186 292 187 293
rect 185 292 186 293
rect 184 292 185 293
rect 183 292 184 293
rect 182 292 183 293
rect 181 292 182 293
rect 180 292 181 293
rect 179 292 180 293
rect 178 292 179 293
rect 177 292 178 293
rect 176 292 177 293
rect 175 292 176 293
rect 174 292 175 293
rect 173 292 174 293
rect 172 292 173 293
rect 171 292 172 293
rect 170 292 171 293
rect 169 292 170 293
rect 168 292 169 293
rect 167 292 168 293
rect 166 292 167 293
rect 165 292 166 293
rect 164 292 165 293
rect 163 292 164 293
rect 162 292 163 293
rect 161 292 162 293
rect 160 292 161 293
rect 159 292 160 293
rect 158 292 159 293
rect 157 292 158 293
rect 156 292 157 293
rect 155 292 156 293
rect 154 292 155 293
rect 153 292 154 293
rect 152 292 153 293
rect 151 292 152 293
rect 150 292 151 293
rect 149 292 150 293
rect 148 292 149 293
rect 147 292 148 293
rect 146 292 147 293
rect 145 292 146 293
rect 144 292 145 293
rect 143 292 144 293
rect 142 292 143 293
rect 141 292 142 293
rect 140 292 141 293
rect 139 292 140 293
rect 138 292 139 293
rect 137 292 138 293
rect 120 292 121 293
rect 119 292 120 293
rect 118 292 119 293
rect 117 292 118 293
rect 116 292 117 293
rect 115 292 116 293
rect 114 292 115 293
rect 113 292 114 293
rect 112 292 113 293
rect 111 292 112 293
rect 110 292 111 293
rect 109 292 110 293
rect 108 292 109 293
rect 107 292 108 293
rect 106 292 107 293
rect 105 292 106 293
rect 104 292 105 293
rect 103 292 104 293
rect 102 292 103 293
rect 101 292 102 293
rect 100 292 101 293
rect 99 292 100 293
rect 98 292 99 293
rect 97 292 98 293
rect 96 292 97 293
rect 95 292 96 293
rect 94 292 95 293
rect 93 292 94 293
rect 92 292 93 293
rect 91 292 92 293
rect 90 292 91 293
rect 89 292 90 293
rect 88 292 89 293
rect 87 292 88 293
rect 86 292 87 293
rect 85 292 86 293
rect 69 292 70 293
rect 68 292 69 293
rect 67 292 68 293
rect 66 292 67 293
rect 65 292 66 293
rect 64 292 65 293
rect 63 292 64 293
rect 62 292 63 293
rect 61 292 62 293
rect 60 292 61 293
rect 59 292 60 293
rect 58 292 59 293
rect 57 292 58 293
rect 56 292 57 293
rect 55 292 56 293
rect 54 292 55 293
rect 53 292 54 293
rect 52 292 53 293
rect 51 292 52 293
rect 50 292 51 293
rect 49 292 50 293
rect 48 292 49 293
rect 47 292 48 293
rect 46 292 47 293
rect 45 292 46 293
rect 44 292 45 293
rect 43 292 44 293
rect 42 292 43 293
rect 41 292 42 293
rect 40 292 41 293
rect 31 292 32 293
rect 30 292 31 293
rect 29 292 30 293
rect 28 292 29 293
rect 27 292 28 293
rect 26 292 27 293
rect 25 292 26 293
rect 24 292 25 293
rect 23 292 24 293
rect 22 292 23 293
rect 21 292 22 293
rect 20 292 21 293
rect 19 292 20 293
rect 18 292 19 293
rect 17 292 18 293
rect 16 292 17 293
rect 15 292 16 293
rect 14 292 15 293
rect 13 292 14 293
rect 12 292 13 293
rect 11 292 12 293
rect 10 292 11 293
rect 9 292 10 293
rect 8 292 9 293
rect 7 292 8 293
rect 6 292 7 293
rect 5 292 6 293
rect 482 293 483 294
rect 481 293 482 294
rect 462 293 463 294
rect 441 293 442 294
rect 440 293 441 294
rect 439 293 440 294
rect 419 293 420 294
rect 418 293 419 294
rect 417 293 418 294
rect 416 293 417 294
rect 399 293 400 294
rect 398 293 399 294
rect 397 293 398 294
rect 281 293 282 294
rect 280 293 281 294
rect 279 293 280 294
rect 278 293 279 294
rect 277 293 278 294
rect 276 293 277 294
rect 275 293 276 294
rect 274 293 275 294
rect 273 293 274 294
rect 272 293 273 294
rect 271 293 272 294
rect 270 293 271 294
rect 269 293 270 294
rect 268 293 269 294
rect 267 293 268 294
rect 266 293 267 294
rect 265 293 266 294
rect 264 293 265 294
rect 263 293 264 294
rect 262 293 263 294
rect 261 293 262 294
rect 260 293 261 294
rect 259 293 260 294
rect 258 293 259 294
rect 257 293 258 294
rect 256 293 257 294
rect 255 293 256 294
rect 254 293 255 294
rect 253 293 254 294
rect 252 293 253 294
rect 251 293 252 294
rect 250 293 251 294
rect 249 293 250 294
rect 248 293 249 294
rect 247 293 248 294
rect 246 293 247 294
rect 245 293 246 294
rect 244 293 245 294
rect 243 293 244 294
rect 242 293 243 294
rect 241 293 242 294
rect 240 293 241 294
rect 239 293 240 294
rect 238 293 239 294
rect 237 293 238 294
rect 236 293 237 294
rect 235 293 236 294
rect 234 293 235 294
rect 233 293 234 294
rect 232 293 233 294
rect 231 293 232 294
rect 230 293 231 294
rect 229 293 230 294
rect 228 293 229 294
rect 227 293 228 294
rect 226 293 227 294
rect 225 293 226 294
rect 224 293 225 294
rect 223 293 224 294
rect 222 293 223 294
rect 221 293 222 294
rect 220 293 221 294
rect 219 293 220 294
rect 218 293 219 294
rect 217 293 218 294
rect 216 293 217 294
rect 193 293 194 294
rect 192 293 193 294
rect 191 293 192 294
rect 190 293 191 294
rect 189 293 190 294
rect 188 293 189 294
rect 187 293 188 294
rect 186 293 187 294
rect 185 293 186 294
rect 184 293 185 294
rect 183 293 184 294
rect 182 293 183 294
rect 181 293 182 294
rect 180 293 181 294
rect 179 293 180 294
rect 178 293 179 294
rect 177 293 178 294
rect 176 293 177 294
rect 175 293 176 294
rect 174 293 175 294
rect 173 293 174 294
rect 172 293 173 294
rect 171 293 172 294
rect 170 293 171 294
rect 169 293 170 294
rect 168 293 169 294
rect 167 293 168 294
rect 166 293 167 294
rect 165 293 166 294
rect 164 293 165 294
rect 163 293 164 294
rect 162 293 163 294
rect 161 293 162 294
rect 160 293 161 294
rect 159 293 160 294
rect 158 293 159 294
rect 157 293 158 294
rect 156 293 157 294
rect 155 293 156 294
rect 154 293 155 294
rect 153 293 154 294
rect 152 293 153 294
rect 151 293 152 294
rect 150 293 151 294
rect 149 293 150 294
rect 148 293 149 294
rect 147 293 148 294
rect 146 293 147 294
rect 145 293 146 294
rect 144 293 145 294
rect 143 293 144 294
rect 142 293 143 294
rect 141 293 142 294
rect 140 293 141 294
rect 139 293 140 294
rect 138 293 139 294
rect 137 293 138 294
rect 120 293 121 294
rect 119 293 120 294
rect 118 293 119 294
rect 117 293 118 294
rect 116 293 117 294
rect 115 293 116 294
rect 114 293 115 294
rect 113 293 114 294
rect 112 293 113 294
rect 111 293 112 294
rect 110 293 111 294
rect 109 293 110 294
rect 108 293 109 294
rect 107 293 108 294
rect 106 293 107 294
rect 105 293 106 294
rect 104 293 105 294
rect 103 293 104 294
rect 102 293 103 294
rect 101 293 102 294
rect 100 293 101 294
rect 99 293 100 294
rect 98 293 99 294
rect 97 293 98 294
rect 96 293 97 294
rect 95 293 96 294
rect 94 293 95 294
rect 93 293 94 294
rect 92 293 93 294
rect 91 293 92 294
rect 90 293 91 294
rect 89 293 90 294
rect 88 293 89 294
rect 87 293 88 294
rect 86 293 87 294
rect 85 293 86 294
rect 69 293 70 294
rect 68 293 69 294
rect 67 293 68 294
rect 66 293 67 294
rect 65 293 66 294
rect 64 293 65 294
rect 63 293 64 294
rect 62 293 63 294
rect 61 293 62 294
rect 60 293 61 294
rect 59 293 60 294
rect 58 293 59 294
rect 57 293 58 294
rect 56 293 57 294
rect 55 293 56 294
rect 54 293 55 294
rect 53 293 54 294
rect 52 293 53 294
rect 51 293 52 294
rect 50 293 51 294
rect 49 293 50 294
rect 48 293 49 294
rect 47 293 48 294
rect 46 293 47 294
rect 45 293 46 294
rect 44 293 45 294
rect 43 293 44 294
rect 42 293 43 294
rect 41 293 42 294
rect 40 293 41 294
rect 31 293 32 294
rect 30 293 31 294
rect 29 293 30 294
rect 28 293 29 294
rect 27 293 28 294
rect 26 293 27 294
rect 25 293 26 294
rect 24 293 25 294
rect 23 293 24 294
rect 22 293 23 294
rect 21 293 22 294
rect 20 293 21 294
rect 19 293 20 294
rect 18 293 19 294
rect 17 293 18 294
rect 16 293 17 294
rect 15 293 16 294
rect 14 293 15 294
rect 13 293 14 294
rect 12 293 13 294
rect 11 293 12 294
rect 10 293 11 294
rect 9 293 10 294
rect 8 293 9 294
rect 7 293 8 294
rect 6 293 7 294
rect 5 293 6 294
rect 482 294 483 295
rect 481 294 482 295
rect 480 294 481 295
rect 479 294 480 295
rect 478 294 479 295
rect 477 294 478 295
rect 476 294 477 295
rect 475 294 476 295
rect 474 294 475 295
rect 473 294 474 295
rect 472 294 473 295
rect 471 294 472 295
rect 470 294 471 295
rect 469 294 470 295
rect 468 294 469 295
rect 467 294 468 295
rect 466 294 467 295
rect 465 294 466 295
rect 464 294 465 295
rect 463 294 464 295
rect 462 294 463 295
rect 441 294 442 295
rect 440 294 441 295
rect 439 294 440 295
rect 419 294 420 295
rect 418 294 419 295
rect 417 294 418 295
rect 416 294 417 295
rect 399 294 400 295
rect 398 294 399 295
rect 397 294 398 295
rect 280 294 281 295
rect 279 294 280 295
rect 278 294 279 295
rect 277 294 278 295
rect 276 294 277 295
rect 275 294 276 295
rect 274 294 275 295
rect 273 294 274 295
rect 272 294 273 295
rect 271 294 272 295
rect 270 294 271 295
rect 269 294 270 295
rect 268 294 269 295
rect 267 294 268 295
rect 266 294 267 295
rect 265 294 266 295
rect 264 294 265 295
rect 263 294 264 295
rect 262 294 263 295
rect 261 294 262 295
rect 260 294 261 295
rect 259 294 260 295
rect 258 294 259 295
rect 257 294 258 295
rect 256 294 257 295
rect 255 294 256 295
rect 254 294 255 295
rect 253 294 254 295
rect 252 294 253 295
rect 251 294 252 295
rect 250 294 251 295
rect 249 294 250 295
rect 248 294 249 295
rect 247 294 248 295
rect 246 294 247 295
rect 245 294 246 295
rect 244 294 245 295
rect 243 294 244 295
rect 242 294 243 295
rect 241 294 242 295
rect 240 294 241 295
rect 239 294 240 295
rect 238 294 239 295
rect 237 294 238 295
rect 236 294 237 295
rect 235 294 236 295
rect 234 294 235 295
rect 233 294 234 295
rect 232 294 233 295
rect 231 294 232 295
rect 230 294 231 295
rect 229 294 230 295
rect 228 294 229 295
rect 227 294 228 295
rect 226 294 227 295
rect 225 294 226 295
rect 224 294 225 295
rect 223 294 224 295
rect 222 294 223 295
rect 221 294 222 295
rect 220 294 221 295
rect 219 294 220 295
rect 218 294 219 295
rect 217 294 218 295
rect 216 294 217 295
rect 215 294 216 295
rect 192 294 193 295
rect 191 294 192 295
rect 190 294 191 295
rect 189 294 190 295
rect 188 294 189 295
rect 187 294 188 295
rect 186 294 187 295
rect 185 294 186 295
rect 184 294 185 295
rect 183 294 184 295
rect 182 294 183 295
rect 181 294 182 295
rect 180 294 181 295
rect 179 294 180 295
rect 178 294 179 295
rect 177 294 178 295
rect 176 294 177 295
rect 175 294 176 295
rect 174 294 175 295
rect 173 294 174 295
rect 172 294 173 295
rect 171 294 172 295
rect 170 294 171 295
rect 169 294 170 295
rect 168 294 169 295
rect 167 294 168 295
rect 166 294 167 295
rect 165 294 166 295
rect 164 294 165 295
rect 163 294 164 295
rect 162 294 163 295
rect 161 294 162 295
rect 160 294 161 295
rect 159 294 160 295
rect 158 294 159 295
rect 157 294 158 295
rect 156 294 157 295
rect 155 294 156 295
rect 154 294 155 295
rect 153 294 154 295
rect 152 294 153 295
rect 151 294 152 295
rect 150 294 151 295
rect 149 294 150 295
rect 148 294 149 295
rect 147 294 148 295
rect 146 294 147 295
rect 145 294 146 295
rect 144 294 145 295
rect 143 294 144 295
rect 142 294 143 295
rect 141 294 142 295
rect 140 294 141 295
rect 139 294 140 295
rect 138 294 139 295
rect 120 294 121 295
rect 119 294 120 295
rect 118 294 119 295
rect 117 294 118 295
rect 116 294 117 295
rect 115 294 116 295
rect 114 294 115 295
rect 113 294 114 295
rect 112 294 113 295
rect 111 294 112 295
rect 110 294 111 295
rect 109 294 110 295
rect 108 294 109 295
rect 107 294 108 295
rect 106 294 107 295
rect 105 294 106 295
rect 104 294 105 295
rect 103 294 104 295
rect 102 294 103 295
rect 101 294 102 295
rect 100 294 101 295
rect 99 294 100 295
rect 98 294 99 295
rect 97 294 98 295
rect 96 294 97 295
rect 95 294 96 295
rect 94 294 95 295
rect 93 294 94 295
rect 92 294 93 295
rect 91 294 92 295
rect 90 294 91 295
rect 89 294 90 295
rect 88 294 89 295
rect 87 294 88 295
rect 86 294 87 295
rect 85 294 86 295
rect 69 294 70 295
rect 68 294 69 295
rect 67 294 68 295
rect 66 294 67 295
rect 65 294 66 295
rect 64 294 65 295
rect 63 294 64 295
rect 62 294 63 295
rect 61 294 62 295
rect 60 294 61 295
rect 59 294 60 295
rect 58 294 59 295
rect 57 294 58 295
rect 56 294 57 295
rect 55 294 56 295
rect 54 294 55 295
rect 53 294 54 295
rect 52 294 53 295
rect 51 294 52 295
rect 50 294 51 295
rect 49 294 50 295
rect 48 294 49 295
rect 47 294 48 295
rect 46 294 47 295
rect 45 294 46 295
rect 44 294 45 295
rect 43 294 44 295
rect 42 294 43 295
rect 41 294 42 295
rect 31 294 32 295
rect 30 294 31 295
rect 29 294 30 295
rect 28 294 29 295
rect 27 294 28 295
rect 26 294 27 295
rect 25 294 26 295
rect 24 294 25 295
rect 23 294 24 295
rect 22 294 23 295
rect 21 294 22 295
rect 20 294 21 295
rect 19 294 20 295
rect 18 294 19 295
rect 17 294 18 295
rect 16 294 17 295
rect 15 294 16 295
rect 14 294 15 295
rect 13 294 14 295
rect 12 294 13 295
rect 11 294 12 295
rect 10 294 11 295
rect 9 294 10 295
rect 8 294 9 295
rect 7 294 8 295
rect 6 294 7 295
rect 5 294 6 295
rect 482 295 483 296
rect 481 295 482 296
rect 480 295 481 296
rect 479 295 480 296
rect 478 295 479 296
rect 477 295 478 296
rect 476 295 477 296
rect 475 295 476 296
rect 474 295 475 296
rect 473 295 474 296
rect 472 295 473 296
rect 471 295 472 296
rect 470 295 471 296
rect 469 295 470 296
rect 468 295 469 296
rect 467 295 468 296
rect 466 295 467 296
rect 465 295 466 296
rect 464 295 465 296
rect 463 295 464 296
rect 462 295 463 296
rect 441 295 442 296
rect 440 295 441 296
rect 439 295 440 296
rect 419 295 420 296
rect 418 295 419 296
rect 417 295 418 296
rect 416 295 417 296
rect 399 295 400 296
rect 398 295 399 296
rect 397 295 398 296
rect 279 295 280 296
rect 278 295 279 296
rect 277 295 278 296
rect 276 295 277 296
rect 275 295 276 296
rect 274 295 275 296
rect 273 295 274 296
rect 272 295 273 296
rect 271 295 272 296
rect 270 295 271 296
rect 269 295 270 296
rect 268 295 269 296
rect 267 295 268 296
rect 266 295 267 296
rect 265 295 266 296
rect 264 295 265 296
rect 263 295 264 296
rect 262 295 263 296
rect 261 295 262 296
rect 260 295 261 296
rect 259 295 260 296
rect 258 295 259 296
rect 257 295 258 296
rect 256 295 257 296
rect 255 295 256 296
rect 254 295 255 296
rect 253 295 254 296
rect 252 295 253 296
rect 251 295 252 296
rect 250 295 251 296
rect 249 295 250 296
rect 248 295 249 296
rect 247 295 248 296
rect 246 295 247 296
rect 245 295 246 296
rect 244 295 245 296
rect 243 295 244 296
rect 242 295 243 296
rect 241 295 242 296
rect 240 295 241 296
rect 239 295 240 296
rect 238 295 239 296
rect 237 295 238 296
rect 236 295 237 296
rect 235 295 236 296
rect 234 295 235 296
rect 233 295 234 296
rect 232 295 233 296
rect 231 295 232 296
rect 230 295 231 296
rect 229 295 230 296
rect 228 295 229 296
rect 227 295 228 296
rect 226 295 227 296
rect 225 295 226 296
rect 224 295 225 296
rect 223 295 224 296
rect 222 295 223 296
rect 221 295 222 296
rect 220 295 221 296
rect 219 295 220 296
rect 218 295 219 296
rect 217 295 218 296
rect 216 295 217 296
rect 215 295 216 296
rect 191 295 192 296
rect 190 295 191 296
rect 189 295 190 296
rect 188 295 189 296
rect 187 295 188 296
rect 186 295 187 296
rect 185 295 186 296
rect 184 295 185 296
rect 183 295 184 296
rect 182 295 183 296
rect 181 295 182 296
rect 180 295 181 296
rect 179 295 180 296
rect 178 295 179 296
rect 177 295 178 296
rect 176 295 177 296
rect 175 295 176 296
rect 174 295 175 296
rect 173 295 174 296
rect 172 295 173 296
rect 171 295 172 296
rect 170 295 171 296
rect 169 295 170 296
rect 168 295 169 296
rect 167 295 168 296
rect 166 295 167 296
rect 165 295 166 296
rect 164 295 165 296
rect 163 295 164 296
rect 162 295 163 296
rect 161 295 162 296
rect 160 295 161 296
rect 159 295 160 296
rect 158 295 159 296
rect 157 295 158 296
rect 156 295 157 296
rect 155 295 156 296
rect 154 295 155 296
rect 153 295 154 296
rect 152 295 153 296
rect 151 295 152 296
rect 150 295 151 296
rect 149 295 150 296
rect 148 295 149 296
rect 147 295 148 296
rect 146 295 147 296
rect 145 295 146 296
rect 144 295 145 296
rect 143 295 144 296
rect 142 295 143 296
rect 141 295 142 296
rect 140 295 141 296
rect 139 295 140 296
rect 121 295 122 296
rect 120 295 121 296
rect 119 295 120 296
rect 118 295 119 296
rect 117 295 118 296
rect 116 295 117 296
rect 115 295 116 296
rect 114 295 115 296
rect 113 295 114 296
rect 112 295 113 296
rect 111 295 112 296
rect 110 295 111 296
rect 109 295 110 296
rect 108 295 109 296
rect 107 295 108 296
rect 106 295 107 296
rect 105 295 106 296
rect 104 295 105 296
rect 103 295 104 296
rect 102 295 103 296
rect 101 295 102 296
rect 100 295 101 296
rect 99 295 100 296
rect 98 295 99 296
rect 97 295 98 296
rect 96 295 97 296
rect 95 295 96 296
rect 94 295 95 296
rect 93 295 94 296
rect 92 295 93 296
rect 91 295 92 296
rect 90 295 91 296
rect 89 295 90 296
rect 88 295 89 296
rect 87 295 88 296
rect 86 295 87 296
rect 70 295 71 296
rect 69 295 70 296
rect 68 295 69 296
rect 67 295 68 296
rect 66 295 67 296
rect 65 295 66 296
rect 64 295 65 296
rect 63 295 64 296
rect 62 295 63 296
rect 61 295 62 296
rect 60 295 61 296
rect 59 295 60 296
rect 58 295 59 296
rect 57 295 58 296
rect 56 295 57 296
rect 55 295 56 296
rect 54 295 55 296
rect 53 295 54 296
rect 52 295 53 296
rect 51 295 52 296
rect 50 295 51 296
rect 49 295 50 296
rect 48 295 49 296
rect 47 295 48 296
rect 46 295 47 296
rect 45 295 46 296
rect 44 295 45 296
rect 43 295 44 296
rect 42 295 43 296
rect 41 295 42 296
rect 31 295 32 296
rect 30 295 31 296
rect 29 295 30 296
rect 28 295 29 296
rect 27 295 28 296
rect 26 295 27 296
rect 25 295 26 296
rect 24 295 25 296
rect 23 295 24 296
rect 22 295 23 296
rect 21 295 22 296
rect 20 295 21 296
rect 19 295 20 296
rect 18 295 19 296
rect 17 295 18 296
rect 16 295 17 296
rect 15 295 16 296
rect 14 295 15 296
rect 13 295 14 296
rect 12 295 13 296
rect 11 295 12 296
rect 10 295 11 296
rect 9 295 10 296
rect 8 295 9 296
rect 7 295 8 296
rect 6 295 7 296
rect 5 295 6 296
rect 482 296 483 297
rect 481 296 482 297
rect 480 296 481 297
rect 479 296 480 297
rect 478 296 479 297
rect 477 296 478 297
rect 476 296 477 297
rect 475 296 476 297
rect 474 296 475 297
rect 473 296 474 297
rect 472 296 473 297
rect 471 296 472 297
rect 470 296 471 297
rect 469 296 470 297
rect 468 296 469 297
rect 467 296 468 297
rect 466 296 467 297
rect 465 296 466 297
rect 464 296 465 297
rect 463 296 464 297
rect 462 296 463 297
rect 441 296 442 297
rect 440 296 441 297
rect 419 296 420 297
rect 418 296 419 297
rect 417 296 418 297
rect 416 296 417 297
rect 399 296 400 297
rect 398 296 399 297
rect 397 296 398 297
rect 278 296 279 297
rect 277 296 278 297
rect 276 296 277 297
rect 275 296 276 297
rect 274 296 275 297
rect 273 296 274 297
rect 272 296 273 297
rect 271 296 272 297
rect 270 296 271 297
rect 269 296 270 297
rect 268 296 269 297
rect 267 296 268 297
rect 266 296 267 297
rect 265 296 266 297
rect 264 296 265 297
rect 263 296 264 297
rect 262 296 263 297
rect 261 296 262 297
rect 260 296 261 297
rect 259 296 260 297
rect 258 296 259 297
rect 257 296 258 297
rect 256 296 257 297
rect 255 296 256 297
rect 254 296 255 297
rect 253 296 254 297
rect 252 296 253 297
rect 251 296 252 297
rect 250 296 251 297
rect 249 296 250 297
rect 248 296 249 297
rect 247 296 248 297
rect 246 296 247 297
rect 245 296 246 297
rect 244 296 245 297
rect 243 296 244 297
rect 242 296 243 297
rect 241 296 242 297
rect 240 296 241 297
rect 239 296 240 297
rect 238 296 239 297
rect 237 296 238 297
rect 236 296 237 297
rect 235 296 236 297
rect 234 296 235 297
rect 233 296 234 297
rect 232 296 233 297
rect 231 296 232 297
rect 230 296 231 297
rect 229 296 230 297
rect 228 296 229 297
rect 227 296 228 297
rect 226 296 227 297
rect 225 296 226 297
rect 224 296 225 297
rect 223 296 224 297
rect 222 296 223 297
rect 221 296 222 297
rect 220 296 221 297
rect 219 296 220 297
rect 218 296 219 297
rect 217 296 218 297
rect 216 296 217 297
rect 215 296 216 297
rect 214 296 215 297
rect 190 296 191 297
rect 189 296 190 297
rect 188 296 189 297
rect 187 296 188 297
rect 186 296 187 297
rect 185 296 186 297
rect 184 296 185 297
rect 183 296 184 297
rect 182 296 183 297
rect 181 296 182 297
rect 180 296 181 297
rect 179 296 180 297
rect 178 296 179 297
rect 177 296 178 297
rect 176 296 177 297
rect 175 296 176 297
rect 174 296 175 297
rect 173 296 174 297
rect 172 296 173 297
rect 171 296 172 297
rect 170 296 171 297
rect 169 296 170 297
rect 168 296 169 297
rect 167 296 168 297
rect 166 296 167 297
rect 165 296 166 297
rect 164 296 165 297
rect 163 296 164 297
rect 162 296 163 297
rect 161 296 162 297
rect 160 296 161 297
rect 159 296 160 297
rect 158 296 159 297
rect 157 296 158 297
rect 156 296 157 297
rect 155 296 156 297
rect 154 296 155 297
rect 153 296 154 297
rect 152 296 153 297
rect 151 296 152 297
rect 150 296 151 297
rect 149 296 150 297
rect 148 296 149 297
rect 147 296 148 297
rect 146 296 147 297
rect 145 296 146 297
rect 144 296 145 297
rect 143 296 144 297
rect 142 296 143 297
rect 141 296 142 297
rect 140 296 141 297
rect 121 296 122 297
rect 120 296 121 297
rect 119 296 120 297
rect 118 296 119 297
rect 117 296 118 297
rect 116 296 117 297
rect 115 296 116 297
rect 114 296 115 297
rect 113 296 114 297
rect 112 296 113 297
rect 111 296 112 297
rect 110 296 111 297
rect 109 296 110 297
rect 108 296 109 297
rect 107 296 108 297
rect 106 296 107 297
rect 105 296 106 297
rect 104 296 105 297
rect 103 296 104 297
rect 102 296 103 297
rect 101 296 102 297
rect 100 296 101 297
rect 99 296 100 297
rect 98 296 99 297
rect 97 296 98 297
rect 96 296 97 297
rect 95 296 96 297
rect 94 296 95 297
rect 93 296 94 297
rect 92 296 93 297
rect 91 296 92 297
rect 90 296 91 297
rect 89 296 90 297
rect 88 296 89 297
rect 87 296 88 297
rect 86 296 87 297
rect 70 296 71 297
rect 69 296 70 297
rect 68 296 69 297
rect 67 296 68 297
rect 66 296 67 297
rect 65 296 66 297
rect 64 296 65 297
rect 63 296 64 297
rect 62 296 63 297
rect 61 296 62 297
rect 60 296 61 297
rect 59 296 60 297
rect 58 296 59 297
rect 57 296 58 297
rect 56 296 57 297
rect 55 296 56 297
rect 54 296 55 297
rect 53 296 54 297
rect 52 296 53 297
rect 51 296 52 297
rect 50 296 51 297
rect 49 296 50 297
rect 48 296 49 297
rect 47 296 48 297
rect 46 296 47 297
rect 45 296 46 297
rect 44 296 45 297
rect 43 296 44 297
rect 42 296 43 297
rect 41 296 42 297
rect 31 296 32 297
rect 30 296 31 297
rect 29 296 30 297
rect 28 296 29 297
rect 27 296 28 297
rect 26 296 27 297
rect 25 296 26 297
rect 24 296 25 297
rect 23 296 24 297
rect 22 296 23 297
rect 21 296 22 297
rect 20 296 21 297
rect 19 296 20 297
rect 18 296 19 297
rect 17 296 18 297
rect 16 296 17 297
rect 15 296 16 297
rect 14 296 15 297
rect 13 296 14 297
rect 12 296 13 297
rect 11 296 12 297
rect 10 296 11 297
rect 9 296 10 297
rect 8 296 9 297
rect 7 296 8 297
rect 6 296 7 297
rect 5 296 6 297
rect 482 297 483 298
rect 481 297 482 298
rect 480 297 481 298
rect 479 297 480 298
rect 478 297 479 298
rect 477 297 478 298
rect 476 297 477 298
rect 475 297 476 298
rect 474 297 475 298
rect 473 297 474 298
rect 472 297 473 298
rect 471 297 472 298
rect 470 297 471 298
rect 469 297 470 298
rect 468 297 469 298
rect 467 297 468 298
rect 466 297 467 298
rect 465 297 466 298
rect 464 297 465 298
rect 463 297 464 298
rect 462 297 463 298
rect 419 297 420 298
rect 418 297 419 298
rect 417 297 418 298
rect 416 297 417 298
rect 277 297 278 298
rect 276 297 277 298
rect 275 297 276 298
rect 274 297 275 298
rect 273 297 274 298
rect 272 297 273 298
rect 271 297 272 298
rect 270 297 271 298
rect 269 297 270 298
rect 268 297 269 298
rect 267 297 268 298
rect 266 297 267 298
rect 265 297 266 298
rect 264 297 265 298
rect 263 297 264 298
rect 262 297 263 298
rect 261 297 262 298
rect 260 297 261 298
rect 259 297 260 298
rect 258 297 259 298
rect 257 297 258 298
rect 256 297 257 298
rect 255 297 256 298
rect 254 297 255 298
rect 253 297 254 298
rect 252 297 253 298
rect 251 297 252 298
rect 250 297 251 298
rect 249 297 250 298
rect 248 297 249 298
rect 247 297 248 298
rect 246 297 247 298
rect 245 297 246 298
rect 244 297 245 298
rect 243 297 244 298
rect 242 297 243 298
rect 241 297 242 298
rect 240 297 241 298
rect 239 297 240 298
rect 238 297 239 298
rect 237 297 238 298
rect 236 297 237 298
rect 235 297 236 298
rect 234 297 235 298
rect 233 297 234 298
rect 232 297 233 298
rect 231 297 232 298
rect 230 297 231 298
rect 229 297 230 298
rect 228 297 229 298
rect 227 297 228 298
rect 226 297 227 298
rect 225 297 226 298
rect 224 297 225 298
rect 223 297 224 298
rect 222 297 223 298
rect 221 297 222 298
rect 220 297 221 298
rect 219 297 220 298
rect 218 297 219 298
rect 217 297 218 298
rect 216 297 217 298
rect 215 297 216 298
rect 214 297 215 298
rect 213 297 214 298
rect 189 297 190 298
rect 188 297 189 298
rect 187 297 188 298
rect 186 297 187 298
rect 185 297 186 298
rect 184 297 185 298
rect 183 297 184 298
rect 182 297 183 298
rect 181 297 182 298
rect 180 297 181 298
rect 179 297 180 298
rect 178 297 179 298
rect 177 297 178 298
rect 176 297 177 298
rect 175 297 176 298
rect 174 297 175 298
rect 173 297 174 298
rect 172 297 173 298
rect 171 297 172 298
rect 170 297 171 298
rect 169 297 170 298
rect 168 297 169 298
rect 167 297 168 298
rect 166 297 167 298
rect 165 297 166 298
rect 164 297 165 298
rect 163 297 164 298
rect 162 297 163 298
rect 161 297 162 298
rect 160 297 161 298
rect 159 297 160 298
rect 158 297 159 298
rect 157 297 158 298
rect 156 297 157 298
rect 155 297 156 298
rect 154 297 155 298
rect 153 297 154 298
rect 152 297 153 298
rect 151 297 152 298
rect 150 297 151 298
rect 149 297 150 298
rect 148 297 149 298
rect 147 297 148 298
rect 146 297 147 298
rect 145 297 146 298
rect 144 297 145 298
rect 143 297 144 298
rect 142 297 143 298
rect 141 297 142 298
rect 122 297 123 298
rect 121 297 122 298
rect 120 297 121 298
rect 119 297 120 298
rect 118 297 119 298
rect 117 297 118 298
rect 116 297 117 298
rect 115 297 116 298
rect 114 297 115 298
rect 113 297 114 298
rect 112 297 113 298
rect 111 297 112 298
rect 110 297 111 298
rect 109 297 110 298
rect 108 297 109 298
rect 107 297 108 298
rect 106 297 107 298
rect 105 297 106 298
rect 104 297 105 298
rect 103 297 104 298
rect 102 297 103 298
rect 101 297 102 298
rect 100 297 101 298
rect 99 297 100 298
rect 98 297 99 298
rect 97 297 98 298
rect 96 297 97 298
rect 95 297 96 298
rect 94 297 95 298
rect 93 297 94 298
rect 92 297 93 298
rect 91 297 92 298
rect 90 297 91 298
rect 89 297 90 298
rect 88 297 89 298
rect 87 297 88 298
rect 86 297 87 298
rect 70 297 71 298
rect 69 297 70 298
rect 68 297 69 298
rect 67 297 68 298
rect 66 297 67 298
rect 65 297 66 298
rect 64 297 65 298
rect 63 297 64 298
rect 62 297 63 298
rect 61 297 62 298
rect 60 297 61 298
rect 59 297 60 298
rect 58 297 59 298
rect 57 297 58 298
rect 56 297 57 298
rect 55 297 56 298
rect 54 297 55 298
rect 53 297 54 298
rect 52 297 53 298
rect 51 297 52 298
rect 50 297 51 298
rect 49 297 50 298
rect 48 297 49 298
rect 47 297 48 298
rect 46 297 47 298
rect 45 297 46 298
rect 44 297 45 298
rect 43 297 44 298
rect 42 297 43 298
rect 41 297 42 298
rect 31 297 32 298
rect 30 297 31 298
rect 29 297 30 298
rect 28 297 29 298
rect 27 297 28 298
rect 26 297 27 298
rect 25 297 26 298
rect 24 297 25 298
rect 23 297 24 298
rect 22 297 23 298
rect 21 297 22 298
rect 20 297 21 298
rect 19 297 20 298
rect 18 297 19 298
rect 17 297 18 298
rect 16 297 17 298
rect 15 297 16 298
rect 14 297 15 298
rect 13 297 14 298
rect 12 297 13 298
rect 11 297 12 298
rect 10 297 11 298
rect 9 297 10 298
rect 8 297 9 298
rect 7 297 8 298
rect 6 297 7 298
rect 5 297 6 298
rect 482 298 483 299
rect 481 298 482 299
rect 480 298 481 299
rect 479 298 480 299
rect 478 298 479 299
rect 477 298 478 299
rect 476 298 477 299
rect 475 298 476 299
rect 474 298 475 299
rect 473 298 474 299
rect 472 298 473 299
rect 471 298 472 299
rect 470 298 471 299
rect 469 298 470 299
rect 468 298 469 299
rect 467 298 468 299
rect 466 298 467 299
rect 465 298 466 299
rect 464 298 465 299
rect 463 298 464 299
rect 462 298 463 299
rect 419 298 420 299
rect 418 298 419 299
rect 417 298 418 299
rect 416 298 417 299
rect 275 298 276 299
rect 274 298 275 299
rect 273 298 274 299
rect 272 298 273 299
rect 271 298 272 299
rect 270 298 271 299
rect 269 298 270 299
rect 268 298 269 299
rect 267 298 268 299
rect 266 298 267 299
rect 265 298 266 299
rect 264 298 265 299
rect 263 298 264 299
rect 262 298 263 299
rect 261 298 262 299
rect 260 298 261 299
rect 259 298 260 299
rect 258 298 259 299
rect 257 298 258 299
rect 256 298 257 299
rect 255 298 256 299
rect 254 298 255 299
rect 253 298 254 299
rect 252 298 253 299
rect 251 298 252 299
rect 250 298 251 299
rect 249 298 250 299
rect 248 298 249 299
rect 247 298 248 299
rect 246 298 247 299
rect 245 298 246 299
rect 244 298 245 299
rect 243 298 244 299
rect 242 298 243 299
rect 241 298 242 299
rect 240 298 241 299
rect 239 298 240 299
rect 238 298 239 299
rect 237 298 238 299
rect 236 298 237 299
rect 235 298 236 299
rect 234 298 235 299
rect 233 298 234 299
rect 232 298 233 299
rect 231 298 232 299
rect 230 298 231 299
rect 229 298 230 299
rect 228 298 229 299
rect 227 298 228 299
rect 226 298 227 299
rect 225 298 226 299
rect 224 298 225 299
rect 223 298 224 299
rect 222 298 223 299
rect 221 298 222 299
rect 220 298 221 299
rect 219 298 220 299
rect 218 298 219 299
rect 217 298 218 299
rect 216 298 217 299
rect 215 298 216 299
rect 214 298 215 299
rect 213 298 214 299
rect 188 298 189 299
rect 187 298 188 299
rect 186 298 187 299
rect 185 298 186 299
rect 184 298 185 299
rect 183 298 184 299
rect 182 298 183 299
rect 181 298 182 299
rect 180 298 181 299
rect 179 298 180 299
rect 178 298 179 299
rect 177 298 178 299
rect 176 298 177 299
rect 175 298 176 299
rect 174 298 175 299
rect 173 298 174 299
rect 172 298 173 299
rect 171 298 172 299
rect 170 298 171 299
rect 169 298 170 299
rect 168 298 169 299
rect 167 298 168 299
rect 166 298 167 299
rect 165 298 166 299
rect 164 298 165 299
rect 163 298 164 299
rect 162 298 163 299
rect 161 298 162 299
rect 160 298 161 299
rect 159 298 160 299
rect 158 298 159 299
rect 157 298 158 299
rect 156 298 157 299
rect 155 298 156 299
rect 154 298 155 299
rect 153 298 154 299
rect 152 298 153 299
rect 151 298 152 299
rect 150 298 151 299
rect 149 298 150 299
rect 148 298 149 299
rect 147 298 148 299
rect 146 298 147 299
rect 145 298 146 299
rect 144 298 145 299
rect 143 298 144 299
rect 142 298 143 299
rect 122 298 123 299
rect 121 298 122 299
rect 120 298 121 299
rect 119 298 120 299
rect 118 298 119 299
rect 117 298 118 299
rect 116 298 117 299
rect 115 298 116 299
rect 114 298 115 299
rect 113 298 114 299
rect 112 298 113 299
rect 111 298 112 299
rect 110 298 111 299
rect 109 298 110 299
rect 108 298 109 299
rect 107 298 108 299
rect 106 298 107 299
rect 105 298 106 299
rect 104 298 105 299
rect 103 298 104 299
rect 102 298 103 299
rect 101 298 102 299
rect 100 298 101 299
rect 99 298 100 299
rect 98 298 99 299
rect 97 298 98 299
rect 96 298 97 299
rect 95 298 96 299
rect 94 298 95 299
rect 93 298 94 299
rect 92 298 93 299
rect 91 298 92 299
rect 90 298 91 299
rect 89 298 90 299
rect 88 298 89 299
rect 87 298 88 299
rect 86 298 87 299
rect 70 298 71 299
rect 69 298 70 299
rect 68 298 69 299
rect 67 298 68 299
rect 66 298 67 299
rect 65 298 66 299
rect 64 298 65 299
rect 63 298 64 299
rect 62 298 63 299
rect 61 298 62 299
rect 60 298 61 299
rect 59 298 60 299
rect 58 298 59 299
rect 57 298 58 299
rect 56 298 57 299
rect 55 298 56 299
rect 54 298 55 299
rect 53 298 54 299
rect 52 298 53 299
rect 51 298 52 299
rect 50 298 51 299
rect 49 298 50 299
rect 48 298 49 299
rect 47 298 48 299
rect 46 298 47 299
rect 45 298 46 299
rect 44 298 45 299
rect 43 298 44 299
rect 42 298 43 299
rect 41 298 42 299
rect 31 298 32 299
rect 30 298 31 299
rect 29 298 30 299
rect 28 298 29 299
rect 27 298 28 299
rect 26 298 27 299
rect 25 298 26 299
rect 24 298 25 299
rect 23 298 24 299
rect 22 298 23 299
rect 21 298 22 299
rect 20 298 21 299
rect 19 298 20 299
rect 18 298 19 299
rect 17 298 18 299
rect 16 298 17 299
rect 15 298 16 299
rect 14 298 15 299
rect 13 298 14 299
rect 12 298 13 299
rect 11 298 12 299
rect 10 298 11 299
rect 9 298 10 299
rect 8 298 9 299
rect 7 298 8 299
rect 6 298 7 299
rect 482 299 483 300
rect 462 299 463 300
rect 419 299 420 300
rect 418 299 419 300
rect 417 299 418 300
rect 416 299 417 300
rect 274 299 275 300
rect 273 299 274 300
rect 272 299 273 300
rect 271 299 272 300
rect 270 299 271 300
rect 269 299 270 300
rect 268 299 269 300
rect 267 299 268 300
rect 266 299 267 300
rect 265 299 266 300
rect 264 299 265 300
rect 263 299 264 300
rect 262 299 263 300
rect 261 299 262 300
rect 260 299 261 300
rect 259 299 260 300
rect 258 299 259 300
rect 257 299 258 300
rect 256 299 257 300
rect 255 299 256 300
rect 254 299 255 300
rect 253 299 254 300
rect 252 299 253 300
rect 251 299 252 300
rect 250 299 251 300
rect 249 299 250 300
rect 248 299 249 300
rect 247 299 248 300
rect 246 299 247 300
rect 245 299 246 300
rect 244 299 245 300
rect 243 299 244 300
rect 242 299 243 300
rect 241 299 242 300
rect 240 299 241 300
rect 239 299 240 300
rect 238 299 239 300
rect 237 299 238 300
rect 236 299 237 300
rect 235 299 236 300
rect 234 299 235 300
rect 233 299 234 300
rect 232 299 233 300
rect 231 299 232 300
rect 230 299 231 300
rect 229 299 230 300
rect 228 299 229 300
rect 227 299 228 300
rect 226 299 227 300
rect 225 299 226 300
rect 224 299 225 300
rect 223 299 224 300
rect 222 299 223 300
rect 221 299 222 300
rect 220 299 221 300
rect 219 299 220 300
rect 218 299 219 300
rect 217 299 218 300
rect 216 299 217 300
rect 215 299 216 300
rect 214 299 215 300
rect 213 299 214 300
rect 212 299 213 300
rect 187 299 188 300
rect 186 299 187 300
rect 185 299 186 300
rect 184 299 185 300
rect 183 299 184 300
rect 182 299 183 300
rect 181 299 182 300
rect 180 299 181 300
rect 179 299 180 300
rect 178 299 179 300
rect 177 299 178 300
rect 176 299 177 300
rect 175 299 176 300
rect 174 299 175 300
rect 173 299 174 300
rect 172 299 173 300
rect 171 299 172 300
rect 170 299 171 300
rect 169 299 170 300
rect 168 299 169 300
rect 167 299 168 300
rect 166 299 167 300
rect 165 299 166 300
rect 164 299 165 300
rect 163 299 164 300
rect 162 299 163 300
rect 161 299 162 300
rect 160 299 161 300
rect 159 299 160 300
rect 158 299 159 300
rect 157 299 158 300
rect 156 299 157 300
rect 155 299 156 300
rect 154 299 155 300
rect 153 299 154 300
rect 152 299 153 300
rect 151 299 152 300
rect 150 299 151 300
rect 149 299 150 300
rect 148 299 149 300
rect 147 299 148 300
rect 146 299 147 300
rect 145 299 146 300
rect 144 299 145 300
rect 143 299 144 300
rect 122 299 123 300
rect 121 299 122 300
rect 120 299 121 300
rect 119 299 120 300
rect 118 299 119 300
rect 117 299 118 300
rect 116 299 117 300
rect 115 299 116 300
rect 114 299 115 300
rect 113 299 114 300
rect 112 299 113 300
rect 111 299 112 300
rect 110 299 111 300
rect 109 299 110 300
rect 108 299 109 300
rect 107 299 108 300
rect 106 299 107 300
rect 105 299 106 300
rect 104 299 105 300
rect 103 299 104 300
rect 102 299 103 300
rect 101 299 102 300
rect 100 299 101 300
rect 99 299 100 300
rect 98 299 99 300
rect 97 299 98 300
rect 96 299 97 300
rect 95 299 96 300
rect 94 299 95 300
rect 93 299 94 300
rect 92 299 93 300
rect 91 299 92 300
rect 90 299 91 300
rect 89 299 90 300
rect 88 299 89 300
rect 87 299 88 300
rect 86 299 87 300
rect 70 299 71 300
rect 69 299 70 300
rect 68 299 69 300
rect 67 299 68 300
rect 66 299 67 300
rect 65 299 66 300
rect 64 299 65 300
rect 63 299 64 300
rect 62 299 63 300
rect 61 299 62 300
rect 60 299 61 300
rect 59 299 60 300
rect 58 299 59 300
rect 57 299 58 300
rect 56 299 57 300
rect 55 299 56 300
rect 54 299 55 300
rect 53 299 54 300
rect 52 299 53 300
rect 51 299 52 300
rect 50 299 51 300
rect 49 299 50 300
rect 48 299 49 300
rect 47 299 48 300
rect 46 299 47 300
rect 45 299 46 300
rect 44 299 45 300
rect 43 299 44 300
rect 42 299 43 300
rect 32 299 33 300
rect 31 299 32 300
rect 30 299 31 300
rect 29 299 30 300
rect 28 299 29 300
rect 27 299 28 300
rect 26 299 27 300
rect 25 299 26 300
rect 24 299 25 300
rect 23 299 24 300
rect 22 299 23 300
rect 21 299 22 300
rect 20 299 21 300
rect 19 299 20 300
rect 18 299 19 300
rect 17 299 18 300
rect 16 299 17 300
rect 15 299 16 300
rect 14 299 15 300
rect 13 299 14 300
rect 12 299 13 300
rect 11 299 12 300
rect 10 299 11 300
rect 9 299 10 300
rect 8 299 9 300
rect 7 299 8 300
rect 6 299 7 300
rect 482 300 483 301
rect 462 300 463 301
rect 419 300 420 301
rect 418 300 419 301
rect 417 300 418 301
rect 416 300 417 301
rect 273 300 274 301
rect 272 300 273 301
rect 271 300 272 301
rect 270 300 271 301
rect 269 300 270 301
rect 268 300 269 301
rect 267 300 268 301
rect 266 300 267 301
rect 265 300 266 301
rect 264 300 265 301
rect 263 300 264 301
rect 262 300 263 301
rect 261 300 262 301
rect 260 300 261 301
rect 259 300 260 301
rect 258 300 259 301
rect 257 300 258 301
rect 256 300 257 301
rect 255 300 256 301
rect 254 300 255 301
rect 253 300 254 301
rect 252 300 253 301
rect 251 300 252 301
rect 250 300 251 301
rect 249 300 250 301
rect 248 300 249 301
rect 247 300 248 301
rect 246 300 247 301
rect 245 300 246 301
rect 244 300 245 301
rect 243 300 244 301
rect 242 300 243 301
rect 241 300 242 301
rect 240 300 241 301
rect 239 300 240 301
rect 238 300 239 301
rect 237 300 238 301
rect 236 300 237 301
rect 235 300 236 301
rect 234 300 235 301
rect 233 300 234 301
rect 232 300 233 301
rect 231 300 232 301
rect 230 300 231 301
rect 229 300 230 301
rect 228 300 229 301
rect 227 300 228 301
rect 226 300 227 301
rect 225 300 226 301
rect 224 300 225 301
rect 223 300 224 301
rect 222 300 223 301
rect 221 300 222 301
rect 220 300 221 301
rect 219 300 220 301
rect 218 300 219 301
rect 217 300 218 301
rect 216 300 217 301
rect 215 300 216 301
rect 214 300 215 301
rect 213 300 214 301
rect 212 300 213 301
rect 211 300 212 301
rect 186 300 187 301
rect 185 300 186 301
rect 184 300 185 301
rect 183 300 184 301
rect 182 300 183 301
rect 181 300 182 301
rect 180 300 181 301
rect 179 300 180 301
rect 178 300 179 301
rect 177 300 178 301
rect 176 300 177 301
rect 175 300 176 301
rect 174 300 175 301
rect 173 300 174 301
rect 172 300 173 301
rect 171 300 172 301
rect 170 300 171 301
rect 169 300 170 301
rect 168 300 169 301
rect 167 300 168 301
rect 166 300 167 301
rect 165 300 166 301
rect 164 300 165 301
rect 163 300 164 301
rect 162 300 163 301
rect 161 300 162 301
rect 160 300 161 301
rect 159 300 160 301
rect 158 300 159 301
rect 157 300 158 301
rect 156 300 157 301
rect 155 300 156 301
rect 154 300 155 301
rect 153 300 154 301
rect 152 300 153 301
rect 151 300 152 301
rect 150 300 151 301
rect 149 300 150 301
rect 148 300 149 301
rect 147 300 148 301
rect 146 300 147 301
rect 145 300 146 301
rect 144 300 145 301
rect 123 300 124 301
rect 122 300 123 301
rect 121 300 122 301
rect 120 300 121 301
rect 119 300 120 301
rect 118 300 119 301
rect 117 300 118 301
rect 116 300 117 301
rect 115 300 116 301
rect 114 300 115 301
rect 113 300 114 301
rect 112 300 113 301
rect 111 300 112 301
rect 110 300 111 301
rect 109 300 110 301
rect 108 300 109 301
rect 107 300 108 301
rect 106 300 107 301
rect 105 300 106 301
rect 104 300 105 301
rect 103 300 104 301
rect 102 300 103 301
rect 101 300 102 301
rect 100 300 101 301
rect 99 300 100 301
rect 98 300 99 301
rect 97 300 98 301
rect 96 300 97 301
rect 95 300 96 301
rect 94 300 95 301
rect 93 300 94 301
rect 92 300 93 301
rect 91 300 92 301
rect 90 300 91 301
rect 89 300 90 301
rect 88 300 89 301
rect 87 300 88 301
rect 70 300 71 301
rect 69 300 70 301
rect 68 300 69 301
rect 67 300 68 301
rect 66 300 67 301
rect 65 300 66 301
rect 64 300 65 301
rect 63 300 64 301
rect 62 300 63 301
rect 61 300 62 301
rect 60 300 61 301
rect 59 300 60 301
rect 58 300 59 301
rect 57 300 58 301
rect 56 300 57 301
rect 55 300 56 301
rect 54 300 55 301
rect 53 300 54 301
rect 52 300 53 301
rect 51 300 52 301
rect 50 300 51 301
rect 49 300 50 301
rect 48 300 49 301
rect 47 300 48 301
rect 46 300 47 301
rect 45 300 46 301
rect 44 300 45 301
rect 43 300 44 301
rect 42 300 43 301
rect 32 300 33 301
rect 31 300 32 301
rect 30 300 31 301
rect 29 300 30 301
rect 28 300 29 301
rect 27 300 28 301
rect 26 300 27 301
rect 25 300 26 301
rect 24 300 25 301
rect 23 300 24 301
rect 22 300 23 301
rect 21 300 22 301
rect 20 300 21 301
rect 19 300 20 301
rect 18 300 19 301
rect 17 300 18 301
rect 16 300 17 301
rect 15 300 16 301
rect 14 300 15 301
rect 13 300 14 301
rect 12 300 13 301
rect 11 300 12 301
rect 10 300 11 301
rect 9 300 10 301
rect 8 300 9 301
rect 7 300 8 301
rect 6 300 7 301
rect 482 301 483 302
rect 462 301 463 302
rect 419 301 420 302
rect 418 301 419 302
rect 417 301 418 302
rect 416 301 417 302
rect 272 301 273 302
rect 271 301 272 302
rect 270 301 271 302
rect 269 301 270 302
rect 268 301 269 302
rect 267 301 268 302
rect 266 301 267 302
rect 265 301 266 302
rect 264 301 265 302
rect 263 301 264 302
rect 262 301 263 302
rect 261 301 262 302
rect 260 301 261 302
rect 259 301 260 302
rect 258 301 259 302
rect 257 301 258 302
rect 256 301 257 302
rect 255 301 256 302
rect 254 301 255 302
rect 253 301 254 302
rect 252 301 253 302
rect 251 301 252 302
rect 250 301 251 302
rect 249 301 250 302
rect 248 301 249 302
rect 247 301 248 302
rect 246 301 247 302
rect 245 301 246 302
rect 244 301 245 302
rect 243 301 244 302
rect 242 301 243 302
rect 241 301 242 302
rect 240 301 241 302
rect 239 301 240 302
rect 238 301 239 302
rect 237 301 238 302
rect 236 301 237 302
rect 235 301 236 302
rect 234 301 235 302
rect 233 301 234 302
rect 232 301 233 302
rect 231 301 232 302
rect 230 301 231 302
rect 229 301 230 302
rect 228 301 229 302
rect 227 301 228 302
rect 226 301 227 302
rect 225 301 226 302
rect 224 301 225 302
rect 223 301 224 302
rect 222 301 223 302
rect 221 301 222 302
rect 220 301 221 302
rect 219 301 220 302
rect 218 301 219 302
rect 217 301 218 302
rect 216 301 217 302
rect 215 301 216 302
rect 214 301 215 302
rect 213 301 214 302
rect 212 301 213 302
rect 211 301 212 302
rect 184 301 185 302
rect 183 301 184 302
rect 182 301 183 302
rect 181 301 182 302
rect 180 301 181 302
rect 179 301 180 302
rect 178 301 179 302
rect 177 301 178 302
rect 176 301 177 302
rect 175 301 176 302
rect 174 301 175 302
rect 173 301 174 302
rect 172 301 173 302
rect 171 301 172 302
rect 170 301 171 302
rect 169 301 170 302
rect 168 301 169 302
rect 167 301 168 302
rect 166 301 167 302
rect 165 301 166 302
rect 164 301 165 302
rect 163 301 164 302
rect 162 301 163 302
rect 161 301 162 302
rect 160 301 161 302
rect 159 301 160 302
rect 158 301 159 302
rect 157 301 158 302
rect 156 301 157 302
rect 155 301 156 302
rect 154 301 155 302
rect 153 301 154 302
rect 152 301 153 302
rect 151 301 152 302
rect 150 301 151 302
rect 149 301 150 302
rect 148 301 149 302
rect 147 301 148 302
rect 146 301 147 302
rect 145 301 146 302
rect 123 301 124 302
rect 122 301 123 302
rect 121 301 122 302
rect 120 301 121 302
rect 119 301 120 302
rect 118 301 119 302
rect 117 301 118 302
rect 116 301 117 302
rect 115 301 116 302
rect 114 301 115 302
rect 113 301 114 302
rect 112 301 113 302
rect 111 301 112 302
rect 110 301 111 302
rect 109 301 110 302
rect 108 301 109 302
rect 107 301 108 302
rect 106 301 107 302
rect 105 301 106 302
rect 104 301 105 302
rect 103 301 104 302
rect 102 301 103 302
rect 101 301 102 302
rect 100 301 101 302
rect 99 301 100 302
rect 98 301 99 302
rect 97 301 98 302
rect 96 301 97 302
rect 95 301 96 302
rect 94 301 95 302
rect 93 301 94 302
rect 92 301 93 302
rect 91 301 92 302
rect 90 301 91 302
rect 89 301 90 302
rect 88 301 89 302
rect 87 301 88 302
rect 71 301 72 302
rect 70 301 71 302
rect 69 301 70 302
rect 68 301 69 302
rect 67 301 68 302
rect 66 301 67 302
rect 65 301 66 302
rect 64 301 65 302
rect 63 301 64 302
rect 62 301 63 302
rect 61 301 62 302
rect 60 301 61 302
rect 59 301 60 302
rect 58 301 59 302
rect 57 301 58 302
rect 56 301 57 302
rect 55 301 56 302
rect 54 301 55 302
rect 53 301 54 302
rect 52 301 53 302
rect 51 301 52 302
rect 50 301 51 302
rect 49 301 50 302
rect 48 301 49 302
rect 47 301 48 302
rect 46 301 47 302
rect 45 301 46 302
rect 44 301 45 302
rect 43 301 44 302
rect 42 301 43 302
rect 32 301 33 302
rect 31 301 32 302
rect 30 301 31 302
rect 29 301 30 302
rect 28 301 29 302
rect 27 301 28 302
rect 26 301 27 302
rect 25 301 26 302
rect 24 301 25 302
rect 23 301 24 302
rect 22 301 23 302
rect 21 301 22 302
rect 20 301 21 302
rect 19 301 20 302
rect 18 301 19 302
rect 17 301 18 302
rect 16 301 17 302
rect 15 301 16 302
rect 14 301 15 302
rect 13 301 14 302
rect 12 301 13 302
rect 11 301 12 302
rect 10 301 11 302
rect 9 301 10 302
rect 8 301 9 302
rect 7 301 8 302
rect 463 302 464 303
rect 462 302 463 303
rect 419 302 420 303
rect 418 302 419 303
rect 417 302 418 303
rect 416 302 417 303
rect 271 302 272 303
rect 270 302 271 303
rect 269 302 270 303
rect 268 302 269 303
rect 267 302 268 303
rect 266 302 267 303
rect 265 302 266 303
rect 264 302 265 303
rect 263 302 264 303
rect 262 302 263 303
rect 261 302 262 303
rect 260 302 261 303
rect 259 302 260 303
rect 258 302 259 303
rect 257 302 258 303
rect 256 302 257 303
rect 255 302 256 303
rect 254 302 255 303
rect 253 302 254 303
rect 252 302 253 303
rect 251 302 252 303
rect 250 302 251 303
rect 249 302 250 303
rect 248 302 249 303
rect 247 302 248 303
rect 246 302 247 303
rect 245 302 246 303
rect 244 302 245 303
rect 243 302 244 303
rect 242 302 243 303
rect 241 302 242 303
rect 240 302 241 303
rect 239 302 240 303
rect 238 302 239 303
rect 237 302 238 303
rect 236 302 237 303
rect 235 302 236 303
rect 234 302 235 303
rect 233 302 234 303
rect 232 302 233 303
rect 231 302 232 303
rect 230 302 231 303
rect 229 302 230 303
rect 228 302 229 303
rect 227 302 228 303
rect 226 302 227 303
rect 225 302 226 303
rect 224 302 225 303
rect 223 302 224 303
rect 222 302 223 303
rect 221 302 222 303
rect 220 302 221 303
rect 219 302 220 303
rect 218 302 219 303
rect 217 302 218 303
rect 216 302 217 303
rect 215 302 216 303
rect 214 302 215 303
rect 213 302 214 303
rect 212 302 213 303
rect 211 302 212 303
rect 210 302 211 303
rect 183 302 184 303
rect 182 302 183 303
rect 181 302 182 303
rect 180 302 181 303
rect 179 302 180 303
rect 178 302 179 303
rect 177 302 178 303
rect 176 302 177 303
rect 175 302 176 303
rect 174 302 175 303
rect 173 302 174 303
rect 172 302 173 303
rect 171 302 172 303
rect 170 302 171 303
rect 169 302 170 303
rect 168 302 169 303
rect 167 302 168 303
rect 166 302 167 303
rect 165 302 166 303
rect 164 302 165 303
rect 163 302 164 303
rect 162 302 163 303
rect 161 302 162 303
rect 160 302 161 303
rect 159 302 160 303
rect 158 302 159 303
rect 157 302 158 303
rect 156 302 157 303
rect 155 302 156 303
rect 154 302 155 303
rect 153 302 154 303
rect 152 302 153 303
rect 151 302 152 303
rect 150 302 151 303
rect 149 302 150 303
rect 148 302 149 303
rect 147 302 148 303
rect 146 302 147 303
rect 123 302 124 303
rect 122 302 123 303
rect 121 302 122 303
rect 120 302 121 303
rect 119 302 120 303
rect 118 302 119 303
rect 117 302 118 303
rect 116 302 117 303
rect 115 302 116 303
rect 114 302 115 303
rect 113 302 114 303
rect 112 302 113 303
rect 111 302 112 303
rect 110 302 111 303
rect 109 302 110 303
rect 108 302 109 303
rect 107 302 108 303
rect 106 302 107 303
rect 105 302 106 303
rect 104 302 105 303
rect 103 302 104 303
rect 102 302 103 303
rect 101 302 102 303
rect 100 302 101 303
rect 99 302 100 303
rect 98 302 99 303
rect 97 302 98 303
rect 96 302 97 303
rect 95 302 96 303
rect 94 302 95 303
rect 93 302 94 303
rect 92 302 93 303
rect 91 302 92 303
rect 90 302 91 303
rect 89 302 90 303
rect 88 302 89 303
rect 87 302 88 303
rect 71 302 72 303
rect 70 302 71 303
rect 69 302 70 303
rect 68 302 69 303
rect 67 302 68 303
rect 66 302 67 303
rect 65 302 66 303
rect 64 302 65 303
rect 63 302 64 303
rect 62 302 63 303
rect 61 302 62 303
rect 60 302 61 303
rect 59 302 60 303
rect 58 302 59 303
rect 57 302 58 303
rect 56 302 57 303
rect 55 302 56 303
rect 54 302 55 303
rect 53 302 54 303
rect 52 302 53 303
rect 51 302 52 303
rect 50 302 51 303
rect 49 302 50 303
rect 48 302 49 303
rect 47 302 48 303
rect 46 302 47 303
rect 45 302 46 303
rect 44 302 45 303
rect 43 302 44 303
rect 42 302 43 303
rect 32 302 33 303
rect 31 302 32 303
rect 30 302 31 303
rect 29 302 30 303
rect 28 302 29 303
rect 27 302 28 303
rect 26 302 27 303
rect 25 302 26 303
rect 24 302 25 303
rect 23 302 24 303
rect 22 302 23 303
rect 21 302 22 303
rect 20 302 21 303
rect 19 302 20 303
rect 18 302 19 303
rect 17 302 18 303
rect 16 302 17 303
rect 15 302 16 303
rect 14 302 15 303
rect 13 302 14 303
rect 12 302 13 303
rect 11 302 12 303
rect 10 302 11 303
rect 9 302 10 303
rect 8 302 9 303
rect 7 302 8 303
rect 464 303 465 304
rect 463 303 464 304
rect 462 303 463 304
rect 419 303 420 304
rect 418 303 419 304
rect 417 303 418 304
rect 416 303 417 304
rect 270 303 271 304
rect 269 303 270 304
rect 268 303 269 304
rect 267 303 268 304
rect 266 303 267 304
rect 265 303 266 304
rect 264 303 265 304
rect 263 303 264 304
rect 262 303 263 304
rect 261 303 262 304
rect 260 303 261 304
rect 259 303 260 304
rect 258 303 259 304
rect 257 303 258 304
rect 256 303 257 304
rect 255 303 256 304
rect 254 303 255 304
rect 253 303 254 304
rect 252 303 253 304
rect 251 303 252 304
rect 250 303 251 304
rect 249 303 250 304
rect 248 303 249 304
rect 247 303 248 304
rect 246 303 247 304
rect 245 303 246 304
rect 244 303 245 304
rect 243 303 244 304
rect 242 303 243 304
rect 241 303 242 304
rect 240 303 241 304
rect 239 303 240 304
rect 238 303 239 304
rect 237 303 238 304
rect 236 303 237 304
rect 235 303 236 304
rect 234 303 235 304
rect 233 303 234 304
rect 232 303 233 304
rect 231 303 232 304
rect 230 303 231 304
rect 229 303 230 304
rect 228 303 229 304
rect 227 303 228 304
rect 226 303 227 304
rect 225 303 226 304
rect 224 303 225 304
rect 223 303 224 304
rect 222 303 223 304
rect 221 303 222 304
rect 220 303 221 304
rect 219 303 220 304
rect 218 303 219 304
rect 217 303 218 304
rect 216 303 217 304
rect 215 303 216 304
rect 214 303 215 304
rect 213 303 214 304
rect 212 303 213 304
rect 211 303 212 304
rect 210 303 211 304
rect 209 303 210 304
rect 182 303 183 304
rect 181 303 182 304
rect 180 303 181 304
rect 179 303 180 304
rect 178 303 179 304
rect 177 303 178 304
rect 176 303 177 304
rect 175 303 176 304
rect 174 303 175 304
rect 173 303 174 304
rect 172 303 173 304
rect 171 303 172 304
rect 170 303 171 304
rect 169 303 170 304
rect 168 303 169 304
rect 167 303 168 304
rect 166 303 167 304
rect 165 303 166 304
rect 164 303 165 304
rect 163 303 164 304
rect 162 303 163 304
rect 161 303 162 304
rect 160 303 161 304
rect 159 303 160 304
rect 158 303 159 304
rect 157 303 158 304
rect 156 303 157 304
rect 155 303 156 304
rect 154 303 155 304
rect 153 303 154 304
rect 152 303 153 304
rect 151 303 152 304
rect 150 303 151 304
rect 149 303 150 304
rect 148 303 149 304
rect 124 303 125 304
rect 123 303 124 304
rect 122 303 123 304
rect 121 303 122 304
rect 120 303 121 304
rect 119 303 120 304
rect 118 303 119 304
rect 117 303 118 304
rect 116 303 117 304
rect 115 303 116 304
rect 114 303 115 304
rect 113 303 114 304
rect 112 303 113 304
rect 111 303 112 304
rect 110 303 111 304
rect 109 303 110 304
rect 108 303 109 304
rect 107 303 108 304
rect 106 303 107 304
rect 105 303 106 304
rect 104 303 105 304
rect 103 303 104 304
rect 102 303 103 304
rect 101 303 102 304
rect 100 303 101 304
rect 99 303 100 304
rect 98 303 99 304
rect 97 303 98 304
rect 96 303 97 304
rect 95 303 96 304
rect 94 303 95 304
rect 93 303 94 304
rect 92 303 93 304
rect 91 303 92 304
rect 90 303 91 304
rect 89 303 90 304
rect 88 303 89 304
rect 87 303 88 304
rect 71 303 72 304
rect 70 303 71 304
rect 69 303 70 304
rect 68 303 69 304
rect 67 303 68 304
rect 66 303 67 304
rect 65 303 66 304
rect 64 303 65 304
rect 63 303 64 304
rect 62 303 63 304
rect 61 303 62 304
rect 60 303 61 304
rect 59 303 60 304
rect 58 303 59 304
rect 57 303 58 304
rect 56 303 57 304
rect 55 303 56 304
rect 54 303 55 304
rect 53 303 54 304
rect 52 303 53 304
rect 51 303 52 304
rect 50 303 51 304
rect 49 303 50 304
rect 48 303 49 304
rect 47 303 48 304
rect 46 303 47 304
rect 45 303 46 304
rect 44 303 45 304
rect 43 303 44 304
rect 32 303 33 304
rect 31 303 32 304
rect 30 303 31 304
rect 29 303 30 304
rect 28 303 29 304
rect 27 303 28 304
rect 26 303 27 304
rect 25 303 26 304
rect 24 303 25 304
rect 23 303 24 304
rect 22 303 23 304
rect 21 303 22 304
rect 20 303 21 304
rect 19 303 20 304
rect 18 303 19 304
rect 17 303 18 304
rect 16 303 17 304
rect 15 303 16 304
rect 14 303 15 304
rect 13 303 14 304
rect 12 303 13 304
rect 11 303 12 304
rect 10 303 11 304
rect 9 303 10 304
rect 8 303 9 304
rect 7 303 8 304
rect 466 304 467 305
rect 465 304 466 305
rect 464 304 465 305
rect 463 304 464 305
rect 462 304 463 305
rect 461 304 462 305
rect 441 304 442 305
rect 440 304 441 305
rect 419 304 420 305
rect 418 304 419 305
rect 417 304 418 305
rect 416 304 417 305
rect 398 304 399 305
rect 397 304 398 305
rect 268 304 269 305
rect 267 304 268 305
rect 266 304 267 305
rect 265 304 266 305
rect 264 304 265 305
rect 263 304 264 305
rect 262 304 263 305
rect 261 304 262 305
rect 260 304 261 305
rect 259 304 260 305
rect 258 304 259 305
rect 257 304 258 305
rect 256 304 257 305
rect 255 304 256 305
rect 254 304 255 305
rect 253 304 254 305
rect 252 304 253 305
rect 251 304 252 305
rect 250 304 251 305
rect 249 304 250 305
rect 248 304 249 305
rect 247 304 248 305
rect 246 304 247 305
rect 245 304 246 305
rect 244 304 245 305
rect 243 304 244 305
rect 242 304 243 305
rect 241 304 242 305
rect 240 304 241 305
rect 239 304 240 305
rect 238 304 239 305
rect 237 304 238 305
rect 236 304 237 305
rect 235 304 236 305
rect 234 304 235 305
rect 233 304 234 305
rect 232 304 233 305
rect 231 304 232 305
rect 230 304 231 305
rect 229 304 230 305
rect 228 304 229 305
rect 227 304 228 305
rect 226 304 227 305
rect 225 304 226 305
rect 224 304 225 305
rect 223 304 224 305
rect 222 304 223 305
rect 221 304 222 305
rect 220 304 221 305
rect 219 304 220 305
rect 218 304 219 305
rect 217 304 218 305
rect 216 304 217 305
rect 215 304 216 305
rect 214 304 215 305
rect 213 304 214 305
rect 212 304 213 305
rect 211 304 212 305
rect 210 304 211 305
rect 209 304 210 305
rect 180 304 181 305
rect 179 304 180 305
rect 178 304 179 305
rect 177 304 178 305
rect 176 304 177 305
rect 175 304 176 305
rect 174 304 175 305
rect 173 304 174 305
rect 172 304 173 305
rect 171 304 172 305
rect 170 304 171 305
rect 169 304 170 305
rect 168 304 169 305
rect 167 304 168 305
rect 166 304 167 305
rect 165 304 166 305
rect 164 304 165 305
rect 163 304 164 305
rect 162 304 163 305
rect 161 304 162 305
rect 160 304 161 305
rect 159 304 160 305
rect 158 304 159 305
rect 157 304 158 305
rect 156 304 157 305
rect 155 304 156 305
rect 154 304 155 305
rect 153 304 154 305
rect 152 304 153 305
rect 151 304 152 305
rect 150 304 151 305
rect 149 304 150 305
rect 124 304 125 305
rect 123 304 124 305
rect 122 304 123 305
rect 121 304 122 305
rect 120 304 121 305
rect 119 304 120 305
rect 118 304 119 305
rect 117 304 118 305
rect 116 304 117 305
rect 115 304 116 305
rect 114 304 115 305
rect 113 304 114 305
rect 112 304 113 305
rect 111 304 112 305
rect 110 304 111 305
rect 109 304 110 305
rect 108 304 109 305
rect 107 304 108 305
rect 106 304 107 305
rect 105 304 106 305
rect 104 304 105 305
rect 103 304 104 305
rect 102 304 103 305
rect 101 304 102 305
rect 100 304 101 305
rect 99 304 100 305
rect 98 304 99 305
rect 97 304 98 305
rect 96 304 97 305
rect 95 304 96 305
rect 94 304 95 305
rect 93 304 94 305
rect 92 304 93 305
rect 91 304 92 305
rect 90 304 91 305
rect 89 304 90 305
rect 88 304 89 305
rect 71 304 72 305
rect 70 304 71 305
rect 69 304 70 305
rect 68 304 69 305
rect 67 304 68 305
rect 66 304 67 305
rect 65 304 66 305
rect 64 304 65 305
rect 63 304 64 305
rect 62 304 63 305
rect 61 304 62 305
rect 60 304 61 305
rect 59 304 60 305
rect 58 304 59 305
rect 57 304 58 305
rect 56 304 57 305
rect 55 304 56 305
rect 54 304 55 305
rect 53 304 54 305
rect 52 304 53 305
rect 51 304 52 305
rect 50 304 51 305
rect 49 304 50 305
rect 48 304 49 305
rect 47 304 48 305
rect 46 304 47 305
rect 45 304 46 305
rect 44 304 45 305
rect 43 304 44 305
rect 32 304 33 305
rect 31 304 32 305
rect 30 304 31 305
rect 29 304 30 305
rect 28 304 29 305
rect 27 304 28 305
rect 26 304 27 305
rect 25 304 26 305
rect 24 304 25 305
rect 23 304 24 305
rect 22 304 23 305
rect 21 304 22 305
rect 20 304 21 305
rect 19 304 20 305
rect 18 304 19 305
rect 17 304 18 305
rect 16 304 17 305
rect 15 304 16 305
rect 14 304 15 305
rect 13 304 14 305
rect 12 304 13 305
rect 11 304 12 305
rect 10 304 11 305
rect 9 304 10 305
rect 8 304 9 305
rect 466 305 467 306
rect 465 305 466 306
rect 464 305 465 306
rect 463 305 464 306
rect 462 305 463 306
rect 461 305 462 306
rect 441 305 442 306
rect 440 305 441 306
rect 439 305 440 306
rect 419 305 420 306
rect 418 305 419 306
rect 417 305 418 306
rect 416 305 417 306
rect 399 305 400 306
rect 398 305 399 306
rect 397 305 398 306
rect 267 305 268 306
rect 266 305 267 306
rect 265 305 266 306
rect 264 305 265 306
rect 263 305 264 306
rect 262 305 263 306
rect 261 305 262 306
rect 260 305 261 306
rect 259 305 260 306
rect 258 305 259 306
rect 257 305 258 306
rect 256 305 257 306
rect 255 305 256 306
rect 254 305 255 306
rect 253 305 254 306
rect 252 305 253 306
rect 251 305 252 306
rect 250 305 251 306
rect 249 305 250 306
rect 248 305 249 306
rect 247 305 248 306
rect 246 305 247 306
rect 245 305 246 306
rect 244 305 245 306
rect 243 305 244 306
rect 242 305 243 306
rect 241 305 242 306
rect 240 305 241 306
rect 239 305 240 306
rect 238 305 239 306
rect 237 305 238 306
rect 236 305 237 306
rect 235 305 236 306
rect 234 305 235 306
rect 233 305 234 306
rect 232 305 233 306
rect 231 305 232 306
rect 230 305 231 306
rect 229 305 230 306
rect 228 305 229 306
rect 227 305 228 306
rect 226 305 227 306
rect 225 305 226 306
rect 224 305 225 306
rect 223 305 224 306
rect 222 305 223 306
rect 221 305 222 306
rect 220 305 221 306
rect 219 305 220 306
rect 218 305 219 306
rect 217 305 218 306
rect 216 305 217 306
rect 215 305 216 306
rect 214 305 215 306
rect 213 305 214 306
rect 212 305 213 306
rect 211 305 212 306
rect 210 305 211 306
rect 209 305 210 306
rect 208 305 209 306
rect 179 305 180 306
rect 178 305 179 306
rect 177 305 178 306
rect 176 305 177 306
rect 175 305 176 306
rect 174 305 175 306
rect 173 305 174 306
rect 172 305 173 306
rect 171 305 172 306
rect 170 305 171 306
rect 169 305 170 306
rect 168 305 169 306
rect 167 305 168 306
rect 166 305 167 306
rect 165 305 166 306
rect 164 305 165 306
rect 163 305 164 306
rect 162 305 163 306
rect 161 305 162 306
rect 160 305 161 306
rect 159 305 160 306
rect 158 305 159 306
rect 157 305 158 306
rect 156 305 157 306
rect 155 305 156 306
rect 154 305 155 306
rect 153 305 154 306
rect 152 305 153 306
rect 151 305 152 306
rect 125 305 126 306
rect 124 305 125 306
rect 123 305 124 306
rect 122 305 123 306
rect 121 305 122 306
rect 120 305 121 306
rect 119 305 120 306
rect 118 305 119 306
rect 117 305 118 306
rect 116 305 117 306
rect 115 305 116 306
rect 114 305 115 306
rect 113 305 114 306
rect 112 305 113 306
rect 111 305 112 306
rect 110 305 111 306
rect 109 305 110 306
rect 108 305 109 306
rect 107 305 108 306
rect 106 305 107 306
rect 105 305 106 306
rect 104 305 105 306
rect 103 305 104 306
rect 102 305 103 306
rect 101 305 102 306
rect 100 305 101 306
rect 99 305 100 306
rect 98 305 99 306
rect 97 305 98 306
rect 96 305 97 306
rect 95 305 96 306
rect 94 305 95 306
rect 93 305 94 306
rect 92 305 93 306
rect 91 305 92 306
rect 90 305 91 306
rect 89 305 90 306
rect 88 305 89 306
rect 72 305 73 306
rect 71 305 72 306
rect 70 305 71 306
rect 69 305 70 306
rect 68 305 69 306
rect 67 305 68 306
rect 66 305 67 306
rect 65 305 66 306
rect 64 305 65 306
rect 63 305 64 306
rect 62 305 63 306
rect 61 305 62 306
rect 60 305 61 306
rect 59 305 60 306
rect 58 305 59 306
rect 57 305 58 306
rect 56 305 57 306
rect 55 305 56 306
rect 54 305 55 306
rect 53 305 54 306
rect 52 305 53 306
rect 51 305 52 306
rect 50 305 51 306
rect 49 305 50 306
rect 48 305 49 306
rect 47 305 48 306
rect 46 305 47 306
rect 45 305 46 306
rect 44 305 45 306
rect 43 305 44 306
rect 33 305 34 306
rect 32 305 33 306
rect 31 305 32 306
rect 30 305 31 306
rect 29 305 30 306
rect 28 305 29 306
rect 27 305 28 306
rect 26 305 27 306
rect 25 305 26 306
rect 24 305 25 306
rect 23 305 24 306
rect 22 305 23 306
rect 21 305 22 306
rect 20 305 21 306
rect 19 305 20 306
rect 18 305 19 306
rect 17 305 18 306
rect 16 305 17 306
rect 15 305 16 306
rect 14 305 15 306
rect 13 305 14 306
rect 12 305 13 306
rect 11 305 12 306
rect 10 305 11 306
rect 9 305 10 306
rect 8 305 9 306
rect 441 306 442 307
rect 440 306 441 307
rect 439 306 440 307
rect 419 306 420 307
rect 418 306 419 307
rect 417 306 418 307
rect 416 306 417 307
rect 399 306 400 307
rect 398 306 399 307
rect 397 306 398 307
rect 266 306 267 307
rect 265 306 266 307
rect 264 306 265 307
rect 263 306 264 307
rect 262 306 263 307
rect 261 306 262 307
rect 260 306 261 307
rect 259 306 260 307
rect 258 306 259 307
rect 257 306 258 307
rect 256 306 257 307
rect 255 306 256 307
rect 254 306 255 307
rect 253 306 254 307
rect 252 306 253 307
rect 251 306 252 307
rect 250 306 251 307
rect 249 306 250 307
rect 248 306 249 307
rect 247 306 248 307
rect 246 306 247 307
rect 245 306 246 307
rect 244 306 245 307
rect 243 306 244 307
rect 242 306 243 307
rect 241 306 242 307
rect 240 306 241 307
rect 239 306 240 307
rect 238 306 239 307
rect 237 306 238 307
rect 236 306 237 307
rect 235 306 236 307
rect 234 306 235 307
rect 233 306 234 307
rect 232 306 233 307
rect 231 306 232 307
rect 230 306 231 307
rect 229 306 230 307
rect 228 306 229 307
rect 227 306 228 307
rect 226 306 227 307
rect 225 306 226 307
rect 224 306 225 307
rect 223 306 224 307
rect 222 306 223 307
rect 221 306 222 307
rect 220 306 221 307
rect 219 306 220 307
rect 218 306 219 307
rect 217 306 218 307
rect 216 306 217 307
rect 215 306 216 307
rect 214 306 215 307
rect 213 306 214 307
rect 212 306 213 307
rect 211 306 212 307
rect 210 306 211 307
rect 209 306 210 307
rect 208 306 209 307
rect 207 306 208 307
rect 177 306 178 307
rect 176 306 177 307
rect 175 306 176 307
rect 174 306 175 307
rect 173 306 174 307
rect 172 306 173 307
rect 171 306 172 307
rect 170 306 171 307
rect 169 306 170 307
rect 168 306 169 307
rect 167 306 168 307
rect 166 306 167 307
rect 165 306 166 307
rect 164 306 165 307
rect 163 306 164 307
rect 162 306 163 307
rect 161 306 162 307
rect 160 306 161 307
rect 159 306 160 307
rect 158 306 159 307
rect 157 306 158 307
rect 156 306 157 307
rect 155 306 156 307
rect 154 306 155 307
rect 153 306 154 307
rect 125 306 126 307
rect 124 306 125 307
rect 123 306 124 307
rect 122 306 123 307
rect 121 306 122 307
rect 120 306 121 307
rect 119 306 120 307
rect 118 306 119 307
rect 117 306 118 307
rect 116 306 117 307
rect 115 306 116 307
rect 114 306 115 307
rect 113 306 114 307
rect 112 306 113 307
rect 111 306 112 307
rect 110 306 111 307
rect 109 306 110 307
rect 108 306 109 307
rect 107 306 108 307
rect 106 306 107 307
rect 105 306 106 307
rect 104 306 105 307
rect 103 306 104 307
rect 102 306 103 307
rect 101 306 102 307
rect 100 306 101 307
rect 99 306 100 307
rect 98 306 99 307
rect 97 306 98 307
rect 96 306 97 307
rect 95 306 96 307
rect 94 306 95 307
rect 93 306 94 307
rect 92 306 93 307
rect 91 306 92 307
rect 90 306 91 307
rect 89 306 90 307
rect 88 306 89 307
rect 72 306 73 307
rect 71 306 72 307
rect 70 306 71 307
rect 69 306 70 307
rect 68 306 69 307
rect 67 306 68 307
rect 66 306 67 307
rect 65 306 66 307
rect 64 306 65 307
rect 63 306 64 307
rect 62 306 63 307
rect 61 306 62 307
rect 60 306 61 307
rect 59 306 60 307
rect 58 306 59 307
rect 57 306 58 307
rect 56 306 57 307
rect 55 306 56 307
rect 54 306 55 307
rect 53 306 54 307
rect 52 306 53 307
rect 51 306 52 307
rect 50 306 51 307
rect 49 306 50 307
rect 48 306 49 307
rect 47 306 48 307
rect 46 306 47 307
rect 45 306 46 307
rect 44 306 45 307
rect 33 306 34 307
rect 32 306 33 307
rect 31 306 32 307
rect 30 306 31 307
rect 29 306 30 307
rect 28 306 29 307
rect 27 306 28 307
rect 26 306 27 307
rect 25 306 26 307
rect 24 306 25 307
rect 23 306 24 307
rect 22 306 23 307
rect 21 306 22 307
rect 20 306 21 307
rect 19 306 20 307
rect 18 306 19 307
rect 17 306 18 307
rect 16 306 17 307
rect 15 306 16 307
rect 14 306 15 307
rect 13 306 14 307
rect 12 306 13 307
rect 11 306 12 307
rect 10 306 11 307
rect 9 306 10 307
rect 441 307 442 308
rect 440 307 441 308
rect 439 307 440 308
rect 419 307 420 308
rect 418 307 419 308
rect 417 307 418 308
rect 416 307 417 308
rect 399 307 400 308
rect 398 307 399 308
rect 397 307 398 308
rect 264 307 265 308
rect 263 307 264 308
rect 262 307 263 308
rect 261 307 262 308
rect 260 307 261 308
rect 259 307 260 308
rect 258 307 259 308
rect 257 307 258 308
rect 256 307 257 308
rect 255 307 256 308
rect 254 307 255 308
rect 253 307 254 308
rect 252 307 253 308
rect 251 307 252 308
rect 250 307 251 308
rect 249 307 250 308
rect 248 307 249 308
rect 247 307 248 308
rect 246 307 247 308
rect 245 307 246 308
rect 244 307 245 308
rect 243 307 244 308
rect 242 307 243 308
rect 241 307 242 308
rect 240 307 241 308
rect 239 307 240 308
rect 238 307 239 308
rect 237 307 238 308
rect 236 307 237 308
rect 235 307 236 308
rect 234 307 235 308
rect 233 307 234 308
rect 232 307 233 308
rect 231 307 232 308
rect 230 307 231 308
rect 229 307 230 308
rect 228 307 229 308
rect 227 307 228 308
rect 226 307 227 308
rect 225 307 226 308
rect 224 307 225 308
rect 223 307 224 308
rect 222 307 223 308
rect 221 307 222 308
rect 220 307 221 308
rect 219 307 220 308
rect 218 307 219 308
rect 217 307 218 308
rect 216 307 217 308
rect 215 307 216 308
rect 214 307 215 308
rect 213 307 214 308
rect 212 307 213 308
rect 211 307 212 308
rect 210 307 211 308
rect 209 307 210 308
rect 208 307 209 308
rect 207 307 208 308
rect 206 307 207 308
rect 175 307 176 308
rect 174 307 175 308
rect 173 307 174 308
rect 172 307 173 308
rect 171 307 172 308
rect 170 307 171 308
rect 169 307 170 308
rect 168 307 169 308
rect 167 307 168 308
rect 166 307 167 308
rect 165 307 166 308
rect 164 307 165 308
rect 163 307 164 308
rect 162 307 163 308
rect 161 307 162 308
rect 160 307 161 308
rect 159 307 160 308
rect 158 307 159 308
rect 157 307 158 308
rect 156 307 157 308
rect 155 307 156 308
rect 126 307 127 308
rect 125 307 126 308
rect 124 307 125 308
rect 123 307 124 308
rect 122 307 123 308
rect 121 307 122 308
rect 120 307 121 308
rect 119 307 120 308
rect 118 307 119 308
rect 117 307 118 308
rect 116 307 117 308
rect 115 307 116 308
rect 114 307 115 308
rect 113 307 114 308
rect 112 307 113 308
rect 111 307 112 308
rect 110 307 111 308
rect 109 307 110 308
rect 108 307 109 308
rect 107 307 108 308
rect 106 307 107 308
rect 105 307 106 308
rect 104 307 105 308
rect 103 307 104 308
rect 102 307 103 308
rect 101 307 102 308
rect 100 307 101 308
rect 99 307 100 308
rect 98 307 99 308
rect 97 307 98 308
rect 96 307 97 308
rect 95 307 96 308
rect 94 307 95 308
rect 93 307 94 308
rect 92 307 93 308
rect 91 307 92 308
rect 90 307 91 308
rect 89 307 90 308
rect 72 307 73 308
rect 71 307 72 308
rect 70 307 71 308
rect 69 307 70 308
rect 68 307 69 308
rect 67 307 68 308
rect 66 307 67 308
rect 65 307 66 308
rect 64 307 65 308
rect 63 307 64 308
rect 62 307 63 308
rect 61 307 62 308
rect 60 307 61 308
rect 59 307 60 308
rect 58 307 59 308
rect 57 307 58 308
rect 56 307 57 308
rect 55 307 56 308
rect 54 307 55 308
rect 53 307 54 308
rect 52 307 53 308
rect 51 307 52 308
rect 50 307 51 308
rect 49 307 50 308
rect 48 307 49 308
rect 47 307 48 308
rect 46 307 47 308
rect 45 307 46 308
rect 44 307 45 308
rect 33 307 34 308
rect 32 307 33 308
rect 31 307 32 308
rect 30 307 31 308
rect 29 307 30 308
rect 28 307 29 308
rect 27 307 28 308
rect 26 307 27 308
rect 25 307 26 308
rect 24 307 25 308
rect 23 307 24 308
rect 22 307 23 308
rect 21 307 22 308
rect 20 307 21 308
rect 19 307 20 308
rect 18 307 19 308
rect 17 307 18 308
rect 16 307 17 308
rect 15 307 16 308
rect 14 307 15 308
rect 13 307 14 308
rect 12 307 13 308
rect 11 307 12 308
rect 10 307 11 308
rect 9 307 10 308
rect 441 308 442 309
rect 440 308 441 309
rect 439 308 440 309
rect 419 308 420 309
rect 418 308 419 309
rect 417 308 418 309
rect 416 308 417 309
rect 399 308 400 309
rect 398 308 399 309
rect 397 308 398 309
rect 263 308 264 309
rect 262 308 263 309
rect 261 308 262 309
rect 260 308 261 309
rect 259 308 260 309
rect 258 308 259 309
rect 257 308 258 309
rect 256 308 257 309
rect 255 308 256 309
rect 254 308 255 309
rect 253 308 254 309
rect 252 308 253 309
rect 251 308 252 309
rect 250 308 251 309
rect 249 308 250 309
rect 248 308 249 309
rect 247 308 248 309
rect 246 308 247 309
rect 245 308 246 309
rect 244 308 245 309
rect 243 308 244 309
rect 242 308 243 309
rect 241 308 242 309
rect 240 308 241 309
rect 239 308 240 309
rect 238 308 239 309
rect 237 308 238 309
rect 236 308 237 309
rect 235 308 236 309
rect 234 308 235 309
rect 233 308 234 309
rect 232 308 233 309
rect 231 308 232 309
rect 230 308 231 309
rect 229 308 230 309
rect 228 308 229 309
rect 227 308 228 309
rect 226 308 227 309
rect 225 308 226 309
rect 224 308 225 309
rect 223 308 224 309
rect 222 308 223 309
rect 221 308 222 309
rect 220 308 221 309
rect 219 308 220 309
rect 218 308 219 309
rect 217 308 218 309
rect 216 308 217 309
rect 215 308 216 309
rect 214 308 215 309
rect 213 308 214 309
rect 212 308 213 309
rect 211 308 212 309
rect 210 308 211 309
rect 209 308 210 309
rect 208 308 209 309
rect 207 308 208 309
rect 206 308 207 309
rect 205 308 206 309
rect 172 308 173 309
rect 171 308 172 309
rect 170 308 171 309
rect 169 308 170 309
rect 168 308 169 309
rect 167 308 168 309
rect 166 308 167 309
rect 165 308 166 309
rect 164 308 165 309
rect 163 308 164 309
rect 162 308 163 309
rect 161 308 162 309
rect 160 308 161 309
rect 159 308 160 309
rect 158 308 159 309
rect 127 308 128 309
rect 126 308 127 309
rect 125 308 126 309
rect 124 308 125 309
rect 123 308 124 309
rect 122 308 123 309
rect 121 308 122 309
rect 120 308 121 309
rect 119 308 120 309
rect 118 308 119 309
rect 117 308 118 309
rect 116 308 117 309
rect 115 308 116 309
rect 114 308 115 309
rect 113 308 114 309
rect 112 308 113 309
rect 111 308 112 309
rect 110 308 111 309
rect 109 308 110 309
rect 108 308 109 309
rect 107 308 108 309
rect 106 308 107 309
rect 105 308 106 309
rect 104 308 105 309
rect 103 308 104 309
rect 102 308 103 309
rect 101 308 102 309
rect 100 308 101 309
rect 99 308 100 309
rect 98 308 99 309
rect 97 308 98 309
rect 96 308 97 309
rect 95 308 96 309
rect 94 308 95 309
rect 93 308 94 309
rect 92 308 93 309
rect 91 308 92 309
rect 90 308 91 309
rect 89 308 90 309
rect 73 308 74 309
rect 72 308 73 309
rect 71 308 72 309
rect 70 308 71 309
rect 69 308 70 309
rect 68 308 69 309
rect 67 308 68 309
rect 66 308 67 309
rect 65 308 66 309
rect 64 308 65 309
rect 63 308 64 309
rect 62 308 63 309
rect 61 308 62 309
rect 60 308 61 309
rect 59 308 60 309
rect 58 308 59 309
rect 57 308 58 309
rect 56 308 57 309
rect 55 308 56 309
rect 54 308 55 309
rect 53 308 54 309
rect 52 308 53 309
rect 51 308 52 309
rect 50 308 51 309
rect 49 308 50 309
rect 48 308 49 309
rect 47 308 48 309
rect 46 308 47 309
rect 45 308 46 309
rect 44 308 45 309
rect 33 308 34 309
rect 32 308 33 309
rect 31 308 32 309
rect 30 308 31 309
rect 29 308 30 309
rect 28 308 29 309
rect 27 308 28 309
rect 26 308 27 309
rect 25 308 26 309
rect 24 308 25 309
rect 23 308 24 309
rect 22 308 23 309
rect 21 308 22 309
rect 20 308 21 309
rect 19 308 20 309
rect 18 308 19 309
rect 17 308 18 309
rect 16 308 17 309
rect 15 308 16 309
rect 14 308 15 309
rect 13 308 14 309
rect 12 308 13 309
rect 11 308 12 309
rect 10 308 11 309
rect 441 309 442 310
rect 440 309 441 310
rect 439 309 440 310
rect 438 309 439 310
rect 419 309 420 310
rect 418 309 419 310
rect 417 309 418 310
rect 416 309 417 310
rect 401 309 402 310
rect 400 309 401 310
rect 399 309 400 310
rect 398 309 399 310
rect 397 309 398 310
rect 261 309 262 310
rect 260 309 261 310
rect 259 309 260 310
rect 258 309 259 310
rect 257 309 258 310
rect 256 309 257 310
rect 255 309 256 310
rect 254 309 255 310
rect 253 309 254 310
rect 252 309 253 310
rect 251 309 252 310
rect 250 309 251 310
rect 249 309 250 310
rect 248 309 249 310
rect 247 309 248 310
rect 246 309 247 310
rect 245 309 246 310
rect 244 309 245 310
rect 243 309 244 310
rect 242 309 243 310
rect 241 309 242 310
rect 240 309 241 310
rect 239 309 240 310
rect 238 309 239 310
rect 237 309 238 310
rect 236 309 237 310
rect 235 309 236 310
rect 234 309 235 310
rect 233 309 234 310
rect 232 309 233 310
rect 231 309 232 310
rect 230 309 231 310
rect 229 309 230 310
rect 228 309 229 310
rect 227 309 228 310
rect 226 309 227 310
rect 225 309 226 310
rect 224 309 225 310
rect 223 309 224 310
rect 222 309 223 310
rect 221 309 222 310
rect 220 309 221 310
rect 219 309 220 310
rect 218 309 219 310
rect 217 309 218 310
rect 216 309 217 310
rect 215 309 216 310
rect 214 309 215 310
rect 213 309 214 310
rect 212 309 213 310
rect 211 309 212 310
rect 210 309 211 310
rect 209 309 210 310
rect 208 309 209 310
rect 207 309 208 310
rect 206 309 207 310
rect 205 309 206 310
rect 166 309 167 310
rect 165 309 166 310
rect 164 309 165 310
rect 127 309 128 310
rect 126 309 127 310
rect 125 309 126 310
rect 124 309 125 310
rect 123 309 124 310
rect 122 309 123 310
rect 121 309 122 310
rect 120 309 121 310
rect 119 309 120 310
rect 118 309 119 310
rect 117 309 118 310
rect 116 309 117 310
rect 115 309 116 310
rect 114 309 115 310
rect 113 309 114 310
rect 112 309 113 310
rect 111 309 112 310
rect 110 309 111 310
rect 109 309 110 310
rect 108 309 109 310
rect 107 309 108 310
rect 106 309 107 310
rect 105 309 106 310
rect 104 309 105 310
rect 103 309 104 310
rect 102 309 103 310
rect 101 309 102 310
rect 100 309 101 310
rect 99 309 100 310
rect 98 309 99 310
rect 97 309 98 310
rect 96 309 97 310
rect 95 309 96 310
rect 94 309 95 310
rect 93 309 94 310
rect 92 309 93 310
rect 91 309 92 310
rect 90 309 91 310
rect 73 309 74 310
rect 72 309 73 310
rect 71 309 72 310
rect 70 309 71 310
rect 69 309 70 310
rect 68 309 69 310
rect 67 309 68 310
rect 66 309 67 310
rect 65 309 66 310
rect 64 309 65 310
rect 63 309 64 310
rect 62 309 63 310
rect 61 309 62 310
rect 60 309 61 310
rect 59 309 60 310
rect 58 309 59 310
rect 57 309 58 310
rect 56 309 57 310
rect 55 309 56 310
rect 54 309 55 310
rect 53 309 54 310
rect 52 309 53 310
rect 51 309 52 310
rect 50 309 51 310
rect 49 309 50 310
rect 48 309 49 310
rect 47 309 48 310
rect 46 309 47 310
rect 45 309 46 310
rect 34 309 35 310
rect 33 309 34 310
rect 32 309 33 310
rect 31 309 32 310
rect 30 309 31 310
rect 29 309 30 310
rect 28 309 29 310
rect 27 309 28 310
rect 26 309 27 310
rect 25 309 26 310
rect 24 309 25 310
rect 23 309 24 310
rect 22 309 23 310
rect 21 309 22 310
rect 20 309 21 310
rect 19 309 20 310
rect 18 309 19 310
rect 17 309 18 310
rect 16 309 17 310
rect 15 309 16 310
rect 14 309 15 310
rect 13 309 14 310
rect 12 309 13 310
rect 11 309 12 310
rect 10 309 11 310
rect 441 310 442 311
rect 440 310 441 311
rect 439 310 440 311
rect 438 310 439 311
rect 437 310 438 311
rect 436 310 437 311
rect 435 310 436 311
rect 434 310 435 311
rect 433 310 434 311
rect 432 310 433 311
rect 431 310 432 311
rect 430 310 431 311
rect 429 310 430 311
rect 428 310 429 311
rect 427 310 428 311
rect 426 310 427 311
rect 425 310 426 311
rect 424 310 425 311
rect 423 310 424 311
rect 422 310 423 311
rect 421 310 422 311
rect 420 310 421 311
rect 419 310 420 311
rect 418 310 419 311
rect 417 310 418 311
rect 416 310 417 311
rect 415 310 416 311
rect 414 310 415 311
rect 413 310 414 311
rect 412 310 413 311
rect 411 310 412 311
rect 410 310 411 311
rect 409 310 410 311
rect 408 310 409 311
rect 407 310 408 311
rect 406 310 407 311
rect 405 310 406 311
rect 404 310 405 311
rect 403 310 404 311
rect 402 310 403 311
rect 401 310 402 311
rect 400 310 401 311
rect 399 310 400 311
rect 398 310 399 311
rect 397 310 398 311
rect 260 310 261 311
rect 259 310 260 311
rect 258 310 259 311
rect 257 310 258 311
rect 256 310 257 311
rect 255 310 256 311
rect 254 310 255 311
rect 253 310 254 311
rect 252 310 253 311
rect 251 310 252 311
rect 250 310 251 311
rect 249 310 250 311
rect 248 310 249 311
rect 247 310 248 311
rect 246 310 247 311
rect 245 310 246 311
rect 244 310 245 311
rect 243 310 244 311
rect 242 310 243 311
rect 241 310 242 311
rect 240 310 241 311
rect 239 310 240 311
rect 238 310 239 311
rect 237 310 238 311
rect 236 310 237 311
rect 235 310 236 311
rect 234 310 235 311
rect 233 310 234 311
rect 232 310 233 311
rect 231 310 232 311
rect 230 310 231 311
rect 229 310 230 311
rect 228 310 229 311
rect 227 310 228 311
rect 226 310 227 311
rect 225 310 226 311
rect 224 310 225 311
rect 223 310 224 311
rect 222 310 223 311
rect 221 310 222 311
rect 220 310 221 311
rect 219 310 220 311
rect 218 310 219 311
rect 217 310 218 311
rect 216 310 217 311
rect 215 310 216 311
rect 214 310 215 311
rect 213 310 214 311
rect 212 310 213 311
rect 211 310 212 311
rect 210 310 211 311
rect 209 310 210 311
rect 208 310 209 311
rect 207 310 208 311
rect 206 310 207 311
rect 205 310 206 311
rect 204 310 205 311
rect 128 310 129 311
rect 127 310 128 311
rect 126 310 127 311
rect 125 310 126 311
rect 124 310 125 311
rect 123 310 124 311
rect 122 310 123 311
rect 121 310 122 311
rect 120 310 121 311
rect 119 310 120 311
rect 118 310 119 311
rect 117 310 118 311
rect 116 310 117 311
rect 115 310 116 311
rect 114 310 115 311
rect 113 310 114 311
rect 112 310 113 311
rect 111 310 112 311
rect 110 310 111 311
rect 109 310 110 311
rect 108 310 109 311
rect 107 310 108 311
rect 106 310 107 311
rect 105 310 106 311
rect 104 310 105 311
rect 103 310 104 311
rect 102 310 103 311
rect 101 310 102 311
rect 100 310 101 311
rect 99 310 100 311
rect 98 310 99 311
rect 97 310 98 311
rect 96 310 97 311
rect 95 310 96 311
rect 94 310 95 311
rect 93 310 94 311
rect 92 310 93 311
rect 91 310 92 311
rect 90 310 91 311
rect 74 310 75 311
rect 73 310 74 311
rect 72 310 73 311
rect 71 310 72 311
rect 70 310 71 311
rect 69 310 70 311
rect 68 310 69 311
rect 67 310 68 311
rect 66 310 67 311
rect 65 310 66 311
rect 64 310 65 311
rect 63 310 64 311
rect 62 310 63 311
rect 61 310 62 311
rect 60 310 61 311
rect 59 310 60 311
rect 58 310 59 311
rect 57 310 58 311
rect 56 310 57 311
rect 55 310 56 311
rect 54 310 55 311
rect 53 310 54 311
rect 52 310 53 311
rect 51 310 52 311
rect 50 310 51 311
rect 49 310 50 311
rect 48 310 49 311
rect 47 310 48 311
rect 46 310 47 311
rect 45 310 46 311
rect 34 310 35 311
rect 33 310 34 311
rect 32 310 33 311
rect 31 310 32 311
rect 30 310 31 311
rect 29 310 30 311
rect 28 310 29 311
rect 27 310 28 311
rect 26 310 27 311
rect 25 310 26 311
rect 24 310 25 311
rect 23 310 24 311
rect 22 310 23 311
rect 21 310 22 311
rect 20 310 21 311
rect 19 310 20 311
rect 18 310 19 311
rect 17 310 18 311
rect 16 310 17 311
rect 15 310 16 311
rect 14 310 15 311
rect 13 310 14 311
rect 12 310 13 311
rect 11 310 12 311
rect 441 311 442 312
rect 440 311 441 312
rect 439 311 440 312
rect 438 311 439 312
rect 437 311 438 312
rect 436 311 437 312
rect 435 311 436 312
rect 434 311 435 312
rect 433 311 434 312
rect 432 311 433 312
rect 431 311 432 312
rect 430 311 431 312
rect 429 311 430 312
rect 428 311 429 312
rect 427 311 428 312
rect 426 311 427 312
rect 425 311 426 312
rect 424 311 425 312
rect 423 311 424 312
rect 422 311 423 312
rect 421 311 422 312
rect 420 311 421 312
rect 419 311 420 312
rect 418 311 419 312
rect 417 311 418 312
rect 416 311 417 312
rect 415 311 416 312
rect 414 311 415 312
rect 413 311 414 312
rect 412 311 413 312
rect 411 311 412 312
rect 410 311 411 312
rect 409 311 410 312
rect 408 311 409 312
rect 407 311 408 312
rect 406 311 407 312
rect 405 311 406 312
rect 404 311 405 312
rect 403 311 404 312
rect 402 311 403 312
rect 401 311 402 312
rect 400 311 401 312
rect 399 311 400 312
rect 398 311 399 312
rect 397 311 398 312
rect 258 311 259 312
rect 257 311 258 312
rect 256 311 257 312
rect 255 311 256 312
rect 254 311 255 312
rect 253 311 254 312
rect 252 311 253 312
rect 251 311 252 312
rect 250 311 251 312
rect 249 311 250 312
rect 248 311 249 312
rect 247 311 248 312
rect 246 311 247 312
rect 245 311 246 312
rect 244 311 245 312
rect 243 311 244 312
rect 242 311 243 312
rect 241 311 242 312
rect 240 311 241 312
rect 239 311 240 312
rect 238 311 239 312
rect 237 311 238 312
rect 236 311 237 312
rect 235 311 236 312
rect 234 311 235 312
rect 233 311 234 312
rect 232 311 233 312
rect 231 311 232 312
rect 230 311 231 312
rect 229 311 230 312
rect 228 311 229 312
rect 227 311 228 312
rect 226 311 227 312
rect 225 311 226 312
rect 224 311 225 312
rect 223 311 224 312
rect 222 311 223 312
rect 221 311 222 312
rect 220 311 221 312
rect 219 311 220 312
rect 218 311 219 312
rect 217 311 218 312
rect 216 311 217 312
rect 215 311 216 312
rect 214 311 215 312
rect 213 311 214 312
rect 212 311 213 312
rect 211 311 212 312
rect 210 311 211 312
rect 209 311 210 312
rect 208 311 209 312
rect 207 311 208 312
rect 206 311 207 312
rect 205 311 206 312
rect 204 311 205 312
rect 203 311 204 312
rect 129 311 130 312
rect 128 311 129 312
rect 127 311 128 312
rect 126 311 127 312
rect 125 311 126 312
rect 124 311 125 312
rect 123 311 124 312
rect 122 311 123 312
rect 121 311 122 312
rect 120 311 121 312
rect 119 311 120 312
rect 118 311 119 312
rect 117 311 118 312
rect 116 311 117 312
rect 115 311 116 312
rect 114 311 115 312
rect 113 311 114 312
rect 112 311 113 312
rect 111 311 112 312
rect 110 311 111 312
rect 109 311 110 312
rect 108 311 109 312
rect 107 311 108 312
rect 106 311 107 312
rect 105 311 106 312
rect 104 311 105 312
rect 103 311 104 312
rect 102 311 103 312
rect 101 311 102 312
rect 100 311 101 312
rect 99 311 100 312
rect 98 311 99 312
rect 97 311 98 312
rect 96 311 97 312
rect 95 311 96 312
rect 94 311 95 312
rect 93 311 94 312
rect 92 311 93 312
rect 91 311 92 312
rect 74 311 75 312
rect 73 311 74 312
rect 72 311 73 312
rect 71 311 72 312
rect 70 311 71 312
rect 69 311 70 312
rect 68 311 69 312
rect 67 311 68 312
rect 66 311 67 312
rect 65 311 66 312
rect 64 311 65 312
rect 63 311 64 312
rect 62 311 63 312
rect 61 311 62 312
rect 60 311 61 312
rect 59 311 60 312
rect 58 311 59 312
rect 57 311 58 312
rect 56 311 57 312
rect 55 311 56 312
rect 54 311 55 312
rect 53 311 54 312
rect 52 311 53 312
rect 51 311 52 312
rect 50 311 51 312
rect 49 311 50 312
rect 48 311 49 312
rect 47 311 48 312
rect 46 311 47 312
rect 45 311 46 312
rect 34 311 35 312
rect 33 311 34 312
rect 32 311 33 312
rect 31 311 32 312
rect 30 311 31 312
rect 29 311 30 312
rect 28 311 29 312
rect 27 311 28 312
rect 26 311 27 312
rect 25 311 26 312
rect 24 311 25 312
rect 23 311 24 312
rect 22 311 23 312
rect 21 311 22 312
rect 20 311 21 312
rect 19 311 20 312
rect 18 311 19 312
rect 17 311 18 312
rect 16 311 17 312
rect 15 311 16 312
rect 14 311 15 312
rect 13 311 14 312
rect 12 311 13 312
rect 441 312 442 313
rect 440 312 441 313
rect 439 312 440 313
rect 438 312 439 313
rect 437 312 438 313
rect 436 312 437 313
rect 435 312 436 313
rect 434 312 435 313
rect 433 312 434 313
rect 432 312 433 313
rect 431 312 432 313
rect 430 312 431 313
rect 429 312 430 313
rect 428 312 429 313
rect 427 312 428 313
rect 426 312 427 313
rect 425 312 426 313
rect 424 312 425 313
rect 423 312 424 313
rect 422 312 423 313
rect 421 312 422 313
rect 420 312 421 313
rect 419 312 420 313
rect 418 312 419 313
rect 417 312 418 313
rect 416 312 417 313
rect 415 312 416 313
rect 414 312 415 313
rect 413 312 414 313
rect 412 312 413 313
rect 411 312 412 313
rect 410 312 411 313
rect 409 312 410 313
rect 408 312 409 313
rect 407 312 408 313
rect 406 312 407 313
rect 405 312 406 313
rect 404 312 405 313
rect 403 312 404 313
rect 402 312 403 313
rect 401 312 402 313
rect 400 312 401 313
rect 399 312 400 313
rect 398 312 399 313
rect 397 312 398 313
rect 256 312 257 313
rect 255 312 256 313
rect 254 312 255 313
rect 253 312 254 313
rect 252 312 253 313
rect 251 312 252 313
rect 250 312 251 313
rect 249 312 250 313
rect 248 312 249 313
rect 247 312 248 313
rect 246 312 247 313
rect 245 312 246 313
rect 244 312 245 313
rect 243 312 244 313
rect 242 312 243 313
rect 241 312 242 313
rect 240 312 241 313
rect 239 312 240 313
rect 238 312 239 313
rect 237 312 238 313
rect 236 312 237 313
rect 235 312 236 313
rect 234 312 235 313
rect 233 312 234 313
rect 232 312 233 313
rect 231 312 232 313
rect 230 312 231 313
rect 229 312 230 313
rect 228 312 229 313
rect 227 312 228 313
rect 226 312 227 313
rect 225 312 226 313
rect 224 312 225 313
rect 223 312 224 313
rect 222 312 223 313
rect 221 312 222 313
rect 220 312 221 313
rect 219 312 220 313
rect 218 312 219 313
rect 217 312 218 313
rect 216 312 217 313
rect 215 312 216 313
rect 214 312 215 313
rect 213 312 214 313
rect 212 312 213 313
rect 211 312 212 313
rect 210 312 211 313
rect 209 312 210 313
rect 208 312 209 313
rect 207 312 208 313
rect 206 312 207 313
rect 205 312 206 313
rect 204 312 205 313
rect 203 312 204 313
rect 202 312 203 313
rect 130 312 131 313
rect 129 312 130 313
rect 128 312 129 313
rect 127 312 128 313
rect 126 312 127 313
rect 125 312 126 313
rect 124 312 125 313
rect 123 312 124 313
rect 122 312 123 313
rect 121 312 122 313
rect 120 312 121 313
rect 119 312 120 313
rect 118 312 119 313
rect 117 312 118 313
rect 116 312 117 313
rect 115 312 116 313
rect 114 312 115 313
rect 113 312 114 313
rect 112 312 113 313
rect 111 312 112 313
rect 110 312 111 313
rect 109 312 110 313
rect 108 312 109 313
rect 107 312 108 313
rect 106 312 107 313
rect 105 312 106 313
rect 104 312 105 313
rect 103 312 104 313
rect 102 312 103 313
rect 101 312 102 313
rect 100 312 101 313
rect 99 312 100 313
rect 98 312 99 313
rect 97 312 98 313
rect 96 312 97 313
rect 95 312 96 313
rect 94 312 95 313
rect 93 312 94 313
rect 92 312 93 313
rect 91 312 92 313
rect 74 312 75 313
rect 73 312 74 313
rect 72 312 73 313
rect 71 312 72 313
rect 70 312 71 313
rect 69 312 70 313
rect 68 312 69 313
rect 67 312 68 313
rect 66 312 67 313
rect 65 312 66 313
rect 64 312 65 313
rect 63 312 64 313
rect 62 312 63 313
rect 61 312 62 313
rect 60 312 61 313
rect 59 312 60 313
rect 58 312 59 313
rect 57 312 58 313
rect 56 312 57 313
rect 55 312 56 313
rect 54 312 55 313
rect 53 312 54 313
rect 52 312 53 313
rect 51 312 52 313
rect 50 312 51 313
rect 49 312 50 313
rect 48 312 49 313
rect 47 312 48 313
rect 46 312 47 313
rect 34 312 35 313
rect 33 312 34 313
rect 32 312 33 313
rect 31 312 32 313
rect 30 312 31 313
rect 29 312 30 313
rect 28 312 29 313
rect 27 312 28 313
rect 26 312 27 313
rect 25 312 26 313
rect 24 312 25 313
rect 23 312 24 313
rect 22 312 23 313
rect 21 312 22 313
rect 20 312 21 313
rect 19 312 20 313
rect 18 312 19 313
rect 17 312 18 313
rect 16 312 17 313
rect 15 312 16 313
rect 14 312 15 313
rect 13 312 14 313
rect 12 312 13 313
rect 441 313 442 314
rect 440 313 441 314
rect 439 313 440 314
rect 438 313 439 314
rect 437 313 438 314
rect 436 313 437 314
rect 435 313 436 314
rect 434 313 435 314
rect 433 313 434 314
rect 432 313 433 314
rect 431 313 432 314
rect 430 313 431 314
rect 429 313 430 314
rect 428 313 429 314
rect 427 313 428 314
rect 426 313 427 314
rect 425 313 426 314
rect 424 313 425 314
rect 423 313 424 314
rect 422 313 423 314
rect 421 313 422 314
rect 420 313 421 314
rect 419 313 420 314
rect 418 313 419 314
rect 417 313 418 314
rect 416 313 417 314
rect 415 313 416 314
rect 414 313 415 314
rect 413 313 414 314
rect 412 313 413 314
rect 411 313 412 314
rect 410 313 411 314
rect 409 313 410 314
rect 408 313 409 314
rect 407 313 408 314
rect 406 313 407 314
rect 405 313 406 314
rect 404 313 405 314
rect 403 313 404 314
rect 402 313 403 314
rect 401 313 402 314
rect 400 313 401 314
rect 399 313 400 314
rect 398 313 399 314
rect 397 313 398 314
rect 255 313 256 314
rect 254 313 255 314
rect 253 313 254 314
rect 252 313 253 314
rect 251 313 252 314
rect 250 313 251 314
rect 249 313 250 314
rect 248 313 249 314
rect 247 313 248 314
rect 246 313 247 314
rect 245 313 246 314
rect 244 313 245 314
rect 243 313 244 314
rect 242 313 243 314
rect 241 313 242 314
rect 240 313 241 314
rect 239 313 240 314
rect 238 313 239 314
rect 237 313 238 314
rect 236 313 237 314
rect 235 313 236 314
rect 234 313 235 314
rect 233 313 234 314
rect 232 313 233 314
rect 231 313 232 314
rect 230 313 231 314
rect 229 313 230 314
rect 228 313 229 314
rect 227 313 228 314
rect 226 313 227 314
rect 225 313 226 314
rect 224 313 225 314
rect 223 313 224 314
rect 222 313 223 314
rect 221 313 222 314
rect 220 313 221 314
rect 219 313 220 314
rect 218 313 219 314
rect 217 313 218 314
rect 216 313 217 314
rect 215 313 216 314
rect 214 313 215 314
rect 213 313 214 314
rect 212 313 213 314
rect 211 313 212 314
rect 210 313 211 314
rect 209 313 210 314
rect 208 313 209 314
rect 207 313 208 314
rect 206 313 207 314
rect 205 313 206 314
rect 204 313 205 314
rect 203 313 204 314
rect 202 313 203 314
rect 201 313 202 314
rect 131 313 132 314
rect 130 313 131 314
rect 129 313 130 314
rect 128 313 129 314
rect 127 313 128 314
rect 126 313 127 314
rect 125 313 126 314
rect 124 313 125 314
rect 123 313 124 314
rect 122 313 123 314
rect 121 313 122 314
rect 120 313 121 314
rect 119 313 120 314
rect 118 313 119 314
rect 117 313 118 314
rect 116 313 117 314
rect 115 313 116 314
rect 114 313 115 314
rect 113 313 114 314
rect 112 313 113 314
rect 111 313 112 314
rect 110 313 111 314
rect 109 313 110 314
rect 108 313 109 314
rect 107 313 108 314
rect 106 313 107 314
rect 105 313 106 314
rect 104 313 105 314
rect 103 313 104 314
rect 102 313 103 314
rect 101 313 102 314
rect 100 313 101 314
rect 99 313 100 314
rect 98 313 99 314
rect 97 313 98 314
rect 96 313 97 314
rect 95 313 96 314
rect 94 313 95 314
rect 93 313 94 314
rect 92 313 93 314
rect 75 313 76 314
rect 74 313 75 314
rect 73 313 74 314
rect 72 313 73 314
rect 71 313 72 314
rect 70 313 71 314
rect 69 313 70 314
rect 68 313 69 314
rect 67 313 68 314
rect 66 313 67 314
rect 65 313 66 314
rect 64 313 65 314
rect 63 313 64 314
rect 62 313 63 314
rect 61 313 62 314
rect 60 313 61 314
rect 59 313 60 314
rect 58 313 59 314
rect 57 313 58 314
rect 56 313 57 314
rect 55 313 56 314
rect 54 313 55 314
rect 53 313 54 314
rect 52 313 53 314
rect 51 313 52 314
rect 50 313 51 314
rect 49 313 50 314
rect 48 313 49 314
rect 47 313 48 314
rect 46 313 47 314
rect 35 313 36 314
rect 34 313 35 314
rect 33 313 34 314
rect 32 313 33 314
rect 31 313 32 314
rect 30 313 31 314
rect 29 313 30 314
rect 28 313 29 314
rect 27 313 28 314
rect 26 313 27 314
rect 25 313 26 314
rect 24 313 25 314
rect 23 313 24 314
rect 22 313 23 314
rect 21 313 22 314
rect 20 313 21 314
rect 19 313 20 314
rect 18 313 19 314
rect 17 313 18 314
rect 16 313 17 314
rect 15 313 16 314
rect 14 313 15 314
rect 13 313 14 314
rect 462 314 463 315
rect 441 314 442 315
rect 440 314 441 315
rect 439 314 440 315
rect 438 314 439 315
rect 437 314 438 315
rect 436 314 437 315
rect 435 314 436 315
rect 434 314 435 315
rect 433 314 434 315
rect 432 314 433 315
rect 431 314 432 315
rect 430 314 431 315
rect 429 314 430 315
rect 428 314 429 315
rect 427 314 428 315
rect 426 314 427 315
rect 425 314 426 315
rect 424 314 425 315
rect 423 314 424 315
rect 422 314 423 315
rect 421 314 422 315
rect 420 314 421 315
rect 419 314 420 315
rect 418 314 419 315
rect 417 314 418 315
rect 416 314 417 315
rect 415 314 416 315
rect 414 314 415 315
rect 413 314 414 315
rect 412 314 413 315
rect 411 314 412 315
rect 410 314 411 315
rect 409 314 410 315
rect 408 314 409 315
rect 407 314 408 315
rect 406 314 407 315
rect 405 314 406 315
rect 404 314 405 315
rect 403 314 404 315
rect 402 314 403 315
rect 401 314 402 315
rect 400 314 401 315
rect 399 314 400 315
rect 398 314 399 315
rect 397 314 398 315
rect 253 314 254 315
rect 252 314 253 315
rect 251 314 252 315
rect 250 314 251 315
rect 249 314 250 315
rect 248 314 249 315
rect 247 314 248 315
rect 246 314 247 315
rect 245 314 246 315
rect 244 314 245 315
rect 243 314 244 315
rect 242 314 243 315
rect 241 314 242 315
rect 240 314 241 315
rect 239 314 240 315
rect 238 314 239 315
rect 237 314 238 315
rect 236 314 237 315
rect 235 314 236 315
rect 234 314 235 315
rect 233 314 234 315
rect 232 314 233 315
rect 231 314 232 315
rect 230 314 231 315
rect 229 314 230 315
rect 228 314 229 315
rect 227 314 228 315
rect 226 314 227 315
rect 225 314 226 315
rect 224 314 225 315
rect 223 314 224 315
rect 222 314 223 315
rect 221 314 222 315
rect 220 314 221 315
rect 219 314 220 315
rect 218 314 219 315
rect 217 314 218 315
rect 216 314 217 315
rect 215 314 216 315
rect 214 314 215 315
rect 213 314 214 315
rect 212 314 213 315
rect 211 314 212 315
rect 210 314 211 315
rect 209 314 210 315
rect 208 314 209 315
rect 207 314 208 315
rect 206 314 207 315
rect 205 314 206 315
rect 204 314 205 315
rect 203 314 204 315
rect 202 314 203 315
rect 201 314 202 315
rect 200 314 201 315
rect 132 314 133 315
rect 131 314 132 315
rect 130 314 131 315
rect 129 314 130 315
rect 128 314 129 315
rect 127 314 128 315
rect 126 314 127 315
rect 125 314 126 315
rect 124 314 125 315
rect 123 314 124 315
rect 122 314 123 315
rect 121 314 122 315
rect 120 314 121 315
rect 119 314 120 315
rect 118 314 119 315
rect 117 314 118 315
rect 116 314 117 315
rect 115 314 116 315
rect 114 314 115 315
rect 113 314 114 315
rect 112 314 113 315
rect 111 314 112 315
rect 110 314 111 315
rect 109 314 110 315
rect 108 314 109 315
rect 107 314 108 315
rect 106 314 107 315
rect 105 314 106 315
rect 104 314 105 315
rect 103 314 104 315
rect 102 314 103 315
rect 101 314 102 315
rect 100 314 101 315
rect 99 314 100 315
rect 98 314 99 315
rect 97 314 98 315
rect 96 314 97 315
rect 95 314 96 315
rect 94 314 95 315
rect 93 314 94 315
rect 75 314 76 315
rect 74 314 75 315
rect 73 314 74 315
rect 72 314 73 315
rect 71 314 72 315
rect 70 314 71 315
rect 69 314 70 315
rect 68 314 69 315
rect 67 314 68 315
rect 66 314 67 315
rect 65 314 66 315
rect 64 314 65 315
rect 63 314 64 315
rect 62 314 63 315
rect 61 314 62 315
rect 60 314 61 315
rect 59 314 60 315
rect 58 314 59 315
rect 57 314 58 315
rect 56 314 57 315
rect 55 314 56 315
rect 54 314 55 315
rect 53 314 54 315
rect 52 314 53 315
rect 51 314 52 315
rect 50 314 51 315
rect 49 314 50 315
rect 48 314 49 315
rect 47 314 48 315
rect 46 314 47 315
rect 35 314 36 315
rect 34 314 35 315
rect 33 314 34 315
rect 32 314 33 315
rect 31 314 32 315
rect 30 314 31 315
rect 29 314 30 315
rect 28 314 29 315
rect 27 314 28 315
rect 26 314 27 315
rect 25 314 26 315
rect 24 314 25 315
rect 23 314 24 315
rect 22 314 23 315
rect 21 314 22 315
rect 20 314 21 315
rect 19 314 20 315
rect 18 314 19 315
rect 17 314 18 315
rect 16 314 17 315
rect 15 314 16 315
rect 14 314 15 315
rect 462 315 463 316
rect 441 315 442 316
rect 440 315 441 316
rect 439 315 440 316
rect 438 315 439 316
rect 437 315 438 316
rect 436 315 437 316
rect 435 315 436 316
rect 434 315 435 316
rect 433 315 434 316
rect 432 315 433 316
rect 431 315 432 316
rect 430 315 431 316
rect 429 315 430 316
rect 428 315 429 316
rect 427 315 428 316
rect 426 315 427 316
rect 425 315 426 316
rect 424 315 425 316
rect 423 315 424 316
rect 422 315 423 316
rect 421 315 422 316
rect 420 315 421 316
rect 419 315 420 316
rect 418 315 419 316
rect 417 315 418 316
rect 416 315 417 316
rect 415 315 416 316
rect 414 315 415 316
rect 413 315 414 316
rect 412 315 413 316
rect 411 315 412 316
rect 410 315 411 316
rect 409 315 410 316
rect 408 315 409 316
rect 407 315 408 316
rect 406 315 407 316
rect 405 315 406 316
rect 404 315 405 316
rect 403 315 404 316
rect 402 315 403 316
rect 401 315 402 316
rect 400 315 401 316
rect 399 315 400 316
rect 398 315 399 316
rect 397 315 398 316
rect 251 315 252 316
rect 250 315 251 316
rect 249 315 250 316
rect 248 315 249 316
rect 247 315 248 316
rect 246 315 247 316
rect 245 315 246 316
rect 244 315 245 316
rect 243 315 244 316
rect 242 315 243 316
rect 241 315 242 316
rect 240 315 241 316
rect 239 315 240 316
rect 238 315 239 316
rect 237 315 238 316
rect 236 315 237 316
rect 235 315 236 316
rect 234 315 235 316
rect 233 315 234 316
rect 232 315 233 316
rect 231 315 232 316
rect 230 315 231 316
rect 229 315 230 316
rect 228 315 229 316
rect 227 315 228 316
rect 226 315 227 316
rect 225 315 226 316
rect 224 315 225 316
rect 223 315 224 316
rect 222 315 223 316
rect 221 315 222 316
rect 220 315 221 316
rect 219 315 220 316
rect 218 315 219 316
rect 217 315 218 316
rect 216 315 217 316
rect 215 315 216 316
rect 214 315 215 316
rect 213 315 214 316
rect 212 315 213 316
rect 211 315 212 316
rect 210 315 211 316
rect 209 315 210 316
rect 208 315 209 316
rect 207 315 208 316
rect 206 315 207 316
rect 205 315 206 316
rect 204 315 205 316
rect 203 315 204 316
rect 202 315 203 316
rect 201 315 202 316
rect 200 315 201 316
rect 199 315 200 316
rect 133 315 134 316
rect 132 315 133 316
rect 131 315 132 316
rect 130 315 131 316
rect 129 315 130 316
rect 128 315 129 316
rect 127 315 128 316
rect 126 315 127 316
rect 125 315 126 316
rect 124 315 125 316
rect 123 315 124 316
rect 122 315 123 316
rect 121 315 122 316
rect 120 315 121 316
rect 119 315 120 316
rect 118 315 119 316
rect 117 315 118 316
rect 116 315 117 316
rect 115 315 116 316
rect 114 315 115 316
rect 113 315 114 316
rect 112 315 113 316
rect 111 315 112 316
rect 110 315 111 316
rect 109 315 110 316
rect 108 315 109 316
rect 107 315 108 316
rect 106 315 107 316
rect 105 315 106 316
rect 104 315 105 316
rect 103 315 104 316
rect 102 315 103 316
rect 101 315 102 316
rect 100 315 101 316
rect 99 315 100 316
rect 98 315 99 316
rect 97 315 98 316
rect 96 315 97 316
rect 95 315 96 316
rect 94 315 95 316
rect 93 315 94 316
rect 76 315 77 316
rect 75 315 76 316
rect 74 315 75 316
rect 73 315 74 316
rect 72 315 73 316
rect 71 315 72 316
rect 70 315 71 316
rect 69 315 70 316
rect 68 315 69 316
rect 67 315 68 316
rect 66 315 67 316
rect 65 315 66 316
rect 64 315 65 316
rect 63 315 64 316
rect 62 315 63 316
rect 61 315 62 316
rect 60 315 61 316
rect 59 315 60 316
rect 58 315 59 316
rect 57 315 58 316
rect 56 315 57 316
rect 55 315 56 316
rect 54 315 55 316
rect 53 315 54 316
rect 52 315 53 316
rect 51 315 52 316
rect 50 315 51 316
rect 49 315 50 316
rect 48 315 49 316
rect 47 315 48 316
rect 35 315 36 316
rect 34 315 35 316
rect 33 315 34 316
rect 32 315 33 316
rect 31 315 32 316
rect 30 315 31 316
rect 29 315 30 316
rect 28 315 29 316
rect 27 315 28 316
rect 26 315 27 316
rect 25 315 26 316
rect 24 315 25 316
rect 23 315 24 316
rect 22 315 23 316
rect 21 315 22 316
rect 20 315 21 316
rect 19 315 20 316
rect 18 315 19 316
rect 17 315 18 316
rect 16 315 17 316
rect 15 315 16 316
rect 14 315 15 316
rect 463 316 464 317
rect 462 316 463 317
rect 441 316 442 317
rect 440 316 441 317
rect 439 316 440 317
rect 438 316 439 317
rect 437 316 438 317
rect 436 316 437 317
rect 435 316 436 317
rect 434 316 435 317
rect 433 316 434 317
rect 432 316 433 317
rect 431 316 432 317
rect 430 316 431 317
rect 429 316 430 317
rect 428 316 429 317
rect 427 316 428 317
rect 426 316 427 317
rect 425 316 426 317
rect 424 316 425 317
rect 423 316 424 317
rect 422 316 423 317
rect 421 316 422 317
rect 420 316 421 317
rect 419 316 420 317
rect 418 316 419 317
rect 417 316 418 317
rect 416 316 417 317
rect 415 316 416 317
rect 414 316 415 317
rect 413 316 414 317
rect 412 316 413 317
rect 411 316 412 317
rect 410 316 411 317
rect 409 316 410 317
rect 408 316 409 317
rect 407 316 408 317
rect 406 316 407 317
rect 405 316 406 317
rect 404 316 405 317
rect 403 316 404 317
rect 402 316 403 317
rect 401 316 402 317
rect 400 316 401 317
rect 399 316 400 317
rect 398 316 399 317
rect 397 316 398 317
rect 249 316 250 317
rect 248 316 249 317
rect 247 316 248 317
rect 246 316 247 317
rect 245 316 246 317
rect 244 316 245 317
rect 243 316 244 317
rect 242 316 243 317
rect 241 316 242 317
rect 240 316 241 317
rect 239 316 240 317
rect 238 316 239 317
rect 237 316 238 317
rect 236 316 237 317
rect 235 316 236 317
rect 234 316 235 317
rect 233 316 234 317
rect 232 316 233 317
rect 231 316 232 317
rect 230 316 231 317
rect 229 316 230 317
rect 228 316 229 317
rect 227 316 228 317
rect 226 316 227 317
rect 225 316 226 317
rect 224 316 225 317
rect 223 316 224 317
rect 222 316 223 317
rect 221 316 222 317
rect 220 316 221 317
rect 219 316 220 317
rect 218 316 219 317
rect 217 316 218 317
rect 216 316 217 317
rect 215 316 216 317
rect 214 316 215 317
rect 213 316 214 317
rect 212 316 213 317
rect 211 316 212 317
rect 210 316 211 317
rect 209 316 210 317
rect 208 316 209 317
rect 207 316 208 317
rect 206 316 207 317
rect 205 316 206 317
rect 204 316 205 317
rect 203 316 204 317
rect 202 316 203 317
rect 201 316 202 317
rect 200 316 201 317
rect 199 316 200 317
rect 198 316 199 317
rect 134 316 135 317
rect 133 316 134 317
rect 132 316 133 317
rect 131 316 132 317
rect 130 316 131 317
rect 129 316 130 317
rect 128 316 129 317
rect 127 316 128 317
rect 126 316 127 317
rect 125 316 126 317
rect 124 316 125 317
rect 123 316 124 317
rect 122 316 123 317
rect 121 316 122 317
rect 120 316 121 317
rect 119 316 120 317
rect 118 316 119 317
rect 117 316 118 317
rect 116 316 117 317
rect 115 316 116 317
rect 114 316 115 317
rect 113 316 114 317
rect 112 316 113 317
rect 111 316 112 317
rect 110 316 111 317
rect 109 316 110 317
rect 108 316 109 317
rect 107 316 108 317
rect 106 316 107 317
rect 105 316 106 317
rect 104 316 105 317
rect 103 316 104 317
rect 102 316 103 317
rect 101 316 102 317
rect 100 316 101 317
rect 99 316 100 317
rect 98 316 99 317
rect 97 316 98 317
rect 96 316 97 317
rect 95 316 96 317
rect 94 316 95 317
rect 76 316 77 317
rect 75 316 76 317
rect 74 316 75 317
rect 73 316 74 317
rect 72 316 73 317
rect 71 316 72 317
rect 70 316 71 317
rect 69 316 70 317
rect 68 316 69 317
rect 67 316 68 317
rect 66 316 67 317
rect 65 316 66 317
rect 64 316 65 317
rect 63 316 64 317
rect 62 316 63 317
rect 61 316 62 317
rect 60 316 61 317
rect 59 316 60 317
rect 58 316 59 317
rect 57 316 58 317
rect 56 316 57 317
rect 55 316 56 317
rect 54 316 55 317
rect 53 316 54 317
rect 52 316 53 317
rect 51 316 52 317
rect 50 316 51 317
rect 49 316 50 317
rect 48 316 49 317
rect 47 316 48 317
rect 35 316 36 317
rect 34 316 35 317
rect 33 316 34 317
rect 32 316 33 317
rect 31 316 32 317
rect 30 316 31 317
rect 29 316 30 317
rect 28 316 29 317
rect 27 316 28 317
rect 26 316 27 317
rect 25 316 26 317
rect 24 316 25 317
rect 23 316 24 317
rect 22 316 23 317
rect 21 316 22 317
rect 20 316 21 317
rect 19 316 20 317
rect 18 316 19 317
rect 17 316 18 317
rect 16 316 17 317
rect 15 316 16 317
rect 465 317 466 318
rect 464 317 465 318
rect 463 317 464 318
rect 462 317 463 318
rect 441 317 442 318
rect 440 317 441 318
rect 439 317 440 318
rect 438 317 439 318
rect 437 317 438 318
rect 436 317 437 318
rect 435 317 436 318
rect 434 317 435 318
rect 433 317 434 318
rect 432 317 433 318
rect 431 317 432 318
rect 430 317 431 318
rect 429 317 430 318
rect 428 317 429 318
rect 427 317 428 318
rect 426 317 427 318
rect 425 317 426 318
rect 424 317 425 318
rect 423 317 424 318
rect 422 317 423 318
rect 421 317 422 318
rect 420 317 421 318
rect 419 317 420 318
rect 418 317 419 318
rect 417 317 418 318
rect 416 317 417 318
rect 415 317 416 318
rect 414 317 415 318
rect 413 317 414 318
rect 412 317 413 318
rect 411 317 412 318
rect 410 317 411 318
rect 409 317 410 318
rect 408 317 409 318
rect 407 317 408 318
rect 406 317 407 318
rect 405 317 406 318
rect 404 317 405 318
rect 403 317 404 318
rect 402 317 403 318
rect 401 317 402 318
rect 400 317 401 318
rect 399 317 400 318
rect 398 317 399 318
rect 397 317 398 318
rect 247 317 248 318
rect 246 317 247 318
rect 245 317 246 318
rect 244 317 245 318
rect 243 317 244 318
rect 242 317 243 318
rect 241 317 242 318
rect 240 317 241 318
rect 239 317 240 318
rect 238 317 239 318
rect 237 317 238 318
rect 236 317 237 318
rect 235 317 236 318
rect 234 317 235 318
rect 233 317 234 318
rect 232 317 233 318
rect 231 317 232 318
rect 230 317 231 318
rect 229 317 230 318
rect 228 317 229 318
rect 227 317 228 318
rect 226 317 227 318
rect 225 317 226 318
rect 224 317 225 318
rect 223 317 224 318
rect 222 317 223 318
rect 221 317 222 318
rect 220 317 221 318
rect 219 317 220 318
rect 218 317 219 318
rect 217 317 218 318
rect 216 317 217 318
rect 215 317 216 318
rect 214 317 215 318
rect 213 317 214 318
rect 212 317 213 318
rect 211 317 212 318
rect 210 317 211 318
rect 209 317 210 318
rect 208 317 209 318
rect 207 317 208 318
rect 206 317 207 318
rect 205 317 206 318
rect 204 317 205 318
rect 203 317 204 318
rect 202 317 203 318
rect 201 317 202 318
rect 200 317 201 318
rect 199 317 200 318
rect 198 317 199 318
rect 197 317 198 318
rect 135 317 136 318
rect 134 317 135 318
rect 133 317 134 318
rect 132 317 133 318
rect 131 317 132 318
rect 130 317 131 318
rect 129 317 130 318
rect 128 317 129 318
rect 127 317 128 318
rect 126 317 127 318
rect 125 317 126 318
rect 124 317 125 318
rect 123 317 124 318
rect 122 317 123 318
rect 121 317 122 318
rect 120 317 121 318
rect 119 317 120 318
rect 118 317 119 318
rect 117 317 118 318
rect 116 317 117 318
rect 115 317 116 318
rect 114 317 115 318
rect 113 317 114 318
rect 112 317 113 318
rect 111 317 112 318
rect 110 317 111 318
rect 109 317 110 318
rect 108 317 109 318
rect 107 317 108 318
rect 106 317 107 318
rect 105 317 106 318
rect 104 317 105 318
rect 103 317 104 318
rect 102 317 103 318
rect 101 317 102 318
rect 100 317 101 318
rect 99 317 100 318
rect 98 317 99 318
rect 97 317 98 318
rect 96 317 97 318
rect 95 317 96 318
rect 94 317 95 318
rect 77 317 78 318
rect 76 317 77 318
rect 75 317 76 318
rect 74 317 75 318
rect 73 317 74 318
rect 72 317 73 318
rect 71 317 72 318
rect 70 317 71 318
rect 69 317 70 318
rect 68 317 69 318
rect 67 317 68 318
rect 66 317 67 318
rect 65 317 66 318
rect 64 317 65 318
rect 63 317 64 318
rect 62 317 63 318
rect 61 317 62 318
rect 60 317 61 318
rect 59 317 60 318
rect 58 317 59 318
rect 57 317 58 318
rect 56 317 57 318
rect 55 317 56 318
rect 54 317 55 318
rect 53 317 54 318
rect 52 317 53 318
rect 51 317 52 318
rect 50 317 51 318
rect 49 317 50 318
rect 48 317 49 318
rect 47 317 48 318
rect 36 317 37 318
rect 35 317 36 318
rect 34 317 35 318
rect 33 317 34 318
rect 32 317 33 318
rect 31 317 32 318
rect 30 317 31 318
rect 29 317 30 318
rect 28 317 29 318
rect 27 317 28 318
rect 26 317 27 318
rect 25 317 26 318
rect 24 317 25 318
rect 23 317 24 318
rect 22 317 23 318
rect 21 317 22 318
rect 20 317 21 318
rect 19 317 20 318
rect 18 317 19 318
rect 17 317 18 318
rect 16 317 17 318
rect 15 317 16 318
rect 467 318 468 319
rect 466 318 467 319
rect 465 318 466 319
rect 464 318 465 319
rect 463 318 464 319
rect 462 318 463 319
rect 441 318 442 319
rect 440 318 441 319
rect 439 318 440 319
rect 438 318 439 319
rect 437 318 438 319
rect 436 318 437 319
rect 435 318 436 319
rect 434 318 435 319
rect 433 318 434 319
rect 432 318 433 319
rect 431 318 432 319
rect 430 318 431 319
rect 429 318 430 319
rect 428 318 429 319
rect 427 318 428 319
rect 426 318 427 319
rect 425 318 426 319
rect 424 318 425 319
rect 423 318 424 319
rect 422 318 423 319
rect 421 318 422 319
rect 420 318 421 319
rect 419 318 420 319
rect 418 318 419 319
rect 417 318 418 319
rect 416 318 417 319
rect 415 318 416 319
rect 414 318 415 319
rect 413 318 414 319
rect 412 318 413 319
rect 411 318 412 319
rect 410 318 411 319
rect 409 318 410 319
rect 408 318 409 319
rect 407 318 408 319
rect 406 318 407 319
rect 405 318 406 319
rect 404 318 405 319
rect 403 318 404 319
rect 402 318 403 319
rect 401 318 402 319
rect 400 318 401 319
rect 399 318 400 319
rect 398 318 399 319
rect 397 318 398 319
rect 244 318 245 319
rect 243 318 244 319
rect 242 318 243 319
rect 241 318 242 319
rect 240 318 241 319
rect 239 318 240 319
rect 238 318 239 319
rect 237 318 238 319
rect 236 318 237 319
rect 235 318 236 319
rect 234 318 235 319
rect 233 318 234 319
rect 232 318 233 319
rect 231 318 232 319
rect 230 318 231 319
rect 229 318 230 319
rect 228 318 229 319
rect 227 318 228 319
rect 226 318 227 319
rect 225 318 226 319
rect 224 318 225 319
rect 223 318 224 319
rect 222 318 223 319
rect 221 318 222 319
rect 220 318 221 319
rect 219 318 220 319
rect 218 318 219 319
rect 217 318 218 319
rect 216 318 217 319
rect 215 318 216 319
rect 214 318 215 319
rect 213 318 214 319
rect 212 318 213 319
rect 211 318 212 319
rect 210 318 211 319
rect 209 318 210 319
rect 208 318 209 319
rect 207 318 208 319
rect 206 318 207 319
rect 205 318 206 319
rect 204 318 205 319
rect 203 318 204 319
rect 202 318 203 319
rect 201 318 202 319
rect 200 318 201 319
rect 199 318 200 319
rect 198 318 199 319
rect 197 318 198 319
rect 196 318 197 319
rect 136 318 137 319
rect 135 318 136 319
rect 134 318 135 319
rect 133 318 134 319
rect 132 318 133 319
rect 131 318 132 319
rect 130 318 131 319
rect 129 318 130 319
rect 128 318 129 319
rect 127 318 128 319
rect 126 318 127 319
rect 125 318 126 319
rect 124 318 125 319
rect 123 318 124 319
rect 122 318 123 319
rect 121 318 122 319
rect 120 318 121 319
rect 119 318 120 319
rect 118 318 119 319
rect 117 318 118 319
rect 116 318 117 319
rect 115 318 116 319
rect 114 318 115 319
rect 113 318 114 319
rect 112 318 113 319
rect 111 318 112 319
rect 110 318 111 319
rect 109 318 110 319
rect 108 318 109 319
rect 107 318 108 319
rect 106 318 107 319
rect 105 318 106 319
rect 104 318 105 319
rect 103 318 104 319
rect 102 318 103 319
rect 101 318 102 319
rect 100 318 101 319
rect 99 318 100 319
rect 98 318 99 319
rect 97 318 98 319
rect 96 318 97 319
rect 95 318 96 319
rect 77 318 78 319
rect 76 318 77 319
rect 75 318 76 319
rect 74 318 75 319
rect 73 318 74 319
rect 72 318 73 319
rect 71 318 72 319
rect 70 318 71 319
rect 69 318 70 319
rect 68 318 69 319
rect 67 318 68 319
rect 66 318 67 319
rect 65 318 66 319
rect 64 318 65 319
rect 63 318 64 319
rect 62 318 63 319
rect 61 318 62 319
rect 60 318 61 319
rect 59 318 60 319
rect 58 318 59 319
rect 57 318 58 319
rect 56 318 57 319
rect 55 318 56 319
rect 54 318 55 319
rect 53 318 54 319
rect 52 318 53 319
rect 51 318 52 319
rect 50 318 51 319
rect 49 318 50 319
rect 48 318 49 319
rect 36 318 37 319
rect 35 318 36 319
rect 34 318 35 319
rect 33 318 34 319
rect 32 318 33 319
rect 31 318 32 319
rect 30 318 31 319
rect 29 318 30 319
rect 28 318 29 319
rect 27 318 28 319
rect 26 318 27 319
rect 25 318 26 319
rect 24 318 25 319
rect 23 318 24 319
rect 22 318 23 319
rect 21 318 22 319
rect 20 318 21 319
rect 19 318 20 319
rect 18 318 19 319
rect 17 318 18 319
rect 16 318 17 319
rect 482 319 483 320
rect 468 319 469 320
rect 467 319 468 320
rect 466 319 467 320
rect 465 319 466 320
rect 464 319 465 320
rect 463 319 464 320
rect 462 319 463 320
rect 441 319 442 320
rect 440 319 441 320
rect 439 319 440 320
rect 438 319 439 320
rect 437 319 438 320
rect 436 319 437 320
rect 435 319 436 320
rect 434 319 435 320
rect 433 319 434 320
rect 432 319 433 320
rect 431 319 432 320
rect 430 319 431 320
rect 429 319 430 320
rect 428 319 429 320
rect 427 319 428 320
rect 426 319 427 320
rect 425 319 426 320
rect 424 319 425 320
rect 423 319 424 320
rect 422 319 423 320
rect 421 319 422 320
rect 420 319 421 320
rect 419 319 420 320
rect 418 319 419 320
rect 417 319 418 320
rect 416 319 417 320
rect 415 319 416 320
rect 414 319 415 320
rect 413 319 414 320
rect 412 319 413 320
rect 411 319 412 320
rect 410 319 411 320
rect 409 319 410 320
rect 408 319 409 320
rect 407 319 408 320
rect 406 319 407 320
rect 405 319 406 320
rect 404 319 405 320
rect 403 319 404 320
rect 402 319 403 320
rect 401 319 402 320
rect 400 319 401 320
rect 399 319 400 320
rect 398 319 399 320
rect 397 319 398 320
rect 242 319 243 320
rect 241 319 242 320
rect 240 319 241 320
rect 239 319 240 320
rect 238 319 239 320
rect 237 319 238 320
rect 236 319 237 320
rect 235 319 236 320
rect 234 319 235 320
rect 233 319 234 320
rect 232 319 233 320
rect 231 319 232 320
rect 230 319 231 320
rect 229 319 230 320
rect 228 319 229 320
rect 227 319 228 320
rect 226 319 227 320
rect 225 319 226 320
rect 224 319 225 320
rect 223 319 224 320
rect 222 319 223 320
rect 221 319 222 320
rect 220 319 221 320
rect 219 319 220 320
rect 218 319 219 320
rect 217 319 218 320
rect 216 319 217 320
rect 215 319 216 320
rect 214 319 215 320
rect 213 319 214 320
rect 212 319 213 320
rect 211 319 212 320
rect 210 319 211 320
rect 209 319 210 320
rect 208 319 209 320
rect 207 319 208 320
rect 206 319 207 320
rect 205 319 206 320
rect 204 319 205 320
rect 203 319 204 320
rect 202 319 203 320
rect 201 319 202 320
rect 200 319 201 320
rect 199 319 200 320
rect 198 319 199 320
rect 197 319 198 320
rect 196 319 197 320
rect 195 319 196 320
rect 138 319 139 320
rect 137 319 138 320
rect 136 319 137 320
rect 135 319 136 320
rect 134 319 135 320
rect 133 319 134 320
rect 132 319 133 320
rect 131 319 132 320
rect 130 319 131 320
rect 129 319 130 320
rect 128 319 129 320
rect 127 319 128 320
rect 126 319 127 320
rect 125 319 126 320
rect 124 319 125 320
rect 123 319 124 320
rect 122 319 123 320
rect 121 319 122 320
rect 120 319 121 320
rect 119 319 120 320
rect 118 319 119 320
rect 117 319 118 320
rect 116 319 117 320
rect 115 319 116 320
rect 114 319 115 320
rect 113 319 114 320
rect 112 319 113 320
rect 111 319 112 320
rect 110 319 111 320
rect 109 319 110 320
rect 108 319 109 320
rect 107 319 108 320
rect 106 319 107 320
rect 105 319 106 320
rect 104 319 105 320
rect 103 319 104 320
rect 102 319 103 320
rect 101 319 102 320
rect 100 319 101 320
rect 99 319 100 320
rect 98 319 99 320
rect 97 319 98 320
rect 96 319 97 320
rect 78 319 79 320
rect 77 319 78 320
rect 76 319 77 320
rect 75 319 76 320
rect 74 319 75 320
rect 73 319 74 320
rect 72 319 73 320
rect 71 319 72 320
rect 70 319 71 320
rect 69 319 70 320
rect 68 319 69 320
rect 67 319 68 320
rect 66 319 67 320
rect 65 319 66 320
rect 64 319 65 320
rect 63 319 64 320
rect 62 319 63 320
rect 61 319 62 320
rect 60 319 61 320
rect 59 319 60 320
rect 58 319 59 320
rect 57 319 58 320
rect 56 319 57 320
rect 55 319 56 320
rect 54 319 55 320
rect 53 319 54 320
rect 52 319 53 320
rect 51 319 52 320
rect 50 319 51 320
rect 49 319 50 320
rect 48 319 49 320
rect 36 319 37 320
rect 35 319 36 320
rect 34 319 35 320
rect 33 319 34 320
rect 32 319 33 320
rect 31 319 32 320
rect 30 319 31 320
rect 29 319 30 320
rect 28 319 29 320
rect 27 319 28 320
rect 26 319 27 320
rect 25 319 26 320
rect 24 319 25 320
rect 23 319 24 320
rect 22 319 23 320
rect 21 319 22 320
rect 20 319 21 320
rect 19 319 20 320
rect 18 319 19 320
rect 17 319 18 320
rect 482 320 483 321
rect 470 320 471 321
rect 469 320 470 321
rect 468 320 469 321
rect 467 320 468 321
rect 466 320 467 321
rect 465 320 466 321
rect 464 320 465 321
rect 463 320 464 321
rect 462 320 463 321
rect 441 320 442 321
rect 440 320 441 321
rect 439 320 440 321
rect 438 320 439 321
rect 400 320 401 321
rect 399 320 400 321
rect 398 320 399 321
rect 397 320 398 321
rect 239 320 240 321
rect 238 320 239 321
rect 237 320 238 321
rect 236 320 237 321
rect 235 320 236 321
rect 234 320 235 321
rect 233 320 234 321
rect 232 320 233 321
rect 231 320 232 321
rect 230 320 231 321
rect 229 320 230 321
rect 228 320 229 321
rect 227 320 228 321
rect 226 320 227 321
rect 225 320 226 321
rect 224 320 225 321
rect 223 320 224 321
rect 222 320 223 321
rect 221 320 222 321
rect 220 320 221 321
rect 219 320 220 321
rect 218 320 219 321
rect 217 320 218 321
rect 216 320 217 321
rect 215 320 216 321
rect 214 320 215 321
rect 213 320 214 321
rect 212 320 213 321
rect 211 320 212 321
rect 210 320 211 321
rect 209 320 210 321
rect 208 320 209 321
rect 207 320 208 321
rect 206 320 207 321
rect 205 320 206 321
rect 204 320 205 321
rect 203 320 204 321
rect 202 320 203 321
rect 201 320 202 321
rect 200 320 201 321
rect 199 320 200 321
rect 198 320 199 321
rect 197 320 198 321
rect 196 320 197 321
rect 195 320 196 321
rect 194 320 195 321
rect 139 320 140 321
rect 138 320 139 321
rect 137 320 138 321
rect 136 320 137 321
rect 135 320 136 321
rect 134 320 135 321
rect 133 320 134 321
rect 132 320 133 321
rect 131 320 132 321
rect 130 320 131 321
rect 129 320 130 321
rect 128 320 129 321
rect 127 320 128 321
rect 126 320 127 321
rect 125 320 126 321
rect 124 320 125 321
rect 123 320 124 321
rect 122 320 123 321
rect 121 320 122 321
rect 120 320 121 321
rect 119 320 120 321
rect 118 320 119 321
rect 117 320 118 321
rect 116 320 117 321
rect 115 320 116 321
rect 114 320 115 321
rect 113 320 114 321
rect 112 320 113 321
rect 111 320 112 321
rect 110 320 111 321
rect 109 320 110 321
rect 108 320 109 321
rect 107 320 108 321
rect 106 320 107 321
rect 105 320 106 321
rect 104 320 105 321
rect 103 320 104 321
rect 102 320 103 321
rect 101 320 102 321
rect 100 320 101 321
rect 99 320 100 321
rect 98 320 99 321
rect 97 320 98 321
rect 96 320 97 321
rect 78 320 79 321
rect 77 320 78 321
rect 76 320 77 321
rect 75 320 76 321
rect 74 320 75 321
rect 73 320 74 321
rect 72 320 73 321
rect 71 320 72 321
rect 70 320 71 321
rect 69 320 70 321
rect 68 320 69 321
rect 67 320 68 321
rect 66 320 67 321
rect 65 320 66 321
rect 64 320 65 321
rect 63 320 64 321
rect 62 320 63 321
rect 61 320 62 321
rect 60 320 61 321
rect 59 320 60 321
rect 58 320 59 321
rect 57 320 58 321
rect 56 320 57 321
rect 55 320 56 321
rect 54 320 55 321
rect 53 320 54 321
rect 52 320 53 321
rect 51 320 52 321
rect 50 320 51 321
rect 49 320 50 321
rect 48 320 49 321
rect 37 320 38 321
rect 36 320 37 321
rect 35 320 36 321
rect 34 320 35 321
rect 33 320 34 321
rect 32 320 33 321
rect 31 320 32 321
rect 30 320 31 321
rect 29 320 30 321
rect 28 320 29 321
rect 27 320 28 321
rect 26 320 27 321
rect 25 320 26 321
rect 24 320 25 321
rect 23 320 24 321
rect 22 320 23 321
rect 21 320 22 321
rect 20 320 21 321
rect 19 320 20 321
rect 18 320 19 321
rect 482 321 483 322
rect 481 321 482 322
rect 472 321 473 322
rect 471 321 472 322
rect 470 321 471 322
rect 469 321 470 322
rect 468 321 469 322
rect 467 321 468 322
rect 466 321 467 322
rect 465 321 466 322
rect 464 321 465 322
rect 463 321 464 322
rect 462 321 463 322
rect 441 321 442 322
rect 440 321 441 322
rect 439 321 440 322
rect 399 321 400 322
rect 398 321 399 322
rect 397 321 398 322
rect 236 321 237 322
rect 235 321 236 322
rect 234 321 235 322
rect 233 321 234 322
rect 232 321 233 322
rect 231 321 232 322
rect 230 321 231 322
rect 229 321 230 322
rect 228 321 229 322
rect 227 321 228 322
rect 226 321 227 322
rect 225 321 226 322
rect 224 321 225 322
rect 223 321 224 322
rect 222 321 223 322
rect 221 321 222 322
rect 220 321 221 322
rect 219 321 220 322
rect 218 321 219 322
rect 217 321 218 322
rect 216 321 217 322
rect 215 321 216 322
rect 214 321 215 322
rect 213 321 214 322
rect 212 321 213 322
rect 211 321 212 322
rect 210 321 211 322
rect 209 321 210 322
rect 208 321 209 322
rect 207 321 208 322
rect 206 321 207 322
rect 205 321 206 322
rect 204 321 205 322
rect 203 321 204 322
rect 202 321 203 322
rect 201 321 202 322
rect 200 321 201 322
rect 199 321 200 322
rect 198 321 199 322
rect 197 321 198 322
rect 196 321 197 322
rect 195 321 196 322
rect 194 321 195 322
rect 193 321 194 322
rect 140 321 141 322
rect 139 321 140 322
rect 138 321 139 322
rect 137 321 138 322
rect 136 321 137 322
rect 135 321 136 322
rect 134 321 135 322
rect 133 321 134 322
rect 132 321 133 322
rect 131 321 132 322
rect 130 321 131 322
rect 129 321 130 322
rect 128 321 129 322
rect 127 321 128 322
rect 126 321 127 322
rect 125 321 126 322
rect 124 321 125 322
rect 123 321 124 322
rect 122 321 123 322
rect 121 321 122 322
rect 120 321 121 322
rect 119 321 120 322
rect 118 321 119 322
rect 117 321 118 322
rect 116 321 117 322
rect 115 321 116 322
rect 114 321 115 322
rect 113 321 114 322
rect 112 321 113 322
rect 111 321 112 322
rect 110 321 111 322
rect 109 321 110 322
rect 108 321 109 322
rect 107 321 108 322
rect 106 321 107 322
rect 105 321 106 322
rect 104 321 105 322
rect 103 321 104 322
rect 102 321 103 322
rect 101 321 102 322
rect 100 321 101 322
rect 99 321 100 322
rect 98 321 99 322
rect 97 321 98 322
rect 79 321 80 322
rect 78 321 79 322
rect 77 321 78 322
rect 76 321 77 322
rect 75 321 76 322
rect 74 321 75 322
rect 73 321 74 322
rect 72 321 73 322
rect 71 321 72 322
rect 70 321 71 322
rect 69 321 70 322
rect 68 321 69 322
rect 67 321 68 322
rect 66 321 67 322
rect 65 321 66 322
rect 64 321 65 322
rect 63 321 64 322
rect 62 321 63 322
rect 61 321 62 322
rect 60 321 61 322
rect 59 321 60 322
rect 58 321 59 322
rect 57 321 58 322
rect 56 321 57 322
rect 55 321 56 322
rect 54 321 55 322
rect 53 321 54 322
rect 52 321 53 322
rect 51 321 52 322
rect 50 321 51 322
rect 49 321 50 322
rect 37 321 38 322
rect 36 321 37 322
rect 35 321 36 322
rect 34 321 35 322
rect 33 321 34 322
rect 32 321 33 322
rect 31 321 32 322
rect 30 321 31 322
rect 29 321 30 322
rect 28 321 29 322
rect 27 321 28 322
rect 26 321 27 322
rect 25 321 26 322
rect 24 321 25 322
rect 23 321 24 322
rect 22 321 23 322
rect 21 321 22 322
rect 20 321 21 322
rect 19 321 20 322
rect 18 321 19 322
rect 482 322 483 323
rect 481 322 482 323
rect 480 322 481 323
rect 479 322 480 323
rect 478 322 479 323
rect 477 322 478 323
rect 476 322 477 323
rect 475 322 476 323
rect 474 322 475 323
rect 473 322 474 323
rect 472 322 473 323
rect 471 322 472 323
rect 470 322 471 323
rect 469 322 470 323
rect 468 322 469 323
rect 467 322 468 323
rect 466 322 467 323
rect 462 322 463 323
rect 441 322 442 323
rect 440 322 441 323
rect 439 322 440 323
rect 399 322 400 323
rect 398 322 399 323
rect 397 322 398 323
rect 232 322 233 323
rect 231 322 232 323
rect 230 322 231 323
rect 229 322 230 323
rect 228 322 229 323
rect 227 322 228 323
rect 226 322 227 323
rect 225 322 226 323
rect 224 322 225 323
rect 223 322 224 323
rect 222 322 223 323
rect 221 322 222 323
rect 220 322 221 323
rect 219 322 220 323
rect 218 322 219 323
rect 217 322 218 323
rect 216 322 217 323
rect 215 322 216 323
rect 214 322 215 323
rect 213 322 214 323
rect 212 322 213 323
rect 211 322 212 323
rect 210 322 211 323
rect 209 322 210 323
rect 208 322 209 323
rect 207 322 208 323
rect 206 322 207 323
rect 205 322 206 323
rect 204 322 205 323
rect 203 322 204 323
rect 202 322 203 323
rect 201 322 202 323
rect 200 322 201 323
rect 199 322 200 323
rect 198 322 199 323
rect 197 322 198 323
rect 196 322 197 323
rect 195 322 196 323
rect 194 322 195 323
rect 193 322 194 323
rect 192 322 193 323
rect 142 322 143 323
rect 141 322 142 323
rect 140 322 141 323
rect 139 322 140 323
rect 138 322 139 323
rect 137 322 138 323
rect 136 322 137 323
rect 135 322 136 323
rect 134 322 135 323
rect 133 322 134 323
rect 132 322 133 323
rect 131 322 132 323
rect 130 322 131 323
rect 129 322 130 323
rect 128 322 129 323
rect 127 322 128 323
rect 126 322 127 323
rect 125 322 126 323
rect 124 322 125 323
rect 123 322 124 323
rect 122 322 123 323
rect 121 322 122 323
rect 120 322 121 323
rect 119 322 120 323
rect 118 322 119 323
rect 117 322 118 323
rect 116 322 117 323
rect 115 322 116 323
rect 114 322 115 323
rect 113 322 114 323
rect 112 322 113 323
rect 111 322 112 323
rect 110 322 111 323
rect 109 322 110 323
rect 108 322 109 323
rect 107 322 108 323
rect 106 322 107 323
rect 105 322 106 323
rect 104 322 105 323
rect 103 322 104 323
rect 102 322 103 323
rect 101 322 102 323
rect 100 322 101 323
rect 99 322 100 323
rect 98 322 99 323
rect 79 322 80 323
rect 78 322 79 323
rect 77 322 78 323
rect 76 322 77 323
rect 75 322 76 323
rect 74 322 75 323
rect 73 322 74 323
rect 72 322 73 323
rect 71 322 72 323
rect 70 322 71 323
rect 69 322 70 323
rect 68 322 69 323
rect 67 322 68 323
rect 66 322 67 323
rect 65 322 66 323
rect 64 322 65 323
rect 63 322 64 323
rect 62 322 63 323
rect 61 322 62 323
rect 60 322 61 323
rect 59 322 60 323
rect 58 322 59 323
rect 57 322 58 323
rect 56 322 57 323
rect 55 322 56 323
rect 54 322 55 323
rect 53 322 54 323
rect 52 322 53 323
rect 51 322 52 323
rect 50 322 51 323
rect 49 322 50 323
rect 37 322 38 323
rect 36 322 37 323
rect 35 322 36 323
rect 34 322 35 323
rect 33 322 34 323
rect 32 322 33 323
rect 31 322 32 323
rect 30 322 31 323
rect 29 322 30 323
rect 28 322 29 323
rect 27 322 28 323
rect 26 322 27 323
rect 25 322 26 323
rect 24 322 25 323
rect 23 322 24 323
rect 22 322 23 323
rect 21 322 22 323
rect 20 322 21 323
rect 19 322 20 323
rect 482 323 483 324
rect 481 323 482 324
rect 480 323 481 324
rect 479 323 480 324
rect 478 323 479 324
rect 477 323 478 324
rect 476 323 477 324
rect 475 323 476 324
rect 474 323 475 324
rect 473 323 474 324
rect 472 323 473 324
rect 471 323 472 324
rect 470 323 471 324
rect 469 323 470 324
rect 468 323 469 324
rect 462 323 463 324
rect 441 323 442 324
rect 440 323 441 324
rect 439 323 440 324
rect 399 323 400 324
rect 398 323 399 324
rect 397 323 398 324
rect 228 323 229 324
rect 227 323 228 324
rect 226 323 227 324
rect 225 323 226 324
rect 224 323 225 324
rect 223 323 224 324
rect 222 323 223 324
rect 221 323 222 324
rect 220 323 221 324
rect 219 323 220 324
rect 218 323 219 324
rect 217 323 218 324
rect 216 323 217 324
rect 215 323 216 324
rect 214 323 215 324
rect 213 323 214 324
rect 212 323 213 324
rect 211 323 212 324
rect 210 323 211 324
rect 209 323 210 324
rect 208 323 209 324
rect 207 323 208 324
rect 206 323 207 324
rect 205 323 206 324
rect 204 323 205 324
rect 203 323 204 324
rect 202 323 203 324
rect 201 323 202 324
rect 200 323 201 324
rect 199 323 200 324
rect 198 323 199 324
rect 197 323 198 324
rect 196 323 197 324
rect 195 323 196 324
rect 144 323 145 324
rect 143 323 144 324
rect 142 323 143 324
rect 141 323 142 324
rect 140 323 141 324
rect 139 323 140 324
rect 138 323 139 324
rect 137 323 138 324
rect 136 323 137 324
rect 135 323 136 324
rect 134 323 135 324
rect 133 323 134 324
rect 132 323 133 324
rect 131 323 132 324
rect 130 323 131 324
rect 129 323 130 324
rect 128 323 129 324
rect 127 323 128 324
rect 126 323 127 324
rect 125 323 126 324
rect 124 323 125 324
rect 123 323 124 324
rect 122 323 123 324
rect 121 323 122 324
rect 120 323 121 324
rect 119 323 120 324
rect 118 323 119 324
rect 117 323 118 324
rect 116 323 117 324
rect 115 323 116 324
rect 114 323 115 324
rect 113 323 114 324
rect 112 323 113 324
rect 111 323 112 324
rect 110 323 111 324
rect 109 323 110 324
rect 108 323 109 324
rect 107 323 108 324
rect 106 323 107 324
rect 105 323 106 324
rect 104 323 105 324
rect 103 323 104 324
rect 102 323 103 324
rect 101 323 102 324
rect 100 323 101 324
rect 99 323 100 324
rect 80 323 81 324
rect 79 323 80 324
rect 78 323 79 324
rect 77 323 78 324
rect 76 323 77 324
rect 75 323 76 324
rect 74 323 75 324
rect 73 323 74 324
rect 72 323 73 324
rect 71 323 72 324
rect 70 323 71 324
rect 69 323 70 324
rect 68 323 69 324
rect 67 323 68 324
rect 66 323 67 324
rect 65 323 66 324
rect 64 323 65 324
rect 63 323 64 324
rect 62 323 63 324
rect 61 323 62 324
rect 60 323 61 324
rect 59 323 60 324
rect 58 323 59 324
rect 57 323 58 324
rect 56 323 57 324
rect 55 323 56 324
rect 54 323 55 324
rect 53 323 54 324
rect 52 323 53 324
rect 51 323 52 324
rect 50 323 51 324
rect 49 323 50 324
rect 37 323 38 324
rect 36 323 37 324
rect 35 323 36 324
rect 34 323 35 324
rect 33 323 34 324
rect 32 323 33 324
rect 31 323 32 324
rect 30 323 31 324
rect 29 323 30 324
rect 28 323 29 324
rect 27 323 28 324
rect 26 323 27 324
rect 25 323 26 324
rect 24 323 25 324
rect 23 323 24 324
rect 22 323 23 324
rect 21 323 22 324
rect 20 323 21 324
rect 482 324 483 325
rect 481 324 482 325
rect 480 324 481 325
rect 479 324 480 325
rect 478 324 479 325
rect 477 324 478 325
rect 476 324 477 325
rect 475 324 476 325
rect 474 324 475 325
rect 473 324 474 325
rect 472 324 473 325
rect 471 324 472 325
rect 470 324 471 325
rect 441 324 442 325
rect 440 324 441 325
rect 439 324 440 325
rect 399 324 400 325
rect 398 324 399 325
rect 397 324 398 325
rect 221 324 222 325
rect 220 324 221 325
rect 219 324 220 325
rect 218 324 219 325
rect 217 324 218 325
rect 216 324 217 325
rect 215 324 216 325
rect 214 324 215 325
rect 213 324 214 325
rect 212 324 213 325
rect 211 324 212 325
rect 210 324 211 325
rect 209 324 210 325
rect 208 324 209 325
rect 207 324 208 325
rect 206 324 207 325
rect 205 324 206 325
rect 204 324 205 325
rect 203 324 204 325
rect 202 324 203 325
rect 145 324 146 325
rect 144 324 145 325
rect 143 324 144 325
rect 142 324 143 325
rect 141 324 142 325
rect 140 324 141 325
rect 139 324 140 325
rect 138 324 139 325
rect 137 324 138 325
rect 136 324 137 325
rect 135 324 136 325
rect 134 324 135 325
rect 133 324 134 325
rect 132 324 133 325
rect 131 324 132 325
rect 130 324 131 325
rect 129 324 130 325
rect 128 324 129 325
rect 127 324 128 325
rect 126 324 127 325
rect 125 324 126 325
rect 124 324 125 325
rect 123 324 124 325
rect 122 324 123 325
rect 121 324 122 325
rect 120 324 121 325
rect 119 324 120 325
rect 118 324 119 325
rect 117 324 118 325
rect 116 324 117 325
rect 115 324 116 325
rect 114 324 115 325
rect 113 324 114 325
rect 112 324 113 325
rect 111 324 112 325
rect 110 324 111 325
rect 109 324 110 325
rect 108 324 109 325
rect 107 324 108 325
rect 106 324 107 325
rect 105 324 106 325
rect 104 324 105 325
rect 103 324 104 325
rect 102 324 103 325
rect 101 324 102 325
rect 100 324 101 325
rect 99 324 100 325
rect 81 324 82 325
rect 80 324 81 325
rect 79 324 80 325
rect 78 324 79 325
rect 77 324 78 325
rect 76 324 77 325
rect 75 324 76 325
rect 74 324 75 325
rect 73 324 74 325
rect 72 324 73 325
rect 71 324 72 325
rect 70 324 71 325
rect 69 324 70 325
rect 68 324 69 325
rect 67 324 68 325
rect 66 324 67 325
rect 65 324 66 325
rect 64 324 65 325
rect 63 324 64 325
rect 62 324 63 325
rect 61 324 62 325
rect 60 324 61 325
rect 59 324 60 325
rect 58 324 59 325
rect 57 324 58 325
rect 56 324 57 325
rect 55 324 56 325
rect 54 324 55 325
rect 53 324 54 325
rect 52 324 53 325
rect 51 324 52 325
rect 50 324 51 325
rect 38 324 39 325
rect 37 324 38 325
rect 36 324 37 325
rect 35 324 36 325
rect 34 324 35 325
rect 33 324 34 325
rect 32 324 33 325
rect 31 324 32 325
rect 30 324 31 325
rect 29 324 30 325
rect 28 324 29 325
rect 27 324 28 325
rect 26 324 27 325
rect 25 324 26 325
rect 24 324 25 325
rect 23 324 24 325
rect 22 324 23 325
rect 21 324 22 325
rect 20 324 21 325
rect 482 325 483 326
rect 481 325 482 326
rect 480 325 481 326
rect 479 325 480 326
rect 478 325 479 326
rect 477 325 478 326
rect 476 325 477 326
rect 475 325 476 326
rect 474 325 475 326
rect 473 325 474 326
rect 472 325 473 326
rect 471 325 472 326
rect 147 325 148 326
rect 146 325 147 326
rect 145 325 146 326
rect 144 325 145 326
rect 143 325 144 326
rect 142 325 143 326
rect 141 325 142 326
rect 140 325 141 326
rect 139 325 140 326
rect 138 325 139 326
rect 137 325 138 326
rect 136 325 137 326
rect 135 325 136 326
rect 134 325 135 326
rect 133 325 134 326
rect 132 325 133 326
rect 131 325 132 326
rect 130 325 131 326
rect 129 325 130 326
rect 128 325 129 326
rect 127 325 128 326
rect 126 325 127 326
rect 125 325 126 326
rect 124 325 125 326
rect 123 325 124 326
rect 122 325 123 326
rect 121 325 122 326
rect 120 325 121 326
rect 119 325 120 326
rect 118 325 119 326
rect 117 325 118 326
rect 116 325 117 326
rect 115 325 116 326
rect 114 325 115 326
rect 113 325 114 326
rect 112 325 113 326
rect 111 325 112 326
rect 110 325 111 326
rect 109 325 110 326
rect 108 325 109 326
rect 107 325 108 326
rect 106 325 107 326
rect 105 325 106 326
rect 104 325 105 326
rect 103 325 104 326
rect 102 325 103 326
rect 101 325 102 326
rect 100 325 101 326
rect 81 325 82 326
rect 80 325 81 326
rect 79 325 80 326
rect 78 325 79 326
rect 77 325 78 326
rect 76 325 77 326
rect 75 325 76 326
rect 74 325 75 326
rect 73 325 74 326
rect 72 325 73 326
rect 71 325 72 326
rect 70 325 71 326
rect 69 325 70 326
rect 68 325 69 326
rect 67 325 68 326
rect 66 325 67 326
rect 65 325 66 326
rect 64 325 65 326
rect 63 325 64 326
rect 62 325 63 326
rect 61 325 62 326
rect 60 325 61 326
rect 59 325 60 326
rect 58 325 59 326
rect 57 325 58 326
rect 56 325 57 326
rect 55 325 56 326
rect 54 325 55 326
rect 53 325 54 326
rect 52 325 53 326
rect 51 325 52 326
rect 50 325 51 326
rect 38 325 39 326
rect 37 325 38 326
rect 36 325 37 326
rect 35 325 36 326
rect 34 325 35 326
rect 33 325 34 326
rect 32 325 33 326
rect 31 325 32 326
rect 30 325 31 326
rect 29 325 30 326
rect 28 325 29 326
rect 27 325 28 326
rect 26 325 27 326
rect 25 325 26 326
rect 24 325 25 326
rect 23 325 24 326
rect 22 325 23 326
rect 21 325 22 326
rect 482 326 483 327
rect 481 326 482 327
rect 480 326 481 327
rect 479 326 480 327
rect 478 326 479 327
rect 477 326 478 327
rect 476 326 477 327
rect 475 326 476 327
rect 474 326 475 327
rect 473 326 474 327
rect 472 326 473 327
rect 471 326 472 327
rect 470 326 471 327
rect 149 326 150 327
rect 148 326 149 327
rect 147 326 148 327
rect 146 326 147 327
rect 145 326 146 327
rect 144 326 145 327
rect 143 326 144 327
rect 142 326 143 327
rect 141 326 142 327
rect 140 326 141 327
rect 139 326 140 327
rect 138 326 139 327
rect 137 326 138 327
rect 136 326 137 327
rect 135 326 136 327
rect 134 326 135 327
rect 133 326 134 327
rect 132 326 133 327
rect 131 326 132 327
rect 130 326 131 327
rect 129 326 130 327
rect 128 326 129 327
rect 127 326 128 327
rect 126 326 127 327
rect 125 326 126 327
rect 124 326 125 327
rect 123 326 124 327
rect 122 326 123 327
rect 121 326 122 327
rect 120 326 121 327
rect 119 326 120 327
rect 118 326 119 327
rect 117 326 118 327
rect 116 326 117 327
rect 115 326 116 327
rect 114 326 115 327
rect 113 326 114 327
rect 112 326 113 327
rect 111 326 112 327
rect 110 326 111 327
rect 109 326 110 327
rect 108 326 109 327
rect 107 326 108 327
rect 106 326 107 327
rect 105 326 106 327
rect 104 326 105 327
rect 103 326 104 327
rect 102 326 103 327
rect 101 326 102 327
rect 82 326 83 327
rect 81 326 82 327
rect 80 326 81 327
rect 79 326 80 327
rect 78 326 79 327
rect 77 326 78 327
rect 76 326 77 327
rect 75 326 76 327
rect 74 326 75 327
rect 73 326 74 327
rect 72 326 73 327
rect 71 326 72 327
rect 70 326 71 327
rect 69 326 70 327
rect 68 326 69 327
rect 67 326 68 327
rect 66 326 67 327
rect 65 326 66 327
rect 64 326 65 327
rect 63 326 64 327
rect 62 326 63 327
rect 61 326 62 327
rect 60 326 61 327
rect 59 326 60 327
rect 58 326 59 327
rect 57 326 58 327
rect 56 326 57 327
rect 55 326 56 327
rect 54 326 55 327
rect 53 326 54 327
rect 52 326 53 327
rect 51 326 52 327
rect 50 326 51 327
rect 38 326 39 327
rect 37 326 38 327
rect 36 326 37 327
rect 35 326 36 327
rect 34 326 35 327
rect 33 326 34 327
rect 32 326 33 327
rect 31 326 32 327
rect 30 326 31 327
rect 29 326 30 327
rect 28 326 29 327
rect 27 326 28 327
rect 26 326 27 327
rect 25 326 26 327
rect 24 326 25 327
rect 23 326 24 327
rect 22 326 23 327
rect 482 327 483 328
rect 471 327 472 328
rect 470 327 471 328
rect 469 327 470 328
rect 468 327 469 328
rect 462 327 463 328
rect 151 327 152 328
rect 150 327 151 328
rect 149 327 150 328
rect 148 327 149 328
rect 147 327 148 328
rect 146 327 147 328
rect 145 327 146 328
rect 144 327 145 328
rect 143 327 144 328
rect 142 327 143 328
rect 141 327 142 328
rect 140 327 141 328
rect 139 327 140 328
rect 138 327 139 328
rect 137 327 138 328
rect 136 327 137 328
rect 135 327 136 328
rect 134 327 135 328
rect 133 327 134 328
rect 132 327 133 328
rect 131 327 132 328
rect 130 327 131 328
rect 129 327 130 328
rect 128 327 129 328
rect 127 327 128 328
rect 126 327 127 328
rect 125 327 126 328
rect 124 327 125 328
rect 123 327 124 328
rect 122 327 123 328
rect 121 327 122 328
rect 120 327 121 328
rect 119 327 120 328
rect 118 327 119 328
rect 117 327 118 328
rect 116 327 117 328
rect 115 327 116 328
rect 114 327 115 328
rect 113 327 114 328
rect 112 327 113 328
rect 111 327 112 328
rect 110 327 111 328
rect 109 327 110 328
rect 108 327 109 328
rect 107 327 108 328
rect 106 327 107 328
rect 105 327 106 328
rect 104 327 105 328
rect 103 327 104 328
rect 102 327 103 328
rect 82 327 83 328
rect 81 327 82 328
rect 80 327 81 328
rect 79 327 80 328
rect 78 327 79 328
rect 77 327 78 328
rect 76 327 77 328
rect 75 327 76 328
rect 74 327 75 328
rect 73 327 74 328
rect 72 327 73 328
rect 71 327 72 328
rect 70 327 71 328
rect 69 327 70 328
rect 68 327 69 328
rect 67 327 68 328
rect 66 327 67 328
rect 65 327 66 328
rect 64 327 65 328
rect 63 327 64 328
rect 62 327 63 328
rect 61 327 62 328
rect 60 327 61 328
rect 59 327 60 328
rect 58 327 59 328
rect 57 327 58 328
rect 56 327 57 328
rect 55 327 56 328
rect 54 327 55 328
rect 53 327 54 328
rect 52 327 53 328
rect 51 327 52 328
rect 39 327 40 328
rect 38 327 39 328
rect 37 327 38 328
rect 36 327 37 328
rect 35 327 36 328
rect 34 327 35 328
rect 33 327 34 328
rect 32 327 33 328
rect 31 327 32 328
rect 30 327 31 328
rect 29 327 30 328
rect 28 327 29 328
rect 27 327 28 328
rect 26 327 27 328
rect 25 327 26 328
rect 24 327 25 328
rect 23 327 24 328
rect 482 328 483 329
rect 469 328 470 329
rect 468 328 469 329
rect 467 328 468 329
rect 466 328 467 329
rect 462 328 463 329
rect 153 328 154 329
rect 152 328 153 329
rect 151 328 152 329
rect 150 328 151 329
rect 149 328 150 329
rect 148 328 149 329
rect 147 328 148 329
rect 146 328 147 329
rect 145 328 146 329
rect 144 328 145 329
rect 143 328 144 329
rect 142 328 143 329
rect 141 328 142 329
rect 140 328 141 329
rect 139 328 140 329
rect 138 328 139 329
rect 137 328 138 329
rect 136 328 137 329
rect 135 328 136 329
rect 134 328 135 329
rect 133 328 134 329
rect 132 328 133 329
rect 131 328 132 329
rect 130 328 131 329
rect 129 328 130 329
rect 128 328 129 329
rect 127 328 128 329
rect 126 328 127 329
rect 125 328 126 329
rect 124 328 125 329
rect 123 328 124 329
rect 122 328 123 329
rect 121 328 122 329
rect 120 328 121 329
rect 119 328 120 329
rect 118 328 119 329
rect 117 328 118 329
rect 116 328 117 329
rect 115 328 116 329
rect 114 328 115 329
rect 113 328 114 329
rect 112 328 113 329
rect 111 328 112 329
rect 110 328 111 329
rect 109 328 110 329
rect 108 328 109 329
rect 107 328 108 329
rect 106 328 107 329
rect 105 328 106 329
rect 104 328 105 329
rect 103 328 104 329
rect 102 328 103 329
rect 83 328 84 329
rect 82 328 83 329
rect 81 328 82 329
rect 80 328 81 329
rect 79 328 80 329
rect 78 328 79 329
rect 77 328 78 329
rect 76 328 77 329
rect 75 328 76 329
rect 74 328 75 329
rect 73 328 74 329
rect 72 328 73 329
rect 71 328 72 329
rect 70 328 71 329
rect 69 328 70 329
rect 68 328 69 329
rect 67 328 68 329
rect 66 328 67 329
rect 65 328 66 329
rect 64 328 65 329
rect 63 328 64 329
rect 62 328 63 329
rect 61 328 62 329
rect 60 328 61 329
rect 59 328 60 329
rect 58 328 59 329
rect 57 328 58 329
rect 56 328 57 329
rect 55 328 56 329
rect 54 328 55 329
rect 53 328 54 329
rect 52 328 53 329
rect 51 328 52 329
rect 39 328 40 329
rect 38 328 39 329
rect 37 328 38 329
rect 36 328 37 329
rect 35 328 36 329
rect 34 328 35 329
rect 33 328 34 329
rect 32 328 33 329
rect 31 328 32 329
rect 30 328 31 329
rect 29 328 30 329
rect 28 328 29 329
rect 27 328 28 329
rect 26 328 27 329
rect 25 328 26 329
rect 24 328 25 329
rect 482 329 483 330
rect 467 329 468 330
rect 466 329 467 330
rect 465 329 466 330
rect 464 329 465 330
rect 463 329 464 330
rect 462 329 463 330
rect 155 329 156 330
rect 154 329 155 330
rect 153 329 154 330
rect 152 329 153 330
rect 151 329 152 330
rect 150 329 151 330
rect 149 329 150 330
rect 148 329 149 330
rect 147 329 148 330
rect 146 329 147 330
rect 145 329 146 330
rect 144 329 145 330
rect 143 329 144 330
rect 142 329 143 330
rect 141 329 142 330
rect 140 329 141 330
rect 139 329 140 330
rect 138 329 139 330
rect 137 329 138 330
rect 136 329 137 330
rect 135 329 136 330
rect 134 329 135 330
rect 133 329 134 330
rect 132 329 133 330
rect 131 329 132 330
rect 130 329 131 330
rect 129 329 130 330
rect 128 329 129 330
rect 127 329 128 330
rect 126 329 127 330
rect 125 329 126 330
rect 124 329 125 330
rect 123 329 124 330
rect 122 329 123 330
rect 121 329 122 330
rect 120 329 121 330
rect 119 329 120 330
rect 118 329 119 330
rect 117 329 118 330
rect 116 329 117 330
rect 115 329 116 330
rect 114 329 115 330
rect 113 329 114 330
rect 112 329 113 330
rect 111 329 112 330
rect 110 329 111 330
rect 109 329 110 330
rect 108 329 109 330
rect 107 329 108 330
rect 106 329 107 330
rect 105 329 106 330
rect 104 329 105 330
rect 103 329 104 330
rect 84 329 85 330
rect 83 329 84 330
rect 82 329 83 330
rect 81 329 82 330
rect 80 329 81 330
rect 79 329 80 330
rect 78 329 79 330
rect 77 329 78 330
rect 76 329 77 330
rect 75 329 76 330
rect 74 329 75 330
rect 73 329 74 330
rect 72 329 73 330
rect 71 329 72 330
rect 70 329 71 330
rect 69 329 70 330
rect 68 329 69 330
rect 67 329 68 330
rect 66 329 67 330
rect 65 329 66 330
rect 64 329 65 330
rect 63 329 64 330
rect 62 329 63 330
rect 61 329 62 330
rect 60 329 61 330
rect 59 329 60 330
rect 58 329 59 330
rect 57 329 58 330
rect 56 329 57 330
rect 55 329 56 330
rect 54 329 55 330
rect 53 329 54 330
rect 52 329 53 330
rect 39 329 40 330
rect 38 329 39 330
rect 37 329 38 330
rect 36 329 37 330
rect 35 329 36 330
rect 34 329 35 330
rect 33 329 34 330
rect 32 329 33 330
rect 31 329 32 330
rect 30 329 31 330
rect 29 329 30 330
rect 28 329 29 330
rect 27 329 28 330
rect 26 329 27 330
rect 25 329 26 330
rect 24 329 25 330
rect 465 330 466 331
rect 464 330 465 331
rect 463 330 464 331
rect 462 330 463 331
rect 158 330 159 331
rect 157 330 158 331
rect 156 330 157 331
rect 155 330 156 331
rect 154 330 155 331
rect 153 330 154 331
rect 152 330 153 331
rect 151 330 152 331
rect 150 330 151 331
rect 149 330 150 331
rect 148 330 149 331
rect 147 330 148 331
rect 146 330 147 331
rect 145 330 146 331
rect 144 330 145 331
rect 143 330 144 331
rect 142 330 143 331
rect 141 330 142 331
rect 140 330 141 331
rect 139 330 140 331
rect 138 330 139 331
rect 137 330 138 331
rect 136 330 137 331
rect 135 330 136 331
rect 134 330 135 331
rect 133 330 134 331
rect 132 330 133 331
rect 131 330 132 331
rect 130 330 131 331
rect 129 330 130 331
rect 128 330 129 331
rect 127 330 128 331
rect 126 330 127 331
rect 125 330 126 331
rect 124 330 125 331
rect 123 330 124 331
rect 122 330 123 331
rect 121 330 122 331
rect 120 330 121 331
rect 119 330 120 331
rect 118 330 119 331
rect 117 330 118 331
rect 116 330 117 331
rect 115 330 116 331
rect 114 330 115 331
rect 113 330 114 331
rect 112 330 113 331
rect 111 330 112 331
rect 110 330 111 331
rect 109 330 110 331
rect 108 330 109 331
rect 107 330 108 331
rect 106 330 107 331
rect 105 330 106 331
rect 104 330 105 331
rect 84 330 85 331
rect 83 330 84 331
rect 82 330 83 331
rect 81 330 82 331
rect 80 330 81 331
rect 79 330 80 331
rect 78 330 79 331
rect 77 330 78 331
rect 76 330 77 331
rect 75 330 76 331
rect 74 330 75 331
rect 73 330 74 331
rect 72 330 73 331
rect 71 330 72 331
rect 70 330 71 331
rect 69 330 70 331
rect 68 330 69 331
rect 67 330 68 331
rect 66 330 67 331
rect 65 330 66 331
rect 64 330 65 331
rect 63 330 64 331
rect 62 330 63 331
rect 61 330 62 331
rect 60 330 61 331
rect 59 330 60 331
rect 58 330 59 331
rect 57 330 58 331
rect 56 330 57 331
rect 55 330 56 331
rect 54 330 55 331
rect 53 330 54 331
rect 52 330 53 331
rect 40 330 41 331
rect 39 330 40 331
rect 38 330 39 331
rect 37 330 38 331
rect 36 330 37 331
rect 35 330 36 331
rect 34 330 35 331
rect 33 330 34 331
rect 32 330 33 331
rect 31 330 32 331
rect 30 330 31 331
rect 29 330 30 331
rect 28 330 29 331
rect 27 330 28 331
rect 26 330 27 331
rect 25 330 26 331
rect 464 331 465 332
rect 463 331 464 332
rect 462 331 463 332
rect 160 331 161 332
rect 159 331 160 332
rect 158 331 159 332
rect 157 331 158 332
rect 156 331 157 332
rect 155 331 156 332
rect 154 331 155 332
rect 153 331 154 332
rect 152 331 153 332
rect 151 331 152 332
rect 150 331 151 332
rect 149 331 150 332
rect 148 331 149 332
rect 147 331 148 332
rect 146 331 147 332
rect 145 331 146 332
rect 144 331 145 332
rect 143 331 144 332
rect 142 331 143 332
rect 141 331 142 332
rect 140 331 141 332
rect 139 331 140 332
rect 138 331 139 332
rect 137 331 138 332
rect 136 331 137 332
rect 135 331 136 332
rect 134 331 135 332
rect 133 331 134 332
rect 132 331 133 332
rect 131 331 132 332
rect 130 331 131 332
rect 129 331 130 332
rect 128 331 129 332
rect 127 331 128 332
rect 126 331 127 332
rect 125 331 126 332
rect 124 331 125 332
rect 123 331 124 332
rect 122 331 123 332
rect 121 331 122 332
rect 120 331 121 332
rect 119 331 120 332
rect 118 331 119 332
rect 117 331 118 332
rect 116 331 117 332
rect 115 331 116 332
rect 114 331 115 332
rect 113 331 114 332
rect 112 331 113 332
rect 111 331 112 332
rect 110 331 111 332
rect 109 331 110 332
rect 108 331 109 332
rect 107 331 108 332
rect 106 331 107 332
rect 105 331 106 332
rect 85 331 86 332
rect 84 331 85 332
rect 83 331 84 332
rect 82 331 83 332
rect 81 331 82 332
rect 80 331 81 332
rect 79 331 80 332
rect 78 331 79 332
rect 77 331 78 332
rect 76 331 77 332
rect 75 331 76 332
rect 74 331 75 332
rect 73 331 74 332
rect 72 331 73 332
rect 71 331 72 332
rect 70 331 71 332
rect 69 331 70 332
rect 68 331 69 332
rect 67 331 68 332
rect 66 331 67 332
rect 65 331 66 332
rect 64 331 65 332
rect 63 331 64 332
rect 62 331 63 332
rect 61 331 62 332
rect 60 331 61 332
rect 59 331 60 332
rect 58 331 59 332
rect 57 331 58 332
rect 56 331 57 332
rect 55 331 56 332
rect 54 331 55 332
rect 53 331 54 332
rect 52 331 53 332
rect 40 331 41 332
rect 39 331 40 332
rect 38 331 39 332
rect 37 331 38 332
rect 36 331 37 332
rect 35 331 36 332
rect 34 331 35 332
rect 33 331 34 332
rect 32 331 33 332
rect 31 331 32 332
rect 30 331 31 332
rect 29 331 30 332
rect 28 331 29 332
rect 27 331 28 332
rect 26 331 27 332
rect 463 332 464 333
rect 462 332 463 333
rect 163 332 164 333
rect 162 332 163 333
rect 161 332 162 333
rect 160 332 161 333
rect 159 332 160 333
rect 158 332 159 333
rect 157 332 158 333
rect 156 332 157 333
rect 155 332 156 333
rect 154 332 155 333
rect 153 332 154 333
rect 152 332 153 333
rect 151 332 152 333
rect 150 332 151 333
rect 149 332 150 333
rect 148 332 149 333
rect 147 332 148 333
rect 146 332 147 333
rect 145 332 146 333
rect 144 332 145 333
rect 143 332 144 333
rect 142 332 143 333
rect 141 332 142 333
rect 140 332 141 333
rect 139 332 140 333
rect 138 332 139 333
rect 137 332 138 333
rect 136 332 137 333
rect 135 332 136 333
rect 134 332 135 333
rect 133 332 134 333
rect 132 332 133 333
rect 131 332 132 333
rect 130 332 131 333
rect 129 332 130 333
rect 128 332 129 333
rect 127 332 128 333
rect 126 332 127 333
rect 125 332 126 333
rect 124 332 125 333
rect 123 332 124 333
rect 122 332 123 333
rect 121 332 122 333
rect 120 332 121 333
rect 119 332 120 333
rect 118 332 119 333
rect 117 332 118 333
rect 116 332 117 333
rect 115 332 116 333
rect 114 332 115 333
rect 113 332 114 333
rect 112 332 113 333
rect 111 332 112 333
rect 110 332 111 333
rect 109 332 110 333
rect 108 332 109 333
rect 107 332 108 333
rect 106 332 107 333
rect 86 332 87 333
rect 85 332 86 333
rect 84 332 85 333
rect 83 332 84 333
rect 82 332 83 333
rect 81 332 82 333
rect 80 332 81 333
rect 79 332 80 333
rect 78 332 79 333
rect 77 332 78 333
rect 76 332 77 333
rect 75 332 76 333
rect 74 332 75 333
rect 73 332 74 333
rect 72 332 73 333
rect 71 332 72 333
rect 70 332 71 333
rect 69 332 70 333
rect 68 332 69 333
rect 67 332 68 333
rect 66 332 67 333
rect 65 332 66 333
rect 64 332 65 333
rect 63 332 64 333
rect 62 332 63 333
rect 61 332 62 333
rect 60 332 61 333
rect 59 332 60 333
rect 58 332 59 333
rect 57 332 58 333
rect 56 332 57 333
rect 55 332 56 333
rect 54 332 55 333
rect 53 332 54 333
rect 41 332 42 333
rect 40 332 41 333
rect 39 332 40 333
rect 38 332 39 333
rect 37 332 38 333
rect 36 332 37 333
rect 35 332 36 333
rect 34 332 35 333
rect 33 332 34 333
rect 32 332 33 333
rect 31 332 32 333
rect 30 332 31 333
rect 29 332 30 333
rect 28 332 29 333
rect 27 332 28 333
rect 462 333 463 334
rect 441 333 442 334
rect 440 333 441 334
rect 439 333 440 334
rect 166 333 167 334
rect 165 333 166 334
rect 164 333 165 334
rect 163 333 164 334
rect 162 333 163 334
rect 161 333 162 334
rect 160 333 161 334
rect 159 333 160 334
rect 158 333 159 334
rect 157 333 158 334
rect 156 333 157 334
rect 155 333 156 334
rect 154 333 155 334
rect 153 333 154 334
rect 152 333 153 334
rect 151 333 152 334
rect 150 333 151 334
rect 149 333 150 334
rect 148 333 149 334
rect 147 333 148 334
rect 146 333 147 334
rect 145 333 146 334
rect 144 333 145 334
rect 143 333 144 334
rect 142 333 143 334
rect 141 333 142 334
rect 140 333 141 334
rect 139 333 140 334
rect 138 333 139 334
rect 137 333 138 334
rect 136 333 137 334
rect 135 333 136 334
rect 134 333 135 334
rect 133 333 134 334
rect 132 333 133 334
rect 131 333 132 334
rect 130 333 131 334
rect 129 333 130 334
rect 128 333 129 334
rect 127 333 128 334
rect 126 333 127 334
rect 125 333 126 334
rect 124 333 125 334
rect 123 333 124 334
rect 122 333 123 334
rect 121 333 122 334
rect 120 333 121 334
rect 119 333 120 334
rect 118 333 119 334
rect 117 333 118 334
rect 116 333 117 334
rect 115 333 116 334
rect 114 333 115 334
rect 113 333 114 334
rect 112 333 113 334
rect 111 333 112 334
rect 110 333 111 334
rect 109 333 110 334
rect 108 333 109 334
rect 107 333 108 334
rect 106 333 107 334
rect 86 333 87 334
rect 85 333 86 334
rect 84 333 85 334
rect 83 333 84 334
rect 82 333 83 334
rect 81 333 82 334
rect 80 333 81 334
rect 79 333 80 334
rect 78 333 79 334
rect 77 333 78 334
rect 76 333 77 334
rect 75 333 76 334
rect 74 333 75 334
rect 73 333 74 334
rect 72 333 73 334
rect 71 333 72 334
rect 70 333 71 334
rect 69 333 70 334
rect 68 333 69 334
rect 67 333 68 334
rect 66 333 67 334
rect 65 333 66 334
rect 64 333 65 334
rect 63 333 64 334
rect 62 333 63 334
rect 61 333 62 334
rect 60 333 61 334
rect 59 333 60 334
rect 58 333 59 334
rect 57 333 58 334
rect 56 333 57 334
rect 55 333 56 334
rect 54 333 55 334
rect 53 333 54 334
rect 41 333 42 334
rect 40 333 41 334
rect 39 333 40 334
rect 38 333 39 334
rect 37 333 38 334
rect 36 333 37 334
rect 35 333 36 334
rect 34 333 35 334
rect 33 333 34 334
rect 32 333 33 334
rect 31 333 32 334
rect 30 333 31 334
rect 29 333 30 334
rect 28 333 29 334
rect 462 334 463 335
rect 441 334 442 335
rect 440 334 441 335
rect 439 334 440 335
rect 399 334 400 335
rect 398 334 399 335
rect 397 334 398 335
rect 169 334 170 335
rect 168 334 169 335
rect 167 334 168 335
rect 166 334 167 335
rect 165 334 166 335
rect 164 334 165 335
rect 163 334 164 335
rect 162 334 163 335
rect 161 334 162 335
rect 160 334 161 335
rect 159 334 160 335
rect 158 334 159 335
rect 157 334 158 335
rect 156 334 157 335
rect 155 334 156 335
rect 154 334 155 335
rect 153 334 154 335
rect 152 334 153 335
rect 151 334 152 335
rect 150 334 151 335
rect 149 334 150 335
rect 148 334 149 335
rect 147 334 148 335
rect 146 334 147 335
rect 145 334 146 335
rect 144 334 145 335
rect 143 334 144 335
rect 142 334 143 335
rect 141 334 142 335
rect 140 334 141 335
rect 139 334 140 335
rect 138 334 139 335
rect 137 334 138 335
rect 136 334 137 335
rect 135 334 136 335
rect 134 334 135 335
rect 133 334 134 335
rect 132 334 133 335
rect 131 334 132 335
rect 130 334 131 335
rect 129 334 130 335
rect 128 334 129 335
rect 127 334 128 335
rect 126 334 127 335
rect 125 334 126 335
rect 124 334 125 335
rect 123 334 124 335
rect 122 334 123 335
rect 121 334 122 335
rect 120 334 121 335
rect 119 334 120 335
rect 118 334 119 335
rect 117 334 118 335
rect 116 334 117 335
rect 115 334 116 335
rect 114 334 115 335
rect 113 334 114 335
rect 112 334 113 335
rect 111 334 112 335
rect 110 334 111 335
rect 109 334 110 335
rect 108 334 109 335
rect 107 334 108 335
rect 87 334 88 335
rect 86 334 87 335
rect 85 334 86 335
rect 84 334 85 335
rect 83 334 84 335
rect 82 334 83 335
rect 81 334 82 335
rect 80 334 81 335
rect 79 334 80 335
rect 78 334 79 335
rect 77 334 78 335
rect 76 334 77 335
rect 75 334 76 335
rect 74 334 75 335
rect 73 334 74 335
rect 72 334 73 335
rect 71 334 72 335
rect 70 334 71 335
rect 69 334 70 335
rect 68 334 69 335
rect 67 334 68 335
rect 66 334 67 335
rect 65 334 66 335
rect 64 334 65 335
rect 63 334 64 335
rect 62 334 63 335
rect 61 334 62 335
rect 60 334 61 335
rect 59 334 60 335
rect 58 334 59 335
rect 57 334 58 335
rect 56 334 57 335
rect 55 334 56 335
rect 54 334 55 335
rect 53 334 54 335
rect 41 334 42 335
rect 40 334 41 335
rect 39 334 40 335
rect 38 334 39 335
rect 37 334 38 335
rect 36 334 37 335
rect 35 334 36 335
rect 34 334 35 335
rect 33 334 34 335
rect 32 334 33 335
rect 31 334 32 335
rect 30 334 31 335
rect 29 334 30 335
rect 441 335 442 336
rect 440 335 441 336
rect 439 335 440 336
rect 399 335 400 336
rect 398 335 399 336
rect 397 335 398 336
rect 172 335 173 336
rect 171 335 172 336
rect 170 335 171 336
rect 169 335 170 336
rect 168 335 169 336
rect 167 335 168 336
rect 166 335 167 336
rect 165 335 166 336
rect 164 335 165 336
rect 163 335 164 336
rect 162 335 163 336
rect 161 335 162 336
rect 160 335 161 336
rect 159 335 160 336
rect 158 335 159 336
rect 157 335 158 336
rect 156 335 157 336
rect 155 335 156 336
rect 154 335 155 336
rect 153 335 154 336
rect 152 335 153 336
rect 151 335 152 336
rect 150 335 151 336
rect 149 335 150 336
rect 148 335 149 336
rect 147 335 148 336
rect 146 335 147 336
rect 145 335 146 336
rect 144 335 145 336
rect 143 335 144 336
rect 142 335 143 336
rect 141 335 142 336
rect 140 335 141 336
rect 139 335 140 336
rect 138 335 139 336
rect 137 335 138 336
rect 136 335 137 336
rect 135 335 136 336
rect 134 335 135 336
rect 133 335 134 336
rect 132 335 133 336
rect 131 335 132 336
rect 130 335 131 336
rect 129 335 130 336
rect 128 335 129 336
rect 127 335 128 336
rect 126 335 127 336
rect 125 335 126 336
rect 124 335 125 336
rect 123 335 124 336
rect 122 335 123 336
rect 121 335 122 336
rect 120 335 121 336
rect 119 335 120 336
rect 118 335 119 336
rect 117 335 118 336
rect 116 335 117 336
rect 115 335 116 336
rect 114 335 115 336
rect 113 335 114 336
rect 112 335 113 336
rect 111 335 112 336
rect 110 335 111 336
rect 109 335 110 336
rect 108 335 109 336
rect 88 335 89 336
rect 87 335 88 336
rect 86 335 87 336
rect 85 335 86 336
rect 84 335 85 336
rect 83 335 84 336
rect 82 335 83 336
rect 81 335 82 336
rect 80 335 81 336
rect 79 335 80 336
rect 78 335 79 336
rect 77 335 78 336
rect 76 335 77 336
rect 75 335 76 336
rect 74 335 75 336
rect 73 335 74 336
rect 72 335 73 336
rect 71 335 72 336
rect 70 335 71 336
rect 69 335 70 336
rect 68 335 69 336
rect 67 335 68 336
rect 66 335 67 336
rect 65 335 66 336
rect 64 335 65 336
rect 63 335 64 336
rect 62 335 63 336
rect 61 335 62 336
rect 60 335 61 336
rect 59 335 60 336
rect 58 335 59 336
rect 57 335 58 336
rect 56 335 57 336
rect 55 335 56 336
rect 54 335 55 336
rect 42 335 43 336
rect 41 335 42 336
rect 40 335 41 336
rect 39 335 40 336
rect 38 335 39 336
rect 37 335 38 336
rect 36 335 37 336
rect 35 335 36 336
rect 34 335 35 336
rect 33 335 34 336
rect 32 335 33 336
rect 31 335 32 336
rect 30 335 31 336
rect 441 336 442 337
rect 440 336 441 337
rect 439 336 440 337
rect 399 336 400 337
rect 398 336 399 337
rect 397 336 398 337
rect 176 336 177 337
rect 175 336 176 337
rect 174 336 175 337
rect 173 336 174 337
rect 172 336 173 337
rect 171 336 172 337
rect 170 336 171 337
rect 169 336 170 337
rect 168 336 169 337
rect 167 336 168 337
rect 166 336 167 337
rect 165 336 166 337
rect 164 336 165 337
rect 163 336 164 337
rect 162 336 163 337
rect 161 336 162 337
rect 160 336 161 337
rect 159 336 160 337
rect 158 336 159 337
rect 157 336 158 337
rect 156 336 157 337
rect 155 336 156 337
rect 154 336 155 337
rect 153 336 154 337
rect 152 336 153 337
rect 151 336 152 337
rect 150 336 151 337
rect 149 336 150 337
rect 148 336 149 337
rect 147 336 148 337
rect 146 336 147 337
rect 145 336 146 337
rect 144 336 145 337
rect 143 336 144 337
rect 142 336 143 337
rect 141 336 142 337
rect 140 336 141 337
rect 139 336 140 337
rect 138 336 139 337
rect 137 336 138 337
rect 136 336 137 337
rect 135 336 136 337
rect 134 336 135 337
rect 133 336 134 337
rect 132 336 133 337
rect 131 336 132 337
rect 130 336 131 337
rect 129 336 130 337
rect 128 336 129 337
rect 127 336 128 337
rect 126 336 127 337
rect 125 336 126 337
rect 124 336 125 337
rect 123 336 124 337
rect 122 336 123 337
rect 121 336 122 337
rect 120 336 121 337
rect 119 336 120 337
rect 118 336 119 337
rect 117 336 118 337
rect 116 336 117 337
rect 115 336 116 337
rect 114 336 115 337
rect 113 336 114 337
rect 112 336 113 337
rect 111 336 112 337
rect 110 336 111 337
rect 109 336 110 337
rect 89 336 90 337
rect 88 336 89 337
rect 87 336 88 337
rect 86 336 87 337
rect 85 336 86 337
rect 84 336 85 337
rect 83 336 84 337
rect 82 336 83 337
rect 81 336 82 337
rect 80 336 81 337
rect 79 336 80 337
rect 78 336 79 337
rect 77 336 78 337
rect 76 336 77 337
rect 75 336 76 337
rect 74 336 75 337
rect 73 336 74 337
rect 72 336 73 337
rect 71 336 72 337
rect 70 336 71 337
rect 69 336 70 337
rect 68 336 69 337
rect 67 336 68 337
rect 66 336 67 337
rect 65 336 66 337
rect 64 336 65 337
rect 63 336 64 337
rect 62 336 63 337
rect 61 336 62 337
rect 60 336 61 337
rect 59 336 60 337
rect 58 336 59 337
rect 57 336 58 337
rect 56 336 57 337
rect 55 336 56 337
rect 54 336 55 337
rect 42 336 43 337
rect 41 336 42 337
rect 40 336 41 337
rect 39 336 40 337
rect 38 336 39 337
rect 37 336 38 337
rect 36 336 37 337
rect 35 336 36 337
rect 34 336 35 337
rect 33 336 34 337
rect 32 336 33 337
rect 31 336 32 337
rect 441 337 442 338
rect 440 337 441 338
rect 439 337 440 338
rect 399 337 400 338
rect 398 337 399 338
rect 397 337 398 338
rect 180 337 181 338
rect 179 337 180 338
rect 178 337 179 338
rect 177 337 178 338
rect 176 337 177 338
rect 175 337 176 338
rect 174 337 175 338
rect 173 337 174 338
rect 172 337 173 338
rect 171 337 172 338
rect 170 337 171 338
rect 169 337 170 338
rect 168 337 169 338
rect 167 337 168 338
rect 166 337 167 338
rect 165 337 166 338
rect 164 337 165 338
rect 163 337 164 338
rect 162 337 163 338
rect 161 337 162 338
rect 160 337 161 338
rect 159 337 160 338
rect 158 337 159 338
rect 157 337 158 338
rect 156 337 157 338
rect 155 337 156 338
rect 154 337 155 338
rect 153 337 154 338
rect 152 337 153 338
rect 151 337 152 338
rect 150 337 151 338
rect 149 337 150 338
rect 148 337 149 338
rect 147 337 148 338
rect 146 337 147 338
rect 145 337 146 338
rect 144 337 145 338
rect 143 337 144 338
rect 142 337 143 338
rect 141 337 142 338
rect 140 337 141 338
rect 139 337 140 338
rect 138 337 139 338
rect 137 337 138 338
rect 136 337 137 338
rect 135 337 136 338
rect 134 337 135 338
rect 133 337 134 338
rect 132 337 133 338
rect 131 337 132 338
rect 130 337 131 338
rect 129 337 130 338
rect 128 337 129 338
rect 127 337 128 338
rect 126 337 127 338
rect 125 337 126 338
rect 124 337 125 338
rect 123 337 124 338
rect 122 337 123 338
rect 121 337 122 338
rect 120 337 121 338
rect 119 337 120 338
rect 118 337 119 338
rect 117 337 118 338
rect 116 337 117 338
rect 115 337 116 338
rect 114 337 115 338
rect 113 337 114 338
rect 112 337 113 338
rect 111 337 112 338
rect 110 337 111 338
rect 89 337 90 338
rect 88 337 89 338
rect 87 337 88 338
rect 86 337 87 338
rect 85 337 86 338
rect 84 337 85 338
rect 83 337 84 338
rect 82 337 83 338
rect 81 337 82 338
rect 80 337 81 338
rect 79 337 80 338
rect 78 337 79 338
rect 77 337 78 338
rect 76 337 77 338
rect 75 337 76 338
rect 74 337 75 338
rect 73 337 74 338
rect 72 337 73 338
rect 71 337 72 338
rect 70 337 71 338
rect 69 337 70 338
rect 68 337 69 338
rect 67 337 68 338
rect 66 337 67 338
rect 65 337 66 338
rect 64 337 65 338
rect 63 337 64 338
rect 62 337 63 338
rect 61 337 62 338
rect 60 337 61 338
rect 59 337 60 338
rect 58 337 59 338
rect 57 337 58 338
rect 56 337 57 338
rect 55 337 56 338
rect 42 337 43 338
rect 41 337 42 338
rect 40 337 41 338
rect 39 337 40 338
rect 38 337 39 338
rect 37 337 38 338
rect 36 337 37 338
rect 35 337 36 338
rect 34 337 35 338
rect 33 337 34 338
rect 32 337 33 338
rect 441 338 442 339
rect 440 338 441 339
rect 439 338 440 339
rect 438 338 439 339
rect 400 338 401 339
rect 399 338 400 339
rect 398 338 399 339
rect 397 338 398 339
rect 179 338 180 339
rect 178 338 179 339
rect 177 338 178 339
rect 176 338 177 339
rect 175 338 176 339
rect 174 338 175 339
rect 173 338 174 339
rect 172 338 173 339
rect 171 338 172 339
rect 170 338 171 339
rect 169 338 170 339
rect 168 338 169 339
rect 167 338 168 339
rect 166 338 167 339
rect 165 338 166 339
rect 164 338 165 339
rect 163 338 164 339
rect 162 338 163 339
rect 161 338 162 339
rect 160 338 161 339
rect 159 338 160 339
rect 158 338 159 339
rect 157 338 158 339
rect 156 338 157 339
rect 155 338 156 339
rect 154 338 155 339
rect 153 338 154 339
rect 152 338 153 339
rect 151 338 152 339
rect 150 338 151 339
rect 149 338 150 339
rect 148 338 149 339
rect 147 338 148 339
rect 146 338 147 339
rect 145 338 146 339
rect 144 338 145 339
rect 143 338 144 339
rect 142 338 143 339
rect 141 338 142 339
rect 140 338 141 339
rect 139 338 140 339
rect 138 338 139 339
rect 137 338 138 339
rect 136 338 137 339
rect 135 338 136 339
rect 134 338 135 339
rect 133 338 134 339
rect 132 338 133 339
rect 131 338 132 339
rect 130 338 131 339
rect 129 338 130 339
rect 128 338 129 339
rect 127 338 128 339
rect 126 338 127 339
rect 125 338 126 339
rect 124 338 125 339
rect 123 338 124 339
rect 122 338 123 339
rect 121 338 122 339
rect 120 338 121 339
rect 119 338 120 339
rect 118 338 119 339
rect 117 338 118 339
rect 116 338 117 339
rect 115 338 116 339
rect 114 338 115 339
rect 113 338 114 339
rect 112 338 113 339
rect 111 338 112 339
rect 90 338 91 339
rect 89 338 90 339
rect 88 338 89 339
rect 87 338 88 339
rect 86 338 87 339
rect 85 338 86 339
rect 84 338 85 339
rect 83 338 84 339
rect 82 338 83 339
rect 81 338 82 339
rect 80 338 81 339
rect 79 338 80 339
rect 78 338 79 339
rect 77 338 78 339
rect 76 338 77 339
rect 75 338 76 339
rect 74 338 75 339
rect 73 338 74 339
rect 72 338 73 339
rect 71 338 72 339
rect 70 338 71 339
rect 69 338 70 339
rect 68 338 69 339
rect 67 338 68 339
rect 66 338 67 339
rect 65 338 66 339
rect 64 338 65 339
rect 63 338 64 339
rect 62 338 63 339
rect 61 338 62 339
rect 60 338 61 339
rect 59 338 60 339
rect 58 338 59 339
rect 57 338 58 339
rect 56 338 57 339
rect 55 338 56 339
rect 43 338 44 339
rect 42 338 43 339
rect 41 338 42 339
rect 40 338 41 339
rect 39 338 40 339
rect 38 338 39 339
rect 37 338 38 339
rect 36 338 37 339
rect 35 338 36 339
rect 34 338 35 339
rect 33 338 34 339
rect 441 339 442 340
rect 440 339 441 340
rect 439 339 440 340
rect 438 339 439 340
rect 437 339 438 340
rect 436 339 437 340
rect 435 339 436 340
rect 434 339 435 340
rect 433 339 434 340
rect 432 339 433 340
rect 431 339 432 340
rect 430 339 431 340
rect 429 339 430 340
rect 428 339 429 340
rect 427 339 428 340
rect 426 339 427 340
rect 425 339 426 340
rect 424 339 425 340
rect 423 339 424 340
rect 422 339 423 340
rect 421 339 422 340
rect 420 339 421 340
rect 419 339 420 340
rect 418 339 419 340
rect 417 339 418 340
rect 416 339 417 340
rect 415 339 416 340
rect 414 339 415 340
rect 413 339 414 340
rect 412 339 413 340
rect 411 339 412 340
rect 410 339 411 340
rect 409 339 410 340
rect 408 339 409 340
rect 407 339 408 340
rect 406 339 407 340
rect 405 339 406 340
rect 404 339 405 340
rect 403 339 404 340
rect 402 339 403 340
rect 401 339 402 340
rect 400 339 401 340
rect 399 339 400 340
rect 398 339 399 340
rect 397 339 398 340
rect 178 339 179 340
rect 177 339 178 340
rect 176 339 177 340
rect 175 339 176 340
rect 174 339 175 340
rect 173 339 174 340
rect 172 339 173 340
rect 171 339 172 340
rect 170 339 171 340
rect 169 339 170 340
rect 168 339 169 340
rect 167 339 168 340
rect 166 339 167 340
rect 165 339 166 340
rect 164 339 165 340
rect 163 339 164 340
rect 162 339 163 340
rect 161 339 162 340
rect 160 339 161 340
rect 159 339 160 340
rect 158 339 159 340
rect 157 339 158 340
rect 156 339 157 340
rect 155 339 156 340
rect 154 339 155 340
rect 153 339 154 340
rect 152 339 153 340
rect 151 339 152 340
rect 150 339 151 340
rect 149 339 150 340
rect 148 339 149 340
rect 147 339 148 340
rect 146 339 147 340
rect 145 339 146 340
rect 144 339 145 340
rect 143 339 144 340
rect 142 339 143 340
rect 141 339 142 340
rect 140 339 141 340
rect 139 339 140 340
rect 138 339 139 340
rect 137 339 138 340
rect 136 339 137 340
rect 135 339 136 340
rect 134 339 135 340
rect 133 339 134 340
rect 132 339 133 340
rect 131 339 132 340
rect 130 339 131 340
rect 129 339 130 340
rect 128 339 129 340
rect 127 339 128 340
rect 126 339 127 340
rect 125 339 126 340
rect 124 339 125 340
rect 123 339 124 340
rect 122 339 123 340
rect 121 339 122 340
rect 120 339 121 340
rect 119 339 120 340
rect 118 339 119 340
rect 117 339 118 340
rect 116 339 117 340
rect 115 339 116 340
rect 114 339 115 340
rect 113 339 114 340
rect 112 339 113 340
rect 91 339 92 340
rect 90 339 91 340
rect 89 339 90 340
rect 88 339 89 340
rect 87 339 88 340
rect 86 339 87 340
rect 85 339 86 340
rect 84 339 85 340
rect 83 339 84 340
rect 82 339 83 340
rect 81 339 82 340
rect 80 339 81 340
rect 79 339 80 340
rect 78 339 79 340
rect 77 339 78 340
rect 76 339 77 340
rect 75 339 76 340
rect 74 339 75 340
rect 73 339 74 340
rect 72 339 73 340
rect 71 339 72 340
rect 70 339 71 340
rect 69 339 70 340
rect 68 339 69 340
rect 67 339 68 340
rect 66 339 67 340
rect 65 339 66 340
rect 64 339 65 340
rect 63 339 64 340
rect 62 339 63 340
rect 61 339 62 340
rect 60 339 61 340
rect 59 339 60 340
rect 58 339 59 340
rect 57 339 58 340
rect 56 339 57 340
rect 55 339 56 340
rect 43 339 44 340
rect 42 339 43 340
rect 41 339 42 340
rect 40 339 41 340
rect 39 339 40 340
rect 38 339 39 340
rect 37 339 38 340
rect 36 339 37 340
rect 35 339 36 340
rect 34 339 35 340
rect 441 340 442 341
rect 440 340 441 341
rect 439 340 440 341
rect 438 340 439 341
rect 437 340 438 341
rect 436 340 437 341
rect 435 340 436 341
rect 434 340 435 341
rect 433 340 434 341
rect 432 340 433 341
rect 431 340 432 341
rect 430 340 431 341
rect 429 340 430 341
rect 428 340 429 341
rect 427 340 428 341
rect 426 340 427 341
rect 425 340 426 341
rect 424 340 425 341
rect 423 340 424 341
rect 422 340 423 341
rect 421 340 422 341
rect 420 340 421 341
rect 419 340 420 341
rect 418 340 419 341
rect 417 340 418 341
rect 416 340 417 341
rect 415 340 416 341
rect 414 340 415 341
rect 413 340 414 341
rect 412 340 413 341
rect 411 340 412 341
rect 410 340 411 341
rect 409 340 410 341
rect 408 340 409 341
rect 407 340 408 341
rect 406 340 407 341
rect 405 340 406 341
rect 404 340 405 341
rect 403 340 404 341
rect 402 340 403 341
rect 401 340 402 341
rect 400 340 401 341
rect 399 340 400 341
rect 398 340 399 341
rect 397 340 398 341
rect 177 340 178 341
rect 176 340 177 341
rect 175 340 176 341
rect 174 340 175 341
rect 173 340 174 341
rect 172 340 173 341
rect 171 340 172 341
rect 170 340 171 341
rect 169 340 170 341
rect 168 340 169 341
rect 167 340 168 341
rect 166 340 167 341
rect 165 340 166 341
rect 164 340 165 341
rect 163 340 164 341
rect 162 340 163 341
rect 161 340 162 341
rect 160 340 161 341
rect 159 340 160 341
rect 158 340 159 341
rect 157 340 158 341
rect 156 340 157 341
rect 155 340 156 341
rect 154 340 155 341
rect 153 340 154 341
rect 152 340 153 341
rect 151 340 152 341
rect 150 340 151 341
rect 149 340 150 341
rect 148 340 149 341
rect 147 340 148 341
rect 146 340 147 341
rect 145 340 146 341
rect 144 340 145 341
rect 143 340 144 341
rect 142 340 143 341
rect 141 340 142 341
rect 140 340 141 341
rect 139 340 140 341
rect 138 340 139 341
rect 137 340 138 341
rect 136 340 137 341
rect 135 340 136 341
rect 134 340 135 341
rect 133 340 134 341
rect 132 340 133 341
rect 131 340 132 341
rect 130 340 131 341
rect 129 340 130 341
rect 128 340 129 341
rect 127 340 128 341
rect 126 340 127 341
rect 125 340 126 341
rect 124 340 125 341
rect 123 340 124 341
rect 122 340 123 341
rect 121 340 122 341
rect 120 340 121 341
rect 119 340 120 341
rect 118 340 119 341
rect 117 340 118 341
rect 116 340 117 341
rect 115 340 116 341
rect 114 340 115 341
rect 113 340 114 341
rect 92 340 93 341
rect 91 340 92 341
rect 90 340 91 341
rect 89 340 90 341
rect 88 340 89 341
rect 87 340 88 341
rect 86 340 87 341
rect 85 340 86 341
rect 84 340 85 341
rect 83 340 84 341
rect 82 340 83 341
rect 81 340 82 341
rect 80 340 81 341
rect 79 340 80 341
rect 78 340 79 341
rect 77 340 78 341
rect 76 340 77 341
rect 75 340 76 341
rect 74 340 75 341
rect 73 340 74 341
rect 72 340 73 341
rect 71 340 72 341
rect 70 340 71 341
rect 69 340 70 341
rect 68 340 69 341
rect 67 340 68 341
rect 66 340 67 341
rect 65 340 66 341
rect 64 340 65 341
rect 63 340 64 341
rect 62 340 63 341
rect 61 340 62 341
rect 60 340 61 341
rect 59 340 60 341
rect 58 340 59 341
rect 57 340 58 341
rect 56 340 57 341
rect 44 340 45 341
rect 43 340 44 341
rect 42 340 43 341
rect 41 340 42 341
rect 40 340 41 341
rect 39 340 40 341
rect 38 340 39 341
rect 37 340 38 341
rect 36 340 37 341
rect 35 340 36 341
rect 441 341 442 342
rect 440 341 441 342
rect 439 341 440 342
rect 438 341 439 342
rect 437 341 438 342
rect 436 341 437 342
rect 435 341 436 342
rect 434 341 435 342
rect 433 341 434 342
rect 432 341 433 342
rect 431 341 432 342
rect 430 341 431 342
rect 429 341 430 342
rect 428 341 429 342
rect 427 341 428 342
rect 426 341 427 342
rect 425 341 426 342
rect 424 341 425 342
rect 423 341 424 342
rect 422 341 423 342
rect 421 341 422 342
rect 420 341 421 342
rect 419 341 420 342
rect 418 341 419 342
rect 417 341 418 342
rect 416 341 417 342
rect 415 341 416 342
rect 414 341 415 342
rect 413 341 414 342
rect 412 341 413 342
rect 411 341 412 342
rect 410 341 411 342
rect 409 341 410 342
rect 408 341 409 342
rect 407 341 408 342
rect 406 341 407 342
rect 405 341 406 342
rect 404 341 405 342
rect 403 341 404 342
rect 402 341 403 342
rect 401 341 402 342
rect 400 341 401 342
rect 399 341 400 342
rect 398 341 399 342
rect 397 341 398 342
rect 176 341 177 342
rect 175 341 176 342
rect 174 341 175 342
rect 173 341 174 342
rect 172 341 173 342
rect 171 341 172 342
rect 170 341 171 342
rect 169 341 170 342
rect 168 341 169 342
rect 167 341 168 342
rect 166 341 167 342
rect 165 341 166 342
rect 164 341 165 342
rect 163 341 164 342
rect 162 341 163 342
rect 161 341 162 342
rect 160 341 161 342
rect 159 341 160 342
rect 158 341 159 342
rect 157 341 158 342
rect 156 341 157 342
rect 155 341 156 342
rect 154 341 155 342
rect 153 341 154 342
rect 152 341 153 342
rect 151 341 152 342
rect 150 341 151 342
rect 149 341 150 342
rect 148 341 149 342
rect 147 341 148 342
rect 146 341 147 342
rect 145 341 146 342
rect 144 341 145 342
rect 143 341 144 342
rect 142 341 143 342
rect 141 341 142 342
rect 140 341 141 342
rect 139 341 140 342
rect 138 341 139 342
rect 137 341 138 342
rect 136 341 137 342
rect 135 341 136 342
rect 134 341 135 342
rect 133 341 134 342
rect 132 341 133 342
rect 131 341 132 342
rect 130 341 131 342
rect 129 341 130 342
rect 128 341 129 342
rect 127 341 128 342
rect 126 341 127 342
rect 125 341 126 342
rect 124 341 125 342
rect 123 341 124 342
rect 122 341 123 342
rect 121 341 122 342
rect 120 341 121 342
rect 119 341 120 342
rect 118 341 119 342
rect 117 341 118 342
rect 116 341 117 342
rect 115 341 116 342
rect 114 341 115 342
rect 93 341 94 342
rect 92 341 93 342
rect 91 341 92 342
rect 90 341 91 342
rect 89 341 90 342
rect 88 341 89 342
rect 87 341 88 342
rect 86 341 87 342
rect 85 341 86 342
rect 84 341 85 342
rect 83 341 84 342
rect 82 341 83 342
rect 81 341 82 342
rect 80 341 81 342
rect 79 341 80 342
rect 78 341 79 342
rect 77 341 78 342
rect 76 341 77 342
rect 75 341 76 342
rect 74 341 75 342
rect 73 341 74 342
rect 72 341 73 342
rect 71 341 72 342
rect 70 341 71 342
rect 69 341 70 342
rect 68 341 69 342
rect 67 341 68 342
rect 66 341 67 342
rect 65 341 66 342
rect 64 341 65 342
rect 63 341 64 342
rect 62 341 63 342
rect 61 341 62 342
rect 60 341 61 342
rect 59 341 60 342
rect 58 341 59 342
rect 57 341 58 342
rect 56 341 57 342
rect 44 341 45 342
rect 43 341 44 342
rect 42 341 43 342
rect 41 341 42 342
rect 40 341 41 342
rect 39 341 40 342
rect 38 341 39 342
rect 37 341 38 342
rect 36 341 37 342
rect 441 342 442 343
rect 440 342 441 343
rect 439 342 440 343
rect 438 342 439 343
rect 437 342 438 343
rect 436 342 437 343
rect 435 342 436 343
rect 434 342 435 343
rect 433 342 434 343
rect 432 342 433 343
rect 431 342 432 343
rect 430 342 431 343
rect 429 342 430 343
rect 428 342 429 343
rect 427 342 428 343
rect 426 342 427 343
rect 425 342 426 343
rect 424 342 425 343
rect 423 342 424 343
rect 422 342 423 343
rect 421 342 422 343
rect 420 342 421 343
rect 419 342 420 343
rect 418 342 419 343
rect 417 342 418 343
rect 416 342 417 343
rect 415 342 416 343
rect 414 342 415 343
rect 413 342 414 343
rect 412 342 413 343
rect 411 342 412 343
rect 410 342 411 343
rect 409 342 410 343
rect 408 342 409 343
rect 407 342 408 343
rect 406 342 407 343
rect 405 342 406 343
rect 404 342 405 343
rect 403 342 404 343
rect 402 342 403 343
rect 401 342 402 343
rect 400 342 401 343
rect 399 342 400 343
rect 398 342 399 343
rect 397 342 398 343
rect 174 342 175 343
rect 173 342 174 343
rect 172 342 173 343
rect 171 342 172 343
rect 170 342 171 343
rect 169 342 170 343
rect 168 342 169 343
rect 167 342 168 343
rect 166 342 167 343
rect 165 342 166 343
rect 164 342 165 343
rect 163 342 164 343
rect 162 342 163 343
rect 161 342 162 343
rect 160 342 161 343
rect 159 342 160 343
rect 158 342 159 343
rect 157 342 158 343
rect 156 342 157 343
rect 155 342 156 343
rect 154 342 155 343
rect 153 342 154 343
rect 152 342 153 343
rect 151 342 152 343
rect 150 342 151 343
rect 149 342 150 343
rect 148 342 149 343
rect 147 342 148 343
rect 146 342 147 343
rect 145 342 146 343
rect 144 342 145 343
rect 143 342 144 343
rect 142 342 143 343
rect 141 342 142 343
rect 140 342 141 343
rect 139 342 140 343
rect 138 342 139 343
rect 137 342 138 343
rect 136 342 137 343
rect 135 342 136 343
rect 134 342 135 343
rect 133 342 134 343
rect 132 342 133 343
rect 131 342 132 343
rect 130 342 131 343
rect 129 342 130 343
rect 128 342 129 343
rect 127 342 128 343
rect 126 342 127 343
rect 125 342 126 343
rect 124 342 125 343
rect 123 342 124 343
rect 122 342 123 343
rect 121 342 122 343
rect 120 342 121 343
rect 119 342 120 343
rect 118 342 119 343
rect 117 342 118 343
rect 116 342 117 343
rect 115 342 116 343
rect 93 342 94 343
rect 92 342 93 343
rect 91 342 92 343
rect 90 342 91 343
rect 89 342 90 343
rect 88 342 89 343
rect 87 342 88 343
rect 86 342 87 343
rect 85 342 86 343
rect 84 342 85 343
rect 83 342 84 343
rect 82 342 83 343
rect 81 342 82 343
rect 80 342 81 343
rect 79 342 80 343
rect 78 342 79 343
rect 77 342 78 343
rect 76 342 77 343
rect 75 342 76 343
rect 74 342 75 343
rect 73 342 74 343
rect 72 342 73 343
rect 71 342 72 343
rect 70 342 71 343
rect 69 342 70 343
rect 68 342 69 343
rect 67 342 68 343
rect 66 342 67 343
rect 65 342 66 343
rect 64 342 65 343
rect 63 342 64 343
rect 62 342 63 343
rect 61 342 62 343
rect 60 342 61 343
rect 59 342 60 343
rect 58 342 59 343
rect 57 342 58 343
rect 45 342 46 343
rect 44 342 45 343
rect 43 342 44 343
rect 42 342 43 343
rect 41 342 42 343
rect 40 342 41 343
rect 39 342 40 343
rect 38 342 39 343
rect 37 342 38 343
rect 441 343 442 344
rect 440 343 441 344
rect 439 343 440 344
rect 438 343 439 344
rect 437 343 438 344
rect 436 343 437 344
rect 435 343 436 344
rect 434 343 435 344
rect 433 343 434 344
rect 432 343 433 344
rect 431 343 432 344
rect 430 343 431 344
rect 429 343 430 344
rect 428 343 429 344
rect 427 343 428 344
rect 426 343 427 344
rect 425 343 426 344
rect 424 343 425 344
rect 423 343 424 344
rect 422 343 423 344
rect 421 343 422 344
rect 420 343 421 344
rect 419 343 420 344
rect 418 343 419 344
rect 417 343 418 344
rect 416 343 417 344
rect 415 343 416 344
rect 414 343 415 344
rect 413 343 414 344
rect 412 343 413 344
rect 411 343 412 344
rect 410 343 411 344
rect 409 343 410 344
rect 408 343 409 344
rect 407 343 408 344
rect 406 343 407 344
rect 405 343 406 344
rect 404 343 405 344
rect 403 343 404 344
rect 402 343 403 344
rect 401 343 402 344
rect 400 343 401 344
rect 399 343 400 344
rect 398 343 399 344
rect 397 343 398 344
rect 172 343 173 344
rect 171 343 172 344
rect 170 343 171 344
rect 169 343 170 344
rect 168 343 169 344
rect 167 343 168 344
rect 166 343 167 344
rect 165 343 166 344
rect 164 343 165 344
rect 163 343 164 344
rect 162 343 163 344
rect 161 343 162 344
rect 160 343 161 344
rect 159 343 160 344
rect 158 343 159 344
rect 157 343 158 344
rect 156 343 157 344
rect 155 343 156 344
rect 154 343 155 344
rect 153 343 154 344
rect 152 343 153 344
rect 151 343 152 344
rect 150 343 151 344
rect 149 343 150 344
rect 148 343 149 344
rect 147 343 148 344
rect 146 343 147 344
rect 145 343 146 344
rect 144 343 145 344
rect 143 343 144 344
rect 142 343 143 344
rect 141 343 142 344
rect 140 343 141 344
rect 139 343 140 344
rect 138 343 139 344
rect 137 343 138 344
rect 136 343 137 344
rect 135 343 136 344
rect 134 343 135 344
rect 133 343 134 344
rect 132 343 133 344
rect 131 343 132 344
rect 130 343 131 344
rect 129 343 130 344
rect 128 343 129 344
rect 127 343 128 344
rect 126 343 127 344
rect 125 343 126 344
rect 124 343 125 344
rect 123 343 124 344
rect 122 343 123 344
rect 121 343 122 344
rect 120 343 121 344
rect 119 343 120 344
rect 118 343 119 344
rect 117 343 118 344
rect 116 343 117 344
rect 94 343 95 344
rect 93 343 94 344
rect 92 343 93 344
rect 91 343 92 344
rect 90 343 91 344
rect 89 343 90 344
rect 88 343 89 344
rect 87 343 88 344
rect 86 343 87 344
rect 85 343 86 344
rect 84 343 85 344
rect 83 343 84 344
rect 82 343 83 344
rect 81 343 82 344
rect 80 343 81 344
rect 79 343 80 344
rect 78 343 79 344
rect 77 343 78 344
rect 76 343 77 344
rect 75 343 76 344
rect 74 343 75 344
rect 73 343 74 344
rect 72 343 73 344
rect 71 343 72 344
rect 70 343 71 344
rect 69 343 70 344
rect 68 343 69 344
rect 67 343 68 344
rect 66 343 67 344
rect 65 343 66 344
rect 64 343 65 344
rect 63 343 64 344
rect 62 343 63 344
rect 61 343 62 344
rect 60 343 61 344
rect 59 343 60 344
rect 58 343 59 344
rect 57 343 58 344
rect 45 343 46 344
rect 44 343 45 344
rect 43 343 44 344
rect 42 343 43 344
rect 41 343 42 344
rect 40 343 41 344
rect 39 343 40 344
rect 441 344 442 345
rect 440 344 441 345
rect 439 344 440 345
rect 438 344 439 345
rect 437 344 438 345
rect 436 344 437 345
rect 435 344 436 345
rect 434 344 435 345
rect 433 344 434 345
rect 432 344 433 345
rect 431 344 432 345
rect 430 344 431 345
rect 429 344 430 345
rect 428 344 429 345
rect 427 344 428 345
rect 426 344 427 345
rect 425 344 426 345
rect 424 344 425 345
rect 423 344 424 345
rect 422 344 423 345
rect 421 344 422 345
rect 420 344 421 345
rect 419 344 420 345
rect 418 344 419 345
rect 417 344 418 345
rect 416 344 417 345
rect 415 344 416 345
rect 414 344 415 345
rect 413 344 414 345
rect 412 344 413 345
rect 411 344 412 345
rect 410 344 411 345
rect 409 344 410 345
rect 408 344 409 345
rect 407 344 408 345
rect 406 344 407 345
rect 405 344 406 345
rect 404 344 405 345
rect 403 344 404 345
rect 402 344 403 345
rect 401 344 402 345
rect 400 344 401 345
rect 399 344 400 345
rect 398 344 399 345
rect 397 344 398 345
rect 170 344 171 345
rect 169 344 170 345
rect 168 344 169 345
rect 167 344 168 345
rect 166 344 167 345
rect 165 344 166 345
rect 164 344 165 345
rect 163 344 164 345
rect 162 344 163 345
rect 161 344 162 345
rect 160 344 161 345
rect 159 344 160 345
rect 158 344 159 345
rect 157 344 158 345
rect 156 344 157 345
rect 155 344 156 345
rect 154 344 155 345
rect 153 344 154 345
rect 152 344 153 345
rect 151 344 152 345
rect 150 344 151 345
rect 149 344 150 345
rect 148 344 149 345
rect 147 344 148 345
rect 146 344 147 345
rect 145 344 146 345
rect 144 344 145 345
rect 143 344 144 345
rect 142 344 143 345
rect 141 344 142 345
rect 140 344 141 345
rect 139 344 140 345
rect 138 344 139 345
rect 137 344 138 345
rect 136 344 137 345
rect 135 344 136 345
rect 134 344 135 345
rect 133 344 134 345
rect 132 344 133 345
rect 131 344 132 345
rect 130 344 131 345
rect 129 344 130 345
rect 128 344 129 345
rect 127 344 128 345
rect 126 344 127 345
rect 125 344 126 345
rect 124 344 125 345
rect 123 344 124 345
rect 122 344 123 345
rect 121 344 122 345
rect 120 344 121 345
rect 119 344 120 345
rect 118 344 119 345
rect 117 344 118 345
rect 95 344 96 345
rect 94 344 95 345
rect 93 344 94 345
rect 92 344 93 345
rect 91 344 92 345
rect 90 344 91 345
rect 89 344 90 345
rect 88 344 89 345
rect 87 344 88 345
rect 86 344 87 345
rect 85 344 86 345
rect 84 344 85 345
rect 83 344 84 345
rect 82 344 83 345
rect 81 344 82 345
rect 80 344 81 345
rect 79 344 80 345
rect 78 344 79 345
rect 77 344 78 345
rect 76 344 77 345
rect 75 344 76 345
rect 74 344 75 345
rect 73 344 74 345
rect 72 344 73 345
rect 71 344 72 345
rect 70 344 71 345
rect 69 344 70 345
rect 68 344 69 345
rect 67 344 68 345
rect 66 344 67 345
rect 65 344 66 345
rect 64 344 65 345
rect 63 344 64 345
rect 62 344 63 345
rect 61 344 62 345
rect 60 344 61 345
rect 59 344 60 345
rect 58 344 59 345
rect 57 344 58 345
rect 46 344 47 345
rect 45 344 46 345
rect 44 344 45 345
rect 43 344 44 345
rect 42 344 43 345
rect 41 344 42 345
rect 40 344 41 345
rect 441 345 442 346
rect 440 345 441 346
rect 439 345 440 346
rect 438 345 439 346
rect 437 345 438 346
rect 436 345 437 346
rect 435 345 436 346
rect 434 345 435 346
rect 433 345 434 346
rect 432 345 433 346
rect 431 345 432 346
rect 430 345 431 346
rect 429 345 430 346
rect 428 345 429 346
rect 427 345 428 346
rect 426 345 427 346
rect 425 345 426 346
rect 424 345 425 346
rect 423 345 424 346
rect 422 345 423 346
rect 421 345 422 346
rect 420 345 421 346
rect 419 345 420 346
rect 418 345 419 346
rect 417 345 418 346
rect 416 345 417 346
rect 415 345 416 346
rect 414 345 415 346
rect 413 345 414 346
rect 412 345 413 346
rect 411 345 412 346
rect 410 345 411 346
rect 409 345 410 346
rect 408 345 409 346
rect 407 345 408 346
rect 406 345 407 346
rect 405 345 406 346
rect 404 345 405 346
rect 403 345 404 346
rect 402 345 403 346
rect 401 345 402 346
rect 400 345 401 346
rect 399 345 400 346
rect 398 345 399 346
rect 397 345 398 346
rect 168 345 169 346
rect 167 345 168 346
rect 166 345 167 346
rect 165 345 166 346
rect 164 345 165 346
rect 163 345 164 346
rect 162 345 163 346
rect 161 345 162 346
rect 160 345 161 346
rect 159 345 160 346
rect 158 345 159 346
rect 157 345 158 346
rect 156 345 157 346
rect 155 345 156 346
rect 154 345 155 346
rect 153 345 154 346
rect 152 345 153 346
rect 151 345 152 346
rect 150 345 151 346
rect 149 345 150 346
rect 148 345 149 346
rect 147 345 148 346
rect 146 345 147 346
rect 145 345 146 346
rect 144 345 145 346
rect 143 345 144 346
rect 142 345 143 346
rect 141 345 142 346
rect 140 345 141 346
rect 139 345 140 346
rect 138 345 139 346
rect 137 345 138 346
rect 136 345 137 346
rect 135 345 136 346
rect 134 345 135 346
rect 133 345 134 346
rect 132 345 133 346
rect 131 345 132 346
rect 130 345 131 346
rect 129 345 130 346
rect 128 345 129 346
rect 127 345 128 346
rect 126 345 127 346
rect 125 345 126 346
rect 124 345 125 346
rect 123 345 124 346
rect 122 345 123 346
rect 121 345 122 346
rect 120 345 121 346
rect 119 345 120 346
rect 96 345 97 346
rect 95 345 96 346
rect 94 345 95 346
rect 93 345 94 346
rect 92 345 93 346
rect 91 345 92 346
rect 90 345 91 346
rect 89 345 90 346
rect 88 345 89 346
rect 87 345 88 346
rect 86 345 87 346
rect 85 345 86 346
rect 84 345 85 346
rect 83 345 84 346
rect 82 345 83 346
rect 81 345 82 346
rect 80 345 81 346
rect 79 345 80 346
rect 78 345 79 346
rect 77 345 78 346
rect 76 345 77 346
rect 75 345 76 346
rect 74 345 75 346
rect 73 345 74 346
rect 72 345 73 346
rect 71 345 72 346
rect 70 345 71 346
rect 69 345 70 346
rect 68 345 69 346
rect 67 345 68 346
rect 66 345 67 346
rect 65 345 66 346
rect 64 345 65 346
rect 63 345 64 346
rect 62 345 63 346
rect 61 345 62 346
rect 60 345 61 346
rect 59 345 60 346
rect 58 345 59 346
rect 46 345 47 346
rect 45 345 46 346
rect 44 345 45 346
rect 43 345 44 346
rect 42 345 43 346
rect 441 346 442 347
rect 440 346 441 347
rect 439 346 440 347
rect 438 346 439 347
rect 437 346 438 347
rect 436 346 437 347
rect 435 346 436 347
rect 434 346 435 347
rect 433 346 434 347
rect 432 346 433 347
rect 431 346 432 347
rect 430 346 431 347
rect 429 346 430 347
rect 428 346 429 347
rect 427 346 428 347
rect 426 346 427 347
rect 425 346 426 347
rect 424 346 425 347
rect 423 346 424 347
rect 422 346 423 347
rect 421 346 422 347
rect 420 346 421 347
rect 419 346 420 347
rect 418 346 419 347
rect 417 346 418 347
rect 416 346 417 347
rect 415 346 416 347
rect 414 346 415 347
rect 413 346 414 347
rect 412 346 413 347
rect 411 346 412 347
rect 410 346 411 347
rect 409 346 410 347
rect 408 346 409 347
rect 407 346 408 347
rect 406 346 407 347
rect 405 346 406 347
rect 404 346 405 347
rect 403 346 404 347
rect 402 346 403 347
rect 401 346 402 347
rect 400 346 401 347
rect 399 346 400 347
rect 398 346 399 347
rect 397 346 398 347
rect 165 346 166 347
rect 164 346 165 347
rect 163 346 164 347
rect 162 346 163 347
rect 161 346 162 347
rect 160 346 161 347
rect 159 346 160 347
rect 158 346 159 347
rect 157 346 158 347
rect 156 346 157 347
rect 155 346 156 347
rect 154 346 155 347
rect 153 346 154 347
rect 152 346 153 347
rect 151 346 152 347
rect 150 346 151 347
rect 149 346 150 347
rect 148 346 149 347
rect 147 346 148 347
rect 146 346 147 347
rect 145 346 146 347
rect 144 346 145 347
rect 143 346 144 347
rect 142 346 143 347
rect 141 346 142 347
rect 140 346 141 347
rect 139 346 140 347
rect 138 346 139 347
rect 137 346 138 347
rect 136 346 137 347
rect 135 346 136 347
rect 134 346 135 347
rect 133 346 134 347
rect 132 346 133 347
rect 131 346 132 347
rect 130 346 131 347
rect 129 346 130 347
rect 128 346 129 347
rect 127 346 128 347
rect 126 346 127 347
rect 125 346 126 347
rect 124 346 125 347
rect 123 346 124 347
rect 122 346 123 347
rect 121 346 122 347
rect 120 346 121 347
rect 97 346 98 347
rect 96 346 97 347
rect 95 346 96 347
rect 94 346 95 347
rect 93 346 94 347
rect 92 346 93 347
rect 91 346 92 347
rect 90 346 91 347
rect 89 346 90 347
rect 88 346 89 347
rect 87 346 88 347
rect 86 346 87 347
rect 85 346 86 347
rect 84 346 85 347
rect 83 346 84 347
rect 82 346 83 347
rect 81 346 82 347
rect 80 346 81 347
rect 79 346 80 347
rect 78 346 79 347
rect 77 346 78 347
rect 76 346 77 347
rect 75 346 76 347
rect 74 346 75 347
rect 73 346 74 347
rect 72 346 73 347
rect 71 346 72 347
rect 70 346 71 347
rect 69 346 70 347
rect 68 346 69 347
rect 67 346 68 347
rect 66 346 67 347
rect 65 346 66 347
rect 64 346 65 347
rect 63 346 64 347
rect 62 346 63 347
rect 61 346 62 347
rect 60 346 61 347
rect 59 346 60 347
rect 58 346 59 347
rect 47 346 48 347
rect 46 346 47 347
rect 45 346 46 347
rect 441 347 442 348
rect 440 347 441 348
rect 439 347 440 348
rect 438 347 439 348
rect 437 347 438 348
rect 436 347 437 348
rect 435 347 436 348
rect 434 347 435 348
rect 433 347 434 348
rect 432 347 433 348
rect 431 347 432 348
rect 430 347 431 348
rect 429 347 430 348
rect 428 347 429 348
rect 427 347 428 348
rect 426 347 427 348
rect 425 347 426 348
rect 424 347 425 348
rect 423 347 424 348
rect 422 347 423 348
rect 421 347 422 348
rect 420 347 421 348
rect 419 347 420 348
rect 418 347 419 348
rect 417 347 418 348
rect 416 347 417 348
rect 415 347 416 348
rect 414 347 415 348
rect 413 347 414 348
rect 412 347 413 348
rect 411 347 412 348
rect 410 347 411 348
rect 409 347 410 348
rect 408 347 409 348
rect 407 347 408 348
rect 406 347 407 348
rect 405 347 406 348
rect 404 347 405 348
rect 403 347 404 348
rect 402 347 403 348
rect 401 347 402 348
rect 400 347 401 348
rect 399 347 400 348
rect 398 347 399 348
rect 397 347 398 348
rect 162 347 163 348
rect 161 347 162 348
rect 160 347 161 348
rect 159 347 160 348
rect 158 347 159 348
rect 157 347 158 348
rect 156 347 157 348
rect 155 347 156 348
rect 154 347 155 348
rect 153 347 154 348
rect 152 347 153 348
rect 151 347 152 348
rect 150 347 151 348
rect 149 347 150 348
rect 148 347 149 348
rect 147 347 148 348
rect 146 347 147 348
rect 145 347 146 348
rect 144 347 145 348
rect 143 347 144 348
rect 142 347 143 348
rect 141 347 142 348
rect 140 347 141 348
rect 139 347 140 348
rect 138 347 139 348
rect 137 347 138 348
rect 136 347 137 348
rect 135 347 136 348
rect 134 347 135 348
rect 133 347 134 348
rect 132 347 133 348
rect 131 347 132 348
rect 130 347 131 348
rect 129 347 130 348
rect 128 347 129 348
rect 127 347 128 348
rect 126 347 127 348
rect 125 347 126 348
rect 124 347 125 348
rect 123 347 124 348
rect 98 347 99 348
rect 97 347 98 348
rect 96 347 97 348
rect 95 347 96 348
rect 94 347 95 348
rect 93 347 94 348
rect 92 347 93 348
rect 91 347 92 348
rect 90 347 91 348
rect 89 347 90 348
rect 88 347 89 348
rect 87 347 88 348
rect 86 347 87 348
rect 85 347 86 348
rect 84 347 85 348
rect 83 347 84 348
rect 82 347 83 348
rect 81 347 82 348
rect 80 347 81 348
rect 79 347 80 348
rect 78 347 79 348
rect 77 347 78 348
rect 76 347 77 348
rect 75 347 76 348
rect 74 347 75 348
rect 73 347 74 348
rect 72 347 73 348
rect 71 347 72 348
rect 70 347 71 348
rect 69 347 70 348
rect 68 347 69 348
rect 67 347 68 348
rect 66 347 67 348
rect 65 347 66 348
rect 64 347 65 348
rect 63 347 64 348
rect 62 347 63 348
rect 61 347 62 348
rect 60 347 61 348
rect 59 347 60 348
rect 441 348 442 349
rect 440 348 441 349
rect 439 348 440 349
rect 438 348 439 349
rect 437 348 438 349
rect 436 348 437 349
rect 435 348 436 349
rect 434 348 435 349
rect 433 348 434 349
rect 432 348 433 349
rect 431 348 432 349
rect 430 348 431 349
rect 429 348 430 349
rect 428 348 429 349
rect 427 348 428 349
rect 426 348 427 349
rect 425 348 426 349
rect 424 348 425 349
rect 423 348 424 349
rect 422 348 423 349
rect 421 348 422 349
rect 420 348 421 349
rect 419 348 420 349
rect 418 348 419 349
rect 417 348 418 349
rect 416 348 417 349
rect 415 348 416 349
rect 414 348 415 349
rect 413 348 414 349
rect 412 348 413 349
rect 411 348 412 349
rect 410 348 411 349
rect 409 348 410 349
rect 408 348 409 349
rect 407 348 408 349
rect 406 348 407 349
rect 405 348 406 349
rect 404 348 405 349
rect 403 348 404 349
rect 402 348 403 349
rect 401 348 402 349
rect 400 348 401 349
rect 399 348 400 349
rect 398 348 399 349
rect 397 348 398 349
rect 158 348 159 349
rect 157 348 158 349
rect 156 348 157 349
rect 155 348 156 349
rect 154 348 155 349
rect 153 348 154 349
rect 152 348 153 349
rect 151 348 152 349
rect 150 348 151 349
rect 149 348 150 349
rect 148 348 149 349
rect 147 348 148 349
rect 146 348 147 349
rect 145 348 146 349
rect 144 348 145 349
rect 143 348 144 349
rect 142 348 143 349
rect 141 348 142 349
rect 140 348 141 349
rect 139 348 140 349
rect 138 348 139 349
rect 137 348 138 349
rect 136 348 137 349
rect 135 348 136 349
rect 134 348 135 349
rect 133 348 134 349
rect 132 348 133 349
rect 131 348 132 349
rect 130 348 131 349
rect 129 348 130 349
rect 128 348 129 349
rect 127 348 128 349
rect 126 348 127 349
rect 99 348 100 349
rect 98 348 99 349
rect 97 348 98 349
rect 96 348 97 349
rect 95 348 96 349
rect 94 348 95 349
rect 93 348 94 349
rect 92 348 93 349
rect 91 348 92 349
rect 90 348 91 349
rect 89 348 90 349
rect 88 348 89 349
rect 87 348 88 349
rect 86 348 87 349
rect 85 348 86 349
rect 84 348 85 349
rect 83 348 84 349
rect 82 348 83 349
rect 81 348 82 349
rect 80 348 81 349
rect 79 348 80 349
rect 78 348 79 349
rect 77 348 78 349
rect 76 348 77 349
rect 75 348 76 349
rect 74 348 75 349
rect 73 348 74 349
rect 72 348 73 349
rect 71 348 72 349
rect 70 348 71 349
rect 69 348 70 349
rect 68 348 69 349
rect 67 348 68 349
rect 66 348 67 349
rect 65 348 66 349
rect 64 348 65 349
rect 63 348 64 349
rect 62 348 63 349
rect 61 348 62 349
rect 60 348 61 349
rect 59 348 60 349
rect 441 349 442 350
rect 440 349 441 350
rect 439 349 440 350
rect 438 349 439 350
rect 420 349 421 350
rect 419 349 420 350
rect 418 349 419 350
rect 417 349 418 350
rect 399 349 400 350
rect 398 349 399 350
rect 397 349 398 350
rect 152 349 153 350
rect 151 349 152 350
rect 150 349 151 350
rect 149 349 150 350
rect 148 349 149 350
rect 147 349 148 350
rect 146 349 147 350
rect 145 349 146 350
rect 144 349 145 350
rect 143 349 144 350
rect 142 349 143 350
rect 141 349 142 350
rect 140 349 141 350
rect 139 349 140 350
rect 138 349 139 350
rect 137 349 138 350
rect 136 349 137 350
rect 135 349 136 350
rect 134 349 135 350
rect 133 349 134 350
rect 132 349 133 350
rect 131 349 132 350
rect 100 349 101 350
rect 99 349 100 350
rect 98 349 99 350
rect 97 349 98 350
rect 96 349 97 350
rect 95 349 96 350
rect 94 349 95 350
rect 93 349 94 350
rect 92 349 93 350
rect 91 349 92 350
rect 90 349 91 350
rect 89 349 90 350
rect 88 349 89 350
rect 87 349 88 350
rect 86 349 87 350
rect 85 349 86 350
rect 84 349 85 350
rect 83 349 84 350
rect 82 349 83 350
rect 81 349 82 350
rect 80 349 81 350
rect 79 349 80 350
rect 78 349 79 350
rect 77 349 78 350
rect 76 349 77 350
rect 75 349 76 350
rect 74 349 75 350
rect 73 349 74 350
rect 72 349 73 350
rect 71 349 72 350
rect 70 349 71 350
rect 69 349 70 350
rect 68 349 69 350
rect 67 349 68 350
rect 66 349 67 350
rect 65 349 66 350
rect 64 349 65 350
rect 63 349 64 350
rect 62 349 63 350
rect 61 349 62 350
rect 60 349 61 350
rect 441 350 442 351
rect 440 350 441 351
rect 439 350 440 351
rect 438 350 439 351
rect 420 350 421 351
rect 419 350 420 351
rect 418 350 419 351
rect 417 350 418 351
rect 399 350 400 351
rect 398 350 399 351
rect 397 350 398 351
rect 101 350 102 351
rect 100 350 101 351
rect 99 350 100 351
rect 98 350 99 351
rect 97 350 98 351
rect 96 350 97 351
rect 95 350 96 351
rect 94 350 95 351
rect 93 350 94 351
rect 92 350 93 351
rect 91 350 92 351
rect 90 350 91 351
rect 89 350 90 351
rect 88 350 89 351
rect 87 350 88 351
rect 86 350 87 351
rect 85 350 86 351
rect 84 350 85 351
rect 83 350 84 351
rect 82 350 83 351
rect 81 350 82 351
rect 80 350 81 351
rect 79 350 80 351
rect 78 350 79 351
rect 77 350 78 351
rect 76 350 77 351
rect 75 350 76 351
rect 74 350 75 351
rect 73 350 74 351
rect 72 350 73 351
rect 71 350 72 351
rect 70 350 71 351
rect 69 350 70 351
rect 68 350 69 351
rect 67 350 68 351
rect 66 350 67 351
rect 65 350 66 351
rect 64 350 65 351
rect 63 350 64 351
rect 62 350 63 351
rect 61 350 62 351
rect 60 350 61 351
rect 441 351 442 352
rect 440 351 441 352
rect 439 351 440 352
rect 420 351 421 352
rect 419 351 420 352
rect 418 351 419 352
rect 417 351 418 352
rect 399 351 400 352
rect 398 351 399 352
rect 397 351 398 352
rect 102 351 103 352
rect 101 351 102 352
rect 100 351 101 352
rect 99 351 100 352
rect 98 351 99 352
rect 97 351 98 352
rect 96 351 97 352
rect 95 351 96 352
rect 94 351 95 352
rect 93 351 94 352
rect 92 351 93 352
rect 91 351 92 352
rect 90 351 91 352
rect 89 351 90 352
rect 88 351 89 352
rect 87 351 88 352
rect 86 351 87 352
rect 85 351 86 352
rect 84 351 85 352
rect 83 351 84 352
rect 82 351 83 352
rect 81 351 82 352
rect 80 351 81 352
rect 79 351 80 352
rect 78 351 79 352
rect 77 351 78 352
rect 76 351 77 352
rect 75 351 76 352
rect 74 351 75 352
rect 73 351 74 352
rect 72 351 73 352
rect 71 351 72 352
rect 70 351 71 352
rect 69 351 70 352
rect 68 351 69 352
rect 67 351 68 352
rect 66 351 67 352
rect 65 351 66 352
rect 64 351 65 352
rect 63 351 64 352
rect 62 351 63 352
rect 61 351 62 352
rect 60 351 61 352
rect 441 352 442 353
rect 440 352 441 353
rect 439 352 440 353
rect 420 352 421 353
rect 419 352 420 353
rect 418 352 419 353
rect 417 352 418 353
rect 399 352 400 353
rect 398 352 399 353
rect 397 352 398 353
rect 103 352 104 353
rect 102 352 103 353
rect 101 352 102 353
rect 100 352 101 353
rect 99 352 100 353
rect 98 352 99 353
rect 97 352 98 353
rect 96 352 97 353
rect 95 352 96 353
rect 94 352 95 353
rect 93 352 94 353
rect 92 352 93 353
rect 91 352 92 353
rect 90 352 91 353
rect 89 352 90 353
rect 88 352 89 353
rect 87 352 88 353
rect 86 352 87 353
rect 85 352 86 353
rect 84 352 85 353
rect 83 352 84 353
rect 82 352 83 353
rect 81 352 82 353
rect 80 352 81 353
rect 79 352 80 353
rect 78 352 79 353
rect 77 352 78 353
rect 76 352 77 353
rect 75 352 76 353
rect 74 352 75 353
rect 73 352 74 353
rect 72 352 73 353
rect 71 352 72 353
rect 70 352 71 353
rect 69 352 70 353
rect 68 352 69 353
rect 67 352 68 353
rect 66 352 67 353
rect 65 352 66 353
rect 64 352 65 353
rect 63 352 64 353
rect 62 352 63 353
rect 61 352 62 353
rect 441 353 442 354
rect 440 353 441 354
rect 439 353 440 354
rect 420 353 421 354
rect 419 353 420 354
rect 418 353 419 354
rect 417 353 418 354
rect 399 353 400 354
rect 398 353 399 354
rect 397 353 398 354
rect 105 353 106 354
rect 104 353 105 354
rect 103 353 104 354
rect 102 353 103 354
rect 101 353 102 354
rect 100 353 101 354
rect 99 353 100 354
rect 98 353 99 354
rect 97 353 98 354
rect 96 353 97 354
rect 95 353 96 354
rect 94 353 95 354
rect 93 353 94 354
rect 92 353 93 354
rect 91 353 92 354
rect 90 353 91 354
rect 89 353 90 354
rect 88 353 89 354
rect 87 353 88 354
rect 86 353 87 354
rect 85 353 86 354
rect 84 353 85 354
rect 83 353 84 354
rect 82 353 83 354
rect 81 353 82 354
rect 80 353 81 354
rect 79 353 80 354
rect 78 353 79 354
rect 77 353 78 354
rect 76 353 77 354
rect 75 353 76 354
rect 74 353 75 354
rect 73 353 74 354
rect 72 353 73 354
rect 71 353 72 354
rect 70 353 71 354
rect 69 353 70 354
rect 68 353 69 354
rect 67 353 68 354
rect 66 353 67 354
rect 65 353 66 354
rect 64 353 65 354
rect 63 353 64 354
rect 62 353 63 354
rect 441 354 442 355
rect 440 354 441 355
rect 439 354 440 355
rect 420 354 421 355
rect 419 354 420 355
rect 418 354 419 355
rect 417 354 418 355
rect 399 354 400 355
rect 398 354 399 355
rect 397 354 398 355
rect 106 354 107 355
rect 105 354 106 355
rect 104 354 105 355
rect 103 354 104 355
rect 102 354 103 355
rect 101 354 102 355
rect 100 354 101 355
rect 99 354 100 355
rect 98 354 99 355
rect 97 354 98 355
rect 96 354 97 355
rect 95 354 96 355
rect 94 354 95 355
rect 93 354 94 355
rect 92 354 93 355
rect 91 354 92 355
rect 90 354 91 355
rect 89 354 90 355
rect 88 354 89 355
rect 87 354 88 355
rect 86 354 87 355
rect 85 354 86 355
rect 84 354 85 355
rect 83 354 84 355
rect 82 354 83 355
rect 81 354 82 355
rect 80 354 81 355
rect 79 354 80 355
rect 78 354 79 355
rect 77 354 78 355
rect 76 354 77 355
rect 75 354 76 355
rect 74 354 75 355
rect 73 354 74 355
rect 72 354 73 355
rect 71 354 72 355
rect 70 354 71 355
rect 69 354 70 355
rect 68 354 69 355
rect 67 354 68 355
rect 66 354 67 355
rect 65 354 66 355
rect 64 354 65 355
rect 63 354 64 355
rect 441 355 442 356
rect 440 355 441 356
rect 439 355 440 356
rect 420 355 421 356
rect 419 355 420 356
rect 418 355 419 356
rect 417 355 418 356
rect 399 355 400 356
rect 398 355 399 356
rect 397 355 398 356
rect 107 355 108 356
rect 106 355 107 356
rect 105 355 106 356
rect 104 355 105 356
rect 103 355 104 356
rect 102 355 103 356
rect 101 355 102 356
rect 100 355 101 356
rect 99 355 100 356
rect 98 355 99 356
rect 97 355 98 356
rect 96 355 97 356
rect 95 355 96 356
rect 94 355 95 356
rect 93 355 94 356
rect 92 355 93 356
rect 91 355 92 356
rect 90 355 91 356
rect 89 355 90 356
rect 88 355 89 356
rect 87 355 88 356
rect 86 355 87 356
rect 85 355 86 356
rect 84 355 85 356
rect 83 355 84 356
rect 82 355 83 356
rect 81 355 82 356
rect 80 355 81 356
rect 79 355 80 356
rect 78 355 79 356
rect 77 355 78 356
rect 76 355 77 356
rect 75 355 76 356
rect 74 355 75 356
rect 73 355 74 356
rect 72 355 73 356
rect 71 355 72 356
rect 70 355 71 356
rect 69 355 70 356
rect 68 355 69 356
rect 67 355 68 356
rect 66 355 67 356
rect 65 355 66 356
rect 64 355 65 356
rect 63 355 64 356
rect 441 356 442 357
rect 440 356 441 357
rect 439 356 440 357
rect 420 356 421 357
rect 419 356 420 357
rect 418 356 419 357
rect 417 356 418 357
rect 399 356 400 357
rect 398 356 399 357
rect 397 356 398 357
rect 109 356 110 357
rect 108 356 109 357
rect 107 356 108 357
rect 106 356 107 357
rect 105 356 106 357
rect 104 356 105 357
rect 103 356 104 357
rect 102 356 103 357
rect 101 356 102 357
rect 100 356 101 357
rect 99 356 100 357
rect 98 356 99 357
rect 97 356 98 357
rect 96 356 97 357
rect 95 356 96 357
rect 94 356 95 357
rect 93 356 94 357
rect 92 356 93 357
rect 91 356 92 357
rect 90 356 91 357
rect 89 356 90 357
rect 88 356 89 357
rect 87 356 88 357
rect 86 356 87 357
rect 85 356 86 357
rect 84 356 85 357
rect 83 356 84 357
rect 82 356 83 357
rect 81 356 82 357
rect 80 356 81 357
rect 79 356 80 357
rect 78 356 79 357
rect 77 356 78 357
rect 76 356 77 357
rect 75 356 76 357
rect 74 356 75 357
rect 73 356 74 357
rect 72 356 73 357
rect 71 356 72 357
rect 70 356 71 357
rect 69 356 70 357
rect 68 356 69 357
rect 67 356 68 357
rect 66 356 67 357
rect 65 356 66 357
rect 441 357 442 358
rect 440 357 441 358
rect 439 357 440 358
rect 420 357 421 358
rect 419 357 420 358
rect 418 357 419 358
rect 417 357 418 358
rect 399 357 400 358
rect 398 357 399 358
rect 397 357 398 358
rect 110 357 111 358
rect 109 357 110 358
rect 108 357 109 358
rect 107 357 108 358
rect 106 357 107 358
rect 105 357 106 358
rect 104 357 105 358
rect 103 357 104 358
rect 102 357 103 358
rect 101 357 102 358
rect 100 357 101 358
rect 99 357 100 358
rect 98 357 99 358
rect 97 357 98 358
rect 96 357 97 358
rect 95 357 96 358
rect 94 357 95 358
rect 93 357 94 358
rect 92 357 93 358
rect 91 357 92 358
rect 90 357 91 358
rect 89 357 90 358
rect 88 357 89 358
rect 87 357 88 358
rect 86 357 87 358
rect 85 357 86 358
rect 84 357 85 358
rect 83 357 84 358
rect 82 357 83 358
rect 81 357 82 358
rect 80 357 81 358
rect 79 357 80 358
rect 78 357 79 358
rect 77 357 78 358
rect 76 357 77 358
rect 75 357 76 358
rect 74 357 75 358
rect 73 357 74 358
rect 72 357 73 358
rect 71 357 72 358
rect 70 357 71 358
rect 69 357 70 358
rect 68 357 69 358
rect 67 357 68 358
rect 66 357 67 358
rect 441 358 442 359
rect 440 358 441 359
rect 439 358 440 359
rect 420 358 421 359
rect 419 358 420 359
rect 418 358 419 359
rect 417 358 418 359
rect 400 358 401 359
rect 399 358 400 359
rect 398 358 399 359
rect 397 358 398 359
rect 112 358 113 359
rect 111 358 112 359
rect 110 358 111 359
rect 109 358 110 359
rect 108 358 109 359
rect 107 358 108 359
rect 106 358 107 359
rect 105 358 106 359
rect 104 358 105 359
rect 103 358 104 359
rect 102 358 103 359
rect 101 358 102 359
rect 100 358 101 359
rect 99 358 100 359
rect 98 358 99 359
rect 97 358 98 359
rect 96 358 97 359
rect 95 358 96 359
rect 94 358 95 359
rect 93 358 94 359
rect 92 358 93 359
rect 91 358 92 359
rect 90 358 91 359
rect 89 358 90 359
rect 88 358 89 359
rect 87 358 88 359
rect 86 358 87 359
rect 85 358 86 359
rect 84 358 85 359
rect 83 358 84 359
rect 82 358 83 359
rect 81 358 82 359
rect 80 358 81 359
rect 79 358 80 359
rect 78 358 79 359
rect 77 358 78 359
rect 76 358 77 359
rect 75 358 76 359
rect 74 358 75 359
rect 73 358 74 359
rect 72 358 73 359
rect 71 358 72 359
rect 70 358 71 359
rect 69 358 70 359
rect 68 358 69 359
rect 67 358 68 359
rect 441 359 442 360
rect 440 359 441 360
rect 439 359 440 360
rect 421 359 422 360
rect 420 359 421 360
rect 419 359 420 360
rect 418 359 419 360
rect 417 359 418 360
rect 416 359 417 360
rect 400 359 401 360
rect 399 359 400 360
rect 398 359 399 360
rect 397 359 398 360
rect 113 359 114 360
rect 112 359 113 360
rect 111 359 112 360
rect 110 359 111 360
rect 109 359 110 360
rect 108 359 109 360
rect 107 359 108 360
rect 106 359 107 360
rect 105 359 106 360
rect 104 359 105 360
rect 103 359 104 360
rect 102 359 103 360
rect 101 359 102 360
rect 100 359 101 360
rect 99 359 100 360
rect 98 359 99 360
rect 97 359 98 360
rect 96 359 97 360
rect 95 359 96 360
rect 94 359 95 360
rect 93 359 94 360
rect 92 359 93 360
rect 91 359 92 360
rect 90 359 91 360
rect 89 359 90 360
rect 88 359 89 360
rect 87 359 88 360
rect 86 359 87 360
rect 85 359 86 360
rect 84 359 85 360
rect 83 359 84 360
rect 82 359 83 360
rect 81 359 82 360
rect 80 359 81 360
rect 79 359 80 360
rect 78 359 79 360
rect 77 359 78 360
rect 76 359 77 360
rect 75 359 76 360
rect 74 359 75 360
rect 73 359 74 360
rect 72 359 73 360
rect 71 359 72 360
rect 70 359 71 360
rect 69 359 70 360
rect 441 360 442 361
rect 440 360 441 361
rect 439 360 440 361
rect 424 360 425 361
rect 423 360 424 361
rect 422 360 423 361
rect 421 360 422 361
rect 420 360 421 361
rect 419 360 420 361
rect 418 360 419 361
rect 417 360 418 361
rect 416 360 417 361
rect 415 360 416 361
rect 414 360 415 361
rect 413 360 414 361
rect 400 360 401 361
rect 399 360 400 361
rect 398 360 399 361
rect 397 360 398 361
rect 115 360 116 361
rect 114 360 115 361
rect 113 360 114 361
rect 112 360 113 361
rect 111 360 112 361
rect 110 360 111 361
rect 109 360 110 361
rect 108 360 109 361
rect 107 360 108 361
rect 106 360 107 361
rect 105 360 106 361
rect 104 360 105 361
rect 103 360 104 361
rect 102 360 103 361
rect 101 360 102 361
rect 100 360 101 361
rect 99 360 100 361
rect 98 360 99 361
rect 97 360 98 361
rect 96 360 97 361
rect 95 360 96 361
rect 94 360 95 361
rect 93 360 94 361
rect 92 360 93 361
rect 91 360 92 361
rect 90 360 91 361
rect 89 360 90 361
rect 88 360 89 361
rect 87 360 88 361
rect 86 360 87 361
rect 85 360 86 361
rect 84 360 85 361
rect 83 360 84 361
rect 82 360 83 361
rect 81 360 82 361
rect 80 360 81 361
rect 79 360 80 361
rect 78 360 79 361
rect 77 360 78 361
rect 76 360 77 361
rect 75 360 76 361
rect 74 360 75 361
rect 73 360 74 361
rect 72 360 73 361
rect 71 360 72 361
rect 441 361 442 362
rect 440 361 441 362
rect 439 361 440 362
rect 438 361 439 362
rect 425 361 426 362
rect 424 361 425 362
rect 423 361 424 362
rect 422 361 423 362
rect 421 361 422 362
rect 420 361 421 362
rect 419 361 420 362
rect 418 361 419 362
rect 417 361 418 362
rect 416 361 417 362
rect 415 361 416 362
rect 414 361 415 362
rect 413 361 414 362
rect 412 361 413 362
rect 401 361 402 362
rect 400 361 401 362
rect 399 361 400 362
rect 398 361 399 362
rect 397 361 398 362
rect 117 361 118 362
rect 116 361 117 362
rect 115 361 116 362
rect 114 361 115 362
rect 113 361 114 362
rect 112 361 113 362
rect 111 361 112 362
rect 110 361 111 362
rect 109 361 110 362
rect 108 361 109 362
rect 107 361 108 362
rect 106 361 107 362
rect 105 361 106 362
rect 104 361 105 362
rect 103 361 104 362
rect 102 361 103 362
rect 101 361 102 362
rect 100 361 101 362
rect 99 361 100 362
rect 98 361 99 362
rect 97 361 98 362
rect 96 361 97 362
rect 95 361 96 362
rect 94 361 95 362
rect 93 361 94 362
rect 92 361 93 362
rect 91 361 92 362
rect 90 361 91 362
rect 89 361 90 362
rect 88 361 89 362
rect 87 361 88 362
rect 86 361 87 362
rect 85 361 86 362
rect 84 361 85 362
rect 83 361 84 362
rect 82 361 83 362
rect 81 361 82 362
rect 80 361 81 362
rect 79 361 80 362
rect 78 361 79 362
rect 77 361 78 362
rect 76 361 77 362
rect 75 361 76 362
rect 74 361 75 362
rect 73 361 74 362
rect 441 362 442 363
rect 440 362 441 363
rect 439 362 440 363
rect 438 362 439 363
rect 425 362 426 363
rect 424 362 425 363
rect 423 362 424 363
rect 422 362 423 363
rect 421 362 422 363
rect 420 362 421 363
rect 419 362 420 363
rect 418 362 419 363
rect 417 362 418 363
rect 416 362 417 363
rect 415 362 416 363
rect 414 362 415 363
rect 413 362 414 363
rect 412 362 413 363
rect 402 362 403 363
rect 401 362 402 363
rect 400 362 401 363
rect 399 362 400 363
rect 398 362 399 363
rect 397 362 398 363
rect 119 362 120 363
rect 118 362 119 363
rect 117 362 118 363
rect 116 362 117 363
rect 115 362 116 363
rect 114 362 115 363
rect 113 362 114 363
rect 112 362 113 363
rect 111 362 112 363
rect 110 362 111 363
rect 109 362 110 363
rect 108 362 109 363
rect 107 362 108 363
rect 106 362 107 363
rect 105 362 106 363
rect 104 362 105 363
rect 103 362 104 363
rect 102 362 103 363
rect 101 362 102 363
rect 100 362 101 363
rect 99 362 100 363
rect 98 362 99 363
rect 97 362 98 363
rect 96 362 97 363
rect 95 362 96 363
rect 94 362 95 363
rect 93 362 94 363
rect 92 362 93 363
rect 91 362 92 363
rect 90 362 91 363
rect 89 362 90 363
rect 88 362 89 363
rect 87 362 88 363
rect 86 362 87 363
rect 85 362 86 363
rect 84 362 85 363
rect 83 362 84 363
rect 82 362 83 363
rect 81 362 82 363
rect 80 362 81 363
rect 79 362 80 363
rect 78 362 79 363
rect 77 362 78 363
rect 76 362 77 363
rect 75 362 76 363
rect 441 363 442 364
rect 440 363 441 364
rect 439 363 440 364
rect 438 363 439 364
rect 437 363 438 364
rect 404 363 405 364
rect 403 363 404 364
rect 402 363 403 364
rect 401 363 402 364
rect 400 363 401 364
rect 399 363 400 364
rect 398 363 399 364
rect 397 363 398 364
rect 118 363 119 364
rect 117 363 118 364
rect 116 363 117 364
rect 115 363 116 364
rect 114 363 115 364
rect 113 363 114 364
rect 112 363 113 364
rect 111 363 112 364
rect 110 363 111 364
rect 109 363 110 364
rect 108 363 109 364
rect 107 363 108 364
rect 106 363 107 364
rect 105 363 106 364
rect 104 363 105 364
rect 103 363 104 364
rect 102 363 103 364
rect 101 363 102 364
rect 100 363 101 364
rect 99 363 100 364
rect 98 363 99 364
rect 97 363 98 364
rect 96 363 97 364
rect 95 363 96 364
rect 94 363 95 364
rect 93 363 94 364
rect 92 363 93 364
rect 91 363 92 364
rect 90 363 91 364
rect 89 363 90 364
rect 88 363 89 364
rect 87 363 88 364
rect 86 363 87 364
rect 85 363 86 364
rect 84 363 85 364
rect 83 363 84 364
rect 82 363 83 364
rect 81 363 82 364
rect 80 363 81 364
rect 79 363 80 364
rect 78 363 79 364
rect 441 364 442 365
rect 440 364 441 365
rect 439 364 440 365
rect 438 364 439 365
rect 437 364 438 365
rect 436 364 437 365
rect 407 364 408 365
rect 406 364 407 365
rect 405 364 406 365
rect 404 364 405 365
rect 403 364 404 365
rect 402 364 403 365
rect 401 364 402 365
rect 400 364 401 365
rect 399 364 400 365
rect 398 364 399 365
rect 397 364 398 365
rect 116 364 117 365
rect 115 364 116 365
rect 114 364 115 365
rect 113 364 114 365
rect 112 364 113 365
rect 111 364 112 365
rect 110 364 111 365
rect 109 364 110 365
rect 108 364 109 365
rect 107 364 108 365
rect 106 364 107 365
rect 105 364 106 365
rect 104 364 105 365
rect 103 364 104 365
rect 102 364 103 365
rect 101 364 102 365
rect 100 364 101 365
rect 99 364 100 365
rect 98 364 99 365
rect 97 364 98 365
rect 96 364 97 365
rect 95 364 96 365
rect 94 364 95 365
rect 93 364 94 365
rect 92 364 93 365
rect 91 364 92 365
rect 90 364 91 365
rect 89 364 90 365
rect 88 364 89 365
rect 87 364 88 365
rect 86 364 87 365
rect 85 364 86 365
rect 84 364 85 365
rect 83 364 84 365
rect 82 364 83 365
rect 441 365 442 366
rect 440 365 441 366
rect 439 365 440 366
rect 438 365 439 366
rect 437 365 438 366
rect 436 365 437 366
rect 435 365 436 366
rect 407 365 408 366
rect 406 365 407 366
rect 405 365 406 366
rect 404 365 405 366
rect 403 365 404 366
rect 402 365 403 366
rect 401 365 402 366
rect 400 365 401 366
rect 399 365 400 366
rect 398 365 399 366
rect 397 365 398 366
rect 113 365 114 366
rect 112 365 113 366
rect 111 365 112 366
rect 110 365 111 366
rect 109 365 110 366
rect 108 365 109 366
rect 107 365 108 366
rect 106 365 107 366
rect 105 365 106 366
rect 104 365 105 366
rect 103 365 104 366
rect 102 365 103 366
rect 101 365 102 366
rect 100 365 101 366
rect 99 365 100 366
rect 98 365 99 366
rect 97 365 98 366
rect 96 365 97 366
rect 95 365 96 366
rect 94 365 95 366
rect 93 365 94 366
rect 92 365 93 366
rect 91 365 92 366
rect 90 365 91 366
rect 89 365 90 366
rect 88 365 89 366
rect 87 365 88 366
rect 86 365 87 366
rect 441 366 442 367
rect 440 366 441 367
rect 439 366 440 367
rect 438 366 439 367
rect 437 366 438 367
rect 436 366 437 367
rect 435 366 436 367
rect 434 366 435 367
rect 433 366 434 367
rect 407 366 408 367
rect 406 366 407 367
rect 405 366 406 367
rect 404 366 405 367
rect 403 366 404 367
rect 402 366 403 367
rect 401 366 402 367
rect 400 366 401 367
rect 399 366 400 367
rect 107 366 108 367
rect 106 366 107 367
rect 105 366 106 367
rect 104 366 105 367
rect 103 366 104 367
rect 102 366 103 367
rect 101 366 102 367
rect 100 366 101 367
rect 99 366 100 367
rect 98 366 99 367
rect 97 366 98 367
rect 96 366 97 367
rect 95 366 96 367
rect 94 366 95 367
rect 93 366 94 367
rect 441 367 442 368
rect 440 367 441 368
rect 439 367 440 368
rect 438 367 439 368
rect 437 367 438 368
rect 436 367 437 368
rect 435 367 436 368
rect 434 367 435 368
rect 433 367 434 368
rect 432 367 433 368
rect 431 367 432 368
rect 440 368 441 369
rect 439 368 440 369
rect 438 368 439 369
rect 437 368 438 369
rect 436 368 437 369
rect 435 368 436 369
rect 434 368 435 369
rect 433 368 434 369
rect 432 368 433 369
rect 431 368 432 369
rect 430 368 431 369
rect 435 369 436 370
rect 434 369 435 370
rect 433 369 434 370
rect 432 369 433 370
rect 431 369 432 370
rect 430 369 431 370
rect 441 376 442 377
rect 440 376 441 377
rect 441 377 442 378
rect 440 377 441 378
rect 439 377 440 378
rect 399 377 400 378
rect 398 377 399 378
rect 397 377 398 378
rect 441 378 442 379
rect 440 378 441 379
rect 439 378 440 379
rect 399 378 400 379
rect 398 378 399 379
rect 397 378 398 379
rect 441 379 442 380
rect 440 379 441 380
rect 439 379 440 380
rect 399 379 400 380
rect 398 379 399 380
rect 397 379 398 380
rect 441 380 442 381
rect 440 380 441 381
rect 439 380 440 381
rect 399 380 400 381
rect 398 380 399 381
rect 397 380 398 381
rect 441 381 442 382
rect 440 381 441 382
rect 439 381 440 382
rect 438 381 439 382
rect 400 381 401 382
rect 399 381 400 382
rect 398 381 399 382
rect 397 381 398 382
rect 441 382 442 383
rect 440 382 441 383
rect 439 382 440 383
rect 438 382 439 383
rect 437 382 438 383
rect 436 382 437 383
rect 435 382 436 383
rect 434 382 435 383
rect 433 382 434 383
rect 432 382 433 383
rect 431 382 432 383
rect 430 382 431 383
rect 429 382 430 383
rect 428 382 429 383
rect 427 382 428 383
rect 426 382 427 383
rect 425 382 426 383
rect 424 382 425 383
rect 423 382 424 383
rect 422 382 423 383
rect 421 382 422 383
rect 420 382 421 383
rect 419 382 420 383
rect 418 382 419 383
rect 417 382 418 383
rect 416 382 417 383
rect 415 382 416 383
rect 414 382 415 383
rect 413 382 414 383
rect 412 382 413 383
rect 411 382 412 383
rect 410 382 411 383
rect 409 382 410 383
rect 408 382 409 383
rect 407 382 408 383
rect 406 382 407 383
rect 405 382 406 383
rect 404 382 405 383
rect 403 382 404 383
rect 402 382 403 383
rect 401 382 402 383
rect 400 382 401 383
rect 399 382 400 383
rect 398 382 399 383
rect 397 382 398 383
rect 441 383 442 384
rect 440 383 441 384
rect 439 383 440 384
rect 438 383 439 384
rect 437 383 438 384
rect 436 383 437 384
rect 435 383 436 384
rect 434 383 435 384
rect 433 383 434 384
rect 432 383 433 384
rect 431 383 432 384
rect 430 383 431 384
rect 429 383 430 384
rect 428 383 429 384
rect 427 383 428 384
rect 426 383 427 384
rect 425 383 426 384
rect 424 383 425 384
rect 423 383 424 384
rect 422 383 423 384
rect 421 383 422 384
rect 420 383 421 384
rect 419 383 420 384
rect 418 383 419 384
rect 417 383 418 384
rect 416 383 417 384
rect 415 383 416 384
rect 414 383 415 384
rect 413 383 414 384
rect 412 383 413 384
rect 411 383 412 384
rect 410 383 411 384
rect 409 383 410 384
rect 408 383 409 384
rect 407 383 408 384
rect 406 383 407 384
rect 405 383 406 384
rect 404 383 405 384
rect 403 383 404 384
rect 402 383 403 384
rect 401 383 402 384
rect 400 383 401 384
rect 399 383 400 384
rect 398 383 399 384
rect 397 383 398 384
rect 441 384 442 385
rect 440 384 441 385
rect 439 384 440 385
rect 438 384 439 385
rect 437 384 438 385
rect 436 384 437 385
rect 435 384 436 385
rect 434 384 435 385
rect 433 384 434 385
rect 432 384 433 385
rect 431 384 432 385
rect 430 384 431 385
rect 429 384 430 385
rect 428 384 429 385
rect 427 384 428 385
rect 426 384 427 385
rect 425 384 426 385
rect 424 384 425 385
rect 423 384 424 385
rect 422 384 423 385
rect 421 384 422 385
rect 420 384 421 385
rect 419 384 420 385
rect 418 384 419 385
rect 417 384 418 385
rect 416 384 417 385
rect 415 384 416 385
rect 414 384 415 385
rect 413 384 414 385
rect 412 384 413 385
rect 411 384 412 385
rect 410 384 411 385
rect 409 384 410 385
rect 408 384 409 385
rect 407 384 408 385
rect 406 384 407 385
rect 405 384 406 385
rect 404 384 405 385
rect 403 384 404 385
rect 402 384 403 385
rect 401 384 402 385
rect 400 384 401 385
rect 399 384 400 385
rect 398 384 399 385
rect 397 384 398 385
rect 441 385 442 386
rect 440 385 441 386
rect 439 385 440 386
rect 438 385 439 386
rect 437 385 438 386
rect 436 385 437 386
rect 435 385 436 386
rect 434 385 435 386
rect 433 385 434 386
rect 432 385 433 386
rect 431 385 432 386
rect 430 385 431 386
rect 429 385 430 386
rect 428 385 429 386
rect 427 385 428 386
rect 426 385 427 386
rect 425 385 426 386
rect 424 385 425 386
rect 423 385 424 386
rect 422 385 423 386
rect 421 385 422 386
rect 420 385 421 386
rect 419 385 420 386
rect 418 385 419 386
rect 417 385 418 386
rect 416 385 417 386
rect 415 385 416 386
rect 414 385 415 386
rect 413 385 414 386
rect 412 385 413 386
rect 411 385 412 386
rect 410 385 411 386
rect 409 385 410 386
rect 408 385 409 386
rect 407 385 408 386
rect 406 385 407 386
rect 405 385 406 386
rect 404 385 405 386
rect 403 385 404 386
rect 402 385 403 386
rect 401 385 402 386
rect 400 385 401 386
rect 399 385 400 386
rect 398 385 399 386
rect 397 385 398 386
rect 441 386 442 387
rect 440 386 441 387
rect 439 386 440 387
rect 438 386 439 387
rect 437 386 438 387
rect 436 386 437 387
rect 435 386 436 387
rect 434 386 435 387
rect 433 386 434 387
rect 432 386 433 387
rect 431 386 432 387
rect 430 386 431 387
rect 429 386 430 387
rect 428 386 429 387
rect 427 386 428 387
rect 426 386 427 387
rect 425 386 426 387
rect 424 386 425 387
rect 423 386 424 387
rect 422 386 423 387
rect 421 386 422 387
rect 420 386 421 387
rect 419 386 420 387
rect 418 386 419 387
rect 417 386 418 387
rect 416 386 417 387
rect 415 386 416 387
rect 414 386 415 387
rect 413 386 414 387
rect 412 386 413 387
rect 411 386 412 387
rect 410 386 411 387
rect 409 386 410 387
rect 408 386 409 387
rect 407 386 408 387
rect 406 386 407 387
rect 405 386 406 387
rect 404 386 405 387
rect 403 386 404 387
rect 402 386 403 387
rect 401 386 402 387
rect 400 386 401 387
rect 399 386 400 387
rect 398 386 399 387
rect 397 386 398 387
rect 441 387 442 388
rect 440 387 441 388
rect 439 387 440 388
rect 438 387 439 388
rect 437 387 438 388
rect 436 387 437 388
rect 435 387 436 388
rect 434 387 435 388
rect 433 387 434 388
rect 432 387 433 388
rect 431 387 432 388
rect 430 387 431 388
rect 429 387 430 388
rect 428 387 429 388
rect 427 387 428 388
rect 426 387 427 388
rect 425 387 426 388
rect 424 387 425 388
rect 423 387 424 388
rect 422 387 423 388
rect 421 387 422 388
rect 420 387 421 388
rect 419 387 420 388
rect 418 387 419 388
rect 417 387 418 388
rect 416 387 417 388
rect 415 387 416 388
rect 414 387 415 388
rect 413 387 414 388
rect 412 387 413 388
rect 411 387 412 388
rect 410 387 411 388
rect 409 387 410 388
rect 408 387 409 388
rect 407 387 408 388
rect 406 387 407 388
rect 405 387 406 388
rect 404 387 405 388
rect 403 387 404 388
rect 402 387 403 388
rect 401 387 402 388
rect 400 387 401 388
rect 399 387 400 388
rect 398 387 399 388
rect 397 387 398 388
rect 441 388 442 389
rect 440 388 441 389
rect 439 388 440 389
rect 438 388 439 389
rect 437 388 438 389
rect 436 388 437 389
rect 435 388 436 389
rect 434 388 435 389
rect 433 388 434 389
rect 432 388 433 389
rect 431 388 432 389
rect 430 388 431 389
rect 429 388 430 389
rect 428 388 429 389
rect 427 388 428 389
rect 426 388 427 389
rect 425 388 426 389
rect 424 388 425 389
rect 423 388 424 389
rect 422 388 423 389
rect 421 388 422 389
rect 420 388 421 389
rect 419 388 420 389
rect 418 388 419 389
rect 417 388 418 389
rect 416 388 417 389
rect 415 388 416 389
rect 414 388 415 389
rect 413 388 414 389
rect 412 388 413 389
rect 411 388 412 389
rect 410 388 411 389
rect 409 388 410 389
rect 408 388 409 389
rect 407 388 408 389
rect 406 388 407 389
rect 405 388 406 389
rect 404 388 405 389
rect 403 388 404 389
rect 402 388 403 389
rect 401 388 402 389
rect 400 388 401 389
rect 399 388 400 389
rect 398 388 399 389
rect 397 388 398 389
rect 441 389 442 390
rect 440 389 441 390
rect 439 389 440 390
rect 438 389 439 390
rect 437 389 438 390
rect 436 389 437 390
rect 435 389 436 390
rect 434 389 435 390
rect 433 389 434 390
rect 432 389 433 390
rect 431 389 432 390
rect 430 389 431 390
rect 429 389 430 390
rect 428 389 429 390
rect 427 389 428 390
rect 426 389 427 390
rect 425 389 426 390
rect 424 389 425 390
rect 423 389 424 390
rect 422 389 423 390
rect 421 389 422 390
rect 420 389 421 390
rect 419 389 420 390
rect 418 389 419 390
rect 417 389 418 390
rect 416 389 417 390
rect 415 389 416 390
rect 414 389 415 390
rect 413 389 414 390
rect 412 389 413 390
rect 411 389 412 390
rect 410 389 411 390
rect 409 389 410 390
rect 408 389 409 390
rect 407 389 408 390
rect 406 389 407 390
rect 405 389 406 390
rect 404 389 405 390
rect 403 389 404 390
rect 402 389 403 390
rect 401 389 402 390
rect 400 389 401 390
rect 399 389 400 390
rect 398 389 399 390
rect 397 389 398 390
rect 441 390 442 391
rect 440 390 441 391
rect 439 390 440 391
rect 438 390 439 391
rect 437 390 438 391
rect 436 390 437 391
rect 435 390 436 391
rect 434 390 435 391
rect 433 390 434 391
rect 432 390 433 391
rect 431 390 432 391
rect 430 390 431 391
rect 429 390 430 391
rect 428 390 429 391
rect 427 390 428 391
rect 426 390 427 391
rect 425 390 426 391
rect 424 390 425 391
rect 423 390 424 391
rect 422 390 423 391
rect 421 390 422 391
rect 420 390 421 391
rect 419 390 420 391
rect 418 390 419 391
rect 417 390 418 391
rect 416 390 417 391
rect 415 390 416 391
rect 414 390 415 391
rect 413 390 414 391
rect 412 390 413 391
rect 411 390 412 391
rect 410 390 411 391
rect 409 390 410 391
rect 408 390 409 391
rect 407 390 408 391
rect 406 390 407 391
rect 405 390 406 391
rect 404 390 405 391
rect 403 390 404 391
rect 402 390 403 391
rect 401 390 402 391
rect 400 390 401 391
rect 399 390 400 391
rect 398 390 399 391
rect 397 390 398 391
rect 441 391 442 392
rect 440 391 441 392
rect 439 391 440 392
rect 438 391 439 392
rect 437 391 438 392
rect 436 391 437 392
rect 435 391 436 392
rect 434 391 435 392
rect 433 391 434 392
rect 432 391 433 392
rect 431 391 432 392
rect 430 391 431 392
rect 429 391 430 392
rect 428 391 429 392
rect 427 391 428 392
rect 426 391 427 392
rect 425 391 426 392
rect 424 391 425 392
rect 423 391 424 392
rect 422 391 423 392
rect 421 391 422 392
rect 420 391 421 392
rect 419 391 420 392
rect 418 391 419 392
rect 417 391 418 392
rect 416 391 417 392
rect 415 391 416 392
rect 414 391 415 392
rect 413 391 414 392
rect 412 391 413 392
rect 411 391 412 392
rect 410 391 411 392
rect 409 391 410 392
rect 408 391 409 392
rect 407 391 408 392
rect 406 391 407 392
rect 405 391 406 392
rect 404 391 405 392
rect 403 391 404 392
rect 402 391 403 392
rect 401 391 402 392
rect 400 391 401 392
rect 399 391 400 392
rect 398 391 399 392
rect 397 391 398 392
rect 441 392 442 393
rect 440 392 441 393
rect 439 392 440 393
rect 438 392 439 393
rect 437 392 438 393
rect 420 392 421 393
rect 419 392 420 393
rect 418 392 419 393
rect 417 392 418 393
rect 400 392 401 393
rect 399 392 400 393
rect 398 392 399 393
rect 397 392 398 393
rect 441 393 442 394
rect 440 393 441 394
rect 439 393 440 394
rect 438 393 439 394
rect 420 393 421 394
rect 419 393 420 394
rect 418 393 419 394
rect 417 393 418 394
rect 399 393 400 394
rect 398 393 399 394
rect 397 393 398 394
rect 441 394 442 395
rect 440 394 441 395
rect 439 394 440 395
rect 420 394 421 395
rect 419 394 420 395
rect 418 394 419 395
rect 417 394 418 395
rect 399 394 400 395
rect 398 394 399 395
rect 397 394 398 395
rect 441 395 442 396
rect 440 395 441 396
rect 439 395 440 396
rect 420 395 421 396
rect 419 395 420 396
rect 418 395 419 396
rect 417 395 418 396
rect 399 395 400 396
rect 398 395 399 396
rect 397 395 398 396
rect 441 396 442 397
rect 440 396 441 397
rect 439 396 440 397
rect 420 396 421 397
rect 419 396 420 397
rect 418 396 419 397
rect 417 396 418 397
rect 399 396 400 397
rect 398 396 399 397
rect 397 396 398 397
rect 441 397 442 398
rect 440 397 441 398
rect 439 397 440 398
rect 420 397 421 398
rect 419 397 420 398
rect 418 397 419 398
rect 417 397 418 398
rect 399 397 400 398
rect 398 397 399 398
rect 397 397 398 398
rect 441 398 442 399
rect 440 398 441 399
rect 439 398 440 399
rect 420 398 421 399
rect 419 398 420 399
rect 418 398 419 399
rect 417 398 418 399
rect 399 398 400 399
rect 398 398 399 399
rect 397 398 398 399
rect 441 399 442 400
rect 440 399 441 400
rect 439 399 440 400
rect 420 399 421 400
rect 419 399 420 400
rect 418 399 419 400
rect 417 399 418 400
rect 399 399 400 400
rect 398 399 399 400
rect 397 399 398 400
rect 441 400 442 401
rect 440 400 441 401
rect 439 400 440 401
rect 420 400 421 401
rect 419 400 420 401
rect 418 400 419 401
rect 417 400 418 401
rect 399 400 400 401
rect 398 400 399 401
rect 397 400 398 401
rect 441 401 442 402
rect 440 401 441 402
rect 439 401 440 402
rect 420 401 421 402
rect 419 401 420 402
rect 418 401 419 402
rect 417 401 418 402
rect 400 401 401 402
rect 399 401 400 402
rect 398 401 399 402
rect 397 401 398 402
rect 441 402 442 403
rect 440 402 441 403
rect 439 402 440 403
rect 421 402 422 403
rect 420 402 421 403
rect 419 402 420 403
rect 418 402 419 403
rect 417 402 418 403
rect 416 402 417 403
rect 400 402 401 403
rect 399 402 400 403
rect 398 402 399 403
rect 397 402 398 403
rect 441 403 442 404
rect 440 403 441 404
rect 439 403 440 404
rect 423 403 424 404
rect 422 403 423 404
rect 421 403 422 404
rect 420 403 421 404
rect 419 403 420 404
rect 418 403 419 404
rect 417 403 418 404
rect 416 403 417 404
rect 415 403 416 404
rect 414 403 415 404
rect 400 403 401 404
rect 399 403 400 404
rect 398 403 399 404
rect 397 403 398 404
rect 441 404 442 405
rect 440 404 441 405
rect 439 404 440 405
rect 438 404 439 405
rect 425 404 426 405
rect 424 404 425 405
rect 423 404 424 405
rect 422 404 423 405
rect 421 404 422 405
rect 420 404 421 405
rect 419 404 420 405
rect 418 404 419 405
rect 417 404 418 405
rect 416 404 417 405
rect 415 404 416 405
rect 414 404 415 405
rect 413 404 414 405
rect 412 404 413 405
rect 401 404 402 405
rect 400 404 401 405
rect 399 404 400 405
rect 398 404 399 405
rect 397 404 398 405
rect 441 405 442 406
rect 440 405 441 406
rect 439 405 440 406
rect 438 405 439 406
rect 425 405 426 406
rect 424 405 425 406
rect 423 405 424 406
rect 422 405 423 406
rect 421 405 422 406
rect 420 405 421 406
rect 419 405 420 406
rect 418 405 419 406
rect 417 405 418 406
rect 416 405 417 406
rect 415 405 416 406
rect 414 405 415 406
rect 413 405 414 406
rect 412 405 413 406
rect 402 405 403 406
rect 401 405 402 406
rect 400 405 401 406
rect 399 405 400 406
rect 398 405 399 406
rect 397 405 398 406
rect 441 406 442 407
rect 440 406 441 407
rect 439 406 440 407
rect 438 406 439 407
rect 437 406 438 407
rect 425 406 426 407
rect 424 406 425 407
rect 423 406 424 407
rect 422 406 423 407
rect 421 406 422 407
rect 420 406 421 407
rect 419 406 420 407
rect 418 406 419 407
rect 417 406 418 407
rect 416 406 417 407
rect 415 406 416 407
rect 414 406 415 407
rect 413 406 414 407
rect 412 406 413 407
rect 404 406 405 407
rect 403 406 404 407
rect 402 406 403 407
rect 401 406 402 407
rect 400 406 401 407
rect 399 406 400 407
rect 398 406 399 407
rect 397 406 398 407
rect 441 407 442 408
rect 440 407 441 408
rect 439 407 440 408
rect 438 407 439 408
rect 437 407 438 408
rect 436 407 437 408
rect 407 407 408 408
rect 406 407 407 408
rect 405 407 406 408
rect 404 407 405 408
rect 403 407 404 408
rect 402 407 403 408
rect 401 407 402 408
rect 400 407 401 408
rect 399 407 400 408
rect 398 407 399 408
rect 397 407 398 408
rect 441 408 442 409
rect 440 408 441 409
rect 439 408 440 409
rect 438 408 439 409
rect 437 408 438 409
rect 436 408 437 409
rect 435 408 436 409
rect 407 408 408 409
rect 406 408 407 409
rect 405 408 406 409
rect 404 408 405 409
rect 403 408 404 409
rect 402 408 403 409
rect 401 408 402 409
rect 400 408 401 409
rect 399 408 400 409
rect 398 408 399 409
rect 397 408 398 409
rect 441 409 442 410
rect 440 409 441 410
rect 439 409 440 410
rect 438 409 439 410
rect 437 409 438 410
rect 436 409 437 410
rect 435 409 436 410
rect 434 409 435 410
rect 433 409 434 410
rect 407 409 408 410
rect 406 409 407 410
rect 405 409 406 410
rect 404 409 405 410
rect 403 409 404 410
rect 402 409 403 410
rect 401 409 402 410
rect 400 409 401 410
rect 399 409 400 410
rect 398 409 399 410
rect 397 409 398 410
rect 441 410 442 411
rect 440 410 441 411
rect 439 410 440 411
rect 438 410 439 411
rect 437 410 438 411
rect 436 410 437 411
rect 435 410 436 411
rect 434 410 435 411
rect 433 410 434 411
rect 432 410 433 411
rect 431 410 432 411
rect 440 411 441 412
rect 439 411 440 412
rect 438 411 439 412
rect 437 411 438 412
rect 436 411 437 412
rect 435 411 436 412
rect 434 411 435 412
rect 433 411 434 412
rect 432 411 433 412
rect 431 411 432 412
rect 430 411 431 412
rect 436 412 437 413
rect 435 412 436 413
rect 434 412 435 413
rect 433 412 434 413
rect 432 412 433 413
rect 431 412 432 413
rect 430 412 431 413
rect 431 413 432 414
rect 430 413 431 414
<< end >>
