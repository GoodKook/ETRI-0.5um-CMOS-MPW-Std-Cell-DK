magic
tech scmos
magscale 1 30
timestamp 1727178509
<< checkpaint >>
rect 18300 186927 44800 197000
rect 13915 181835 44800 186927
rect 46919 186419 142100 190000
rect 46919 181835 143266 186419
rect 6771 176042 185015 181835
rect 6771 175958 328570 176042
rect 205 167042 328570 175958
rect 205 160774 185015 167042
rect 6771 143081 185015 160774
rect 0 142100 185015 143081
rect 0 102896 190000 142100
rect -13866 102380 190000 102896
rect -25613 89180 190000 102380
rect -24170 89077 190000 89180
rect -17472 83925 190000 89077
rect 0 47900 190000 83925
rect 6771 46919 190000 47900
rect 6771 32547 185015 46919
rect 6771 31724 186496 32547
rect -4457 10781 186496 31724
rect -4457 8670 185015 10781
rect -4457 7765 35955 8670
rect 205 1458 35955 7765
rect -600 -600 630 630
rect 46919 0 142100 8670
<< metal1 >>
rect 51100 145800 57800 145900
rect 48500 142000 57800 144500
rect 142400 131900 144600 140200
rect 44800 129600 47500 129800
rect 45600 127200 45700 128900
rect 44100 51200 44200 57800
rect 45400 51200 48700 57800
<< m2contact >>
rect 51100 144500 57800 145800
rect 144600 131900 145800 140200
rect 44800 129800 47500 130100
rect 45300 127200 45600 128900
rect 46400 127500 46700 128300
rect 44200 51200 45400 57800
<< metal2 >>
rect 51100 145800 57800 145900
rect 73300 143000 73700 145900
rect 86800 143600 87200 145900
rect 100300 144200 100700 145900
rect 113800 144800 114200 145900
rect 127300 145400 127700 145900
rect 140800 145400 141200 145900
rect 100300 143900 107500 144200
rect 118100 143900 124100 144200
rect 96500 143300 105100 143600
rect 116800 143300 122600 143600
rect 74200 142700 81100 143000
rect 92800 142700 99700 143000
rect 122200 142700 122600 143300
rect 123700 142700 124100 143900
rect 126100 142700 126500 144500
rect 136600 142700 137000 145100
rect 137200 145100 141200 145400
rect 137200 142700 137600 145100
rect 138100 143800 143900 144200
rect 138100 142700 138500 143800
rect 139400 143100 143300 143500
rect 139400 142700 139800 143100
rect 44200 131400 45300 136100
rect 145800 131900 145900 140200
rect 44800 130100 45300 131400
rect 45300 122600 45600 127200
rect 44100 117900 45600 122600
rect 46400 109100 46700 127500
rect 144200 126300 144500 130600
rect 144800 127700 145100 131200
rect 144800 127300 145900 127700
rect 144200 126000 145100 126300
rect 44100 104400 46700 109100
rect 44100 100100 47400 100500
rect 47100 90300 47400 100100
rect 142600 99300 142900 113200
rect 143200 109300 143500 119700
rect 143800 110900 144100 121200
rect 144800 114200 145100 126000
rect 144800 113800 145900 114200
rect 144100 100300 145900 100700
rect 143200 87200 143500 96500
rect 44100 86600 45700 87000
rect 143200 86800 145900 87200
rect 45400 82100 45700 86600
rect 142600 73700 142900 82500
rect 44100 73100 45600 73500
rect 142600 73300 145900 73700
rect 45300 66600 45600 73100
rect 143600 59800 145900 60200
rect 44100 51200 44200 57800
rect 64500 47700 77300 48000
rect 93300 47700 104600 48000
rect 49000 44100 49400 47700
rect 125000 47400 125400 47900
rect 63400 47100 76900 47400
rect 92300 47100 105800 47400
rect 117900 47100 125400 47400
rect 62500 44100 62900 47100
rect 130400 46800 130800 48000
rect 76900 46500 90400 46800
rect 91300 46500 104900 46800
rect 118800 46500 130800 46800
rect 76000 44100 76400 46500
rect 132500 46200 132800 48000
rect 90400 45900 103900 46200
rect 120200 45900 132800 46200
rect 89500 44100 89900 45900
rect 134500 45600 134800 48000
rect 103900 45300 115300 45600
rect 132300 45300 134800 45600
rect 103000 44100 103400 45300
rect 136300 45000 136600 48000
rect 142700 47000 143000 55000
rect 116500 44700 123600 45000
rect 124500 44700 135700 45000
rect 116500 44100 116900 44700
rect 140800 44100 141300 46100
<< m3contact >>
rect 127300 145100 128100 145400
rect 136200 145100 137000 145400
rect 113800 144500 114700 144800
rect 125700 144500 126500 144800
rect 107500 143900 108400 144200
rect 117200 143900 118100 144200
rect 86800 143300 87700 143600
rect 95600 143300 96500 143600
rect 105100 143300 106000 143600
rect 115900 143300 116800 143600
rect 73300 142700 74200 143000
rect 81100 142700 82000 143000
rect 91900 142700 92800 143000
rect 143300 142600 143600 143500
rect 143900 143300 144200 144200
rect 143900 131200 145100 131500
rect 143300 130600 144500 130900
rect 143800 121200 144100 122100
rect 143200 119700 143500 120600
rect 142600 113200 142900 114100
rect 143800 110000 144100 110900
rect 143200 108400 143500 109300
rect 143800 100300 144100 101200
rect 142600 98400 142900 99300
rect 47100 89300 47400 90300
rect 143200 96500 143500 97400
rect 45400 81100 45700 82100
rect 142600 82500 142900 83400
rect 45300 65700 45600 66600
rect 143300 59800 143600 60600
rect 142700 55000 143000 55800
rect 49000 47700 49900 48000
rect 63600 47700 64500 48000
rect 77300 47700 78200 48000
rect 92400 47700 93300 48000
rect 104600 47700 105500 48000
rect 118900 47700 119700 48000
rect 62500 47100 63400 47400
rect 76900 47100 77800 47400
rect 91400 47100 92300 47400
rect 105800 47100 106700 47400
rect 117000 47100 117900 47400
rect 76000 46500 76900 46800
rect 90400 46500 91300 46800
rect 104900 46500 105800 46800
rect 117900 46500 118800 46800
rect 89500 45900 90400 46200
rect 103900 45900 104800 46200
rect 119300 45900 120200 46200
rect 103000 45300 103900 45600
rect 115300 45300 116200 45600
rect 131400 45300 132300 45600
rect 123600 44700 124500 45000
rect 135700 44700 136600 45000
rect 140800 46100 141700 46600
rect 142700 46100 143000 47000
<< metal3 >>
rect 128100 145100 136200 145400
rect 114700 144500 125700 144800
rect 108400 143900 117200 144200
rect 87700 143300 95600 143600
rect 106000 143300 115900 143600
rect 82000 142700 91900 143000
rect 143300 130900 143600 142600
rect 143900 131500 144200 143300
rect 142100 129600 144100 130000
rect 142500 127300 143500 127600
rect 142600 114100 142900 126100
rect 143200 120600 143500 127300
rect 143800 122100 144100 129600
rect 47100 82400 47400 89300
rect 142600 83400 142900 98400
rect 143200 97400 143500 108400
rect 143800 101200 144100 110000
rect 47100 82000 49200 82400
rect 45700 81100 49200 81500
rect 142500 69100 143600 69400
rect 45600 65700 49200 66100
rect 142100 61900 143000 62200
rect 142700 55800 143000 61900
rect 143300 60600 143600 69100
rect 49900 47700 63600 48000
rect 78200 47700 92400 48000
rect 105500 47700 118900 48000
rect 77800 47100 91400 47400
rect 106700 47100 117000 47400
rect 105800 46500 117900 46800
rect 104800 45900 119300 46200
rect 141700 46100 142700 46600
rect 116200 45300 131400 45600
use PIC  ABCMD_I_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use PIC  ABCMD_I_1
timestamp 1555589239
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use PIC  ABCMD_I_2
timestamp 1555589239
transform 0 -1 171100 1 0 89000
box -100 -9150 12100 25300
use PIC  ABCMD_I_3
timestamp 1555589239
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use PIC  ABCMD_I_4
timestamp 1555589239
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use PIC  ABCMD_I_5
timestamp 1555589239
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use PIC  ABCMD_I_6
timestamp 1555589239
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use PIC  ABCMD_I_7
timestamp 1555589239
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use POB8  ACC_O_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 0 1 18900 -1 0 101000
box -100 -9150 12100 25300
use POB8  ACC_O_1
timestamp 1555589239
transform 0 1 18900 -1 0 87500
box -100 -9150 12100 25300
use POB8  ACC_O_2
timestamp 1555589239
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use POB8  ACC_O_3
timestamp 1555589239
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use POB8  ACC_O_4
timestamp 1555589239
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use POB8  ACC_O_5
timestamp 1555589239
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use POB8  ACC_O_6
timestamp 1555589239
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use POB8  ACC_O_7
timestamp 1555589239
transform 1 0 48500 0 1 18900
box -100 -9150 12100 25300
use ALU_wrapper_Core  ALU_wrapper_Core_0
timestamp 1727158408
transform 1 0 49445 0 1 48260
box -945 -360 93165 94560
use PIC  CLK
timestamp 1555589239
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
use POB8  DONE_O
timestamp 1555589239
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI050
timestamp 1725930584
transform 0 -1 171100 -1 0 75646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_1
timestamp 1725930584
transform 0 -1 171098 -1 0 62146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_2
timestamp 1725930584
transform 0 -1 171100 -1 0 102646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_3
timestamp 1725930584
transform 0 -1 171100 -1 0 89146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_4
timestamp 1725930584
transform 0 -1 171102 -1 0 129646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_5
timestamp 1725930584
transform 0 -1 171100 -1 0 116146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_6
timestamp 1725930584
transform 1 0 73845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_7
timestamp 1725930584
transform 1 0 60345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_8
timestamp 1725930584
transform 1 0 100845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_9
timestamp 1725930584
transform 1 0 87345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_10
timestamp 1725930584
transform 1 0 127845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_11
timestamp 1725930584
transform 1 0 114345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_12
timestamp 1725930584
transform 0 1 18899 -1 0 75655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_13
timestamp 1725930584
transform 0 1 18899 -1 0 62155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_14
timestamp 1725930584
transform 0 1 18900 -1 0 102655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_15
timestamp 1725930584
transform 0 1 18900 -1 0 89155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_16
timestamp 1725930584
transform 1 0 73845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_17
timestamp 1725930584
transform 0 1 18897 -1 0 116155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_18
timestamp 1725930584
transform 0 1 18900 -1 0 129655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_19
timestamp 1725930584
transform 1 0 60345 0 -1 171101
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_20
timestamp 1725930584
transform 1 0 100845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_21
timestamp 1725930584
transform 1 0 87344 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_22
timestamp 1725930584
transform 1 0 127845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_23
timestamp 1725930584
transform 1 0 114345 0 -1 171100
box -60 0 1860 25060
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 1 0 43621 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1555589239
transform 1 0 141360 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1555589239
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1555589239
transform 1 0 43638 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1555589239
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1555589239
transform 0 1 18900 -1 0 146379
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1555589239
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1555589239
transform 0 -1 171100 -1 0 146346
box -35 0 5035 25060
use PIC  LOADA_I
timestamp 1555589239
transform 0 -1 171100 1 0 102500
box -100 -9150 12100 25300
use PIC  LOADB_I
timestamp 1555589239
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use PIC  LOADCMD_I
timestamp 1555589239
transform 1 0 129500 0 -1 171100
box -100 -9150 12100 25300
use MY_LOGO  MY_LOGO_0
timestamp 1700409309
transform 1 0 144900 0 1 10300
box 0 0 20340 7290
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1555589239
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1555589239
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1555589239
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use pnp5  pnp5_0 ~/ETRI050_DesignKit/analog_ETRI/GDS_Magic
timestamp 1555596690
transform 1 0 44350 0 1 125850
box 450 450 3950 3950
use PANA  PNP_B ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use PANA  PNP_C
timestamp 1555589239
transform 0 1 18900 -1 0 141500
box -100 -9150 12100 25300
use PANA  PNP_E
timestamp 1555589239
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use PIC  RESET
timestamp 1555589239
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
use PVDD  VDD_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 1 0 48500 0 -1 171100
box -100 -9150 12100 25300
use PVDD  VDD_1
timestamp 1555589239
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use PVSS  VSS_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1555589239
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
<< end >>
