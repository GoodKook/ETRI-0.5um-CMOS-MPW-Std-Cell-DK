magic
tech scmos
magscale 1 2
timestamp 1727268294
<< nwell >>
rect -12 154 112 272
<< ntransistor >>
rect 24 14 28 54
rect 34 14 38 54
rect 54 14 58 34
<< ptransistor >>
rect 20 166 24 246
rect 40 166 44 246
rect 60 166 64 246
<< ndiffusion >>
rect 22 14 24 54
rect 28 14 34 54
rect 38 34 49 54
rect 38 14 40 34
rect 52 14 54 34
rect 58 14 60 34
<< pdiffusion >>
rect 18 174 20 246
rect 6 166 20 174
rect 24 178 26 246
rect 38 178 40 246
rect 24 166 40 178
rect 44 166 46 246
rect 58 166 60 246
rect 64 166 66 246
<< ndcontact >>
rect 10 14 22 54
rect 40 14 52 34
rect 60 14 72 34
<< pdcontact >>
rect 6 174 18 246
rect 26 178 38 246
rect 46 166 58 246
rect 66 166 78 246
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 254 106 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 20 152 24 166
rect 40 152 44 166
rect 9 146 24 152
rect 30 146 44 152
rect 9 123 15 146
rect 30 129 36 146
rect 60 123 64 166
rect 10 64 16 111
rect 30 82 36 117
rect 56 111 64 123
rect 30 72 38 82
rect 10 58 28 64
rect 24 54 28 58
rect 34 54 38 72
rect 54 34 58 111
rect 24 10 28 14
rect 34 10 38 14
rect 54 10 58 14
<< polycontact >>
rect 4 111 16 123
rect 24 117 36 129
rect 44 111 56 123
<< metal1 >>
rect -6 266 106 268
rect -6 252 106 254
rect 26 246 38 252
rect 6 172 18 174
rect 6 166 46 172
rect 68 117 74 166
rect 68 54 74 103
rect 40 46 74 54
rect 40 34 52 46
rect 10 8 22 14
rect 60 8 72 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m2contact >>
rect 3 123 17 137
rect 43 123 57 137
rect 23 103 37 117
rect 63 103 77 117
<< metal2 >>
rect 6 137 14 154
rect 46 137 54 154
rect 26 86 34 103
rect 66 86 74 103
<< m1p >>
rect -6 252 106 268
rect -6 -8 106 8
<< m2p >>
rect 6 137 14 154
rect 46 137 54 154
rect 26 86 34 103
rect 66 86 74 103
<< labels >>
rlabel metal1 -6 252 86 268 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -6 -8 86 8 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal2 30 91 30 91 1 B
port 2 n signal input
rlabel metal2 70 89 70 89 1 Y
port 4 n signal output
rlabel metal2 10 151 10 151 1 A
port 1 n signal input
rlabel metal2 50 151 50 151 1 C
port 3 n signal input
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
