VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO counter16
  CLASS BLOCK ;
  FOREIGN counter16 ;
  ORIGIN 6.000 6.000 ;
  SIZE 375.000 BY 366.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 351.300 372.450 353.700 ;
        RECT 363.450 275.700 372.450 351.300 ;
        RECT 0.600 273.300 372.450 275.700 ;
        RECT 363.450 197.700 372.450 273.300 ;
        RECT 0.600 195.300 372.450 197.700 ;
        RECT 363.450 119.700 372.450 195.300 ;
        RECT 0.600 117.300 372.450 119.700 ;
        RECT 363.450 41.700 372.450 117.300 ;
        RECT 0.600 39.300 372.450 41.700 ;
        RECT 363.450 0.300 372.450 39.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.450 314.700 -0.450 353.700 ;
        RECT 358.950 314.700 361.050 316.050 ;
        RECT -9.450 312.300 362.400 314.700 ;
        RECT -9.450 236.700 -0.450 312.300 ;
        RECT 70.950 310.950 73.050 312.300 ;
        RECT 272.550 310.050 273.450 312.300 ;
        RECT 268.950 308.550 273.450 310.050 ;
        RECT 268.950 307.950 273.000 308.550 ;
        RECT 277.950 246.450 280.050 247.050 ;
        RECT 286.950 246.450 289.050 247.050 ;
        RECT 277.950 245.550 289.050 246.450 ;
        RECT 277.950 244.950 280.050 245.550 ;
        RECT 286.950 244.950 289.050 245.550 ;
        RECT -9.450 234.300 362.400 236.700 ;
        RECT -9.450 158.700 -0.450 234.300 ;
        RECT 28.950 232.950 31.050 234.300 ;
        RECT 127.950 232.950 130.050 234.300 ;
        RECT 187.950 232.950 190.050 234.300 ;
        RECT 229.950 232.950 232.050 234.300 ;
        RECT 310.950 232.950 313.050 234.300 ;
        RECT -9.450 156.300 362.400 158.700 ;
        RECT -9.450 80.700 -0.450 156.300 ;
        RECT 100.950 154.950 103.050 156.300 ;
        RECT 151.950 154.950 154.050 156.300 ;
        RECT 172.950 154.950 175.050 156.300 ;
        RECT 205.950 154.950 208.050 156.300 ;
        RECT 244.950 154.950 247.050 156.300 ;
        RECT 358.950 154.950 361.050 156.300 ;
        RECT -9.450 78.300 362.400 80.700 ;
        RECT -9.450 2.700 -0.450 78.300 ;
        RECT 133.950 76.950 136.050 78.300 ;
        RECT 253.950 76.950 256.050 78.300 ;
        RECT 358.950 76.950 361.050 78.300 ;
        RECT 134.550 73.050 135.450 76.950 ;
        RECT 133.950 70.950 136.050 73.050 ;
        RECT 133.950 61.950 136.050 64.050 ;
        RECT 134.550 45.900 135.450 61.950 ;
        RECT 133.950 43.800 136.050 45.900 ;
        RECT 82.950 2.700 85.500 4.050 ;
        RECT 232.950 2.700 235.500 4.050 ;
        RECT 328.950 2.700 331.500 4.050 ;
        RECT -9.450 0.300 362.400 2.700 ;
      LAYER metal2 ;
        RECT 280.950 349.950 283.050 352.050 ;
        RECT 358.950 349.950 361.050 352.050 ;
        RECT 281.400 336.600 282.450 349.950 ;
        RECT 11.400 336.450 12.600 336.600 ;
        RECT 80.400 336.450 81.600 336.600 ;
        RECT 11.400 335.400 15.450 336.450 ;
        RECT 11.400 334.350 12.600 335.400 ;
        RECT 14.400 313.050 15.450 335.400 ;
        RECT 80.400 335.400 84.450 336.450 ;
        RECT 80.400 334.350 81.600 335.400 ;
        RECT 83.400 319.050 84.450 335.400 ;
        RECT 281.400 334.350 282.600 336.600 ;
        RECT 67.950 316.950 70.050 319.050 ;
        RECT 82.950 316.950 85.050 319.050 ;
        RECT 68.400 313.050 69.450 316.950 ;
        RECT 359.400 316.050 360.450 349.950 ;
        RECT 358.950 313.950 361.050 316.050 ;
        RECT 13.950 310.950 16.050 313.050 ;
        RECT 67.950 310.950 73.050 313.050 ;
        RECT 11.400 291.450 12.600 292.650 ;
        RECT 14.400 291.450 15.450 310.950 ;
        RECT 265.950 307.950 271.050 310.050 ;
        RECT 295.950 307.950 298.050 310.050 ;
        RECT 11.400 290.400 15.450 291.450 ;
        RECT 293.400 291.450 294.600 292.650 ;
        RECT 296.400 291.450 297.450 307.950 ;
        RECT 293.400 290.400 297.450 291.450 ;
        RECT 296.400 276.450 297.450 290.400 ;
        RECT 296.400 275.400 300.450 276.450 ;
        RECT 127.950 260.100 130.050 262.200 ;
        RECT 299.400 261.600 300.450 275.400 ;
        RECT 128.400 259.350 129.600 260.100 ;
        RECT 299.400 259.350 300.600 261.600 ;
        RECT 26.400 258.450 27.600 258.600 ;
        RECT 26.400 257.400 30.450 258.450 ;
        RECT 26.400 256.350 27.600 257.400 ;
        RECT 29.400 235.050 30.450 257.400 ;
        RECT 155.400 254.400 156.600 256.650 ;
        RECT 233.400 254.400 234.600 256.650 ;
        RECT 272.400 254.400 273.600 256.650 ;
        RECT 278.400 254.400 279.600 256.650 ;
        RECT 302.400 254.400 303.600 256.650 ;
        RECT 127.950 250.950 130.050 253.050 ;
        RECT 128.400 235.050 129.450 250.950 ;
        RECT 155.400 237.450 156.450 254.400 ;
        RECT 233.400 238.050 234.450 254.400 ;
        RECT 272.400 243.450 273.450 254.400 ;
        RECT 278.400 247.050 279.450 254.400 ;
        RECT 277.950 244.950 280.050 247.050 ;
        RECT 286.950 244.950 289.050 247.050 ;
        RECT 269.400 242.400 273.450 243.450 ;
        RECT 269.400 238.050 270.450 242.400 ;
        RECT 287.400 241.050 288.450 244.950 ;
        RECT 302.400 241.050 303.450 254.400 ;
        RECT 286.950 238.950 289.050 241.050 ;
        RECT 301.950 238.950 304.050 241.050 ;
        RECT 310.950 238.950 313.050 241.050 ;
        RECT 155.400 236.400 159.450 237.450 ;
        RECT 28.950 232.950 31.050 235.050 ;
        RECT 127.950 232.950 130.050 235.050 ;
        RECT 158.400 226.050 159.450 236.400 ;
        RECT 232.950 235.050 235.050 238.050 ;
        RECT 268.950 235.950 271.050 238.050 ;
        RECT 311.400 235.050 312.450 238.950 ;
        RECT 187.950 232.950 190.050 235.050 ;
        RECT 229.950 234.000 235.050 235.050 ;
        RECT 229.950 233.400 234.450 234.000 ;
        RECT 229.950 232.950 234.000 233.400 ;
        RECT 310.950 232.950 313.050 235.050 ;
        RECT 188.400 226.050 189.450 232.950 ;
        RECT 157.950 223.950 160.050 226.050 ;
        RECT 166.950 223.950 169.050 226.050 ;
        RECT 187.950 223.950 190.050 226.050 ;
        RECT 167.400 220.200 168.450 223.950 ;
        RECT 166.950 218.100 169.050 220.200 ;
        RECT 161.400 210.900 162.600 211.650 ;
        RECT 160.950 208.800 163.050 210.900 ;
        RECT 154.950 182.100 157.050 184.200 ;
        RECT 155.400 181.350 156.600 182.100 ;
        RECT 10.950 179.100 13.050 181.200 ;
        RECT 11.400 178.350 12.600 179.100 ;
        RECT 25.800 178.950 27.900 181.050 ;
        RECT 203.400 180.450 204.600 180.600 ;
        RECT 203.400 179.400 207.450 180.450 ;
        RECT 26.400 172.050 27.450 178.950 ;
        RECT 170.400 176.400 171.600 178.650 ;
        RECT 191.400 176.400 192.600 178.650 ;
        RECT 203.400 178.350 204.600 179.400 ;
        RECT 25.950 169.950 28.050 172.050 ;
        RECT 61.950 169.950 64.050 172.050 ;
        RECT 151.950 169.950 154.050 172.050 ;
        RECT 62.400 163.050 63.450 169.950 ;
        RECT 61.950 160.950 64.050 163.050 ;
        RECT 100.950 160.950 103.050 163.050 ;
        RECT 62.400 142.050 63.450 160.950 ;
        RECT 101.400 157.050 102.450 160.950 ;
        RECT 152.400 157.050 153.450 169.950 ;
        RECT 170.400 157.050 171.450 176.400 ;
        RECT 191.400 163.050 192.450 176.400 ;
        RECT 206.400 163.050 207.450 179.400 ;
        RECT 190.950 160.950 193.050 163.050 ;
        RECT 205.950 160.950 208.050 163.050 ;
        RECT 206.400 157.050 207.450 160.950 ;
        RECT 100.950 154.950 103.050 157.050 ;
        RECT 151.950 154.950 154.050 157.050 ;
        RECT 170.400 155.400 175.050 157.050 ;
        RECT 171.000 154.950 175.050 155.400 ;
        RECT 205.950 154.950 208.050 157.050 ;
        RECT 244.950 156.450 249.000 157.050 ;
        RECT 244.950 154.950 249.450 156.450 ;
        RECT 358.950 154.950 361.050 157.050 ;
        RECT 61.950 139.950 64.050 142.050 ;
        RECT 248.400 138.600 249.450 154.950 ;
        RECT 11.400 135.900 12.600 136.650 ;
        RECT 248.400 136.350 249.600 138.600 ;
        RECT 10.950 133.800 13.050 135.900 ;
        RECT 299.400 134.400 300.600 136.650 ;
        RECT 251.400 132.900 252.600 133.650 ;
        RECT 250.950 130.800 253.050 132.900 ;
        RECT 268.950 127.650 271.050 129.750 ;
        RECT 115.950 101.100 118.050 103.200 ;
        RECT 269.400 103.050 270.450 127.650 ;
        RECT 299.400 127.050 300.450 134.400 ;
        RECT 359.400 132.450 360.450 154.950 ;
        RECT 356.400 131.400 360.450 132.450 ;
        RECT 356.400 127.050 357.450 131.400 ;
        RECT 298.950 124.950 301.050 127.050 ;
        RECT 355.950 124.950 358.050 127.050 ;
        RECT 116.400 100.350 117.600 101.100 ;
        RECT 130.800 100.950 132.900 103.050 ;
        RECT 268.950 100.950 271.050 103.050 ;
        RECT 271.950 101.100 274.050 103.200 ;
        RECT 131.400 93.450 132.450 100.950 ;
        RECT 212.400 98.400 213.600 100.650 ;
        RECT 272.400 100.350 273.600 101.100 ;
        RECT 131.400 92.400 135.450 93.450 ;
        RECT 134.400 79.050 135.450 92.400 ;
        RECT 212.400 82.050 213.450 98.400 ;
        RECT 256.950 94.950 259.050 97.050 ;
        RECT 211.950 79.950 214.050 82.050 ;
        RECT 253.950 81.450 256.050 82.050 ;
        RECT 257.400 81.450 258.450 94.950 ;
        RECT 253.950 80.400 258.450 81.450 ;
        RECT 133.950 76.950 136.050 79.050 ;
        RECT 253.950 76.950 256.050 80.400 ;
        RECT 358.950 76.950 361.050 79.050 ;
        RECT 133.950 70.950 136.050 73.050 ;
        RECT 134.400 64.050 135.450 70.950 ;
        RECT 133.950 61.950 136.050 64.050 ;
        RECT 41.400 56.400 42.600 58.650 ;
        RECT 293.400 56.400 294.600 58.650 ;
        RECT 41.400 40.050 42.450 56.400 ;
        RECT 173.400 53.400 174.600 55.650 ;
        RECT 173.400 46.050 174.450 53.400 ;
        RECT 293.400 52.050 294.450 56.400 ;
        RECT 359.400 52.050 360.450 76.950 ;
        RECT 292.950 49.950 295.050 52.050 ;
        RECT 358.950 49.950 361.050 52.050 ;
        RECT 135.000 45.900 138.000 46.050 ;
        RECT 133.950 43.950 139.050 45.900 ;
        RECT 172.950 43.950 175.050 46.050 ;
        RECT 133.950 43.800 136.050 43.950 ;
        RECT 136.950 43.800 139.050 43.950 ;
        RECT 40.950 37.950 43.050 40.050 ;
        RECT 70.950 34.950 73.050 37.050 ;
        RECT 22.800 23.100 24.900 25.200 ;
        RECT 23.400 22.350 24.600 23.100 ;
        RECT 25.950 19.800 28.050 21.900 ;
        RECT 26.400 4.050 27.450 19.800 ;
        RECT 71.400 4.050 72.450 34.950 ;
        RECT 268.950 23.100 271.050 25.200 ;
        RECT 227.400 21.900 228.600 22.650 ;
        RECT 269.400 22.350 270.600 23.100 ;
        RECT 328.950 22.950 331.050 25.050 ;
        RECT 226.950 19.800 229.050 21.900 ;
        RECT 232.950 16.950 235.050 19.050 ;
        RECT 233.400 4.050 234.450 16.950 ;
        RECT 329.400 4.050 330.450 22.950 ;
        RECT 25.950 1.950 28.050 4.050 ;
        RECT 70.950 1.950 73.050 4.050 ;
        RECT 79.950 1.950 85.050 4.050 ;
        RECT 232.950 1.950 235.050 4.050 ;
        RECT 328.950 1.950 331.050 4.050 ;
      LAYER metal3 ;
        RECT 280.950 351.600 283.050 352.050 ;
        RECT 358.950 351.600 361.050 352.050 ;
        RECT 280.950 350.400 361.050 351.600 ;
        RECT 280.950 349.950 283.050 350.400 ;
        RECT 358.950 349.950 361.050 350.400 ;
        RECT 67.950 318.600 70.050 319.050 ;
        RECT 82.950 318.600 85.050 319.050 ;
        RECT 67.950 317.400 85.050 318.600 ;
        RECT 67.950 316.950 70.050 317.400 ;
        RECT 82.950 316.950 85.050 317.400 ;
        RECT 13.950 312.600 16.050 313.050 ;
        RECT 67.950 312.600 70.050 313.050 ;
        RECT 13.950 311.400 70.050 312.600 ;
        RECT 13.950 310.950 16.050 311.400 ;
        RECT 67.950 310.950 70.050 311.400 ;
        RECT 265.950 309.600 268.050 310.050 ;
        RECT 295.950 309.600 298.050 310.050 ;
        RECT 265.950 308.400 298.050 309.600 ;
        RECT 265.950 307.950 268.050 308.400 ;
        RECT 295.950 307.950 298.050 308.400 ;
        RECT 127.950 261.600 130.050 262.200 ;
        RECT 125.400 260.400 130.050 261.600 ;
        RECT 125.400 253.050 126.600 260.400 ;
        RECT 127.950 260.100 130.050 260.400 ;
        RECT 125.400 251.400 130.050 253.050 ;
        RECT 126.000 250.950 130.050 251.400 ;
        RECT 286.950 240.600 289.050 241.050 ;
        RECT 301.950 240.600 304.050 241.050 ;
        RECT 310.950 240.600 313.050 241.050 ;
        RECT 286.950 239.400 313.050 240.600 ;
        RECT 286.950 238.950 289.050 239.400 ;
        RECT 301.950 238.950 304.050 239.400 ;
        RECT 310.950 238.950 313.050 239.400 ;
        RECT 232.950 237.600 235.050 238.050 ;
        RECT 268.950 237.600 271.050 238.050 ;
        RECT 232.950 236.400 271.050 237.600 ;
        RECT 232.950 235.950 235.050 236.400 ;
        RECT 268.950 235.950 271.050 236.400 ;
        RECT 157.950 225.600 160.050 226.050 ;
        RECT 166.950 225.600 169.050 226.050 ;
        RECT 187.950 225.600 190.050 226.050 ;
        RECT 157.950 224.400 190.050 225.600 ;
        RECT 157.950 223.950 160.050 224.400 ;
        RECT 166.950 223.950 169.050 224.400 ;
        RECT 187.950 223.950 190.050 224.400 ;
        RECT 166.950 220.050 169.050 220.200 ;
        RECT 165.000 219.600 169.050 220.050 ;
        RECT 164.400 218.100 169.050 219.600 ;
        RECT 164.400 217.950 168.000 218.100 ;
        RECT 160.950 210.600 163.050 210.900 ;
        RECT 164.400 210.600 165.600 217.950 ;
        RECT 160.950 209.400 165.600 210.600 ;
        RECT 160.950 208.800 163.050 209.400 ;
        RECT 154.950 182.100 157.050 184.200 ;
        RECT 10.950 180.600 13.050 181.200 ;
        RECT 25.800 180.600 27.900 181.050 ;
        RECT 155.400 180.600 156.600 182.100 ;
        RECT 10.950 179.400 27.900 180.600 ;
        RECT 10.950 179.100 13.050 179.400 ;
        RECT 25.800 178.950 27.900 179.400 ;
        RECT 152.400 179.400 156.600 180.600 ;
        RECT 152.400 172.050 153.600 179.400 ;
        RECT 25.950 171.600 28.050 172.050 ;
        RECT 61.950 171.600 64.050 172.050 ;
        RECT 25.950 170.400 64.050 171.600 ;
        RECT 25.950 169.950 28.050 170.400 ;
        RECT 61.950 169.950 64.050 170.400 ;
        RECT 151.950 169.950 154.050 172.050 ;
        RECT 61.950 162.600 64.050 163.050 ;
        RECT 100.950 162.600 103.050 163.050 ;
        RECT 61.950 161.400 103.050 162.600 ;
        RECT 61.950 160.950 64.050 161.400 ;
        RECT 100.950 160.950 103.050 161.400 ;
        RECT 190.950 162.600 193.050 163.050 ;
        RECT 205.950 162.600 208.050 163.050 ;
        RECT 190.950 161.400 208.050 162.600 ;
        RECT 190.950 160.950 193.050 161.400 ;
        RECT 205.950 160.950 208.050 161.400 ;
        RECT 61.950 141.600 64.050 142.050 ;
        RECT 23.400 140.400 64.050 141.600 ;
        RECT 23.400 138.600 24.600 140.400 ;
        RECT 61.950 139.950 64.050 140.400 ;
        RECT 20.400 137.400 24.600 138.600 ;
        RECT 10.950 135.600 13.050 135.900 ;
        RECT 20.400 135.600 21.600 137.400 ;
        RECT 10.950 134.400 21.600 135.600 ;
        RECT 10.950 133.800 13.050 134.400 ;
        RECT 250.950 132.600 253.050 132.900 ;
        RECT 250.950 131.400 255.600 132.600 ;
        RECT 250.950 130.800 253.050 131.400 ;
        RECT 254.400 129.600 255.600 131.400 ;
        RECT 268.950 129.600 271.050 129.750 ;
        RECT 254.400 128.400 271.050 129.600 ;
        RECT 268.950 127.650 271.050 128.400 ;
        RECT 298.950 126.600 301.050 127.050 ;
        RECT 355.950 126.600 358.050 127.050 ;
        RECT 298.950 125.400 358.050 126.600 ;
        RECT 298.950 124.950 301.050 125.400 ;
        RECT 355.950 124.950 358.050 125.400 ;
        RECT 115.950 102.600 118.050 103.200 ;
        RECT 130.800 102.600 132.900 103.050 ;
        RECT 268.950 102.600 271.050 103.050 ;
        RECT 271.950 102.600 274.050 103.200 ;
        RECT 115.950 101.400 132.900 102.600 ;
        RECT 115.950 101.100 118.050 101.400 ;
        RECT 130.800 100.950 132.900 101.400 ;
        RECT 257.400 101.400 274.050 102.600 ;
        RECT 257.400 97.050 258.600 101.400 ;
        RECT 268.950 100.950 271.050 101.400 ;
        RECT 271.950 101.100 274.050 101.400 ;
        RECT 256.950 94.950 259.050 97.050 ;
        RECT 211.950 81.600 214.050 82.050 ;
        RECT 253.950 81.600 256.050 82.050 ;
        RECT 211.950 80.400 256.050 81.600 ;
        RECT 211.950 79.950 214.050 80.400 ;
        RECT 253.950 79.950 256.050 80.400 ;
        RECT 292.950 51.600 295.050 52.050 ;
        RECT 358.950 51.600 361.050 52.050 ;
        RECT 292.950 50.400 361.050 51.600 ;
        RECT 292.950 49.950 295.050 50.400 ;
        RECT 358.950 49.950 361.050 50.400 ;
        RECT 136.950 45.600 139.050 45.900 ;
        RECT 172.950 45.600 175.050 46.050 ;
        RECT 136.950 44.400 175.050 45.600 ;
        RECT 136.950 43.800 139.050 44.400 ;
        RECT 172.950 43.950 175.050 44.400 ;
        RECT 40.950 39.600 43.050 40.050 ;
        RECT 40.950 38.400 69.600 39.600 ;
        RECT 40.950 37.950 43.050 38.400 ;
        RECT 68.400 37.050 69.600 38.400 ;
        RECT 68.400 35.400 73.050 37.050 ;
        RECT 69.000 34.950 73.050 35.400 ;
        RECT 22.800 23.100 24.900 25.200 ;
        RECT 268.950 24.600 271.050 25.200 ;
        RECT 328.950 24.600 331.050 25.050 ;
        RECT 268.950 23.400 331.050 24.600 ;
        RECT 268.950 23.100 271.050 23.400 ;
        RECT 23.400 22.050 24.600 23.100 ;
        RECT 328.950 22.950 331.050 23.400 ;
        RECT 23.400 21.900 27.000 22.050 ;
        RECT 23.400 20.400 28.050 21.900 ;
        RECT 24.000 19.950 28.050 20.400 ;
        RECT 25.950 19.800 28.050 19.950 ;
        RECT 226.950 21.600 229.050 21.900 ;
        RECT 226.950 20.400 231.600 21.600 ;
        RECT 226.950 19.800 229.050 20.400 ;
        RECT 230.400 19.050 231.600 20.400 ;
        RECT 230.400 17.400 235.050 19.050 ;
        RECT 231.000 16.950 235.050 17.400 ;
        RECT 25.950 3.600 28.050 4.050 ;
        RECT 70.950 3.600 73.050 4.050 ;
        RECT 79.950 3.600 82.050 4.050 ;
        RECT 25.950 2.400 82.050 3.600 ;
        RECT 25.950 1.950 28.050 2.400 ;
        RECT 70.950 1.950 73.050 2.400 ;
        RECT 79.950 1.950 82.050 2.400 ;
    END
  END vdd
  PIN CLK
    PORT
      LAYER metal2 ;
        RECT 55.950 340.950 58.050 343.050 ;
        RECT 124.950 340.950 127.050 343.050 ;
        RECT 56.400 337.200 57.450 340.950 ;
        RECT 49.950 335.100 52.050 337.200 ;
        RECT 55.950 335.100 58.050 337.200 ;
        RECT 125.400 336.600 126.450 340.950 ;
        RECT 50.400 286.050 51.450 335.100 ;
        RECT 56.400 334.350 57.600 335.100 ;
        RECT 125.400 334.350 126.600 336.600 ;
        RECT 323.400 336.450 324.450 360.450 ;
        RECT 325.950 336.450 328.050 337.200 ;
        RECT 323.400 335.400 328.050 336.450 ;
        RECT 325.950 335.100 328.050 335.400 ;
        RECT 340.950 335.100 343.050 337.200 ;
        RECT 326.400 334.350 327.600 335.100 ;
        RECT 56.400 290.400 57.600 292.650 ;
        RECT 338.400 291.450 339.600 292.650 ;
        RECT 341.400 291.450 342.450 335.100 ;
        RECT 338.400 290.400 342.450 291.450 ;
        RECT 56.400 286.050 57.450 290.400 ;
        RECT 49.950 283.950 52.050 286.050 ;
        RECT 55.950 283.950 58.050 286.050 ;
        RECT 64.950 283.950 67.050 286.050 ;
        RECT 65.400 259.200 66.450 283.950 ;
        RECT 338.400 280.050 339.450 290.400 ;
        RECT 337.950 277.950 340.050 280.050 ;
        RECT 301.950 274.950 304.050 277.050 ;
        RECT 302.400 265.050 303.450 274.950 ;
        RECT 301.950 262.950 304.050 265.050 ;
        RECT 64.950 257.100 67.050 259.200 ;
        RECT 70.950 257.100 73.050 259.200 ;
        RECT 65.400 220.050 66.450 257.100 ;
        RECT 71.400 256.350 72.600 257.100 ;
        RECT 316.950 250.950 319.050 253.050 ;
        RECT 317.400 238.050 318.450 250.950 ;
        RECT 316.950 235.950 319.050 238.050 ;
        RECT 334.950 235.950 337.050 238.050 ;
        RECT 64.950 217.950 67.050 220.050 ;
        RECT 335.400 217.050 336.450 235.950 ;
        RECT 334.950 214.950 337.050 217.050 ;
        RECT 337.950 208.950 340.050 211.050 ;
        RECT 70.950 199.950 73.050 202.050 ;
        RECT 71.400 192.450 72.450 199.950 ;
        RECT 65.400 191.400 72.450 192.450 ;
        RECT 65.400 183.450 66.450 191.400 ;
        RECT 62.400 183.000 66.450 183.450 ;
        RECT 61.950 182.400 66.450 183.000 ;
        RECT 61.950 181.200 64.050 182.400 ;
        RECT 55.950 179.100 58.050 181.200 ;
        RECT 61.800 180.000 64.050 181.200 ;
        RECT 61.800 179.100 63.900 180.000 ;
        RECT 56.400 178.350 57.600 179.100 ;
        RECT 71.400 157.050 72.450 191.400 ;
        RECT 248.400 180.450 249.600 180.600 ;
        RECT 248.400 179.400 252.450 180.450 ;
        RECT 248.400 178.350 249.600 179.400 ;
        RECT 251.400 178.050 252.450 179.400 ;
        RECT 250.950 175.950 253.050 178.050 ;
        RECT 193.950 172.950 196.050 175.050 ;
        RECT 251.400 174.450 252.450 175.950 ;
        RECT 251.400 173.400 255.450 174.450 ;
        RECT 58.950 154.950 61.050 157.050 ;
        RECT 70.950 154.950 73.050 157.050 ;
        RECT 56.400 135.450 57.600 136.650 ;
        RECT 59.400 135.450 60.450 154.950 ;
        RECT 194.400 142.050 195.450 172.950 ;
        RECT 254.400 151.050 255.450 173.400 ;
        RECT 253.950 148.950 256.050 151.050 ;
        RECT 338.400 148.050 339.450 208.950 ;
        RECT 337.950 145.950 340.050 148.050 ;
        RECT 193.950 139.950 196.050 142.050 ;
        RECT 338.400 136.050 339.450 145.950 ;
        RECT 56.400 134.400 60.450 135.450 ;
        RECT 56.400 106.050 57.450 134.400 ;
        RECT 337.950 133.950 340.050 136.050 ;
        RECT 344.400 135.900 345.600 136.650 ;
        RECT 343.950 133.800 346.050 135.900 ;
        RECT 172.950 130.950 175.050 133.050 ;
        RECT 173.400 124.050 174.450 130.950 ;
        RECT 160.950 121.950 163.050 124.050 ;
        RECT 172.950 121.950 175.050 124.050 ;
        RECT 55.950 103.950 58.050 106.050 ;
        RECT 161.400 102.600 162.450 121.950 ;
        RECT 344.400 109.050 345.450 133.800 ;
        RECT 316.950 106.950 319.050 109.050 ;
        RECT 331.950 106.950 334.050 109.050 ;
        RECT 343.950 106.950 346.050 109.050 ;
        RECT 317.400 102.600 318.450 106.950 ;
        RECT 161.400 100.350 162.600 102.600 ;
        RECT 317.400 100.350 318.600 102.600 ;
        RECT 43.950 94.950 46.050 97.050 ;
        RECT 44.400 55.050 45.450 94.950 ;
        RECT 86.400 56.400 87.600 58.650 ;
        RECT 86.400 55.050 87.450 56.400 ;
        RECT 332.400 55.050 333.450 106.950 ;
        RECT 338.400 57.000 339.600 58.650 ;
        RECT 43.950 52.950 46.050 55.050 ;
        RECT 85.950 52.950 88.050 55.050 ;
        RECT 331.950 52.950 334.050 55.050 ;
        RECT 337.950 52.950 340.050 57.000 ;
        RECT 86.400 43.050 87.450 52.950 ;
        RECT 67.950 40.950 70.050 43.050 ;
        RECT 85.950 40.950 88.050 43.050 ;
        RECT 68.400 24.600 69.450 40.950 ;
        RECT 68.400 22.350 69.600 24.600 ;
        RECT 86.400 13.050 87.450 40.950 ;
        RECT 332.400 40.050 333.450 52.950 ;
        RECT 307.950 37.950 310.050 40.050 ;
        RECT 313.950 37.950 316.050 40.050 ;
        RECT 331.950 37.950 334.050 40.050 ;
        RECT 85.950 10.950 88.050 13.050 ;
        RECT 308.400 10.050 309.450 37.950 ;
        RECT 314.400 24.600 315.450 37.950 ;
        RECT 314.400 22.350 315.600 24.600 ;
        RECT 307.950 7.950 310.050 10.050 ;
      LAYER metal3 ;
        RECT 55.950 342.600 58.050 343.050 ;
        RECT 124.950 342.600 127.050 343.050 ;
        RECT 55.950 341.400 127.050 342.600 ;
        RECT 55.950 340.950 58.050 341.400 ;
        RECT 124.950 340.950 127.050 341.400 ;
        RECT 49.950 336.750 52.050 337.200 ;
        RECT 55.950 336.750 58.050 337.200 ;
        RECT 49.950 335.550 58.050 336.750 ;
        RECT 49.950 335.100 52.050 335.550 ;
        RECT 55.950 335.100 58.050 335.550 ;
        RECT 325.950 336.750 328.050 337.200 ;
        RECT 340.950 336.750 343.050 337.200 ;
        RECT 325.950 335.550 343.050 336.750 ;
        RECT 325.950 335.100 328.050 335.550 ;
        RECT 340.950 335.100 343.050 335.550 ;
        RECT 49.950 285.600 52.050 286.050 ;
        RECT 55.950 285.600 58.050 286.050 ;
        RECT 64.950 285.600 67.050 286.050 ;
        RECT 49.950 284.400 67.050 285.600 ;
        RECT 49.950 283.950 52.050 284.400 ;
        RECT 55.950 283.950 58.050 284.400 ;
        RECT 64.950 283.950 67.050 284.400 ;
        RECT 301.950 276.600 304.050 277.050 ;
        RECT 337.950 276.600 340.050 280.050 ;
        RECT 301.950 276.000 340.050 276.600 ;
        RECT 301.950 275.400 339.600 276.000 ;
        RECT 301.950 274.950 304.050 275.400 ;
        RECT 300.000 264.600 304.050 265.050 ;
        RECT 299.400 262.950 304.050 264.600 ;
        RECT 64.950 258.750 67.050 259.200 ;
        RECT 70.950 258.750 73.050 259.200 ;
        RECT 64.950 257.550 73.050 258.750 ;
        RECT 64.950 257.100 67.050 257.550 ;
        RECT 70.950 257.100 73.050 257.550 ;
        RECT 299.400 252.600 300.600 262.950 ;
        RECT 316.950 252.600 319.050 253.050 ;
        RECT 299.400 251.400 319.050 252.600 ;
        RECT 316.950 250.950 319.050 251.400 ;
        RECT 316.950 237.600 319.050 238.050 ;
        RECT 334.950 237.600 337.050 238.050 ;
        RECT 316.950 236.400 337.050 237.600 ;
        RECT 316.950 235.950 319.050 236.400 ;
        RECT 334.950 235.950 337.050 236.400 ;
        RECT 64.950 219.600 67.050 220.050 ;
        RECT 64.950 218.400 72.600 219.600 ;
        RECT 64.950 217.950 67.050 218.400 ;
        RECT 71.400 213.600 72.600 218.400 ;
        RECT 334.950 214.950 337.050 217.050 ;
        RECT 68.400 212.400 72.600 213.600 ;
        RECT 68.400 202.050 69.600 212.400 ;
        RECT 335.400 211.050 336.600 214.950 ;
        RECT 335.400 209.400 340.050 211.050 ;
        RECT 336.000 208.950 340.050 209.400 ;
        RECT 68.400 200.400 73.050 202.050 ;
        RECT 69.000 199.950 73.050 200.400 ;
        RECT 55.950 180.750 58.050 181.200 ;
        RECT 61.800 180.750 63.900 181.200 ;
        RECT 55.950 179.550 63.900 180.750 ;
        RECT 55.950 179.100 58.050 179.550 ;
        RECT 61.800 179.100 63.900 179.550 ;
        RECT 250.950 177.600 253.050 178.050 ;
        RECT 194.400 177.000 253.050 177.600 ;
        RECT 193.950 176.400 253.050 177.000 ;
        RECT 193.950 172.950 196.050 176.400 ;
        RECT 250.950 175.950 253.050 176.400 ;
        RECT 58.950 156.600 61.050 157.050 ;
        RECT 70.950 156.600 73.050 157.050 ;
        RECT 58.950 155.400 73.050 156.600 ;
        RECT 58.950 154.950 61.050 155.400 ;
        RECT 70.950 154.950 73.050 155.400 ;
        RECT 253.950 150.600 256.050 151.050 ;
        RECT 253.950 149.400 285.600 150.600 ;
        RECT 253.950 148.950 256.050 149.400 ;
        RECT 284.400 147.600 285.600 149.400 ;
        RECT 337.950 147.600 340.050 148.050 ;
        RECT 284.400 146.400 340.050 147.600 ;
        RECT 337.950 145.950 340.050 146.400 ;
        RECT 193.950 139.950 196.050 142.050 ;
        RECT 194.400 135.600 195.600 139.950 ;
        RECT 182.400 134.400 195.600 135.600 ;
        RECT 337.950 135.600 340.050 136.050 ;
        RECT 343.950 135.600 346.050 135.900 ;
        RECT 337.950 134.400 346.050 135.600 ;
        RECT 172.950 132.600 175.050 133.050 ;
        RECT 182.400 132.600 183.600 134.400 ;
        RECT 337.950 133.950 340.050 134.400 ;
        RECT 343.950 133.800 346.050 134.400 ;
        RECT 172.950 131.400 183.600 132.600 ;
        RECT 172.950 130.950 175.050 131.400 ;
        RECT 160.950 123.600 163.050 124.050 ;
        RECT 172.950 123.600 175.050 124.050 ;
        RECT 160.950 122.400 175.050 123.600 ;
        RECT 160.950 121.950 163.050 122.400 ;
        RECT 172.950 121.950 175.050 122.400 ;
        RECT 316.950 108.600 319.050 109.050 ;
        RECT 331.950 108.600 334.050 109.050 ;
        RECT 343.950 108.600 346.050 109.050 ;
        RECT 316.950 107.400 346.050 108.600 ;
        RECT 316.950 106.950 319.050 107.400 ;
        RECT 331.950 106.950 334.050 107.400 ;
        RECT 343.950 106.950 346.050 107.400 ;
        RECT 55.950 103.950 58.050 106.050 ;
        RECT 56.400 99.600 57.600 103.950 ;
        RECT 50.400 98.400 57.600 99.600 ;
        RECT 43.950 96.600 46.050 97.050 ;
        RECT 50.400 96.600 51.600 98.400 ;
        RECT 43.950 95.400 51.600 96.600 ;
        RECT 43.950 94.950 46.050 95.400 ;
        RECT 43.950 54.600 46.050 55.050 ;
        RECT 85.950 54.600 88.050 55.050 ;
        RECT 43.950 53.400 88.050 54.600 ;
        RECT 43.950 52.950 46.050 53.400 ;
        RECT 85.950 52.950 88.050 53.400 ;
        RECT 331.950 54.600 334.050 55.050 ;
        RECT 337.950 54.600 340.050 55.050 ;
        RECT 331.950 53.400 340.050 54.600 ;
        RECT 331.950 52.950 334.050 53.400 ;
        RECT 337.950 52.950 340.050 53.400 ;
        RECT 67.950 42.600 70.050 43.050 ;
        RECT 85.950 42.600 88.050 43.050 ;
        RECT 67.950 41.400 88.050 42.600 ;
        RECT 67.950 40.950 70.050 41.400 ;
        RECT 85.950 40.950 88.050 41.400 ;
        RECT 307.950 39.600 310.050 40.050 ;
        RECT 313.950 39.600 316.050 40.050 ;
        RECT 331.950 39.600 334.050 40.050 ;
        RECT 307.950 38.400 334.050 39.600 ;
        RECT 307.950 37.950 310.050 38.400 ;
        RECT 313.950 37.950 316.050 38.400 ;
        RECT 331.950 37.950 334.050 38.400 ;
        RECT 85.950 12.600 90.000 13.050 ;
        RECT 85.950 10.950 90.600 12.600 ;
        RECT 89.400 9.600 90.600 10.950 ;
        RECT 307.950 9.600 310.050 10.050 ;
        RECT 89.400 8.400 310.050 9.600 ;
        RECT 307.950 7.950 310.050 8.400 ;
    END
  END CLK
  PIN Din[3]
    PORT
      LAYER metal2 ;
        RECT 221.400 346.050 222.450 360.450 ;
        RECT 187.950 343.950 190.050 346.050 ;
        RECT 220.950 343.950 223.050 346.050 ;
        RECT 188.400 325.050 189.450 343.950 ;
        RECT 187.950 322.950 190.050 325.050 ;
        RECT 220.950 322.950 223.050 325.050 ;
        RECT 221.400 295.200 222.450 322.950 ;
        RECT 220.950 293.100 223.050 295.200 ;
        RECT 221.400 292.350 222.600 293.100 ;
        RECT 223.950 286.950 226.050 289.050 ;
        RECT 224.400 274.050 225.450 286.950 ;
        RECT 208.950 271.950 211.050 274.050 ;
        RECT 223.950 271.950 226.050 274.050 ;
        RECT 209.400 250.050 210.450 271.950 ;
        RECT 136.950 247.950 139.050 250.050 ;
        RECT 137.400 219.450 138.450 247.950 ;
        RECT 202.950 247.800 205.050 249.900 ;
        RECT 208.950 247.950 211.050 250.050 ;
        RECT 137.400 218.400 141.450 219.450 ;
        RECT 140.400 216.600 141.450 218.400 ;
        RECT 140.400 214.350 141.600 216.600 ;
        RECT 203.400 187.050 204.450 247.800 ;
        RECT 202.800 184.950 204.900 187.050 ;
        RECT 181.950 175.950 184.050 178.050 ;
        RECT 266.400 176.400 267.600 178.650 ;
        RECT 182.400 151.050 183.450 175.950 ;
        RECT 266.400 169.050 267.450 176.400 ;
        RECT 199.950 166.950 202.050 169.050 ;
        RECT 265.950 166.950 268.050 169.050 ;
        RECT 200.400 151.050 201.450 166.950 ;
        RECT 181.950 148.950 184.050 151.050 ;
        RECT 199.950 148.950 202.050 151.050 ;
        RECT 182.400 138.600 183.450 148.950 ;
        RECT 182.400 136.350 183.600 138.600 ;
      LAYER metal3 ;
        RECT 187.950 345.600 190.050 346.050 ;
        RECT 220.950 345.600 223.050 346.050 ;
        RECT 187.950 344.400 223.050 345.600 ;
        RECT 187.950 343.950 190.050 344.400 ;
        RECT 220.950 343.950 223.050 344.400 ;
        RECT 187.950 324.600 190.050 325.050 ;
        RECT 220.950 324.600 223.050 325.050 ;
        RECT 187.950 323.400 223.050 324.600 ;
        RECT 187.950 322.950 190.050 323.400 ;
        RECT 220.950 322.950 223.050 323.400 ;
        RECT 220.950 293.100 223.050 295.200 ;
        RECT 221.400 289.050 222.600 293.100 ;
        RECT 221.400 287.400 226.050 289.050 ;
        RECT 222.000 286.950 226.050 287.400 ;
        RECT 208.950 273.600 211.050 274.050 ;
        RECT 223.950 273.600 226.050 274.050 ;
        RECT 208.950 272.400 226.050 273.600 ;
        RECT 208.950 271.950 211.050 272.400 ;
        RECT 223.950 271.950 226.050 272.400 ;
        RECT 136.950 249.600 139.050 250.050 ;
        RECT 202.950 249.600 205.050 249.900 ;
        RECT 208.950 249.600 211.050 250.050 ;
        RECT 136.950 248.400 211.050 249.600 ;
        RECT 136.950 247.950 139.050 248.400 ;
        RECT 202.950 247.800 205.050 248.400 ;
        RECT 208.950 247.950 211.050 248.400 ;
        RECT 202.800 186.600 204.900 187.050 ;
        RECT 197.400 185.400 204.900 186.600 ;
        RECT 197.400 183.600 198.600 185.400 ;
        RECT 202.800 184.950 204.900 185.400 ;
        RECT 185.400 182.400 198.600 183.600 ;
        RECT 185.400 178.050 186.600 182.400 ;
        RECT 181.950 176.400 186.600 178.050 ;
        RECT 181.950 175.950 186.000 176.400 ;
        RECT 199.950 168.600 202.050 169.050 ;
        RECT 265.950 168.600 268.050 169.050 ;
        RECT 199.950 167.400 268.050 168.600 ;
        RECT 199.950 166.950 202.050 167.400 ;
        RECT 265.950 166.950 268.050 167.400 ;
        RECT 181.950 150.600 184.050 151.050 ;
        RECT 199.950 150.600 202.050 151.050 ;
        RECT 181.950 149.400 202.050 150.600 ;
        RECT 181.950 148.950 184.050 149.400 ;
        RECT 199.950 148.950 202.050 149.400 ;
    END
  END Din[3]
  PIN Din[2]
    PORT
      LAYER metal2 ;
        RECT 110.400 352.050 111.450 360.450 ;
        RECT 109.950 349.950 112.050 352.050 ;
        RECT 127.950 349.950 130.050 352.050 ;
        RECT 128.400 319.050 129.450 349.950 ;
        RECT 103.950 316.950 106.050 319.050 ;
        RECT 127.950 316.950 130.050 319.050 ;
        RECT 104.400 295.050 105.450 316.950 ;
        RECT 103.950 294.600 108.000 295.050 ;
        RECT 103.950 292.950 108.600 294.600 ;
        RECT 107.400 292.350 108.600 292.950 ;
        RECT 100.950 286.950 103.050 289.050 ;
        RECT 101.400 262.050 102.450 286.950 ;
        RECT 100.950 259.950 103.050 262.050 ;
        RECT 100.950 253.950 103.050 256.050 ;
        RECT 101.400 234.450 102.450 253.950 ;
        RECT 98.400 233.400 102.450 234.450 ;
        RECT 98.400 223.050 99.450 233.400 ;
        RECT 79.950 220.950 82.050 223.050 ;
        RECT 97.950 220.950 100.050 223.050 ;
        RECT 80.400 217.050 81.450 220.950 ;
        RECT 79.950 214.950 82.050 217.050 ;
        RECT 79.950 208.950 82.050 211.050 ;
        RECT 80.400 196.050 81.450 208.950 ;
        RECT 58.950 193.950 61.050 196.050 ;
        RECT 79.950 193.950 82.050 196.050 ;
        RECT 59.400 166.050 60.450 193.950 ;
        RECT 131.400 176.400 132.600 178.650 ;
        RECT 131.400 174.450 132.450 176.400 ;
        RECT 131.400 173.400 135.450 174.450 ;
        RECT 134.400 169.050 135.450 173.400 ;
        RECT 133.950 166.950 136.050 169.050 ;
        RECT 178.950 166.950 181.050 169.050 ;
        RECT 58.950 163.950 61.050 166.050 ;
        RECT 112.950 163.950 115.050 166.050 ;
        RECT 113.400 160.050 114.450 163.950 ;
        RECT 134.400 160.050 135.450 166.950 ;
        RECT 179.400 160.050 180.450 166.950 ;
        RECT 112.950 157.950 115.050 160.050 ;
        RECT 133.950 157.950 136.050 160.050 ;
        RECT 178.950 157.950 181.050 160.050 ;
        RECT 214.950 157.950 217.050 160.050 ;
        RECT 215.400 145.050 216.450 157.950 ;
        RECT 214.950 142.950 217.050 145.050 ;
        RECT 235.950 142.950 238.050 145.050 ;
        RECT 215.400 138.600 216.450 142.950 ;
        RECT 236.400 138.600 237.450 142.950 ;
        RECT 215.400 136.350 216.600 138.600 ;
        RECT 236.400 136.350 237.600 138.600 ;
      LAYER metal3 ;
        RECT 109.950 351.600 112.050 352.050 ;
        RECT 127.950 351.600 130.050 352.050 ;
        RECT 109.950 350.400 130.050 351.600 ;
        RECT 109.950 349.950 112.050 350.400 ;
        RECT 127.950 349.950 130.050 350.400 ;
        RECT 103.950 318.600 106.050 319.050 ;
        RECT 127.950 318.600 130.050 319.050 ;
        RECT 103.950 317.400 130.050 318.600 ;
        RECT 103.950 316.950 106.050 317.400 ;
        RECT 127.950 316.950 130.050 317.400 ;
        RECT 103.950 292.950 106.050 295.050 ;
        RECT 104.400 289.050 105.600 292.950 ;
        RECT 100.950 287.400 105.600 289.050 ;
        RECT 100.950 286.950 105.000 287.400 ;
        RECT 100.950 259.950 103.050 262.050 ;
        RECT 101.400 256.050 102.600 259.950 ;
        RECT 100.950 253.950 103.050 256.050 ;
        RECT 79.950 222.600 82.050 223.050 ;
        RECT 97.950 222.600 100.050 223.050 ;
        RECT 79.950 221.400 100.050 222.600 ;
        RECT 79.950 220.950 82.050 221.400 ;
        RECT 97.950 220.950 100.050 221.400 ;
        RECT 79.950 214.950 82.050 217.050 ;
        RECT 80.400 211.050 81.600 214.950 ;
        RECT 79.950 208.950 82.050 211.050 ;
        RECT 58.950 195.600 61.050 196.050 ;
        RECT 79.950 195.600 82.050 196.050 ;
        RECT 58.950 194.400 82.050 195.600 ;
        RECT 58.950 193.950 61.050 194.400 ;
        RECT 79.950 193.950 82.050 194.400 ;
        RECT 133.950 168.600 136.050 169.050 ;
        RECT 178.950 168.600 181.050 169.050 ;
        RECT 133.950 167.400 181.050 168.600 ;
        RECT 133.950 166.950 136.050 167.400 ;
        RECT 178.950 166.950 181.050 167.400 ;
        RECT 58.950 165.600 61.050 166.050 ;
        RECT 112.950 165.600 115.050 166.050 ;
        RECT 58.950 164.400 115.050 165.600 ;
        RECT 58.950 163.950 61.050 164.400 ;
        RECT 112.950 163.950 115.050 164.400 ;
        RECT 112.950 159.600 115.050 160.050 ;
        RECT 133.950 159.600 136.050 160.050 ;
        RECT 112.950 158.400 136.050 159.600 ;
        RECT 112.950 157.950 115.050 158.400 ;
        RECT 133.950 157.950 136.050 158.400 ;
        RECT 178.950 159.600 181.050 160.050 ;
        RECT 214.950 159.600 217.050 160.050 ;
        RECT 178.950 158.400 217.050 159.600 ;
        RECT 178.950 157.950 181.050 158.400 ;
        RECT 214.950 157.950 217.050 158.400 ;
        RECT 214.950 144.600 217.050 145.050 ;
        RECT 235.950 144.600 238.050 145.050 ;
        RECT 214.950 143.400 238.050 144.600 ;
        RECT 214.950 142.950 217.050 143.400 ;
        RECT 235.950 142.950 238.050 143.400 ;
    END
  END Din[2]
  PIN Din[1]
    PORT
      LAYER metal1 ;
        RECT 184.950 216.450 189.000 217.050 ;
        RECT 184.950 214.950 189.450 216.450 ;
        RECT 188.550 211.050 189.450 214.950 ;
        RECT 184.950 209.550 189.450 211.050 ;
        RECT 184.950 208.950 189.000 209.550 ;
        RECT 184.950 138.450 189.000 139.050 ;
        RECT 184.950 136.950 189.450 138.450 ;
        RECT 188.550 133.050 189.450 136.950 ;
        RECT 184.950 131.550 189.450 133.050 ;
        RECT 184.950 130.950 189.000 131.550 ;
      LAYER metal2 ;
        RECT 170.400 254.400 171.600 256.650 ;
        RECT 350.400 254.400 351.600 256.650 ;
        RECT 170.400 246.450 171.450 254.400 ;
        RECT 170.400 245.400 174.450 246.450 ;
        RECT 173.400 232.050 174.450 245.400 ;
        RECT 350.400 244.050 351.450 254.400 ;
        RECT 361.950 253.950 364.050 256.050 ;
        RECT 362.400 244.050 363.450 253.950 ;
        RECT 349.950 241.950 352.050 244.050 ;
        RECT 361.950 241.950 364.050 244.050 ;
        RECT 274.950 232.950 277.050 235.050 ;
        RECT 301.950 232.950 304.050 235.050 ;
        RECT 172.950 229.950 175.050 232.050 ;
        RECT 184.950 229.950 187.050 232.050 ;
        RECT 268.950 229.950 271.050 232.050 ;
        RECT 185.400 217.050 186.450 229.950 ;
        RECT 269.400 220.050 270.450 229.950 ;
        RECT 275.400 220.050 276.450 232.950 ;
        RECT 302.400 229.050 303.450 232.950 ;
        RECT 350.400 229.050 351.450 241.950 ;
        RECT 301.950 226.950 304.050 229.050 ;
        RECT 349.950 226.950 352.050 229.050 ;
        RECT 268.950 217.950 271.050 220.050 ;
        RECT 274.950 217.950 277.050 220.050 ;
        RECT 184.950 214.950 187.050 217.050 ;
        RECT 184.950 208.950 187.050 211.050 ;
        RECT 185.400 187.050 186.450 208.950 ;
        RECT 184.950 184.950 187.050 187.050 ;
        RECT 163.950 175.950 166.050 178.050 ;
        RECT 164.400 148.050 165.450 175.950 ;
        RECT 142.950 145.950 145.050 148.050 ;
        RECT 163.950 145.950 166.050 148.050 ;
        RECT 184.950 145.950 187.050 148.050 ;
        RECT 143.400 138.600 144.450 145.950 ;
        RECT 185.400 139.050 186.450 145.950 ;
        RECT 143.400 136.350 144.600 138.600 ;
        RECT 184.950 136.950 187.050 139.050 ;
        RECT 184.950 127.950 187.050 133.050 ;
        RECT 241.950 127.950 244.050 130.050 ;
        RECT 242.400 109.050 243.450 127.950 ;
        RECT 241.950 106.950 244.050 109.050 ;
        RECT 241.950 94.950 244.050 97.050 ;
        RECT 242.400 60.600 243.450 94.950 ;
        RECT 242.400 58.350 243.600 60.600 ;
      LAYER metal3 ;
        RECT 361.950 255.600 364.050 256.050 ;
        RECT 361.950 254.400 369.600 255.600 ;
        RECT 361.950 253.950 364.050 254.400 ;
        RECT 349.950 243.600 352.050 244.050 ;
        RECT 361.950 243.600 364.050 244.050 ;
        RECT 349.950 242.400 364.050 243.600 ;
        RECT 349.950 241.950 352.050 242.400 ;
        RECT 361.950 241.950 364.050 242.400 ;
        RECT 274.950 234.600 277.050 235.050 ;
        RECT 301.950 234.600 304.050 235.050 ;
        RECT 274.950 233.400 304.050 234.600 ;
        RECT 274.950 232.950 277.050 233.400 ;
        RECT 301.950 232.950 304.050 233.400 ;
        RECT 172.950 231.600 175.050 232.050 ;
        RECT 184.950 231.600 187.050 232.050 ;
        RECT 268.950 231.600 271.050 232.050 ;
        RECT 172.950 230.400 271.050 231.600 ;
        RECT 172.950 229.950 175.050 230.400 ;
        RECT 184.950 229.950 187.050 230.400 ;
        RECT 268.950 229.950 271.050 230.400 ;
        RECT 301.950 228.600 304.050 229.050 ;
        RECT 349.950 228.600 352.050 229.050 ;
        RECT 301.950 227.400 352.050 228.600 ;
        RECT 301.950 226.950 304.050 227.400 ;
        RECT 349.950 226.950 352.050 227.400 ;
        RECT 268.950 219.600 271.050 220.050 ;
        RECT 274.950 219.600 277.050 220.050 ;
        RECT 268.950 218.400 277.050 219.600 ;
        RECT 268.950 217.950 271.050 218.400 ;
        RECT 274.950 217.950 277.050 218.400 ;
        RECT 184.950 186.600 187.050 187.050 ;
        RECT 176.400 185.400 187.050 186.600 ;
        RECT 176.400 180.600 177.600 185.400 ;
        RECT 184.950 184.950 187.050 185.400 ;
        RECT 164.400 180.000 177.600 180.600 ;
        RECT 163.950 179.400 177.600 180.000 ;
        RECT 163.950 175.950 166.050 179.400 ;
        RECT 142.950 147.600 145.050 148.050 ;
        RECT 163.950 147.600 166.050 148.050 ;
        RECT 184.950 147.600 187.050 148.050 ;
        RECT 142.950 146.400 187.050 147.600 ;
        RECT 142.950 145.950 145.050 146.400 ;
        RECT 163.950 145.950 166.050 146.400 ;
        RECT 184.950 145.950 187.050 146.400 ;
        RECT 184.950 129.600 187.050 130.050 ;
        RECT 241.950 129.600 244.050 130.050 ;
        RECT 184.950 128.400 244.050 129.600 ;
        RECT 184.950 127.950 187.050 128.400 ;
        RECT 241.950 127.950 244.050 128.400 ;
        RECT 241.950 106.950 244.050 109.050 ;
        RECT 242.400 97.050 243.600 106.950 ;
        RECT 241.950 94.950 244.050 97.050 ;
    END
  END Din[1]
  PIN Din[0]
    PORT
      LAYER metal1 ;
        RECT 151.950 186.450 154.050 187.050 ;
        RECT 160.950 186.450 163.050 187.050 ;
        RECT 151.950 185.550 163.050 186.450 ;
        RECT 151.950 184.950 154.050 185.550 ;
        RECT 160.950 184.950 163.050 185.550 ;
      LAYER metal2 ;
        RECT 116.400 209.400 117.600 211.650 ;
        RECT 116.400 199.050 117.450 209.400 ;
        RECT 241.950 202.950 244.050 205.050 ;
        RECT 253.950 202.950 256.050 205.050 ;
        RECT 106.950 196.950 109.050 199.050 ;
        RECT 115.950 196.950 118.050 199.050 ;
        RECT 160.950 196.950 163.050 199.050 ;
        RECT 175.950 196.950 178.050 199.050 ;
        RECT 107.400 184.050 108.450 196.950 ;
        RECT 151.950 193.950 154.050 196.050 ;
        RECT 152.400 187.050 153.450 193.950 ;
        RECT 161.400 187.050 162.450 196.950 ;
        RECT 176.400 190.050 177.450 196.950 ;
        RECT 242.400 190.050 243.450 202.950 ;
        RECT 254.400 193.050 255.450 202.950 ;
        RECT 253.950 190.950 256.050 193.050 ;
        RECT 274.950 190.950 277.050 193.050 ;
        RECT 175.950 187.950 178.050 190.050 ;
        RECT 241.950 187.950 244.050 190.050 ;
        RECT 151.950 184.950 154.050 187.050 ;
        RECT 160.950 184.950 163.050 187.050 ;
        RECT 275.400 184.050 276.450 190.950 ;
        RECT 106.950 181.950 109.050 184.050 ;
        RECT 274.950 181.950 277.050 184.050 ;
        RECT 283.800 182.100 285.900 184.200 ;
        RECT 284.400 181.350 285.600 182.100 ;
        RECT 106.950 175.950 109.050 178.050 ;
        RECT 107.400 147.450 108.450 175.950 ;
        RECT 104.400 146.400 108.450 147.450 ;
        RECT 104.400 139.050 105.450 146.400 ;
        RECT 103.950 136.950 106.050 139.050 ;
        RECT 100.950 130.950 103.050 133.050 ;
        RECT 101.400 106.200 102.450 130.950 ;
        RECT 100.950 104.100 103.050 106.200 ;
        RECT 101.400 103.350 102.600 104.100 ;
        RECT 97.950 97.950 100.050 100.050 ;
        RECT 98.400 72.450 99.450 97.950 ;
        RECT 95.400 72.000 99.450 72.450 ;
        RECT 94.950 71.400 99.450 72.000 ;
        RECT 94.950 70.050 97.050 71.400 ;
        RECT 88.950 67.950 91.050 70.050 ;
        RECT 94.800 69.000 97.050 70.050 ;
        RECT 94.800 67.950 96.900 69.000 ;
        RECT 89.400 37.050 90.450 67.950 ;
        RECT 88.950 34.950 91.050 37.050 ;
        RECT 103.950 36.450 106.050 37.050 ;
        RECT 101.400 35.400 106.050 36.450 ;
        RECT 101.400 -2.550 102.450 35.400 ;
        RECT 103.950 34.950 106.050 35.400 ;
        RECT 104.400 30.450 105.450 34.950 ;
        RECT 104.400 29.400 108.450 30.450 ;
        RECT 107.400 27.600 108.450 29.400 ;
        RECT 107.400 25.350 108.600 27.600 ;
        RECT 101.400 -3.600 105.450 -2.550 ;
      LAYER metal3 ;
        RECT 241.950 204.600 244.050 205.050 ;
        RECT 253.950 204.600 256.050 205.050 ;
        RECT 241.950 203.400 256.050 204.600 ;
        RECT 241.950 202.950 244.050 203.400 ;
        RECT 253.950 202.950 256.050 203.400 ;
        RECT 106.950 198.600 109.050 199.050 ;
        RECT 115.950 198.600 118.050 199.050 ;
        RECT 160.950 198.600 163.050 199.050 ;
        RECT 175.950 198.600 178.050 199.050 ;
        RECT 106.950 197.400 135.600 198.600 ;
        RECT 106.950 196.950 109.050 197.400 ;
        RECT 115.950 196.950 118.050 197.400 ;
        RECT 134.400 195.600 135.600 197.400 ;
        RECT 160.950 197.400 178.050 198.600 ;
        RECT 160.950 196.950 163.050 197.400 ;
        RECT 175.950 196.950 178.050 197.400 ;
        RECT 151.950 195.600 154.050 196.050 ;
        RECT 134.400 194.400 154.050 195.600 ;
        RECT 151.950 193.950 154.050 194.400 ;
        RECT 253.950 192.600 256.050 193.050 ;
        RECT 274.950 192.600 277.050 193.050 ;
        RECT 253.950 191.400 277.050 192.600 ;
        RECT 253.950 190.950 256.050 191.400 ;
        RECT 274.950 190.950 277.050 191.400 ;
        RECT 175.950 189.600 178.050 190.050 ;
        RECT 241.950 189.600 244.050 190.050 ;
        RECT 175.950 188.400 244.050 189.600 ;
        RECT 175.950 187.950 178.050 188.400 ;
        RECT 241.950 187.950 244.050 188.400 ;
        RECT 106.950 181.950 109.050 184.050 ;
        RECT 274.950 183.600 277.050 184.050 ;
        RECT 283.800 183.600 285.900 184.200 ;
        RECT 274.950 182.400 285.900 183.600 ;
        RECT 274.950 181.950 277.050 182.400 ;
        RECT 283.800 182.100 285.900 182.400 ;
        RECT 107.400 178.050 108.600 181.950 ;
        RECT 106.950 175.950 109.050 178.050 ;
        RECT 102.000 138.600 106.050 139.050 ;
        RECT 101.400 136.950 106.050 138.600 ;
        RECT 101.400 133.050 102.600 136.950 ;
        RECT 100.950 130.950 103.050 133.050 ;
        RECT 100.950 105.600 103.050 106.200 ;
        RECT 98.400 104.400 103.050 105.600 ;
        RECT 98.400 100.050 99.600 104.400 ;
        RECT 100.950 104.100 103.050 104.400 ;
        RECT 97.950 97.950 100.050 100.050 ;
        RECT 88.950 69.600 91.050 70.050 ;
        RECT 94.800 69.600 96.900 70.050 ;
        RECT 88.950 68.400 96.900 69.600 ;
        RECT 88.950 67.950 91.050 68.400 ;
        RECT 94.800 67.950 96.900 68.400 ;
        RECT 88.950 36.600 91.050 37.050 ;
        RECT 103.950 36.600 106.050 37.050 ;
        RECT 88.950 35.400 106.050 36.600 ;
        RECT 88.950 34.950 91.050 35.400 ;
        RECT 103.950 34.950 106.050 35.400 ;
    END
  END Din[0]
  PIN Dout[15]
    PORT
      LAYER metal2 ;
        RECT 128.400 20.400 129.600 22.650 ;
        RECT 128.400 -2.550 129.450 20.400 ;
        RECT 128.400 -3.600 132.450 -2.550 ;
    END
  END Dout[15]
  PIN Dout[14]
    PORT
      LAYER metal2 ;
        RECT 341.400 20.400 342.600 22.650 ;
        RECT 341.400 -2.550 342.450 20.400 ;
        RECT 338.400 -3.600 342.450 -2.550 ;
    END
  END Dout[14]
  PIN Dout[13]
    PORT
      LAYER metal2 ;
        RECT 353.400 21.900 354.600 22.650 ;
        RECT 352.950 19.800 355.050 21.900 ;
      LAYER metal3 ;
        RECT 352.950 21.600 355.050 21.900 ;
        RECT 352.950 20.400 369.600 21.600 ;
        RECT 352.950 19.800 355.050 20.400 ;
    END
  END Dout[13]
  PIN Dout[12]
    PORT
      LAYER metal2 ;
        RECT 89.400 20.400 90.600 22.650 ;
        RECT 89.400 -2.550 90.450 20.400 ;
        RECT 89.400 -3.600 93.450 -2.550 ;
    END
  END Dout[12]
  PIN Dout[11]
    PORT
      LAYER metal2 ;
        RECT 266.400 355.050 267.450 360.450 ;
        RECT 265.950 352.950 268.050 355.050 ;
        RECT 271.950 352.950 274.050 355.050 ;
        RECT 272.400 337.050 273.450 352.950 ;
        RECT 271.950 334.950 274.050 337.050 ;
        RECT 269.400 333.900 270.600 334.650 ;
        RECT 268.950 331.800 271.050 333.900 ;
      LAYER metal3 ;
        RECT 265.950 354.600 268.050 355.050 ;
        RECT 271.950 354.600 274.050 355.050 ;
        RECT 265.950 353.400 274.050 354.600 ;
        RECT 265.950 352.950 268.050 353.400 ;
        RECT 271.950 352.950 274.050 353.400 ;
        RECT 268.950 333.600 271.050 333.900 ;
        RECT 271.950 333.600 274.050 337.050 ;
        RECT 268.950 333.000 274.050 333.600 ;
        RECT 268.950 332.400 273.600 333.000 ;
        RECT 268.950 331.800 271.050 332.400 ;
    END
  END Dout[11]
  PIN Dout[10]
    PORT
      LAYER metal2 ;
        RECT 149.400 352.050 150.450 360.450 ;
        RECT 142.950 349.950 145.050 352.050 ;
        RECT 148.950 349.950 151.050 352.050 ;
        RECT 143.400 334.050 144.450 349.950 ;
        RECT 142.950 331.950 145.050 334.050 ;
        RECT 152.400 333.900 153.600 334.650 ;
        RECT 151.950 331.800 154.050 333.900 ;
      LAYER metal3 ;
        RECT 142.950 351.600 145.050 352.050 ;
        RECT 148.950 351.600 151.050 352.050 ;
        RECT 142.950 350.400 151.050 351.600 ;
        RECT 142.950 349.950 145.050 350.400 ;
        RECT 148.950 349.950 151.050 350.400 ;
        RECT 142.950 333.600 145.050 334.050 ;
        RECT 151.950 333.600 154.050 333.900 ;
        RECT 142.950 332.400 154.050 333.600 ;
        RECT 142.950 331.950 145.050 332.400 ;
        RECT 151.950 331.800 154.050 332.400 ;
    END
  END Dout[10]
  PIN Dout[9]
    PORT
      LAYER metal2 ;
        RECT 194.400 343.050 195.450 360.450 ;
        RECT 193.950 340.950 196.050 343.050 ;
        RECT 197.400 333.900 198.600 334.650 ;
        RECT 196.950 331.800 199.050 333.900 ;
      LAYER metal3 ;
        RECT 193.950 340.950 196.050 343.050 ;
        RECT 194.400 333.600 195.600 340.950 ;
        RECT 196.950 333.600 199.050 333.900 ;
        RECT 194.400 332.400 199.050 333.600 ;
        RECT 196.950 331.800 199.050 332.400 ;
    END
  END Dout[9]
  PIN Dout[8]
    PORT
      LAYER metal2 ;
        RECT 179.400 343.050 180.450 360.450 ;
        RECT 178.950 340.950 181.050 343.050 ;
        RECT 176.400 333.900 177.600 334.650 ;
        RECT 175.950 331.800 178.050 333.900 ;
      LAYER metal3 ;
        RECT 178.950 340.950 181.050 343.050 ;
        RECT 175.950 333.600 178.050 333.900 ;
        RECT 179.400 333.600 180.600 340.950 ;
        RECT 175.950 332.400 180.600 333.600 ;
        RECT 175.950 331.800 178.050 332.400 ;
    END
  END Dout[8]
  PIN Dout[7]
    PORT
      LAYER metal2 ;
        RECT 8.400 254.400 9.600 256.650 ;
        RECT 8.400 250.050 9.450 254.400 ;
        RECT 7.950 247.950 10.050 250.050 ;
      LAYER metal3 ;
        RECT -3.600 258.600 -2.400 261.600 ;
        RECT -6.600 257.400 -2.400 258.600 ;
        RECT -6.600 249.600 -5.400 257.400 ;
        RECT 7.950 249.600 10.050 250.050 ;
        RECT -6.600 248.400 10.050 249.600 ;
        RECT 7.950 247.950 10.050 248.400 ;
    END
  END Dout[7]
  PIN Dout[6]
    PORT
      LAYER metal2 ;
        RECT 20.400 98.400 21.600 100.650 ;
        RECT 20.400 94.050 21.450 98.400 ;
        RECT 19.950 91.950 22.050 94.050 ;
      LAYER metal3 ;
        RECT -3.600 93.600 -2.400 99.600 ;
        RECT 19.950 93.600 22.050 94.050 ;
        RECT -3.600 92.400 22.050 93.600 ;
        RECT 19.950 91.950 22.050 92.400 ;
    END
  END Dout[6]
  PIN Dout[5]
    PORT
      LAYER metal2 ;
        RECT 8.400 99.900 9.600 100.650 ;
        RECT 7.950 97.800 10.050 99.900 ;
      LAYER metal3 ;
        RECT -3.600 102.600 -2.400 105.600 ;
        RECT -3.600 101.400 0.600 102.600 ;
        RECT -0.600 99.600 0.600 101.400 ;
        RECT 7.950 99.600 10.050 99.900 ;
        RECT -0.600 98.400 10.050 99.600 ;
        RECT 7.950 97.800 10.050 98.400 ;
    END
  END Dout[5]
  PIN Dout[4]
    PORT
      LAYER metal2 ;
        RECT 5.400 21.900 6.600 22.650 ;
        RECT 4.950 19.800 7.050 21.900 ;
      LAYER metal3 ;
        RECT 4.950 21.600 7.050 21.900 ;
        RECT -3.600 20.400 7.050 21.600 ;
        RECT 4.950 19.800 7.050 20.400 ;
    END
  END Dout[4]
  PIN Dout[3]
    PORT
      LAYER metal2 ;
        RECT 347.400 177.900 348.600 178.650 ;
        RECT 346.950 175.800 349.050 177.900 ;
      LAYER metal3 ;
        RECT 368.400 180.600 369.600 183.600 ;
        RECT 356.400 179.400 369.600 180.600 ;
        RECT 346.950 177.600 349.050 177.900 ;
        RECT 356.400 177.600 357.600 179.400 ;
        RECT 346.950 176.400 357.600 177.600 ;
        RECT 346.950 175.800 349.050 176.400 ;
    END
  END Dout[3]
  PIN Dout[2]
    PORT
      LAYER metal2 ;
        RECT 361.950 103.950 364.050 106.050 ;
        RECT 359.400 99.450 360.600 100.650 ;
        RECT 362.400 99.450 363.450 103.950 ;
        RECT 359.400 98.400 363.450 99.450 ;
      LAYER metal3 ;
        RECT 361.950 105.600 364.050 106.050 ;
        RECT 361.950 104.400 369.600 105.600 ;
        RECT 361.950 103.950 364.050 104.400 ;
    END
  END Dout[2]
  PIN Dout[1]
    PORT
      LAYER metal2 ;
        RECT 359.400 177.900 360.600 178.650 ;
        RECT 358.950 175.800 361.050 177.900 ;
      LAYER metal3 ;
        RECT 358.950 177.600 361.050 177.900 ;
        RECT 358.950 176.400 369.600 177.600 ;
        RECT 358.950 175.800 361.050 176.400 ;
    END
  END Dout[1]
  PIN Dout[0]
    PORT
      LAYER metal2 ;
        RECT 344.400 99.900 345.600 100.650 ;
        RECT 343.950 97.800 346.050 99.900 ;
      LAYER metal3 ;
        RECT 343.950 99.600 346.050 99.900 ;
        RECT 343.950 98.400 369.600 99.600 ;
        RECT 343.950 97.800 346.050 98.400 ;
    END
  END Dout[0]
  PIN RCO
    PORT
      LAYER metal2 ;
        RECT 188.400 20.400 189.600 22.650 ;
        RECT 188.400 -2.550 189.450 20.400 ;
        RECT 185.400 -3.600 189.450 -2.550 ;
    END
  END RCO
  PIN nCLR
    PORT
      LAYER metal1 ;
        RECT 163.950 327.450 166.050 328.050 ;
        RECT 172.950 327.450 175.050 331.050 ;
        RECT 163.950 327.000 175.050 327.450 ;
        RECT 163.950 326.550 174.450 327.000 ;
        RECT 163.950 325.950 166.050 326.550 ;
      LAYER metal2 ;
        RECT 5.400 330.900 6.600 331.650 ;
        RECT 74.400 330.900 75.600 331.650 ;
        RECT 4.950 328.800 7.050 330.900 ;
        RECT 73.950 328.800 76.050 330.900 ;
        RECT 5.400 298.200 6.450 328.800 ;
        RECT 163.950 325.950 166.050 330.750 ;
        RECT 172.950 325.950 175.050 331.050 ;
        RECT 275.400 329.400 276.600 331.650 ;
        RECT 226.950 325.950 229.050 328.050 ;
        RECT 227.400 301.050 228.450 325.950 ;
        RECT 275.400 325.050 276.450 329.400 ;
        RECT 259.950 322.950 262.050 325.050 ;
        RECT 274.950 322.950 277.050 325.050 ;
        RECT 260.400 301.050 261.450 322.950 ;
        RECT 226.950 298.950 229.050 301.050 ;
        RECT 259.950 298.950 262.050 301.050 ;
        RECT 275.400 298.200 276.450 322.950 ;
        RECT 4.950 296.100 7.050 298.200 ;
        RECT 274.950 296.100 277.050 298.200 ;
        RECT 286.950 296.100 289.050 298.200 ;
        RECT 5.400 295.350 6.600 296.100 ;
        RECT 287.400 295.350 288.600 296.100 ;
        RECT 4.950 286.950 7.050 289.050 ;
        RECT 5.400 253.050 6.450 286.950 ;
        RECT 4.950 250.950 7.050 253.050 ;
        RECT 13.950 250.950 16.050 253.050 ;
        RECT 20.400 251.400 21.600 253.650 ;
        RECT 14.400 247.050 15.450 250.950 ;
        RECT 20.400 247.050 21.450 251.400 ;
        RECT 13.950 244.950 16.050 247.050 ;
        RECT 19.950 244.950 22.050 247.050 ;
        RECT 14.400 217.050 15.450 244.950 ;
        RECT 13.950 214.950 16.050 217.050 ;
        RECT 13.950 208.950 16.050 211.050 ;
        RECT 5.400 173.400 6.600 175.650 ;
        RECT 5.400 166.050 6.450 173.400 ;
        RECT 14.400 171.450 15.450 208.950 ;
        RECT 11.400 170.400 15.450 171.450 ;
        RECT 197.400 173.400 198.600 175.650 ;
        RECT 11.400 166.050 12.450 170.400 ;
        RECT 197.400 166.050 198.450 173.400 ;
        RECT 4.950 163.950 7.050 166.050 ;
        RECT 10.950 163.950 13.050 166.050 ;
        RECT 196.950 163.950 199.050 166.050 ;
        RECT 256.950 163.950 259.050 166.050 ;
        RECT 5.400 142.200 6.450 163.950 ;
        RECT 257.400 154.050 258.450 163.950 ;
        RECT 256.950 151.950 259.050 154.050 ;
        RECT 292.950 151.950 295.050 154.050 ;
        RECT 293.400 142.200 294.450 151.950 ;
        RECT 4.950 140.100 7.050 142.200 ;
        RECT 292.950 140.100 295.050 142.200 ;
        RECT 5.400 139.350 6.600 140.100 ;
        RECT 293.400 139.350 294.600 140.100 ;
        RECT 1.950 133.950 4.050 136.050 ;
        RECT 295.950 133.950 298.050 136.050 ;
        RECT 2.400 82.050 3.450 133.950 ;
        RECT 296.400 118.050 297.450 133.950 ;
        RECT 274.950 115.950 277.050 118.050 ;
        RECT 295.950 115.950 298.050 118.050 ;
        RECT 110.400 96.900 111.600 97.650 ;
        RECT 91.950 94.800 94.050 96.900 ;
        RECT 109.950 94.800 112.050 96.900 ;
        RECT 266.400 95.400 267.600 97.650 ;
        RECT 92.400 82.050 93.450 94.800 ;
        RECT 266.400 85.050 267.450 95.400 ;
        RECT 275.400 85.050 276.450 115.950 ;
        RECT 265.950 82.950 268.050 85.050 ;
        RECT 274.950 82.950 277.050 85.050 ;
        RECT 286.950 82.950 289.050 85.050 ;
        RECT 1.950 79.950 4.050 82.050 ;
        RECT 34.950 79.950 37.050 82.050 ;
        RECT 91.950 79.950 94.050 82.050 ;
        RECT 35.400 64.200 36.450 79.950 ;
        RECT 287.400 64.200 288.450 82.950 ;
        RECT 34.950 62.100 37.050 64.200 ;
        RECT 286.950 62.100 289.050 64.200 ;
        RECT 35.400 61.350 36.600 62.100 ;
        RECT 287.400 61.350 288.600 62.100 ;
        RECT 295.950 61.950 298.050 64.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 38.400 43.050 39.450 55.950 ;
        RECT 37.950 40.950 40.050 43.050 ;
        RECT 61.950 40.950 64.050 43.050 ;
        RECT 17.400 17.400 18.600 19.650 ;
        RECT 17.400 10.050 18.450 17.400 ;
        RECT 62.400 10.050 63.450 40.950 ;
        RECT 296.400 40.050 297.450 61.950 ;
        RECT 271.950 37.950 274.050 40.050 ;
        RECT 295.950 37.950 298.050 40.050 ;
        RECT 263.400 18.900 264.600 19.650 ;
        RECT 272.400 18.900 273.450 37.950 ;
        RECT 262.950 16.800 265.050 18.900 ;
        RECT 271.950 16.800 274.050 18.900 ;
        RECT 16.950 7.950 19.050 10.050 ;
        RECT 61.950 7.950 64.050 10.050 ;
        RECT 263.400 7.050 264.450 16.800 ;
        RECT 262.950 4.950 265.050 7.050 ;
      LAYER metal3 ;
        RECT 4.950 330.600 7.050 330.900 ;
        RECT 73.950 330.600 76.050 330.900 ;
        RECT 163.950 330.600 166.050 330.750 ;
        RECT 4.950 329.400 166.050 330.600 ;
        RECT 4.950 328.800 7.050 329.400 ;
        RECT 73.950 328.800 76.050 329.400 ;
        RECT 163.950 328.650 166.050 329.400 ;
        RECT 172.950 327.600 175.050 328.050 ;
        RECT 226.950 327.600 229.050 328.050 ;
        RECT 172.950 326.400 229.050 327.600 ;
        RECT 172.950 325.950 175.050 326.400 ;
        RECT 226.950 325.950 229.050 326.400 ;
        RECT 259.950 324.600 262.050 325.050 ;
        RECT 274.950 324.600 277.050 325.050 ;
        RECT 259.950 323.400 277.050 324.600 ;
        RECT 259.950 322.950 262.050 323.400 ;
        RECT 274.950 322.950 277.050 323.400 ;
        RECT 226.950 300.600 229.050 301.050 ;
        RECT 259.950 300.600 262.050 301.050 ;
        RECT 226.950 299.400 262.050 300.600 ;
        RECT 226.950 298.950 229.050 299.400 ;
        RECT 259.950 298.950 262.050 299.400 ;
        RECT 4.950 296.100 7.050 298.200 ;
        RECT 274.950 297.750 277.050 298.200 ;
        RECT 286.950 297.750 289.050 298.200 ;
        RECT 274.950 296.550 289.050 297.750 ;
        RECT 274.950 296.100 277.050 296.550 ;
        RECT 286.950 296.100 289.050 296.550 ;
        RECT 5.400 289.050 6.600 296.100 ;
        RECT 4.950 286.950 7.050 289.050 ;
        RECT -3.600 252.600 -2.400 255.600 ;
        RECT 4.950 252.600 7.050 253.050 ;
        RECT 13.950 252.600 16.050 253.050 ;
        RECT -3.600 251.400 16.050 252.600 ;
        RECT 4.950 250.950 7.050 251.400 ;
        RECT 13.950 250.950 16.050 251.400 ;
        RECT 13.950 246.600 16.050 247.050 ;
        RECT 19.950 246.600 22.050 247.050 ;
        RECT 13.950 245.400 22.050 246.600 ;
        RECT 13.950 244.950 16.050 245.400 ;
        RECT 19.950 244.950 22.050 245.400 ;
        RECT 13.950 214.950 16.050 217.050 ;
        RECT 14.400 211.050 15.600 214.950 ;
        RECT 13.950 208.950 16.050 211.050 ;
        RECT 4.950 165.600 7.050 166.050 ;
        RECT 10.950 165.600 13.050 166.050 ;
        RECT 4.950 164.400 13.050 165.600 ;
        RECT 4.950 163.950 7.050 164.400 ;
        RECT 10.950 163.950 13.050 164.400 ;
        RECT 196.950 165.600 199.050 166.050 ;
        RECT 256.950 165.600 259.050 166.050 ;
        RECT 196.950 164.400 259.050 165.600 ;
        RECT 196.950 163.950 199.050 164.400 ;
        RECT 256.950 163.950 259.050 164.400 ;
        RECT 256.950 153.600 259.050 154.050 ;
        RECT 292.950 153.600 295.050 154.050 ;
        RECT 256.950 152.400 295.050 153.600 ;
        RECT 256.950 151.950 259.050 152.400 ;
        RECT 292.950 151.950 295.050 152.400 ;
        RECT 4.950 140.100 7.050 142.200 ;
        RECT 292.950 140.100 295.050 142.200 ;
        RECT 5.400 136.050 6.600 140.100 ;
        RECT 1.950 134.400 6.600 136.050 ;
        RECT 293.400 136.050 294.600 140.100 ;
        RECT 293.400 134.400 298.050 136.050 ;
        RECT 1.950 133.950 6.000 134.400 ;
        RECT 294.000 133.950 298.050 134.400 ;
        RECT 274.950 117.600 277.050 118.050 ;
        RECT 295.950 117.600 298.050 118.050 ;
        RECT 274.950 116.400 298.050 117.600 ;
        RECT 274.950 115.950 277.050 116.400 ;
        RECT 295.950 115.950 298.050 116.400 ;
        RECT 91.950 96.450 94.050 96.900 ;
        RECT 109.950 96.450 112.050 96.900 ;
        RECT 91.950 95.250 112.050 96.450 ;
        RECT 91.950 94.800 94.050 95.250 ;
        RECT 109.950 94.800 112.050 95.250 ;
        RECT 265.950 84.600 268.050 85.050 ;
        RECT 274.950 84.600 277.050 85.050 ;
        RECT 286.950 84.600 289.050 85.050 ;
        RECT 265.950 83.400 289.050 84.600 ;
        RECT 265.950 82.950 268.050 83.400 ;
        RECT 274.950 82.950 277.050 83.400 ;
        RECT 286.950 82.950 289.050 83.400 ;
        RECT 1.950 81.600 4.050 82.050 ;
        RECT 34.950 81.600 37.050 82.050 ;
        RECT 91.950 81.600 94.050 82.050 ;
        RECT 1.950 80.400 94.050 81.600 ;
        RECT 1.950 79.950 4.050 80.400 ;
        RECT 34.950 79.950 37.050 80.400 ;
        RECT 91.950 79.950 94.050 80.400 ;
        RECT 34.950 62.100 37.050 64.200 ;
        RECT 286.950 63.600 289.050 64.200 ;
        RECT 295.950 63.600 298.050 64.050 ;
        RECT 286.950 62.400 298.050 63.600 ;
        RECT 286.950 62.100 289.050 62.400 ;
        RECT 35.400 58.050 36.600 62.100 ;
        RECT 295.950 61.950 298.050 62.400 ;
        RECT 35.400 56.400 40.050 58.050 ;
        RECT 36.000 55.950 40.050 56.400 ;
        RECT 37.950 42.600 40.050 43.050 ;
        RECT 61.950 42.600 64.050 43.050 ;
        RECT 37.950 41.400 64.050 42.600 ;
        RECT 37.950 40.950 40.050 41.400 ;
        RECT 61.950 40.950 64.050 41.400 ;
        RECT 271.950 39.600 274.050 40.050 ;
        RECT 295.950 39.600 298.050 40.050 ;
        RECT 271.950 38.400 298.050 39.600 ;
        RECT 271.950 37.950 274.050 38.400 ;
        RECT 295.950 37.950 298.050 38.400 ;
        RECT 262.950 18.450 265.050 18.900 ;
        RECT 271.950 18.450 274.050 18.900 ;
        RECT 262.950 17.250 274.050 18.450 ;
        RECT 262.950 16.800 265.050 17.250 ;
        RECT 271.950 16.800 274.050 17.250 ;
        RECT 16.950 9.600 19.050 10.050 ;
        RECT 61.950 9.600 64.050 10.050 ;
        RECT 16.950 8.400 84.600 9.600 ;
        RECT 16.950 7.950 19.050 8.400 ;
        RECT 61.950 7.950 64.050 8.400 ;
        RECT 83.400 6.600 84.600 8.400 ;
        RECT 262.950 6.600 265.050 7.050 ;
        RECT 83.400 5.400 265.050 6.600 ;
        RECT 262.950 4.950 265.050 5.400 ;
    END
  END nCLR
  PIN nLOAD
    PORT
      LAYER metal2 ;
        RECT 275.400 343.050 276.450 360.450 ;
        RECT 274.950 340.950 277.050 343.050 ;
        RECT 283.950 340.950 286.050 343.050 ;
        RECT 284.400 331.050 285.450 340.950 ;
        RECT 271.950 328.950 274.050 331.050 ;
        RECT 283.950 328.950 286.050 331.050 ;
        RECT 272.400 288.450 273.450 328.950 ;
        RECT 275.400 288.450 276.600 289.650 ;
        RECT 272.400 287.400 276.600 288.450 ;
        RECT 275.400 274.050 276.450 287.400 ;
        RECT 244.950 271.950 247.050 274.050 ;
        RECT 274.950 271.950 277.050 274.050 ;
        RECT 245.400 261.600 246.450 271.950 ;
        RECT 245.400 261.450 246.600 261.600 ;
        RECT 245.400 260.400 249.450 261.450 ;
        RECT 245.400 259.350 246.600 260.400 ;
        RECT 248.400 216.450 249.450 260.400 ;
        RECT 248.400 215.400 252.450 216.450 ;
        RECT 251.400 196.050 252.450 215.400 ;
        RECT 244.950 193.950 247.050 196.050 ;
        RECT 250.950 193.950 253.050 196.050 ;
        RECT 245.400 183.450 246.450 193.950 ;
        RECT 242.400 182.400 246.450 183.450 ;
        RECT 242.400 163.050 243.450 182.400 ;
        RECT 220.950 160.950 223.050 163.050 ;
        RECT 241.950 160.950 244.050 163.050 ;
        RECT 221.400 132.900 222.450 160.950 ;
        RECT 230.400 132.900 231.600 133.650 ;
        RECT 220.950 130.800 223.050 132.900 ;
        RECT 229.950 130.800 232.050 132.900 ;
        RECT 230.400 115.050 231.450 130.800 ;
        RECT 229.950 112.950 232.050 115.050 ;
        RECT 244.950 112.950 247.050 115.050 ;
        RECT 245.400 105.600 246.450 112.950 ;
        RECT 245.400 103.350 246.600 105.600 ;
      LAYER metal3 ;
        RECT 274.950 342.600 277.050 343.050 ;
        RECT 283.950 342.600 286.050 343.050 ;
        RECT 274.950 341.400 286.050 342.600 ;
        RECT 274.950 340.950 277.050 341.400 ;
        RECT 283.950 340.950 286.050 341.400 ;
        RECT 271.950 330.600 274.050 331.050 ;
        RECT 283.950 330.600 286.050 331.050 ;
        RECT 271.950 329.400 286.050 330.600 ;
        RECT 271.950 328.950 274.050 329.400 ;
        RECT 283.950 328.950 286.050 329.400 ;
        RECT 244.950 273.600 247.050 274.050 ;
        RECT 274.950 273.600 277.050 274.050 ;
        RECT 244.950 272.400 277.050 273.600 ;
        RECT 244.950 271.950 247.050 272.400 ;
        RECT 274.950 271.950 277.050 272.400 ;
        RECT 244.950 195.600 247.050 196.050 ;
        RECT 250.950 195.600 253.050 196.050 ;
        RECT 244.950 194.400 253.050 195.600 ;
        RECT 244.950 193.950 247.050 194.400 ;
        RECT 250.950 193.950 253.050 194.400 ;
        RECT 220.950 162.600 223.050 163.050 ;
        RECT 241.950 162.600 244.050 163.050 ;
        RECT 220.950 161.400 244.050 162.600 ;
        RECT 220.950 160.950 223.050 161.400 ;
        RECT 241.950 160.950 244.050 161.400 ;
        RECT 220.950 132.450 223.050 132.900 ;
        RECT 229.950 132.450 232.050 132.900 ;
        RECT 220.950 131.250 232.050 132.450 ;
        RECT 220.950 130.800 223.050 131.250 ;
        RECT 229.950 130.800 232.050 131.250 ;
        RECT 229.950 114.600 232.050 115.050 ;
        RECT 244.950 114.600 247.050 115.050 ;
        RECT 229.950 113.400 247.050 114.600 ;
        RECT 229.950 112.950 232.050 113.400 ;
        RECT 244.950 112.950 247.050 113.400 ;
    END
  END nLOAD
  OBS
      LAYER metal1 ;
        RECT 2.700 344.400 4.500 350.400 ;
        RECT 8.100 344.400 9.900 351.000 ;
        RECT 13.500 344.400 15.300 350.400 ;
        RECT 17.700 347.400 19.500 350.400 ;
        RECT 20.700 347.400 22.500 350.400 ;
        RECT 23.700 347.400 25.500 350.400 ;
        RECT 26.700 347.400 28.500 351.000 ;
        RECT 17.700 345.300 19.800 347.400 ;
        RECT 20.700 345.300 22.800 347.400 ;
        RECT 23.700 345.300 25.800 347.400 ;
        RECT 31.200 346.500 33.000 350.400 ;
        RECT 34.200 347.400 36.000 351.000 ;
        RECT 37.200 347.400 39.000 350.400 ;
        RECT 40.200 347.400 42.000 350.400 ;
        RECT 43.200 347.400 45.000 350.400 ;
        RECT 46.200 347.400 48.000 350.400 ;
        RECT 27.600 345.600 29.400 346.500 ;
        RECT 26.700 344.400 29.400 345.600 ;
        RECT 31.200 344.400 33.900 346.500 ;
        RECT 37.200 345.300 39.300 347.400 ;
        RECT 40.200 345.300 42.300 347.400 ;
        RECT 43.200 345.300 45.300 347.400 ;
        RECT 46.200 345.300 48.300 347.400 ;
        RECT 50.400 345.600 52.200 350.400 ;
        RECT 50.400 344.400 54.600 345.600 ;
        RECT 55.500 344.400 57.300 351.000 ;
        RECT 60.900 344.400 62.700 350.400 ;
        RECT 2.700 340.800 3.900 344.400 ;
        RECT 13.800 343.500 15.300 344.400 ;
        RECT 22.800 343.800 24.600 344.400 ;
        RECT 26.700 343.800 27.600 344.400 ;
        RECT 6.900 342.300 15.300 343.500 ;
        RECT 20.400 342.600 27.600 343.800 ;
        RECT 42.300 342.600 48.900 344.400 ;
        RECT 6.900 341.700 8.700 342.300 ;
        RECT 17.400 340.800 19.500 341.700 ;
        RECT 2.700 339.600 19.500 340.800 ;
        RECT 20.400 339.600 21.300 342.600 ;
        RECT 25.800 339.900 27.600 340.800 ;
        RECT 35.100 340.500 36.900 342.300 ;
        RECT 53.100 341.100 54.600 344.400 ;
        RECT 28.800 339.900 30.900 340.050 ;
        RECT 2.700 323.400 3.900 339.600 ;
        RECT 20.400 337.800 22.200 339.600 ;
        RECT 25.800 339.000 30.900 339.900 ;
        RECT 28.800 337.950 30.900 339.000 ;
        RECT 35.100 339.900 37.200 340.500 ;
        RECT 35.100 338.400 52.200 339.900 ;
        RECT 53.100 339.300 60.900 341.100 ;
        RECT 50.700 336.900 57.300 338.400 ;
        RECT 5.100 335.700 49.500 336.900 ;
        RECT 5.100 334.050 6.900 335.700 ;
        RECT 4.800 331.950 6.900 334.050 ;
        RECT 10.800 333.750 12.900 334.050 ;
        RECT 23.400 333.900 25.200 334.500 ;
        RECT 32.400 333.900 45.900 334.800 ;
        RECT 10.800 331.950 14.700 333.750 ;
        RECT 23.400 332.700 34.500 333.900 ;
        RECT 12.900 331.200 14.700 331.950 ;
        RECT 32.400 331.800 34.500 332.700 ;
        RECT 36.000 331.200 39.900 333.000 ;
        RECT 45.000 332.700 45.900 333.900 ;
        RECT 12.900 330.300 26.400 331.200 ;
        RECT 37.800 330.900 39.900 331.200 ;
        RECT 44.100 330.900 45.900 332.700 ;
        RECT 48.600 334.200 49.500 335.700 ;
        RECT 48.600 332.400 53.700 334.200 ;
        RECT 55.800 334.050 57.300 336.900 ;
        RECT 55.800 331.950 57.900 334.050 ;
        RECT 25.200 329.700 26.400 330.300 ;
        RECT 59.100 329.700 60.900 330.300 ;
        RECT 20.400 328.500 22.500 328.800 ;
        RECT 25.200 328.500 60.900 329.700 ;
        RECT 10.500 327.300 22.500 328.500 ;
        RECT 61.800 327.600 62.700 344.400 ;
        RECT 10.500 326.700 12.300 327.300 ;
        RECT 20.400 326.700 22.500 327.300 ;
        RECT 25.200 326.400 42.900 327.600 ;
        RECT 7.200 325.800 9.000 326.100 ;
        RECT 25.200 325.800 26.400 326.400 ;
        RECT 7.200 324.600 26.400 325.800 ;
        RECT 40.800 325.500 42.900 326.400 ;
        RECT 46.200 326.700 62.700 327.600 ;
        RECT 46.200 325.500 48.300 326.700 ;
        RECT 7.200 324.300 9.000 324.600 ;
        RECT 2.700 322.500 6.300 323.400 ;
        RECT 5.400 321.600 6.300 322.500 ;
        RECT 2.700 315.000 4.500 321.600 ;
        RECT 5.400 320.700 7.500 321.600 ;
        RECT 5.700 315.600 7.500 320.700 ;
        RECT 8.700 315.000 10.500 321.600 ;
        RECT 11.700 315.600 13.500 324.600 ;
        RECT 23.700 321.600 25.800 323.700 ;
        RECT 31.200 323.100 34.500 325.200 ;
        RECT 14.700 315.000 16.500 321.600 ;
        RECT 18.300 318.600 20.400 320.700 ;
        RECT 21.300 318.600 23.400 320.700 ;
        RECT 18.300 315.600 20.100 318.600 ;
        RECT 21.300 315.600 23.100 318.600 ;
        RECT 24.300 315.600 26.100 321.600 ;
        RECT 27.300 315.000 29.100 321.600 ;
        RECT 31.200 315.600 33.000 323.100 ;
        RECT 37.200 321.600 39.900 325.500 ;
        RECT 52.200 324.600 57.900 325.800 ;
        RECT 49.500 323.700 51.300 324.300 ;
        RECT 43.200 322.500 51.300 323.700 ;
        RECT 43.200 321.600 45.300 322.500 ;
        RECT 52.200 321.600 53.400 324.600 ;
        RECT 56.100 324.000 57.900 324.600 ;
        RECT 61.800 323.400 62.700 326.700 ;
        RECT 58.800 322.500 62.700 323.400 ;
        RECT 64.500 347.400 66.300 350.400 ;
        RECT 67.500 347.400 69.300 351.000 ;
        RECT 64.500 334.050 66.000 347.400 ;
        RECT 71.700 344.400 73.500 350.400 ;
        RECT 77.100 344.400 78.900 351.000 ;
        RECT 82.500 344.400 84.300 350.400 ;
        RECT 86.700 347.400 88.500 350.400 ;
        RECT 89.700 347.400 91.500 350.400 ;
        RECT 92.700 347.400 94.500 350.400 ;
        RECT 95.700 347.400 97.500 351.000 ;
        RECT 86.700 345.300 88.800 347.400 ;
        RECT 89.700 345.300 91.800 347.400 ;
        RECT 92.700 345.300 94.800 347.400 ;
        RECT 100.200 346.500 102.000 350.400 ;
        RECT 103.200 347.400 105.000 351.000 ;
        RECT 106.200 347.400 108.000 350.400 ;
        RECT 109.200 347.400 111.000 350.400 ;
        RECT 112.200 347.400 114.000 350.400 ;
        RECT 115.200 347.400 117.000 350.400 ;
        RECT 96.600 345.600 98.400 346.500 ;
        RECT 95.700 344.400 98.400 345.600 ;
        RECT 100.200 344.400 102.900 346.500 ;
        RECT 106.200 345.300 108.300 347.400 ;
        RECT 109.200 345.300 111.300 347.400 ;
        RECT 112.200 345.300 114.300 347.400 ;
        RECT 115.200 345.300 117.300 347.400 ;
        RECT 119.400 345.600 121.200 350.400 ;
        RECT 119.400 344.400 123.600 345.600 ;
        RECT 124.500 344.400 126.300 351.000 ;
        RECT 129.900 344.400 131.700 350.400 ;
        RECT 71.700 340.800 72.900 344.400 ;
        RECT 82.800 343.500 84.300 344.400 ;
        RECT 91.800 343.800 93.600 344.400 ;
        RECT 95.700 343.800 96.600 344.400 ;
        RECT 75.900 342.300 84.300 343.500 ;
        RECT 89.400 342.600 96.600 343.800 ;
        RECT 111.300 342.600 117.900 344.400 ;
        RECT 75.900 341.700 77.700 342.300 ;
        RECT 86.400 340.800 88.500 341.700 ;
        RECT 71.700 339.600 88.500 340.800 ;
        RECT 89.400 339.600 90.300 342.600 ;
        RECT 94.800 339.900 96.600 340.800 ;
        RECT 104.100 340.500 105.900 342.300 ;
        RECT 122.100 341.100 123.600 344.400 ;
        RECT 97.800 339.900 99.900 340.050 ;
        RECT 64.500 331.950 66.900 334.050 ;
        RECT 58.800 321.600 60.000 322.500 ;
        RECT 64.500 321.600 66.000 331.950 ;
        RECT 71.700 323.400 72.900 339.600 ;
        RECT 89.400 337.800 91.200 339.600 ;
        RECT 94.800 339.000 99.900 339.900 ;
        RECT 97.800 337.950 99.900 339.000 ;
        RECT 104.100 339.900 106.200 340.500 ;
        RECT 104.100 338.400 121.200 339.900 ;
        RECT 122.100 339.300 129.900 341.100 ;
        RECT 119.700 336.900 126.300 338.400 ;
        RECT 74.100 335.700 118.500 336.900 ;
        RECT 74.100 334.050 75.900 335.700 ;
        RECT 73.800 331.950 75.900 334.050 ;
        RECT 79.800 333.750 81.900 334.050 ;
        RECT 92.400 333.900 94.200 334.500 ;
        RECT 101.400 333.900 114.900 334.800 ;
        RECT 79.800 331.950 83.700 333.750 ;
        RECT 92.400 332.700 103.500 333.900 ;
        RECT 81.900 331.200 83.700 331.950 ;
        RECT 101.400 331.800 103.500 332.700 ;
        RECT 105.000 331.200 108.900 333.000 ;
        RECT 114.000 332.700 114.900 333.900 ;
        RECT 81.900 330.300 95.400 331.200 ;
        RECT 106.800 330.900 108.900 331.200 ;
        RECT 113.100 330.900 114.900 332.700 ;
        RECT 117.600 334.200 118.500 335.700 ;
        RECT 117.600 332.400 122.700 334.200 ;
        RECT 124.800 334.050 126.300 336.900 ;
        RECT 124.800 331.950 126.900 334.050 ;
        RECT 94.200 329.700 95.400 330.300 ;
        RECT 128.100 329.700 129.900 330.300 ;
        RECT 89.400 328.500 91.500 328.800 ;
        RECT 94.200 328.500 129.900 329.700 ;
        RECT 79.500 327.300 91.500 328.500 ;
        RECT 130.800 327.600 131.700 344.400 ;
        RECT 79.500 326.700 81.300 327.300 ;
        RECT 89.400 326.700 91.500 327.300 ;
        RECT 94.200 326.400 111.900 327.600 ;
        RECT 76.200 325.800 78.000 326.100 ;
        RECT 94.200 325.800 95.400 326.400 ;
        RECT 76.200 324.600 95.400 325.800 ;
        RECT 109.800 325.500 111.900 326.400 ;
        RECT 115.200 326.700 131.700 327.600 ;
        RECT 115.200 325.500 117.300 326.700 ;
        RECT 76.200 324.300 78.000 324.600 ;
        RECT 71.700 322.500 75.300 323.400 ;
        RECT 74.400 321.600 75.300 322.500 ;
        RECT 34.200 315.000 36.000 321.600 ;
        RECT 37.200 315.600 39.000 321.600 ;
        RECT 40.200 318.600 42.300 320.700 ;
        RECT 43.200 318.600 45.300 320.700 ;
        RECT 46.200 318.600 48.300 320.700 ;
        RECT 40.200 315.600 42.000 318.600 ;
        RECT 43.200 315.600 45.000 318.600 ;
        RECT 46.200 315.600 48.000 318.600 ;
        RECT 49.200 315.000 51.000 321.600 ;
        RECT 52.200 315.600 54.000 321.600 ;
        RECT 55.200 315.000 57.000 321.600 ;
        RECT 58.200 315.600 60.000 321.600 ;
        RECT 61.200 315.000 63.000 321.600 ;
        RECT 64.500 315.600 66.300 321.600 ;
        RECT 67.500 315.000 69.300 321.600 ;
        RECT 71.700 315.000 73.500 321.600 ;
        RECT 74.400 320.700 76.500 321.600 ;
        RECT 74.700 315.600 76.500 320.700 ;
        RECT 77.700 315.000 79.500 321.600 ;
        RECT 80.700 315.600 82.500 324.600 ;
        RECT 92.700 321.600 94.800 323.700 ;
        RECT 100.200 323.100 103.500 325.200 ;
        RECT 83.700 315.000 85.500 321.600 ;
        RECT 87.300 318.600 89.400 320.700 ;
        RECT 90.300 318.600 92.400 320.700 ;
        RECT 87.300 315.600 89.100 318.600 ;
        RECT 90.300 315.600 92.100 318.600 ;
        RECT 93.300 315.600 95.100 321.600 ;
        RECT 96.300 315.000 98.100 321.600 ;
        RECT 100.200 315.600 102.000 323.100 ;
        RECT 106.200 321.600 108.900 325.500 ;
        RECT 121.200 324.600 126.900 325.800 ;
        RECT 118.500 323.700 120.300 324.300 ;
        RECT 112.200 322.500 120.300 323.700 ;
        RECT 112.200 321.600 114.300 322.500 ;
        RECT 121.200 321.600 122.400 324.600 ;
        RECT 125.100 324.000 126.900 324.600 ;
        RECT 130.800 323.400 131.700 326.700 ;
        RECT 127.800 322.500 131.700 323.400 ;
        RECT 133.500 347.400 135.300 350.400 ;
        RECT 136.500 347.400 138.300 351.000 ;
        RECT 146.100 347.400 147.900 350.400 ;
        RECT 133.500 334.050 135.000 347.400 ;
        RECT 146.100 343.500 147.300 347.400 ;
        RECT 149.100 344.400 150.900 351.000 ;
        RECT 152.100 344.400 153.900 350.400 ;
        RECT 146.100 342.600 151.800 343.500 ;
        RECT 150.000 341.700 151.800 342.600 ;
        RECT 146.400 334.950 148.500 337.050 ;
        RECT 133.500 331.950 135.900 334.050 ;
        RECT 146.400 333.150 148.200 334.950 ;
        RECT 127.800 321.600 129.000 322.500 ;
        RECT 133.500 321.600 135.000 331.950 ;
        RECT 150.000 330.300 150.900 341.700 ;
        RECT 152.700 337.050 153.900 344.400 ;
        RECT 163.500 342.000 165.300 350.400 ;
        RECT 162.000 340.800 165.300 342.000 ;
        RECT 170.100 341.400 171.900 351.000 ;
        RECT 176.100 344.400 177.900 350.400 ;
        RECT 179.100 344.400 180.900 351.000 ;
        RECT 182.100 347.400 183.900 350.400 ;
        RECT 162.000 337.050 162.900 340.800 ;
        RECT 164.100 337.050 165.900 338.850 ;
        RECT 170.100 337.050 171.900 338.850 ;
        RECT 176.100 337.050 177.300 344.400 ;
        RECT 182.700 343.500 183.900 347.400 ;
        RECT 178.200 342.600 183.900 343.500 ;
        RECT 191.100 347.400 192.900 350.400 ;
        RECT 191.100 343.500 192.300 347.400 ;
        RECT 194.100 344.400 195.900 351.000 ;
        RECT 197.100 344.400 198.900 350.400 ;
        RECT 206.100 344.400 207.900 350.400 ;
        RECT 191.100 342.600 196.800 343.500 ;
        RECT 178.200 341.700 180.000 342.600 ;
        RECT 151.800 334.950 153.900 337.050 ;
        RECT 160.950 334.950 163.050 337.050 ;
        RECT 163.950 334.950 166.050 337.050 ;
        RECT 166.950 334.950 169.050 337.050 ;
        RECT 169.950 334.950 172.050 337.050 ;
        RECT 176.100 334.950 178.200 337.050 ;
        RECT 150.000 329.400 151.800 330.300 ;
        RECT 146.100 328.500 151.800 329.400 ;
        RECT 146.100 321.600 147.300 328.500 ;
        RECT 152.700 327.600 153.900 334.950 ;
        RECT 103.200 315.000 105.000 321.600 ;
        RECT 106.200 315.600 108.000 321.600 ;
        RECT 109.200 318.600 111.300 320.700 ;
        RECT 112.200 318.600 114.300 320.700 ;
        RECT 115.200 318.600 117.300 320.700 ;
        RECT 109.200 315.600 111.000 318.600 ;
        RECT 112.200 315.600 114.000 318.600 ;
        RECT 115.200 315.600 117.000 318.600 ;
        RECT 118.200 315.000 120.000 321.600 ;
        RECT 121.200 315.600 123.000 321.600 ;
        RECT 124.200 315.000 126.000 321.600 ;
        RECT 127.200 315.600 129.000 321.600 ;
        RECT 130.200 315.000 132.000 321.600 ;
        RECT 133.500 315.600 135.300 321.600 ;
        RECT 136.500 315.000 138.300 321.600 ;
        RECT 146.100 315.600 147.900 321.600 ;
        RECT 149.100 315.000 150.900 325.800 ;
        RECT 152.100 315.600 153.900 327.600 ;
        RECT 162.000 322.800 162.900 334.950 ;
        RECT 167.100 333.150 168.900 334.950 ;
        RECT 176.100 327.600 177.300 334.950 ;
        RECT 179.100 330.300 180.000 341.700 ;
        RECT 195.000 341.700 196.800 342.600 ;
        RECT 181.500 334.950 183.600 337.050 ;
        RECT 181.800 333.150 183.600 334.950 ;
        RECT 191.400 334.950 193.500 337.050 ;
        RECT 191.400 333.150 193.200 334.950 ;
        RECT 178.200 329.400 180.000 330.300 ;
        RECT 195.000 330.300 195.900 341.700 ;
        RECT 197.700 337.050 198.900 344.400 ;
        RECT 206.700 342.300 207.900 344.400 ;
        RECT 209.100 345.300 210.900 350.400 ;
        RECT 212.100 346.200 213.900 351.000 ;
        RECT 215.100 345.300 216.900 350.400 ;
        RECT 221.100 347.400 222.900 351.000 ;
        RECT 224.100 347.400 225.900 350.400 ;
        RECT 227.100 347.400 228.900 351.000 ;
        RECT 209.100 343.950 216.900 345.300 ;
        RECT 206.700 341.400 210.300 342.300 ;
        RECT 206.100 337.050 207.900 338.850 ;
        RECT 209.100 337.050 210.300 341.400 ;
        RECT 212.100 337.050 213.900 338.850 ;
        RECT 224.700 337.050 225.600 347.400 ;
        RECT 233.100 342.600 234.900 350.400 ;
        RECT 237.600 344.400 239.400 351.000 ;
        RECT 240.600 346.200 242.400 350.400 ;
        RECT 240.600 344.400 243.300 346.200 ;
        RECT 239.700 342.600 241.500 343.500 ;
        RECT 233.100 341.700 241.500 342.600 ;
        RECT 233.250 337.050 235.050 338.850 ;
        RECT 196.800 334.950 198.900 337.050 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 211.950 334.950 214.050 337.050 ;
        RECT 214.950 334.950 217.050 337.050 ;
        RECT 220.950 334.950 223.050 337.050 ;
        RECT 223.950 334.950 226.050 337.050 ;
        RECT 226.950 334.950 229.050 337.050 ;
        RECT 233.100 334.950 235.200 337.050 ;
        RECT 195.000 329.400 196.800 330.300 ;
        RECT 178.200 328.500 183.900 329.400 ;
        RECT 162.000 321.900 168.600 322.800 ;
        RECT 162.000 321.600 162.900 321.900 ;
        RECT 161.100 315.600 162.900 321.600 ;
        RECT 167.100 321.600 168.600 321.900 ;
        RECT 164.100 315.000 165.900 321.000 ;
        RECT 167.100 315.600 168.900 321.600 ;
        RECT 170.100 315.000 171.900 321.600 ;
        RECT 176.100 315.600 177.900 327.600 ;
        RECT 179.100 315.000 180.900 325.800 ;
        RECT 182.700 321.600 183.900 328.500 ;
        RECT 182.100 315.600 183.900 321.600 ;
        RECT 191.100 328.500 196.800 329.400 ;
        RECT 191.100 321.600 192.300 328.500 ;
        RECT 197.700 327.600 198.900 334.950 ;
        RECT 191.100 315.600 192.900 321.600 ;
        RECT 194.100 315.000 195.900 325.800 ;
        RECT 197.100 315.600 198.900 327.600 ;
        RECT 209.100 327.600 210.300 334.950 ;
        RECT 215.100 333.150 216.900 334.950 ;
        RECT 221.100 333.150 222.900 334.950 ;
        RECT 224.700 327.600 225.600 334.950 ;
        RECT 226.950 333.150 228.750 334.950 ;
        RECT 209.100 326.100 211.500 327.600 ;
        RECT 207.000 323.100 208.800 324.900 ;
        RECT 206.700 315.000 208.500 321.600 ;
        RECT 209.700 315.600 211.500 326.100 ;
        RECT 214.800 315.000 216.600 327.600 ;
        RECT 222.000 326.400 225.600 327.600 ;
        RECT 222.000 315.600 223.800 326.400 ;
        RECT 227.100 315.000 228.900 327.600 ;
        RECT 236.100 321.600 237.000 341.700 ;
        RECT 242.400 337.050 243.300 344.400 ;
        RECT 248.100 345.300 249.900 350.400 ;
        RECT 251.100 346.200 252.900 351.000 ;
        RECT 254.100 345.300 255.900 350.400 ;
        RECT 248.100 343.950 255.900 345.300 ;
        RECT 257.100 344.400 258.900 350.400 ;
        RECT 263.100 347.400 264.900 350.400 ;
        RECT 257.100 342.300 258.300 344.400 ;
        RECT 263.100 343.500 264.300 347.400 ;
        RECT 266.100 344.400 267.900 351.000 ;
        RECT 269.100 344.400 270.900 350.400 ;
        RECT 263.100 342.600 268.800 343.500 ;
        RECT 254.700 341.400 258.300 342.300 ;
        RECT 267.000 341.700 268.800 342.600 ;
        RECT 251.100 337.050 252.900 338.850 ;
        RECT 254.700 337.050 255.900 341.400 ;
        RECT 257.100 337.050 258.900 338.850 ;
        RECT 238.500 334.950 240.600 337.050 ;
        RECT 241.800 334.950 243.900 337.050 ;
        RECT 247.950 334.950 250.050 337.050 ;
        RECT 250.950 334.950 253.050 337.050 ;
        RECT 253.950 334.950 256.050 337.050 ;
        RECT 256.950 334.950 259.050 337.050 ;
        RECT 263.400 334.950 265.500 337.050 ;
        RECT 238.200 333.150 240.000 334.950 ;
        RECT 242.400 327.600 243.300 334.950 ;
        RECT 248.100 333.150 249.900 334.950 ;
        RECT 254.700 327.600 255.900 334.950 ;
        RECT 263.400 333.150 265.200 334.950 ;
        RECT 267.000 330.300 267.900 341.700 ;
        RECT 269.700 337.050 270.900 344.400 ;
        RECT 268.800 334.950 270.900 337.050 ;
        RECT 267.000 329.400 268.800 330.300 ;
        RECT 233.100 315.000 234.900 321.600 ;
        RECT 236.100 315.600 237.900 321.600 ;
        RECT 239.100 315.000 240.900 327.000 ;
        RECT 242.100 315.600 243.900 327.600 ;
        RECT 248.400 315.000 250.200 327.600 ;
        RECT 253.500 326.100 255.900 327.600 ;
        RECT 263.100 328.500 268.800 329.400 ;
        RECT 253.500 315.600 255.300 326.100 ;
        RECT 256.200 323.100 258.000 324.900 ;
        RECT 263.100 321.600 264.300 328.500 ;
        RECT 269.700 327.600 270.900 334.950 ;
        RECT 256.500 315.000 258.300 321.600 ;
        RECT 263.100 315.600 264.900 321.600 ;
        RECT 266.100 315.000 267.900 325.800 ;
        RECT 269.100 315.600 270.900 327.600 ;
        RECT 272.700 344.400 274.500 350.400 ;
        RECT 278.100 344.400 279.900 351.000 ;
        RECT 283.500 344.400 285.300 350.400 ;
        RECT 287.700 347.400 289.500 350.400 ;
        RECT 290.700 347.400 292.500 350.400 ;
        RECT 293.700 347.400 295.500 350.400 ;
        RECT 296.700 347.400 298.500 351.000 ;
        RECT 287.700 345.300 289.800 347.400 ;
        RECT 290.700 345.300 292.800 347.400 ;
        RECT 293.700 345.300 295.800 347.400 ;
        RECT 301.200 346.500 303.000 350.400 ;
        RECT 304.200 347.400 306.000 351.000 ;
        RECT 307.200 347.400 309.000 350.400 ;
        RECT 310.200 347.400 312.000 350.400 ;
        RECT 313.200 347.400 315.000 350.400 ;
        RECT 316.200 347.400 318.000 350.400 ;
        RECT 297.600 345.600 299.400 346.500 ;
        RECT 296.700 344.400 299.400 345.600 ;
        RECT 301.200 344.400 303.900 346.500 ;
        RECT 307.200 345.300 309.300 347.400 ;
        RECT 310.200 345.300 312.300 347.400 ;
        RECT 313.200 345.300 315.300 347.400 ;
        RECT 316.200 345.300 318.300 347.400 ;
        RECT 320.400 345.600 322.200 350.400 ;
        RECT 320.400 344.400 324.600 345.600 ;
        RECT 325.500 344.400 327.300 351.000 ;
        RECT 330.900 344.400 332.700 350.400 ;
        RECT 272.700 340.800 273.900 344.400 ;
        RECT 283.800 343.500 285.300 344.400 ;
        RECT 292.800 343.800 294.600 344.400 ;
        RECT 296.700 343.800 297.600 344.400 ;
        RECT 276.900 342.300 285.300 343.500 ;
        RECT 290.400 342.600 297.600 343.800 ;
        RECT 312.300 342.600 318.900 344.400 ;
        RECT 276.900 341.700 278.700 342.300 ;
        RECT 287.400 340.800 289.500 341.700 ;
        RECT 272.700 339.600 289.500 340.800 ;
        RECT 290.400 339.600 291.300 342.600 ;
        RECT 295.800 339.900 297.600 340.800 ;
        RECT 305.100 340.500 306.900 342.300 ;
        RECT 323.100 341.100 324.600 344.400 ;
        RECT 298.800 339.900 300.900 340.050 ;
        RECT 272.700 323.400 273.900 339.600 ;
        RECT 290.400 337.800 292.200 339.600 ;
        RECT 295.800 339.000 300.900 339.900 ;
        RECT 298.800 337.950 300.900 339.000 ;
        RECT 305.100 339.900 307.200 340.500 ;
        RECT 305.100 338.400 322.200 339.900 ;
        RECT 323.100 339.300 330.900 341.100 ;
        RECT 320.700 336.900 327.300 338.400 ;
        RECT 275.100 335.700 319.500 336.900 ;
        RECT 275.100 334.050 276.900 335.700 ;
        RECT 274.800 331.950 276.900 334.050 ;
        RECT 280.800 333.750 282.900 334.050 ;
        RECT 293.400 333.900 295.200 334.500 ;
        RECT 302.400 333.900 315.900 334.800 ;
        RECT 280.800 331.950 284.700 333.750 ;
        RECT 293.400 332.700 304.500 333.900 ;
        RECT 282.900 331.200 284.700 331.950 ;
        RECT 302.400 331.800 304.500 332.700 ;
        RECT 306.000 331.200 309.900 333.000 ;
        RECT 315.000 332.700 315.900 333.900 ;
        RECT 282.900 330.300 296.400 331.200 ;
        RECT 307.800 330.900 309.900 331.200 ;
        RECT 314.100 330.900 315.900 332.700 ;
        RECT 318.600 334.200 319.500 335.700 ;
        RECT 318.600 332.400 323.700 334.200 ;
        RECT 325.800 334.050 327.300 336.900 ;
        RECT 325.800 331.950 327.900 334.050 ;
        RECT 295.200 329.700 296.400 330.300 ;
        RECT 329.100 329.700 330.900 330.300 ;
        RECT 290.400 328.500 292.500 328.800 ;
        RECT 295.200 328.500 330.900 329.700 ;
        RECT 280.500 327.300 292.500 328.500 ;
        RECT 331.800 327.600 332.700 344.400 ;
        RECT 280.500 326.700 282.300 327.300 ;
        RECT 290.400 326.700 292.500 327.300 ;
        RECT 295.200 326.400 312.900 327.600 ;
        RECT 277.200 325.800 279.000 326.100 ;
        RECT 295.200 325.800 296.400 326.400 ;
        RECT 277.200 324.600 296.400 325.800 ;
        RECT 310.800 325.500 312.900 326.400 ;
        RECT 316.200 326.700 332.700 327.600 ;
        RECT 316.200 325.500 318.300 326.700 ;
        RECT 277.200 324.300 279.000 324.600 ;
        RECT 272.700 322.500 276.300 323.400 ;
        RECT 275.400 321.600 276.300 322.500 ;
        RECT 272.700 315.000 274.500 321.600 ;
        RECT 275.400 320.700 277.500 321.600 ;
        RECT 275.700 315.600 277.500 320.700 ;
        RECT 278.700 315.000 280.500 321.600 ;
        RECT 281.700 315.600 283.500 324.600 ;
        RECT 293.700 321.600 295.800 323.700 ;
        RECT 301.200 323.100 304.500 325.200 ;
        RECT 284.700 315.000 286.500 321.600 ;
        RECT 288.300 318.600 290.400 320.700 ;
        RECT 291.300 318.600 293.400 320.700 ;
        RECT 288.300 315.600 290.100 318.600 ;
        RECT 291.300 315.600 293.100 318.600 ;
        RECT 294.300 315.600 296.100 321.600 ;
        RECT 297.300 315.000 299.100 321.600 ;
        RECT 301.200 315.600 303.000 323.100 ;
        RECT 307.200 321.600 309.900 325.500 ;
        RECT 322.200 324.600 327.900 325.800 ;
        RECT 319.500 323.700 321.300 324.300 ;
        RECT 313.200 322.500 321.300 323.700 ;
        RECT 313.200 321.600 315.300 322.500 ;
        RECT 322.200 321.600 323.400 324.600 ;
        RECT 326.100 324.000 327.900 324.600 ;
        RECT 331.800 323.400 332.700 326.700 ;
        RECT 328.800 322.500 332.700 323.400 ;
        RECT 334.500 347.400 336.300 350.400 ;
        RECT 337.500 347.400 339.300 351.000 ;
        RECT 334.500 334.050 336.000 347.400 ;
        RECT 347.700 343.200 349.500 350.400 ;
        RECT 352.800 344.400 354.600 351.000 ;
        RECT 347.700 342.300 351.900 343.200 ;
        RECT 347.100 337.050 348.900 338.850 ;
        RECT 350.700 337.050 351.900 342.300 ;
        RECT 352.950 337.050 354.750 338.850 ;
        RECT 346.950 334.950 349.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 352.950 334.950 355.050 337.050 ;
        RECT 334.500 331.950 336.900 334.050 ;
        RECT 328.800 321.600 330.000 322.500 ;
        RECT 334.500 321.600 336.000 331.950 ;
        RECT 350.700 321.600 351.900 334.950 ;
        RECT 304.200 315.000 306.000 321.600 ;
        RECT 307.200 315.600 309.000 321.600 ;
        RECT 310.200 318.600 312.300 320.700 ;
        RECT 313.200 318.600 315.300 320.700 ;
        RECT 316.200 318.600 318.300 320.700 ;
        RECT 310.200 315.600 312.000 318.600 ;
        RECT 313.200 315.600 315.000 318.600 ;
        RECT 316.200 315.600 318.000 318.600 ;
        RECT 319.200 315.000 321.000 321.600 ;
        RECT 322.200 315.600 324.000 321.600 ;
        RECT 325.200 315.000 327.000 321.600 ;
        RECT 328.200 315.600 330.000 321.600 ;
        RECT 331.200 315.000 333.000 321.600 ;
        RECT 334.500 315.600 336.300 321.600 ;
        RECT 337.500 315.000 339.300 321.600 ;
        RECT 347.100 315.000 348.900 321.600 ;
        RECT 350.100 315.600 351.900 321.600 ;
        RECT 353.100 315.000 354.900 321.600 ;
        RECT 2.700 305.400 4.500 312.000 ;
        RECT 5.700 306.300 7.500 311.400 ;
        RECT 5.400 305.400 7.500 306.300 ;
        RECT 8.700 305.400 10.500 312.000 ;
        RECT 5.400 304.500 6.300 305.400 ;
        RECT 2.700 303.600 6.300 304.500 ;
        RECT 2.700 287.400 3.900 303.600 ;
        RECT 7.200 302.400 9.000 302.700 ;
        RECT 11.700 302.400 13.500 311.400 ;
        RECT 14.700 305.400 16.500 312.000 ;
        RECT 18.300 308.400 20.100 311.400 ;
        RECT 21.300 308.400 23.100 311.400 ;
        RECT 18.300 306.300 20.400 308.400 ;
        RECT 21.300 306.300 23.400 308.400 ;
        RECT 24.300 305.400 26.100 311.400 ;
        RECT 27.300 305.400 29.100 312.000 ;
        RECT 23.700 303.300 25.800 305.400 ;
        RECT 31.200 303.900 33.000 311.400 ;
        RECT 34.200 305.400 36.000 312.000 ;
        RECT 37.200 305.400 39.000 311.400 ;
        RECT 40.200 308.400 42.000 311.400 ;
        RECT 43.200 308.400 45.000 311.400 ;
        RECT 46.200 308.400 48.000 311.400 ;
        RECT 40.200 306.300 42.300 308.400 ;
        RECT 43.200 306.300 45.300 308.400 ;
        RECT 46.200 306.300 48.300 308.400 ;
        RECT 49.200 305.400 51.000 312.000 ;
        RECT 52.200 305.400 54.000 311.400 ;
        RECT 55.200 305.400 57.000 312.000 ;
        RECT 58.200 305.400 60.000 311.400 ;
        RECT 61.200 305.400 63.000 312.000 ;
        RECT 64.500 305.400 66.300 311.400 ;
        RECT 67.500 305.400 69.300 312.000 ;
        RECT 77.100 305.400 78.900 311.400 ;
        RECT 80.100 306.000 81.900 312.000 ;
        RECT 7.200 301.200 26.400 302.400 ;
        RECT 31.200 301.800 34.500 303.900 ;
        RECT 37.200 301.500 39.900 305.400 ;
        RECT 43.200 304.500 45.300 305.400 ;
        RECT 43.200 303.300 51.300 304.500 ;
        RECT 49.500 302.700 51.300 303.300 ;
        RECT 52.200 302.400 53.400 305.400 ;
        RECT 58.800 304.500 60.000 305.400 ;
        RECT 58.800 303.600 62.700 304.500 ;
        RECT 56.100 302.400 57.900 303.000 ;
        RECT 7.200 300.900 9.000 301.200 ;
        RECT 25.200 300.600 26.400 301.200 ;
        RECT 40.800 300.600 42.900 301.500 ;
        RECT 10.500 299.700 12.300 300.300 ;
        RECT 20.400 299.700 22.500 300.300 ;
        RECT 10.500 298.500 22.500 299.700 ;
        RECT 25.200 299.400 42.900 300.600 ;
        RECT 46.200 300.300 48.300 301.500 ;
        RECT 52.200 301.200 57.900 302.400 ;
        RECT 61.800 300.300 62.700 303.600 ;
        RECT 46.200 299.400 62.700 300.300 ;
        RECT 20.400 298.200 22.500 298.500 ;
        RECT 25.200 297.300 60.900 298.500 ;
        RECT 25.200 296.700 26.400 297.300 ;
        RECT 59.100 296.700 60.900 297.300 ;
        RECT 12.900 295.800 26.400 296.700 ;
        RECT 37.800 295.800 39.900 296.100 ;
        RECT 12.900 295.050 14.700 295.800 ;
        RECT 4.800 292.950 6.900 295.050 ;
        RECT 10.800 293.250 14.700 295.050 ;
        RECT 32.400 294.300 34.500 295.200 ;
        RECT 10.800 292.950 12.900 293.250 ;
        RECT 23.400 293.100 34.500 294.300 ;
        RECT 36.000 294.000 39.900 295.800 ;
        RECT 44.100 294.300 45.900 296.100 ;
        RECT 45.000 293.100 45.900 294.300 ;
        RECT 5.100 291.300 6.900 292.950 ;
        RECT 23.400 292.500 25.200 293.100 ;
        RECT 32.400 292.200 45.900 293.100 ;
        RECT 48.600 292.800 53.700 294.600 ;
        RECT 55.800 292.950 57.900 295.050 ;
        RECT 48.600 291.300 49.500 292.800 ;
        RECT 5.100 290.100 49.500 291.300 ;
        RECT 55.800 290.100 57.300 292.950 ;
        RECT 20.400 287.400 22.200 289.200 ;
        RECT 28.800 288.000 30.900 289.050 ;
        RECT 50.700 288.600 57.300 290.100 ;
        RECT 2.700 286.200 19.500 287.400 ;
        RECT 2.700 282.600 3.900 286.200 ;
        RECT 17.400 285.300 19.500 286.200 ;
        RECT 6.900 284.700 8.700 285.300 ;
        RECT 6.900 283.500 15.300 284.700 ;
        RECT 13.800 282.600 15.300 283.500 ;
        RECT 20.400 284.400 21.300 287.400 ;
        RECT 25.800 287.100 30.900 288.000 ;
        RECT 25.800 286.200 27.600 287.100 ;
        RECT 28.800 286.950 30.900 287.100 ;
        RECT 35.100 287.100 52.200 288.600 ;
        RECT 35.100 286.500 37.200 287.100 ;
        RECT 35.100 284.700 36.900 286.500 ;
        RECT 53.100 285.900 60.900 287.700 ;
        RECT 20.400 283.200 27.600 284.400 ;
        RECT 22.800 282.600 24.600 283.200 ;
        RECT 26.700 282.600 27.600 283.200 ;
        RECT 42.300 282.600 48.900 284.400 ;
        RECT 53.100 282.600 54.600 285.900 ;
        RECT 61.800 282.600 62.700 299.400 ;
        RECT 2.700 276.600 4.500 282.600 ;
        RECT 8.100 276.000 9.900 282.600 ;
        RECT 13.500 276.600 15.300 282.600 ;
        RECT 17.700 279.600 19.800 281.700 ;
        RECT 20.700 279.600 22.800 281.700 ;
        RECT 23.700 279.600 25.800 281.700 ;
        RECT 26.700 281.400 29.400 282.600 ;
        RECT 27.600 280.500 29.400 281.400 ;
        RECT 31.200 280.500 33.900 282.600 ;
        RECT 17.700 276.600 19.500 279.600 ;
        RECT 20.700 276.600 22.500 279.600 ;
        RECT 23.700 276.600 25.500 279.600 ;
        RECT 26.700 276.000 28.500 279.600 ;
        RECT 31.200 276.600 33.000 280.500 ;
        RECT 37.200 279.600 39.300 281.700 ;
        RECT 40.200 279.600 42.300 281.700 ;
        RECT 43.200 279.600 45.300 281.700 ;
        RECT 46.200 279.600 48.300 281.700 ;
        RECT 50.400 281.400 54.600 282.600 ;
        RECT 34.200 276.000 36.000 279.600 ;
        RECT 37.200 276.600 39.000 279.600 ;
        RECT 40.200 276.600 42.000 279.600 ;
        RECT 43.200 276.600 45.000 279.600 ;
        RECT 46.200 276.600 48.000 279.600 ;
        RECT 50.400 276.600 52.200 281.400 ;
        RECT 55.500 276.000 57.300 282.600 ;
        RECT 60.900 276.600 62.700 282.600 ;
        RECT 64.500 295.050 66.000 305.400 ;
        RECT 78.000 305.100 78.900 305.400 ;
        RECT 83.100 305.400 84.900 311.400 ;
        RECT 86.100 305.400 87.900 312.000 ;
        RECT 92.100 305.400 93.900 312.000 ;
        RECT 95.100 305.400 96.900 311.400 ;
        RECT 98.100 305.400 99.900 312.000 ;
        RECT 107.100 305.400 108.900 312.000 ;
        RECT 110.100 305.400 111.900 311.400 ;
        RECT 113.100 305.400 114.900 312.000 ;
        RECT 119.100 305.400 120.900 312.000 ;
        RECT 122.100 305.400 123.900 311.400 ;
        RECT 131.700 305.400 133.500 312.000 ;
        RECT 83.100 305.100 84.600 305.400 ;
        RECT 78.000 304.200 84.600 305.100 ;
        RECT 64.500 292.950 66.900 295.050 ;
        RECT 64.500 279.600 66.000 292.950 ;
        RECT 78.000 292.050 78.900 304.200 ;
        RECT 83.100 292.050 84.900 293.850 ;
        RECT 95.100 292.050 96.300 305.400 ;
        RECT 110.100 292.050 111.300 305.400 ;
        RECT 119.100 292.050 120.900 293.850 ;
        RECT 122.100 292.050 123.300 305.400 ;
        RECT 132.000 302.100 133.800 303.900 ;
        RECT 134.700 300.900 136.500 311.400 ;
        RECT 134.100 299.400 136.500 300.900 ;
        RECT 139.800 299.400 141.600 312.000 ;
        RECT 146.100 305.400 147.900 311.400 ;
        RECT 149.100 306.000 150.900 312.000 ;
        RECT 147.000 305.100 147.900 305.400 ;
        RECT 152.100 305.400 153.900 311.400 ;
        RECT 155.100 305.400 156.900 312.000 ;
        RECT 164.100 305.400 165.900 311.400 ;
        RECT 167.100 305.400 168.900 312.000 ;
        RECT 152.100 305.100 153.600 305.400 ;
        RECT 147.000 304.200 153.600 305.100 ;
        RECT 134.100 292.050 135.300 299.400 ;
        RECT 140.100 292.050 141.900 293.850 ;
        RECT 147.000 292.050 147.900 304.200 ;
        RECT 152.100 292.050 153.900 293.850 ;
        RECT 164.700 292.050 165.900 305.400 ;
        RECT 173.100 299.400 174.900 311.400 ;
        RECT 176.100 300.300 177.900 311.400 ;
        RECT 179.100 301.200 180.900 312.000 ;
        RECT 182.100 300.300 183.900 311.400 ;
        RECT 188.100 305.400 189.900 311.400 ;
        RECT 191.100 305.400 192.900 312.000 ;
        RECT 176.100 299.400 183.900 300.300 ;
        RECT 167.100 292.050 168.900 293.850 ;
        RECT 173.400 292.050 174.300 299.400 ;
        RECT 178.950 292.050 180.750 293.850 ;
        RECT 188.700 292.050 189.900 305.400 ;
        RECT 197.400 299.400 199.200 312.000 ;
        RECT 202.500 300.900 204.300 311.400 ;
        RECT 205.500 305.400 207.300 312.000 ;
        RECT 215.100 305.400 216.900 312.000 ;
        RECT 218.100 305.400 219.900 311.400 ;
        RECT 221.100 305.400 222.900 312.000 ;
        RECT 230.100 305.400 231.900 312.000 ;
        RECT 233.100 305.400 234.900 311.400 ;
        RECT 236.100 305.400 237.900 312.000 ;
        RECT 205.200 302.100 207.000 303.900 ;
        RECT 202.500 299.400 204.900 300.900 ;
        RECT 191.100 292.050 192.900 293.850 ;
        RECT 197.100 292.050 198.900 293.850 ;
        RECT 203.700 292.050 204.900 299.400 ;
        RECT 218.700 292.050 219.900 305.400 ;
        RECT 233.700 292.050 234.900 305.400 ;
        RECT 242.100 299.400 243.900 311.400 ;
        RECT 245.100 300.000 246.900 312.000 ;
        RECT 248.100 305.400 249.900 311.400 ;
        RECT 251.100 305.400 252.900 312.000 ;
        RECT 257.100 305.400 258.900 311.400 ;
        RECT 260.100 306.000 261.900 312.000 ;
        RECT 242.700 292.050 243.600 299.400 ;
        RECT 246.000 292.050 247.800 293.850 ;
        RECT 76.950 289.950 79.050 292.050 ;
        RECT 79.950 289.950 82.050 292.050 ;
        RECT 82.950 289.950 85.050 292.050 ;
        RECT 85.950 289.950 88.050 292.050 ;
        RECT 91.950 289.950 94.050 292.050 ;
        RECT 94.950 289.950 97.050 292.050 ;
        RECT 97.950 289.950 100.050 292.050 ;
        RECT 106.950 289.950 109.050 292.050 ;
        RECT 109.950 289.950 112.050 292.050 ;
        RECT 112.950 289.950 115.050 292.050 ;
        RECT 118.950 289.950 121.050 292.050 ;
        RECT 121.950 289.950 124.050 292.050 ;
        RECT 130.950 289.950 133.050 292.050 ;
        RECT 133.950 289.950 136.050 292.050 ;
        RECT 136.950 289.950 139.050 292.050 ;
        RECT 139.950 289.950 142.050 292.050 ;
        RECT 145.950 289.950 148.050 292.050 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 154.950 289.950 157.050 292.050 ;
        RECT 163.950 289.950 166.050 292.050 ;
        RECT 166.950 289.950 169.050 292.050 ;
        RECT 172.950 289.950 175.050 292.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 178.950 289.950 181.050 292.050 ;
        RECT 181.950 289.950 184.050 292.050 ;
        RECT 187.950 289.950 190.050 292.050 ;
        RECT 190.950 289.950 193.050 292.050 ;
        RECT 196.950 289.950 199.050 292.050 ;
        RECT 199.950 289.950 202.050 292.050 ;
        RECT 202.950 289.950 205.050 292.050 ;
        RECT 205.950 289.950 208.050 292.050 ;
        RECT 214.950 289.950 217.050 292.050 ;
        RECT 217.950 289.950 220.050 292.050 ;
        RECT 220.950 289.950 223.050 292.050 ;
        RECT 229.950 289.950 232.050 292.050 ;
        RECT 232.950 289.950 235.050 292.050 ;
        RECT 235.950 289.950 238.050 292.050 ;
        RECT 242.100 289.950 244.200 292.050 ;
        RECT 245.400 289.950 247.500 292.050 ;
        RECT 78.000 286.200 78.900 289.950 ;
        RECT 80.100 288.150 81.900 289.950 ;
        RECT 86.100 288.150 87.900 289.950 ;
        RECT 92.250 288.150 94.050 289.950 ;
        RECT 78.000 285.000 81.300 286.200 ;
        RECT 64.500 276.600 66.300 279.600 ;
        RECT 67.500 276.000 69.300 279.600 ;
        RECT 79.500 276.600 81.300 285.000 ;
        RECT 86.100 276.000 87.900 285.600 ;
        RECT 95.100 284.700 96.300 289.950 ;
        RECT 98.100 288.150 99.900 289.950 ;
        RECT 107.250 288.150 109.050 289.950 ;
        RECT 110.100 284.700 111.300 289.950 ;
        RECT 113.100 288.150 114.900 289.950 ;
        RECT 95.100 283.800 99.300 284.700 ;
        RECT 110.100 283.800 114.300 284.700 ;
        RECT 92.400 276.000 94.200 282.600 ;
        RECT 97.500 276.600 99.300 283.800 ;
        RECT 107.400 276.000 109.200 282.600 ;
        RECT 112.500 276.600 114.300 283.800 ;
        RECT 122.100 279.600 123.300 289.950 ;
        RECT 131.100 288.150 132.900 289.950 ;
        RECT 134.100 285.600 135.300 289.950 ;
        RECT 137.100 288.150 138.900 289.950 ;
        RECT 131.700 284.700 135.300 285.600 ;
        RECT 147.000 286.200 147.900 289.950 ;
        RECT 149.100 288.150 150.900 289.950 ;
        RECT 155.100 288.150 156.900 289.950 ;
        RECT 147.000 285.000 150.300 286.200 ;
        RECT 131.700 282.600 132.900 284.700 ;
        RECT 119.100 276.000 120.900 279.600 ;
        RECT 122.100 276.600 123.900 279.600 ;
        RECT 131.100 276.600 132.900 282.600 ;
        RECT 134.100 281.700 141.900 283.050 ;
        RECT 134.100 276.600 135.900 281.700 ;
        RECT 137.100 276.000 138.900 280.800 ;
        RECT 140.100 276.600 141.900 281.700 ;
        RECT 148.500 276.600 150.300 285.000 ;
        RECT 155.100 276.000 156.900 285.600 ;
        RECT 164.700 279.600 165.900 289.950 ;
        RECT 173.400 282.600 174.300 289.950 ;
        RECT 175.950 288.150 177.750 289.950 ;
        RECT 182.100 288.150 183.900 289.950 ;
        RECT 173.400 281.400 178.500 282.600 ;
        RECT 164.100 276.600 165.900 279.600 ;
        RECT 167.100 276.000 168.900 279.600 ;
        RECT 173.700 276.000 175.500 279.600 ;
        RECT 176.700 276.600 178.500 281.400 ;
        RECT 181.200 276.000 183.000 282.600 ;
        RECT 188.700 279.600 189.900 289.950 ;
        RECT 200.100 288.150 201.900 289.950 ;
        RECT 203.700 285.600 204.900 289.950 ;
        RECT 206.100 288.150 207.900 289.950 ;
        RECT 215.100 288.150 216.900 289.950 ;
        RECT 203.700 284.700 207.300 285.600 ;
        RECT 218.700 284.700 219.900 289.950 ;
        RECT 220.950 288.150 222.750 289.950 ;
        RECT 230.100 288.150 231.900 289.950 ;
        RECT 233.700 284.700 234.900 289.950 ;
        RECT 235.950 288.150 237.750 289.950 ;
        RECT 197.100 281.700 204.900 283.050 ;
        RECT 188.100 276.600 189.900 279.600 ;
        RECT 191.100 276.000 192.900 279.600 ;
        RECT 197.100 276.600 198.900 281.700 ;
        RECT 200.100 276.000 201.900 280.800 ;
        RECT 203.100 276.600 204.900 281.700 ;
        RECT 206.100 282.600 207.300 284.700 ;
        RECT 215.700 283.800 219.900 284.700 ;
        RECT 230.700 283.800 234.900 284.700 ;
        RECT 206.100 276.600 207.900 282.600 ;
        RECT 215.700 276.600 217.500 283.800 ;
        RECT 220.800 276.000 222.600 282.600 ;
        RECT 230.700 276.600 232.500 283.800 ;
        RECT 242.700 282.600 243.600 289.950 ;
        RECT 249.000 285.300 249.900 305.400 ;
        RECT 258.000 305.100 258.900 305.400 ;
        RECT 263.100 305.400 264.900 311.400 ;
        RECT 266.100 305.400 267.900 312.000 ;
        RECT 275.100 305.400 276.900 311.400 ;
        RECT 263.100 305.100 264.600 305.400 ;
        RECT 258.000 304.200 264.600 305.100 ;
        RECT 258.000 292.050 258.900 304.200 ;
        RECT 275.100 298.500 276.300 305.400 ;
        RECT 278.100 301.200 279.900 312.000 ;
        RECT 281.100 299.400 282.900 311.400 ;
        RECT 284.700 305.400 286.500 312.000 ;
        RECT 287.700 306.300 289.500 311.400 ;
        RECT 287.400 305.400 289.500 306.300 ;
        RECT 290.700 305.400 292.500 312.000 ;
        RECT 287.400 304.500 288.300 305.400 ;
        RECT 275.100 297.600 280.800 298.500 ;
        RECT 279.000 296.700 280.800 297.600 ;
        RECT 263.100 292.050 264.900 293.850 ;
        RECT 275.400 292.050 277.200 293.850 ;
        RECT 250.800 289.950 252.900 292.050 ;
        RECT 256.950 289.950 259.050 292.050 ;
        RECT 259.950 289.950 262.050 292.050 ;
        RECT 262.950 289.950 265.050 292.050 ;
        RECT 265.950 289.950 268.050 292.050 ;
        RECT 275.400 289.950 277.500 292.050 ;
        RECT 250.950 288.150 252.750 289.950 ;
        RECT 258.000 286.200 258.900 289.950 ;
        RECT 260.100 288.150 261.900 289.950 ;
        RECT 266.100 288.150 267.900 289.950 ;
        RECT 244.500 284.400 252.900 285.300 ;
        RECT 258.000 285.000 261.300 286.200 ;
        RECT 244.500 283.500 246.300 284.400 ;
        RECT 235.800 276.000 237.600 282.600 ;
        RECT 242.700 280.800 245.400 282.600 ;
        RECT 243.600 276.600 245.400 280.800 ;
        RECT 246.600 276.000 248.400 282.600 ;
        RECT 251.100 276.600 252.900 284.400 ;
        RECT 259.500 276.600 261.300 285.000 ;
        RECT 266.100 276.000 267.900 285.600 ;
        RECT 279.000 285.300 279.900 296.700 ;
        RECT 281.700 292.050 282.900 299.400 ;
        RECT 280.800 289.950 282.900 292.050 ;
        RECT 279.000 284.400 280.800 285.300 ;
        RECT 275.100 283.500 280.800 284.400 ;
        RECT 275.100 279.600 276.300 283.500 ;
        RECT 281.700 282.600 282.900 289.950 ;
        RECT 275.100 276.600 276.900 279.600 ;
        RECT 278.100 276.000 279.900 282.600 ;
        RECT 281.100 276.600 282.900 282.600 ;
        RECT 284.700 303.600 288.300 304.500 ;
        RECT 284.700 287.400 285.900 303.600 ;
        RECT 289.200 302.400 291.000 302.700 ;
        RECT 293.700 302.400 295.500 311.400 ;
        RECT 296.700 305.400 298.500 312.000 ;
        RECT 300.300 308.400 302.100 311.400 ;
        RECT 303.300 308.400 305.100 311.400 ;
        RECT 300.300 306.300 302.400 308.400 ;
        RECT 303.300 306.300 305.400 308.400 ;
        RECT 306.300 305.400 308.100 311.400 ;
        RECT 309.300 305.400 311.100 312.000 ;
        RECT 305.700 303.300 307.800 305.400 ;
        RECT 313.200 303.900 315.000 311.400 ;
        RECT 316.200 305.400 318.000 312.000 ;
        RECT 319.200 305.400 321.000 311.400 ;
        RECT 322.200 308.400 324.000 311.400 ;
        RECT 325.200 308.400 327.000 311.400 ;
        RECT 328.200 308.400 330.000 311.400 ;
        RECT 322.200 306.300 324.300 308.400 ;
        RECT 325.200 306.300 327.300 308.400 ;
        RECT 328.200 306.300 330.300 308.400 ;
        RECT 331.200 305.400 333.000 312.000 ;
        RECT 334.200 305.400 336.000 311.400 ;
        RECT 337.200 305.400 339.000 312.000 ;
        RECT 340.200 305.400 342.000 311.400 ;
        RECT 343.200 305.400 345.000 312.000 ;
        RECT 346.500 305.400 348.300 311.400 ;
        RECT 349.500 305.400 351.300 312.000 ;
        RECT 289.200 301.200 308.400 302.400 ;
        RECT 313.200 301.800 316.500 303.900 ;
        RECT 319.200 301.500 321.900 305.400 ;
        RECT 325.200 304.500 327.300 305.400 ;
        RECT 325.200 303.300 333.300 304.500 ;
        RECT 331.500 302.700 333.300 303.300 ;
        RECT 334.200 302.400 335.400 305.400 ;
        RECT 340.800 304.500 342.000 305.400 ;
        RECT 340.800 303.600 344.700 304.500 ;
        RECT 338.100 302.400 339.900 303.000 ;
        RECT 289.200 300.900 291.000 301.200 ;
        RECT 307.200 300.600 308.400 301.200 ;
        RECT 322.800 300.600 324.900 301.500 ;
        RECT 292.500 299.700 294.300 300.300 ;
        RECT 302.400 299.700 304.500 300.300 ;
        RECT 292.500 298.500 304.500 299.700 ;
        RECT 307.200 299.400 324.900 300.600 ;
        RECT 328.200 300.300 330.300 301.500 ;
        RECT 334.200 301.200 339.900 302.400 ;
        RECT 343.800 300.300 344.700 303.600 ;
        RECT 328.200 299.400 344.700 300.300 ;
        RECT 302.400 298.200 304.500 298.500 ;
        RECT 307.200 297.300 342.900 298.500 ;
        RECT 307.200 296.700 308.400 297.300 ;
        RECT 341.100 296.700 342.900 297.300 ;
        RECT 294.900 295.800 308.400 296.700 ;
        RECT 319.800 295.800 321.900 296.100 ;
        RECT 294.900 295.050 296.700 295.800 ;
        RECT 286.800 292.950 288.900 295.050 ;
        RECT 292.800 293.250 296.700 295.050 ;
        RECT 314.400 294.300 316.500 295.200 ;
        RECT 292.800 292.950 294.900 293.250 ;
        RECT 305.400 293.100 316.500 294.300 ;
        RECT 318.000 294.000 321.900 295.800 ;
        RECT 326.100 294.300 327.900 296.100 ;
        RECT 327.000 293.100 327.900 294.300 ;
        RECT 287.100 291.300 288.900 292.950 ;
        RECT 305.400 292.500 307.200 293.100 ;
        RECT 314.400 292.200 327.900 293.100 ;
        RECT 330.600 292.800 335.700 294.600 ;
        RECT 337.800 292.950 339.900 295.050 ;
        RECT 330.600 291.300 331.500 292.800 ;
        RECT 287.100 290.100 331.500 291.300 ;
        RECT 337.800 290.100 339.300 292.950 ;
        RECT 302.400 287.400 304.200 289.200 ;
        RECT 310.800 288.000 312.900 289.050 ;
        RECT 332.700 288.600 339.300 290.100 ;
        RECT 284.700 286.200 301.500 287.400 ;
        RECT 284.700 282.600 285.900 286.200 ;
        RECT 299.400 285.300 301.500 286.200 ;
        RECT 288.900 284.700 290.700 285.300 ;
        RECT 288.900 283.500 297.300 284.700 ;
        RECT 295.800 282.600 297.300 283.500 ;
        RECT 302.400 284.400 303.300 287.400 ;
        RECT 307.800 287.100 312.900 288.000 ;
        RECT 307.800 286.200 309.600 287.100 ;
        RECT 310.800 286.950 312.900 287.100 ;
        RECT 317.100 287.100 334.200 288.600 ;
        RECT 317.100 286.500 319.200 287.100 ;
        RECT 317.100 284.700 318.900 286.500 ;
        RECT 335.100 285.900 342.900 287.700 ;
        RECT 302.400 283.200 309.600 284.400 ;
        RECT 304.800 282.600 306.600 283.200 ;
        RECT 308.700 282.600 309.600 283.200 ;
        RECT 324.300 282.600 330.900 284.400 ;
        RECT 335.100 282.600 336.600 285.900 ;
        RECT 343.800 282.600 344.700 299.400 ;
        RECT 284.700 276.600 286.500 282.600 ;
        RECT 290.100 276.000 291.900 282.600 ;
        RECT 295.500 276.600 297.300 282.600 ;
        RECT 299.700 279.600 301.800 281.700 ;
        RECT 302.700 279.600 304.800 281.700 ;
        RECT 305.700 279.600 307.800 281.700 ;
        RECT 308.700 281.400 311.400 282.600 ;
        RECT 309.600 280.500 311.400 281.400 ;
        RECT 313.200 280.500 315.900 282.600 ;
        RECT 299.700 276.600 301.500 279.600 ;
        RECT 302.700 276.600 304.500 279.600 ;
        RECT 305.700 276.600 307.500 279.600 ;
        RECT 308.700 276.000 310.500 279.600 ;
        RECT 313.200 276.600 315.000 280.500 ;
        RECT 319.200 279.600 321.300 281.700 ;
        RECT 322.200 279.600 324.300 281.700 ;
        RECT 325.200 279.600 327.300 281.700 ;
        RECT 328.200 279.600 330.300 281.700 ;
        RECT 332.400 281.400 336.600 282.600 ;
        RECT 316.200 276.000 318.000 279.600 ;
        RECT 319.200 276.600 321.000 279.600 ;
        RECT 322.200 276.600 324.000 279.600 ;
        RECT 325.200 276.600 327.000 279.600 ;
        RECT 328.200 276.600 330.000 279.600 ;
        RECT 332.400 276.600 334.200 281.400 ;
        RECT 337.500 276.000 339.300 282.600 ;
        RECT 342.900 276.600 344.700 282.600 ;
        RECT 346.500 295.050 348.000 305.400 ;
        RECT 346.500 292.950 348.900 295.050 ;
        RECT 346.500 279.600 348.000 292.950 ;
        RECT 346.500 276.600 348.300 279.600 ;
        RECT 349.500 276.000 351.300 279.600 ;
        RECT 8.100 266.400 9.900 272.400 ;
        RECT 11.100 266.400 12.900 273.000 ;
        RECT 14.100 269.400 15.900 272.400 ;
        RECT 8.100 259.050 9.300 266.400 ;
        RECT 14.700 265.500 15.900 269.400 ;
        RECT 10.200 264.600 15.900 265.500 ;
        RECT 17.700 266.400 19.500 272.400 ;
        RECT 23.100 266.400 24.900 273.000 ;
        RECT 28.500 266.400 30.300 272.400 ;
        RECT 32.700 269.400 34.500 272.400 ;
        RECT 35.700 269.400 37.500 272.400 ;
        RECT 38.700 269.400 40.500 272.400 ;
        RECT 41.700 269.400 43.500 273.000 ;
        RECT 32.700 267.300 34.800 269.400 ;
        RECT 35.700 267.300 37.800 269.400 ;
        RECT 38.700 267.300 40.800 269.400 ;
        RECT 46.200 268.500 48.000 272.400 ;
        RECT 49.200 269.400 51.000 273.000 ;
        RECT 52.200 269.400 54.000 272.400 ;
        RECT 55.200 269.400 57.000 272.400 ;
        RECT 58.200 269.400 60.000 272.400 ;
        RECT 61.200 269.400 63.000 272.400 ;
        RECT 42.600 267.600 44.400 268.500 ;
        RECT 41.700 266.400 44.400 267.600 ;
        RECT 46.200 266.400 48.900 268.500 ;
        RECT 52.200 267.300 54.300 269.400 ;
        RECT 55.200 267.300 57.300 269.400 ;
        RECT 58.200 267.300 60.300 269.400 ;
        RECT 61.200 267.300 63.300 269.400 ;
        RECT 65.400 267.600 67.200 272.400 ;
        RECT 65.400 266.400 69.600 267.600 ;
        RECT 70.500 266.400 72.300 273.000 ;
        RECT 75.900 266.400 77.700 272.400 ;
        RECT 10.200 263.700 12.000 264.600 ;
        RECT 8.100 256.950 10.200 259.050 ;
        RECT 8.100 249.600 9.300 256.950 ;
        RECT 11.100 252.300 12.000 263.700 ;
        RECT 17.700 262.800 18.900 266.400 ;
        RECT 28.800 265.500 30.300 266.400 ;
        RECT 37.800 265.800 39.600 266.400 ;
        RECT 41.700 265.800 42.600 266.400 ;
        RECT 21.900 264.300 30.300 265.500 ;
        RECT 35.400 264.600 42.600 265.800 ;
        RECT 57.300 264.600 63.900 266.400 ;
        RECT 21.900 263.700 23.700 264.300 ;
        RECT 32.400 262.800 34.500 263.700 ;
        RECT 17.700 261.600 34.500 262.800 ;
        RECT 35.400 261.600 36.300 264.600 ;
        RECT 40.800 261.900 42.600 262.800 ;
        RECT 50.100 262.500 51.900 264.300 ;
        RECT 68.100 263.100 69.600 266.400 ;
        RECT 43.800 261.900 45.900 262.050 ;
        RECT 13.500 256.950 15.600 259.050 ;
        RECT 13.800 255.150 15.600 256.950 ;
        RECT 10.200 251.400 12.000 252.300 ;
        RECT 10.200 250.500 15.900 251.400 ;
        RECT 8.100 237.600 9.900 249.600 ;
        RECT 11.100 237.000 12.900 247.800 ;
        RECT 14.700 243.600 15.900 250.500 ;
        RECT 17.700 245.400 18.900 261.600 ;
        RECT 35.400 259.800 37.200 261.600 ;
        RECT 40.800 261.000 45.900 261.900 ;
        RECT 43.800 259.950 45.900 261.000 ;
        RECT 50.100 261.900 52.200 262.500 ;
        RECT 50.100 260.400 67.200 261.900 ;
        RECT 68.100 261.300 75.900 263.100 ;
        RECT 65.700 258.900 72.300 260.400 ;
        RECT 20.100 257.700 64.500 258.900 ;
        RECT 20.100 256.050 21.900 257.700 ;
        RECT 19.800 253.950 21.900 256.050 ;
        RECT 25.800 255.750 27.900 256.050 ;
        RECT 38.400 255.900 40.200 256.500 ;
        RECT 47.400 255.900 60.900 256.800 ;
        RECT 25.800 253.950 29.700 255.750 ;
        RECT 38.400 254.700 49.500 255.900 ;
        RECT 27.900 253.200 29.700 253.950 ;
        RECT 47.400 253.800 49.500 254.700 ;
        RECT 51.000 253.200 54.900 255.000 ;
        RECT 60.000 254.700 60.900 255.900 ;
        RECT 27.900 252.300 41.400 253.200 ;
        RECT 52.800 252.900 54.900 253.200 ;
        RECT 59.100 252.900 60.900 254.700 ;
        RECT 63.600 256.200 64.500 257.700 ;
        RECT 63.600 254.400 68.700 256.200 ;
        RECT 70.800 256.050 72.300 258.900 ;
        RECT 70.800 253.950 72.900 256.050 ;
        RECT 40.200 251.700 41.400 252.300 ;
        RECT 74.100 251.700 75.900 252.300 ;
        RECT 35.400 250.500 37.500 250.800 ;
        RECT 40.200 250.500 75.900 251.700 ;
        RECT 25.500 249.300 37.500 250.500 ;
        RECT 76.800 249.600 77.700 266.400 ;
        RECT 25.500 248.700 27.300 249.300 ;
        RECT 35.400 248.700 37.500 249.300 ;
        RECT 40.200 248.400 57.900 249.600 ;
        RECT 22.200 247.800 24.000 248.100 ;
        RECT 40.200 247.800 41.400 248.400 ;
        RECT 22.200 246.600 41.400 247.800 ;
        RECT 55.800 247.500 57.900 248.400 ;
        RECT 61.200 248.700 77.700 249.600 ;
        RECT 61.200 247.500 63.300 248.700 ;
        RECT 22.200 246.300 24.000 246.600 ;
        RECT 17.700 244.500 21.300 245.400 ;
        RECT 20.400 243.600 21.300 244.500 ;
        RECT 14.100 237.600 15.900 243.600 ;
        RECT 17.700 237.000 19.500 243.600 ;
        RECT 20.400 242.700 22.500 243.600 ;
        RECT 20.700 237.600 22.500 242.700 ;
        RECT 23.700 237.000 25.500 243.600 ;
        RECT 26.700 237.600 28.500 246.600 ;
        RECT 38.700 243.600 40.800 245.700 ;
        RECT 46.200 245.100 49.500 247.200 ;
        RECT 29.700 237.000 31.500 243.600 ;
        RECT 33.300 240.600 35.400 242.700 ;
        RECT 36.300 240.600 38.400 242.700 ;
        RECT 33.300 237.600 35.100 240.600 ;
        RECT 36.300 237.600 38.100 240.600 ;
        RECT 39.300 237.600 41.100 243.600 ;
        RECT 42.300 237.000 44.100 243.600 ;
        RECT 46.200 237.600 48.000 245.100 ;
        RECT 52.200 243.600 54.900 247.500 ;
        RECT 67.200 246.600 72.900 247.800 ;
        RECT 64.500 245.700 66.300 246.300 ;
        RECT 58.200 244.500 66.300 245.700 ;
        RECT 58.200 243.600 60.300 244.500 ;
        RECT 67.200 243.600 68.400 246.600 ;
        RECT 71.100 246.000 72.900 246.600 ;
        RECT 76.800 245.400 77.700 248.700 ;
        RECT 73.800 244.500 77.700 245.400 ;
        RECT 79.500 269.400 81.300 272.400 ;
        RECT 82.500 269.400 84.300 273.000 ;
        RECT 79.500 256.050 81.000 269.400 ;
        RECT 89.400 266.400 91.200 273.000 ;
        RECT 94.500 265.200 96.300 272.400 ;
        RECT 104.100 266.400 105.900 272.400 ;
        RECT 92.100 264.300 96.300 265.200 ;
        RECT 104.700 264.300 105.900 266.400 ;
        RECT 107.100 267.300 108.900 272.400 ;
        RECT 110.100 268.200 111.900 273.000 ;
        RECT 113.100 267.300 114.900 272.400 ;
        RECT 122.700 269.400 124.500 273.000 ;
        RECT 125.700 267.600 127.500 272.400 ;
        RECT 107.100 265.950 114.900 267.300 ;
        RECT 122.400 266.400 127.500 267.600 ;
        RECT 130.200 266.400 132.000 273.000 ;
        RECT 140.100 269.400 141.900 272.400 ;
        RECT 143.100 269.400 144.900 273.000 ;
        RECT 89.250 259.050 91.050 260.850 ;
        RECT 92.100 259.050 93.300 264.300 ;
        RECT 104.700 263.400 108.300 264.300 ;
        RECT 95.100 259.050 96.900 260.850 ;
        RECT 104.100 259.050 105.900 260.850 ;
        RECT 107.100 259.050 108.300 263.400 ;
        RECT 110.100 259.050 111.900 260.850 ;
        RECT 122.400 259.050 123.300 266.400 ;
        RECT 124.950 259.050 126.750 260.850 ;
        RECT 131.100 259.050 132.900 260.850 ;
        RECT 140.700 259.050 141.900 269.400 ;
        RECT 149.100 263.400 150.900 273.000 ;
        RECT 155.700 264.000 157.500 272.400 ;
        RECT 167.100 267.000 168.900 272.400 ;
        RECT 170.100 267.900 171.900 273.000 ;
        RECT 173.100 271.500 180.900 272.400 ;
        RECT 173.100 267.000 174.900 271.500 ;
        RECT 167.100 266.100 174.900 267.000 ;
        RECT 176.100 266.400 177.900 270.600 ;
        RECT 179.100 266.400 180.900 271.500 ;
        RECT 160.950 264.450 163.050 265.050 ;
        RECT 176.400 264.900 177.300 266.400 ;
        RECT 188.700 265.200 190.500 272.400 ;
        RECT 193.800 266.400 195.600 273.000 ;
        RECT 200.100 269.400 201.900 272.400 ;
        RECT 203.100 269.400 204.900 273.000 ;
        RECT 166.950 264.450 169.050 264.900 ;
        RECT 155.700 262.800 159.000 264.000 ;
        RECT 160.950 263.550 169.050 264.450 ;
        RECT 160.950 262.950 163.050 263.550 ;
        RECT 166.950 262.800 169.050 263.550 ;
        RECT 172.950 263.700 177.300 264.900 ;
        RECT 178.950 264.450 181.050 265.050 ;
        RECT 184.950 264.450 187.050 265.050 ;
        RECT 149.100 259.050 150.900 260.850 ;
        RECT 155.100 259.050 156.900 260.850 ;
        RECT 158.100 259.050 159.000 262.800 ;
        RECT 170.250 259.050 172.050 260.850 ;
        RECT 88.950 256.950 91.050 259.050 ;
        RECT 91.950 256.950 94.050 259.050 ;
        RECT 94.950 256.950 97.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 109.950 256.950 112.050 259.050 ;
        RECT 112.950 256.950 115.050 259.050 ;
        RECT 121.950 256.950 124.050 259.050 ;
        RECT 124.950 256.950 127.050 259.050 ;
        RECT 127.950 256.950 130.050 259.050 ;
        RECT 130.950 256.950 133.050 259.050 ;
        RECT 139.950 256.950 142.050 259.050 ;
        RECT 142.950 256.950 145.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 151.950 256.950 154.050 259.050 ;
        RECT 154.950 256.950 157.050 259.050 ;
        RECT 157.950 256.950 160.050 259.050 ;
        RECT 166.950 256.950 169.050 259.050 ;
        RECT 169.950 256.950 172.050 259.050 ;
        RECT 172.950 259.050 174.000 263.700 ;
        RECT 178.950 263.550 187.050 264.450 ;
        RECT 188.700 264.300 192.900 265.200 ;
        RECT 178.950 262.950 181.050 263.550 ;
        RECT 184.950 262.950 187.050 263.550 ;
        RECT 175.950 259.050 177.750 260.850 ;
        RECT 188.100 259.050 189.900 260.850 ;
        RECT 191.700 259.050 192.900 264.300 ;
        RECT 193.950 259.050 195.750 260.850 ;
        RECT 200.700 259.050 201.900 269.400 ;
        RECT 212.100 264.600 213.900 272.400 ;
        RECT 216.600 266.400 218.400 273.000 ;
        RECT 219.600 268.200 221.400 272.400 ;
        RECT 219.600 266.400 222.300 268.200 ;
        RECT 227.400 266.400 229.200 273.000 ;
        RECT 218.700 264.600 220.500 265.500 ;
        RECT 212.100 263.700 220.500 264.600 ;
        RECT 205.950 261.450 210.000 262.050 ;
        RECT 205.950 259.950 210.450 261.450 ;
        RECT 172.950 256.950 175.050 259.050 ;
        RECT 175.950 256.950 178.050 259.050 ;
        RECT 178.950 256.950 181.050 259.050 ;
        RECT 187.950 256.950 190.050 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 193.950 256.950 196.050 259.050 ;
        RECT 199.950 256.950 202.050 259.050 ;
        RECT 202.950 256.950 205.050 259.050 ;
        RECT 79.500 253.950 81.900 256.050 ;
        RECT 73.800 243.600 75.000 244.500 ;
        RECT 79.500 243.600 81.000 253.950 ;
        RECT 92.100 243.600 93.300 256.950 ;
        RECT 107.100 249.600 108.300 256.950 ;
        RECT 113.100 255.150 114.900 256.950 ;
        RECT 122.400 249.600 123.300 256.950 ;
        RECT 127.950 255.150 129.750 256.950 ;
        RECT 107.100 248.100 109.500 249.600 ;
        RECT 105.000 245.100 106.800 246.900 ;
        RECT 49.200 237.000 51.000 243.600 ;
        RECT 52.200 237.600 54.000 243.600 ;
        RECT 55.200 240.600 57.300 242.700 ;
        RECT 58.200 240.600 60.300 242.700 ;
        RECT 61.200 240.600 63.300 242.700 ;
        RECT 55.200 237.600 57.000 240.600 ;
        RECT 58.200 237.600 60.000 240.600 ;
        RECT 61.200 237.600 63.000 240.600 ;
        RECT 64.200 237.000 66.000 243.600 ;
        RECT 67.200 237.600 69.000 243.600 ;
        RECT 70.200 237.000 72.000 243.600 ;
        RECT 73.200 237.600 75.000 243.600 ;
        RECT 76.200 237.000 78.000 243.600 ;
        RECT 79.500 237.600 81.300 243.600 ;
        RECT 82.500 237.000 84.300 243.600 ;
        RECT 89.100 237.000 90.900 243.600 ;
        RECT 92.100 237.600 93.900 243.600 ;
        RECT 95.100 237.000 96.900 243.600 ;
        RECT 104.700 237.000 106.500 243.600 ;
        RECT 107.700 237.600 109.500 248.100 ;
        RECT 112.800 237.000 114.600 249.600 ;
        RECT 122.100 237.600 123.900 249.600 ;
        RECT 125.100 248.700 132.900 249.600 ;
        RECT 125.100 237.600 126.900 248.700 ;
        RECT 128.100 237.000 129.900 247.800 ;
        RECT 131.100 237.600 132.900 248.700 ;
        RECT 140.700 243.600 141.900 256.950 ;
        RECT 143.100 255.150 144.900 256.950 ;
        RECT 152.100 255.150 153.900 256.950 ;
        RECT 158.100 244.800 159.000 256.950 ;
        RECT 167.100 255.150 168.900 256.950 ;
        RECT 172.950 249.600 174.000 256.950 ;
        RECT 178.950 255.150 180.750 256.950 ;
        RECT 152.400 243.900 159.000 244.800 ;
        RECT 152.400 243.600 153.900 243.900 ;
        RECT 140.100 237.600 141.900 243.600 ;
        RECT 143.100 237.000 144.900 243.600 ;
        RECT 149.100 237.000 150.900 243.600 ;
        RECT 152.100 237.600 153.900 243.600 ;
        RECT 158.100 243.600 159.000 243.900 ;
        RECT 155.100 237.000 156.900 243.000 ;
        RECT 158.100 237.600 159.900 243.600 ;
        RECT 167.100 237.000 168.900 249.600 ;
        RECT 171.600 237.600 174.900 249.600 ;
        RECT 177.600 237.000 179.400 249.600 ;
        RECT 191.700 243.600 192.900 256.950 ;
        RECT 200.700 243.600 201.900 256.950 ;
        RECT 203.100 255.150 204.900 256.950 ;
        RECT 202.950 252.450 205.050 253.050 ;
        RECT 209.550 252.450 210.450 259.950 ;
        RECT 212.250 259.050 214.050 260.850 ;
        RECT 212.100 256.950 214.200 259.050 ;
        RECT 202.950 251.550 210.450 252.450 ;
        RECT 202.950 250.950 205.050 251.550 ;
        RECT 215.100 243.600 216.000 263.700 ;
        RECT 221.400 259.050 222.300 266.400 ;
        RECT 232.500 265.200 234.300 272.400 ;
        RECT 230.100 264.300 234.300 265.200 ;
        RECT 239.100 266.400 240.900 272.400 ;
        RECT 242.100 266.400 243.900 273.000 ;
        RECT 245.100 269.400 246.900 272.400 ;
        RECT 254.100 269.400 255.900 273.000 ;
        RECT 257.100 269.400 258.900 272.400 ;
        RECT 263.100 269.400 264.900 273.000 ;
        RECT 266.100 269.400 267.900 272.400 ;
        RECT 227.250 259.050 229.050 260.850 ;
        RECT 230.100 259.050 231.300 264.300 ;
        RECT 233.100 259.050 234.900 260.850 ;
        RECT 239.100 259.050 240.300 266.400 ;
        RECT 245.700 265.500 246.900 269.400 ;
        RECT 241.200 264.600 246.900 265.500 ;
        RECT 241.200 263.700 243.000 264.600 ;
        RECT 217.500 256.950 219.600 259.050 ;
        RECT 220.800 256.950 222.900 259.050 ;
        RECT 226.950 256.950 229.050 259.050 ;
        RECT 229.950 256.950 232.050 259.050 ;
        RECT 232.950 256.950 235.050 259.050 ;
        RECT 239.100 256.950 241.200 259.050 ;
        RECT 217.200 255.150 219.000 256.950 ;
        RECT 221.400 249.600 222.300 256.950 ;
        RECT 188.100 237.000 189.900 243.600 ;
        RECT 191.100 237.600 192.900 243.600 ;
        RECT 194.100 237.000 195.900 243.600 ;
        RECT 200.100 237.600 201.900 243.600 ;
        RECT 203.100 237.000 204.900 243.600 ;
        RECT 212.100 237.000 213.900 243.600 ;
        RECT 215.100 237.600 216.900 243.600 ;
        RECT 218.100 237.000 219.900 249.000 ;
        RECT 221.100 237.600 222.900 249.600 ;
        RECT 230.100 243.600 231.300 256.950 ;
        RECT 239.100 249.600 240.300 256.950 ;
        RECT 242.100 252.300 243.000 263.700 ;
        RECT 257.100 259.050 258.300 269.400 ;
        RECT 266.100 259.050 267.300 269.400 ;
        RECT 272.400 266.400 274.200 273.000 ;
        RECT 277.500 265.200 279.300 272.400 ;
        RECT 275.100 264.300 279.300 265.200 ;
        RECT 287.700 265.200 289.500 272.400 ;
        RECT 292.800 266.400 294.600 273.000 ;
        RECT 287.700 264.300 291.900 265.200 ;
        RECT 272.250 259.050 274.050 260.850 ;
        RECT 275.100 259.050 276.300 264.300 ;
        RECT 278.100 259.050 279.900 260.850 ;
        RECT 287.100 259.050 288.900 260.850 ;
        RECT 290.700 259.050 291.900 264.300 ;
        RECT 296.100 263.400 297.900 273.000 ;
        RECT 302.700 264.000 304.500 272.400 ;
        RECT 311.100 267.300 312.900 272.400 ;
        RECT 314.100 268.200 315.900 273.000 ;
        RECT 317.100 267.300 318.900 272.400 ;
        RECT 311.100 265.950 318.900 267.300 ;
        RECT 320.100 266.400 321.900 272.400 ;
        RECT 330.000 266.400 331.800 273.000 ;
        RECT 334.500 267.600 336.300 272.400 ;
        RECT 337.500 269.400 339.300 273.000 ;
        RECT 334.500 266.400 339.600 267.600 ;
        RECT 320.100 264.300 321.300 266.400 ;
        RECT 302.700 262.800 306.000 264.000 ;
        RECT 292.950 259.050 294.750 260.850 ;
        RECT 296.100 259.050 297.900 260.850 ;
        RECT 302.100 259.050 303.900 260.850 ;
        RECT 305.100 259.050 306.000 262.800 ;
        RECT 317.700 263.400 321.300 264.300 ;
        RECT 314.100 259.050 315.900 260.850 ;
        RECT 317.700 259.050 318.900 263.400 ;
        RECT 320.100 259.050 321.900 260.850 ;
        RECT 329.100 259.050 330.900 260.850 ;
        RECT 335.250 259.050 337.050 260.850 ;
        RECT 338.700 259.050 339.600 266.400 ;
        RECT 347.100 267.000 348.900 272.400 ;
        RECT 350.100 267.900 351.900 273.000 ;
        RECT 353.100 271.500 360.900 272.400 ;
        RECT 353.100 267.000 354.900 271.500 ;
        RECT 347.100 266.100 354.900 267.000 ;
        RECT 356.100 266.400 357.900 270.600 ;
        RECT 359.100 266.400 360.900 271.500 ;
        RECT 356.400 264.900 357.300 266.400 ;
        RECT 352.950 263.700 357.300 264.900 ;
        RECT 350.250 259.050 352.050 260.850 ;
        RECT 244.500 256.950 246.600 259.050 ;
        RECT 253.950 256.950 256.050 259.050 ;
        RECT 256.950 256.950 259.050 259.050 ;
        RECT 262.950 256.950 265.050 259.050 ;
        RECT 265.950 256.950 268.050 259.050 ;
        RECT 271.950 256.950 274.050 259.050 ;
        RECT 274.950 256.950 277.050 259.050 ;
        RECT 277.950 256.950 280.050 259.050 ;
        RECT 286.950 256.950 289.050 259.050 ;
        RECT 289.950 256.950 292.050 259.050 ;
        RECT 292.950 256.950 295.050 259.050 ;
        RECT 295.950 256.950 298.050 259.050 ;
        RECT 298.950 256.950 301.050 259.050 ;
        RECT 301.950 256.950 304.050 259.050 ;
        RECT 304.950 256.950 307.050 259.050 ;
        RECT 310.950 256.950 313.050 259.050 ;
        RECT 313.950 256.950 316.050 259.050 ;
        RECT 316.950 256.950 319.050 259.050 ;
        RECT 319.950 256.950 322.050 259.050 ;
        RECT 328.950 256.950 331.050 259.050 ;
        RECT 331.950 256.950 334.050 259.050 ;
        RECT 334.950 256.950 337.050 259.050 ;
        RECT 337.950 256.950 340.050 259.050 ;
        RECT 346.950 256.950 349.050 259.050 ;
        RECT 349.950 256.950 352.050 259.050 ;
        RECT 352.950 259.050 354.000 263.700 ;
        RECT 355.950 259.050 357.750 260.850 ;
        RECT 352.950 256.950 355.050 259.050 ;
        RECT 355.950 256.950 358.050 259.050 ;
        RECT 358.950 256.950 361.050 259.050 ;
        RECT 244.800 255.150 246.600 256.950 ;
        RECT 254.100 255.150 255.900 256.950 ;
        RECT 241.200 251.400 243.000 252.300 ;
        RECT 241.200 250.500 246.900 251.400 ;
        RECT 227.100 237.000 228.900 243.600 ;
        RECT 230.100 237.600 231.900 243.600 ;
        RECT 233.100 237.000 234.900 243.600 ;
        RECT 239.100 237.600 240.900 249.600 ;
        RECT 242.100 237.000 243.900 247.800 ;
        RECT 245.700 243.600 246.900 250.500 ;
        RECT 257.100 243.600 258.300 256.950 ;
        RECT 263.100 255.150 264.900 256.950 ;
        RECT 266.100 243.600 267.300 256.950 ;
        RECT 275.100 243.600 276.300 256.950 ;
        RECT 280.950 252.450 283.050 253.050 ;
        RECT 286.950 252.450 289.050 253.050 ;
        RECT 280.950 251.550 289.050 252.450 ;
        RECT 280.950 250.950 283.050 251.550 ;
        RECT 286.950 250.950 289.050 251.550 ;
        RECT 290.700 243.600 291.900 256.950 ;
        RECT 299.100 255.150 300.900 256.950 ;
        RECT 305.100 244.800 306.000 256.950 ;
        RECT 311.100 255.150 312.900 256.950 ;
        RECT 317.700 249.600 318.900 256.950 ;
        RECT 332.250 255.150 334.050 256.950 ;
        RECT 338.700 249.600 339.600 256.950 ;
        RECT 347.100 255.150 348.900 256.950 ;
        RECT 352.950 249.600 354.000 256.950 ;
        RECT 358.950 255.150 360.750 256.950 ;
        RECT 299.400 243.900 306.000 244.800 ;
        RECT 299.400 243.600 300.900 243.900 ;
        RECT 245.100 237.600 246.900 243.600 ;
        RECT 254.100 237.000 255.900 243.600 ;
        RECT 257.100 237.600 258.900 243.600 ;
        RECT 263.100 237.000 264.900 243.600 ;
        RECT 266.100 237.600 267.900 243.600 ;
        RECT 272.100 237.000 273.900 243.600 ;
        RECT 275.100 237.600 276.900 243.600 ;
        RECT 278.100 237.000 279.900 243.600 ;
        RECT 287.100 237.000 288.900 243.600 ;
        RECT 290.100 237.600 291.900 243.600 ;
        RECT 293.100 237.000 294.900 243.600 ;
        RECT 296.100 237.000 297.900 243.600 ;
        RECT 299.100 237.600 300.900 243.600 ;
        RECT 305.100 243.600 306.000 243.900 ;
        RECT 302.100 237.000 303.900 243.000 ;
        RECT 305.100 237.600 306.900 243.600 ;
        RECT 311.400 237.000 313.200 249.600 ;
        RECT 316.500 248.100 318.900 249.600 ;
        RECT 329.100 248.700 336.900 249.600 ;
        RECT 316.500 237.600 318.300 248.100 ;
        RECT 319.200 245.100 321.000 246.900 ;
        RECT 319.500 237.000 321.300 243.600 ;
        RECT 329.100 237.600 330.900 248.700 ;
        RECT 332.100 237.000 333.900 247.800 ;
        RECT 335.100 237.600 336.900 248.700 ;
        RECT 338.100 237.600 339.900 249.600 ;
        RECT 347.100 237.000 348.900 249.600 ;
        RECT 351.600 237.600 354.900 249.600 ;
        RECT 357.600 237.000 359.400 249.600 ;
        RECT 8.100 227.400 9.900 233.400 ;
        RECT 11.100 227.400 12.900 234.000 ;
        RECT 8.700 214.050 9.900 227.400 ;
        RECT 17.100 221.400 18.900 233.400 ;
        RECT 20.100 222.000 21.900 234.000 ;
        RECT 23.100 227.400 24.900 233.400 ;
        RECT 26.100 227.400 27.900 234.000 ;
        RECT 11.100 214.050 12.900 215.850 ;
        RECT 17.700 214.050 18.600 221.400 ;
        RECT 21.000 214.050 22.800 215.850 ;
        RECT 7.950 211.950 10.050 214.050 ;
        RECT 10.950 211.950 13.050 214.050 ;
        RECT 17.100 211.950 19.200 214.050 ;
        RECT 20.400 211.950 22.500 214.050 ;
        RECT 8.700 201.600 9.900 211.950 ;
        RECT 17.700 204.600 18.600 211.950 ;
        RECT 24.000 207.300 24.900 227.400 ;
        RECT 35.400 221.400 37.200 234.000 ;
        RECT 40.500 222.900 42.300 233.400 ;
        RECT 43.500 227.400 45.300 234.000 ;
        RECT 43.200 224.100 45.000 225.900 ;
        RECT 40.500 221.400 42.900 222.900 ;
        RECT 53.400 221.400 55.200 234.000 ;
        RECT 58.500 222.900 60.300 233.400 ;
        RECT 61.500 227.400 63.300 234.000 ;
        RECT 61.200 224.100 63.000 225.900 ;
        RECT 58.500 221.400 60.900 222.900 ;
        RECT 71.100 221.400 72.900 234.000 ;
        RECT 76.200 222.600 78.000 233.400 ;
        RECT 74.400 221.400 78.000 222.600 ;
        RECT 83.100 221.400 84.900 233.400 ;
        RECT 86.100 222.000 87.900 234.000 ;
        RECT 89.100 227.400 90.900 233.400 ;
        RECT 92.100 227.400 93.900 234.000 ;
        RECT 98.100 227.400 99.900 233.400 ;
        RECT 101.100 228.000 102.900 234.000 ;
        RECT 30.000 216.450 34.050 217.050 ;
        RECT 29.550 214.950 34.050 216.450 ;
        RECT 25.800 211.950 27.900 214.050 ;
        RECT 25.950 210.150 27.750 211.950 ;
        RECT 29.550 210.900 30.450 214.950 ;
        RECT 35.100 214.050 36.900 215.850 ;
        RECT 41.700 214.050 42.900 221.400 ;
        RECT 53.100 214.050 54.900 215.850 ;
        RECT 59.700 214.050 60.900 221.400 ;
        RECT 71.250 214.050 73.050 215.850 ;
        RECT 74.400 214.050 75.300 221.400 ;
        RECT 77.100 214.050 78.900 215.850 ;
        RECT 83.700 214.050 84.600 221.400 ;
        RECT 87.000 214.050 88.800 215.850 ;
        RECT 34.950 211.950 37.050 214.050 ;
        RECT 37.950 211.950 40.050 214.050 ;
        RECT 40.950 211.950 43.050 214.050 ;
        RECT 43.950 211.950 46.050 214.050 ;
        RECT 52.950 211.950 55.050 214.050 ;
        RECT 55.950 211.950 58.050 214.050 ;
        RECT 58.950 211.950 61.050 214.050 ;
        RECT 61.950 211.950 64.050 214.050 ;
        RECT 70.950 211.950 73.050 214.050 ;
        RECT 73.950 211.950 76.050 214.050 ;
        RECT 76.950 211.950 79.050 214.050 ;
        RECT 83.100 211.950 85.200 214.050 ;
        RECT 86.400 211.950 88.500 214.050 ;
        RECT 28.950 208.800 31.050 210.900 ;
        RECT 38.100 210.150 39.900 211.950 ;
        RECT 41.700 207.600 42.900 211.950 ;
        RECT 44.100 210.150 45.900 211.950 ;
        RECT 56.100 210.150 57.900 211.950 ;
        RECT 59.700 207.600 60.900 211.950 ;
        RECT 62.100 210.150 63.900 211.950 ;
        RECT 19.500 206.400 27.900 207.300 ;
        RECT 41.700 206.700 45.300 207.600 ;
        RECT 59.700 206.700 63.300 207.600 ;
        RECT 19.500 205.500 21.300 206.400 ;
        RECT 17.700 202.800 20.400 204.600 ;
        RECT 8.100 198.600 9.900 201.600 ;
        RECT 11.100 198.000 12.900 201.600 ;
        RECT 18.600 198.600 20.400 202.800 ;
        RECT 21.600 198.000 23.400 204.600 ;
        RECT 26.100 198.600 27.900 206.400 ;
        RECT 35.100 203.700 42.900 205.050 ;
        RECT 35.100 198.600 36.900 203.700 ;
        RECT 38.100 198.000 39.900 202.800 ;
        RECT 41.100 198.600 42.900 203.700 ;
        RECT 44.100 204.600 45.300 206.700 ;
        RECT 44.100 198.600 45.900 204.600 ;
        RECT 53.100 203.700 60.900 205.050 ;
        RECT 53.100 198.600 54.900 203.700 ;
        RECT 56.100 198.000 57.900 202.800 ;
        RECT 59.100 198.600 60.900 203.700 ;
        RECT 62.100 204.600 63.300 206.700 ;
        RECT 64.950 207.450 67.050 208.050 ;
        RECT 70.950 207.450 73.050 208.050 ;
        RECT 64.950 206.550 73.050 207.450 ;
        RECT 64.950 205.950 67.050 206.550 ;
        RECT 70.950 205.950 73.050 206.550 ;
        RECT 62.100 198.600 63.900 204.600 ;
        RECT 74.400 201.600 75.300 211.950 ;
        RECT 83.700 204.600 84.600 211.950 ;
        RECT 90.000 207.300 90.900 227.400 ;
        RECT 99.000 227.100 99.900 227.400 ;
        RECT 104.100 227.400 105.900 233.400 ;
        RECT 107.100 227.400 108.900 234.000 ;
        RECT 104.100 227.100 105.600 227.400 ;
        RECT 99.000 226.200 105.600 227.100 ;
        RECT 113.100 226.200 114.900 232.200 ;
        RECT 99.000 214.050 99.900 226.200 ;
        RECT 113.100 221.100 114.000 226.200 ;
        RECT 116.100 222.000 117.900 234.000 ;
        RECT 120.600 222.900 122.400 233.400 ;
        RECT 120.600 222.000 122.700 222.900 ;
        RECT 113.100 220.200 120.900 221.100 ;
        RECT 119.700 215.850 120.900 220.200 ;
        RECT 104.100 214.050 105.900 215.850 ;
        RECT 116.100 214.050 117.900 215.850 ;
        RECT 119.100 214.050 120.900 215.850 ;
        RECT 121.800 214.050 122.700 222.000 ;
        RECT 125.100 221.400 126.900 234.000 ;
        RECT 134.100 227.400 135.900 234.000 ;
        RECT 137.100 227.400 138.900 233.400 ;
        RECT 140.100 227.400 141.900 234.000 ;
        RECT 143.100 227.400 144.900 234.000 ;
        RECT 146.100 227.400 147.900 233.400 ;
        RECT 129.000 216.450 133.050 217.050 ;
        RECT 124.800 214.050 126.600 215.850 ;
        RECT 128.550 214.950 133.050 216.450 ;
        RECT 91.800 211.950 93.900 214.050 ;
        RECT 97.950 211.950 100.050 214.050 ;
        RECT 100.950 211.950 103.050 214.050 ;
        RECT 103.950 211.950 106.050 214.050 ;
        RECT 106.950 211.950 109.050 214.050 ;
        RECT 113.100 211.950 115.200 214.050 ;
        RECT 116.100 211.950 118.200 214.050 ;
        RECT 91.950 210.150 93.750 211.950 ;
        RECT 99.000 208.200 99.900 211.950 ;
        RECT 101.100 210.150 102.900 211.950 ;
        RECT 107.100 210.150 108.900 211.950 ;
        RECT 113.100 210.150 114.900 211.950 ;
        RECT 85.500 206.400 93.900 207.300 ;
        RECT 99.000 207.000 102.300 208.200 ;
        RECT 85.500 205.500 87.300 206.400 ;
        RECT 83.700 202.800 86.400 204.600 ;
        RECT 71.100 198.000 72.900 201.600 ;
        RECT 74.100 198.600 75.900 201.600 ;
        RECT 77.100 198.000 78.900 201.600 ;
        RECT 84.600 198.600 86.400 202.800 ;
        RECT 87.600 198.000 89.400 204.600 ;
        RECT 92.100 198.600 93.900 206.400 ;
        RECT 100.500 198.600 102.300 207.000 ;
        RECT 107.100 198.000 108.900 207.600 ;
        RECT 119.100 207.000 120.300 214.050 ;
        RECT 113.100 206.100 120.300 207.000 ;
        RECT 121.800 211.950 123.900 214.050 ;
        RECT 124.800 211.950 126.900 214.050 ;
        RECT 113.100 202.800 114.000 206.100 ;
        RECT 121.800 205.200 122.700 211.950 ;
        RECT 128.550 211.050 129.450 214.950 ;
        RECT 137.700 214.050 138.900 227.400 ;
        RECT 133.950 211.950 136.050 214.050 ;
        RECT 136.950 211.950 139.050 214.050 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 143.100 211.950 145.200 214.050 ;
        RECT 128.550 209.550 133.050 211.050 ;
        RECT 134.100 210.150 135.900 211.950 ;
        RECT 129.000 208.950 133.050 209.550 ;
        RECT 137.700 206.700 138.900 211.950 ;
        RECT 139.950 210.150 141.750 211.950 ;
        RECT 143.250 210.150 145.050 211.950 ;
        RECT 146.100 207.300 147.000 227.400 ;
        RECT 149.100 222.000 150.900 234.000 ;
        RECT 152.100 221.400 153.900 233.400 ;
        RECT 158.100 221.400 159.900 233.400 ;
        RECT 161.100 222.000 162.900 234.000 ;
        RECT 164.100 227.400 165.900 233.400 ;
        RECT 167.100 227.400 168.900 234.000 ;
        RECT 148.200 214.050 150.000 215.850 ;
        RECT 152.400 214.050 153.300 221.400 ;
        RECT 158.700 214.050 159.600 221.400 ;
        RECT 162.000 214.050 163.800 215.850 ;
        RECT 148.500 211.950 150.600 214.050 ;
        RECT 151.800 211.950 153.900 214.050 ;
        RECT 158.100 211.950 160.200 214.050 ;
        RECT 161.400 211.950 163.500 214.050 ;
        RECT 134.700 205.800 138.900 206.700 ;
        RECT 143.100 206.400 151.500 207.300 ;
        RECT 113.100 199.800 114.900 202.800 ;
        RECT 116.100 200.400 117.900 205.200 ;
        RECT 120.600 204.300 122.700 205.200 ;
        RECT 116.100 198.000 117.300 200.400 ;
        RECT 120.600 199.800 122.400 204.300 ;
        RECT 125.100 199.800 126.900 205.800 ;
        RECT 125.100 198.000 126.300 199.800 ;
        RECT 134.700 198.600 136.500 205.800 ;
        RECT 139.800 198.000 141.600 204.600 ;
        RECT 143.100 198.600 144.900 206.400 ;
        RECT 149.700 205.500 151.500 206.400 ;
        RECT 152.400 204.600 153.300 211.950 ;
        RECT 147.600 198.000 149.400 204.600 ;
        RECT 150.600 202.800 153.300 204.600 ;
        RECT 158.700 204.600 159.600 211.950 ;
        RECT 165.000 207.300 165.900 227.400 ;
        RECT 177.000 222.600 178.800 233.400 ;
        RECT 177.000 221.400 180.600 222.600 ;
        RECT 182.100 221.400 183.900 234.000 ;
        RECT 191.100 227.400 192.900 234.000 ;
        RECT 194.100 227.400 195.900 233.400 ;
        RECT 176.100 214.050 177.900 215.850 ;
        RECT 179.700 214.050 180.600 221.400 ;
        RECT 181.950 214.050 183.750 215.850 ;
        RECT 166.800 211.950 168.900 214.050 ;
        RECT 175.950 211.950 178.050 214.050 ;
        RECT 178.950 211.950 181.050 214.050 ;
        RECT 181.950 211.950 184.050 214.050 ;
        RECT 191.100 211.950 193.200 214.050 ;
        RECT 166.950 210.150 168.750 211.950 ;
        RECT 169.950 207.450 172.050 208.050 ;
        RECT 175.950 207.450 178.050 208.050 ;
        RECT 160.500 206.400 168.900 207.300 ;
        RECT 160.500 205.500 162.300 206.400 ;
        RECT 158.700 202.800 161.400 204.600 ;
        RECT 150.600 198.600 152.400 202.800 ;
        RECT 159.600 198.600 161.400 202.800 ;
        RECT 162.600 198.000 164.400 204.600 ;
        RECT 167.100 198.600 168.900 206.400 ;
        RECT 169.950 206.550 178.050 207.450 ;
        RECT 169.950 205.950 172.050 206.550 ;
        RECT 175.950 205.950 178.050 206.550 ;
        RECT 179.700 201.600 180.600 211.950 ;
        RECT 191.250 210.150 193.050 211.950 ;
        RECT 194.100 207.300 195.000 227.400 ;
        RECT 197.100 222.000 198.900 234.000 ;
        RECT 200.100 221.400 201.900 233.400 ;
        RECT 209.100 227.400 210.900 233.400 ;
        RECT 212.100 227.400 213.900 234.000 ;
        RECT 196.200 214.050 198.000 215.850 ;
        RECT 200.400 214.050 201.300 221.400 ;
        RECT 209.700 214.050 210.900 227.400 ;
        RECT 218.400 221.400 220.200 234.000 ;
        RECT 223.500 222.900 225.300 233.400 ;
        RECT 226.500 227.400 228.300 234.000 ;
        RECT 236.100 227.400 237.900 234.000 ;
        RECT 239.100 227.400 240.900 233.400 ;
        RECT 242.100 228.000 243.900 234.000 ;
        RECT 239.400 227.100 240.900 227.400 ;
        RECT 245.100 227.400 246.900 233.400 ;
        RECT 254.100 227.400 255.900 234.000 ;
        RECT 257.100 227.400 258.900 233.400 ;
        RECT 245.100 227.100 246.000 227.400 ;
        RECT 239.400 226.200 246.000 227.100 ;
        RECT 226.200 224.100 228.000 225.900 ;
        RECT 223.500 221.400 225.900 222.900 ;
        RECT 214.950 219.450 217.050 220.050 ;
        RECT 220.950 219.450 223.050 220.200 ;
        RECT 214.950 218.550 223.050 219.450 ;
        RECT 214.950 217.950 217.050 218.550 ;
        RECT 220.950 218.100 223.050 218.550 ;
        RECT 212.100 214.050 213.900 215.850 ;
        RECT 218.100 214.050 219.900 215.850 ;
        RECT 224.700 214.050 225.900 221.400 ;
        RECT 239.100 214.050 240.900 215.850 ;
        RECT 245.100 214.050 246.000 226.200 ;
        RECT 196.500 211.950 198.600 214.050 ;
        RECT 199.800 211.950 201.900 214.050 ;
        RECT 208.950 211.950 211.050 214.050 ;
        RECT 211.950 211.950 214.050 214.050 ;
        RECT 217.950 211.950 220.050 214.050 ;
        RECT 220.950 211.950 223.050 214.050 ;
        RECT 223.950 211.950 226.050 214.050 ;
        RECT 226.950 211.950 229.050 214.050 ;
        RECT 235.950 211.950 238.050 214.050 ;
        RECT 238.950 211.950 241.050 214.050 ;
        RECT 241.950 211.950 244.050 214.050 ;
        RECT 244.950 211.950 247.050 214.050 ;
        RECT 254.100 211.950 256.200 214.050 ;
        RECT 191.100 206.400 199.500 207.300 ;
        RECT 176.100 198.000 177.900 201.600 ;
        RECT 179.100 198.600 180.900 201.600 ;
        RECT 182.100 198.000 183.900 201.600 ;
        RECT 191.100 198.600 192.900 206.400 ;
        RECT 197.700 205.500 199.500 206.400 ;
        RECT 200.400 204.600 201.300 211.950 ;
        RECT 195.600 198.000 197.400 204.600 ;
        RECT 198.600 202.800 201.300 204.600 ;
        RECT 198.600 198.600 200.400 202.800 ;
        RECT 209.700 201.600 210.900 211.950 ;
        RECT 221.100 210.150 222.900 211.950 ;
        RECT 224.700 207.600 225.900 211.950 ;
        RECT 227.100 210.150 228.900 211.950 ;
        RECT 236.100 210.150 237.900 211.950 ;
        RECT 242.100 210.150 243.900 211.950 ;
        RECT 245.100 208.200 246.000 211.950 ;
        RECT 254.250 210.150 256.050 211.950 ;
        RECT 224.700 206.700 228.300 207.600 ;
        RECT 218.100 203.700 225.900 205.050 ;
        RECT 209.100 198.600 210.900 201.600 ;
        RECT 212.100 198.000 213.900 201.600 ;
        RECT 218.100 198.600 219.900 203.700 ;
        RECT 221.100 198.000 222.900 202.800 ;
        RECT 224.100 198.600 225.900 203.700 ;
        RECT 227.100 204.600 228.300 206.700 ;
        RECT 227.100 198.600 228.900 204.600 ;
        RECT 236.100 198.000 237.900 207.600 ;
        RECT 242.700 207.000 246.000 208.200 ;
        RECT 257.100 207.300 258.000 227.400 ;
        RECT 260.100 222.000 261.900 234.000 ;
        RECT 263.100 221.400 264.900 233.400 ;
        RECT 269.400 221.400 271.200 234.000 ;
        RECT 274.500 222.900 276.300 233.400 ;
        RECT 277.500 227.400 279.300 234.000 ;
        RECT 287.100 227.400 288.900 233.400 ;
        RECT 290.100 228.000 291.900 234.000 ;
        RECT 288.000 227.100 288.900 227.400 ;
        RECT 293.100 227.400 294.900 233.400 ;
        RECT 296.100 227.400 297.900 234.000 ;
        RECT 302.100 227.400 303.900 233.400 ;
        RECT 305.100 227.400 306.900 234.000 ;
        RECT 314.100 227.400 315.900 234.000 ;
        RECT 317.100 227.400 318.900 233.400 ;
        RECT 323.700 227.400 325.500 234.000 ;
        RECT 293.100 227.100 294.600 227.400 ;
        RECT 288.000 226.200 294.600 227.100 ;
        RECT 277.200 224.100 279.000 225.900 ;
        RECT 274.500 221.400 276.900 222.900 ;
        RECT 259.200 214.050 261.000 215.850 ;
        RECT 263.400 214.050 264.300 221.400 ;
        RECT 269.100 214.050 270.900 215.850 ;
        RECT 275.700 214.050 276.900 221.400 ;
        RECT 288.000 214.050 288.900 226.200 ;
        RECT 293.100 214.050 294.900 215.850 ;
        RECT 302.700 214.050 303.900 227.400 ;
        RECT 305.100 214.050 306.900 215.850 ;
        RECT 314.100 214.050 315.900 215.850 ;
        RECT 317.100 214.050 318.300 227.400 ;
        RECT 324.000 224.100 325.800 225.900 ;
        RECT 326.700 222.900 328.500 233.400 ;
        RECT 326.100 221.400 328.500 222.900 ;
        RECT 331.800 221.400 333.600 234.000 ;
        RECT 341.100 227.400 342.900 233.400 ;
        RECT 344.100 227.400 345.900 234.000 ;
        RECT 350.100 227.400 351.900 233.400 ;
        RECT 353.100 228.000 354.900 234.000 ;
        RECT 326.100 214.050 327.300 221.400 ;
        RECT 332.100 214.050 333.900 215.850 ;
        RECT 341.700 214.050 342.900 227.400 ;
        RECT 351.000 227.100 351.900 227.400 ;
        RECT 356.100 227.400 357.900 233.400 ;
        RECT 359.100 227.400 360.900 234.000 ;
        RECT 356.100 227.100 357.600 227.400 ;
        RECT 351.000 226.200 357.600 227.100 ;
        RECT 344.100 214.050 345.900 215.850 ;
        RECT 351.000 214.050 351.900 226.200 ;
        RECT 356.100 214.050 357.900 215.850 ;
        RECT 259.500 211.950 261.600 214.050 ;
        RECT 262.800 211.950 264.900 214.050 ;
        RECT 268.950 211.950 271.050 214.050 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 277.950 211.950 280.050 214.050 ;
        RECT 286.950 211.950 289.050 214.050 ;
        RECT 289.950 211.950 292.050 214.050 ;
        RECT 292.950 211.950 295.050 214.050 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 301.950 211.950 304.050 214.050 ;
        RECT 304.950 211.950 307.050 214.050 ;
        RECT 313.950 211.950 316.050 214.050 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 322.950 211.950 325.050 214.050 ;
        RECT 325.950 211.950 328.050 214.050 ;
        RECT 328.950 211.950 331.050 214.050 ;
        RECT 331.950 211.950 334.050 214.050 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 343.950 211.950 346.050 214.050 ;
        RECT 349.950 211.950 352.050 214.050 ;
        RECT 352.950 211.950 355.050 214.050 ;
        RECT 355.950 211.950 358.050 214.050 ;
        RECT 358.950 211.950 361.050 214.050 ;
        RECT 242.700 198.600 244.500 207.000 ;
        RECT 254.100 206.400 262.500 207.300 ;
        RECT 254.100 198.600 255.900 206.400 ;
        RECT 260.700 205.500 262.500 206.400 ;
        RECT 263.400 204.600 264.300 211.950 ;
        RECT 272.100 210.150 273.900 211.950 ;
        RECT 275.700 207.600 276.900 211.950 ;
        RECT 278.100 210.150 279.900 211.950 ;
        RECT 288.000 208.200 288.900 211.950 ;
        RECT 290.100 210.150 291.900 211.950 ;
        RECT 296.100 210.150 297.900 211.950 ;
        RECT 275.700 206.700 279.300 207.600 ;
        RECT 288.000 207.000 291.300 208.200 ;
        RECT 258.600 198.000 260.400 204.600 ;
        RECT 261.600 202.800 264.300 204.600 ;
        RECT 269.100 203.700 276.900 205.050 ;
        RECT 261.600 198.600 263.400 202.800 ;
        RECT 269.100 198.600 270.900 203.700 ;
        RECT 272.100 198.000 273.900 202.800 ;
        RECT 275.100 198.600 276.900 203.700 ;
        RECT 278.100 204.600 279.300 206.700 ;
        RECT 278.100 198.600 279.900 204.600 ;
        RECT 289.500 198.600 291.300 207.000 ;
        RECT 296.100 198.000 297.900 207.600 ;
        RECT 302.700 201.600 303.900 211.950 ;
        RECT 317.100 201.600 318.300 211.950 ;
        RECT 323.100 210.150 324.900 211.950 ;
        RECT 326.100 207.600 327.300 211.950 ;
        RECT 329.100 210.150 330.900 211.950 ;
        RECT 323.700 206.700 327.300 207.600 ;
        RECT 323.700 204.600 324.900 206.700 ;
        RECT 302.100 198.600 303.900 201.600 ;
        RECT 305.100 198.000 306.900 201.600 ;
        RECT 314.100 198.000 315.900 201.600 ;
        RECT 317.100 198.600 318.900 201.600 ;
        RECT 323.100 198.600 324.900 204.600 ;
        RECT 326.100 203.700 333.900 205.050 ;
        RECT 326.100 198.600 327.900 203.700 ;
        RECT 329.100 198.000 330.900 202.800 ;
        RECT 332.100 198.600 333.900 203.700 ;
        RECT 341.700 201.600 342.900 211.950 ;
        RECT 351.000 208.200 351.900 211.950 ;
        RECT 353.100 210.150 354.900 211.950 ;
        RECT 359.100 210.150 360.900 211.950 ;
        RECT 351.000 207.000 354.300 208.200 ;
        RECT 341.100 198.600 342.900 201.600 ;
        RECT 344.100 198.000 345.900 201.600 ;
        RECT 352.500 198.600 354.300 207.000 ;
        RECT 359.100 198.000 360.900 207.600 ;
        RECT 2.700 188.400 4.500 194.400 ;
        RECT 8.100 188.400 9.900 195.000 ;
        RECT 13.500 188.400 15.300 194.400 ;
        RECT 17.700 191.400 19.500 194.400 ;
        RECT 20.700 191.400 22.500 194.400 ;
        RECT 23.700 191.400 25.500 194.400 ;
        RECT 26.700 191.400 28.500 195.000 ;
        RECT 17.700 189.300 19.800 191.400 ;
        RECT 20.700 189.300 22.800 191.400 ;
        RECT 23.700 189.300 25.800 191.400 ;
        RECT 31.200 190.500 33.000 194.400 ;
        RECT 34.200 191.400 36.000 195.000 ;
        RECT 37.200 191.400 39.000 194.400 ;
        RECT 40.200 191.400 42.000 194.400 ;
        RECT 43.200 191.400 45.000 194.400 ;
        RECT 46.200 191.400 48.000 194.400 ;
        RECT 27.600 189.600 29.400 190.500 ;
        RECT 26.700 188.400 29.400 189.600 ;
        RECT 31.200 188.400 33.900 190.500 ;
        RECT 37.200 189.300 39.300 191.400 ;
        RECT 40.200 189.300 42.300 191.400 ;
        RECT 43.200 189.300 45.300 191.400 ;
        RECT 46.200 189.300 48.300 191.400 ;
        RECT 50.400 189.600 52.200 194.400 ;
        RECT 50.400 188.400 54.600 189.600 ;
        RECT 55.500 188.400 57.300 195.000 ;
        RECT 60.900 188.400 62.700 194.400 ;
        RECT 2.700 184.800 3.900 188.400 ;
        RECT 13.800 187.500 15.300 188.400 ;
        RECT 22.800 187.800 24.600 188.400 ;
        RECT 26.700 187.800 27.600 188.400 ;
        RECT 6.900 186.300 15.300 187.500 ;
        RECT 20.400 186.600 27.600 187.800 ;
        RECT 42.300 186.600 48.900 188.400 ;
        RECT 6.900 185.700 8.700 186.300 ;
        RECT 17.400 184.800 19.500 185.700 ;
        RECT 2.700 183.600 19.500 184.800 ;
        RECT 20.400 183.600 21.300 186.600 ;
        RECT 25.800 183.900 27.600 184.800 ;
        RECT 35.100 184.500 36.900 186.300 ;
        RECT 53.100 185.100 54.600 188.400 ;
        RECT 28.800 183.900 30.900 184.050 ;
        RECT 2.700 167.400 3.900 183.600 ;
        RECT 20.400 181.800 22.200 183.600 ;
        RECT 25.800 183.000 30.900 183.900 ;
        RECT 28.800 181.950 30.900 183.000 ;
        RECT 35.100 183.900 37.200 184.500 ;
        RECT 35.100 182.400 52.200 183.900 ;
        RECT 53.100 183.300 60.900 185.100 ;
        RECT 50.700 180.900 57.300 182.400 ;
        RECT 5.100 179.700 49.500 180.900 ;
        RECT 5.100 178.050 6.900 179.700 ;
        RECT 4.800 175.950 6.900 178.050 ;
        RECT 10.800 177.750 12.900 178.050 ;
        RECT 23.400 177.900 25.200 178.500 ;
        RECT 32.400 177.900 45.900 178.800 ;
        RECT 10.800 175.950 14.700 177.750 ;
        RECT 23.400 176.700 34.500 177.900 ;
        RECT 12.900 175.200 14.700 175.950 ;
        RECT 32.400 175.800 34.500 176.700 ;
        RECT 36.000 175.200 39.900 177.000 ;
        RECT 45.000 176.700 45.900 177.900 ;
        RECT 12.900 174.300 26.400 175.200 ;
        RECT 37.800 174.900 39.900 175.200 ;
        RECT 44.100 174.900 45.900 176.700 ;
        RECT 48.600 178.200 49.500 179.700 ;
        RECT 48.600 176.400 53.700 178.200 ;
        RECT 55.800 178.050 57.300 180.900 ;
        RECT 55.800 175.950 57.900 178.050 ;
        RECT 25.200 173.700 26.400 174.300 ;
        RECT 59.100 173.700 60.900 174.300 ;
        RECT 20.400 172.500 22.500 172.800 ;
        RECT 25.200 172.500 60.900 173.700 ;
        RECT 10.500 171.300 22.500 172.500 ;
        RECT 61.800 171.600 62.700 188.400 ;
        RECT 10.500 170.700 12.300 171.300 ;
        RECT 20.400 170.700 22.500 171.300 ;
        RECT 25.200 170.400 42.900 171.600 ;
        RECT 7.200 169.800 9.000 170.100 ;
        RECT 25.200 169.800 26.400 170.400 ;
        RECT 7.200 168.600 26.400 169.800 ;
        RECT 40.800 169.500 42.900 170.400 ;
        RECT 46.200 170.700 62.700 171.600 ;
        RECT 46.200 169.500 48.300 170.700 ;
        RECT 7.200 168.300 9.000 168.600 ;
        RECT 2.700 166.500 6.300 167.400 ;
        RECT 5.400 165.600 6.300 166.500 ;
        RECT 2.700 159.000 4.500 165.600 ;
        RECT 5.400 164.700 7.500 165.600 ;
        RECT 5.700 159.600 7.500 164.700 ;
        RECT 8.700 159.000 10.500 165.600 ;
        RECT 11.700 159.600 13.500 168.600 ;
        RECT 23.700 165.600 25.800 167.700 ;
        RECT 31.200 167.100 34.500 169.200 ;
        RECT 14.700 159.000 16.500 165.600 ;
        RECT 18.300 162.600 20.400 164.700 ;
        RECT 21.300 162.600 23.400 164.700 ;
        RECT 18.300 159.600 20.100 162.600 ;
        RECT 21.300 159.600 23.100 162.600 ;
        RECT 24.300 159.600 26.100 165.600 ;
        RECT 27.300 159.000 29.100 165.600 ;
        RECT 31.200 159.600 33.000 167.100 ;
        RECT 37.200 165.600 39.900 169.500 ;
        RECT 52.200 168.600 57.900 169.800 ;
        RECT 49.500 167.700 51.300 168.300 ;
        RECT 43.200 166.500 51.300 167.700 ;
        RECT 43.200 165.600 45.300 166.500 ;
        RECT 52.200 165.600 53.400 168.600 ;
        RECT 56.100 168.000 57.900 168.600 ;
        RECT 61.800 167.400 62.700 170.700 ;
        RECT 58.800 166.500 62.700 167.400 ;
        RECT 64.500 191.400 66.300 194.400 ;
        RECT 67.500 191.400 69.300 195.000 ;
        RECT 64.500 178.050 66.000 191.400 ;
        RECT 77.100 185.400 78.900 195.000 ;
        RECT 83.700 186.000 85.500 194.400 ;
        RECT 97.500 186.000 99.300 194.400 ;
        RECT 83.700 184.800 87.000 186.000 ;
        RECT 77.100 181.050 78.900 182.850 ;
        RECT 83.100 181.050 84.900 182.850 ;
        RECT 86.100 181.050 87.000 184.800 ;
        RECT 96.000 184.800 99.300 186.000 ;
        RECT 104.100 185.400 105.900 195.000 ;
        RECT 113.400 188.400 115.200 195.000 ;
        RECT 118.500 187.200 120.300 194.400 ;
        RECT 116.100 186.300 120.300 187.200 ;
        RECT 125.700 187.200 127.500 194.400 ;
        RECT 130.800 188.400 132.600 195.000 ;
        RECT 137.100 191.400 138.900 194.400 ;
        RECT 140.100 191.400 141.900 195.000 ;
        RECT 149.700 191.400 151.500 195.000 ;
        RECT 125.700 186.300 129.900 187.200 ;
        RECT 96.000 181.050 96.900 184.800 ;
        RECT 98.100 181.050 99.900 182.850 ;
        RECT 104.100 181.050 105.900 182.850 ;
        RECT 113.250 181.050 115.050 182.850 ;
        RECT 116.100 181.050 117.300 186.300 ;
        RECT 119.100 181.050 120.900 182.850 ;
        RECT 125.100 181.050 126.900 182.850 ;
        RECT 128.700 181.050 129.900 186.300 ;
        RECT 130.950 181.050 132.750 182.850 ;
        RECT 137.700 181.050 138.900 191.400 ;
        RECT 152.700 189.600 154.500 194.400 ;
        RECT 149.400 188.400 154.500 189.600 ;
        RECT 157.200 188.400 159.000 195.000 ;
        RECT 149.400 181.050 150.300 188.400 ;
        RECT 169.500 186.000 171.300 194.400 ;
        RECT 168.000 184.800 171.300 186.000 ;
        RECT 176.100 185.400 177.900 195.000 ;
        RECT 185.400 188.400 187.200 195.000 ;
        RECT 190.500 187.200 192.300 194.400 ;
        RECT 188.100 186.300 192.300 187.200 ;
        RECT 194.700 188.400 196.500 194.400 ;
        RECT 200.100 188.400 201.900 195.000 ;
        RECT 205.500 188.400 207.300 194.400 ;
        RECT 209.700 191.400 211.500 194.400 ;
        RECT 212.700 191.400 214.500 194.400 ;
        RECT 215.700 191.400 217.500 194.400 ;
        RECT 218.700 191.400 220.500 195.000 ;
        RECT 209.700 189.300 211.800 191.400 ;
        RECT 212.700 189.300 214.800 191.400 ;
        RECT 215.700 189.300 217.800 191.400 ;
        RECT 223.200 190.500 225.000 194.400 ;
        RECT 226.200 191.400 228.000 195.000 ;
        RECT 229.200 191.400 231.000 194.400 ;
        RECT 232.200 191.400 234.000 194.400 ;
        RECT 235.200 191.400 237.000 194.400 ;
        RECT 238.200 191.400 240.000 194.400 ;
        RECT 219.600 189.600 221.400 190.500 ;
        RECT 218.700 188.400 221.400 189.600 ;
        RECT 223.200 188.400 225.900 190.500 ;
        RECT 229.200 189.300 231.300 191.400 ;
        RECT 232.200 189.300 234.300 191.400 ;
        RECT 235.200 189.300 237.300 191.400 ;
        RECT 238.200 189.300 240.300 191.400 ;
        RECT 242.400 189.600 244.200 194.400 ;
        RECT 242.400 188.400 246.600 189.600 ;
        RECT 247.500 188.400 249.300 195.000 ;
        RECT 252.900 188.400 254.700 194.400 ;
        RECT 151.950 181.050 153.750 182.850 ;
        RECT 158.100 181.050 159.900 182.850 ;
        RECT 168.000 181.050 168.900 184.800 ;
        RECT 170.100 181.050 171.900 182.850 ;
        RECT 176.100 181.050 177.900 182.850 ;
        RECT 185.250 181.050 187.050 182.850 ;
        RECT 188.100 181.050 189.300 186.300 ;
        RECT 194.700 184.800 195.900 188.400 ;
        RECT 205.800 187.500 207.300 188.400 ;
        RECT 214.800 187.800 216.600 188.400 ;
        RECT 218.700 187.800 219.600 188.400 ;
        RECT 198.900 186.300 207.300 187.500 ;
        RECT 212.400 186.600 219.600 187.800 ;
        RECT 234.300 186.600 240.900 188.400 ;
        RECT 198.900 185.700 200.700 186.300 ;
        RECT 209.400 184.800 211.500 185.700 ;
        RECT 194.700 183.600 211.500 184.800 ;
        RECT 212.400 183.600 213.300 186.600 ;
        RECT 217.800 183.900 219.600 184.800 ;
        RECT 227.100 184.500 228.900 186.300 ;
        RECT 245.100 185.100 246.600 188.400 ;
        RECT 220.800 183.900 222.900 184.050 ;
        RECT 191.100 181.050 192.900 182.850 ;
        RECT 76.950 178.950 79.050 181.050 ;
        RECT 79.950 178.950 82.050 181.050 ;
        RECT 82.950 178.950 85.050 181.050 ;
        RECT 85.950 178.950 88.050 181.050 ;
        RECT 94.950 178.950 97.050 181.050 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 100.950 178.950 103.050 181.050 ;
        RECT 103.950 178.950 106.050 181.050 ;
        RECT 112.950 178.950 115.050 181.050 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 118.950 178.950 121.050 181.050 ;
        RECT 124.950 178.950 127.050 181.050 ;
        RECT 127.950 178.950 130.050 181.050 ;
        RECT 130.950 178.950 133.050 181.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 148.950 178.950 151.050 181.050 ;
        RECT 151.950 178.950 154.050 181.050 ;
        RECT 154.950 178.950 157.050 181.050 ;
        RECT 157.950 178.950 160.050 181.050 ;
        RECT 166.950 178.950 169.050 181.050 ;
        RECT 169.950 178.950 172.050 181.050 ;
        RECT 172.950 178.950 175.050 181.050 ;
        RECT 175.950 178.950 178.050 181.050 ;
        RECT 184.950 178.950 187.050 181.050 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 190.950 178.950 193.050 181.050 ;
        RECT 64.500 175.950 66.900 178.050 ;
        RECT 67.950 177.450 70.050 178.050 ;
        RECT 73.950 177.450 76.050 178.050 ;
        RECT 67.950 176.550 76.050 177.450 ;
        RECT 80.100 177.150 81.900 178.950 ;
        RECT 67.950 175.950 70.050 176.550 ;
        RECT 73.950 175.950 76.050 176.550 ;
        RECT 58.800 165.600 60.000 166.500 ;
        RECT 64.500 165.600 66.000 175.950 ;
        RECT 67.950 174.450 70.050 174.900 ;
        RECT 82.950 174.450 85.050 175.050 ;
        RECT 67.950 173.550 85.050 174.450 ;
        RECT 67.950 172.800 70.050 173.550 ;
        RECT 82.950 172.950 85.050 173.550 ;
        RECT 86.100 166.800 87.000 178.950 ;
        RECT 80.400 165.900 87.000 166.800 ;
        RECT 80.400 165.600 81.900 165.900 ;
        RECT 34.200 159.000 36.000 165.600 ;
        RECT 37.200 159.600 39.000 165.600 ;
        RECT 40.200 162.600 42.300 164.700 ;
        RECT 43.200 162.600 45.300 164.700 ;
        RECT 46.200 162.600 48.300 164.700 ;
        RECT 40.200 159.600 42.000 162.600 ;
        RECT 43.200 159.600 45.000 162.600 ;
        RECT 46.200 159.600 48.000 162.600 ;
        RECT 49.200 159.000 51.000 165.600 ;
        RECT 52.200 159.600 54.000 165.600 ;
        RECT 55.200 159.000 57.000 165.600 ;
        RECT 58.200 159.600 60.000 165.600 ;
        RECT 61.200 159.000 63.000 165.600 ;
        RECT 64.500 159.600 66.300 165.600 ;
        RECT 67.500 159.000 69.300 165.600 ;
        RECT 77.100 159.000 78.900 165.600 ;
        RECT 80.100 159.600 81.900 165.600 ;
        RECT 86.100 165.600 87.000 165.900 ;
        RECT 96.000 166.800 96.900 178.950 ;
        RECT 101.100 177.150 102.900 178.950 ;
        RECT 96.000 165.900 102.600 166.800 ;
        RECT 96.000 165.600 96.900 165.900 ;
        RECT 83.100 159.000 84.900 165.000 ;
        RECT 86.100 159.600 87.900 165.600 ;
        RECT 95.100 159.600 96.900 165.600 ;
        RECT 101.100 165.600 102.600 165.900 ;
        RECT 116.100 165.600 117.300 178.950 ;
        RECT 128.700 165.600 129.900 178.950 ;
        RECT 133.950 174.450 136.050 178.050 ;
        RECT 131.550 174.000 136.050 174.450 ;
        RECT 130.950 173.550 135.450 174.000 ;
        RECT 130.950 169.950 133.050 173.550 ;
        RECT 137.700 165.600 138.900 178.950 ;
        RECT 140.100 177.150 141.900 178.950 ;
        RECT 149.400 171.600 150.300 178.950 ;
        RECT 154.950 177.150 156.750 178.950 ;
        RECT 98.100 159.000 99.900 165.000 ;
        RECT 101.100 159.600 102.900 165.600 ;
        RECT 104.100 159.000 105.900 165.600 ;
        RECT 113.100 159.000 114.900 165.600 ;
        RECT 116.100 159.600 117.900 165.600 ;
        RECT 119.100 159.000 120.900 165.600 ;
        RECT 125.100 159.000 126.900 165.600 ;
        RECT 128.100 159.600 129.900 165.600 ;
        RECT 131.100 159.000 132.900 165.600 ;
        RECT 137.100 159.600 138.900 165.600 ;
        RECT 140.100 159.000 141.900 165.600 ;
        RECT 149.100 159.600 150.900 171.600 ;
        RECT 152.100 170.700 159.900 171.600 ;
        RECT 152.100 159.600 153.900 170.700 ;
        RECT 155.100 159.000 156.900 169.800 ;
        RECT 158.100 159.600 159.900 170.700 ;
        RECT 168.000 166.800 168.900 178.950 ;
        RECT 173.100 177.150 174.900 178.950 ;
        RECT 168.000 165.900 174.600 166.800 ;
        RECT 168.000 165.600 168.900 165.900 ;
        RECT 167.100 159.600 168.900 165.600 ;
        RECT 173.100 165.600 174.600 165.900 ;
        RECT 188.100 165.600 189.300 178.950 ;
        RECT 194.700 167.400 195.900 183.600 ;
        RECT 212.400 181.800 214.200 183.600 ;
        RECT 217.800 183.000 222.900 183.900 ;
        RECT 220.800 181.950 222.900 183.000 ;
        RECT 227.100 183.900 229.200 184.500 ;
        RECT 227.100 182.400 244.200 183.900 ;
        RECT 245.100 183.300 252.900 185.100 ;
        RECT 242.700 180.900 249.300 182.400 ;
        RECT 197.100 179.700 241.500 180.900 ;
        RECT 197.100 178.050 198.900 179.700 ;
        RECT 196.800 175.950 198.900 178.050 ;
        RECT 202.800 177.750 204.900 178.050 ;
        RECT 215.400 177.900 217.200 178.500 ;
        RECT 224.400 177.900 237.900 178.800 ;
        RECT 202.800 175.950 206.700 177.750 ;
        RECT 215.400 176.700 226.500 177.900 ;
        RECT 204.900 175.200 206.700 175.950 ;
        RECT 224.400 175.800 226.500 176.700 ;
        RECT 228.000 175.200 231.900 177.000 ;
        RECT 237.000 176.700 237.900 177.900 ;
        RECT 204.900 174.300 218.400 175.200 ;
        RECT 229.800 174.900 231.900 175.200 ;
        RECT 236.100 174.900 237.900 176.700 ;
        RECT 240.600 178.200 241.500 179.700 ;
        RECT 240.600 176.400 245.700 178.200 ;
        RECT 247.800 178.050 249.300 180.900 ;
        RECT 247.800 175.950 249.900 178.050 ;
        RECT 217.200 173.700 218.400 174.300 ;
        RECT 251.100 173.700 252.900 174.300 ;
        RECT 212.400 172.500 214.500 172.800 ;
        RECT 217.200 172.500 252.900 173.700 ;
        RECT 202.500 171.300 214.500 172.500 ;
        RECT 253.800 171.600 254.700 188.400 ;
        RECT 202.500 170.700 204.300 171.300 ;
        RECT 212.400 170.700 214.500 171.300 ;
        RECT 217.200 170.400 234.900 171.600 ;
        RECT 199.200 169.800 201.000 170.100 ;
        RECT 217.200 169.800 218.400 170.400 ;
        RECT 199.200 168.600 218.400 169.800 ;
        RECT 232.800 169.500 234.900 170.400 ;
        RECT 238.200 170.700 254.700 171.600 ;
        RECT 238.200 169.500 240.300 170.700 ;
        RECT 199.200 168.300 201.000 168.600 ;
        RECT 194.700 166.500 198.300 167.400 ;
        RECT 197.400 165.600 198.300 166.500 ;
        RECT 170.100 159.000 171.900 165.000 ;
        RECT 173.100 159.600 174.900 165.600 ;
        RECT 176.100 159.000 177.900 165.600 ;
        RECT 185.100 159.000 186.900 165.600 ;
        RECT 188.100 159.600 189.900 165.600 ;
        RECT 191.100 159.000 192.900 165.600 ;
        RECT 194.700 159.000 196.500 165.600 ;
        RECT 197.400 164.700 199.500 165.600 ;
        RECT 197.700 159.600 199.500 164.700 ;
        RECT 200.700 159.000 202.500 165.600 ;
        RECT 203.700 159.600 205.500 168.600 ;
        RECT 215.700 165.600 217.800 167.700 ;
        RECT 223.200 167.100 226.500 169.200 ;
        RECT 206.700 159.000 208.500 165.600 ;
        RECT 210.300 162.600 212.400 164.700 ;
        RECT 213.300 162.600 215.400 164.700 ;
        RECT 210.300 159.600 212.100 162.600 ;
        RECT 213.300 159.600 215.100 162.600 ;
        RECT 216.300 159.600 218.100 165.600 ;
        RECT 219.300 159.000 221.100 165.600 ;
        RECT 223.200 159.600 225.000 167.100 ;
        RECT 229.200 165.600 231.900 169.500 ;
        RECT 244.200 168.600 249.900 169.800 ;
        RECT 241.500 167.700 243.300 168.300 ;
        RECT 235.200 166.500 243.300 167.700 ;
        RECT 235.200 165.600 237.300 166.500 ;
        RECT 244.200 165.600 245.400 168.600 ;
        RECT 248.100 168.000 249.900 168.600 ;
        RECT 253.800 167.400 254.700 170.700 ;
        RECT 250.800 166.500 254.700 167.400 ;
        RECT 256.500 191.400 258.300 194.400 ;
        RECT 259.500 191.400 261.300 195.000 ;
        RECT 256.500 178.050 258.000 191.400 ;
        RECT 266.400 188.400 268.200 195.000 ;
        RECT 271.500 187.200 273.300 194.400 ;
        RECT 269.100 186.300 273.300 187.200 ;
        RECT 281.100 190.200 282.900 193.200 ;
        RECT 284.100 192.600 285.300 195.000 ;
        RECT 293.100 193.200 294.300 195.000 ;
        RECT 281.100 186.900 282.000 190.200 ;
        RECT 284.100 187.800 285.900 192.600 ;
        RECT 288.600 188.700 290.400 193.200 ;
        RECT 288.600 187.800 290.700 188.700 ;
        RECT 266.250 181.050 268.050 182.850 ;
        RECT 269.100 181.050 270.300 186.300 ;
        RECT 281.100 186.000 288.300 186.900 ;
        RECT 272.100 181.050 273.900 182.850 ;
        RECT 281.100 181.050 282.900 182.850 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 268.950 178.950 271.050 181.050 ;
        RECT 271.950 178.950 274.050 181.050 ;
        RECT 281.100 178.950 283.200 181.050 ;
        RECT 284.100 178.950 286.200 181.050 ;
        RECT 287.100 178.950 288.300 186.000 ;
        RECT 289.800 181.050 290.700 187.800 ;
        RECT 293.100 187.200 294.900 193.200 ;
        RECT 299.100 189.300 300.900 194.400 ;
        RECT 302.100 190.200 303.900 195.000 ;
        RECT 305.100 189.300 306.900 194.400 ;
        RECT 299.100 187.950 306.900 189.300 ;
        RECT 308.100 188.400 309.900 194.400 ;
        RECT 308.100 186.300 309.300 188.400 ;
        RECT 317.700 187.200 319.500 194.400 ;
        RECT 322.800 188.400 324.600 195.000 ;
        RECT 329.100 191.400 330.900 195.000 ;
        RECT 332.100 191.400 333.900 194.400 ;
        RECT 341.100 191.400 342.900 194.400 ;
        RECT 317.700 186.300 321.900 187.200 ;
        RECT 305.700 185.400 309.300 186.300 ;
        RECT 302.100 181.050 303.900 182.850 ;
        RECT 305.700 181.050 306.900 185.400 ;
        RECT 308.100 181.050 309.900 182.850 ;
        RECT 317.100 181.050 318.900 182.850 ;
        RECT 320.700 181.050 321.900 186.300 ;
        RECT 322.950 181.050 324.750 182.850 ;
        RECT 332.100 181.050 333.300 191.400 ;
        RECT 341.100 187.500 342.300 191.400 ;
        RECT 344.100 188.400 345.900 195.000 ;
        RECT 347.100 188.400 348.900 194.400 ;
        RECT 341.100 186.600 346.800 187.500 ;
        RECT 345.000 185.700 346.800 186.600 ;
        RECT 289.800 178.950 291.900 181.050 ;
        RECT 292.800 178.950 294.900 181.050 ;
        RECT 298.950 178.950 301.050 181.050 ;
        RECT 301.950 178.950 304.050 181.050 ;
        RECT 304.950 178.950 307.050 181.050 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 316.950 178.950 319.050 181.050 ;
        RECT 319.950 178.950 322.050 181.050 ;
        RECT 322.950 178.950 325.050 181.050 ;
        RECT 328.950 178.950 331.050 181.050 ;
        RECT 331.950 178.950 334.050 181.050 ;
        RECT 341.400 178.950 343.500 181.050 ;
        RECT 256.500 175.950 258.900 178.050 ;
        RECT 250.800 165.600 252.000 166.500 ;
        RECT 256.500 165.600 258.000 175.950 ;
        RECT 269.100 165.600 270.300 178.950 ;
        RECT 284.100 177.150 285.900 178.950 ;
        RECT 287.100 177.150 288.900 178.950 ;
        RECT 287.700 172.800 288.900 177.150 ;
        RECT 281.100 171.900 288.900 172.800 ;
        RECT 281.100 166.800 282.000 171.900 ;
        RECT 289.800 171.000 290.700 178.950 ;
        RECT 292.800 177.150 294.600 178.950 ;
        RECT 299.100 177.150 300.900 178.950 ;
        RECT 292.950 174.450 295.050 175.050 ;
        RECT 301.950 174.450 304.050 175.050 ;
        RECT 292.950 173.550 304.050 174.450 ;
        RECT 292.950 172.950 295.050 173.550 ;
        RECT 301.950 172.950 304.050 173.550 ;
        RECT 305.700 171.600 306.900 178.950 ;
        RECT 226.200 159.000 228.000 165.600 ;
        RECT 229.200 159.600 231.000 165.600 ;
        RECT 232.200 162.600 234.300 164.700 ;
        RECT 235.200 162.600 237.300 164.700 ;
        RECT 238.200 162.600 240.300 164.700 ;
        RECT 232.200 159.600 234.000 162.600 ;
        RECT 235.200 159.600 237.000 162.600 ;
        RECT 238.200 159.600 240.000 162.600 ;
        RECT 241.200 159.000 243.000 165.600 ;
        RECT 244.200 159.600 246.000 165.600 ;
        RECT 247.200 159.000 249.000 165.600 ;
        RECT 250.200 159.600 252.000 165.600 ;
        RECT 253.200 159.000 255.000 165.600 ;
        RECT 256.500 159.600 258.300 165.600 ;
        RECT 259.500 159.000 261.300 165.600 ;
        RECT 266.100 159.000 267.900 165.600 ;
        RECT 269.100 159.600 270.900 165.600 ;
        RECT 272.100 159.000 273.900 165.600 ;
        RECT 281.100 160.800 282.900 166.800 ;
        RECT 284.100 159.000 285.900 171.000 ;
        RECT 288.600 170.100 290.700 171.000 ;
        RECT 288.600 159.600 290.400 170.100 ;
        RECT 293.100 159.000 294.900 171.600 ;
        RECT 299.400 159.000 301.200 171.600 ;
        RECT 304.500 170.100 306.900 171.600 ;
        RECT 304.500 159.600 306.300 170.100 ;
        RECT 307.200 167.100 309.000 168.900 ;
        RECT 320.700 165.600 321.900 178.950 ;
        RECT 329.100 177.150 330.900 178.950 ;
        RECT 332.100 165.600 333.300 178.950 ;
        RECT 341.400 177.150 343.200 178.950 ;
        RECT 345.000 174.300 345.900 185.700 ;
        RECT 347.700 181.050 348.900 188.400 ;
        RECT 353.100 191.400 354.900 194.400 ;
        RECT 353.100 187.500 354.300 191.400 ;
        RECT 356.100 188.400 357.900 195.000 ;
        RECT 359.100 188.400 360.900 194.400 ;
        RECT 353.100 186.600 358.800 187.500 ;
        RECT 357.000 185.700 358.800 186.600 ;
        RECT 346.800 178.950 348.900 181.050 ;
        RECT 345.000 173.400 346.800 174.300 ;
        RECT 341.100 172.500 346.800 173.400 ;
        RECT 341.100 165.600 342.300 172.500 ;
        RECT 347.700 171.600 348.900 178.950 ;
        RECT 353.400 178.950 355.500 181.050 ;
        RECT 353.400 177.150 355.200 178.950 ;
        RECT 357.000 174.300 357.900 185.700 ;
        RECT 359.700 181.050 360.900 188.400 ;
        RECT 358.800 178.950 360.900 181.050 ;
        RECT 357.000 173.400 358.800 174.300 ;
        RECT 307.500 159.000 309.300 165.600 ;
        RECT 317.100 159.000 318.900 165.600 ;
        RECT 320.100 159.600 321.900 165.600 ;
        RECT 323.100 159.000 324.900 165.600 ;
        RECT 329.100 159.000 330.900 165.600 ;
        RECT 332.100 159.600 333.900 165.600 ;
        RECT 341.100 159.600 342.900 165.600 ;
        RECT 344.100 159.000 345.900 169.800 ;
        RECT 347.100 159.600 348.900 171.600 ;
        RECT 353.100 172.500 358.800 173.400 ;
        RECT 353.100 165.600 354.300 172.500 ;
        RECT 359.700 171.600 360.900 178.950 ;
        RECT 353.100 159.600 354.900 165.600 ;
        RECT 356.100 159.000 357.900 169.800 ;
        RECT 359.100 159.600 360.900 171.600 ;
        RECT 2.700 149.400 4.500 156.000 ;
        RECT 5.700 150.300 7.500 155.400 ;
        RECT 5.400 149.400 7.500 150.300 ;
        RECT 8.700 149.400 10.500 156.000 ;
        RECT 5.400 148.500 6.300 149.400 ;
        RECT 2.700 147.600 6.300 148.500 ;
        RECT 2.700 131.400 3.900 147.600 ;
        RECT 7.200 146.400 9.000 146.700 ;
        RECT 11.700 146.400 13.500 155.400 ;
        RECT 14.700 149.400 16.500 156.000 ;
        RECT 18.300 152.400 20.100 155.400 ;
        RECT 21.300 152.400 23.100 155.400 ;
        RECT 18.300 150.300 20.400 152.400 ;
        RECT 21.300 150.300 23.400 152.400 ;
        RECT 24.300 149.400 26.100 155.400 ;
        RECT 27.300 149.400 29.100 156.000 ;
        RECT 23.700 147.300 25.800 149.400 ;
        RECT 31.200 147.900 33.000 155.400 ;
        RECT 34.200 149.400 36.000 156.000 ;
        RECT 37.200 149.400 39.000 155.400 ;
        RECT 40.200 152.400 42.000 155.400 ;
        RECT 43.200 152.400 45.000 155.400 ;
        RECT 46.200 152.400 48.000 155.400 ;
        RECT 40.200 150.300 42.300 152.400 ;
        RECT 43.200 150.300 45.300 152.400 ;
        RECT 46.200 150.300 48.300 152.400 ;
        RECT 49.200 149.400 51.000 156.000 ;
        RECT 52.200 149.400 54.000 155.400 ;
        RECT 55.200 149.400 57.000 156.000 ;
        RECT 58.200 149.400 60.000 155.400 ;
        RECT 61.200 149.400 63.000 156.000 ;
        RECT 64.500 149.400 66.300 155.400 ;
        RECT 67.500 149.400 69.300 156.000 ;
        RECT 74.100 149.400 75.900 156.000 ;
        RECT 77.100 149.400 78.900 155.400 ;
        RECT 80.100 149.400 81.900 156.000 ;
        RECT 7.200 145.200 26.400 146.400 ;
        RECT 31.200 145.800 34.500 147.900 ;
        RECT 37.200 145.500 39.900 149.400 ;
        RECT 43.200 148.500 45.300 149.400 ;
        RECT 43.200 147.300 51.300 148.500 ;
        RECT 49.500 146.700 51.300 147.300 ;
        RECT 52.200 146.400 53.400 149.400 ;
        RECT 58.800 148.500 60.000 149.400 ;
        RECT 58.800 147.600 62.700 148.500 ;
        RECT 56.100 146.400 57.900 147.000 ;
        RECT 7.200 144.900 9.000 145.200 ;
        RECT 25.200 144.600 26.400 145.200 ;
        RECT 40.800 144.600 42.900 145.500 ;
        RECT 10.500 143.700 12.300 144.300 ;
        RECT 20.400 143.700 22.500 144.300 ;
        RECT 10.500 142.500 22.500 143.700 ;
        RECT 25.200 143.400 42.900 144.600 ;
        RECT 46.200 144.300 48.300 145.500 ;
        RECT 52.200 145.200 57.900 146.400 ;
        RECT 61.800 144.300 62.700 147.600 ;
        RECT 46.200 143.400 62.700 144.300 ;
        RECT 20.400 142.200 22.500 142.500 ;
        RECT 25.200 141.300 60.900 142.500 ;
        RECT 25.200 140.700 26.400 141.300 ;
        RECT 59.100 140.700 60.900 141.300 ;
        RECT 12.900 139.800 26.400 140.700 ;
        RECT 37.800 139.800 39.900 140.100 ;
        RECT 12.900 139.050 14.700 139.800 ;
        RECT 4.800 136.950 6.900 139.050 ;
        RECT 10.800 137.250 14.700 139.050 ;
        RECT 32.400 138.300 34.500 139.200 ;
        RECT 10.800 136.950 12.900 137.250 ;
        RECT 23.400 137.100 34.500 138.300 ;
        RECT 36.000 138.000 39.900 139.800 ;
        RECT 44.100 138.300 45.900 140.100 ;
        RECT 45.000 137.100 45.900 138.300 ;
        RECT 5.100 135.300 6.900 136.950 ;
        RECT 23.400 136.500 25.200 137.100 ;
        RECT 32.400 136.200 45.900 137.100 ;
        RECT 48.600 136.800 53.700 138.600 ;
        RECT 55.800 136.950 57.900 139.050 ;
        RECT 48.600 135.300 49.500 136.800 ;
        RECT 5.100 134.100 49.500 135.300 ;
        RECT 55.800 134.100 57.300 136.950 ;
        RECT 20.400 131.400 22.200 133.200 ;
        RECT 28.800 132.000 30.900 133.050 ;
        RECT 50.700 132.600 57.300 134.100 ;
        RECT 2.700 130.200 19.500 131.400 ;
        RECT 2.700 126.600 3.900 130.200 ;
        RECT 17.400 129.300 19.500 130.200 ;
        RECT 6.900 128.700 8.700 129.300 ;
        RECT 6.900 127.500 15.300 128.700 ;
        RECT 13.800 126.600 15.300 127.500 ;
        RECT 20.400 128.400 21.300 131.400 ;
        RECT 25.800 131.100 30.900 132.000 ;
        RECT 25.800 130.200 27.600 131.100 ;
        RECT 28.800 130.950 30.900 131.100 ;
        RECT 35.100 131.100 52.200 132.600 ;
        RECT 35.100 130.500 37.200 131.100 ;
        RECT 35.100 128.700 36.900 130.500 ;
        RECT 53.100 129.900 60.900 131.700 ;
        RECT 20.400 127.200 27.600 128.400 ;
        RECT 22.800 126.600 24.600 127.200 ;
        RECT 26.700 126.600 27.600 127.200 ;
        RECT 42.300 126.600 48.900 128.400 ;
        RECT 53.100 126.600 54.600 129.900 ;
        RECT 61.800 126.600 62.700 143.400 ;
        RECT 2.700 120.600 4.500 126.600 ;
        RECT 8.100 120.000 9.900 126.600 ;
        RECT 13.500 120.600 15.300 126.600 ;
        RECT 17.700 123.600 19.800 125.700 ;
        RECT 20.700 123.600 22.800 125.700 ;
        RECT 23.700 123.600 25.800 125.700 ;
        RECT 26.700 125.400 29.400 126.600 ;
        RECT 27.600 124.500 29.400 125.400 ;
        RECT 31.200 124.500 33.900 126.600 ;
        RECT 17.700 120.600 19.500 123.600 ;
        RECT 20.700 120.600 22.500 123.600 ;
        RECT 23.700 120.600 25.500 123.600 ;
        RECT 26.700 120.000 28.500 123.600 ;
        RECT 31.200 120.600 33.000 124.500 ;
        RECT 37.200 123.600 39.300 125.700 ;
        RECT 40.200 123.600 42.300 125.700 ;
        RECT 43.200 123.600 45.300 125.700 ;
        RECT 46.200 123.600 48.300 125.700 ;
        RECT 50.400 125.400 54.600 126.600 ;
        RECT 34.200 120.000 36.000 123.600 ;
        RECT 37.200 120.600 39.000 123.600 ;
        RECT 40.200 120.600 42.000 123.600 ;
        RECT 43.200 120.600 45.000 123.600 ;
        RECT 46.200 120.600 48.000 123.600 ;
        RECT 50.400 120.600 52.200 125.400 ;
        RECT 55.500 120.000 57.300 126.600 ;
        RECT 60.900 120.600 62.700 126.600 ;
        RECT 64.500 139.050 66.000 149.400 ;
        RECT 64.500 136.950 66.900 139.050 ;
        RECT 64.500 123.600 66.000 136.950 ;
        RECT 77.700 136.050 78.900 149.400 ;
        RECT 89.100 143.400 90.900 155.400 ;
        RECT 92.100 144.300 93.900 155.400 ;
        RECT 95.100 145.200 96.900 156.000 ;
        RECT 98.100 144.300 99.900 155.400 ;
        RECT 107.700 149.400 109.500 156.000 ;
        RECT 108.000 146.100 109.800 147.900 ;
        RECT 110.700 144.900 112.500 155.400 ;
        RECT 92.100 143.400 99.900 144.300 ;
        RECT 110.100 143.400 112.500 144.900 ;
        RECT 115.800 143.400 117.600 156.000 ;
        RECT 122.100 149.400 123.900 156.000 ;
        RECT 125.100 149.400 126.900 155.400 ;
        RECT 128.100 149.400 129.900 156.000 ;
        RECT 89.400 136.050 90.300 143.400 ;
        RECT 94.950 136.050 96.750 137.850 ;
        RECT 110.100 136.050 111.300 143.400 ;
        RECT 116.100 136.050 117.900 137.850 ;
        RECT 125.700 136.050 126.900 149.400 ;
        RECT 135.600 143.400 137.400 156.000 ;
        RECT 140.100 143.400 143.400 155.400 ;
        RECT 146.100 143.400 147.900 156.000 ;
        RECT 155.100 149.400 156.900 155.400 ;
        RECT 158.100 149.400 159.900 156.000 ;
        RECT 167.100 149.400 168.900 156.000 ;
        RECT 170.100 149.400 171.900 155.400 ;
        RECT 176.100 149.400 177.900 156.000 ;
        RECT 179.100 149.400 180.900 155.400 ;
        RECT 182.100 149.400 183.900 156.000 ;
        RECT 134.250 136.050 136.050 137.850 ;
        RECT 141.000 136.050 142.050 143.400 ;
        RECT 146.100 136.050 147.900 137.850 ;
        RECT 155.700 136.050 156.900 149.400 ;
        RECT 158.100 136.050 159.900 137.850 ;
        RECT 167.100 136.050 168.900 137.850 ;
        RECT 170.100 136.050 171.300 149.400 ;
        RECT 179.700 136.050 180.900 149.400 ;
        RECT 191.100 143.400 192.900 155.400 ;
        RECT 194.100 144.000 195.900 156.000 ;
        RECT 197.100 149.400 198.900 155.400 ;
        RECT 200.100 149.400 201.900 156.000 ;
        RECT 209.100 149.400 210.900 156.000 ;
        RECT 212.100 149.400 213.900 155.400 ;
        RECT 215.100 149.400 216.900 156.000 ;
        RECT 191.700 136.050 192.600 143.400 ;
        RECT 195.000 136.050 196.800 137.850 ;
        RECT 73.950 133.950 76.050 136.050 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 88.950 133.950 91.050 136.050 ;
        RECT 91.950 133.950 94.050 136.050 ;
        RECT 94.950 133.950 97.050 136.050 ;
        RECT 97.950 133.950 100.050 136.050 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 109.950 133.950 112.050 136.050 ;
        RECT 112.950 133.950 115.050 136.050 ;
        RECT 115.950 133.950 118.050 136.050 ;
        RECT 121.950 133.950 124.050 136.050 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 133.950 133.950 136.050 136.050 ;
        RECT 136.950 133.950 139.050 136.050 ;
        RECT 139.950 133.950 142.050 136.050 ;
        RECT 74.100 132.150 75.900 133.950 ;
        RECT 77.700 128.700 78.900 133.950 ;
        RECT 79.950 132.150 81.750 133.950 ;
        RECT 74.700 127.800 78.900 128.700 ;
        RECT 64.500 120.600 66.300 123.600 ;
        RECT 67.500 120.000 69.300 123.600 ;
        RECT 74.700 120.600 76.500 127.800 ;
        RECT 89.400 126.600 90.300 133.950 ;
        RECT 91.950 132.150 93.750 133.950 ;
        RECT 98.100 132.150 99.900 133.950 ;
        RECT 107.100 132.150 108.900 133.950 ;
        RECT 110.100 129.600 111.300 133.950 ;
        RECT 113.100 132.150 114.900 133.950 ;
        RECT 122.100 132.150 123.900 133.950 ;
        RECT 107.700 128.700 111.300 129.600 ;
        RECT 125.700 128.700 126.900 133.950 ;
        RECT 127.950 132.150 129.750 133.950 ;
        RECT 137.250 132.150 139.050 133.950 ;
        RECT 141.000 129.300 142.050 133.950 ;
        RECT 142.950 133.950 145.050 136.050 ;
        RECT 145.950 133.950 148.050 136.050 ;
        RECT 154.950 133.950 157.050 136.050 ;
        RECT 157.950 133.950 160.050 136.050 ;
        RECT 166.950 133.950 169.050 136.050 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 175.950 133.950 178.050 136.050 ;
        RECT 178.950 133.950 181.050 136.050 ;
        RECT 181.950 133.950 184.050 136.050 ;
        RECT 191.100 133.950 193.200 136.050 ;
        RECT 194.400 133.950 196.500 136.050 ;
        RECT 142.950 132.150 144.750 133.950 ;
        RECT 107.700 126.600 108.900 128.700 ;
        RECT 122.700 127.800 126.900 128.700 ;
        RECT 137.700 128.100 142.050 129.300 ;
        RECT 79.800 120.000 81.600 126.600 ;
        RECT 89.400 125.400 94.500 126.600 ;
        RECT 89.700 120.000 91.500 123.600 ;
        RECT 92.700 120.600 94.500 125.400 ;
        RECT 97.200 120.000 99.000 126.600 ;
        RECT 107.100 120.600 108.900 126.600 ;
        RECT 110.100 125.700 117.900 127.050 ;
        RECT 110.100 120.600 111.900 125.700 ;
        RECT 113.100 120.000 114.900 124.800 ;
        RECT 116.100 120.600 117.900 125.700 ;
        RECT 122.700 120.600 124.500 127.800 ;
        RECT 137.700 126.600 138.600 128.100 ;
        RECT 127.800 120.000 129.600 126.600 ;
        RECT 134.100 121.500 135.900 126.600 ;
        RECT 137.100 122.400 138.900 126.600 ;
        RECT 140.100 126.000 147.900 126.900 ;
        RECT 140.100 121.500 141.900 126.000 ;
        RECT 134.100 120.600 141.900 121.500 ;
        RECT 143.100 120.000 144.900 125.100 ;
        RECT 146.100 120.600 147.900 126.000 ;
        RECT 155.700 123.600 156.900 133.950 ;
        RECT 170.100 123.600 171.300 133.950 ;
        RECT 176.100 132.150 177.900 133.950 ;
        RECT 179.700 128.700 180.900 133.950 ;
        RECT 181.950 132.150 183.750 133.950 ;
        RECT 176.700 127.800 180.900 128.700 ;
        RECT 155.100 120.600 156.900 123.600 ;
        RECT 158.100 120.000 159.900 123.600 ;
        RECT 167.100 120.000 168.900 123.600 ;
        RECT 170.100 120.600 171.900 123.600 ;
        RECT 176.700 120.600 178.500 127.800 ;
        RECT 191.700 126.600 192.600 133.950 ;
        RECT 198.000 129.300 198.900 149.400 ;
        RECT 212.700 136.050 213.900 149.400 ;
        RECT 224.100 143.400 225.900 155.400 ;
        RECT 227.100 145.200 228.900 156.000 ;
        RECT 230.100 149.400 231.900 155.400 ;
        RECT 236.100 149.400 237.900 156.000 ;
        RECT 239.100 149.400 240.900 155.400 ;
        RECT 242.100 149.400 243.900 156.000 ;
        RECT 224.100 136.050 225.300 143.400 ;
        RECT 230.700 142.500 231.900 149.400 ;
        RECT 226.200 141.600 231.900 142.500 ;
        RECT 226.200 140.700 228.000 141.600 ;
        RECT 199.800 133.950 201.900 136.050 ;
        RECT 208.950 133.950 211.050 136.050 ;
        RECT 211.950 133.950 214.050 136.050 ;
        RECT 214.950 133.950 217.050 136.050 ;
        RECT 224.100 133.950 226.200 136.050 ;
        RECT 199.950 132.150 201.750 133.950 ;
        RECT 209.100 132.150 210.900 133.950 ;
        RECT 193.500 128.400 201.900 129.300 ;
        RECT 212.700 128.700 213.900 133.950 ;
        RECT 214.950 132.150 216.750 133.950 ;
        RECT 193.500 127.500 195.300 128.400 ;
        RECT 181.800 120.000 183.600 126.600 ;
        RECT 191.700 124.800 194.400 126.600 ;
        RECT 192.600 120.600 194.400 124.800 ;
        RECT 195.600 120.000 197.400 126.600 ;
        RECT 200.100 120.600 201.900 128.400 ;
        RECT 209.700 127.800 213.900 128.700 ;
        RECT 209.700 120.600 211.500 127.800 ;
        RECT 224.100 126.600 225.300 133.950 ;
        RECT 227.100 129.300 228.000 140.700 ;
        RECT 229.800 136.050 231.600 137.850 ;
        RECT 239.100 136.050 240.300 149.400 ;
        RECT 248.100 144.300 249.900 155.400 ;
        RECT 251.100 145.200 252.900 156.000 ;
        RECT 254.100 144.300 255.900 155.400 ;
        RECT 248.100 143.400 255.900 144.300 ;
        RECT 257.100 143.400 258.900 155.400 ;
        RECT 266.100 149.400 267.900 156.000 ;
        RECT 269.100 149.400 270.900 155.400 ;
        RECT 272.100 149.400 273.900 156.000 ;
        RECT 278.100 149.400 279.900 156.000 ;
        RECT 281.100 149.400 282.900 155.400 ;
        RECT 284.100 150.000 285.900 156.000 ;
        RECT 251.250 136.050 253.050 137.850 ;
        RECT 257.700 136.050 258.600 143.400 ;
        RECT 269.700 136.050 270.900 149.400 ;
        RECT 281.400 149.100 282.900 149.400 ;
        RECT 287.100 149.400 288.900 155.400 ;
        RECT 290.700 149.400 292.500 156.000 ;
        RECT 293.700 150.300 295.500 155.400 ;
        RECT 293.400 149.400 295.500 150.300 ;
        RECT 296.700 149.400 298.500 156.000 ;
        RECT 287.100 149.100 288.000 149.400 ;
        RECT 281.400 148.200 288.000 149.100 ;
        RECT 293.400 148.500 294.300 149.400 ;
        RECT 281.100 136.050 282.900 137.850 ;
        RECT 287.100 136.050 288.000 148.200 ;
        RECT 290.700 147.600 294.300 148.500 ;
        RECT 229.500 133.950 231.600 136.050 ;
        RECT 235.950 133.950 238.050 136.050 ;
        RECT 238.950 133.950 241.050 136.050 ;
        RECT 241.950 133.950 244.050 136.050 ;
        RECT 247.950 133.950 250.050 136.050 ;
        RECT 250.950 133.950 253.050 136.050 ;
        RECT 253.950 133.950 256.050 136.050 ;
        RECT 256.950 133.950 259.050 136.050 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 268.950 133.950 271.050 136.050 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 277.950 133.950 280.050 136.050 ;
        RECT 280.950 133.950 283.050 136.050 ;
        RECT 283.950 133.950 286.050 136.050 ;
        RECT 286.950 133.950 289.050 136.050 ;
        RECT 236.250 132.150 238.050 133.950 ;
        RECT 226.200 128.400 228.000 129.300 ;
        RECT 239.100 128.700 240.300 133.950 ;
        RECT 242.100 132.150 243.900 133.950 ;
        RECT 248.100 132.150 249.900 133.950 ;
        RECT 254.250 132.150 256.050 133.950 ;
        RECT 226.200 127.500 231.900 128.400 ;
        RECT 239.100 127.800 243.300 128.700 ;
        RECT 214.800 120.000 216.600 126.600 ;
        RECT 224.100 120.600 225.900 126.600 ;
        RECT 227.100 120.000 228.900 126.600 ;
        RECT 230.700 123.600 231.900 127.500 ;
        RECT 230.100 120.600 231.900 123.600 ;
        RECT 236.400 120.000 238.200 126.600 ;
        RECT 241.500 120.600 243.300 127.800 ;
        RECT 257.700 126.600 258.600 133.950 ;
        RECT 266.100 132.150 267.900 133.950 ;
        RECT 269.700 128.700 270.900 133.950 ;
        RECT 271.950 132.150 273.750 133.950 ;
        RECT 278.100 132.150 279.900 133.950 ;
        RECT 284.100 132.150 285.900 133.950 ;
        RECT 287.100 130.200 288.000 133.950 ;
        RECT 249.000 120.000 250.800 126.600 ;
        RECT 253.500 125.400 258.600 126.600 ;
        RECT 266.700 127.800 270.900 128.700 ;
        RECT 253.500 120.600 255.300 125.400 ;
        RECT 256.500 120.000 258.300 123.600 ;
        RECT 266.700 120.600 268.500 127.800 ;
        RECT 271.800 120.000 273.600 126.600 ;
        RECT 278.100 120.000 279.900 129.600 ;
        RECT 284.700 129.000 288.000 130.200 ;
        RECT 290.700 131.400 291.900 147.600 ;
        RECT 295.200 146.400 297.000 146.700 ;
        RECT 299.700 146.400 301.500 155.400 ;
        RECT 302.700 149.400 304.500 156.000 ;
        RECT 306.300 152.400 308.100 155.400 ;
        RECT 309.300 152.400 311.100 155.400 ;
        RECT 306.300 150.300 308.400 152.400 ;
        RECT 309.300 150.300 311.400 152.400 ;
        RECT 312.300 149.400 314.100 155.400 ;
        RECT 315.300 149.400 317.100 156.000 ;
        RECT 311.700 147.300 313.800 149.400 ;
        RECT 319.200 147.900 321.000 155.400 ;
        RECT 322.200 149.400 324.000 156.000 ;
        RECT 325.200 149.400 327.000 155.400 ;
        RECT 328.200 152.400 330.000 155.400 ;
        RECT 331.200 152.400 333.000 155.400 ;
        RECT 334.200 152.400 336.000 155.400 ;
        RECT 328.200 150.300 330.300 152.400 ;
        RECT 331.200 150.300 333.300 152.400 ;
        RECT 334.200 150.300 336.300 152.400 ;
        RECT 337.200 149.400 339.000 156.000 ;
        RECT 340.200 149.400 342.000 155.400 ;
        RECT 343.200 149.400 345.000 156.000 ;
        RECT 346.200 149.400 348.000 155.400 ;
        RECT 349.200 149.400 351.000 156.000 ;
        RECT 352.500 149.400 354.300 155.400 ;
        RECT 355.500 149.400 357.300 156.000 ;
        RECT 295.200 145.200 314.400 146.400 ;
        RECT 319.200 145.800 322.500 147.900 ;
        RECT 325.200 145.500 327.900 149.400 ;
        RECT 331.200 148.500 333.300 149.400 ;
        RECT 331.200 147.300 339.300 148.500 ;
        RECT 337.500 146.700 339.300 147.300 ;
        RECT 340.200 146.400 341.400 149.400 ;
        RECT 346.800 148.500 348.000 149.400 ;
        RECT 346.800 147.600 350.700 148.500 ;
        RECT 344.100 146.400 345.900 147.000 ;
        RECT 295.200 144.900 297.000 145.200 ;
        RECT 313.200 144.600 314.400 145.200 ;
        RECT 328.800 144.600 330.900 145.500 ;
        RECT 298.500 143.700 300.300 144.300 ;
        RECT 308.400 143.700 310.500 144.300 ;
        RECT 298.500 142.500 310.500 143.700 ;
        RECT 313.200 143.400 330.900 144.600 ;
        RECT 334.200 144.300 336.300 145.500 ;
        RECT 340.200 145.200 345.900 146.400 ;
        RECT 349.800 144.300 350.700 147.600 ;
        RECT 334.200 143.400 350.700 144.300 ;
        RECT 308.400 142.200 310.500 142.500 ;
        RECT 313.200 141.300 348.900 142.500 ;
        RECT 313.200 140.700 314.400 141.300 ;
        RECT 347.100 140.700 348.900 141.300 ;
        RECT 300.900 139.800 314.400 140.700 ;
        RECT 325.800 139.800 327.900 140.100 ;
        RECT 300.900 139.050 302.700 139.800 ;
        RECT 292.800 136.950 294.900 139.050 ;
        RECT 298.800 137.250 302.700 139.050 ;
        RECT 320.400 138.300 322.500 139.200 ;
        RECT 298.800 136.950 300.900 137.250 ;
        RECT 311.400 137.100 322.500 138.300 ;
        RECT 324.000 138.000 327.900 139.800 ;
        RECT 332.100 138.300 333.900 140.100 ;
        RECT 333.000 137.100 333.900 138.300 ;
        RECT 293.100 135.300 294.900 136.950 ;
        RECT 311.400 136.500 313.200 137.100 ;
        RECT 320.400 136.200 333.900 137.100 ;
        RECT 336.600 136.800 341.700 138.600 ;
        RECT 343.800 136.950 345.900 139.050 ;
        RECT 336.600 135.300 337.500 136.800 ;
        RECT 293.100 134.100 337.500 135.300 ;
        RECT 343.800 134.100 345.300 136.950 ;
        RECT 308.400 131.400 310.200 133.200 ;
        RECT 316.800 132.000 318.900 133.050 ;
        RECT 338.700 132.600 345.300 134.100 ;
        RECT 290.700 130.200 307.500 131.400 ;
        RECT 284.700 120.600 286.500 129.000 ;
        RECT 290.700 126.600 291.900 130.200 ;
        RECT 305.400 129.300 307.500 130.200 ;
        RECT 294.900 128.700 296.700 129.300 ;
        RECT 294.900 127.500 303.300 128.700 ;
        RECT 301.800 126.600 303.300 127.500 ;
        RECT 308.400 128.400 309.300 131.400 ;
        RECT 313.800 131.100 318.900 132.000 ;
        RECT 313.800 130.200 315.600 131.100 ;
        RECT 316.800 130.950 318.900 131.100 ;
        RECT 323.100 131.100 340.200 132.600 ;
        RECT 323.100 130.500 325.200 131.100 ;
        RECT 323.100 128.700 324.900 130.500 ;
        RECT 341.100 129.900 348.900 131.700 ;
        RECT 308.400 127.200 315.600 128.400 ;
        RECT 310.800 126.600 312.600 127.200 ;
        RECT 314.700 126.600 315.600 127.200 ;
        RECT 330.300 126.600 336.900 128.400 ;
        RECT 341.100 126.600 342.600 129.900 ;
        RECT 349.800 126.600 350.700 143.400 ;
        RECT 290.700 120.600 292.500 126.600 ;
        RECT 296.100 120.000 297.900 126.600 ;
        RECT 301.500 120.600 303.300 126.600 ;
        RECT 305.700 123.600 307.800 125.700 ;
        RECT 308.700 123.600 310.800 125.700 ;
        RECT 311.700 123.600 313.800 125.700 ;
        RECT 314.700 125.400 317.400 126.600 ;
        RECT 315.600 124.500 317.400 125.400 ;
        RECT 319.200 124.500 321.900 126.600 ;
        RECT 305.700 120.600 307.500 123.600 ;
        RECT 308.700 120.600 310.500 123.600 ;
        RECT 311.700 120.600 313.500 123.600 ;
        RECT 314.700 120.000 316.500 123.600 ;
        RECT 319.200 120.600 321.000 124.500 ;
        RECT 325.200 123.600 327.300 125.700 ;
        RECT 328.200 123.600 330.300 125.700 ;
        RECT 331.200 123.600 333.300 125.700 ;
        RECT 334.200 123.600 336.300 125.700 ;
        RECT 338.400 125.400 342.600 126.600 ;
        RECT 322.200 120.000 324.000 123.600 ;
        RECT 325.200 120.600 327.000 123.600 ;
        RECT 328.200 120.600 330.000 123.600 ;
        RECT 331.200 120.600 333.000 123.600 ;
        RECT 334.200 120.600 336.000 123.600 ;
        RECT 338.400 120.600 340.200 125.400 ;
        RECT 343.500 120.000 345.300 126.600 ;
        RECT 348.900 120.600 350.700 126.600 ;
        RECT 352.500 139.050 354.000 149.400 ;
        RECT 352.500 136.950 354.900 139.050 ;
        RECT 352.500 123.600 354.000 136.950 ;
        RECT 352.500 120.600 354.300 123.600 ;
        RECT 355.500 120.000 357.300 123.600 ;
        RECT 8.100 110.400 9.900 116.400 ;
        RECT 11.100 110.400 12.900 117.000 ;
        RECT 14.100 113.400 15.900 116.400 ;
        RECT 8.100 103.050 9.300 110.400 ;
        RECT 14.700 109.500 15.900 113.400 ;
        RECT 10.200 108.600 15.900 109.500 ;
        RECT 20.100 110.400 21.900 116.400 ;
        RECT 23.100 110.400 24.900 117.000 ;
        RECT 26.100 113.400 27.900 116.400 ;
        RECT 10.200 107.700 12.000 108.600 ;
        RECT 8.100 100.950 10.200 103.050 ;
        RECT 8.100 93.600 9.300 100.950 ;
        RECT 11.100 96.300 12.000 107.700 ;
        RECT 20.100 103.050 21.300 110.400 ;
        RECT 26.700 109.500 27.900 113.400 ;
        RECT 22.200 108.600 27.900 109.500 ;
        RECT 22.200 107.700 24.000 108.600 ;
        RECT 34.500 108.000 36.300 116.400 ;
        RECT 13.500 100.950 15.600 103.050 ;
        RECT 13.800 99.150 15.600 100.950 ;
        RECT 20.100 100.950 22.200 103.050 ;
        RECT 10.200 95.400 12.000 96.300 ;
        RECT 10.200 94.500 15.900 95.400 ;
        RECT 8.100 81.600 9.900 93.600 ;
        RECT 11.100 81.000 12.900 91.800 ;
        RECT 14.700 87.600 15.900 94.500 ;
        RECT 14.100 81.600 15.900 87.600 ;
        RECT 20.100 93.600 21.300 100.950 ;
        RECT 23.100 96.300 24.000 107.700 ;
        RECT 33.000 106.800 36.300 108.000 ;
        RECT 41.100 107.400 42.900 117.000 ;
        RECT 50.100 113.400 51.900 117.000 ;
        RECT 53.100 113.400 54.900 116.400 ;
        RECT 59.100 113.400 60.900 117.000 ;
        RECT 62.100 113.400 63.900 116.400 ;
        RECT 33.000 103.050 33.900 106.800 ;
        RECT 35.100 103.050 36.900 104.850 ;
        RECT 41.100 103.050 42.900 104.850 ;
        RECT 53.100 103.050 54.300 113.400 ;
        RECT 62.100 103.050 63.300 113.400 ;
        RECT 65.100 110.400 66.900 116.400 ;
        RECT 65.700 108.300 66.900 110.400 ;
        RECT 68.100 111.300 69.900 116.400 ;
        RECT 71.100 112.200 72.900 117.000 ;
        RECT 74.100 111.300 75.900 116.400 ;
        RECT 83.100 113.400 84.900 116.400 ;
        RECT 86.100 113.400 87.900 117.000 ;
        RECT 92.700 115.200 93.900 117.000 ;
        RECT 68.100 109.950 75.900 111.300 ;
        RECT 65.700 107.400 69.300 108.300 ;
        RECT 65.100 103.050 66.900 104.850 ;
        RECT 68.100 103.050 69.300 107.400 ;
        RECT 71.100 103.050 72.900 104.850 ;
        RECT 83.700 103.050 84.900 113.400 ;
        RECT 92.100 109.200 93.900 115.200 ;
        RECT 96.600 110.700 98.400 115.200 ;
        RECT 101.700 114.600 102.900 117.000 ;
        RECT 96.300 109.800 98.400 110.700 ;
        RECT 101.100 109.800 102.900 114.600 ;
        RECT 104.100 112.200 105.900 115.200 ;
        RECT 96.300 103.050 97.200 109.800 ;
        RECT 105.000 108.900 105.900 112.200 ;
        RECT 25.500 100.950 27.600 103.050 ;
        RECT 31.950 100.950 34.050 103.050 ;
        RECT 34.950 100.950 37.050 103.050 ;
        RECT 37.950 100.950 40.050 103.050 ;
        RECT 40.950 100.950 43.050 103.050 ;
        RECT 49.950 100.950 52.050 103.050 ;
        RECT 52.950 100.950 55.050 103.050 ;
        RECT 58.950 100.950 61.050 103.050 ;
        RECT 61.950 100.950 64.050 103.050 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 70.950 100.950 73.050 103.050 ;
        RECT 73.950 100.950 76.050 103.050 ;
        RECT 82.950 100.950 85.050 103.050 ;
        RECT 85.950 100.950 88.050 103.050 ;
        RECT 92.100 100.950 94.200 103.050 ;
        RECT 95.100 100.950 97.200 103.050 ;
        RECT 98.700 108.000 105.900 108.900 ;
        RECT 107.700 110.400 109.500 116.400 ;
        RECT 113.100 110.400 114.900 117.000 ;
        RECT 118.500 110.400 120.300 116.400 ;
        RECT 122.700 113.400 124.500 116.400 ;
        RECT 125.700 113.400 127.500 116.400 ;
        RECT 128.700 113.400 130.500 116.400 ;
        RECT 131.700 113.400 133.500 117.000 ;
        RECT 122.700 111.300 124.800 113.400 ;
        RECT 125.700 111.300 127.800 113.400 ;
        RECT 128.700 111.300 130.800 113.400 ;
        RECT 136.200 112.500 138.000 116.400 ;
        RECT 139.200 113.400 141.000 117.000 ;
        RECT 142.200 113.400 144.000 116.400 ;
        RECT 145.200 113.400 147.000 116.400 ;
        RECT 148.200 113.400 150.000 116.400 ;
        RECT 151.200 113.400 153.000 116.400 ;
        RECT 132.600 111.600 134.400 112.500 ;
        RECT 131.700 110.400 134.400 111.600 ;
        RECT 136.200 110.400 138.900 112.500 ;
        RECT 142.200 111.300 144.300 113.400 ;
        RECT 145.200 111.300 147.300 113.400 ;
        RECT 148.200 111.300 150.300 113.400 ;
        RECT 151.200 111.300 153.300 113.400 ;
        RECT 155.400 111.600 157.200 116.400 ;
        RECT 155.400 110.400 159.600 111.600 ;
        RECT 160.500 110.400 162.300 117.000 ;
        RECT 165.900 110.400 167.700 116.400 ;
        RECT 98.700 100.950 99.900 108.000 ;
        RECT 107.700 106.800 108.900 110.400 ;
        RECT 118.800 109.500 120.300 110.400 ;
        RECT 127.800 109.800 129.600 110.400 ;
        RECT 131.700 109.800 132.600 110.400 ;
        RECT 111.900 108.300 120.300 109.500 ;
        RECT 125.400 108.600 132.600 109.800 ;
        RECT 147.300 108.600 153.900 110.400 ;
        RECT 111.900 107.700 113.700 108.300 ;
        RECT 122.400 106.800 124.500 107.700 ;
        RECT 107.700 105.600 124.500 106.800 ;
        RECT 125.400 105.600 126.300 108.600 ;
        RECT 130.800 105.900 132.600 106.800 ;
        RECT 140.100 106.500 141.900 108.300 ;
        RECT 158.100 107.100 159.600 110.400 ;
        RECT 133.800 105.900 135.900 106.050 ;
        RECT 104.100 103.050 105.900 104.850 ;
        RECT 100.800 100.950 102.900 103.050 ;
        RECT 103.800 100.950 105.900 103.050 ;
        RECT 25.800 99.150 27.600 100.950 ;
        RECT 22.200 95.400 24.000 96.300 ;
        RECT 22.200 94.500 27.900 95.400 ;
        RECT 20.100 81.600 21.900 93.600 ;
        RECT 23.100 81.000 24.900 91.800 ;
        RECT 26.700 87.600 27.900 94.500 ;
        RECT 33.000 88.800 33.900 100.950 ;
        RECT 38.100 99.150 39.900 100.950 ;
        RECT 50.100 99.150 51.900 100.950 ;
        RECT 33.000 87.900 39.600 88.800 ;
        RECT 33.000 87.600 33.900 87.900 ;
        RECT 26.100 81.600 27.900 87.600 ;
        RECT 32.100 81.600 33.900 87.600 ;
        RECT 38.100 87.600 39.600 87.900 ;
        RECT 53.100 87.600 54.300 100.950 ;
        RECT 59.100 99.150 60.900 100.950 ;
        RECT 62.100 87.600 63.300 100.950 ;
        RECT 68.100 93.600 69.300 100.950 ;
        RECT 74.100 99.150 75.900 100.950 ;
        RECT 68.100 92.100 70.500 93.600 ;
        RECT 66.000 89.100 67.800 90.900 ;
        RECT 35.100 81.000 36.900 87.000 ;
        RECT 38.100 81.600 39.900 87.600 ;
        RECT 41.100 81.000 42.900 87.600 ;
        RECT 50.100 81.000 51.900 87.600 ;
        RECT 53.100 81.600 54.900 87.600 ;
        RECT 59.100 81.000 60.900 87.600 ;
        RECT 62.100 81.600 63.900 87.600 ;
        RECT 65.700 81.000 67.500 87.600 ;
        RECT 68.700 81.600 70.500 92.100 ;
        RECT 73.800 81.000 75.600 93.600 ;
        RECT 83.700 87.600 84.900 100.950 ;
        RECT 86.100 99.150 87.900 100.950 ;
        RECT 92.400 99.150 94.200 100.950 ;
        RECT 83.100 81.600 84.900 87.600 ;
        RECT 86.100 81.000 87.900 87.600 ;
        RECT 92.100 81.000 93.900 93.600 ;
        RECT 96.300 93.000 97.200 100.950 ;
        RECT 98.100 99.150 99.900 100.950 ;
        RECT 101.100 99.150 102.900 100.950 ;
        RECT 98.100 94.800 99.300 99.150 ;
        RECT 98.100 93.900 105.900 94.800 ;
        RECT 96.300 92.100 98.400 93.000 ;
        RECT 96.600 81.600 98.400 92.100 ;
        RECT 101.100 81.000 102.900 93.000 ;
        RECT 105.000 88.800 105.900 93.900 ;
        RECT 104.100 82.800 105.900 88.800 ;
        RECT 107.700 89.400 108.900 105.600 ;
        RECT 125.400 103.800 127.200 105.600 ;
        RECT 130.800 105.000 135.900 105.900 ;
        RECT 133.800 103.950 135.900 105.000 ;
        RECT 140.100 105.900 142.200 106.500 ;
        RECT 140.100 104.400 157.200 105.900 ;
        RECT 158.100 105.300 165.900 107.100 ;
        RECT 155.700 102.900 162.300 104.400 ;
        RECT 110.100 101.700 154.500 102.900 ;
        RECT 110.100 100.050 111.900 101.700 ;
        RECT 109.800 97.950 111.900 100.050 ;
        RECT 115.800 99.750 117.900 100.050 ;
        RECT 128.400 99.900 130.200 100.500 ;
        RECT 137.400 99.900 150.900 100.800 ;
        RECT 115.800 97.950 119.700 99.750 ;
        RECT 128.400 98.700 139.500 99.900 ;
        RECT 117.900 97.200 119.700 97.950 ;
        RECT 137.400 97.800 139.500 98.700 ;
        RECT 141.000 97.200 144.900 99.000 ;
        RECT 150.000 98.700 150.900 99.900 ;
        RECT 117.900 96.300 131.400 97.200 ;
        RECT 142.800 96.900 144.900 97.200 ;
        RECT 149.100 96.900 150.900 98.700 ;
        RECT 153.600 100.200 154.500 101.700 ;
        RECT 153.600 98.400 158.700 100.200 ;
        RECT 160.800 100.050 162.300 102.900 ;
        RECT 160.800 97.950 162.900 100.050 ;
        RECT 130.200 95.700 131.400 96.300 ;
        RECT 164.100 95.700 165.900 96.300 ;
        RECT 125.400 94.500 127.500 94.800 ;
        RECT 130.200 94.500 165.900 95.700 ;
        RECT 115.500 93.300 127.500 94.500 ;
        RECT 166.800 93.600 167.700 110.400 ;
        RECT 115.500 92.700 117.300 93.300 ;
        RECT 125.400 92.700 127.500 93.300 ;
        RECT 130.200 92.400 147.900 93.600 ;
        RECT 112.200 91.800 114.000 92.100 ;
        RECT 130.200 91.800 131.400 92.400 ;
        RECT 112.200 90.600 131.400 91.800 ;
        RECT 145.800 91.500 147.900 92.400 ;
        RECT 151.200 92.700 167.700 93.600 ;
        RECT 151.200 91.500 153.300 92.700 ;
        RECT 112.200 90.300 114.000 90.600 ;
        RECT 107.700 88.500 111.300 89.400 ;
        RECT 110.400 87.600 111.300 88.500 ;
        RECT 107.700 81.000 109.500 87.600 ;
        RECT 110.400 86.700 112.500 87.600 ;
        RECT 110.700 81.600 112.500 86.700 ;
        RECT 113.700 81.000 115.500 87.600 ;
        RECT 116.700 81.600 118.500 90.600 ;
        RECT 128.700 87.600 130.800 89.700 ;
        RECT 136.200 89.100 139.500 91.200 ;
        RECT 119.700 81.000 121.500 87.600 ;
        RECT 123.300 84.600 125.400 86.700 ;
        RECT 126.300 84.600 128.400 86.700 ;
        RECT 123.300 81.600 125.100 84.600 ;
        RECT 126.300 81.600 128.100 84.600 ;
        RECT 129.300 81.600 131.100 87.600 ;
        RECT 132.300 81.000 134.100 87.600 ;
        RECT 136.200 81.600 138.000 89.100 ;
        RECT 142.200 87.600 144.900 91.500 ;
        RECT 157.200 90.600 162.900 91.800 ;
        RECT 154.500 89.700 156.300 90.300 ;
        RECT 148.200 88.500 156.300 89.700 ;
        RECT 148.200 87.600 150.300 88.500 ;
        RECT 157.200 87.600 158.400 90.600 ;
        RECT 161.100 90.000 162.900 90.600 ;
        RECT 166.800 89.400 167.700 92.700 ;
        RECT 163.800 88.500 167.700 89.400 ;
        RECT 169.500 113.400 171.300 116.400 ;
        RECT 172.500 113.400 174.300 117.000 ;
        RECT 169.500 100.050 171.000 113.400 ;
        RECT 179.100 111.300 180.900 116.400 ;
        RECT 182.100 112.200 183.900 117.000 ;
        RECT 185.100 111.300 186.900 116.400 ;
        RECT 179.100 109.950 186.900 111.300 ;
        RECT 188.100 110.400 189.900 116.400 ;
        RECT 188.100 108.300 189.300 110.400 ;
        RECT 185.700 107.400 189.300 108.300 ;
        RECT 197.100 107.400 198.900 117.000 ;
        RECT 203.700 108.000 205.500 116.400 ;
        RECT 212.700 109.200 214.500 116.400 ;
        RECT 217.800 110.400 219.600 117.000 ;
        RECT 227.700 109.200 229.500 116.400 ;
        RECT 232.800 110.400 234.600 117.000 ;
        RECT 239.100 110.400 240.900 116.400 ;
        RECT 242.100 110.400 243.900 117.000 ;
        RECT 245.100 113.400 246.900 116.400 ;
        RECT 212.700 108.300 216.900 109.200 ;
        RECT 227.700 108.300 231.900 109.200 ;
        RECT 182.100 103.050 183.900 104.850 ;
        RECT 185.700 103.050 186.900 107.400 ;
        RECT 203.700 106.800 207.000 108.000 ;
        RECT 188.100 103.050 189.900 104.850 ;
        RECT 197.100 103.050 198.900 104.850 ;
        RECT 203.100 103.050 204.900 104.850 ;
        RECT 206.100 103.050 207.000 106.800 ;
        RECT 212.100 103.050 213.900 104.850 ;
        RECT 215.700 103.050 216.900 108.300 ;
        RECT 217.950 103.050 219.750 104.850 ;
        RECT 227.100 103.050 228.900 104.850 ;
        RECT 230.700 103.050 231.900 108.300 ;
        RECT 232.950 103.050 234.750 104.850 ;
        RECT 239.100 103.050 240.300 110.400 ;
        RECT 245.700 109.500 246.900 113.400 ;
        RECT 251.100 111.300 252.900 116.400 ;
        RECT 254.100 112.200 255.900 117.000 ;
        RECT 257.100 111.300 258.900 116.400 ;
        RECT 251.100 109.950 258.900 111.300 ;
        RECT 260.100 110.400 261.900 116.400 ;
        RECT 263.700 110.400 265.500 116.400 ;
        RECT 269.100 110.400 270.900 117.000 ;
        RECT 274.500 110.400 276.300 116.400 ;
        RECT 278.700 113.400 280.500 116.400 ;
        RECT 281.700 113.400 283.500 116.400 ;
        RECT 284.700 113.400 286.500 116.400 ;
        RECT 287.700 113.400 289.500 117.000 ;
        RECT 278.700 111.300 280.800 113.400 ;
        RECT 281.700 111.300 283.800 113.400 ;
        RECT 284.700 111.300 286.800 113.400 ;
        RECT 292.200 112.500 294.000 116.400 ;
        RECT 295.200 113.400 297.000 117.000 ;
        RECT 298.200 113.400 300.000 116.400 ;
        RECT 301.200 113.400 303.000 116.400 ;
        RECT 304.200 113.400 306.000 116.400 ;
        RECT 307.200 113.400 309.000 116.400 ;
        RECT 288.600 111.600 290.400 112.500 ;
        RECT 287.700 110.400 290.400 111.600 ;
        RECT 292.200 110.400 294.900 112.500 ;
        RECT 298.200 111.300 300.300 113.400 ;
        RECT 301.200 111.300 303.300 113.400 ;
        RECT 304.200 111.300 306.300 113.400 ;
        RECT 307.200 111.300 309.300 113.400 ;
        RECT 311.400 111.600 313.200 116.400 ;
        RECT 311.400 110.400 315.600 111.600 ;
        RECT 316.500 110.400 318.300 117.000 ;
        RECT 321.900 110.400 323.700 116.400 ;
        RECT 241.200 108.600 246.900 109.500 ;
        RECT 241.200 107.700 243.000 108.600 ;
        RECT 260.100 108.300 261.300 110.400 ;
        RECT 178.950 100.950 181.050 103.050 ;
        RECT 181.950 100.950 184.050 103.050 ;
        RECT 184.950 100.950 187.050 103.050 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 196.950 100.950 199.050 103.050 ;
        RECT 199.950 100.950 202.050 103.050 ;
        RECT 202.950 100.950 205.050 103.050 ;
        RECT 205.950 100.950 208.050 103.050 ;
        RECT 211.950 100.950 214.050 103.050 ;
        RECT 214.950 100.950 217.050 103.050 ;
        RECT 217.950 100.950 220.050 103.050 ;
        RECT 226.950 100.950 229.050 103.050 ;
        RECT 229.950 100.950 232.050 103.050 ;
        RECT 232.950 100.950 235.050 103.050 ;
        RECT 239.100 100.950 241.200 103.050 ;
        RECT 169.500 97.950 171.900 100.050 ;
        RECT 179.100 99.150 180.900 100.950 ;
        RECT 163.800 87.600 165.000 88.500 ;
        RECT 169.500 87.600 171.000 97.950 ;
        RECT 185.700 93.600 186.900 100.950 ;
        RECT 200.100 99.150 201.900 100.950 ;
        RECT 139.200 81.000 141.000 87.600 ;
        RECT 142.200 81.600 144.000 87.600 ;
        RECT 145.200 84.600 147.300 86.700 ;
        RECT 148.200 84.600 150.300 86.700 ;
        RECT 151.200 84.600 153.300 86.700 ;
        RECT 145.200 81.600 147.000 84.600 ;
        RECT 148.200 81.600 150.000 84.600 ;
        RECT 151.200 81.600 153.000 84.600 ;
        RECT 154.200 81.000 156.000 87.600 ;
        RECT 157.200 81.600 159.000 87.600 ;
        RECT 160.200 81.000 162.000 87.600 ;
        RECT 163.200 81.600 165.000 87.600 ;
        RECT 166.200 81.000 168.000 87.600 ;
        RECT 169.500 81.600 171.300 87.600 ;
        RECT 172.500 81.000 174.300 87.600 ;
        RECT 179.400 81.000 181.200 93.600 ;
        RECT 184.500 92.100 186.900 93.600 ;
        RECT 184.500 81.600 186.300 92.100 ;
        RECT 187.200 89.100 189.000 90.900 ;
        RECT 206.100 88.800 207.000 100.950 ;
        RECT 200.400 87.900 207.000 88.800 ;
        RECT 200.400 87.600 201.900 87.900 ;
        RECT 187.500 81.000 189.300 87.600 ;
        RECT 197.100 81.000 198.900 87.600 ;
        RECT 200.100 81.600 201.900 87.600 ;
        RECT 206.100 87.600 207.000 87.900 ;
        RECT 215.700 87.600 216.900 100.950 ;
        RECT 230.700 87.600 231.900 100.950 ;
        RECT 239.100 93.600 240.300 100.950 ;
        RECT 242.100 96.300 243.000 107.700 ;
        RECT 257.700 107.400 261.300 108.300 ;
        RECT 254.100 103.050 255.900 104.850 ;
        RECT 257.700 103.050 258.900 107.400 ;
        RECT 263.700 106.800 264.900 110.400 ;
        RECT 274.800 109.500 276.300 110.400 ;
        RECT 283.800 109.800 285.600 110.400 ;
        RECT 287.700 109.800 288.600 110.400 ;
        RECT 267.900 108.300 276.300 109.500 ;
        RECT 281.400 108.600 288.600 109.800 ;
        RECT 303.300 108.600 309.900 110.400 ;
        RECT 267.900 107.700 269.700 108.300 ;
        RECT 278.400 106.800 280.500 107.700 ;
        RECT 263.700 105.600 280.500 106.800 ;
        RECT 281.400 105.600 282.300 108.600 ;
        RECT 286.800 105.900 288.600 106.800 ;
        RECT 296.100 106.500 297.900 108.300 ;
        RECT 314.100 107.100 315.600 110.400 ;
        RECT 289.800 105.900 291.900 106.050 ;
        RECT 260.100 103.050 261.900 104.850 ;
        RECT 244.500 100.950 246.600 103.050 ;
        RECT 250.950 100.950 253.050 103.050 ;
        RECT 253.950 100.950 256.050 103.050 ;
        RECT 256.950 100.950 259.050 103.050 ;
        RECT 259.950 100.950 262.050 103.050 ;
        RECT 244.800 99.150 246.600 100.950 ;
        RECT 251.100 99.150 252.900 100.950 ;
        RECT 241.200 95.400 243.000 96.300 ;
        RECT 241.200 94.500 246.900 95.400 ;
        RECT 203.100 81.000 204.900 87.000 ;
        RECT 206.100 81.600 207.900 87.600 ;
        RECT 212.100 81.000 213.900 87.600 ;
        RECT 215.100 81.600 216.900 87.600 ;
        RECT 218.100 81.000 219.900 87.600 ;
        RECT 227.100 81.000 228.900 87.600 ;
        RECT 230.100 81.600 231.900 87.600 ;
        RECT 233.100 81.000 234.900 87.600 ;
        RECT 239.100 81.600 240.900 93.600 ;
        RECT 242.100 81.000 243.900 91.800 ;
        RECT 245.700 87.600 246.900 94.500 ;
        RECT 257.700 93.600 258.900 100.950 ;
        RECT 245.100 81.600 246.900 87.600 ;
        RECT 251.400 81.000 253.200 93.600 ;
        RECT 256.500 92.100 258.900 93.600 ;
        RECT 256.500 81.600 258.300 92.100 ;
        RECT 259.200 89.100 261.000 90.900 ;
        RECT 263.700 89.400 264.900 105.600 ;
        RECT 281.400 103.800 283.200 105.600 ;
        RECT 286.800 105.000 291.900 105.900 ;
        RECT 289.800 103.950 291.900 105.000 ;
        RECT 296.100 105.900 298.200 106.500 ;
        RECT 296.100 104.400 313.200 105.900 ;
        RECT 314.100 105.300 321.900 107.100 ;
        RECT 311.700 102.900 318.300 104.400 ;
        RECT 266.100 101.700 310.500 102.900 ;
        RECT 266.100 100.050 267.900 101.700 ;
        RECT 265.800 97.950 267.900 100.050 ;
        RECT 271.800 99.750 273.900 100.050 ;
        RECT 284.400 99.900 286.200 100.500 ;
        RECT 293.400 99.900 306.900 100.800 ;
        RECT 271.800 97.950 275.700 99.750 ;
        RECT 284.400 98.700 295.500 99.900 ;
        RECT 273.900 97.200 275.700 97.950 ;
        RECT 293.400 97.800 295.500 98.700 ;
        RECT 297.000 97.200 300.900 99.000 ;
        RECT 306.000 98.700 306.900 99.900 ;
        RECT 273.900 96.300 287.400 97.200 ;
        RECT 298.800 96.900 300.900 97.200 ;
        RECT 305.100 96.900 306.900 98.700 ;
        RECT 309.600 100.200 310.500 101.700 ;
        RECT 309.600 98.400 314.700 100.200 ;
        RECT 316.800 100.050 318.300 102.900 ;
        RECT 316.800 97.950 318.900 100.050 ;
        RECT 286.200 95.700 287.400 96.300 ;
        RECT 320.100 95.700 321.900 96.300 ;
        RECT 281.400 94.500 283.500 94.800 ;
        RECT 286.200 94.500 321.900 95.700 ;
        RECT 271.500 93.300 283.500 94.500 ;
        RECT 322.800 93.600 323.700 110.400 ;
        RECT 271.500 92.700 273.300 93.300 ;
        RECT 281.400 92.700 283.500 93.300 ;
        RECT 286.200 92.400 303.900 93.600 ;
        RECT 268.200 91.800 270.000 92.100 ;
        RECT 286.200 91.800 287.400 92.400 ;
        RECT 268.200 90.600 287.400 91.800 ;
        RECT 301.800 91.500 303.900 92.400 ;
        RECT 307.200 92.700 323.700 93.600 ;
        RECT 307.200 91.500 309.300 92.700 ;
        RECT 268.200 90.300 270.000 90.600 ;
        RECT 263.700 88.500 267.300 89.400 ;
        RECT 266.400 87.600 267.300 88.500 ;
        RECT 259.500 81.000 261.300 87.600 ;
        RECT 263.700 81.000 265.500 87.600 ;
        RECT 266.400 86.700 268.500 87.600 ;
        RECT 266.700 81.600 268.500 86.700 ;
        RECT 269.700 81.000 271.500 87.600 ;
        RECT 272.700 81.600 274.500 90.600 ;
        RECT 284.700 87.600 286.800 89.700 ;
        RECT 292.200 89.100 295.500 91.200 ;
        RECT 275.700 81.000 277.500 87.600 ;
        RECT 279.300 84.600 281.400 86.700 ;
        RECT 282.300 84.600 284.400 86.700 ;
        RECT 279.300 81.600 281.100 84.600 ;
        RECT 282.300 81.600 284.100 84.600 ;
        RECT 285.300 81.600 287.100 87.600 ;
        RECT 288.300 81.000 290.100 87.600 ;
        RECT 292.200 81.600 294.000 89.100 ;
        RECT 298.200 87.600 300.900 91.500 ;
        RECT 313.200 90.600 318.900 91.800 ;
        RECT 310.500 89.700 312.300 90.300 ;
        RECT 304.200 88.500 312.300 89.700 ;
        RECT 304.200 87.600 306.300 88.500 ;
        RECT 313.200 87.600 314.400 90.600 ;
        RECT 317.100 90.000 318.900 90.600 ;
        RECT 322.800 89.400 323.700 92.700 ;
        RECT 319.800 88.500 323.700 89.400 ;
        RECT 325.500 113.400 327.300 116.400 ;
        RECT 328.500 113.400 330.300 117.000 ;
        RECT 338.100 113.400 339.900 116.400 ;
        RECT 325.500 100.050 327.000 113.400 ;
        RECT 338.100 109.500 339.300 113.400 ;
        RECT 341.100 110.400 342.900 117.000 ;
        RECT 344.100 110.400 345.900 116.400 ;
        RECT 338.100 108.600 343.800 109.500 ;
        RECT 342.000 107.700 343.800 108.600 ;
        RECT 338.400 100.950 340.500 103.050 ;
        RECT 325.500 97.950 327.900 100.050 ;
        RECT 338.400 99.150 340.200 100.950 ;
        RECT 319.800 87.600 321.000 88.500 ;
        RECT 325.500 87.600 327.000 97.950 ;
        RECT 342.000 96.300 342.900 107.700 ;
        RECT 344.700 103.050 345.900 110.400 ;
        RECT 353.100 113.400 354.900 116.400 ;
        RECT 353.100 109.500 354.300 113.400 ;
        RECT 356.100 110.400 357.900 117.000 ;
        RECT 359.100 110.400 360.900 116.400 ;
        RECT 353.100 108.600 358.800 109.500 ;
        RECT 357.000 107.700 358.800 108.600 ;
        RECT 343.800 100.950 345.900 103.050 ;
        RECT 342.000 95.400 343.800 96.300 ;
        RECT 338.100 94.500 343.800 95.400 ;
        RECT 338.100 87.600 339.300 94.500 ;
        RECT 344.700 93.600 345.900 100.950 ;
        RECT 353.400 100.950 355.500 103.050 ;
        RECT 353.400 99.150 355.200 100.950 ;
        RECT 357.000 96.300 357.900 107.700 ;
        RECT 359.700 103.050 360.900 110.400 ;
        RECT 358.800 100.950 360.900 103.050 ;
        RECT 357.000 95.400 358.800 96.300 ;
        RECT 295.200 81.000 297.000 87.600 ;
        RECT 298.200 81.600 300.000 87.600 ;
        RECT 301.200 84.600 303.300 86.700 ;
        RECT 304.200 84.600 306.300 86.700 ;
        RECT 307.200 84.600 309.300 86.700 ;
        RECT 301.200 81.600 303.000 84.600 ;
        RECT 304.200 81.600 306.000 84.600 ;
        RECT 307.200 81.600 309.000 84.600 ;
        RECT 310.200 81.000 312.000 87.600 ;
        RECT 313.200 81.600 315.000 87.600 ;
        RECT 316.200 81.000 318.000 87.600 ;
        RECT 319.200 81.600 321.000 87.600 ;
        RECT 322.200 81.000 324.000 87.600 ;
        RECT 325.500 81.600 327.300 87.600 ;
        RECT 328.500 81.000 330.300 87.600 ;
        RECT 338.100 81.600 339.900 87.600 ;
        RECT 341.100 81.000 342.900 91.800 ;
        RECT 344.100 81.600 345.900 93.600 ;
        RECT 353.100 94.500 358.800 95.400 ;
        RECT 353.100 87.600 354.300 94.500 ;
        RECT 359.700 93.600 360.900 100.950 ;
        RECT 353.100 81.600 354.900 87.600 ;
        RECT 356.100 81.000 357.900 91.800 ;
        RECT 359.100 81.600 360.900 93.600 ;
        RECT 5.100 71.400 6.900 78.000 ;
        RECT 8.100 71.400 9.900 77.400 ;
        RECT 11.100 71.400 12.900 78.000 ;
        RECT 20.700 71.400 22.500 78.000 ;
        RECT 8.100 58.050 9.300 71.400 ;
        RECT 21.000 68.100 22.800 69.900 ;
        RECT 23.700 66.900 25.500 77.400 ;
        RECT 23.100 65.400 25.500 66.900 ;
        RECT 28.800 65.400 30.600 78.000 ;
        RECT 32.700 71.400 34.500 78.000 ;
        RECT 35.700 72.300 37.500 77.400 ;
        RECT 35.400 71.400 37.500 72.300 ;
        RECT 38.700 71.400 40.500 78.000 ;
        RECT 35.400 70.500 36.300 71.400 ;
        RECT 32.700 69.600 36.300 70.500 ;
        RECT 23.100 58.050 24.300 65.400 ;
        RECT 29.100 58.050 30.900 59.850 ;
        RECT 4.950 55.950 7.050 58.050 ;
        RECT 7.950 55.950 10.050 58.050 ;
        RECT 10.950 55.950 13.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 22.950 55.950 25.050 58.050 ;
        RECT 25.950 55.950 28.050 58.050 ;
        RECT 28.950 55.950 31.050 58.050 ;
        RECT 5.250 54.150 7.050 55.950 ;
        RECT 8.100 50.700 9.300 55.950 ;
        RECT 11.100 54.150 12.900 55.950 ;
        RECT 20.100 54.150 21.900 55.950 ;
        RECT 23.100 51.600 24.300 55.950 ;
        RECT 26.100 54.150 27.900 55.950 ;
        RECT 20.700 50.700 24.300 51.600 ;
        RECT 32.700 53.400 33.900 69.600 ;
        RECT 37.200 68.400 39.000 68.700 ;
        RECT 41.700 68.400 43.500 77.400 ;
        RECT 44.700 71.400 46.500 78.000 ;
        RECT 48.300 74.400 50.100 77.400 ;
        RECT 51.300 74.400 53.100 77.400 ;
        RECT 48.300 72.300 50.400 74.400 ;
        RECT 51.300 72.300 53.400 74.400 ;
        RECT 54.300 71.400 56.100 77.400 ;
        RECT 57.300 71.400 59.100 78.000 ;
        RECT 53.700 69.300 55.800 71.400 ;
        RECT 61.200 69.900 63.000 77.400 ;
        RECT 64.200 71.400 66.000 78.000 ;
        RECT 67.200 71.400 69.000 77.400 ;
        RECT 70.200 74.400 72.000 77.400 ;
        RECT 73.200 74.400 75.000 77.400 ;
        RECT 76.200 74.400 78.000 77.400 ;
        RECT 70.200 72.300 72.300 74.400 ;
        RECT 73.200 72.300 75.300 74.400 ;
        RECT 76.200 72.300 78.300 74.400 ;
        RECT 79.200 71.400 81.000 78.000 ;
        RECT 82.200 71.400 84.000 77.400 ;
        RECT 85.200 71.400 87.000 78.000 ;
        RECT 88.200 71.400 90.000 77.400 ;
        RECT 91.200 71.400 93.000 78.000 ;
        RECT 94.500 71.400 96.300 77.400 ;
        RECT 97.500 71.400 99.300 78.000 ;
        RECT 104.700 71.400 106.500 78.000 ;
        RECT 37.200 67.200 56.400 68.400 ;
        RECT 61.200 67.800 64.500 69.900 ;
        RECT 67.200 67.500 69.900 71.400 ;
        RECT 73.200 70.500 75.300 71.400 ;
        RECT 73.200 69.300 81.300 70.500 ;
        RECT 79.500 68.700 81.300 69.300 ;
        RECT 82.200 68.400 83.400 71.400 ;
        RECT 88.800 70.500 90.000 71.400 ;
        RECT 88.800 69.600 92.700 70.500 ;
        RECT 86.100 68.400 87.900 69.000 ;
        RECT 37.200 66.900 39.000 67.200 ;
        RECT 55.200 66.600 56.400 67.200 ;
        RECT 70.800 66.600 72.900 67.500 ;
        RECT 40.500 65.700 42.300 66.300 ;
        RECT 50.400 65.700 52.500 66.300 ;
        RECT 40.500 64.500 52.500 65.700 ;
        RECT 55.200 65.400 72.900 66.600 ;
        RECT 76.200 66.300 78.300 67.500 ;
        RECT 82.200 67.200 87.900 68.400 ;
        RECT 91.800 66.300 92.700 69.600 ;
        RECT 76.200 65.400 92.700 66.300 ;
        RECT 50.400 64.200 52.500 64.500 ;
        RECT 55.200 63.300 90.900 64.500 ;
        RECT 55.200 62.700 56.400 63.300 ;
        RECT 89.100 62.700 90.900 63.300 ;
        RECT 42.900 61.800 56.400 62.700 ;
        RECT 67.800 61.800 69.900 62.100 ;
        RECT 42.900 61.050 44.700 61.800 ;
        RECT 34.800 58.950 36.900 61.050 ;
        RECT 40.800 59.250 44.700 61.050 ;
        RECT 62.400 60.300 64.500 61.200 ;
        RECT 40.800 58.950 42.900 59.250 ;
        RECT 53.400 59.100 64.500 60.300 ;
        RECT 66.000 60.000 69.900 61.800 ;
        RECT 74.100 60.300 75.900 62.100 ;
        RECT 75.000 59.100 75.900 60.300 ;
        RECT 35.100 57.300 36.900 58.950 ;
        RECT 53.400 58.500 55.200 59.100 ;
        RECT 62.400 58.200 75.900 59.100 ;
        RECT 78.600 58.800 83.700 60.600 ;
        RECT 85.800 58.950 87.900 61.050 ;
        RECT 78.600 57.300 79.500 58.800 ;
        RECT 35.100 56.100 79.500 57.300 ;
        RECT 85.800 56.100 87.300 58.950 ;
        RECT 50.400 53.400 52.200 55.200 ;
        RECT 58.800 54.000 60.900 55.050 ;
        RECT 80.700 54.600 87.300 56.100 ;
        RECT 32.700 52.200 49.500 53.400 ;
        RECT 8.100 49.800 12.300 50.700 ;
        RECT 5.400 42.000 7.200 48.600 ;
        RECT 10.500 42.600 12.300 49.800 ;
        RECT 20.700 48.600 21.900 50.700 ;
        RECT 20.100 42.600 21.900 48.600 ;
        RECT 23.100 47.700 30.900 49.050 ;
        RECT 23.100 42.600 24.900 47.700 ;
        RECT 26.100 42.000 27.900 46.800 ;
        RECT 29.100 42.600 30.900 47.700 ;
        RECT 32.700 48.600 33.900 52.200 ;
        RECT 47.400 51.300 49.500 52.200 ;
        RECT 36.900 50.700 38.700 51.300 ;
        RECT 36.900 49.500 45.300 50.700 ;
        RECT 43.800 48.600 45.300 49.500 ;
        RECT 50.400 50.400 51.300 53.400 ;
        RECT 55.800 53.100 60.900 54.000 ;
        RECT 55.800 52.200 57.600 53.100 ;
        RECT 58.800 52.950 60.900 53.100 ;
        RECT 65.100 53.100 82.200 54.600 ;
        RECT 65.100 52.500 67.200 53.100 ;
        RECT 65.100 50.700 66.900 52.500 ;
        RECT 83.100 51.900 90.900 53.700 ;
        RECT 50.400 49.200 57.600 50.400 ;
        RECT 52.800 48.600 54.600 49.200 ;
        RECT 56.700 48.600 57.600 49.200 ;
        RECT 72.300 48.600 78.900 50.400 ;
        RECT 83.100 48.600 84.600 51.900 ;
        RECT 91.800 48.600 92.700 65.400 ;
        RECT 32.700 42.600 34.500 48.600 ;
        RECT 38.100 42.000 39.900 48.600 ;
        RECT 43.500 42.600 45.300 48.600 ;
        RECT 47.700 45.600 49.800 47.700 ;
        RECT 50.700 45.600 52.800 47.700 ;
        RECT 53.700 45.600 55.800 47.700 ;
        RECT 56.700 47.400 59.400 48.600 ;
        RECT 57.600 46.500 59.400 47.400 ;
        RECT 61.200 46.500 63.900 48.600 ;
        RECT 47.700 42.600 49.500 45.600 ;
        RECT 50.700 42.600 52.500 45.600 ;
        RECT 53.700 42.600 55.500 45.600 ;
        RECT 56.700 42.000 58.500 45.600 ;
        RECT 61.200 42.600 63.000 46.500 ;
        RECT 67.200 45.600 69.300 47.700 ;
        RECT 70.200 45.600 72.300 47.700 ;
        RECT 73.200 45.600 75.300 47.700 ;
        RECT 76.200 45.600 78.300 47.700 ;
        RECT 80.400 47.400 84.600 48.600 ;
        RECT 64.200 42.000 66.000 45.600 ;
        RECT 67.200 42.600 69.000 45.600 ;
        RECT 70.200 42.600 72.000 45.600 ;
        RECT 73.200 42.600 75.000 45.600 ;
        RECT 76.200 42.600 78.000 45.600 ;
        RECT 80.400 42.600 82.200 47.400 ;
        RECT 85.500 42.000 87.300 48.600 ;
        RECT 90.900 42.600 92.700 48.600 ;
        RECT 94.500 61.050 96.000 71.400 ;
        RECT 105.000 68.100 106.800 69.900 ;
        RECT 107.700 66.900 109.500 77.400 ;
        RECT 107.100 65.400 109.500 66.900 ;
        RECT 112.800 65.400 114.600 78.000 ;
        RECT 122.100 71.400 123.900 78.000 ;
        RECT 125.100 71.400 126.900 77.400 ;
        RECT 128.100 71.400 129.900 78.000 ;
        RECT 137.100 71.400 138.900 78.000 ;
        RECT 140.100 71.400 141.900 77.400 ;
        RECT 94.500 58.950 96.900 61.050 ;
        RECT 94.500 45.600 96.000 58.950 ;
        RECT 107.100 58.050 108.300 65.400 ;
        RECT 113.100 58.050 114.900 59.850 ;
        RECT 125.100 58.050 126.300 71.400 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 112.950 55.950 115.050 58.050 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 137.100 55.950 139.200 58.050 ;
        RECT 104.100 54.150 105.900 55.950 ;
        RECT 107.100 51.600 108.300 55.950 ;
        RECT 110.100 54.150 111.900 55.950 ;
        RECT 122.250 54.150 124.050 55.950 ;
        RECT 104.700 50.700 108.300 51.600 ;
        RECT 125.100 50.700 126.300 55.950 ;
        RECT 128.100 54.150 129.900 55.950 ;
        RECT 137.250 54.150 139.050 55.950 ;
        RECT 140.100 51.300 141.000 71.400 ;
        RECT 143.100 66.000 144.900 78.000 ;
        RECT 146.100 65.400 147.900 77.400 ;
        RECT 152.400 65.400 154.200 78.000 ;
        RECT 157.500 66.900 159.300 77.400 ;
        RECT 160.500 71.400 162.300 78.000 ;
        RECT 160.200 68.100 162.000 69.900 ;
        RECT 157.500 65.400 159.900 66.900 ;
        RECT 167.100 65.400 168.900 77.400 ;
        RECT 170.100 66.300 171.900 77.400 ;
        RECT 173.100 67.200 174.900 78.000 ;
        RECT 176.100 66.300 177.900 77.400 ;
        RECT 179.100 71.400 180.900 78.000 ;
        RECT 182.100 71.400 183.900 77.400 ;
        RECT 185.100 71.400 186.900 78.000 ;
        RECT 194.100 71.400 195.900 78.000 ;
        RECT 197.100 71.400 198.900 77.400 ;
        RECT 200.100 72.000 201.900 78.000 ;
        RECT 170.100 65.400 177.900 66.300 ;
        RECT 142.200 58.050 144.000 59.850 ;
        RECT 146.400 58.050 147.300 65.400 ;
        RECT 152.100 58.050 153.900 59.850 ;
        RECT 158.700 58.050 159.900 65.400 ;
        RECT 167.400 58.050 168.300 65.400 ;
        RECT 172.950 58.050 174.750 59.850 ;
        RECT 182.700 58.050 183.900 71.400 ;
        RECT 197.400 71.100 198.900 71.400 ;
        RECT 203.100 71.400 204.900 77.400 ;
        RECT 209.100 71.400 210.900 78.000 ;
        RECT 212.100 71.400 213.900 77.400 ;
        RECT 215.100 72.000 216.900 78.000 ;
        RECT 203.100 71.100 204.000 71.400 ;
        RECT 197.400 70.200 204.000 71.100 ;
        RECT 212.400 71.100 213.900 71.400 ;
        RECT 218.100 71.400 219.900 77.400 ;
        RECT 227.100 71.400 228.900 77.400 ;
        RECT 230.100 71.400 231.900 78.000 ;
        RECT 218.100 71.100 219.000 71.400 ;
        RECT 212.400 70.200 219.000 71.100 ;
        RECT 197.100 58.050 198.900 59.850 ;
        RECT 203.100 58.050 204.000 70.200 ;
        RECT 212.100 58.050 213.900 59.850 ;
        RECT 218.100 58.050 219.000 70.200 ;
        RECT 227.700 58.050 228.900 71.400 ;
        RECT 239.100 65.400 240.900 78.000 ;
        RECT 243.600 65.400 246.900 77.400 ;
        RECT 249.600 65.400 251.400 78.000 ;
        RECT 260.100 71.400 261.900 78.000 ;
        RECT 263.100 71.400 264.900 77.400 ;
        RECT 266.100 71.400 267.900 78.000 ;
        RECT 230.100 58.050 231.900 59.850 ;
        RECT 239.100 58.050 240.900 59.850 ;
        RECT 244.950 58.050 246.000 65.400 ;
        RECT 250.950 58.050 252.750 59.850 ;
        RECT 263.100 58.050 264.300 71.400 ;
        RECT 272.100 66.300 273.900 77.400 ;
        RECT 275.100 67.200 276.900 78.000 ;
        RECT 278.100 66.300 279.900 77.400 ;
        RECT 272.100 65.400 279.900 66.300 ;
        RECT 281.100 65.400 282.900 77.400 ;
        RECT 284.700 71.400 286.500 78.000 ;
        RECT 287.700 72.300 289.500 77.400 ;
        RECT 287.400 71.400 289.500 72.300 ;
        RECT 290.700 71.400 292.500 78.000 ;
        RECT 287.400 70.500 288.300 71.400 ;
        RECT 284.700 69.600 288.300 70.500 ;
        RECT 275.250 58.050 277.050 59.850 ;
        RECT 281.700 58.050 282.600 65.400 ;
        RECT 142.500 55.950 144.600 58.050 ;
        RECT 145.800 55.950 147.900 58.050 ;
        RECT 151.950 55.950 154.050 58.050 ;
        RECT 154.950 55.950 157.050 58.050 ;
        RECT 157.950 55.950 160.050 58.050 ;
        RECT 160.950 55.950 163.050 58.050 ;
        RECT 166.950 55.950 169.050 58.050 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 172.950 55.950 175.050 58.050 ;
        RECT 175.950 55.950 178.050 58.050 ;
        RECT 178.950 55.950 181.050 58.050 ;
        RECT 181.950 55.950 184.050 58.050 ;
        RECT 184.950 55.950 187.050 58.050 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 196.950 55.950 199.050 58.050 ;
        RECT 199.950 55.950 202.050 58.050 ;
        RECT 202.950 55.950 205.050 58.050 ;
        RECT 208.950 55.950 211.050 58.050 ;
        RECT 211.950 55.950 214.050 58.050 ;
        RECT 214.950 55.950 217.050 58.050 ;
        RECT 217.950 55.950 220.050 58.050 ;
        RECT 226.950 55.950 229.050 58.050 ;
        RECT 229.950 55.950 232.050 58.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 241.950 55.950 244.050 58.050 ;
        RECT 104.700 48.600 105.900 50.700 ;
        RECT 125.100 49.800 129.300 50.700 ;
        RECT 94.500 42.600 96.300 45.600 ;
        RECT 97.500 42.000 99.300 45.600 ;
        RECT 104.100 42.600 105.900 48.600 ;
        RECT 107.100 47.700 114.900 49.050 ;
        RECT 107.100 42.600 108.900 47.700 ;
        RECT 110.100 42.000 111.900 46.800 ;
        RECT 113.100 42.600 114.900 47.700 ;
        RECT 122.400 42.000 124.200 48.600 ;
        RECT 127.500 42.600 129.300 49.800 ;
        RECT 137.100 50.400 145.500 51.300 ;
        RECT 137.100 42.600 138.900 50.400 ;
        RECT 143.700 49.500 145.500 50.400 ;
        RECT 146.400 48.600 147.300 55.950 ;
        RECT 155.100 54.150 156.900 55.950 ;
        RECT 158.700 51.600 159.900 55.950 ;
        RECT 161.100 54.150 162.900 55.950 ;
        RECT 158.700 50.700 162.300 51.600 ;
        RECT 141.600 42.000 143.400 48.600 ;
        RECT 144.600 46.800 147.300 48.600 ;
        RECT 152.100 47.700 159.900 49.050 ;
        RECT 144.600 42.600 146.400 46.800 ;
        RECT 152.100 42.600 153.900 47.700 ;
        RECT 155.100 42.000 156.900 46.800 ;
        RECT 158.100 42.600 159.900 47.700 ;
        RECT 161.100 48.600 162.300 50.700 ;
        RECT 167.400 48.600 168.300 55.950 ;
        RECT 169.950 54.150 171.750 55.950 ;
        RECT 176.100 54.150 177.900 55.950 ;
        RECT 179.100 54.150 180.900 55.950 ;
        RECT 182.700 50.700 183.900 55.950 ;
        RECT 184.950 54.150 186.750 55.950 ;
        RECT 194.100 54.150 195.900 55.950 ;
        RECT 200.100 54.150 201.900 55.950 ;
        RECT 203.100 52.200 204.000 55.950 ;
        RECT 209.100 54.150 210.900 55.950 ;
        RECT 215.100 54.150 216.900 55.950 ;
        RECT 218.100 52.200 219.000 55.950 ;
        RECT 179.700 49.800 183.900 50.700 ;
        RECT 161.100 42.600 162.900 48.600 ;
        RECT 167.400 47.400 172.500 48.600 ;
        RECT 167.700 42.000 169.500 45.600 ;
        RECT 170.700 42.600 172.500 47.400 ;
        RECT 175.200 42.000 177.000 48.600 ;
        RECT 179.700 42.600 181.500 49.800 ;
        RECT 184.800 42.000 186.600 48.600 ;
        RECT 194.100 42.000 195.900 51.600 ;
        RECT 200.700 51.000 204.000 52.200 ;
        RECT 200.700 42.600 202.500 51.000 ;
        RECT 209.100 42.000 210.900 51.600 ;
        RECT 215.700 51.000 219.000 52.200 ;
        RECT 215.700 42.600 217.500 51.000 ;
        RECT 227.700 45.600 228.900 55.950 ;
        RECT 242.250 54.150 244.050 55.950 ;
        RECT 244.950 55.950 247.050 58.050 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 250.950 55.950 253.050 58.050 ;
        RECT 259.950 55.950 262.050 58.050 ;
        RECT 262.950 55.950 265.050 58.050 ;
        RECT 265.950 55.950 268.050 58.050 ;
        RECT 271.950 55.950 274.050 58.050 ;
        RECT 274.950 55.950 277.050 58.050 ;
        RECT 277.950 55.950 280.050 58.050 ;
        RECT 280.950 55.950 283.050 58.050 ;
        RECT 244.950 51.300 246.000 55.950 ;
        RECT 247.950 54.150 249.750 55.950 ;
        RECT 260.250 54.150 262.050 55.950 ;
        RECT 250.950 51.450 253.050 52.050 ;
        RECT 259.950 51.450 262.050 52.050 ;
        RECT 244.950 50.100 249.300 51.300 ;
        RECT 239.100 48.000 246.900 48.900 ;
        RECT 248.400 48.600 249.300 50.100 ;
        RECT 250.950 50.550 262.050 51.450 ;
        RECT 250.950 49.950 253.050 50.550 ;
        RECT 259.950 49.950 262.050 50.550 ;
        RECT 263.100 50.700 264.300 55.950 ;
        RECT 266.100 54.150 267.900 55.950 ;
        RECT 272.100 54.150 273.900 55.950 ;
        RECT 278.250 54.150 280.050 55.950 ;
        RECT 263.100 49.800 267.300 50.700 ;
        RECT 227.100 42.600 228.900 45.600 ;
        RECT 230.100 42.000 231.900 45.600 ;
        RECT 239.100 42.600 240.900 48.000 ;
        RECT 242.100 42.000 243.900 47.100 ;
        RECT 245.100 43.500 246.900 48.000 ;
        RECT 248.100 44.400 249.900 48.600 ;
        RECT 251.100 43.500 252.900 48.600 ;
        RECT 245.100 42.600 252.900 43.500 ;
        RECT 260.400 42.000 262.200 48.600 ;
        RECT 265.500 42.600 267.300 49.800 ;
        RECT 281.700 48.600 282.600 55.950 ;
        RECT 273.000 42.000 274.800 48.600 ;
        RECT 277.500 47.400 282.600 48.600 ;
        RECT 284.700 53.400 285.900 69.600 ;
        RECT 289.200 68.400 291.000 68.700 ;
        RECT 293.700 68.400 295.500 77.400 ;
        RECT 296.700 71.400 298.500 78.000 ;
        RECT 300.300 74.400 302.100 77.400 ;
        RECT 303.300 74.400 305.100 77.400 ;
        RECT 300.300 72.300 302.400 74.400 ;
        RECT 303.300 72.300 305.400 74.400 ;
        RECT 306.300 71.400 308.100 77.400 ;
        RECT 309.300 71.400 311.100 78.000 ;
        RECT 305.700 69.300 307.800 71.400 ;
        RECT 313.200 69.900 315.000 77.400 ;
        RECT 316.200 71.400 318.000 78.000 ;
        RECT 319.200 71.400 321.000 77.400 ;
        RECT 322.200 74.400 324.000 77.400 ;
        RECT 325.200 74.400 327.000 77.400 ;
        RECT 328.200 74.400 330.000 77.400 ;
        RECT 322.200 72.300 324.300 74.400 ;
        RECT 325.200 72.300 327.300 74.400 ;
        RECT 328.200 72.300 330.300 74.400 ;
        RECT 331.200 71.400 333.000 78.000 ;
        RECT 334.200 71.400 336.000 77.400 ;
        RECT 337.200 71.400 339.000 78.000 ;
        RECT 340.200 71.400 342.000 77.400 ;
        RECT 343.200 71.400 345.000 78.000 ;
        RECT 346.500 71.400 348.300 77.400 ;
        RECT 349.500 71.400 351.300 78.000 ;
        RECT 289.200 67.200 308.400 68.400 ;
        RECT 313.200 67.800 316.500 69.900 ;
        RECT 319.200 67.500 321.900 71.400 ;
        RECT 325.200 70.500 327.300 71.400 ;
        RECT 325.200 69.300 333.300 70.500 ;
        RECT 331.500 68.700 333.300 69.300 ;
        RECT 334.200 68.400 335.400 71.400 ;
        RECT 340.800 70.500 342.000 71.400 ;
        RECT 340.800 69.600 344.700 70.500 ;
        RECT 338.100 68.400 339.900 69.000 ;
        RECT 289.200 66.900 291.000 67.200 ;
        RECT 307.200 66.600 308.400 67.200 ;
        RECT 322.800 66.600 324.900 67.500 ;
        RECT 292.500 65.700 294.300 66.300 ;
        RECT 302.400 65.700 304.500 66.300 ;
        RECT 292.500 64.500 304.500 65.700 ;
        RECT 307.200 65.400 324.900 66.600 ;
        RECT 328.200 66.300 330.300 67.500 ;
        RECT 334.200 67.200 339.900 68.400 ;
        RECT 343.800 66.300 344.700 69.600 ;
        RECT 328.200 65.400 344.700 66.300 ;
        RECT 302.400 64.200 304.500 64.500 ;
        RECT 307.200 63.300 342.900 64.500 ;
        RECT 307.200 62.700 308.400 63.300 ;
        RECT 341.100 62.700 342.900 63.300 ;
        RECT 294.900 61.800 308.400 62.700 ;
        RECT 319.800 61.800 321.900 62.100 ;
        RECT 294.900 61.050 296.700 61.800 ;
        RECT 286.800 58.950 288.900 61.050 ;
        RECT 292.800 59.250 296.700 61.050 ;
        RECT 314.400 60.300 316.500 61.200 ;
        RECT 292.800 58.950 294.900 59.250 ;
        RECT 305.400 59.100 316.500 60.300 ;
        RECT 318.000 60.000 321.900 61.800 ;
        RECT 326.100 60.300 327.900 62.100 ;
        RECT 327.000 59.100 327.900 60.300 ;
        RECT 287.100 57.300 288.900 58.950 ;
        RECT 305.400 58.500 307.200 59.100 ;
        RECT 314.400 58.200 327.900 59.100 ;
        RECT 330.600 58.800 335.700 60.600 ;
        RECT 337.800 58.950 339.900 61.050 ;
        RECT 330.600 57.300 331.500 58.800 ;
        RECT 287.100 56.100 331.500 57.300 ;
        RECT 337.800 56.100 339.300 58.950 ;
        RECT 302.400 53.400 304.200 55.200 ;
        RECT 310.800 54.000 312.900 55.050 ;
        RECT 332.700 54.600 339.300 56.100 ;
        RECT 284.700 52.200 301.500 53.400 ;
        RECT 284.700 48.600 285.900 52.200 ;
        RECT 299.400 51.300 301.500 52.200 ;
        RECT 288.900 50.700 290.700 51.300 ;
        RECT 288.900 49.500 297.300 50.700 ;
        RECT 295.800 48.600 297.300 49.500 ;
        RECT 302.400 50.400 303.300 53.400 ;
        RECT 307.800 53.100 312.900 54.000 ;
        RECT 307.800 52.200 309.600 53.100 ;
        RECT 310.800 52.950 312.900 53.100 ;
        RECT 317.100 53.100 334.200 54.600 ;
        RECT 317.100 52.500 319.200 53.100 ;
        RECT 317.100 50.700 318.900 52.500 ;
        RECT 335.100 51.900 342.900 53.700 ;
        RECT 302.400 49.200 309.600 50.400 ;
        RECT 304.800 48.600 306.600 49.200 ;
        RECT 308.700 48.600 309.600 49.200 ;
        RECT 324.300 48.600 330.900 50.400 ;
        RECT 335.100 48.600 336.600 51.900 ;
        RECT 343.800 48.600 344.700 65.400 ;
        RECT 277.500 42.600 279.300 47.400 ;
        RECT 280.500 42.000 282.300 45.600 ;
        RECT 284.700 42.600 286.500 48.600 ;
        RECT 290.100 42.000 291.900 48.600 ;
        RECT 295.500 42.600 297.300 48.600 ;
        RECT 299.700 45.600 301.800 47.700 ;
        RECT 302.700 45.600 304.800 47.700 ;
        RECT 305.700 45.600 307.800 47.700 ;
        RECT 308.700 47.400 311.400 48.600 ;
        RECT 309.600 46.500 311.400 47.400 ;
        RECT 313.200 46.500 315.900 48.600 ;
        RECT 299.700 42.600 301.500 45.600 ;
        RECT 302.700 42.600 304.500 45.600 ;
        RECT 305.700 42.600 307.500 45.600 ;
        RECT 308.700 42.000 310.500 45.600 ;
        RECT 313.200 42.600 315.000 46.500 ;
        RECT 319.200 45.600 321.300 47.700 ;
        RECT 322.200 45.600 324.300 47.700 ;
        RECT 325.200 45.600 327.300 47.700 ;
        RECT 328.200 45.600 330.300 47.700 ;
        RECT 332.400 47.400 336.600 48.600 ;
        RECT 316.200 42.000 318.000 45.600 ;
        RECT 319.200 42.600 321.000 45.600 ;
        RECT 322.200 42.600 324.000 45.600 ;
        RECT 325.200 42.600 327.000 45.600 ;
        RECT 328.200 42.600 330.000 45.600 ;
        RECT 332.400 42.600 334.200 47.400 ;
        RECT 337.500 42.000 339.300 48.600 ;
        RECT 342.900 42.600 344.700 48.600 ;
        RECT 346.500 61.050 348.000 71.400 ;
        RECT 346.500 58.950 348.900 61.050 ;
        RECT 346.500 45.600 348.000 58.950 ;
        RECT 346.500 42.600 348.300 45.600 ;
        RECT 349.500 42.000 351.300 45.600 ;
        RECT 5.100 32.400 6.900 38.400 ;
        RECT 8.100 32.400 9.900 39.000 ;
        RECT 11.100 35.400 12.900 38.400 ;
        RECT 5.100 25.050 6.300 32.400 ;
        RECT 11.700 31.500 12.900 35.400 ;
        RECT 7.200 30.600 12.900 31.500 ;
        RECT 14.700 32.400 16.500 38.400 ;
        RECT 20.100 32.400 21.900 39.000 ;
        RECT 25.500 32.400 27.300 38.400 ;
        RECT 29.700 35.400 31.500 38.400 ;
        RECT 32.700 35.400 34.500 38.400 ;
        RECT 35.700 35.400 37.500 38.400 ;
        RECT 38.700 35.400 40.500 39.000 ;
        RECT 29.700 33.300 31.800 35.400 ;
        RECT 32.700 33.300 34.800 35.400 ;
        RECT 35.700 33.300 37.800 35.400 ;
        RECT 43.200 34.500 45.000 38.400 ;
        RECT 46.200 35.400 48.000 39.000 ;
        RECT 49.200 35.400 51.000 38.400 ;
        RECT 52.200 35.400 54.000 38.400 ;
        RECT 55.200 35.400 57.000 38.400 ;
        RECT 58.200 35.400 60.000 38.400 ;
        RECT 39.600 33.600 41.400 34.500 ;
        RECT 38.700 32.400 41.400 33.600 ;
        RECT 43.200 32.400 45.900 34.500 ;
        RECT 49.200 33.300 51.300 35.400 ;
        RECT 52.200 33.300 54.300 35.400 ;
        RECT 55.200 33.300 57.300 35.400 ;
        RECT 58.200 33.300 60.300 35.400 ;
        RECT 62.400 33.600 64.200 38.400 ;
        RECT 62.400 32.400 66.600 33.600 ;
        RECT 67.500 32.400 69.300 39.000 ;
        RECT 72.900 32.400 74.700 38.400 ;
        RECT 7.200 29.700 9.000 30.600 ;
        RECT 5.100 22.950 7.200 25.050 ;
        RECT 5.100 15.600 6.300 22.950 ;
        RECT 8.100 18.300 9.000 29.700 ;
        RECT 14.700 28.800 15.900 32.400 ;
        RECT 25.800 31.500 27.300 32.400 ;
        RECT 34.800 31.800 36.600 32.400 ;
        RECT 38.700 31.800 39.600 32.400 ;
        RECT 18.900 30.300 27.300 31.500 ;
        RECT 32.400 30.600 39.600 31.800 ;
        RECT 54.300 30.600 60.900 32.400 ;
        RECT 18.900 29.700 20.700 30.300 ;
        RECT 29.400 28.800 31.500 29.700 ;
        RECT 14.700 27.600 31.500 28.800 ;
        RECT 32.400 27.600 33.300 30.600 ;
        RECT 37.800 27.900 39.600 28.800 ;
        RECT 47.100 28.500 48.900 30.300 ;
        RECT 65.100 29.100 66.600 32.400 ;
        RECT 40.800 27.900 42.900 28.050 ;
        RECT 10.500 22.950 12.600 25.050 ;
        RECT 10.800 21.150 12.600 22.950 ;
        RECT 7.200 17.400 9.000 18.300 ;
        RECT 7.200 16.500 12.900 17.400 ;
        RECT 5.100 3.600 6.900 15.600 ;
        RECT 8.100 3.000 9.900 13.800 ;
        RECT 11.700 9.600 12.900 16.500 ;
        RECT 14.700 11.400 15.900 27.600 ;
        RECT 32.400 25.800 34.200 27.600 ;
        RECT 37.800 27.000 42.900 27.900 ;
        RECT 40.800 25.950 42.900 27.000 ;
        RECT 47.100 27.900 49.200 28.500 ;
        RECT 47.100 26.400 64.200 27.900 ;
        RECT 65.100 27.300 72.900 29.100 ;
        RECT 62.700 24.900 69.300 26.400 ;
        RECT 17.100 23.700 61.500 24.900 ;
        RECT 17.100 22.050 18.900 23.700 ;
        RECT 16.800 19.950 18.900 22.050 ;
        RECT 22.800 21.750 24.900 22.050 ;
        RECT 35.400 21.900 37.200 22.500 ;
        RECT 44.400 21.900 57.900 22.800 ;
        RECT 22.800 19.950 26.700 21.750 ;
        RECT 35.400 20.700 46.500 21.900 ;
        RECT 24.900 19.200 26.700 19.950 ;
        RECT 44.400 19.800 46.500 20.700 ;
        RECT 48.000 19.200 51.900 21.000 ;
        RECT 57.000 20.700 57.900 21.900 ;
        RECT 24.900 18.300 38.400 19.200 ;
        RECT 49.800 18.900 51.900 19.200 ;
        RECT 56.100 18.900 57.900 20.700 ;
        RECT 60.600 22.200 61.500 23.700 ;
        RECT 60.600 20.400 65.700 22.200 ;
        RECT 67.800 22.050 69.300 24.900 ;
        RECT 67.800 19.950 69.900 22.050 ;
        RECT 37.200 17.700 38.400 18.300 ;
        RECT 71.100 17.700 72.900 18.300 ;
        RECT 32.400 16.500 34.500 16.800 ;
        RECT 37.200 16.500 72.900 17.700 ;
        RECT 22.500 15.300 34.500 16.500 ;
        RECT 73.800 15.600 74.700 32.400 ;
        RECT 22.500 14.700 24.300 15.300 ;
        RECT 32.400 14.700 34.500 15.300 ;
        RECT 37.200 14.400 54.900 15.600 ;
        RECT 19.200 13.800 21.000 14.100 ;
        RECT 37.200 13.800 38.400 14.400 ;
        RECT 19.200 12.600 38.400 13.800 ;
        RECT 52.800 13.500 54.900 14.400 ;
        RECT 58.200 14.700 74.700 15.600 ;
        RECT 58.200 13.500 60.300 14.700 ;
        RECT 19.200 12.300 21.000 12.600 ;
        RECT 14.700 10.500 18.300 11.400 ;
        RECT 17.400 9.600 18.300 10.500 ;
        RECT 11.100 3.600 12.900 9.600 ;
        RECT 14.700 3.000 16.500 9.600 ;
        RECT 17.400 8.700 19.500 9.600 ;
        RECT 17.700 3.600 19.500 8.700 ;
        RECT 20.700 3.000 22.500 9.600 ;
        RECT 23.700 3.600 25.500 12.600 ;
        RECT 35.700 9.600 37.800 11.700 ;
        RECT 43.200 11.100 46.500 13.200 ;
        RECT 26.700 3.000 28.500 9.600 ;
        RECT 30.300 6.600 32.400 8.700 ;
        RECT 33.300 6.600 35.400 8.700 ;
        RECT 30.300 3.600 32.100 6.600 ;
        RECT 33.300 3.600 35.100 6.600 ;
        RECT 36.300 3.600 38.100 9.600 ;
        RECT 39.300 3.000 41.100 9.600 ;
        RECT 43.200 3.600 45.000 11.100 ;
        RECT 49.200 9.600 51.900 13.500 ;
        RECT 64.200 12.600 69.900 13.800 ;
        RECT 61.500 11.700 63.300 12.300 ;
        RECT 55.200 10.500 63.300 11.700 ;
        RECT 55.200 9.600 57.300 10.500 ;
        RECT 64.200 9.600 65.400 12.600 ;
        RECT 68.100 12.000 69.900 12.600 ;
        RECT 73.800 11.400 74.700 14.700 ;
        RECT 70.800 10.500 74.700 11.400 ;
        RECT 76.500 35.400 78.300 38.400 ;
        RECT 79.500 35.400 81.300 39.000 ;
        RECT 76.500 22.050 78.000 35.400 ;
        RECT 89.100 32.400 90.900 38.400 ;
        RECT 92.100 32.400 93.900 39.000 ;
        RECT 95.100 35.400 96.900 38.400 ;
        RECT 89.100 25.050 90.300 32.400 ;
        RECT 95.700 31.500 96.900 35.400 ;
        RECT 91.200 30.600 96.900 31.500 ;
        RECT 104.100 34.200 105.900 37.200 ;
        RECT 107.100 36.600 108.300 39.000 ;
        RECT 116.100 37.200 117.300 39.000 ;
        RECT 104.100 30.900 105.000 34.200 ;
        RECT 107.100 31.800 108.900 36.600 ;
        RECT 111.600 32.700 113.400 37.200 ;
        RECT 111.600 31.800 113.700 32.700 ;
        RECT 91.200 29.700 93.000 30.600 ;
        RECT 104.100 30.000 111.300 30.900 ;
        RECT 89.100 22.950 91.200 25.050 ;
        RECT 76.500 19.950 78.900 22.050 ;
        RECT 70.800 9.600 72.000 10.500 ;
        RECT 76.500 9.600 78.000 19.950 ;
        RECT 89.100 15.600 90.300 22.950 ;
        RECT 92.100 18.300 93.000 29.700 ;
        RECT 104.100 25.050 105.900 26.850 ;
        RECT 94.500 22.950 96.600 25.050 ;
        RECT 104.100 22.950 106.200 25.050 ;
        RECT 107.100 22.950 109.200 25.050 ;
        RECT 110.100 22.950 111.300 30.000 ;
        RECT 112.800 25.050 113.700 31.800 ;
        RECT 116.100 31.200 117.900 37.200 ;
        RECT 122.100 35.400 123.900 38.400 ;
        RECT 125.100 35.400 126.900 39.000 ;
        RECT 122.700 25.050 123.900 35.400 ;
        RECT 128.100 32.400 129.900 38.400 ;
        RECT 131.100 32.400 132.900 39.000 ;
        RECT 134.100 35.400 135.900 38.400 ;
        RECT 143.100 35.400 144.900 39.000 ;
        RECT 146.100 35.400 147.900 38.400 ;
        RECT 155.100 35.400 156.900 39.000 ;
        RECT 158.100 35.400 159.900 38.400 ;
        RECT 161.100 35.400 162.900 39.000 ;
        RECT 128.100 25.050 129.300 32.400 ;
        RECT 134.700 31.500 135.900 35.400 ;
        RECT 130.200 30.600 135.900 31.500 ;
        RECT 130.200 29.700 132.000 30.600 ;
        RECT 112.800 22.950 114.900 25.050 ;
        RECT 115.800 22.950 117.900 25.050 ;
        RECT 121.950 22.950 124.050 25.050 ;
        RECT 124.950 22.950 127.050 25.050 ;
        RECT 128.100 22.950 130.200 25.050 ;
        RECT 94.800 21.150 96.600 22.950 ;
        RECT 107.100 21.150 108.900 22.950 ;
        RECT 110.100 21.150 111.900 22.950 ;
        RECT 91.200 17.400 93.000 18.300 ;
        RECT 91.200 16.500 96.900 17.400 ;
        RECT 110.700 16.800 111.900 21.150 ;
        RECT 46.200 3.000 48.000 9.600 ;
        RECT 49.200 3.600 51.000 9.600 ;
        RECT 52.200 6.600 54.300 8.700 ;
        RECT 55.200 6.600 57.300 8.700 ;
        RECT 58.200 6.600 60.300 8.700 ;
        RECT 52.200 3.600 54.000 6.600 ;
        RECT 55.200 3.600 57.000 6.600 ;
        RECT 58.200 3.600 60.000 6.600 ;
        RECT 61.200 3.000 63.000 9.600 ;
        RECT 64.200 3.600 66.000 9.600 ;
        RECT 67.200 3.000 69.000 9.600 ;
        RECT 70.200 3.600 72.000 9.600 ;
        RECT 73.200 3.000 75.000 9.600 ;
        RECT 76.500 3.600 78.300 9.600 ;
        RECT 79.500 3.000 81.300 9.600 ;
        RECT 89.100 3.600 90.900 15.600 ;
        RECT 92.100 3.000 93.900 13.800 ;
        RECT 95.700 9.600 96.900 16.500 ;
        RECT 95.100 3.600 96.900 9.600 ;
        RECT 104.100 15.900 111.900 16.800 ;
        RECT 104.100 10.800 105.000 15.900 ;
        RECT 112.800 15.000 113.700 22.950 ;
        RECT 115.800 21.150 117.600 22.950 ;
        RECT 104.100 4.800 105.900 10.800 ;
        RECT 107.100 3.000 108.900 15.000 ;
        RECT 111.600 14.100 113.700 15.000 ;
        RECT 111.600 3.600 113.400 14.100 ;
        RECT 116.100 3.000 117.900 15.600 ;
        RECT 122.700 9.600 123.900 22.950 ;
        RECT 125.100 21.150 126.900 22.950 ;
        RECT 128.100 15.600 129.300 22.950 ;
        RECT 131.100 18.300 132.000 29.700 ;
        RECT 146.100 25.050 147.300 35.400 ;
        RECT 158.400 25.050 159.300 35.400 ;
        RECT 167.100 30.600 168.900 38.400 ;
        RECT 171.600 32.400 173.400 39.000 ;
        RECT 174.600 34.200 176.400 38.400 ;
        RECT 182.100 35.400 183.900 38.400 ;
        RECT 174.600 32.400 177.300 34.200 ;
        RECT 173.700 30.600 175.500 31.500 ;
        RECT 167.100 29.700 175.500 30.600 ;
        RECT 167.250 25.050 169.050 26.850 ;
        RECT 133.500 22.950 135.600 25.050 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 145.950 22.950 148.050 25.050 ;
        RECT 154.950 22.950 157.050 25.050 ;
        RECT 157.950 22.950 160.050 25.050 ;
        RECT 160.950 22.950 163.050 25.050 ;
        RECT 167.100 22.950 169.200 25.050 ;
        RECT 133.800 21.150 135.600 22.950 ;
        RECT 143.100 21.150 144.900 22.950 ;
        RECT 130.200 17.400 132.000 18.300 ;
        RECT 130.200 16.500 135.900 17.400 ;
        RECT 122.100 3.600 123.900 9.600 ;
        RECT 125.100 3.000 126.900 9.600 ;
        RECT 128.100 3.600 129.900 15.600 ;
        RECT 131.100 3.000 132.900 13.800 ;
        RECT 134.700 9.600 135.900 16.500 ;
        RECT 146.100 9.600 147.300 22.950 ;
        RECT 155.250 21.150 157.050 22.950 ;
        RECT 158.400 15.600 159.300 22.950 ;
        RECT 161.100 21.150 162.900 22.950 ;
        RECT 134.100 3.600 135.900 9.600 ;
        RECT 143.100 3.000 144.900 9.600 ;
        RECT 146.100 3.600 147.900 9.600 ;
        RECT 155.100 3.000 156.900 15.600 ;
        RECT 158.400 14.400 162.000 15.600 ;
        RECT 160.200 3.600 162.000 14.400 ;
        RECT 170.100 9.600 171.000 29.700 ;
        RECT 176.400 25.050 177.300 32.400 ;
        RECT 182.100 31.500 183.300 35.400 ;
        RECT 185.100 32.400 186.900 39.000 ;
        RECT 188.100 32.400 189.900 38.400 ;
        RECT 182.100 30.600 187.800 31.500 ;
        RECT 186.000 29.700 187.800 30.600 ;
        RECT 172.500 22.950 174.600 25.050 ;
        RECT 175.800 22.950 177.900 25.050 ;
        RECT 182.400 22.950 184.500 25.050 ;
        RECT 172.200 21.150 174.000 22.950 ;
        RECT 176.400 15.600 177.300 22.950 ;
        RECT 182.400 21.150 184.200 22.950 ;
        RECT 186.000 18.300 186.900 29.700 ;
        RECT 188.700 25.050 189.900 32.400 ;
        RECT 194.100 33.300 195.900 38.400 ;
        RECT 197.100 34.200 198.900 39.000 ;
        RECT 200.100 33.300 201.900 38.400 ;
        RECT 194.100 31.950 201.900 33.300 ;
        RECT 203.100 32.400 204.900 38.400 ;
        RECT 212.100 35.400 213.900 38.400 ;
        RECT 215.100 35.400 216.900 39.000 ;
        RECT 203.100 30.300 204.300 32.400 ;
        RECT 200.700 29.400 204.300 30.300 ;
        RECT 197.100 25.050 198.900 26.850 ;
        RECT 200.700 25.050 201.900 29.400 ;
        RECT 203.100 25.050 204.900 26.850 ;
        RECT 212.700 25.050 213.900 35.400 ;
        RECT 221.100 29.400 222.900 39.000 ;
        RECT 227.700 30.000 229.500 38.400 ;
        RECT 238.500 30.000 240.300 38.400 ;
        RECT 227.700 28.800 231.000 30.000 ;
        RECT 221.100 25.050 222.900 26.850 ;
        RECT 227.100 25.050 228.900 26.850 ;
        RECT 230.100 25.050 231.000 28.800 ;
        RECT 237.000 28.800 240.300 30.000 ;
        RECT 245.100 29.400 246.900 39.000 ;
        RECT 254.100 35.400 255.900 38.400 ;
        RECT 257.100 35.400 258.900 39.000 ;
        RECT 237.000 25.050 237.900 28.800 ;
        RECT 239.100 25.050 240.900 26.850 ;
        RECT 245.100 25.050 246.900 26.850 ;
        RECT 254.700 25.050 255.900 35.400 ;
        RECT 260.700 32.400 262.500 38.400 ;
        RECT 266.100 32.400 267.900 39.000 ;
        RECT 271.500 32.400 273.300 38.400 ;
        RECT 275.700 35.400 277.500 38.400 ;
        RECT 278.700 35.400 280.500 38.400 ;
        RECT 281.700 35.400 283.500 38.400 ;
        RECT 284.700 35.400 286.500 39.000 ;
        RECT 275.700 33.300 277.800 35.400 ;
        RECT 278.700 33.300 280.800 35.400 ;
        RECT 281.700 33.300 283.800 35.400 ;
        RECT 289.200 34.500 291.000 38.400 ;
        RECT 292.200 35.400 294.000 39.000 ;
        RECT 295.200 35.400 297.000 38.400 ;
        RECT 298.200 35.400 300.000 38.400 ;
        RECT 301.200 35.400 303.000 38.400 ;
        RECT 304.200 35.400 306.000 38.400 ;
        RECT 285.600 33.600 287.400 34.500 ;
        RECT 284.700 32.400 287.400 33.600 ;
        RECT 289.200 32.400 291.900 34.500 ;
        RECT 295.200 33.300 297.300 35.400 ;
        RECT 298.200 33.300 300.300 35.400 ;
        RECT 301.200 33.300 303.300 35.400 ;
        RECT 304.200 33.300 306.300 35.400 ;
        RECT 308.400 33.600 310.200 38.400 ;
        RECT 308.400 32.400 312.600 33.600 ;
        RECT 313.500 32.400 315.300 39.000 ;
        RECT 318.900 32.400 320.700 38.400 ;
        RECT 260.700 28.800 261.900 32.400 ;
        RECT 271.800 31.500 273.300 32.400 ;
        RECT 280.800 31.800 282.600 32.400 ;
        RECT 284.700 31.800 285.600 32.400 ;
        RECT 264.900 30.300 273.300 31.500 ;
        RECT 278.400 30.600 285.600 31.800 ;
        RECT 300.300 30.600 306.900 32.400 ;
        RECT 264.900 29.700 266.700 30.300 ;
        RECT 275.400 28.800 277.500 29.700 ;
        RECT 260.700 27.600 277.500 28.800 ;
        RECT 278.400 27.600 279.300 30.600 ;
        RECT 283.800 27.900 285.600 28.800 ;
        RECT 293.100 28.500 294.900 30.300 ;
        RECT 311.100 29.100 312.600 32.400 ;
        RECT 286.800 27.900 288.900 28.050 ;
        RECT 187.800 22.950 189.900 25.050 ;
        RECT 193.950 22.950 196.050 25.050 ;
        RECT 196.950 22.950 199.050 25.050 ;
        RECT 199.950 22.950 202.050 25.050 ;
        RECT 202.950 22.950 205.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 220.950 22.950 223.050 25.050 ;
        RECT 223.950 22.950 226.050 25.050 ;
        RECT 226.950 22.950 229.050 25.050 ;
        RECT 229.950 22.950 232.050 25.050 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 238.950 22.950 241.050 25.050 ;
        RECT 241.950 22.950 244.050 25.050 ;
        RECT 244.950 22.950 247.050 25.050 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 186.000 17.400 187.800 18.300 ;
        RECT 182.100 16.500 187.800 17.400 ;
        RECT 167.100 3.000 168.900 9.600 ;
        RECT 170.100 3.600 171.900 9.600 ;
        RECT 173.100 3.000 174.900 15.000 ;
        RECT 176.100 3.600 177.900 15.600 ;
        RECT 182.100 9.600 183.300 16.500 ;
        RECT 188.700 15.600 189.900 22.950 ;
        RECT 194.100 21.150 195.900 22.950 ;
        RECT 200.700 15.600 201.900 22.950 ;
        RECT 182.100 3.600 183.900 9.600 ;
        RECT 185.100 3.000 186.900 13.800 ;
        RECT 188.100 3.600 189.900 15.600 ;
        RECT 194.400 3.000 196.200 15.600 ;
        RECT 199.500 14.100 201.900 15.600 ;
        RECT 199.500 3.600 201.300 14.100 ;
        RECT 202.200 11.100 204.000 12.900 ;
        RECT 212.700 9.600 213.900 22.950 ;
        RECT 215.100 21.150 216.900 22.950 ;
        RECT 224.100 21.150 225.900 22.950 ;
        RECT 230.100 10.800 231.000 22.950 ;
        RECT 224.400 9.900 231.000 10.800 ;
        RECT 224.400 9.600 225.900 9.900 ;
        RECT 202.500 3.000 204.300 9.600 ;
        RECT 212.100 3.600 213.900 9.600 ;
        RECT 215.100 3.000 216.900 9.600 ;
        RECT 221.100 3.000 222.900 9.600 ;
        RECT 224.100 3.600 225.900 9.600 ;
        RECT 230.100 9.600 231.000 9.900 ;
        RECT 237.000 10.800 237.900 22.950 ;
        RECT 242.100 21.150 243.900 22.950 ;
        RECT 237.000 9.900 243.600 10.800 ;
        RECT 237.000 9.600 237.900 9.900 ;
        RECT 227.100 3.000 228.900 9.000 ;
        RECT 230.100 3.600 231.900 9.600 ;
        RECT 236.100 3.600 237.900 9.600 ;
        RECT 242.100 9.600 243.600 9.900 ;
        RECT 254.700 9.600 255.900 22.950 ;
        RECT 257.100 21.150 258.900 22.950 ;
        RECT 260.700 11.400 261.900 27.600 ;
        RECT 278.400 25.800 280.200 27.600 ;
        RECT 283.800 27.000 288.900 27.900 ;
        RECT 286.800 25.950 288.900 27.000 ;
        RECT 293.100 27.900 295.200 28.500 ;
        RECT 293.100 26.400 310.200 27.900 ;
        RECT 311.100 27.300 318.900 29.100 ;
        RECT 308.700 24.900 315.300 26.400 ;
        RECT 263.100 23.700 307.500 24.900 ;
        RECT 263.100 22.050 264.900 23.700 ;
        RECT 262.800 19.950 264.900 22.050 ;
        RECT 268.800 21.750 270.900 22.050 ;
        RECT 281.400 21.900 283.200 22.500 ;
        RECT 290.400 21.900 303.900 22.800 ;
        RECT 268.800 19.950 272.700 21.750 ;
        RECT 281.400 20.700 292.500 21.900 ;
        RECT 270.900 19.200 272.700 19.950 ;
        RECT 290.400 19.800 292.500 20.700 ;
        RECT 294.000 19.200 297.900 21.000 ;
        RECT 303.000 20.700 303.900 21.900 ;
        RECT 270.900 18.300 284.400 19.200 ;
        RECT 295.800 18.900 297.900 19.200 ;
        RECT 302.100 18.900 303.900 20.700 ;
        RECT 306.600 22.200 307.500 23.700 ;
        RECT 306.600 20.400 311.700 22.200 ;
        RECT 313.800 22.050 315.300 24.900 ;
        RECT 313.800 19.950 315.900 22.050 ;
        RECT 283.200 17.700 284.400 18.300 ;
        RECT 317.100 17.700 318.900 18.300 ;
        RECT 278.400 16.500 280.500 16.800 ;
        RECT 283.200 16.500 318.900 17.700 ;
        RECT 268.500 15.300 280.500 16.500 ;
        RECT 319.800 15.600 320.700 32.400 ;
        RECT 268.500 14.700 270.300 15.300 ;
        RECT 278.400 14.700 280.500 15.300 ;
        RECT 283.200 14.400 300.900 15.600 ;
        RECT 265.200 13.800 267.000 14.100 ;
        RECT 283.200 13.800 284.400 14.400 ;
        RECT 265.200 12.600 284.400 13.800 ;
        RECT 298.800 13.500 300.900 14.400 ;
        RECT 304.200 14.700 320.700 15.600 ;
        RECT 304.200 13.500 306.300 14.700 ;
        RECT 265.200 12.300 267.000 12.600 ;
        RECT 260.700 10.500 264.300 11.400 ;
        RECT 263.400 9.600 264.300 10.500 ;
        RECT 239.100 3.000 240.900 9.000 ;
        RECT 242.100 3.600 243.900 9.600 ;
        RECT 245.100 3.000 246.900 9.600 ;
        RECT 254.100 3.600 255.900 9.600 ;
        RECT 257.100 3.000 258.900 9.600 ;
        RECT 260.700 3.000 262.500 9.600 ;
        RECT 263.400 8.700 265.500 9.600 ;
        RECT 263.700 3.600 265.500 8.700 ;
        RECT 266.700 3.000 268.500 9.600 ;
        RECT 269.700 3.600 271.500 12.600 ;
        RECT 281.700 9.600 283.800 11.700 ;
        RECT 289.200 11.100 292.500 13.200 ;
        RECT 272.700 3.000 274.500 9.600 ;
        RECT 276.300 6.600 278.400 8.700 ;
        RECT 279.300 6.600 281.400 8.700 ;
        RECT 276.300 3.600 278.100 6.600 ;
        RECT 279.300 3.600 281.100 6.600 ;
        RECT 282.300 3.600 284.100 9.600 ;
        RECT 285.300 3.000 287.100 9.600 ;
        RECT 289.200 3.600 291.000 11.100 ;
        RECT 295.200 9.600 297.900 13.500 ;
        RECT 310.200 12.600 315.900 13.800 ;
        RECT 307.500 11.700 309.300 12.300 ;
        RECT 301.200 10.500 309.300 11.700 ;
        RECT 301.200 9.600 303.300 10.500 ;
        RECT 310.200 9.600 311.400 12.600 ;
        RECT 314.100 12.000 315.900 12.600 ;
        RECT 319.800 11.400 320.700 14.700 ;
        RECT 316.800 10.500 320.700 11.400 ;
        RECT 322.500 35.400 324.300 38.400 ;
        RECT 325.500 35.400 327.300 39.000 ;
        RECT 335.100 35.400 336.900 38.400 ;
        RECT 322.500 22.050 324.000 35.400 ;
        RECT 335.100 31.500 336.300 35.400 ;
        RECT 338.100 32.400 339.900 39.000 ;
        RECT 341.100 32.400 342.900 38.400 ;
        RECT 335.100 30.600 340.800 31.500 ;
        RECT 339.000 29.700 340.800 30.600 ;
        RECT 335.400 22.950 337.500 25.050 ;
        RECT 322.500 19.950 324.900 22.050 ;
        RECT 335.400 21.150 337.200 22.950 ;
        RECT 316.800 9.600 318.000 10.500 ;
        RECT 322.500 9.600 324.000 19.950 ;
        RECT 339.000 18.300 339.900 29.700 ;
        RECT 341.700 25.050 342.900 32.400 ;
        RECT 347.100 35.400 348.900 38.400 ;
        RECT 347.100 31.500 348.300 35.400 ;
        RECT 350.100 32.400 351.900 39.000 ;
        RECT 353.100 32.400 354.900 38.400 ;
        RECT 347.100 30.600 352.800 31.500 ;
        RECT 351.000 29.700 352.800 30.600 ;
        RECT 340.800 22.950 342.900 25.050 ;
        RECT 339.000 17.400 340.800 18.300 ;
        RECT 335.100 16.500 340.800 17.400 ;
        RECT 335.100 9.600 336.300 16.500 ;
        RECT 341.700 15.600 342.900 22.950 ;
        RECT 347.400 22.950 349.500 25.050 ;
        RECT 347.400 21.150 349.200 22.950 ;
        RECT 351.000 18.300 351.900 29.700 ;
        RECT 353.700 25.050 354.900 32.400 ;
        RECT 352.800 22.950 354.900 25.050 ;
        RECT 351.000 17.400 352.800 18.300 ;
        RECT 292.200 3.000 294.000 9.600 ;
        RECT 295.200 3.600 297.000 9.600 ;
        RECT 298.200 6.600 300.300 8.700 ;
        RECT 301.200 6.600 303.300 8.700 ;
        RECT 304.200 6.600 306.300 8.700 ;
        RECT 298.200 3.600 300.000 6.600 ;
        RECT 301.200 3.600 303.000 6.600 ;
        RECT 304.200 3.600 306.000 6.600 ;
        RECT 307.200 3.000 309.000 9.600 ;
        RECT 310.200 3.600 312.000 9.600 ;
        RECT 313.200 3.000 315.000 9.600 ;
        RECT 316.200 3.600 318.000 9.600 ;
        RECT 319.200 3.000 321.000 9.600 ;
        RECT 322.500 3.600 324.300 9.600 ;
        RECT 325.500 3.000 327.300 9.600 ;
        RECT 335.100 3.600 336.900 9.600 ;
        RECT 338.100 3.000 339.900 13.800 ;
        RECT 341.100 3.600 342.900 15.600 ;
        RECT 347.100 16.500 352.800 17.400 ;
        RECT 347.100 9.600 348.300 16.500 ;
        RECT 353.700 15.600 354.900 22.950 ;
        RECT 347.100 3.600 348.900 9.600 ;
        RECT 350.100 3.000 351.900 13.800 ;
        RECT 353.100 3.600 354.900 15.600 ;
      LAYER metal2 ;
        RECT 139.950 352.950 142.050 355.050 ;
        RECT 160.950 352.950 163.050 355.050 ;
        RECT 166.950 352.950 169.050 355.050 ;
        RECT 190.950 352.950 193.050 355.050 ;
        RECT 17.700 345.300 19.800 347.400 ;
        RECT 20.700 345.300 22.800 347.400 ;
        RECT 23.700 345.300 25.800 347.400 ;
        RECT 18.300 341.700 19.500 345.300 ;
        RECT 17.400 339.600 19.500 341.700 ;
        RECT 4.800 331.950 6.900 334.050 ;
        RECT 10.800 331.950 12.900 334.050 ;
        RECT 17.400 320.700 18.900 339.600 ;
        RECT 21.300 328.800 22.500 345.300 ;
        RECT 20.400 326.700 22.500 328.800 ;
        RECT 21.300 320.700 22.500 326.700 ;
        RECT 23.700 323.700 24.900 345.300 ;
        RECT 31.800 344.400 33.900 346.500 ;
        RECT 37.200 345.300 39.300 347.400 ;
        RECT 40.200 345.300 42.300 347.400 ;
        RECT 43.200 345.300 45.300 347.400 ;
        RECT 28.800 337.950 30.900 340.050 ;
        RECT 29.400 335.400 30.600 337.650 ;
        RECT 29.400 328.050 30.450 335.400 ;
        RECT 32.400 333.900 33.300 344.400 ;
        RECT 35.100 338.400 37.200 340.500 ;
        RECT 32.400 331.800 34.500 333.900 ;
        RECT 38.100 333.000 39.300 345.300 ;
        RECT 28.950 325.950 31.050 328.050 ;
        RECT 32.400 325.200 33.300 331.800 ;
        RECT 37.800 330.900 39.900 333.000 ;
        RECT 23.700 321.600 25.800 323.700 ;
        RECT 32.400 323.100 34.500 325.200 ;
        RECT 38.100 323.700 39.300 330.900 ;
        RECT 40.800 327.600 42.300 345.300 ;
        RECT 40.800 325.500 42.900 327.600 ;
        RECT 37.800 321.600 39.900 323.700 ;
        RECT 40.800 320.700 42.300 325.500 ;
        RECT 44.100 323.700 45.300 345.300 ;
        RECT 17.400 318.600 20.400 320.700 ;
        RECT 21.300 318.600 23.400 320.700 ;
        RECT 40.200 318.600 42.300 320.700 ;
        RECT 43.200 318.600 45.300 323.700 ;
        RECT 46.200 345.300 48.300 347.400 ;
        RECT 86.700 345.300 88.800 347.400 ;
        RECT 89.700 345.300 91.800 347.400 ;
        RECT 92.700 345.300 94.800 347.400 ;
        RECT 46.200 327.600 47.700 345.300 ;
        RECT 87.300 341.700 88.500 345.300 ;
        RECT 86.400 339.600 88.500 341.700 ;
        RECT 65.400 336.450 66.600 336.600 ;
        RECT 65.400 335.400 69.450 336.450 ;
        RECT 65.400 334.350 66.600 335.400 ;
        RECT 55.800 331.950 57.900 334.050 ;
        RECT 64.800 331.950 66.900 334.050 ;
        RECT 46.200 325.500 48.300 327.600 ;
        RECT 52.950 325.950 55.050 328.050 ;
        RECT 46.200 320.700 47.700 325.500 ;
        RECT 46.200 318.600 48.300 320.700 ;
        RECT 17.400 306.300 20.400 308.400 ;
        RECT 21.300 306.300 23.400 308.400 ;
        RECT 40.200 306.300 42.300 308.400 ;
        RECT 4.800 292.950 6.900 295.050 ;
        RECT 10.800 292.950 12.900 295.050 ;
        RECT 17.400 287.400 18.900 306.300 ;
        RECT 21.300 300.300 22.500 306.300 ;
        RECT 20.400 298.200 22.500 300.300 ;
        RECT 17.400 285.300 19.500 287.400 ;
        RECT 18.300 281.700 19.500 285.300 ;
        RECT 21.300 281.700 22.500 298.200 ;
        RECT 23.700 303.300 25.800 305.400 ;
        RECT 23.700 281.700 24.900 303.300 ;
        RECT 32.400 301.800 34.500 303.900 ;
        RECT 37.800 303.300 39.900 305.400 ;
        RECT 28.950 298.950 31.050 301.050 ;
        RECT 29.400 291.600 30.450 298.950 ;
        RECT 32.400 295.200 33.300 301.800 ;
        RECT 38.100 296.100 39.300 303.300 ;
        RECT 40.800 301.500 42.300 306.300 ;
        RECT 43.200 303.300 45.300 308.400 ;
        RECT 40.800 299.400 42.900 301.500 ;
        RECT 32.400 293.100 34.500 295.200 ;
        RECT 37.800 294.000 39.900 296.100 ;
        RECT 29.400 289.350 30.600 291.600 ;
        RECT 28.800 286.950 30.900 289.050 ;
        RECT 32.400 282.600 33.300 293.100 ;
        RECT 35.100 286.500 37.200 288.600 ;
        RECT 17.700 279.600 19.800 281.700 ;
        RECT 20.700 279.600 22.800 281.700 ;
        RECT 23.700 279.600 25.800 281.700 ;
        RECT 31.800 280.500 33.900 282.600 ;
        RECT 38.100 281.700 39.300 294.000 ;
        RECT 40.800 281.700 42.300 299.400 ;
        RECT 44.100 281.700 45.300 303.300 ;
        RECT 37.200 279.600 39.300 281.700 ;
        RECT 40.200 279.600 42.300 281.700 ;
        RECT 43.200 279.600 45.300 281.700 ;
        RECT 46.200 306.300 48.300 308.400 ;
        RECT 46.200 301.500 47.700 306.300 ;
        RECT 46.200 299.400 48.300 301.500 ;
        RECT 46.200 281.700 47.700 299.400 ;
        RECT 53.400 298.050 54.450 325.950 ;
        RECT 68.400 325.050 69.450 335.400 ;
        RECT 73.800 331.950 75.900 334.050 ;
        RECT 79.800 331.950 81.900 334.050 ;
        RECT 58.950 322.950 61.050 325.050 ;
        RECT 67.950 322.950 70.050 325.050 ;
        RECT 52.950 295.950 55.050 298.050 ;
        RECT 55.800 292.950 57.900 295.050 ;
        RECT 46.200 279.600 48.300 281.700 ;
        RECT 59.400 274.050 60.450 322.950 ;
        RECT 86.400 320.700 87.900 339.600 ;
        RECT 90.300 328.800 91.500 345.300 ;
        RECT 89.400 326.700 91.500 328.800 ;
        RECT 90.300 320.700 91.500 326.700 ;
        RECT 92.700 323.700 93.900 345.300 ;
        RECT 100.800 344.400 102.900 346.500 ;
        RECT 106.200 345.300 108.300 347.400 ;
        RECT 109.200 345.300 111.300 347.400 ;
        RECT 112.200 345.300 114.300 347.400 ;
        RECT 97.800 337.950 99.900 340.050 ;
        RECT 98.400 335.400 99.600 337.650 ;
        RECT 92.700 321.600 94.800 323.700 ;
        RECT 98.400 322.050 99.450 335.400 ;
        RECT 101.400 333.900 102.300 344.400 ;
        RECT 104.100 338.400 106.200 340.500 ;
        RECT 101.400 331.800 103.500 333.900 ;
        RECT 107.100 333.000 108.300 345.300 ;
        RECT 101.400 325.200 102.300 331.800 ;
        RECT 106.800 330.900 108.900 333.000 ;
        RECT 101.400 323.100 103.500 325.200 ;
        RECT 107.100 323.700 108.300 330.900 ;
        RECT 109.800 327.600 111.300 345.300 ;
        RECT 109.800 325.500 111.900 327.600 ;
        RECT 86.400 318.600 89.400 320.700 ;
        RECT 90.300 318.600 92.400 320.700 ;
        RECT 97.950 319.950 100.050 322.050 ;
        RECT 106.800 321.600 108.900 323.700 ;
        RECT 109.800 320.700 111.300 325.500 ;
        RECT 113.100 323.700 114.300 345.300 ;
        RECT 109.200 318.600 111.300 320.700 ;
        RECT 112.200 318.600 114.300 323.700 ;
        RECT 115.200 345.300 117.300 347.400 ;
        RECT 115.200 327.600 116.700 345.300 ;
        RECT 133.950 343.950 136.050 346.050 ;
        RECT 118.950 334.950 121.050 337.050 ;
        RECT 134.400 336.600 135.450 343.950 ;
        RECT 115.200 325.500 117.300 327.600 ;
        RECT 115.200 320.700 116.700 325.500 ;
        RECT 115.200 318.600 117.300 320.700 ;
        RECT 94.950 307.950 97.050 310.050 ;
        RECT 115.950 307.950 118.050 310.050 ;
        RECT 70.950 304.950 73.050 307.050 ;
        RECT 91.950 304.950 94.050 307.050 ;
        RECT 67.950 298.950 70.050 301.050 ;
        RECT 64.800 292.950 66.900 295.050 ;
        RECT 65.400 291.900 66.600 292.650 ;
        RECT 64.950 289.800 67.050 291.900 ;
        RECT 68.400 283.050 69.450 298.950 ;
        RECT 71.400 291.900 72.450 304.950 ;
        RECT 79.950 298.950 82.050 301.050 ;
        RECT 80.400 294.600 81.450 298.950 ;
        RECT 80.400 292.350 81.600 294.600 ;
        RECT 85.950 294.000 88.050 298.050 ;
        RECT 92.400 294.600 93.450 304.950 ;
        RECT 95.400 301.050 96.450 307.950 ;
        RECT 112.950 301.950 115.050 304.050 ;
        RECT 94.950 298.950 97.050 301.050 ;
        RECT 86.400 292.350 87.600 294.000 ;
        RECT 92.400 292.350 93.600 294.600 ;
        RECT 97.950 293.100 100.050 295.200 ;
        RECT 113.400 294.600 114.450 301.950 ;
        RECT 116.400 295.050 117.450 307.950 ;
        RECT 119.400 307.050 120.450 334.950 ;
        RECT 134.400 334.350 135.600 336.600 ;
        RECT 124.800 331.950 126.900 334.050 ;
        RECT 133.800 331.950 135.900 334.050 ;
        RECT 133.950 316.950 136.050 319.050 ;
        RECT 118.950 304.950 121.050 307.050 ;
        RECT 134.400 304.050 135.450 316.950 ;
        RECT 140.400 313.050 141.450 352.950 ;
        RECT 154.950 343.950 157.050 346.050 ;
        RECT 145.950 338.100 148.050 340.200 ;
        RECT 146.400 337.350 147.600 338.100 ;
        RECT 146.400 334.950 148.500 337.050 ;
        RECT 151.800 334.950 153.900 337.050 ;
        RECT 155.400 321.450 156.450 343.950 ;
        RECT 161.400 339.600 162.450 352.950 ;
        RECT 167.400 346.050 168.450 352.950 ;
        RECT 166.950 343.950 169.050 346.050 ;
        RECT 167.400 339.600 168.450 343.950 ;
        RECT 191.400 339.600 192.450 352.950 ;
        RECT 253.950 346.950 256.050 349.050 ;
        RECT 277.950 346.950 280.050 349.050 ;
        RECT 161.400 337.350 162.600 339.600 ;
        RECT 167.400 337.350 168.600 339.600 ;
        RECT 182.400 339.450 183.600 339.600 ;
        RECT 182.400 338.400 186.450 339.450 ;
        RECT 182.400 337.350 183.600 338.400 ;
        RECT 160.950 334.950 163.050 337.050 ;
        RECT 163.950 334.950 166.050 337.050 ;
        RECT 166.950 334.950 169.050 337.050 ;
        RECT 169.950 334.950 172.050 337.050 ;
        RECT 176.100 334.950 178.200 337.050 ;
        RECT 181.500 334.950 183.600 337.050 ;
        RECT 164.400 333.900 165.600 334.650 ;
        RECT 163.950 331.800 166.050 333.900 ;
        RECT 170.400 333.000 171.600 334.650 ;
        RECT 169.950 328.950 172.050 333.000 ;
        RECT 185.400 331.050 186.450 338.400 ;
        RECT 191.400 337.350 192.600 339.600 ;
        RECT 199.950 337.950 202.050 340.050 ;
        RECT 208.950 338.100 211.050 340.200 ;
        RECT 214.950 338.100 217.050 340.200 ;
        RECT 220.950 339.000 223.050 342.900 ;
        RECT 191.400 334.950 193.500 337.050 ;
        RECT 196.800 334.950 198.900 337.050 ;
        RECT 184.950 328.950 187.050 331.050 ;
        RECT 190.950 328.950 193.050 331.050 ;
        RECT 170.400 325.050 171.450 328.950 ;
        RECT 169.950 322.950 172.050 325.050 ;
        RECT 155.400 320.400 159.450 321.450 ;
        RECT 139.950 310.950 142.050 313.050 ;
        RECT 154.950 310.950 157.050 313.050 ;
        RECT 133.950 301.950 136.050 304.050 ;
        RECT 136.950 298.950 139.050 301.050 ;
        RECT 98.400 292.350 99.600 293.100 ;
        RECT 113.400 292.350 114.600 294.600 ;
        RECT 115.950 292.950 118.050 295.050 ;
        RECT 121.950 293.100 124.050 295.200 ;
        RECT 130.950 293.100 133.050 295.200 ;
        RECT 137.400 294.600 138.450 298.950 ;
        RECT 122.400 292.350 123.600 293.100 ;
        RECT 131.400 292.350 132.600 293.100 ;
        RECT 137.400 292.350 138.600 294.600 ;
        RECT 148.950 293.100 151.050 295.200 ;
        RECT 155.400 294.600 156.450 310.950 ;
        RECT 158.400 295.050 159.450 320.400 ;
        RECT 169.950 319.800 172.050 321.900 ;
        RECT 163.950 307.950 166.050 310.050 ;
        RECT 164.400 298.050 165.450 307.950 ;
        RECT 163.950 295.950 166.050 298.050 ;
        RECT 149.400 292.350 150.600 293.100 ;
        RECT 155.400 292.350 156.600 294.600 ;
        RECT 157.950 292.950 160.050 295.050 ;
        RECT 164.400 294.600 165.450 295.950 ;
        RECT 170.400 295.050 171.450 319.800 ;
        RECT 185.400 298.050 186.450 328.950 ;
        RECT 191.400 313.050 192.450 328.950 ;
        RECT 200.400 319.050 201.450 337.950 ;
        RECT 209.400 337.350 210.600 338.100 ;
        RECT 215.400 337.350 216.600 338.100 ;
        RECT 221.400 337.350 222.600 339.000 ;
        RECT 226.950 338.100 229.050 340.200 ;
        RECT 238.950 338.100 241.050 340.200 ;
        RECT 247.950 338.100 250.050 340.200 ;
        RECT 254.400 339.600 255.450 346.950 ;
        RECT 227.400 337.350 228.600 338.100 ;
        RECT 239.400 337.350 240.600 338.100 ;
        RECT 248.400 337.350 249.600 338.100 ;
        RECT 254.400 337.350 255.600 339.600 ;
        RECT 262.950 338.100 265.050 340.200 ;
        RECT 263.400 337.350 264.600 338.100 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 211.950 334.950 214.050 337.050 ;
        RECT 214.950 334.950 217.050 337.050 ;
        RECT 220.950 334.950 223.050 337.050 ;
        RECT 223.950 334.950 226.050 337.050 ;
        RECT 226.950 334.950 229.050 337.050 ;
        RECT 233.100 334.950 235.200 337.050 ;
        RECT 238.500 334.950 240.600 337.050 ;
        RECT 241.800 334.950 243.900 337.050 ;
        RECT 247.950 334.950 250.050 337.050 ;
        RECT 250.950 334.950 253.050 337.050 ;
        RECT 253.950 334.950 256.050 337.050 ;
        RECT 256.950 334.950 259.050 337.050 ;
        RECT 263.400 334.950 265.500 337.050 ;
        RECT 268.800 334.950 270.900 337.050 ;
        RECT 278.400 336.900 279.450 346.950 ;
        RECT 287.700 345.300 289.800 347.400 ;
        RECT 290.700 345.300 292.800 347.400 ;
        RECT 293.700 345.300 295.800 347.400 ;
        RECT 288.300 341.700 289.500 345.300 ;
        RECT 287.400 339.600 289.500 341.700 ;
        RECT 277.950 334.800 280.050 336.900 ;
        RECT 206.400 332.400 207.600 334.650 ;
        RECT 212.400 333.900 213.600 334.650 ;
        RECT 199.950 316.950 202.050 319.050 ;
        RECT 193.950 313.950 196.050 316.050 ;
        RECT 190.950 310.950 193.050 313.050 ;
        RECT 187.950 298.950 190.050 301.050 ;
        RECT 184.950 295.950 187.050 298.050 ;
        RECT 164.400 292.350 165.600 294.600 ;
        RECT 169.950 292.950 172.050 295.050 ;
        RECT 175.950 293.100 178.050 295.200 ;
        RECT 181.950 293.100 184.050 295.200 ;
        RECT 188.400 294.600 189.450 298.950 ;
        RECT 194.400 295.050 195.450 313.950 ;
        RECT 206.400 310.050 207.450 332.400 ;
        RECT 211.950 328.950 214.050 333.900 ;
        RECT 224.400 332.400 225.600 334.650 ;
        RECT 212.400 322.050 213.450 328.950 ;
        RECT 211.950 319.950 214.050 322.050 ;
        RECT 214.950 313.950 217.050 316.050 ;
        RECT 205.950 307.950 208.050 310.050 ;
        RECT 208.950 298.950 211.050 301.050 ;
        RECT 176.400 292.350 177.600 293.100 ;
        RECT 182.400 292.350 183.600 293.100 ;
        RECT 188.400 292.350 189.600 294.600 ;
        RECT 193.950 292.950 196.050 295.050 ;
        RECT 199.950 294.000 202.050 298.050 ;
        RECT 200.400 292.350 201.600 294.000 ;
        RECT 205.800 293.100 207.900 295.200 ;
        RECT 209.400 295.050 210.450 298.950 ;
        RECT 206.400 292.350 207.600 293.100 ;
        RECT 208.950 292.950 211.050 295.050 ;
        RECT 215.400 294.600 216.450 313.950 ;
        RECT 224.400 304.050 225.450 332.400 ;
        RECT 229.950 331.950 232.050 334.050 ;
        RECT 233.400 332.400 234.600 334.650 ;
        RECT 242.400 333.900 243.600 334.650 ;
        RECT 230.400 318.450 231.450 331.950 ;
        RECT 233.400 322.050 234.450 332.400 ;
        RECT 241.950 331.800 244.050 333.900 ;
        RECT 251.400 332.400 252.600 334.650 ;
        RECT 257.400 332.400 258.600 334.650 ;
        RECT 241.950 325.950 244.050 328.050 ;
        RECT 232.950 319.950 235.050 322.050 ;
        RECT 230.400 317.400 234.450 318.450 ;
        RECT 217.950 301.950 220.050 304.050 ;
        RECT 223.950 301.950 226.050 304.050 ;
        RECT 229.950 301.950 232.050 304.050 ;
        RECT 218.400 298.050 219.450 301.950 ;
        RECT 217.950 295.950 220.050 298.050 ;
        RECT 230.400 295.200 231.450 301.950 ;
        RECT 233.400 298.050 234.450 317.400 ;
        RECT 235.950 304.950 238.050 307.050 ;
        RECT 232.950 295.950 235.050 298.050 ;
        RECT 215.400 292.350 216.600 294.600 ;
        RECT 229.950 293.100 232.050 295.200 ;
        RECT 236.400 294.600 237.450 304.950 ;
        RECT 242.400 294.600 243.450 325.950 ;
        RECT 251.400 319.050 252.450 332.400 ;
        RECT 257.400 328.050 258.450 332.400 ;
        RECT 274.800 331.950 276.900 334.050 ;
        RECT 280.800 331.950 282.900 334.050 ;
        RECT 262.950 328.950 265.050 331.050 ;
        RECT 256.950 325.950 259.050 328.050 ;
        RECT 250.950 316.950 253.050 319.050 ;
        RECT 263.400 316.050 264.450 328.950 ;
        RECT 287.400 320.700 288.900 339.600 ;
        RECT 291.300 328.800 292.500 345.300 ;
        RECT 290.400 326.700 292.500 328.800 ;
        RECT 291.300 320.700 292.500 326.700 ;
        RECT 293.700 323.700 294.900 345.300 ;
        RECT 301.800 344.400 303.900 346.500 ;
        RECT 307.200 345.300 309.300 347.400 ;
        RECT 310.200 345.300 312.300 347.400 ;
        RECT 313.200 345.300 315.300 347.400 ;
        RECT 298.800 337.950 300.900 340.050 ;
        RECT 299.400 336.900 300.600 337.650 ;
        RECT 298.950 334.800 301.050 336.900 ;
        RECT 302.400 333.900 303.300 344.400 ;
        RECT 305.100 338.400 307.200 340.500 ;
        RECT 302.400 331.800 304.500 333.900 ;
        RECT 308.100 333.000 309.300 345.300 ;
        RECT 302.400 325.200 303.300 331.800 ;
        RECT 307.800 330.900 309.900 333.000 ;
        RECT 293.700 321.600 295.800 323.700 ;
        RECT 302.400 323.100 304.500 325.200 ;
        RECT 308.100 323.700 309.300 330.900 ;
        RECT 310.800 327.600 312.300 345.300 ;
        RECT 310.800 325.500 312.900 327.600 ;
        RECT 307.800 321.600 309.900 323.700 ;
        RECT 310.800 320.700 312.300 325.500 ;
        RECT 314.100 323.700 315.300 345.300 ;
        RECT 287.400 318.600 290.400 320.700 ;
        RECT 291.300 318.600 293.400 320.700 ;
        RECT 310.200 318.600 312.300 320.700 ;
        RECT 313.200 318.600 315.300 323.700 ;
        RECT 316.200 345.300 318.300 347.400 ;
        RECT 316.200 327.600 317.700 345.300 ;
        RECT 349.950 338.100 352.050 340.200 ;
        RECT 350.400 337.350 351.600 338.100 ;
        RECT 335.400 336.450 336.600 336.600 ;
        RECT 335.400 335.400 339.450 336.450 ;
        RECT 335.400 334.350 336.600 335.400 ;
        RECT 325.800 331.950 327.900 334.050 ;
        RECT 334.800 331.950 336.900 334.050 ;
        RECT 316.200 325.500 318.300 327.600 ;
        RECT 316.200 320.700 317.700 325.500 ;
        RECT 316.200 318.600 318.300 320.700 ;
        RECT 338.400 316.050 339.450 335.400 ;
        RECT 346.950 334.950 349.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 352.950 334.950 355.050 337.050 ;
        RECT 347.400 332.400 348.600 334.650 ;
        RECT 353.400 332.400 354.600 334.650 ;
        RECT 347.400 330.450 348.450 332.400 ;
        RECT 347.400 329.400 351.450 330.450 ;
        RECT 262.950 313.950 265.050 316.050 ;
        RECT 310.950 313.950 313.050 316.050 ;
        RECT 337.950 313.950 340.050 316.050 ;
        RECT 253.950 304.950 256.050 307.050 ;
        RECT 299.400 306.300 302.400 308.400 ;
        RECT 303.300 306.300 305.400 308.400 ;
        RECT 254.400 298.050 255.450 304.950 ;
        RECT 256.950 301.950 259.050 304.050 ;
        RECT 265.950 301.950 268.050 304.050 ;
        RECT 280.950 301.950 283.050 304.050 ;
        RECT 253.950 295.950 256.050 298.050 ;
        RECT 257.400 297.450 258.450 301.950 ;
        RECT 257.400 296.400 261.450 297.450 ;
        RECT 230.400 292.350 231.600 293.100 ;
        RECT 236.400 292.350 237.600 294.600 ;
        RECT 242.400 292.350 243.600 294.600 ;
        RECT 250.950 293.100 253.050 295.200 ;
        RECT 260.400 294.600 261.450 296.400 ;
        RECT 266.400 295.200 267.450 301.950 ;
        RECT 251.400 292.350 252.600 293.100 ;
        RECT 260.400 292.350 261.600 294.600 ;
        RECT 265.950 293.100 268.050 295.200 ;
        RECT 281.400 294.600 282.450 301.950 ;
        RECT 266.400 292.350 267.600 293.100 ;
        RECT 281.400 292.350 282.600 294.600 ;
        RECT 286.800 292.950 288.900 295.050 ;
        RECT 292.800 292.950 294.900 295.050 ;
        RECT 70.950 289.800 73.050 291.900 ;
        RECT 76.950 289.950 79.050 292.050 ;
        RECT 79.950 289.950 82.050 292.050 ;
        RECT 82.950 289.950 85.050 292.050 ;
        RECT 85.950 289.950 88.050 292.050 ;
        RECT 91.950 289.950 94.050 292.050 ;
        RECT 94.950 289.950 97.050 292.050 ;
        RECT 97.950 289.950 100.050 292.050 ;
        RECT 106.950 289.950 109.050 292.050 ;
        RECT 109.950 289.950 112.050 292.050 ;
        RECT 112.950 289.950 115.050 292.050 ;
        RECT 118.950 289.950 121.050 292.050 ;
        RECT 121.950 289.950 124.050 292.050 ;
        RECT 130.950 289.950 133.050 292.050 ;
        RECT 133.950 289.950 136.050 292.050 ;
        RECT 136.950 289.950 139.050 292.050 ;
        RECT 139.950 289.950 142.050 292.050 ;
        RECT 145.950 289.950 148.050 292.050 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 154.950 289.950 157.050 292.050 ;
        RECT 163.950 289.950 166.050 292.050 ;
        RECT 166.950 289.950 169.050 292.050 ;
        RECT 172.950 289.950 175.050 292.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 178.950 289.950 181.050 292.050 ;
        RECT 181.950 289.950 184.050 292.050 ;
        RECT 187.950 289.950 190.050 292.050 ;
        RECT 190.950 289.950 193.050 292.050 ;
        RECT 196.950 289.950 199.050 292.050 ;
        RECT 199.950 289.950 202.050 292.050 ;
        RECT 202.950 289.950 205.050 292.050 ;
        RECT 205.950 289.950 208.050 292.050 ;
        RECT 214.950 289.950 217.050 292.050 ;
        RECT 217.950 289.950 220.050 292.050 ;
        RECT 220.950 289.950 223.050 292.050 ;
        RECT 229.950 289.950 232.050 292.050 ;
        RECT 232.950 289.950 235.050 292.050 ;
        RECT 235.950 289.950 238.050 292.050 ;
        RECT 242.100 289.950 244.200 292.050 ;
        RECT 245.400 289.950 247.500 292.050 ;
        RECT 250.800 289.950 252.900 292.050 ;
        RECT 256.950 289.950 259.050 292.050 ;
        RECT 259.950 289.950 262.050 292.050 ;
        RECT 262.950 289.950 265.050 292.050 ;
        RECT 265.950 289.950 268.050 292.050 ;
        RECT 275.400 289.950 277.500 292.050 ;
        RECT 280.800 289.950 282.900 292.050 ;
        RECT 67.950 280.950 70.050 283.050 ;
        RECT 58.950 271.950 61.050 274.050 ;
        RECT 32.700 267.300 34.800 269.400 ;
        RECT 35.700 267.300 37.800 269.400 ;
        RECT 38.700 267.300 40.800 269.400 ;
        RECT 33.300 263.700 34.500 267.300 ;
        RECT 1.950 260.100 4.050 262.200 ;
        RECT 13.950 260.100 16.050 262.200 ;
        RECT 32.400 261.600 34.500 263.700 ;
        RECT 2.400 241.050 3.450 260.100 ;
        RECT 14.400 259.350 15.600 260.100 ;
        RECT 8.100 256.950 10.200 259.050 ;
        RECT 13.500 256.950 15.600 259.050 ;
        RECT 19.800 253.950 21.900 256.050 ;
        RECT 25.800 253.950 27.900 256.050 ;
        RECT 32.400 242.700 33.900 261.600 ;
        RECT 36.300 250.800 37.500 267.300 ;
        RECT 35.400 248.700 37.500 250.800 ;
        RECT 36.300 242.700 37.500 248.700 ;
        RECT 38.700 245.700 39.900 267.300 ;
        RECT 46.800 266.400 48.900 268.500 ;
        RECT 52.200 267.300 54.300 269.400 ;
        RECT 55.200 267.300 57.300 269.400 ;
        RECT 58.200 267.300 60.300 269.400 ;
        RECT 43.800 259.950 45.900 262.050 ;
        RECT 44.400 257.400 45.600 259.650 ;
        RECT 38.700 243.600 40.800 245.700 ;
        RECT 1.950 238.950 4.050 241.050 ;
        RECT 32.400 240.600 35.400 242.700 ;
        RECT 36.300 240.600 38.400 242.700 ;
        RECT 2.400 199.050 3.450 238.950 ;
        RECT 44.400 238.050 45.450 257.400 ;
        RECT 47.400 255.900 48.300 266.400 ;
        RECT 50.100 260.400 52.200 262.500 ;
        RECT 47.400 253.800 49.500 255.900 ;
        RECT 53.100 255.000 54.300 267.300 ;
        RECT 47.400 247.200 48.300 253.800 ;
        RECT 52.800 252.900 54.900 255.000 ;
        RECT 47.400 245.100 49.500 247.200 ;
        RECT 53.100 245.700 54.300 252.900 ;
        RECT 55.800 249.600 57.300 267.300 ;
        RECT 55.800 247.500 57.900 249.600 ;
        RECT 52.800 243.600 54.900 245.700 ;
        RECT 55.800 242.700 57.300 247.500 ;
        RECT 59.100 245.700 60.300 267.300 ;
        RECT 55.200 240.600 57.300 242.700 ;
        RECT 58.200 240.600 60.300 245.700 ;
        RECT 61.200 267.300 63.300 269.400 ;
        RECT 71.400 268.050 72.450 289.800 ;
        RECT 77.400 287.400 78.600 289.650 ;
        RECT 83.400 288.900 84.600 289.650 ;
        RECT 95.400 288.900 96.600 289.650 ;
        RECT 110.400 288.900 111.600 289.650 ;
        RECT 77.400 283.050 78.450 287.400 ;
        RECT 82.950 286.800 85.050 288.900 ;
        RECT 94.950 286.800 97.050 288.900 ;
        RECT 109.950 286.800 112.050 288.900 ;
        RECT 119.400 287.400 120.600 289.650 ;
        RECT 134.400 288.900 135.600 289.650 ;
        RECT 79.950 283.950 82.050 286.050 ;
        RECT 97.950 283.950 100.050 286.050 ;
        RECT 112.950 283.950 115.050 286.050 ;
        RECT 76.950 280.950 79.050 283.050 ;
        RECT 73.950 277.950 76.050 280.050 ;
        RECT 74.400 274.050 75.450 277.950 ;
        RECT 80.400 277.050 81.450 283.950 ;
        RECT 79.950 274.950 82.050 277.050 ;
        RECT 73.950 271.950 76.050 274.050 ;
        RECT 61.200 249.600 62.700 267.300 ;
        RECT 70.950 265.950 73.050 268.050 ;
        RECT 70.800 253.950 72.900 256.050 ;
        RECT 61.200 247.500 63.300 249.600 ;
        RECT 61.200 242.700 62.700 247.500 ;
        RECT 61.200 240.600 63.300 242.700 ;
        RECT 74.400 238.050 75.450 271.950 ;
        RECT 91.950 260.100 94.050 262.200 ;
        RECT 98.400 262.050 99.450 283.950 ;
        RECT 106.950 274.950 109.050 277.050 ;
        RECT 92.400 259.350 93.600 260.100 ;
        RECT 97.800 259.950 99.900 262.050 ;
        RECT 107.400 261.600 108.450 274.950 ;
        RECT 113.400 262.200 114.450 283.950 ;
        RECT 119.400 268.050 120.450 287.400 ;
        RECT 133.950 286.800 136.050 288.900 ;
        RECT 140.400 288.450 141.600 289.650 ;
        RECT 140.400 287.400 144.450 288.450 ;
        RECT 146.400 288.000 147.600 289.650 ;
        RECT 152.400 288.900 153.600 289.650 ;
        RECT 139.950 277.950 142.050 280.050 ;
        RECT 143.400 279.450 144.450 287.400 ;
        RECT 145.950 283.950 148.050 288.000 ;
        RECT 151.950 286.800 154.050 288.900 ;
        RECT 160.950 286.950 163.050 289.050 ;
        RECT 167.400 287.400 168.600 289.650 ;
        RECT 173.400 288.900 174.600 289.650 ;
        RECT 157.950 280.950 160.050 283.050 ;
        RECT 143.400 278.400 147.450 279.450 ;
        RECT 140.400 270.450 141.450 277.950 ;
        RECT 140.400 269.400 144.450 270.450 ;
        RECT 118.950 265.950 121.050 268.050 ;
        RECT 107.400 259.350 108.600 261.600 ;
        RECT 112.950 260.100 115.050 262.200 ;
        RECT 121.950 260.100 124.050 262.200 ;
        RECT 143.400 261.600 144.450 269.400 ;
        RECT 146.400 262.050 147.450 278.400 ;
        RECT 113.400 259.350 114.600 260.100 ;
        RECT 122.400 259.350 123.600 260.100 ;
        RECT 143.400 259.350 144.600 261.600 ;
        RECT 145.950 259.950 148.050 262.050 ;
        RECT 151.950 260.100 154.050 262.200 ;
        RECT 158.400 261.600 159.450 280.950 ;
        RECT 161.400 265.050 162.450 286.950 ;
        RECT 167.400 283.050 168.450 287.400 ;
        RECT 172.950 286.800 175.050 288.900 ;
        RECT 179.400 287.400 180.600 289.650 ;
        RECT 174.000 285.450 178.050 286.050 ;
        RECT 173.400 283.950 178.050 285.450 ;
        RECT 166.950 280.950 169.050 283.050 ;
        RECT 167.400 268.050 168.450 280.950 ;
        RECT 169.950 268.950 172.050 271.050 ;
        RECT 166.950 265.950 169.050 268.050 ;
        RECT 170.400 265.050 171.450 268.950 ;
        RECT 160.950 262.950 163.050 265.050 ;
        RECT 168.000 264.900 171.450 265.050 ;
        RECT 166.950 263.400 171.450 264.900 ;
        RECT 166.950 262.950 171.000 263.400 ;
        RECT 166.950 262.800 169.050 262.950 ;
        RECT 152.400 259.350 153.600 260.100 ;
        RECT 158.400 259.350 159.600 261.600 ;
        RECT 166.950 259.950 169.050 262.050 ;
        RECT 173.400 261.600 174.450 283.950 ;
        RECT 179.400 283.050 180.450 287.400 ;
        RECT 184.950 286.950 187.050 289.050 ;
        RECT 191.400 287.400 192.600 289.650 ;
        RECT 197.400 288.900 198.600 289.650 ;
        RECT 178.950 280.950 181.050 283.050 ;
        RECT 185.400 280.050 186.450 286.950 ;
        RECT 175.950 277.950 178.050 280.050 ;
        RECT 184.950 277.950 187.050 280.050 ;
        RECT 176.400 268.050 177.450 277.950 ;
        RECT 191.400 271.050 192.450 287.400 ;
        RECT 196.950 286.800 199.050 288.900 ;
        RECT 203.400 287.400 204.600 289.650 ;
        RECT 197.400 285.450 198.450 286.800 ;
        RECT 197.400 284.400 201.450 285.450 ;
        RECT 200.400 271.050 201.450 284.400 ;
        RECT 203.400 280.050 204.450 287.400 ;
        RECT 208.950 286.950 211.050 289.050 ;
        RECT 218.400 287.400 219.600 289.650 ;
        RECT 233.400 287.400 234.600 289.650 ;
        RECT 245.400 287.400 246.600 289.650 ;
        RECT 257.400 288.900 258.600 289.650 ;
        RECT 263.400 288.900 264.600 289.650 ;
        RECT 205.800 283.950 207.900 286.050 ;
        RECT 202.950 277.950 205.050 280.050 ;
        RECT 206.400 277.050 207.450 283.950 ;
        RECT 209.400 283.050 210.450 286.950 ;
        RECT 214.950 283.950 217.050 286.050 ;
        RECT 208.950 280.950 211.050 283.050 ;
        RECT 205.950 274.950 208.050 277.050 ;
        RECT 181.950 268.950 184.050 271.050 ;
        RECT 190.950 268.950 193.050 271.050 ;
        RECT 199.950 268.950 202.050 271.050 ;
        RECT 205.950 268.950 208.050 271.050 ;
        RECT 175.950 265.950 178.050 268.050 ;
        RECT 167.400 259.350 168.600 259.950 ;
        RECT 173.400 259.350 174.600 261.600 ;
        RECT 178.950 261.000 181.050 265.050 ;
        RECT 182.400 262.050 183.450 268.950 ;
        RECT 196.950 265.950 199.050 268.050 ;
        RECT 184.950 262.950 190.050 265.050 ;
        RECT 179.400 259.350 180.600 261.000 ;
        RECT 181.950 259.950 184.050 262.050 ;
        RECT 190.950 261.000 193.050 265.050 ;
        RECT 197.400 262.050 198.450 265.950 ;
        RECT 191.400 259.350 192.600 261.000 ;
        RECT 196.950 259.950 199.050 262.050 ;
        RECT 202.950 260.100 205.050 262.200 ;
        RECT 206.400 262.050 207.450 268.950 ;
        RECT 215.400 265.050 216.450 283.950 ;
        RECT 218.400 280.050 219.450 287.400 ;
        RECT 229.950 283.950 232.050 286.050 ;
        RECT 217.950 277.950 220.050 280.050 ;
        RECT 214.950 262.950 217.050 265.050 ;
        RECT 203.400 259.350 204.600 260.100 ;
        RECT 205.950 259.950 208.050 262.050 ;
        RECT 217.950 260.100 220.050 262.200 ;
        RECT 230.400 261.600 231.450 283.950 ;
        RECT 233.400 277.050 234.450 287.400 ;
        RECT 235.950 283.950 238.050 286.050 ;
        RECT 232.950 274.950 235.050 277.050 ;
        RECT 236.400 262.050 237.450 283.950 ;
        RECT 245.400 280.050 246.450 287.400 ;
        RECT 256.950 286.800 259.050 288.900 ;
        RECT 262.950 286.800 265.050 288.900 ;
        RECT 299.400 287.400 300.900 306.300 ;
        RECT 303.300 300.300 304.500 306.300 ;
        RECT 302.400 298.200 304.500 300.300 ;
        RECT 244.950 277.950 247.050 280.050 ;
        RECT 256.950 264.450 259.050 268.050 ;
        RECT 254.400 264.000 259.050 264.450 ;
        RECT 254.400 263.400 258.450 264.000 ;
        RECT 218.400 259.350 219.600 260.100 ;
        RECT 230.400 259.350 231.600 261.600 ;
        RECT 235.950 259.950 238.050 262.050 ;
        RECT 254.400 261.600 255.450 263.400 ;
        RECT 263.400 261.600 264.450 286.800 ;
        RECT 299.400 285.300 301.500 287.400 ;
        RECT 300.300 281.700 301.500 285.300 ;
        RECT 303.300 281.700 304.500 298.200 ;
        RECT 305.700 303.300 307.800 305.400 ;
        RECT 305.700 281.700 306.900 303.300 ;
        RECT 311.400 300.450 312.450 313.950 ;
        RECT 322.200 306.300 324.300 308.400 ;
        RECT 308.400 299.400 312.450 300.450 ;
        RECT 314.400 301.800 316.500 303.900 ;
        RECT 319.800 303.300 321.900 305.400 ;
        RECT 308.400 292.050 309.450 299.400 ;
        RECT 314.400 295.200 315.300 301.800 ;
        RECT 320.100 296.100 321.300 303.300 ;
        RECT 322.800 301.500 324.300 306.300 ;
        RECT 325.200 303.300 327.300 308.400 ;
        RECT 322.800 299.400 324.900 301.500 ;
        RECT 314.400 293.100 316.500 295.200 ;
        RECT 319.800 294.000 321.900 296.100 ;
        RECT 307.800 289.950 309.900 292.050 ;
        RECT 310.950 290.100 313.050 292.200 ;
        RECT 311.400 289.350 312.600 290.100 ;
        RECT 310.800 286.950 312.900 289.050 ;
        RECT 314.400 282.600 315.300 293.100 ;
        RECT 317.100 286.500 319.200 288.600 ;
        RECT 299.700 279.600 301.800 281.700 ;
        RECT 302.700 279.600 304.800 281.700 ;
        RECT 305.700 279.600 307.800 281.700 ;
        RECT 313.800 280.500 315.900 282.600 ;
        RECT 320.100 281.700 321.300 294.000 ;
        RECT 322.800 281.700 324.300 299.400 ;
        RECT 326.100 281.700 327.300 303.300 ;
        RECT 319.200 279.600 321.300 281.700 ;
        RECT 322.200 279.600 324.300 281.700 ;
        RECT 325.200 279.600 327.300 281.700 ;
        RECT 328.200 306.300 330.300 308.400 ;
        RECT 328.200 301.500 329.700 306.300 ;
        RECT 331.950 301.950 334.050 304.050 ;
        RECT 328.200 299.400 330.300 301.500 ;
        RECT 328.200 281.700 329.700 299.400 ;
        RECT 328.200 279.600 330.300 281.700 ;
        RECT 268.950 268.950 271.050 271.050 ;
        RECT 310.950 268.950 313.050 271.050 ;
        RECT 269.400 262.050 270.450 268.950 ;
        RECT 254.400 259.350 255.600 261.600 ;
        RECT 263.400 259.350 264.600 261.600 ;
        RECT 268.950 259.950 271.050 262.050 ;
        RECT 274.950 260.100 277.050 262.200 ;
        RECT 289.950 260.100 292.050 262.200 ;
        RECT 304.950 260.100 307.050 262.200 ;
        RECT 311.400 261.600 312.450 268.950 ;
        RECT 332.400 268.050 333.450 301.950 ;
        RECT 337.800 292.950 339.900 295.050 ;
        RECT 346.800 292.950 348.900 295.050 ;
        RECT 334.950 290.100 337.050 292.200 ;
        RECT 347.400 291.450 348.600 292.650 ;
        RECT 350.400 291.450 351.450 329.400 ;
        RECT 344.400 290.400 351.450 291.450 ;
        RECT 335.400 276.450 336.450 290.100 ;
        RECT 335.400 275.400 339.450 276.450 ;
        RECT 331.950 265.950 334.050 268.050 ;
        RECT 275.400 259.350 276.600 260.100 ;
        RECT 290.400 259.350 291.600 260.100 ;
        RECT 305.400 259.350 306.600 260.100 ;
        RECT 311.400 259.350 312.600 261.600 ;
        RECT 316.950 260.100 319.050 262.200 ;
        RECT 331.950 260.100 334.050 262.200 ;
        RECT 338.400 261.600 339.450 275.400 ;
        RECT 344.400 262.050 345.450 290.400 ;
        RECT 346.950 265.950 349.050 268.050 ;
        RECT 317.400 259.350 318.600 260.100 ;
        RECT 332.400 259.350 333.600 260.100 ;
        RECT 338.400 259.350 339.600 261.600 ;
        RECT 343.950 259.950 346.050 262.050 ;
        RECT 347.400 261.600 348.450 265.950 ;
        RECT 353.400 265.200 354.450 332.400 ;
        RECT 355.950 331.950 358.050 334.050 ;
        RECT 352.950 263.100 355.050 265.200 ;
        RECT 356.400 264.450 357.450 331.950 ;
        RECT 356.400 263.400 360.450 264.450 ;
        RECT 347.400 259.350 348.600 261.600 ;
        RECT 352.950 259.950 355.050 262.050 ;
        RECT 359.400 261.600 360.450 263.400 ;
        RECT 353.400 259.350 354.600 259.950 ;
        RECT 359.400 259.350 360.600 261.600 ;
        RECT 80.400 258.450 81.600 258.600 ;
        RECT 80.400 257.400 84.450 258.450 ;
        RECT 80.400 256.350 81.600 257.400 ;
        RECT 79.800 253.950 81.900 256.050 ;
        RECT 83.400 241.050 84.450 257.400 ;
        RECT 88.950 256.950 91.050 259.050 ;
        RECT 91.950 256.950 94.050 259.050 ;
        RECT 94.950 256.950 97.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 109.950 256.950 112.050 259.050 ;
        RECT 112.950 256.950 115.050 259.050 ;
        RECT 121.950 256.950 124.050 259.050 ;
        RECT 124.950 256.950 127.050 259.050 ;
        RECT 127.950 256.950 130.050 259.050 ;
        RECT 130.950 256.950 133.050 259.050 ;
        RECT 139.950 256.950 142.050 259.050 ;
        RECT 142.950 256.950 145.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 151.950 256.950 154.050 259.050 ;
        RECT 154.950 256.950 157.050 259.050 ;
        RECT 157.950 256.950 160.050 259.050 ;
        RECT 166.950 256.950 169.050 259.050 ;
        RECT 169.950 256.950 172.050 259.050 ;
        RECT 172.950 256.950 175.050 259.050 ;
        RECT 175.950 256.950 178.050 259.050 ;
        RECT 178.950 256.950 181.050 259.050 ;
        RECT 187.950 256.950 190.050 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 193.950 256.950 196.050 259.050 ;
        RECT 199.950 256.950 202.050 259.050 ;
        RECT 202.950 256.950 205.050 259.050 ;
        RECT 212.100 256.950 214.200 259.050 ;
        RECT 217.500 256.950 219.600 259.050 ;
        RECT 220.800 256.950 222.900 259.050 ;
        RECT 226.950 256.950 229.050 259.050 ;
        RECT 229.950 256.950 232.050 259.050 ;
        RECT 232.950 256.950 235.050 259.050 ;
        RECT 239.100 256.950 241.200 259.050 ;
        RECT 244.500 256.950 246.600 259.050 ;
        RECT 253.950 256.950 256.050 259.050 ;
        RECT 256.950 256.950 259.050 259.050 ;
        RECT 262.950 256.950 265.050 259.050 ;
        RECT 265.950 256.950 268.050 259.050 ;
        RECT 271.950 256.950 274.050 259.050 ;
        RECT 274.950 256.950 277.050 259.050 ;
        RECT 277.950 256.950 280.050 259.050 ;
        RECT 286.950 256.950 289.050 259.050 ;
        RECT 289.950 256.950 292.050 259.050 ;
        RECT 292.950 256.950 295.050 259.050 ;
        RECT 295.950 256.950 298.050 259.050 ;
        RECT 298.950 256.950 301.050 259.050 ;
        RECT 301.950 256.950 304.050 259.050 ;
        RECT 304.950 256.950 307.050 259.050 ;
        RECT 310.950 256.950 313.050 259.050 ;
        RECT 313.950 256.950 316.050 259.050 ;
        RECT 316.950 256.950 319.050 259.050 ;
        RECT 319.950 256.950 322.050 259.050 ;
        RECT 328.950 256.950 331.050 259.050 ;
        RECT 331.950 256.950 334.050 259.050 ;
        RECT 334.950 256.950 337.050 259.050 ;
        RECT 337.950 256.950 340.050 259.050 ;
        RECT 346.950 256.950 349.050 259.050 ;
        RECT 349.950 256.950 352.050 259.050 ;
        RECT 352.950 256.950 355.050 259.050 ;
        RECT 355.950 256.950 358.050 259.050 ;
        RECT 358.950 256.950 361.050 259.050 ;
        RECT 85.950 253.950 88.050 256.050 ;
        RECT 89.400 254.400 90.600 256.650 ;
        RECT 95.400 255.900 96.600 256.650 ;
        RECT 86.400 250.050 87.450 253.950 ;
        RECT 85.950 247.950 88.050 250.050 ;
        RECT 82.950 238.950 85.050 241.050 ;
        RECT 89.400 238.050 90.450 254.400 ;
        RECT 94.950 253.800 97.050 255.900 ;
        RECT 104.400 254.400 105.600 256.650 ;
        RECT 110.400 255.000 111.600 256.650 ;
        RECT 104.400 250.050 105.450 254.400 ;
        RECT 109.950 250.950 112.050 255.000 ;
        RECT 125.400 254.400 126.600 256.650 ;
        RECT 131.400 254.400 132.600 256.650 ;
        RECT 140.400 255.900 141.600 256.650 ;
        RECT 149.400 255.900 150.600 256.650 ;
        RECT 121.950 250.950 124.050 253.050 ;
        RECT 103.950 247.950 106.050 250.050 ;
        RECT 94.950 238.950 97.050 241.050 ;
        RECT 34.950 235.950 37.050 238.050 ;
        RECT 43.950 235.950 46.050 238.050 ;
        RECT 73.950 235.950 76.050 238.050 ;
        RECT 88.950 235.950 91.050 238.050 ;
        RECT 35.400 231.450 36.450 235.950 ;
        RECT 32.400 230.400 36.450 231.450 ;
        RECT 7.950 215.100 10.050 217.200 ;
        RECT 16.950 216.000 19.050 220.050 ;
        RECT 32.400 217.050 33.450 230.400 ;
        RECT 55.950 229.950 58.050 232.050 ;
        RECT 76.950 229.950 79.050 232.050 ;
        RECT 43.950 226.950 46.050 229.050 ;
        RECT 37.950 220.950 40.050 223.050 ;
        RECT 26.400 216.450 27.600 216.600 ;
        RECT 26.400 216.000 30.450 216.450 ;
        RECT 8.400 214.350 9.600 215.100 ;
        RECT 17.400 214.350 18.600 216.000 ;
        RECT 26.400 215.400 31.050 216.000 ;
        RECT 26.400 214.350 27.600 215.400 ;
        RECT 7.950 211.950 10.050 214.050 ;
        RECT 10.950 211.950 13.050 214.050 ;
        RECT 17.100 211.950 19.200 214.050 ;
        RECT 20.400 211.950 22.500 214.050 ;
        RECT 25.800 211.950 27.900 214.050 ;
        RECT 28.950 211.950 31.050 215.400 ;
        RECT 31.950 214.950 34.050 217.050 ;
        RECT 38.400 216.600 39.450 220.950 ;
        RECT 44.400 216.600 45.450 226.950 ;
        RECT 56.400 217.200 57.450 229.950 ;
        RECT 73.950 223.950 76.050 226.050 ;
        RECT 38.400 214.350 39.600 216.600 ;
        RECT 44.400 214.350 45.600 216.600 ;
        RECT 55.950 215.100 58.050 217.200 ;
        RECT 63.000 216.900 66.000 217.050 ;
        RECT 63.000 216.600 67.050 216.900 ;
        RECT 56.400 214.350 57.600 215.100 ;
        RECT 62.400 214.950 67.050 216.600 ;
        RECT 62.400 214.350 63.600 214.950 ;
        RECT 64.950 214.800 67.050 214.950 ;
        RECT 74.400 216.600 75.450 223.950 ;
        RECT 77.400 220.050 78.450 229.950 ;
        RECT 82.950 226.950 85.050 229.050 ;
        RECT 76.950 217.950 79.050 220.050 ;
        RECT 83.400 216.600 84.450 226.950 ;
        RECT 74.400 214.350 75.600 216.600 ;
        RECT 83.400 214.350 84.600 216.600 ;
        RECT 91.800 215.100 93.900 217.200 ;
        RECT 95.400 217.050 96.450 238.950 ;
        RECT 103.950 235.950 106.050 238.050 ;
        RECT 100.950 226.950 103.050 229.050 ;
        RECT 92.400 214.350 93.600 215.100 ;
        RECT 94.950 214.950 97.050 217.050 ;
        RECT 101.400 216.600 102.450 226.950 ;
        RECT 104.400 226.050 105.450 235.950 ;
        RECT 103.950 223.950 106.050 226.050 ;
        RECT 106.950 220.950 109.050 223.050 ;
        RECT 112.950 220.950 115.050 223.050 ;
        RECT 107.400 216.600 108.450 220.950 ;
        RECT 113.400 216.600 114.450 220.950 ;
        RECT 122.400 216.600 123.450 250.950 ;
        RECT 125.400 247.050 126.450 254.400 ;
        RECT 124.950 244.950 127.050 247.050 ;
        RECT 131.400 244.050 132.450 254.400 ;
        RECT 139.950 253.800 142.050 255.900 ;
        RECT 148.950 253.800 151.050 255.900 ;
        RECT 160.800 253.950 162.900 256.050 ;
        RECT 176.400 255.900 177.600 256.650 ;
        RECT 188.400 255.900 189.600 256.650 ;
        RECT 194.400 255.900 195.600 256.650 ;
        RECT 130.950 241.950 133.050 244.050 ;
        RECT 140.400 232.050 141.450 253.800 ;
        RECT 145.950 250.950 148.050 253.050 ;
        RECT 142.950 235.950 145.050 238.050 ;
        RECT 130.950 229.950 133.050 232.050 ;
        RECT 139.950 229.950 142.050 232.050 ;
        RECT 101.400 214.350 102.600 216.600 ;
        RECT 107.400 214.350 108.600 216.600 ;
        RECT 113.400 214.350 114.600 216.600 ;
        RECT 122.400 214.350 123.600 216.600 ;
        RECT 127.950 215.100 130.050 217.200 ;
        RECT 131.400 217.050 132.450 229.950 ;
        RECT 34.950 211.950 37.050 214.050 ;
        RECT 37.950 211.950 40.050 214.050 ;
        RECT 40.950 211.950 43.050 214.050 ;
        RECT 43.950 211.950 46.050 214.050 ;
        RECT 52.950 211.950 55.050 214.050 ;
        RECT 55.950 211.950 58.050 214.050 ;
        RECT 58.950 211.950 61.050 214.050 ;
        RECT 61.950 211.950 64.050 214.050 ;
        RECT 70.950 211.950 73.050 214.050 ;
        RECT 73.950 211.950 76.050 214.050 ;
        RECT 76.950 211.950 79.050 214.050 ;
        RECT 83.100 211.950 85.200 214.050 ;
        RECT 86.400 211.950 88.500 214.050 ;
        RECT 91.800 211.950 93.900 214.050 ;
        RECT 97.950 211.950 100.050 214.050 ;
        RECT 100.950 211.950 103.050 214.050 ;
        RECT 103.950 211.950 106.050 214.050 ;
        RECT 106.950 211.950 109.050 214.050 ;
        RECT 113.100 211.950 115.200 214.050 ;
        RECT 116.100 211.950 118.200 214.050 ;
        RECT 121.800 211.950 123.900 214.050 ;
        RECT 124.800 211.950 126.900 214.050 ;
        RECT 4.950 208.950 7.050 211.050 ;
        RECT 11.400 209.400 12.600 211.650 ;
        RECT 20.400 209.400 21.600 211.650 ;
        RECT 35.400 210.900 36.600 211.650 ;
        RECT 5.400 205.050 6.450 208.950 ;
        RECT 4.950 202.950 7.050 205.050 ;
        RECT 11.400 199.050 12.450 209.400 ;
        RECT 20.400 205.050 21.450 209.400 ;
        RECT 28.950 208.800 31.050 210.900 ;
        RECT 34.950 208.800 37.050 210.900 ;
        RECT 41.400 209.400 42.600 211.650 ;
        RECT 19.950 202.950 22.050 205.050 ;
        RECT 29.400 202.050 30.450 208.800 ;
        RECT 41.400 202.050 42.450 209.400 ;
        RECT 49.950 208.950 52.050 211.050 ;
        RECT 53.400 209.400 54.600 211.650 ;
        RECT 59.400 210.900 60.600 211.650 ;
        RECT 28.950 199.950 31.050 202.050 ;
        RECT 40.950 199.950 43.050 202.050 ;
        RECT 1.950 196.950 4.050 199.050 ;
        RECT 10.950 196.950 13.050 199.050 ;
        RECT 1.950 187.950 4.050 190.050 ;
        RECT 17.700 189.300 19.800 191.400 ;
        RECT 20.700 189.300 22.800 191.400 ;
        RECT 23.700 189.300 25.800 191.400 ;
        RECT 2.400 181.050 3.450 187.950 ;
        RECT 18.300 185.700 19.500 189.300 ;
        RECT 17.400 183.600 19.500 185.700 ;
        RECT 1.950 178.950 4.050 181.050 ;
        RECT 4.800 175.950 6.900 178.050 ;
        RECT 10.800 175.950 12.900 178.050 ;
        RECT 1.950 172.950 4.050 175.050 ;
        RECT 2.400 157.050 3.450 172.950 ;
        RECT 17.400 164.700 18.900 183.600 ;
        RECT 21.300 172.800 22.500 189.300 ;
        RECT 20.400 170.700 22.500 172.800 ;
        RECT 21.300 164.700 22.500 170.700 ;
        RECT 23.700 167.700 24.900 189.300 ;
        RECT 31.800 188.400 33.900 190.500 ;
        RECT 37.200 189.300 39.300 191.400 ;
        RECT 40.200 189.300 42.300 191.400 ;
        RECT 43.200 189.300 45.300 191.400 ;
        RECT 28.800 181.950 30.900 184.050 ;
        RECT 29.400 180.900 30.600 181.650 ;
        RECT 28.950 178.800 31.050 180.900 ;
        RECT 32.400 177.900 33.300 188.400 ;
        RECT 35.100 182.400 37.200 184.500 ;
        RECT 32.400 175.800 34.500 177.900 ;
        RECT 38.100 177.000 39.300 189.300 ;
        RECT 32.400 169.200 33.300 175.800 ;
        RECT 37.800 174.900 39.900 177.000 ;
        RECT 23.700 165.600 25.800 167.700 ;
        RECT 28.950 166.950 31.050 169.050 ;
        RECT 32.400 167.100 34.500 169.200 ;
        RECT 38.100 167.700 39.300 174.900 ;
        RECT 40.800 171.600 42.300 189.300 ;
        RECT 40.800 169.500 42.900 171.600 ;
        RECT 17.400 162.600 20.400 164.700 ;
        RECT 21.300 162.600 23.400 164.700 ;
        RECT 1.950 154.950 4.050 157.050 ;
        RECT 13.950 154.950 16.050 157.050 ;
        RECT 14.400 148.050 15.450 154.950 ;
        RECT 17.400 150.300 20.400 152.400 ;
        RECT 21.300 150.300 23.400 152.400 ;
        RECT 13.950 145.950 16.050 148.050 ;
        RECT 4.800 136.950 6.900 139.050 ;
        RECT 10.800 136.950 12.900 139.050 ;
        RECT 4.950 118.950 7.050 121.050 ;
        RECT 14.400 120.450 15.450 145.950 ;
        RECT 17.400 131.400 18.900 150.300 ;
        RECT 21.300 144.300 22.500 150.300 ;
        RECT 20.400 142.200 22.500 144.300 ;
        RECT 17.400 129.300 19.500 131.400 ;
        RECT 18.300 125.700 19.500 129.300 ;
        RECT 21.300 125.700 22.500 142.200 ;
        RECT 23.700 147.300 25.800 149.400 ;
        RECT 23.700 125.700 24.900 147.300 ;
        RECT 29.400 139.050 30.450 166.950 ;
        RECT 37.800 165.600 39.900 167.700 ;
        RECT 40.800 164.700 42.300 169.500 ;
        RECT 44.100 167.700 45.300 189.300 ;
        RECT 40.200 162.600 42.300 164.700 ;
        RECT 43.200 162.600 45.300 167.700 ;
        RECT 46.200 189.300 48.300 191.400 ;
        RECT 50.400 190.050 51.450 208.950 ;
        RECT 53.400 205.050 54.450 209.400 ;
        RECT 58.950 208.800 61.050 210.900 ;
        RECT 71.400 210.000 72.600 211.650 ;
        RECT 77.400 210.000 78.600 211.650 ;
        RECT 61.950 205.950 64.050 208.050 ;
        RECT 64.950 205.950 67.050 208.050 ;
        RECT 70.950 205.950 73.050 210.000 ;
        RECT 76.950 205.950 79.050 210.000 ;
        RECT 86.400 209.400 87.600 211.650 ;
        RECT 98.400 210.900 99.600 211.650 ;
        RECT 104.400 210.900 105.600 211.650 ;
        RECT 86.400 207.450 87.450 209.400 ;
        RECT 97.950 208.800 100.050 210.900 ;
        RECT 103.950 208.800 106.050 210.900 ;
        RECT 125.400 209.400 126.600 211.650 ;
        RECT 86.400 207.000 90.450 207.450 ;
        RECT 86.400 206.400 91.050 207.000 ;
        RECT 52.950 202.950 55.050 205.050 ;
        RECT 52.950 190.950 55.050 193.050 ;
        RECT 46.200 171.600 47.700 189.300 ;
        RECT 49.950 187.950 52.050 190.050 ;
        RECT 53.400 180.900 54.450 190.950 ;
        RECT 62.400 190.050 63.450 205.950 ;
        RECT 65.400 202.050 66.450 205.950 ;
        RECT 88.950 202.950 91.050 206.400 ;
        RECT 125.400 204.450 126.450 209.400 ;
        RECT 128.400 208.050 129.450 215.100 ;
        RECT 130.950 214.950 133.050 217.050 ;
        RECT 133.950 215.100 136.050 217.200 ;
        RECT 143.400 216.600 144.450 235.950 ;
        RECT 146.400 223.050 147.450 250.950 ;
        RECT 161.400 244.050 162.450 253.950 ;
        RECT 175.950 253.800 178.050 255.900 ;
        RECT 187.950 253.800 190.050 255.900 ;
        RECT 193.950 253.800 196.050 255.900 ;
        RECT 200.400 254.400 201.600 256.650 ;
        RECT 200.400 253.050 201.450 254.400 ;
        RECT 205.950 253.950 208.050 256.050 ;
        RECT 212.400 255.900 213.600 256.650 ;
        RECT 163.950 250.950 166.050 253.050 ;
        RECT 200.400 250.950 205.050 253.050 ;
        RECT 164.400 244.050 165.450 250.950 ;
        RECT 200.400 247.050 201.450 250.950 ;
        RECT 199.950 244.950 202.050 247.050 ;
        RECT 206.400 244.050 207.450 253.950 ;
        RECT 211.950 253.800 214.050 255.900 ;
        RECT 221.400 254.400 222.600 256.650 ;
        RECT 227.400 255.900 228.600 256.650 ;
        RECT 151.950 241.950 154.050 244.050 ;
        RECT 160.800 241.950 162.900 244.050 ;
        RECT 163.950 241.950 166.050 244.050 ;
        RECT 205.950 241.950 208.050 244.050 ;
        RECT 148.950 226.950 151.050 229.050 ;
        RECT 145.950 220.950 148.050 223.050 ;
        RECT 149.400 220.050 150.450 226.950 ;
        RECT 148.950 217.950 151.050 220.050 ;
        RECT 152.400 216.600 153.450 241.950 ;
        RECT 161.400 238.050 162.450 241.950 ;
        RECT 169.950 238.950 172.050 241.050 ;
        RECT 190.950 238.950 193.050 241.050 ;
        RECT 160.950 235.950 163.050 238.050 ;
        RECT 134.400 214.350 135.600 215.100 ;
        RECT 143.400 214.350 144.600 216.600 ;
        RECT 152.400 214.350 153.600 216.600 ;
        RECT 158.400 216.450 159.600 216.600 ;
        RECT 155.400 215.400 159.600 216.450 ;
        RECT 133.950 211.950 136.050 214.050 ;
        RECT 136.950 211.950 139.050 214.050 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 143.100 211.950 145.200 214.050 ;
        RECT 148.500 211.950 150.600 214.050 ;
        RECT 151.800 211.950 153.900 214.050 ;
        RECT 130.950 208.950 133.050 211.050 ;
        RECT 137.400 209.400 138.600 211.650 ;
        RECT 149.400 209.400 150.600 211.650 ;
        RECT 127.950 205.950 130.050 208.050 ;
        RECT 131.400 204.450 132.450 208.950 ;
        RECT 133.950 205.950 136.050 208.050 ;
        RECT 125.400 203.400 132.450 204.450 ;
        RECT 64.950 199.950 67.050 202.050 ;
        RECT 104.400 200.400 111.450 201.450 ;
        RECT 104.400 195.450 105.450 200.400 ;
        RECT 101.400 194.400 105.450 195.450 ;
        RECT 94.950 190.950 97.050 193.050 ;
        RECT 61.950 187.950 64.050 190.050 ;
        RECT 67.950 187.950 70.050 190.050 ;
        RECT 68.400 184.200 69.450 187.950 ;
        RECT 67.950 182.100 70.050 184.200 ;
        RECT 79.950 182.100 82.050 184.200 ;
        RECT 85.950 182.100 88.050 184.200 ;
        RECT 95.400 183.600 96.450 190.950 ;
        RECT 101.400 183.600 102.450 194.400 ;
        RECT 103.950 190.950 106.050 193.050 ;
        RECT 104.400 187.050 105.450 190.950 ;
        RECT 110.400 190.050 111.450 200.400 ;
        RECT 118.950 190.950 121.050 193.050 ;
        RECT 130.950 192.450 133.050 193.050 ;
        RECT 125.400 191.400 133.050 192.450 ;
        RECT 109.950 187.950 112.050 190.050 ;
        RECT 115.950 187.950 118.050 190.050 ;
        RECT 103.800 184.950 105.900 187.050 ;
        RECT 116.400 183.600 117.450 187.950 ;
        RECT 119.400 187.050 120.450 190.950 ;
        RECT 118.950 184.950 121.050 187.050 ;
        RECT 125.400 186.450 126.450 191.400 ;
        RECT 130.950 190.950 133.050 191.400 ;
        RECT 122.400 186.000 126.450 186.450 ;
        RECT 121.950 185.400 126.450 186.000 ;
        RECT 52.800 178.800 54.900 180.900 ;
        RECT 64.950 179.100 67.050 181.200 ;
        RECT 65.400 178.350 66.600 179.100 ;
        RECT 68.400 178.050 69.450 182.100 ;
        RECT 80.400 181.350 81.600 182.100 ;
        RECT 86.400 181.350 87.600 182.100 ;
        RECT 95.400 181.350 96.600 183.600 ;
        RECT 101.400 181.350 102.600 183.600 ;
        RECT 116.400 181.350 117.600 183.600 ;
        RECT 121.950 181.950 124.050 185.400 ;
        RECT 127.950 183.000 130.050 187.050 ;
        RECT 134.400 184.050 135.450 205.950 ;
        RECT 137.400 202.050 138.450 209.400 ;
        RECT 139.950 205.950 142.050 208.050 ;
        RECT 136.950 199.950 139.050 202.050 ;
        RECT 140.400 193.050 141.450 205.950 ;
        RECT 149.400 205.050 150.450 209.400 ;
        RECT 155.400 205.050 156.450 215.400 ;
        RECT 158.400 214.350 159.600 215.400 ;
        RECT 166.950 214.950 169.050 217.050 ;
        RECT 167.400 214.350 168.600 214.950 ;
        RECT 158.100 211.950 160.200 214.050 ;
        RECT 161.400 211.950 163.500 214.050 ;
        RECT 166.800 211.950 168.900 214.050 ;
        RECT 170.400 208.050 171.450 238.950 ;
        RECT 187.950 217.950 190.050 220.050 ;
        RECT 178.950 215.100 181.050 217.200 ;
        RECT 179.400 214.350 180.600 215.100 ;
        RECT 175.950 211.950 178.050 214.050 ;
        RECT 178.950 211.950 181.050 214.050 ;
        RECT 181.950 211.950 184.050 214.050 ;
        RECT 176.400 210.000 177.600 211.650 ;
        RECT 182.400 210.900 183.600 211.650 ;
        RECT 157.950 205.950 160.050 208.050 ;
        RECT 169.950 205.950 172.050 208.050 ;
        RECT 175.950 205.950 178.050 210.000 ;
        RECT 181.950 208.800 184.050 210.900 ;
        RECT 148.950 202.950 151.050 205.050 ;
        RECT 154.950 202.950 157.050 205.050 ;
        RECT 155.400 193.050 156.450 202.950 ;
        RECT 158.400 202.050 159.450 205.950 ;
        RECT 188.400 205.050 189.450 217.950 ;
        RECT 191.400 216.600 192.450 238.950 ;
        RECT 206.400 229.050 207.450 241.950 ;
        RECT 205.950 226.950 208.050 229.050 ;
        RECT 221.400 220.200 222.450 254.400 ;
        RECT 226.950 253.800 229.050 255.900 ;
        RECT 235.950 253.950 238.050 256.050 ;
        RECT 239.400 254.400 240.600 256.650 ;
        RECT 257.400 255.900 258.600 256.650 ;
        RECT 227.400 238.050 228.450 253.800 ;
        RECT 236.400 250.050 237.450 253.950 ;
        RECT 235.950 247.950 238.050 250.050 ;
        RECT 226.950 235.950 229.050 238.050 ;
        RECT 239.400 229.050 240.450 254.400 ;
        RECT 256.950 253.800 259.050 255.900 ;
        RECT 266.400 254.400 267.600 256.650 ;
        RECT 259.950 250.950 262.050 253.050 ;
        RECT 238.950 226.950 241.050 229.050 ;
        RECT 226.950 220.950 229.050 223.050 ;
        RECT 191.400 214.350 192.600 216.600 ;
        RECT 199.950 216.000 202.050 220.050 ;
        RECT 200.400 214.350 201.600 216.000 ;
        RECT 208.950 215.100 211.050 217.200 ;
        RECT 209.400 214.350 210.600 215.100 ;
        RECT 214.950 214.950 217.050 220.050 ;
        RECT 220.950 218.100 223.050 220.200 ;
        RECT 220.950 214.950 223.050 217.050 ;
        RECT 227.400 216.600 228.450 220.950 ;
        RECT 239.400 219.450 240.450 226.950 ;
        RECT 260.400 220.050 261.450 250.950 ;
        RECT 266.400 250.050 267.450 254.400 ;
        RECT 268.950 253.950 271.050 256.050 ;
        RECT 280.800 255.000 282.900 256.050 ;
        RECT 280.800 253.950 283.050 255.000 ;
        RECT 283.950 253.950 286.050 256.050 ;
        RECT 287.400 255.000 288.600 256.650 ;
        RECT 293.400 255.900 294.600 256.650 ;
        RECT 296.400 255.900 297.600 256.650 ;
        RECT 265.950 247.950 268.050 250.050 ;
        RECT 269.400 246.450 270.450 253.950 ;
        RECT 280.950 250.950 283.050 253.950 ;
        RECT 266.400 245.400 270.450 246.450 ;
        RECT 262.950 220.950 265.050 223.050 ;
        RECT 236.400 218.400 240.450 219.450 ;
        RECT 236.400 216.600 237.450 218.400 ;
        RECT 221.400 214.350 222.600 214.950 ;
        RECT 227.400 214.350 228.600 216.600 ;
        RECT 236.400 214.350 237.600 216.600 ;
        RECT 241.950 216.000 244.050 220.050 ;
        RECT 259.950 217.950 262.050 220.050 ;
        RECT 242.400 214.350 243.600 216.000 ;
        RECT 253.950 215.100 256.050 217.200 ;
        RECT 263.400 216.600 264.450 220.950 ;
        RECT 266.400 217.050 267.450 245.400 ;
        RECT 284.400 244.050 285.450 253.950 ;
        RECT 286.950 250.950 289.050 255.000 ;
        RECT 292.950 253.800 295.050 255.900 ;
        RECT 295.950 253.800 298.050 255.900 ;
        RECT 314.400 254.400 315.600 256.650 ;
        RECT 320.400 254.400 321.600 256.650 ;
        RECT 283.950 241.950 286.050 244.050 ;
        RECT 271.950 238.950 274.050 241.050 ;
        RECT 272.400 229.050 273.450 238.950 ;
        RECT 314.400 235.050 315.450 254.400 ;
        RECT 320.400 244.050 321.450 254.400 ;
        RECT 325.800 253.950 327.900 256.050 ;
        RECT 329.400 255.900 330.600 256.650 ;
        RECT 326.400 250.050 327.450 253.950 ;
        RECT 328.950 253.800 331.050 255.900 ;
        RECT 335.400 254.400 336.600 256.650 ;
        RECT 325.950 247.950 328.050 250.050 ;
        RECT 319.950 241.950 322.050 244.050 ;
        RECT 313.950 232.950 316.050 235.050 ;
        RECT 326.400 232.050 327.450 247.950 ;
        RECT 335.400 247.050 336.450 254.400 ;
        RECT 340.800 253.950 342.900 256.050 ;
        RECT 343.950 253.950 346.050 256.050 ;
        RECT 356.400 254.400 357.600 256.650 ;
        RECT 334.950 244.950 337.050 247.050 ;
        RECT 307.950 229.950 310.050 232.050 ;
        RECT 325.950 229.950 328.050 232.050 ;
        RECT 271.950 226.950 274.050 229.050 ;
        RECT 295.950 226.950 298.050 229.050 ;
        RECT 254.400 214.350 255.600 215.100 ;
        RECT 263.400 214.350 264.600 216.600 ;
        RECT 265.950 214.950 268.050 217.050 ;
        RECT 272.400 216.600 273.450 226.950 ;
        RECT 277.950 220.950 280.050 223.050 ;
        RECT 278.400 216.600 279.450 220.950 ;
        RECT 296.400 217.200 297.450 226.950 ;
        RECT 301.950 220.950 304.050 223.050 ;
        RECT 272.400 214.350 273.600 216.600 ;
        RECT 278.400 214.350 279.600 216.600 ;
        RECT 289.950 215.100 292.050 217.200 ;
        RECT 295.950 215.100 298.050 217.200 ;
        RECT 302.400 216.600 303.450 220.950 ;
        RECT 308.400 217.050 309.450 229.950 ;
        RECT 341.400 226.050 342.450 253.950 ;
        RECT 344.400 246.450 345.450 253.950 ;
        RECT 352.950 250.950 355.050 253.050 ;
        RECT 353.400 247.050 354.450 250.950 ;
        RECT 356.400 250.050 357.450 254.400 ;
        RECT 358.950 250.950 361.050 253.050 ;
        RECT 355.950 247.950 358.050 250.050 ;
        RECT 344.400 245.400 348.450 246.450 ;
        RECT 328.950 223.950 331.050 226.050 ;
        RECT 340.950 223.950 343.050 226.050 ;
        RECT 290.400 214.350 291.600 215.100 ;
        RECT 296.400 214.350 297.600 215.100 ;
        RECT 302.400 214.350 303.600 216.600 ;
        RECT 307.950 214.950 310.050 217.050 ;
        RECT 329.400 216.600 330.450 223.950 ;
        RECT 341.400 216.600 342.450 223.950 ;
        RECT 347.400 217.050 348.450 245.400 ;
        RECT 352.950 244.950 355.050 247.050 ;
        RECT 359.400 235.050 360.450 250.950 ;
        RECT 358.950 232.950 361.050 235.050 ;
        RECT 352.950 220.950 355.050 223.050 ;
        RECT 317.400 216.450 318.600 216.600 ;
        RECT 323.400 216.450 324.600 216.600 ;
        RECT 317.400 215.400 324.600 216.450 ;
        RECT 317.400 214.350 318.600 215.400 ;
        RECT 323.400 214.350 324.600 215.400 ;
        RECT 329.400 214.350 330.600 216.600 ;
        RECT 341.400 214.350 342.600 216.600 ;
        RECT 346.950 214.950 349.050 217.050 ;
        RECT 353.400 216.600 354.450 220.950 ;
        RECT 359.400 220.050 360.450 232.950 ;
        RECT 358.950 217.950 361.050 220.050 ;
        RECT 359.400 216.600 360.450 217.950 ;
        RECT 353.400 214.350 354.600 216.600 ;
        RECT 359.400 214.350 360.600 216.600 ;
        RECT 191.100 211.950 193.200 214.050 ;
        RECT 196.500 211.950 198.600 214.050 ;
        RECT 199.800 211.950 201.900 214.050 ;
        RECT 208.950 211.950 211.050 214.050 ;
        RECT 211.950 211.950 214.050 214.050 ;
        RECT 217.950 211.950 220.050 214.050 ;
        RECT 220.950 211.950 223.050 214.050 ;
        RECT 223.950 211.950 226.050 214.050 ;
        RECT 226.950 211.950 229.050 214.050 ;
        RECT 235.950 211.950 238.050 214.050 ;
        RECT 238.950 211.950 241.050 214.050 ;
        RECT 241.950 211.950 244.050 214.050 ;
        RECT 244.950 211.950 247.050 214.050 ;
        RECT 254.100 211.950 256.200 214.050 ;
        RECT 259.500 211.950 261.600 214.050 ;
        RECT 262.800 211.950 264.900 214.050 ;
        RECT 268.950 211.950 271.050 214.050 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 277.950 211.950 280.050 214.050 ;
        RECT 286.950 211.950 289.050 214.050 ;
        RECT 289.950 211.950 292.050 214.050 ;
        RECT 292.950 211.950 295.050 214.050 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 301.950 211.950 304.050 214.050 ;
        RECT 304.950 211.950 307.050 214.050 ;
        RECT 313.950 211.950 316.050 214.050 ;
        RECT 316.950 211.950 319.050 214.050 ;
        RECT 322.950 211.950 325.050 214.050 ;
        RECT 325.950 211.950 328.050 214.050 ;
        RECT 328.950 211.950 331.050 214.050 ;
        RECT 331.950 211.950 334.050 214.050 ;
        RECT 340.950 211.950 343.050 214.050 ;
        RECT 343.950 211.950 346.050 214.050 ;
        RECT 349.950 211.950 352.050 214.050 ;
        RECT 352.950 211.950 355.050 214.050 ;
        RECT 355.950 211.950 358.050 214.050 ;
        RECT 358.950 211.950 361.050 214.050 ;
        RECT 197.400 210.900 198.600 211.650 ;
        RECT 196.950 208.800 199.050 210.900 ;
        RECT 205.950 208.950 208.050 211.050 ;
        RECT 212.400 210.000 213.600 211.650 ;
        RECT 187.950 202.950 190.050 205.050 ;
        RECT 157.950 199.950 160.050 202.050 ;
        RECT 187.950 199.800 190.050 201.900 ;
        RECT 199.950 199.950 202.050 202.050 ;
        RECT 139.950 190.950 142.050 193.050 ;
        RECT 154.950 190.950 157.050 193.050 ;
        RECT 172.950 190.950 175.050 193.050 ;
        RECT 139.950 187.800 142.050 189.900 ;
        RECT 166.950 187.950 169.050 190.050 ;
        RECT 140.400 184.200 141.450 187.800 ;
        RECT 128.400 181.350 129.600 183.000 ;
        RECT 133.950 181.950 136.050 184.050 ;
        RECT 139.950 182.100 142.050 184.200 ;
        RECT 148.950 182.100 151.050 184.200 ;
        RECT 167.400 183.600 168.450 187.950 ;
        RECT 173.400 184.200 174.450 190.950 ;
        RECT 140.400 181.350 141.600 182.100 ;
        RECT 149.400 181.350 150.600 182.100 ;
        RECT 167.400 181.350 168.600 183.600 ;
        RECT 172.950 182.100 175.050 184.200 ;
        RECT 188.400 183.600 189.450 199.800 ;
        RECT 173.400 181.350 174.600 182.100 ;
        RECT 188.400 181.350 189.600 183.600 ;
        RECT 200.400 181.050 201.450 199.950 ;
        RECT 206.400 199.050 207.450 208.950 ;
        RECT 211.950 205.950 214.050 210.000 ;
        RECT 214.950 208.950 217.050 211.050 ;
        RECT 218.400 209.400 219.600 211.650 ;
        RECT 224.400 209.400 225.600 211.650 ;
        RECT 215.400 202.050 216.450 208.950 ;
        RECT 218.400 205.050 219.450 209.400 ;
        RECT 217.950 202.950 220.050 205.050 ;
        RECT 214.950 199.950 217.050 202.050 ;
        RECT 205.950 196.950 208.050 199.050 ;
        RECT 224.400 196.050 225.450 209.400 ;
        RECT 229.950 208.950 232.050 211.050 ;
        RECT 239.400 210.000 240.600 211.650 ;
        RECT 245.400 210.900 246.600 211.650 ;
        RECT 230.400 202.050 231.450 208.950 ;
        RECT 238.950 205.950 241.050 210.000 ;
        RECT 244.950 208.800 247.050 210.900 ;
        RECT 260.400 209.400 261.600 211.650 ;
        RECT 256.950 205.950 259.050 208.050 ;
        RECT 229.950 199.950 232.050 202.050 ;
        RECT 205.950 193.800 208.050 195.900 ;
        RECT 223.950 193.950 226.050 196.050 ;
        RECT 206.400 187.050 207.450 193.800 ;
        RECT 209.700 189.300 211.800 191.400 ;
        RECT 212.700 189.300 214.800 191.400 ;
        RECT 215.700 189.300 217.800 191.400 ;
        RECT 205.950 184.950 208.050 187.050 ;
        RECT 210.300 185.700 211.500 189.300 ;
        RECT 209.400 183.600 211.500 185.700 ;
        RECT 76.950 178.950 79.050 181.050 ;
        RECT 79.950 178.950 82.050 181.050 ;
        RECT 82.950 178.950 85.050 181.050 ;
        RECT 85.950 178.950 88.050 181.050 ;
        RECT 94.950 178.950 97.050 181.050 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 100.950 178.950 103.050 181.050 ;
        RECT 103.950 178.950 106.050 181.050 ;
        RECT 112.950 178.950 115.050 181.050 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 118.950 178.950 121.050 181.050 ;
        RECT 124.950 178.950 127.050 181.050 ;
        RECT 127.950 178.950 130.050 181.050 ;
        RECT 130.950 178.950 133.050 181.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 148.950 178.950 151.050 181.050 ;
        RECT 151.950 178.950 154.050 181.050 ;
        RECT 154.950 178.950 157.050 181.050 ;
        RECT 157.950 178.950 160.050 181.050 ;
        RECT 166.950 178.950 169.050 181.050 ;
        RECT 169.950 178.950 172.050 181.050 ;
        RECT 172.950 178.950 175.050 181.050 ;
        RECT 175.950 178.950 178.050 181.050 ;
        RECT 184.950 178.950 187.050 181.050 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 190.950 178.950 193.050 181.050 ;
        RECT 199.950 178.950 202.050 181.050 ;
        RECT 49.950 175.950 52.050 178.050 ;
        RECT 55.800 175.950 57.900 178.050 ;
        RECT 64.800 175.950 66.900 178.050 ;
        RECT 67.950 175.950 70.050 178.050 ;
        RECT 46.200 169.500 48.300 171.600 ;
        RECT 46.200 164.700 47.700 169.500 ;
        RECT 46.200 162.600 48.300 164.700 ;
        RECT 40.200 150.300 42.300 152.400 ;
        RECT 32.400 145.800 34.500 147.900 ;
        RECT 37.800 147.300 39.900 149.400 ;
        RECT 32.400 139.200 33.300 145.800 ;
        RECT 38.100 140.100 39.300 147.300 ;
        RECT 40.800 145.500 42.300 150.300 ;
        RECT 43.200 147.300 45.300 152.400 ;
        RECT 40.800 143.400 42.900 145.500 ;
        RECT 28.950 136.950 31.050 139.050 ;
        RECT 32.400 137.100 34.500 139.200 ;
        RECT 37.800 138.000 39.900 140.100 ;
        RECT 25.950 135.600 30.000 136.050 ;
        RECT 25.950 133.950 30.600 135.600 ;
        RECT 29.400 133.350 30.600 133.950 ;
        RECT 28.800 130.950 30.900 133.050 ;
        RECT 32.400 126.600 33.300 137.100 ;
        RECT 35.100 130.500 37.200 132.600 ;
        RECT 17.700 123.600 19.800 125.700 ;
        RECT 20.700 123.600 22.800 125.700 ;
        RECT 23.700 123.600 25.800 125.700 ;
        RECT 31.800 124.500 33.900 126.600 ;
        RECT 38.100 125.700 39.300 138.000 ;
        RECT 40.800 125.700 42.300 143.400 ;
        RECT 44.100 125.700 45.300 147.300 ;
        RECT 37.200 123.600 39.300 125.700 ;
        RECT 40.200 123.600 42.300 125.700 ;
        RECT 43.200 123.600 45.300 125.700 ;
        RECT 46.200 150.300 48.300 152.400 ;
        RECT 46.200 145.500 47.700 150.300 ;
        RECT 46.200 143.400 48.300 145.500 ;
        RECT 46.200 125.700 47.700 143.400 ;
        RECT 46.200 123.600 48.300 125.700 ;
        RECT 14.400 119.400 18.450 120.450 ;
        RECT 1.950 73.950 4.050 76.050 ;
        RECT 2.400 60.450 3.450 73.950 ;
        RECT 5.400 67.050 6.450 118.950 ;
        RECT 13.950 112.950 16.050 115.050 ;
        RECT 14.400 105.600 15.450 112.950 ;
        RECT 17.400 112.050 18.450 119.400 ;
        RECT 50.400 118.050 51.450 175.950 ;
        RECT 67.950 172.800 70.050 174.900 ;
        RECT 73.950 172.950 76.050 178.050 ;
        RECT 77.400 176.400 78.600 178.650 ;
        RECT 83.400 177.000 84.600 178.650 ;
        RECT 55.800 136.950 57.900 139.050 ;
        RECT 64.800 136.950 66.900 139.050 ;
        RECT 52.950 133.950 55.050 136.050 ;
        RECT 65.400 135.900 66.600 136.650 ;
        RECT 53.400 124.050 54.450 133.950 ;
        RECT 64.950 133.800 67.050 135.900 ;
        RECT 65.400 124.050 66.450 133.800 ;
        RECT 52.950 121.950 55.050 124.050 ;
        RECT 58.950 121.950 61.050 124.050 ;
        RECT 64.950 121.950 67.050 124.050 ;
        RECT 25.950 115.950 28.050 118.050 ;
        RECT 49.950 115.950 52.050 118.050 ;
        RECT 16.950 109.950 19.050 112.050 ;
        RECT 26.400 106.200 27.450 115.950 ;
        RECT 37.950 112.950 40.050 115.050 ;
        RECT 31.950 109.950 34.050 112.050 ;
        RECT 14.400 103.350 15.600 105.600 ;
        RECT 25.950 104.100 28.050 106.200 ;
        RECT 32.400 105.600 33.450 109.950 ;
        RECT 38.400 105.600 39.450 112.950 ;
        RECT 46.950 109.950 49.050 112.050 ;
        RECT 47.400 106.050 48.450 109.950 ;
        RECT 26.400 103.350 27.600 104.100 ;
        RECT 32.400 103.350 33.600 105.600 ;
        RECT 38.400 103.350 39.600 105.600 ;
        RECT 46.950 103.950 49.050 106.050 ;
        RECT 50.400 105.600 51.450 115.950 ;
        RECT 59.400 115.050 60.450 121.950 ;
        RECT 58.950 112.950 61.050 115.050 ;
        RECT 59.400 105.600 60.450 112.950 ;
        RECT 68.400 105.600 69.450 172.800 ;
        RECT 77.400 165.450 78.450 176.400 ;
        RECT 82.950 172.950 85.050 177.000 ;
        RECT 88.950 175.950 91.050 178.050 ;
        RECT 98.400 177.900 99.600 178.650 ;
        RECT 104.400 177.900 105.600 178.650 ;
        RECT 89.400 169.050 90.450 175.950 ;
        RECT 97.950 175.800 100.050 177.900 ;
        RECT 103.800 175.800 105.900 177.900 ;
        RECT 113.400 177.450 114.600 178.650 ;
        RECT 110.400 176.400 114.600 177.450 ;
        RECT 119.400 176.400 120.600 178.650 ;
        RECT 91.950 172.950 94.050 175.050 ;
        RECT 88.950 166.950 91.050 169.050 ;
        RECT 74.400 164.400 78.450 165.450 ;
        RECT 74.400 148.050 75.450 164.400 ;
        RECT 92.400 154.050 93.450 172.950 ;
        RECT 110.400 169.050 111.450 176.400 ;
        RECT 119.400 172.050 120.450 176.400 ;
        RECT 121.950 175.950 124.050 178.050 ;
        RECT 125.400 176.400 126.600 178.650 ;
        RECT 137.400 178.050 138.600 178.650 ;
        RECT 133.950 176.400 138.600 178.050 ;
        RECT 152.400 176.400 153.600 178.650 ;
        RECT 158.400 177.900 159.600 178.650 ;
        RECT 118.950 169.950 121.050 172.050 ;
        RECT 109.950 166.950 112.050 169.050 ;
        RECT 119.400 157.050 120.450 169.950 ;
        RECT 118.950 154.950 121.050 157.050 ;
        RECT 91.950 151.950 94.050 154.050 ;
        RECT 73.950 145.950 76.050 148.050 ;
        RECT 97.950 145.950 100.050 148.050 ;
        RECT 118.950 145.950 121.050 148.050 ;
        RECT 73.950 137.100 76.050 139.200 ;
        RECT 79.950 137.100 82.050 142.050 ;
        RECT 91.950 137.100 94.050 139.200 ;
        RECT 98.400 138.600 99.450 145.950 ;
        RECT 106.950 142.950 109.050 145.050 ;
        RECT 107.400 138.600 108.450 142.950 ;
        RECT 74.400 136.350 75.600 137.100 ;
        RECT 80.400 136.350 81.600 137.100 ;
        RECT 92.400 136.350 93.600 137.100 ;
        RECT 98.400 136.350 99.600 138.600 ;
        RECT 107.400 136.350 108.600 138.600 ;
        RECT 112.950 138.000 115.050 142.050 ;
        RECT 119.400 139.050 120.450 145.950 ;
        RECT 113.400 136.350 114.600 138.000 ;
        RECT 118.950 136.950 121.050 139.050 ;
        RECT 122.400 138.600 123.450 175.950 ;
        RECT 125.400 168.450 126.450 176.400 ;
        RECT 133.950 175.950 138.000 176.400 ;
        RECT 127.950 172.950 130.050 175.050 ;
        RECT 136.950 172.950 139.050 175.050 ;
        RECT 145.950 172.950 148.050 175.050 ;
        RECT 152.400 174.450 153.450 176.400 ;
        RECT 157.950 175.800 160.050 177.900 ;
        RECT 176.400 176.400 177.600 178.650 ;
        RECT 185.400 176.400 186.600 178.650 ;
        RECT 152.400 173.400 156.450 174.450 ;
        RECT 128.400 168.450 129.450 172.950 ;
        RECT 130.950 169.950 133.050 172.050 ;
        RECT 125.400 168.000 129.450 168.450 ;
        RECT 125.400 167.400 130.050 168.000 ;
        RECT 127.950 163.950 130.050 167.400 ;
        RECT 127.950 154.950 130.050 157.050 ;
        RECT 128.400 142.050 129.450 154.950 ;
        RECT 131.400 154.050 132.450 169.950 ;
        RECT 130.950 151.950 133.050 154.050 ;
        RECT 130.950 142.950 133.050 145.050 ;
        RECT 127.950 139.950 130.050 142.050 ;
        RECT 122.400 136.350 123.600 138.600 ;
        RECT 128.400 138.450 129.600 138.600 ;
        RECT 131.400 138.450 132.450 142.950 ;
        RECT 128.400 137.400 132.450 138.450 ;
        RECT 137.400 138.600 138.450 172.950 ;
        RECT 139.950 154.950 142.050 157.050 ;
        RECT 140.400 145.050 141.450 154.950 ;
        RECT 139.950 142.950 142.050 145.050 ;
        RECT 146.400 142.050 147.450 172.950 ;
        RECT 155.400 166.050 156.450 173.400 ;
        RECT 158.400 172.050 159.450 175.800 ;
        RECT 157.950 169.950 160.050 172.050 ;
        RECT 154.950 163.950 157.050 166.050 ;
        RECT 145.950 139.950 148.050 142.050 ;
        RECT 155.400 139.200 156.450 163.950 ;
        RECT 176.400 157.050 177.450 176.400 ;
        RECT 185.400 172.050 186.450 176.400 ;
        RECT 196.800 175.950 198.900 178.050 ;
        RECT 202.800 175.950 204.900 178.050 ;
        RECT 187.950 172.950 190.050 175.050 ;
        RECT 184.950 169.950 187.050 172.050 ;
        RECT 160.950 154.950 163.050 157.050 ;
        RECT 175.950 154.950 178.050 157.050 ;
        RECT 128.400 136.350 129.600 137.400 ;
        RECT 137.400 136.350 138.600 138.600 ;
        RECT 154.950 137.100 157.050 139.200 ;
        RECT 161.400 139.050 162.450 154.950 ;
        RECT 175.950 142.950 178.050 145.050 ;
        RECT 176.400 139.200 177.450 142.950 ;
        RECT 155.400 136.350 156.600 137.100 ;
        RECT 160.950 136.950 163.050 139.050 ;
        RECT 169.950 137.100 172.050 139.200 ;
        RECT 175.950 137.100 178.050 139.200 ;
        RECT 170.400 136.350 171.600 137.100 ;
        RECT 176.400 136.350 177.600 137.100 ;
        RECT 73.950 133.950 76.050 136.050 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 88.950 133.950 91.050 136.050 ;
        RECT 91.950 133.950 94.050 136.050 ;
        RECT 94.950 133.950 97.050 136.050 ;
        RECT 97.950 133.950 100.050 136.050 ;
        RECT 106.950 133.950 109.050 136.050 ;
        RECT 109.950 133.950 112.050 136.050 ;
        RECT 112.950 133.950 115.050 136.050 ;
        RECT 115.950 133.950 118.050 136.050 ;
        RECT 121.950 133.950 124.050 136.050 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 133.950 133.950 136.050 136.050 ;
        RECT 136.950 133.950 139.050 136.050 ;
        RECT 139.950 133.950 142.050 136.050 ;
        RECT 142.950 133.950 145.050 136.050 ;
        RECT 145.950 133.950 148.050 136.050 ;
        RECT 154.950 133.950 157.050 136.050 ;
        RECT 157.950 133.950 160.050 136.050 ;
        RECT 166.950 133.950 169.050 136.050 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 175.950 133.950 178.050 136.050 ;
        RECT 178.950 133.950 181.050 136.050 ;
        RECT 181.950 133.950 184.050 136.050 ;
        RECT 77.400 131.400 78.600 133.650 ;
        RECT 70.950 127.950 73.050 130.050 ;
        RECT 71.400 109.050 72.450 127.950 ;
        RECT 77.400 118.050 78.450 131.400 ;
        RECT 85.950 130.950 88.050 133.050 ;
        RECT 89.400 131.400 90.600 133.650 ;
        RECT 95.400 131.400 96.600 133.650 ;
        RECT 110.400 132.900 111.600 133.650 ;
        RECT 76.950 115.950 79.050 118.050 ;
        RECT 86.400 115.050 87.450 130.950 ;
        RECT 89.400 127.050 90.450 131.400 ;
        RECT 95.400 130.050 96.450 131.400 ;
        RECT 109.950 130.800 112.050 132.900 ;
        RECT 116.400 132.000 117.600 133.650 ;
        RECT 125.400 132.900 126.600 133.650 ;
        RECT 91.950 128.400 96.450 130.050 ;
        RECT 91.950 127.950 96.000 128.400 ;
        RECT 97.950 127.950 100.050 130.050 ;
        RECT 115.950 127.950 118.050 132.000 ;
        RECT 124.950 130.800 127.050 132.900 ;
        RECT 134.400 131.400 135.600 133.650 ;
        RECT 140.400 131.400 141.600 133.650 ;
        RECT 146.400 131.400 147.600 133.650 ;
        RECT 158.400 132.900 159.600 133.650 ;
        RECT 88.950 124.950 91.050 127.050 ;
        RECT 98.400 124.050 99.450 127.950 ;
        RECT 97.950 121.950 100.050 124.050 ;
        RECT 103.950 121.950 106.050 124.050 ;
        RECT 121.950 121.950 124.050 124.050 ;
        RECT 97.950 115.950 100.050 118.050 ;
        RECT 85.950 112.950 88.050 115.050 ;
        RECT 70.950 106.950 73.050 109.050 ;
        RECT 50.400 103.350 51.600 105.600 ;
        RECT 59.400 103.350 60.600 105.600 ;
        RECT 68.400 103.350 69.600 105.600 ;
        RECT 73.950 104.100 76.050 106.200 ;
        RECT 86.400 105.600 87.450 112.950 ;
        RECT 98.400 109.050 99.450 115.950 ;
        RECT 104.400 112.050 105.450 121.950 ;
        RECT 112.950 118.950 115.050 121.050 ;
        RECT 103.950 109.950 106.050 112.050 ;
        RECT 113.400 109.050 114.450 118.950 ;
        RECT 122.400 117.450 123.450 121.950 ;
        RECT 134.400 121.050 135.450 131.400 ;
        RECT 140.400 124.050 141.450 131.400 ;
        RECT 146.400 127.050 147.450 131.400 ;
        RECT 157.950 127.950 160.050 132.900 ;
        RECT 163.950 130.950 166.050 133.050 ;
        RECT 167.400 132.000 168.600 133.650 ;
        RECT 145.950 124.950 148.050 127.050 ;
        RECT 139.950 121.950 142.050 124.050 ;
        RECT 133.950 118.950 136.050 121.050 ;
        RECT 157.950 118.950 160.050 121.050 ;
        RECT 116.400 116.400 123.450 117.450 ;
        RECT 116.400 112.050 117.450 116.400 ;
        RECT 115.950 109.950 118.050 112.050 ;
        RECT 122.700 111.300 124.800 113.400 ;
        RECT 125.700 111.300 127.800 113.400 ;
        RECT 128.700 111.300 130.800 113.400 ;
        RECT 97.950 106.950 100.050 109.050 ;
        RECT 112.950 106.950 115.050 109.050 ;
        RECT 123.300 107.700 124.500 111.300 ;
        RECT 74.400 103.350 75.600 104.100 ;
        RECT 86.400 103.350 87.600 105.600 ;
        RECT 91.950 104.100 94.050 106.200 ;
        RECT 122.400 105.600 124.500 107.700 ;
        RECT 92.400 103.350 93.600 104.100 ;
        RECT 8.100 100.950 10.200 103.050 ;
        RECT 13.500 100.950 15.600 103.050 ;
        RECT 20.100 100.950 22.200 103.050 ;
        RECT 25.500 100.950 27.600 103.050 ;
        RECT 31.950 100.950 34.050 103.050 ;
        RECT 34.950 100.950 37.050 103.050 ;
        RECT 37.950 100.950 40.050 103.050 ;
        RECT 40.950 100.950 43.050 103.050 ;
        RECT 49.950 100.950 52.050 103.050 ;
        RECT 52.950 100.950 55.050 103.050 ;
        RECT 58.950 100.950 61.050 103.050 ;
        RECT 61.950 100.950 64.050 103.050 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 70.950 100.950 73.050 103.050 ;
        RECT 73.950 100.950 76.050 103.050 ;
        RECT 82.950 100.950 85.050 103.050 ;
        RECT 85.950 100.950 88.050 103.050 ;
        RECT 92.100 100.950 94.200 103.050 ;
        RECT 95.100 100.950 97.200 103.050 ;
        RECT 100.800 100.950 102.900 103.050 ;
        RECT 103.800 100.950 105.900 103.050 ;
        RECT 35.400 99.900 36.600 100.650 ;
        RECT 41.400 99.900 42.600 100.650 ;
        RECT 34.950 97.800 37.050 99.900 ;
        RECT 40.950 97.800 43.050 99.900 ;
        RECT 53.400 98.400 54.600 100.650 ;
        RECT 62.400 99.900 63.600 100.650 ;
        RECT 25.950 85.950 28.050 88.050 ;
        RECT 16.950 70.950 19.050 73.050 ;
        RECT 4.950 64.950 7.050 67.050 ;
        RECT 10.950 66.450 13.050 67.050 ;
        RECT 10.950 65.400 15.450 66.450 ;
        RECT 10.950 64.950 13.050 65.400 ;
        RECT 4.950 60.450 7.050 61.200 ;
        RECT 2.400 59.400 7.050 60.450 ;
        RECT 4.950 59.100 7.050 59.400 ;
        RECT 11.400 60.600 12.450 64.950 ;
        RECT 14.400 61.050 15.450 65.400 ;
        RECT 5.400 58.350 6.600 59.100 ;
        RECT 11.400 58.350 12.600 60.600 ;
        RECT 13.950 58.950 16.050 61.050 ;
        RECT 17.400 60.450 18.450 70.950 ;
        RECT 26.400 60.600 27.450 85.950 ;
        RECT 41.400 76.050 42.450 97.800 ;
        RECT 53.400 94.050 54.450 98.400 ;
        RECT 61.950 97.800 64.050 99.900 ;
        RECT 65.400 98.400 66.600 100.650 ;
        RECT 71.400 99.900 72.600 100.650 ;
        RECT 83.400 99.900 84.600 100.650 ;
        RECT 65.400 94.050 66.450 98.400 ;
        RECT 70.950 97.800 73.050 99.900 ;
        RECT 82.950 97.800 85.050 99.900 ;
        RECT 95.400 98.400 96.600 100.650 ;
        RECT 104.400 98.400 105.600 100.650 ;
        RECT 52.950 91.950 55.050 94.050 ;
        RECT 64.950 91.950 67.050 94.050 ;
        RECT 95.400 88.050 96.450 98.400 ;
        RECT 104.400 88.050 105.450 98.400 ;
        RECT 109.800 97.950 111.900 100.050 ;
        RECT 115.800 97.950 117.900 100.050 ;
        RECT 94.950 85.950 97.050 88.050 ;
        RECT 103.950 85.950 106.050 88.050 ;
        RECT 122.400 86.700 123.900 105.600 ;
        RECT 126.300 94.800 127.500 111.300 ;
        RECT 125.400 92.700 127.500 94.800 ;
        RECT 126.300 86.700 127.500 92.700 ;
        RECT 128.700 89.700 129.900 111.300 ;
        RECT 136.800 110.400 138.900 112.500 ;
        RECT 142.200 111.300 144.300 113.400 ;
        RECT 145.200 111.300 147.300 113.400 ;
        RECT 148.200 111.300 150.300 113.400 ;
        RECT 133.800 103.950 135.900 106.050 ;
        RECT 134.400 102.900 135.600 103.650 ;
        RECT 133.950 100.800 136.050 102.900 ;
        RECT 137.400 99.900 138.300 110.400 ;
        RECT 140.100 104.400 142.200 106.500 ;
        RECT 137.400 97.800 139.500 99.900 ;
        RECT 143.100 99.000 144.300 111.300 ;
        RECT 137.400 91.200 138.300 97.800 ;
        RECT 142.800 96.900 144.900 99.000 ;
        RECT 128.700 87.600 130.800 89.700 ;
        RECT 137.400 89.100 139.500 91.200 ;
        RECT 143.100 89.700 144.300 96.900 ;
        RECT 145.800 93.600 147.300 111.300 ;
        RECT 145.800 91.500 147.900 93.600 ;
        RECT 142.800 87.600 144.900 89.700 ;
        RECT 145.800 86.700 147.300 91.500 ;
        RECT 149.100 89.700 150.300 111.300 ;
        RECT 40.950 73.950 43.050 76.050 ;
        RECT 47.400 72.300 50.400 74.400 ;
        RECT 51.300 72.300 53.400 74.400 ;
        RECT 70.200 72.300 72.300 74.400 ;
        RECT 20.400 60.450 21.600 60.600 ;
        RECT 17.400 59.400 21.600 60.450 ;
        RECT 20.400 58.350 21.600 59.400 ;
        RECT 26.400 58.350 27.600 60.600 ;
        RECT 34.800 58.950 36.900 61.050 ;
        RECT 40.800 58.950 42.900 61.050 ;
        RECT 4.950 55.950 7.050 58.050 ;
        RECT 7.950 55.950 10.050 58.050 ;
        RECT 10.950 55.950 13.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 22.950 55.950 25.050 58.050 ;
        RECT 25.950 55.950 28.050 58.050 ;
        RECT 28.950 55.950 31.050 58.050 ;
        RECT 8.400 54.900 9.600 55.650 ;
        RECT 7.950 52.800 10.050 54.900 ;
        RECT 23.400 53.400 24.600 55.650 ;
        RECT 29.400 55.050 30.600 55.650 ;
        RECT 29.400 53.400 34.050 55.050 ;
        RECT 10.950 49.950 13.050 52.050 ;
        RECT 11.400 28.200 12.450 49.950 ;
        RECT 10.950 26.100 13.050 28.200 ;
        RECT 23.400 27.450 24.450 53.400 ;
        RECT 30.000 52.950 34.050 53.400 ;
        RECT 47.400 53.400 48.900 72.300 ;
        RECT 51.300 66.300 52.500 72.300 ;
        RECT 50.400 64.200 52.500 66.300 ;
        RECT 47.400 51.300 49.500 53.400 ;
        RECT 48.300 47.700 49.500 51.300 ;
        RECT 51.300 47.700 52.500 64.200 ;
        RECT 53.700 69.300 55.800 71.400 ;
        RECT 53.700 47.700 54.900 69.300 ;
        RECT 62.400 67.800 64.500 69.900 ;
        RECT 67.800 69.300 69.900 71.400 ;
        RECT 58.950 61.950 61.050 64.050 ;
        RECT 59.400 57.600 60.450 61.950 ;
        RECT 62.400 61.200 63.300 67.800 ;
        RECT 68.100 62.100 69.300 69.300 ;
        RECT 70.800 67.500 72.300 72.300 ;
        RECT 73.200 69.300 75.300 74.400 ;
        RECT 70.800 65.400 72.900 67.500 ;
        RECT 62.400 59.100 64.500 61.200 ;
        RECT 67.800 60.000 69.900 62.100 ;
        RECT 59.400 55.350 60.600 57.600 ;
        RECT 58.800 52.950 60.900 55.050 ;
        RECT 62.400 48.600 63.300 59.100 ;
        RECT 65.100 52.500 67.200 54.600 ;
        RECT 47.700 45.600 49.800 47.700 ;
        RECT 50.700 45.600 52.800 47.700 ;
        RECT 53.700 45.600 55.800 47.700 ;
        RECT 61.800 46.500 63.900 48.600 ;
        RECT 68.100 47.700 69.300 60.000 ;
        RECT 70.800 47.700 72.300 65.400 ;
        RECT 74.100 47.700 75.300 69.300 ;
        RECT 67.200 45.600 69.300 47.700 ;
        RECT 70.200 45.600 72.300 47.700 ;
        RECT 73.200 45.600 75.300 47.700 ;
        RECT 76.200 72.300 78.300 74.400 ;
        RECT 76.200 67.500 77.700 72.300 ;
        RECT 97.950 67.950 100.050 70.050 ;
        RECT 76.200 65.400 78.300 67.500 ;
        RECT 76.200 47.700 77.700 65.400 ;
        RECT 79.950 61.950 82.050 64.050 ;
        RECT 76.200 45.600 78.300 47.700 ;
        RECT 80.400 40.050 81.450 61.950 ;
        RECT 85.800 58.950 87.900 61.050 ;
        RECT 94.800 58.950 96.900 61.050 ;
        RECT 82.950 55.950 85.050 58.050 ;
        RECT 95.400 56.400 96.600 58.650 ;
        RECT 79.950 37.950 82.050 40.050 ;
        RECT 29.700 33.300 31.800 35.400 ;
        RECT 32.700 33.300 34.800 35.400 ;
        RECT 35.700 33.300 37.800 35.400 ;
        RECT 30.300 29.700 31.500 33.300 ;
        RECT 29.400 27.600 31.500 29.700 ;
        RECT 23.400 27.000 27.450 27.450 ;
        RECT 23.400 26.400 28.050 27.000 ;
        RECT 11.400 25.350 12.600 26.100 ;
        RECT 5.100 22.950 7.200 25.050 ;
        RECT 10.500 22.950 12.600 25.050 ;
        RECT 25.950 22.950 28.050 26.400 ;
        RECT 16.800 19.950 18.900 22.050 ;
        RECT 22.800 19.950 24.900 22.050 ;
        RECT 29.400 8.700 30.900 27.600 ;
        RECT 33.300 16.800 34.500 33.300 ;
        RECT 32.400 14.700 34.500 16.800 ;
        RECT 33.300 8.700 34.500 14.700 ;
        RECT 35.700 11.700 36.900 33.300 ;
        RECT 43.800 32.400 45.900 34.500 ;
        RECT 49.200 33.300 51.300 35.400 ;
        RECT 52.200 33.300 54.300 35.400 ;
        RECT 55.200 33.300 57.300 35.400 ;
        RECT 40.800 25.950 42.900 28.050 ;
        RECT 41.400 24.900 42.600 25.650 ;
        RECT 40.950 22.800 43.050 24.900 ;
        RECT 44.400 21.900 45.300 32.400 ;
        RECT 47.100 26.400 49.200 28.500 ;
        RECT 44.400 19.800 46.500 21.900 ;
        RECT 50.100 21.000 51.300 33.300 ;
        RECT 44.400 13.200 45.300 19.800 ;
        RECT 49.800 18.900 51.900 21.000 ;
        RECT 35.700 9.600 37.800 11.700 ;
        RECT 44.400 11.100 46.500 13.200 ;
        RECT 50.100 11.700 51.300 18.900 ;
        RECT 52.800 15.600 54.300 33.300 ;
        RECT 52.800 13.500 54.900 15.600 ;
        RECT 49.800 9.600 51.900 11.700 ;
        RECT 52.800 8.700 54.300 13.500 ;
        RECT 56.100 11.700 57.300 33.300 ;
        RECT 29.400 6.600 32.400 8.700 ;
        RECT 33.300 6.600 35.400 8.700 ;
        RECT 52.200 6.600 54.300 8.700 ;
        RECT 55.200 6.600 57.300 11.700 ;
        RECT 58.200 33.300 60.300 35.400 ;
        RECT 58.200 15.600 59.700 33.300 ;
        RECT 76.950 24.000 79.050 28.050 ;
        RECT 77.400 22.350 78.600 24.000 ;
        RECT 67.800 19.950 69.900 22.050 ;
        RECT 76.800 19.950 78.900 22.050 ;
        RECT 83.400 19.050 84.450 55.950 ;
        RECT 95.400 28.200 96.450 56.400 ;
        RECT 98.400 54.900 99.450 67.950 ;
        RECT 104.400 67.050 105.450 85.950 ;
        RECT 122.400 84.600 125.400 86.700 ;
        RECT 126.300 84.600 128.400 86.700 ;
        RECT 145.200 84.600 147.300 86.700 ;
        RECT 148.200 84.600 150.300 89.700 ;
        RECT 151.200 111.300 153.300 113.400 ;
        RECT 154.950 112.950 157.050 115.050 ;
        RECT 151.200 93.600 152.700 111.300 ;
        RECT 151.200 91.500 153.300 93.600 ;
        RECT 151.200 86.700 152.700 91.500 ;
        RECT 151.200 84.600 153.300 86.700 ;
        RECT 155.400 82.050 156.450 112.950 ;
        RECT 158.400 102.900 159.450 118.950 ;
        RECT 164.400 106.050 165.450 130.950 ;
        RECT 166.950 127.950 169.050 132.000 ;
        RECT 179.400 131.400 180.600 133.650 ;
        RECT 179.400 127.050 180.450 131.400 ;
        RECT 178.950 124.950 181.050 127.050 ;
        RECT 184.950 118.950 187.050 121.050 ;
        RECT 169.950 114.450 172.050 115.050 ;
        RECT 169.950 113.400 177.450 114.450 ;
        RECT 169.950 112.950 172.050 113.400 ;
        RECT 172.950 109.950 175.050 112.050 ;
        RECT 169.950 106.950 172.050 109.050 ;
        RECT 163.950 103.950 166.050 106.050 ;
        RECT 170.400 103.200 171.450 106.950 ;
        RECT 157.950 100.800 160.050 102.900 ;
        RECT 163.950 100.800 166.050 102.900 ;
        RECT 169.950 101.100 172.050 103.200 ;
        RECT 160.800 97.950 162.900 100.050 ;
        RECT 145.950 79.950 148.050 82.050 ;
        RECT 154.950 79.950 157.050 82.050 ;
        RECT 121.950 70.950 124.050 73.050 ;
        RECT 103.800 64.950 105.900 67.050 ;
        RECT 106.950 63.450 109.050 67.050 ;
        RECT 115.950 64.950 118.050 67.050 ;
        RECT 104.400 63.000 109.050 63.450 ;
        RECT 104.400 62.400 108.450 63.000 ;
        RECT 104.400 60.600 105.450 62.400 ;
        RECT 104.400 58.350 105.600 60.600 ;
        RECT 109.950 59.100 112.050 61.200 ;
        RECT 116.400 61.050 117.450 64.950 ;
        RECT 110.400 58.350 111.600 59.100 ;
        RECT 115.950 58.950 118.050 61.050 ;
        RECT 122.400 60.600 123.450 70.950 ;
        RECT 127.950 67.950 130.050 70.050 ;
        RECT 128.400 60.600 129.450 67.950 ;
        RECT 146.400 60.600 147.450 79.950 ;
        RECT 148.950 76.950 151.050 79.050 ;
        RECT 149.400 61.050 150.450 76.950 ;
        RECT 157.950 70.950 160.050 73.050 ;
        RECT 158.400 64.050 159.450 70.950 ;
        RECT 160.950 64.950 163.050 67.050 ;
        RECT 157.950 61.950 160.050 64.050 ;
        RECT 122.400 58.350 123.600 60.600 ;
        RECT 128.400 58.350 129.600 60.600 ;
        RECT 137.400 60.450 138.600 60.600 ;
        RECT 134.400 59.400 138.600 60.450 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 112.950 55.950 115.050 58.050 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 97.950 52.800 100.050 54.900 ;
        RECT 107.400 53.400 108.600 55.650 ;
        RECT 113.400 54.900 114.600 55.650 ;
        RECT 107.400 40.050 108.450 53.400 ;
        RECT 112.800 52.800 114.900 54.900 ;
        RECT 115.950 52.950 118.050 55.050 ;
        RECT 125.400 54.900 126.600 55.650 ;
        RECT 106.950 37.950 109.050 40.050 ;
        RECT 109.950 34.950 112.050 37.050 ;
        RECT 110.400 28.200 111.450 34.950 ;
        RECT 116.400 34.050 117.450 52.950 ;
        RECT 124.950 52.800 127.050 54.900 ;
        RECT 130.950 52.950 133.050 55.050 ;
        RECT 127.950 49.950 130.050 52.050 ;
        RECT 128.400 37.050 129.450 49.950 ;
        RECT 131.400 40.050 132.450 52.950 ;
        RECT 134.400 49.050 135.450 59.400 ;
        RECT 137.400 58.350 138.600 59.400 ;
        RECT 146.400 58.350 147.600 60.600 ;
        RECT 148.950 58.950 151.050 61.050 ;
        RECT 154.950 59.100 157.050 61.200 ;
        RECT 161.400 60.600 162.450 64.950 ;
        RECT 164.400 61.050 165.450 100.800 ;
        RECT 170.400 100.350 171.600 101.100 ;
        RECT 169.800 97.950 171.900 100.050 ;
        RECT 173.400 63.450 174.450 109.950 ;
        RECT 176.400 105.450 177.450 113.400 ;
        RECT 185.400 105.600 186.450 118.950 ;
        RECT 188.400 108.450 189.450 172.950 ;
        RECT 209.400 164.700 210.900 183.600 ;
        RECT 213.300 172.800 214.500 189.300 ;
        RECT 212.400 170.700 214.500 172.800 ;
        RECT 213.300 164.700 214.500 170.700 ;
        RECT 215.700 167.700 216.900 189.300 ;
        RECT 223.800 188.400 225.900 190.500 ;
        RECT 229.200 189.300 231.300 191.400 ;
        RECT 232.200 189.300 234.300 191.400 ;
        RECT 235.200 189.300 237.300 191.400 ;
        RECT 220.800 181.950 222.900 184.050 ;
        RECT 221.400 180.900 222.600 181.650 ;
        RECT 220.950 178.800 223.050 180.900 ;
        RECT 224.400 177.900 225.300 188.400 ;
        RECT 227.100 182.400 229.200 184.500 ;
        RECT 224.400 175.800 226.500 177.900 ;
        RECT 230.100 177.000 231.300 189.300 ;
        RECT 224.400 169.200 225.300 175.800 ;
        RECT 229.800 174.900 231.900 177.000 ;
        RECT 215.700 165.600 217.800 167.700 ;
        RECT 224.400 167.100 226.500 169.200 ;
        RECT 230.100 167.700 231.300 174.900 ;
        RECT 232.800 171.600 234.300 189.300 ;
        RECT 232.800 169.500 234.900 171.600 ;
        RECT 229.800 165.600 231.900 167.700 ;
        RECT 232.800 164.700 234.300 169.500 ;
        RECT 236.100 167.700 237.300 189.300 ;
        RECT 209.400 162.600 212.400 164.700 ;
        RECT 213.300 162.600 215.400 164.700 ;
        RECT 232.200 162.600 234.300 164.700 ;
        RECT 235.200 162.600 237.300 167.700 ;
        RECT 238.200 189.300 240.300 191.400 ;
        RECT 238.200 171.600 239.700 189.300 ;
        RECT 257.400 180.600 258.450 205.950 ;
        RECT 260.400 198.450 261.450 209.400 ;
        RECT 265.950 208.950 268.050 211.050 ;
        RECT 269.400 209.400 270.600 211.650 ;
        RECT 275.400 209.400 276.600 211.650 ;
        RECT 260.400 197.400 264.450 198.450 ;
        RECT 263.400 187.050 264.450 197.400 ;
        RECT 266.400 190.050 267.450 208.950 ;
        RECT 269.400 199.050 270.450 209.400 ;
        RECT 275.400 202.050 276.450 209.400 ;
        RECT 283.950 208.950 286.050 211.050 ;
        RECT 287.400 209.400 288.600 211.650 ;
        RECT 293.400 210.900 294.600 211.650 ;
        RECT 305.400 210.900 306.600 211.650 ;
        RECT 314.400 210.900 315.600 211.650 ;
        RECT 280.950 205.950 283.050 208.050 ;
        RECT 281.400 202.050 282.450 205.950 ;
        RECT 274.950 199.950 277.050 202.050 ;
        RECT 280.950 199.950 283.050 202.050 ;
        RECT 284.400 199.050 285.450 208.950 ;
        RECT 268.950 196.950 271.050 199.050 ;
        RECT 283.950 196.950 286.050 199.050 ;
        RECT 265.950 187.950 268.050 190.050 ;
        RECT 277.950 187.950 280.050 190.050 ;
        RECT 262.950 184.950 265.050 187.050 ;
        RECT 268.950 183.000 271.050 187.050 ;
        RECT 269.400 181.350 270.600 183.000 ;
        RECT 257.400 178.350 258.600 180.600 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 268.950 178.950 271.050 181.050 ;
        RECT 271.950 178.950 274.050 181.050 ;
        RECT 247.800 175.950 249.900 178.050 ;
        RECT 256.800 175.950 258.900 178.050 ;
        RECT 272.400 177.900 273.600 178.650 ;
        RECT 278.400 177.900 279.450 187.950 ;
        RECT 287.400 184.050 288.450 209.400 ;
        RECT 292.950 208.800 295.050 210.900 ;
        RECT 304.950 208.800 307.050 210.900 ;
        RECT 313.950 208.800 316.050 210.900 ;
        RECT 326.400 209.400 327.600 211.650 ;
        RECT 332.400 209.400 333.600 211.650 ;
        RECT 344.400 210.900 345.600 211.650 ;
        RECT 301.950 205.950 304.050 208.050 ;
        RECT 292.950 193.950 295.050 196.050 ;
        RECT 286.950 181.950 289.050 184.050 ;
        RECT 293.400 183.600 294.450 193.950 ;
        RECT 302.400 193.050 303.450 205.950 ;
        RECT 314.400 202.050 315.450 208.800 ;
        RECT 304.950 199.950 307.050 202.050 ;
        RECT 313.950 199.950 316.050 202.050 ;
        RECT 301.950 190.950 304.050 193.050 ;
        RECT 305.400 190.050 306.450 199.950 ;
        RECT 326.400 199.050 327.450 209.400 ;
        RECT 328.950 205.950 331.050 208.050 ;
        RECT 325.950 196.950 328.050 199.050 ;
        RECT 304.950 187.950 307.050 190.050 ;
        RECT 329.400 184.200 330.450 205.950 ;
        RECT 332.400 196.050 333.450 209.400 ;
        RECT 343.950 208.800 346.050 210.900 ;
        RECT 350.400 209.400 351.600 211.650 ;
        RECT 356.400 210.900 357.600 211.650 ;
        RECT 346.950 199.950 349.050 202.050 ;
        RECT 331.950 193.950 334.050 196.050 ;
        RECT 332.400 187.050 333.450 193.950 ;
        RECT 340.950 187.950 343.050 190.050 ;
        RECT 331.950 184.950 334.050 187.050 ;
        RECT 293.400 181.350 294.600 183.600 ;
        RECT 298.950 182.100 301.050 184.200 ;
        RECT 304.950 182.100 307.050 184.200 ;
        RECT 319.950 182.100 322.050 184.200 ;
        RECT 328.950 182.100 331.050 184.200 ;
        RECT 341.400 183.600 342.450 187.950 ;
        RECT 347.400 186.450 348.450 199.950 ;
        RECT 350.400 193.050 351.450 209.400 ;
        RECT 355.950 208.800 358.050 210.900 ;
        RECT 349.950 190.950 352.050 193.050 ;
        RECT 356.400 186.450 357.450 208.800 ;
        RECT 347.400 185.400 351.450 186.450 ;
        RECT 299.400 181.350 300.600 182.100 ;
        RECT 305.400 181.350 306.600 182.100 ;
        RECT 320.400 181.350 321.600 182.100 ;
        RECT 329.400 181.350 330.600 182.100 ;
        RECT 341.400 181.350 342.600 183.600 ;
        RECT 281.100 178.950 283.200 181.050 ;
        RECT 284.100 178.950 286.200 181.050 ;
        RECT 289.800 178.950 291.900 181.050 ;
        RECT 292.800 178.950 294.900 181.050 ;
        RECT 298.950 178.950 301.050 181.050 ;
        RECT 301.950 178.950 304.050 181.050 ;
        RECT 304.950 178.950 307.050 181.050 ;
        RECT 307.950 178.950 310.050 181.050 ;
        RECT 316.950 178.950 319.050 181.050 ;
        RECT 319.950 178.950 322.050 181.050 ;
        RECT 322.950 178.950 325.050 181.050 ;
        RECT 328.950 178.950 331.050 181.050 ;
        RECT 331.950 178.950 334.050 181.050 ;
        RECT 341.400 178.950 343.500 181.050 ;
        RECT 346.800 178.950 348.900 181.050 ;
        RECT 271.950 175.800 274.050 177.900 ;
        RECT 277.950 177.450 280.050 177.900 ;
        RECT 275.400 176.400 280.050 177.450 ;
        RECT 238.200 169.500 240.300 171.600 ;
        RECT 238.200 164.700 239.700 169.500 ;
        RECT 271.950 166.950 274.050 169.050 ;
        RECT 238.200 162.600 240.300 164.700 ;
        RECT 265.950 160.950 268.050 163.050 ;
        RECT 223.950 154.950 226.050 157.050 ;
        RECT 232.950 154.950 235.050 157.050 ;
        RECT 202.950 142.950 205.050 145.050 ;
        RECT 208.950 142.950 211.050 145.050 ;
        RECT 190.950 137.100 193.050 139.200 ;
        RECT 199.950 137.100 202.050 139.200 ;
        RECT 191.400 136.350 192.600 137.100 ;
        RECT 200.400 136.350 201.600 137.100 ;
        RECT 191.100 133.950 193.200 136.050 ;
        RECT 194.400 133.950 196.500 136.050 ;
        RECT 199.800 133.950 201.900 136.050 ;
        RECT 194.400 131.400 195.600 133.650 ;
        RECT 194.400 127.050 195.450 131.400 ;
        RECT 193.950 124.950 196.050 127.050 ;
        RECT 203.400 112.050 204.450 142.950 ;
        RECT 209.400 138.600 210.450 142.950 ;
        RECT 224.400 138.600 225.450 154.950 ;
        RECT 233.400 139.050 234.450 154.950 ;
        RECT 241.950 151.950 244.050 154.050 ;
        RECT 242.400 148.050 243.450 151.950 ;
        RECT 241.950 145.950 244.050 148.050 ;
        RECT 253.950 142.950 256.050 145.050 ;
        RECT 254.400 139.200 255.450 142.950 ;
        RECT 266.400 139.200 267.450 160.950 ;
        RECT 209.400 136.350 210.600 138.600 ;
        RECT 224.400 136.350 225.600 138.600 ;
        RECT 232.950 136.950 235.050 139.050 ;
        RECT 241.950 137.100 244.050 139.200 ;
        RECT 253.950 137.100 256.050 139.200 ;
        RECT 265.950 137.100 268.050 139.200 ;
        RECT 272.400 138.600 273.450 166.950 ;
        RECT 275.400 145.050 276.450 176.400 ;
        RECT 277.950 175.800 280.050 176.400 ;
        RECT 281.400 176.400 282.600 178.650 ;
        RECT 277.950 154.950 280.050 157.050 ;
        RECT 274.950 142.950 277.050 145.050 ;
        RECT 278.400 138.600 279.450 154.950 ;
        RECT 281.400 148.050 282.450 176.400 ;
        RECT 286.950 175.950 289.050 178.050 ;
        RECT 290.400 176.400 291.600 178.650 ;
        RECT 302.400 177.000 303.600 178.650 ;
        RECT 308.400 177.900 309.600 178.650 ;
        RECT 280.950 145.950 283.050 148.050 ;
        RECT 287.400 141.450 288.450 175.950 ;
        RECT 290.400 175.050 291.450 176.400 ;
        RECT 290.400 173.400 295.050 175.050 ;
        RECT 291.000 172.950 295.050 173.400 ;
        RECT 301.950 172.950 304.050 177.000 ;
        RECT 307.950 175.800 310.050 177.900 ;
        RECT 317.400 176.400 318.600 178.650 ;
        RECT 323.400 177.900 324.600 178.650 ;
        RECT 332.400 177.900 333.600 178.650 ;
        RECT 317.400 172.050 318.450 176.400 ;
        RECT 322.950 175.800 325.050 177.900 ;
        RECT 331.950 175.800 334.050 177.900 ;
        RECT 298.950 169.950 301.050 172.050 ;
        RECT 316.950 169.950 319.050 172.050 ;
        RECT 295.950 166.950 298.050 169.050 ;
        RECT 296.400 145.050 297.450 166.950 ;
        RECT 295.950 142.950 298.050 145.050 ;
        RECT 299.400 144.450 300.450 169.950 ;
        RECT 317.400 163.050 318.450 169.950 ;
        RECT 316.950 160.950 319.050 163.050 ;
        RECT 323.400 157.050 324.450 175.800 ;
        RECT 322.950 154.950 325.050 157.050 ;
        RECT 346.950 154.950 349.050 157.050 ;
        RECT 305.400 150.300 308.400 152.400 ;
        RECT 309.300 150.300 311.400 152.400 ;
        RECT 328.200 150.300 330.300 152.400 ;
        RECT 299.400 143.400 303.450 144.450 ;
        RECT 284.400 140.400 288.450 141.450 ;
        RECT 284.400 138.600 285.450 140.400 ;
        RECT 242.400 136.350 243.600 137.100 ;
        RECT 254.400 136.350 255.600 137.100 ;
        RECT 266.400 136.350 267.600 137.100 ;
        RECT 272.400 136.350 273.600 138.600 ;
        RECT 278.400 136.350 279.600 138.600 ;
        RECT 284.400 136.350 285.600 138.600 ;
        RECT 292.800 136.950 294.900 139.050 ;
        RECT 298.800 136.950 300.900 139.050 ;
        RECT 208.950 133.950 211.050 136.050 ;
        RECT 211.950 133.950 214.050 136.050 ;
        RECT 214.950 133.950 217.050 136.050 ;
        RECT 224.100 133.950 226.200 136.050 ;
        RECT 229.500 133.950 231.600 136.050 ;
        RECT 235.950 133.950 238.050 136.050 ;
        RECT 238.950 133.950 241.050 136.050 ;
        RECT 241.950 133.950 244.050 136.050 ;
        RECT 247.950 133.950 250.050 136.050 ;
        RECT 250.950 133.950 253.050 136.050 ;
        RECT 253.950 133.950 256.050 136.050 ;
        RECT 256.950 133.950 259.050 136.050 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 268.950 133.950 271.050 136.050 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 277.950 133.950 280.050 136.050 ;
        RECT 280.950 133.950 283.050 136.050 ;
        RECT 283.950 133.950 286.050 136.050 ;
        RECT 286.950 133.950 289.050 136.050 ;
        RECT 205.950 130.950 208.050 133.050 ;
        RECT 212.400 131.400 213.600 133.650 ;
        RECT 239.400 132.900 240.600 133.650 ;
        RECT 257.400 132.900 258.600 133.650 ;
        RECT 269.400 132.900 270.600 133.650 ;
        RECT 281.400 132.900 282.600 133.650 ;
        RECT 287.400 132.900 288.600 133.650 ;
        RECT 202.950 109.950 205.050 112.050 ;
        RECT 188.400 108.000 192.450 108.450 ;
        RECT 188.400 107.400 193.050 108.000 ;
        RECT 179.400 105.450 180.600 105.600 ;
        RECT 176.400 104.400 180.600 105.450 ;
        RECT 179.400 103.350 180.600 104.400 ;
        RECT 185.400 103.350 186.600 105.600 ;
        RECT 190.950 103.950 193.050 107.400 ;
        RECT 199.950 105.000 202.050 109.050 ;
        RECT 206.400 105.600 207.450 130.950 ;
        RECT 212.400 109.050 213.450 131.400 ;
        RECT 238.950 130.800 241.050 132.900 ;
        RECT 256.950 130.800 259.050 132.900 ;
        RECT 268.950 130.800 271.050 132.900 ;
        RECT 280.950 130.800 283.050 132.900 ;
        RECT 286.950 130.800 289.050 132.900 ;
        RECT 302.400 118.050 303.450 143.400 ;
        RECT 305.400 131.400 306.900 150.300 ;
        RECT 309.300 144.300 310.500 150.300 ;
        RECT 308.400 142.200 310.500 144.300 ;
        RECT 305.400 129.300 307.500 131.400 ;
        RECT 306.300 125.700 307.500 129.300 ;
        RECT 309.300 125.700 310.500 142.200 ;
        RECT 311.700 147.300 313.800 149.400 ;
        RECT 311.700 125.700 312.900 147.300 ;
        RECT 320.400 145.800 322.500 147.900 ;
        RECT 325.800 147.300 327.900 149.400 ;
        RECT 320.400 139.200 321.300 145.800 ;
        RECT 326.100 140.100 327.300 147.300 ;
        RECT 328.800 145.500 330.300 150.300 ;
        RECT 331.200 147.300 333.300 152.400 ;
        RECT 328.800 143.400 330.900 145.500 ;
        RECT 320.400 137.100 322.500 139.200 ;
        RECT 325.800 138.000 327.900 140.100 ;
        RECT 316.950 134.100 319.050 136.200 ;
        RECT 317.400 133.350 318.600 134.100 ;
        RECT 316.800 130.950 318.900 133.050 ;
        RECT 320.400 126.600 321.300 137.100 ;
        RECT 323.100 130.500 325.200 132.600 ;
        RECT 305.700 123.600 307.800 125.700 ;
        RECT 308.700 123.600 310.800 125.700 ;
        RECT 311.700 123.600 313.800 125.700 ;
        RECT 319.800 124.500 321.900 126.600 ;
        RECT 326.100 125.700 327.300 138.000 ;
        RECT 328.800 125.700 330.300 143.400 ;
        RECT 332.100 125.700 333.300 147.300 ;
        RECT 325.200 123.600 327.300 125.700 ;
        RECT 328.200 123.600 330.300 125.700 ;
        RECT 331.200 123.600 333.300 125.700 ;
        RECT 334.200 150.300 336.300 152.400 ;
        RECT 334.200 145.500 335.700 150.300 ;
        RECT 334.200 143.400 336.300 145.500 ;
        RECT 334.200 125.700 335.700 143.400 ;
        RECT 343.800 136.950 345.900 139.050 ;
        RECT 334.200 123.600 336.300 125.700 ;
        RECT 301.950 115.950 304.050 118.050 ;
        RECT 310.950 115.950 313.050 118.050 ;
        RECT 250.950 109.950 253.050 112.050 ;
        RECT 278.700 111.300 280.800 113.400 ;
        RECT 281.700 111.300 283.800 113.400 ;
        RECT 284.700 111.300 286.800 113.400 ;
        RECT 211.950 106.950 214.050 109.050 ;
        RECT 200.400 103.350 201.600 105.000 ;
        RECT 206.400 103.350 207.600 105.600 ;
        RECT 214.950 104.100 217.050 106.200 ;
        RECT 229.950 104.100 232.050 106.200 ;
        RECT 251.400 105.600 252.450 109.950 ;
        RECT 279.300 107.700 280.500 111.300 ;
        RECT 215.400 103.350 216.600 104.100 ;
        RECT 230.400 103.350 231.600 104.100 ;
        RECT 251.400 103.350 252.600 105.600 ;
        RECT 256.950 104.100 259.050 106.200 ;
        RECT 278.400 105.600 280.500 107.700 ;
        RECT 257.400 103.350 258.600 104.100 ;
        RECT 178.950 100.950 181.050 103.050 ;
        RECT 181.950 100.950 184.050 103.050 ;
        RECT 184.950 100.950 187.050 103.050 ;
        RECT 187.950 100.950 190.050 103.050 ;
        RECT 196.950 100.950 199.050 103.050 ;
        RECT 199.950 100.950 202.050 103.050 ;
        RECT 202.950 100.950 205.050 103.050 ;
        RECT 205.950 100.950 208.050 103.050 ;
        RECT 211.950 100.950 214.050 103.050 ;
        RECT 214.950 100.950 217.050 103.050 ;
        RECT 217.950 100.950 220.050 103.050 ;
        RECT 226.950 100.950 229.050 103.050 ;
        RECT 229.950 100.950 232.050 103.050 ;
        RECT 232.950 100.950 235.050 103.050 ;
        RECT 239.100 100.950 241.200 103.050 ;
        RECT 244.500 100.950 246.600 103.050 ;
        RECT 250.950 100.950 253.050 103.050 ;
        RECT 253.950 100.950 256.050 103.050 ;
        RECT 256.950 100.950 259.050 103.050 ;
        RECT 259.950 100.950 262.050 103.050 ;
        RECT 182.400 98.400 183.600 100.650 ;
        RECT 188.400 99.900 189.600 100.650 ;
        RECT 175.950 91.950 178.050 94.050 ;
        RECT 170.400 62.400 174.450 63.450 ;
        RECT 155.400 58.350 156.600 59.100 ;
        RECT 161.400 58.350 162.600 60.600 ;
        RECT 163.950 58.950 166.050 61.050 ;
        RECT 170.400 60.600 171.450 62.400 ;
        RECT 176.400 60.600 177.450 91.950 ;
        RECT 182.400 79.050 183.450 98.400 ;
        RECT 187.950 97.800 190.050 99.900 ;
        RECT 193.950 97.950 196.050 100.050 ;
        RECT 197.400 98.400 198.600 100.650 ;
        RECT 203.400 99.000 204.600 100.650 ;
        RECT 194.400 94.050 195.450 97.950 ;
        RECT 193.950 91.950 196.050 94.050 ;
        RECT 197.400 88.050 198.450 98.400 ;
        RECT 202.950 94.950 205.050 99.000 ;
        RECT 208.950 97.950 211.050 100.050 ;
        RECT 218.400 98.400 219.600 100.650 ;
        RECT 227.400 99.900 228.600 100.650 ;
        RECT 196.950 85.950 199.050 88.050 ;
        RECT 197.400 79.050 198.450 85.950 ;
        RECT 181.950 76.950 184.050 79.050 ;
        RECT 196.950 76.950 199.050 79.050 ;
        RECT 178.950 67.950 181.050 70.050 ;
        RECT 184.950 67.950 187.050 70.050 ;
        RECT 205.950 67.950 208.050 70.050 ;
        RECT 179.400 61.200 180.450 67.950 ;
        RECT 170.400 58.350 171.600 60.600 ;
        RECT 176.400 58.350 177.600 60.600 ;
        RECT 178.950 59.100 181.050 61.200 ;
        RECT 185.400 60.600 186.450 67.950 ;
        RECT 187.950 64.950 190.050 67.050 ;
        RECT 188.400 61.050 189.450 64.950 ;
        RECT 179.400 58.350 180.600 59.100 ;
        RECT 185.400 58.350 186.600 60.600 ;
        RECT 187.950 58.950 190.050 61.050 ;
        RECT 193.950 59.100 196.050 61.200 ;
        RECT 199.950 59.100 202.050 61.200 ;
        RECT 206.400 61.050 207.450 67.950 ;
        RECT 194.400 58.350 195.600 59.100 ;
        RECT 200.400 58.350 201.600 59.100 ;
        RECT 205.950 58.950 208.050 61.050 ;
        RECT 209.400 60.600 210.450 97.950 ;
        RECT 218.400 94.050 219.450 98.400 ;
        RECT 226.950 97.800 229.050 99.900 ;
        RECT 233.400 98.400 234.600 100.650 ;
        RECT 217.950 91.950 220.050 94.050 ;
        RECT 229.950 91.950 232.050 94.050 ;
        RECT 218.400 71.400 228.450 72.450 ;
        RECT 218.400 67.050 219.450 71.400 ;
        RECT 220.950 67.950 223.050 70.050 ;
        RECT 217.950 64.950 220.050 67.050 ;
        RECT 209.400 58.350 210.600 60.600 ;
        RECT 214.950 59.100 217.050 61.200 ;
        RECT 221.400 61.050 222.450 67.950 ;
        RECT 215.400 58.350 216.600 59.100 ;
        RECT 220.950 58.950 223.050 61.050 ;
        RECT 227.400 60.600 228.450 71.400 ;
        RECT 230.400 64.050 231.450 91.950 ;
        RECT 233.400 88.050 234.450 98.400 ;
        RECT 235.950 97.950 238.050 100.050 ;
        RECT 239.400 98.400 240.600 100.650 ;
        RECT 236.400 94.050 237.450 97.950 ;
        RECT 235.950 91.950 238.050 94.050 ;
        RECT 239.400 88.050 240.450 98.400 ;
        RECT 247.950 97.950 250.050 100.050 ;
        RECT 254.400 98.400 255.600 100.650 ;
        RECT 260.400 98.400 261.600 100.650 ;
        RECT 232.950 85.950 235.050 88.050 ;
        RECT 238.950 85.950 241.050 88.050 ;
        RECT 233.400 79.050 234.450 85.950 ;
        RECT 232.950 76.950 235.050 79.050 ;
        RECT 229.950 61.950 232.050 64.050 ;
        RECT 233.400 61.050 234.450 76.950 ;
        RECT 244.950 67.950 247.050 70.050 ;
        RECT 245.400 63.450 246.450 67.950 ;
        RECT 248.400 67.050 249.450 97.950 ;
        RECT 254.400 91.050 255.450 98.400 ;
        RECT 260.400 94.050 261.450 98.400 ;
        RECT 265.800 97.950 267.900 100.050 ;
        RECT 271.800 97.950 273.900 100.050 ;
        RECT 259.950 91.950 262.050 94.050 ;
        RECT 253.950 88.950 256.050 91.050 ;
        RECT 259.950 88.800 262.050 90.900 ;
        RECT 260.400 73.050 261.450 88.800 ;
        RECT 278.400 86.700 279.900 105.600 ;
        RECT 282.300 94.800 283.500 111.300 ;
        RECT 281.400 92.700 283.500 94.800 ;
        RECT 282.300 86.700 283.500 92.700 ;
        RECT 284.700 89.700 285.900 111.300 ;
        RECT 292.800 110.400 294.900 112.500 ;
        RECT 298.200 111.300 300.300 113.400 ;
        RECT 301.200 111.300 303.300 113.400 ;
        RECT 304.200 111.300 306.300 113.400 ;
        RECT 289.800 103.950 291.900 106.050 ;
        RECT 290.400 102.900 291.600 103.650 ;
        RECT 289.950 100.800 292.050 102.900 ;
        RECT 293.400 99.900 294.300 110.400 ;
        RECT 296.100 104.400 298.200 106.500 ;
        RECT 293.400 97.800 295.500 99.900 ;
        RECT 299.100 99.000 300.300 111.300 ;
        RECT 293.400 91.200 294.300 97.800 ;
        RECT 298.800 96.900 300.900 99.000 ;
        RECT 284.700 87.600 286.800 89.700 ;
        RECT 293.400 89.100 295.500 91.200 ;
        RECT 299.100 89.700 300.300 96.900 ;
        RECT 301.800 93.600 303.300 111.300 ;
        RECT 301.800 91.500 303.900 93.600 ;
        RECT 298.800 87.600 300.900 89.700 ;
        RECT 301.800 86.700 303.300 91.500 ;
        RECT 305.100 89.700 306.300 111.300 ;
        RECT 278.400 84.600 281.400 86.700 ;
        RECT 282.300 84.600 284.400 86.700 ;
        RECT 301.200 84.600 303.300 86.700 ;
        RECT 304.200 84.600 306.300 89.700 ;
        RECT 307.200 111.300 309.300 113.400 ;
        RECT 307.200 93.600 308.700 111.300 ;
        RECT 311.400 102.900 312.450 115.950 ;
        RECT 347.400 115.050 348.450 154.950 ;
        RECT 350.400 142.050 351.450 185.400 ;
        RECT 353.400 185.400 357.450 186.450 ;
        RECT 353.400 183.600 354.450 185.400 ;
        RECT 353.400 181.350 354.600 183.600 ;
        RECT 353.400 178.950 355.500 181.050 ;
        RECT 358.800 178.950 360.900 181.050 ;
        RECT 349.950 139.950 352.050 142.050 ;
        RECT 355.950 139.950 358.050 142.050 ;
        RECT 352.800 136.950 354.900 139.050 ;
        RECT 353.400 135.450 354.600 136.650 ;
        RECT 356.400 135.450 357.450 139.950 ;
        RECT 353.400 134.400 357.450 135.450 ;
        RECT 325.950 112.950 328.050 115.050 ;
        RECT 337.950 112.950 340.050 115.050 ;
        RECT 346.950 112.950 349.050 115.050 ;
        RECT 310.950 100.800 313.050 102.900 ;
        RECT 326.400 102.600 327.450 112.950 ;
        RECT 338.400 105.600 339.450 112.950 ;
        RECT 353.400 105.600 354.450 134.400 ;
        RECT 338.400 103.350 339.600 105.600 ;
        RECT 353.400 103.350 354.600 105.600 ;
        RECT 326.400 100.350 327.600 102.600 ;
        RECT 338.400 100.950 340.500 103.050 ;
        RECT 343.800 100.950 345.900 103.050 ;
        RECT 353.400 100.950 355.500 103.050 ;
        RECT 358.800 100.950 360.900 103.050 ;
        RECT 316.800 97.950 318.900 100.050 ;
        RECT 325.800 97.950 327.900 100.050 ;
        RECT 307.200 91.500 309.300 93.600 ;
        RECT 307.200 86.700 308.700 91.500 ;
        RECT 307.200 84.600 309.300 86.700 ;
        RECT 259.950 70.950 262.050 73.050 ;
        RECT 299.400 72.300 302.400 74.400 ;
        RECT 303.300 72.300 305.400 74.400 ;
        RECT 322.200 72.300 324.300 74.400 ;
        RECT 247.950 64.950 250.050 67.050 ;
        RECT 245.400 62.400 249.450 63.450 ;
        RECT 227.400 58.350 228.600 60.600 ;
        RECT 232.950 58.950 235.050 61.050 ;
        RECT 248.400 60.600 249.450 62.400 ;
        RECT 260.400 61.200 261.450 70.950 ;
        RECT 271.950 64.950 274.050 67.050 ;
        RECT 248.400 58.350 249.600 60.600 ;
        RECT 259.950 59.100 262.050 61.200 ;
        RECT 265.950 59.100 268.050 61.200 ;
        RECT 272.400 60.600 273.450 64.950 ;
        RECT 260.400 58.350 261.600 59.100 ;
        RECT 266.400 58.350 267.600 59.100 ;
        RECT 272.400 58.350 273.600 60.600 ;
        RECT 277.950 60.000 280.050 64.050 ;
        RECT 278.400 58.350 279.600 60.000 ;
        RECT 286.800 58.950 288.900 61.050 ;
        RECT 292.800 58.950 294.900 61.050 ;
        RECT 137.100 55.950 139.200 58.050 ;
        RECT 142.500 55.950 144.600 58.050 ;
        RECT 145.800 55.950 147.900 58.050 ;
        RECT 151.950 55.950 154.050 58.050 ;
        RECT 154.950 55.950 157.050 58.050 ;
        RECT 157.950 55.950 160.050 58.050 ;
        RECT 160.950 55.950 163.050 58.050 ;
        RECT 166.950 55.950 169.050 58.050 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 172.950 55.950 175.050 58.050 ;
        RECT 175.950 55.950 178.050 58.050 ;
        RECT 178.950 55.950 181.050 58.050 ;
        RECT 181.950 55.950 184.050 58.050 ;
        RECT 184.950 55.950 187.050 58.050 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 196.950 55.950 199.050 58.050 ;
        RECT 199.950 55.950 202.050 58.050 ;
        RECT 202.950 55.950 205.050 58.050 ;
        RECT 208.950 55.950 211.050 58.050 ;
        RECT 211.950 55.950 214.050 58.050 ;
        RECT 214.950 55.950 217.050 58.050 ;
        RECT 217.950 55.950 220.050 58.050 ;
        RECT 226.950 55.950 229.050 58.050 ;
        RECT 229.950 55.950 232.050 58.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 241.950 55.950 244.050 58.050 ;
        RECT 244.950 55.950 247.050 58.050 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 250.950 55.950 253.050 58.050 ;
        RECT 259.950 55.950 262.050 58.050 ;
        RECT 262.950 55.950 265.050 58.050 ;
        RECT 265.950 55.950 268.050 58.050 ;
        RECT 271.950 55.950 274.050 58.050 ;
        RECT 274.950 55.950 277.050 58.050 ;
        RECT 277.950 55.950 280.050 58.050 ;
        RECT 280.950 55.950 283.050 58.050 ;
        RECT 143.400 53.400 144.600 55.650 ;
        RECT 133.950 46.950 136.050 49.050 ;
        RECT 143.400 43.050 144.450 53.400 ;
        RECT 148.950 52.950 151.050 55.050 ;
        RECT 152.400 53.400 153.600 55.650 ;
        RECT 158.400 53.400 159.600 55.650 ;
        RECT 149.400 49.050 150.450 52.950 ;
        RECT 148.950 46.950 151.050 49.050 ;
        RECT 152.400 43.050 153.450 53.400 ;
        RECT 142.950 40.950 145.050 43.050 ;
        RECT 151.950 40.950 154.050 43.050 ;
        RECT 130.950 37.950 133.050 40.050 ;
        RECT 127.950 34.950 130.050 37.050 ;
        RECT 115.950 31.950 118.050 34.050 ;
        RECT 128.400 30.450 129.450 34.950 ;
        RECT 130.950 33.450 133.050 34.050 ;
        RECT 130.950 32.400 138.450 33.450 ;
        RECT 130.950 31.950 133.050 32.400 ;
        RECT 125.400 29.400 129.450 30.450 ;
        RECT 94.950 26.100 97.050 28.200 ;
        RECT 109.950 26.100 112.050 28.200 ;
        RECT 115.950 26.100 118.050 28.200 ;
        RECT 125.400 27.600 126.450 29.400 ;
        RECT 95.400 25.350 96.600 26.100 ;
        RECT 116.400 25.350 117.600 26.100 ;
        RECT 125.400 25.350 126.600 27.600 ;
        RECT 133.950 26.100 136.050 28.200 ;
        RECT 134.400 25.350 135.600 26.100 ;
        RECT 89.100 22.950 91.200 25.050 ;
        RECT 94.500 22.950 96.600 25.050 ;
        RECT 104.100 22.950 106.200 25.050 ;
        RECT 107.100 22.950 109.200 25.050 ;
        RECT 112.800 22.950 114.900 25.050 ;
        RECT 115.800 22.950 117.900 25.050 ;
        RECT 121.950 22.950 124.050 25.050 ;
        RECT 124.950 22.950 127.050 25.050 ;
        RECT 128.100 22.950 130.200 25.050 ;
        RECT 133.500 22.950 135.600 25.050 ;
        RECT 104.400 21.000 105.600 22.650 ;
        RECT 82.950 16.950 85.050 19.050 ;
        RECT 103.950 16.950 106.050 21.000 ;
        RECT 113.400 20.400 114.600 22.650 ;
        RECT 122.400 21.900 123.600 22.650 ;
        RECT 58.200 13.500 60.300 15.600 ;
        RECT 58.200 8.700 59.700 13.500 ;
        RECT 113.400 13.050 114.450 20.400 ;
        RECT 121.950 19.800 124.050 21.900 ;
        RECT 122.400 16.050 123.450 19.800 ;
        RECT 121.950 13.950 124.050 16.050 ;
        RECT 137.400 13.050 138.450 32.400 ;
        RECT 142.950 26.100 145.050 31.050 ;
        RECT 152.400 27.450 153.450 40.950 ;
        RECT 158.400 40.050 159.450 53.400 ;
        RECT 163.800 52.950 165.900 55.050 ;
        RECT 167.400 54.900 168.600 55.650 ;
        RECT 160.950 46.950 163.050 49.050 ;
        RECT 157.950 37.950 160.050 40.050 ;
        RECT 161.400 37.050 162.450 46.950 ;
        RECT 160.950 34.950 163.050 37.050 ;
        RECT 154.950 27.450 157.050 28.200 ;
        RECT 152.400 26.400 157.050 27.450 ;
        RECT 154.950 26.100 157.050 26.400 ;
        RECT 161.400 27.600 162.450 34.950 ;
        RECT 164.400 31.050 165.450 52.950 ;
        RECT 166.950 52.800 169.050 54.900 ;
        RECT 182.400 53.400 183.600 55.650 ;
        RECT 178.950 43.950 181.050 46.050 ;
        RECT 179.400 37.050 180.450 43.950 ;
        RECT 182.400 43.050 183.450 53.400 ;
        RECT 190.950 52.950 193.050 55.050 ;
        RECT 197.400 54.000 198.600 55.650 ;
        RECT 203.400 54.000 204.600 55.650 ;
        RECT 184.950 49.950 187.050 52.050 ;
        RECT 181.950 40.950 184.050 43.050 ;
        RECT 185.400 40.050 186.450 49.950 ;
        RECT 191.400 46.050 192.450 52.950 ;
        RECT 196.950 49.950 199.050 54.000 ;
        RECT 202.950 49.950 205.050 54.000 ;
        RECT 205.950 52.950 208.050 55.050 ;
        RECT 212.400 53.400 213.600 55.650 ;
        RECT 218.400 53.400 219.600 55.650 ;
        RECT 190.950 43.950 193.050 46.050 ;
        RECT 184.950 37.950 187.050 40.050 ;
        RECT 199.950 37.950 202.050 40.050 ;
        RECT 178.950 34.950 181.050 37.050 ;
        RECT 172.950 31.950 175.050 34.050 ;
        RECT 163.950 28.950 166.050 31.050 ;
        RECT 173.400 27.600 174.450 31.950 ;
        RECT 143.400 25.350 144.600 26.100 ;
        RECT 155.400 25.350 156.600 26.100 ;
        RECT 161.400 25.350 162.600 27.600 ;
        RECT 173.400 25.350 174.600 27.600 ;
        RECT 181.950 26.100 184.050 28.200 ;
        RECT 193.950 26.100 196.050 28.200 ;
        RECT 200.400 27.600 201.450 37.950 ;
        RECT 206.400 37.050 207.450 52.950 ;
        RECT 212.400 43.050 213.450 53.400 ;
        RECT 211.950 40.950 214.050 43.050 ;
        RECT 205.950 34.950 208.050 37.050 ;
        RECT 214.950 34.950 217.050 37.050 ;
        RECT 215.400 27.600 216.450 34.950 ;
        RECT 218.400 28.050 219.450 53.400 ;
        RECT 220.800 52.950 222.900 55.050 ;
        RECT 223.950 52.950 226.050 55.050 ;
        RECT 230.400 53.400 231.600 55.650 ;
        RECT 239.400 54.900 240.600 55.650 ;
        RECT 245.400 54.900 246.600 55.650 ;
        RECT 221.400 49.050 222.450 52.950 ;
        RECT 220.950 46.950 223.050 49.050 ;
        RECT 224.400 34.050 225.450 52.950 ;
        RECT 230.400 49.050 231.450 53.400 ;
        RECT 238.950 52.800 241.050 54.900 ;
        RECT 244.950 52.800 247.050 54.900 ;
        RECT 251.400 54.000 252.600 55.650 ;
        RECT 229.950 46.950 232.050 49.050 ;
        RECT 223.950 31.950 226.050 34.050 ;
        RECT 182.400 25.350 183.600 26.100 ;
        RECT 194.400 25.350 195.600 26.100 ;
        RECT 200.400 25.350 201.600 27.600 ;
        RECT 215.400 25.350 216.600 27.600 ;
        RECT 217.950 25.950 220.050 28.050 ;
        RECT 224.400 27.600 225.450 31.950 ;
        RECT 230.400 27.600 231.450 46.950 ;
        RECT 235.950 43.950 238.050 46.050 ;
        RECT 232.950 34.950 235.050 37.050 ;
        RECT 233.400 28.050 234.450 34.950 ;
        RECT 224.400 25.350 225.600 27.600 ;
        RECT 230.400 25.350 231.600 27.600 ;
        RECT 232.950 25.950 235.050 28.050 ;
        RECT 236.400 27.600 237.450 43.950 ;
        RECT 239.400 31.050 240.450 52.800 ;
        RECT 247.950 49.950 250.050 52.050 ;
        RECT 250.950 49.950 253.050 54.000 ;
        RECT 263.400 53.400 264.600 55.650 ;
        RECT 263.400 52.050 264.450 53.400 ;
        RECT 268.950 52.950 271.050 55.050 ;
        RECT 275.400 53.400 276.600 55.650 ;
        RECT 281.400 54.900 282.600 55.650 ;
        RECT 259.950 50.400 264.450 52.050 ;
        RECT 259.950 49.950 264.000 50.400 ;
        RECT 241.950 31.950 244.050 34.050 ;
        RECT 238.950 28.950 241.050 31.050 ;
        RECT 242.400 27.600 243.450 31.950 ;
        RECT 248.400 28.050 249.450 49.950 ;
        RECT 265.950 43.950 268.050 46.050 ;
        RECT 253.800 34.950 255.900 37.050 ;
        RECT 254.400 31.050 255.450 34.950 ;
        RECT 256.950 31.950 259.050 34.050 ;
        RECT 253.950 28.950 256.050 31.050 ;
        RECT 236.400 25.350 237.600 27.600 ;
        RECT 242.400 25.350 243.600 27.600 ;
        RECT 247.950 25.950 250.050 28.050 ;
        RECT 257.400 27.600 258.450 31.950 ;
        RECT 266.400 28.050 267.450 43.950 ;
        RECT 269.400 37.050 270.450 52.950 ;
        RECT 275.400 46.050 276.450 53.400 ;
        RECT 280.950 52.800 283.050 54.900 ;
        RECT 299.400 53.400 300.900 72.300 ;
        RECT 303.300 66.300 304.500 72.300 ;
        RECT 302.400 64.200 304.500 66.300 ;
        RECT 299.400 51.300 301.500 53.400 ;
        RECT 300.300 47.700 301.500 51.300 ;
        RECT 303.300 47.700 304.500 64.200 ;
        RECT 305.700 69.300 307.800 71.400 ;
        RECT 305.700 47.700 306.900 69.300 ;
        RECT 314.400 67.800 316.500 69.900 ;
        RECT 319.800 69.300 321.900 71.400 ;
        RECT 314.400 61.200 315.300 67.800 ;
        RECT 320.100 62.100 321.300 69.300 ;
        RECT 322.800 67.500 324.300 72.300 ;
        RECT 325.200 69.300 327.300 74.400 ;
        RECT 322.800 65.400 324.900 67.500 ;
        RECT 314.400 59.100 316.500 61.200 ;
        RECT 319.800 60.000 321.900 62.100 ;
        RECT 307.950 57.600 312.000 58.050 ;
        RECT 307.950 55.950 312.600 57.600 ;
        RECT 311.400 55.350 312.600 55.950 ;
        RECT 310.800 52.950 312.900 55.050 ;
        RECT 314.400 48.600 315.300 59.100 ;
        RECT 317.100 52.500 319.200 54.600 ;
        RECT 274.950 43.950 277.050 46.050 ;
        RECT 299.700 45.600 301.800 47.700 ;
        RECT 302.700 45.600 304.800 47.700 ;
        RECT 305.700 45.600 307.800 47.700 ;
        RECT 313.800 46.500 315.900 48.600 ;
        RECT 320.100 47.700 321.300 60.000 ;
        RECT 322.800 47.700 324.300 65.400 ;
        RECT 326.100 47.700 327.300 69.300 ;
        RECT 319.200 45.600 321.300 47.700 ;
        RECT 322.200 45.600 324.300 47.700 ;
        RECT 325.200 45.600 327.300 47.700 ;
        RECT 328.200 72.300 330.300 74.400 ;
        RECT 328.200 67.500 329.700 72.300 ;
        RECT 328.200 65.400 330.300 67.500 ;
        RECT 328.200 47.700 329.700 65.400 ;
        RECT 337.800 58.950 339.900 61.050 ;
        RECT 346.800 58.950 348.900 61.050 ;
        RECT 347.400 56.400 348.600 58.650 ;
        RECT 328.200 45.600 330.300 47.700 ;
        RECT 347.400 37.050 348.450 56.400 ;
        RECT 268.950 34.950 271.050 37.050 ;
        RECT 275.700 33.300 277.800 35.400 ;
        RECT 278.700 33.300 280.800 35.400 ;
        RECT 281.700 33.300 283.800 35.400 ;
        RECT 276.300 29.700 277.500 33.300 ;
        RECT 257.400 25.350 258.600 27.600 ;
        RECT 265.950 25.950 268.050 28.050 ;
        RECT 275.400 27.600 277.500 29.700 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 145.950 22.950 148.050 25.050 ;
        RECT 154.950 22.950 157.050 25.050 ;
        RECT 157.950 22.950 160.050 25.050 ;
        RECT 160.950 22.950 163.050 25.050 ;
        RECT 167.100 22.950 169.200 25.050 ;
        RECT 172.500 22.950 174.600 25.050 ;
        RECT 175.800 22.950 177.900 25.050 ;
        RECT 178.950 22.950 181.050 25.050 ;
        RECT 182.400 22.950 184.500 25.050 ;
        RECT 187.800 22.950 189.900 25.050 ;
        RECT 193.950 22.950 196.050 25.050 ;
        RECT 196.950 22.950 199.050 25.050 ;
        RECT 199.950 22.950 202.050 25.050 ;
        RECT 202.950 22.950 205.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 220.950 22.950 223.050 25.050 ;
        RECT 223.950 22.950 226.050 25.050 ;
        RECT 226.950 22.950 229.050 25.050 ;
        RECT 229.950 22.950 232.050 25.050 ;
        RECT 235.950 22.950 238.050 25.050 ;
        RECT 238.950 22.950 241.050 25.050 ;
        RECT 241.950 22.950 244.050 25.050 ;
        RECT 244.950 22.950 247.050 25.050 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 146.400 21.900 147.600 22.650 ;
        RECT 158.400 21.900 159.600 22.650 ;
        RECT 167.400 21.900 168.600 22.650 ;
        RECT 176.400 21.900 177.600 22.650 ;
        RECT 145.950 19.800 148.050 21.900 ;
        RECT 157.950 19.800 160.050 21.900 ;
        RECT 166.950 19.800 169.050 21.900 ;
        RECT 175.950 19.800 178.050 21.900 ;
        RECT 179.400 16.050 180.450 22.950 ;
        RECT 197.400 20.400 198.600 22.650 ;
        RECT 203.400 21.900 204.600 22.650 ;
        RECT 212.400 21.900 213.600 22.650 ;
        RECT 178.950 13.950 181.050 16.050 ;
        RECT 112.950 10.950 115.050 13.050 ;
        RECT 136.950 10.950 139.050 13.050 ;
        RECT 58.200 6.600 60.300 8.700 ;
        RECT 197.400 4.050 198.450 20.400 ;
        RECT 202.950 19.800 205.050 21.900 ;
        RECT 211.950 19.800 214.050 21.900 ;
        RECT 217.950 19.950 220.050 22.050 ;
        RECT 221.400 21.000 222.600 22.650 ;
        RECT 239.400 21.900 240.600 22.650 ;
        RECT 245.400 21.900 246.600 22.650 ;
        RECT 254.400 21.900 255.600 22.650 ;
        RECT 218.400 13.050 219.450 19.950 ;
        RECT 220.950 16.950 223.050 21.000 ;
        RECT 238.950 19.800 241.050 21.900 ;
        RECT 244.950 19.800 247.050 21.900 ;
        RECT 253.950 19.800 256.050 21.900 ;
        RECT 262.800 19.950 264.900 22.050 ;
        RECT 268.800 19.950 270.900 22.050 ;
        RECT 217.950 10.950 220.050 13.050 ;
        RECT 254.400 4.050 255.450 19.800 ;
        RECT 275.400 8.700 276.900 27.600 ;
        RECT 279.300 16.800 280.500 33.300 ;
        RECT 278.400 14.700 280.500 16.800 ;
        RECT 279.300 8.700 280.500 14.700 ;
        RECT 281.700 11.700 282.900 33.300 ;
        RECT 289.800 32.400 291.900 34.500 ;
        RECT 295.200 33.300 297.300 35.400 ;
        RECT 298.200 33.300 300.300 35.400 ;
        RECT 301.200 33.300 303.300 35.400 ;
        RECT 286.800 25.950 288.900 28.050 ;
        RECT 287.400 23.400 288.600 25.650 ;
        RECT 287.400 13.050 288.450 23.400 ;
        RECT 290.400 21.900 291.300 32.400 ;
        RECT 293.100 26.400 295.200 28.500 ;
        RECT 290.400 19.800 292.500 21.900 ;
        RECT 296.100 21.000 297.300 33.300 ;
        RECT 290.400 13.200 291.300 19.800 ;
        RECT 295.800 18.900 297.900 21.000 ;
        RECT 281.700 9.600 283.800 11.700 ;
        RECT 286.950 10.950 289.050 13.050 ;
        RECT 290.400 11.100 292.500 13.200 ;
        RECT 296.100 11.700 297.300 18.900 ;
        RECT 298.800 15.600 300.300 33.300 ;
        RECT 298.800 13.500 300.900 15.600 ;
        RECT 295.800 9.600 297.900 11.700 ;
        RECT 298.800 8.700 300.300 13.500 ;
        RECT 302.100 11.700 303.300 33.300 ;
        RECT 275.400 6.600 278.400 8.700 ;
        RECT 279.300 6.600 281.400 8.700 ;
        RECT 298.200 6.600 300.300 8.700 ;
        RECT 301.200 6.600 303.300 11.700 ;
        RECT 304.200 33.300 306.300 35.400 ;
        RECT 346.950 34.950 349.050 37.050 ;
        RECT 304.200 15.600 305.700 33.300 ;
        RECT 334.950 31.950 337.050 34.050 ;
        RECT 322.950 28.950 325.050 31.050 ;
        RECT 323.400 24.600 324.450 28.950 ;
        RECT 335.400 27.600 336.450 31.950 ;
        RECT 347.400 27.600 348.450 34.950 ;
        RECT 335.400 25.350 336.600 27.600 ;
        RECT 347.400 25.350 348.600 27.600 ;
        RECT 323.400 22.350 324.600 24.600 ;
        RECT 335.400 22.950 337.500 25.050 ;
        RECT 340.800 22.950 342.900 25.050 ;
        RECT 347.400 22.950 349.500 25.050 ;
        RECT 352.800 22.950 354.900 25.050 ;
        RECT 313.800 19.950 315.900 22.050 ;
        RECT 322.800 19.950 324.900 22.050 ;
        RECT 304.200 13.500 306.300 15.600 ;
        RECT 304.200 8.700 305.700 13.500 ;
        RECT 304.200 6.600 306.300 8.700 ;
        RECT 196.950 1.950 199.050 4.050 ;
        RECT 253.950 1.950 256.050 4.050 ;
      LAYER metal3 ;
        RECT 139.950 354.600 142.050 355.050 ;
        RECT 160.950 354.600 163.050 355.050 ;
        RECT 139.950 353.400 163.050 354.600 ;
        RECT 139.950 352.950 142.050 353.400 ;
        RECT 160.950 352.950 163.050 353.400 ;
        RECT 166.950 354.600 169.050 355.050 ;
        RECT 190.950 354.600 193.050 355.050 ;
        RECT 166.950 353.400 193.050 354.600 ;
        RECT 166.950 352.950 169.050 353.400 ;
        RECT 190.950 352.950 193.050 353.400 ;
        RECT 253.950 348.600 256.050 349.050 ;
        RECT 277.950 348.600 280.050 349.050 ;
        RECT 253.950 347.400 280.050 348.600 ;
        RECT 253.950 346.950 256.050 347.400 ;
        RECT 277.950 346.950 280.050 347.400 ;
        RECT 133.950 345.600 136.050 346.050 ;
        RECT 154.950 345.600 157.050 346.050 ;
        RECT 166.950 345.600 169.050 346.050 ;
        RECT 133.950 344.400 169.050 345.600 ;
        RECT 133.950 343.950 136.050 344.400 ;
        RECT 154.950 343.950 157.050 344.400 ;
        RECT 166.950 343.950 169.050 344.400 ;
        RECT 220.950 342.600 223.050 342.900 ;
        RECT 212.400 341.400 223.050 342.600 ;
        RECT 145.950 338.100 148.050 340.200 ;
        RECT 199.950 339.600 202.050 340.050 ;
        RECT 208.950 339.600 211.050 340.200 ;
        RECT 199.950 338.400 211.050 339.600 ;
        RECT 118.950 336.600 121.050 337.050 ;
        RECT 146.400 336.600 147.600 338.100 ;
        RECT 199.950 337.950 202.050 338.400 ;
        RECT 208.950 338.100 211.050 338.400 ;
        RECT 118.950 335.400 156.600 336.600 ;
        RECT 118.950 334.950 121.050 335.400 ;
        RECT 155.400 333.600 156.600 335.400 ;
        RECT 212.400 333.900 213.600 341.400 ;
        RECT 220.950 340.800 223.050 341.400 ;
        RECT 214.950 339.600 217.050 340.200 ;
        RECT 226.950 339.600 229.050 340.200 ;
        RECT 238.950 339.600 241.050 340.200 ;
        RECT 214.950 338.400 241.050 339.600 ;
        RECT 214.950 338.100 217.050 338.400 ;
        RECT 226.950 338.100 229.050 338.400 ;
        RECT 238.950 338.100 241.050 338.400 ;
        RECT 247.950 338.100 250.050 340.200 ;
        RECT 262.950 338.100 265.050 340.200 ;
        RECT 349.950 339.600 352.050 340.200 ;
        RECT 349.950 338.400 357.600 339.600 ;
        RECT 349.950 338.100 352.050 338.400 ;
        RECT 227.400 334.050 228.600 338.100 ;
        RECT 163.950 333.600 166.050 333.900 ;
        RECT 155.400 332.400 166.050 333.600 ;
        RECT 163.950 331.800 166.050 332.400 ;
        RECT 211.950 331.800 214.050 333.900 ;
        RECT 227.400 332.400 232.050 334.050 ;
        RECT 228.000 331.950 232.050 332.400 ;
        RECT 241.950 333.600 244.050 333.900 ;
        RECT 248.400 333.600 249.600 338.100 ;
        RECT 241.950 332.400 249.600 333.600 ;
        RECT 241.950 331.800 244.050 332.400 ;
        RECT 263.400 331.050 264.600 338.100 ;
        RECT 277.950 336.450 280.050 336.900 ;
        RECT 298.950 336.450 301.050 336.900 ;
        RECT 277.950 335.250 301.050 336.450 ;
        RECT 277.950 334.800 280.050 335.250 ;
        RECT 298.950 334.800 301.050 335.250 ;
        RECT 356.400 334.050 357.600 338.400 ;
        RECT 355.950 331.950 358.050 334.050 ;
        RECT 169.950 330.600 172.050 331.050 ;
        RECT 184.950 330.600 187.050 331.050 ;
        RECT 169.950 329.400 187.050 330.600 ;
        RECT 169.950 328.950 172.050 329.400 ;
        RECT 184.950 328.950 187.050 329.400 ;
        RECT 190.950 330.600 193.050 331.050 ;
        RECT 211.950 330.600 214.050 331.050 ;
        RECT 190.950 329.400 214.050 330.600 ;
        RECT 190.950 328.950 193.050 329.400 ;
        RECT 211.950 328.950 214.050 329.400 ;
        RECT 262.950 328.950 265.050 331.050 ;
        RECT 28.950 327.600 31.050 328.050 ;
        RECT 52.950 327.600 55.050 328.050 ;
        RECT 28.950 326.400 55.050 327.600 ;
        RECT 28.950 325.950 31.050 326.400 ;
        RECT 52.950 325.950 55.050 326.400 ;
        RECT 241.950 327.600 244.050 328.050 ;
        RECT 256.950 327.600 259.050 328.050 ;
        RECT 241.950 326.400 259.050 327.600 ;
        RECT 241.950 325.950 244.050 326.400 ;
        RECT 256.950 325.950 259.050 326.400 ;
        RECT 58.950 324.600 61.050 325.050 ;
        RECT 67.950 324.600 70.050 325.050 ;
        RECT 169.950 324.600 172.050 325.050 ;
        RECT 58.950 323.400 172.050 324.600 ;
        RECT 58.950 322.950 61.050 323.400 ;
        RECT 67.950 322.950 70.050 323.400 ;
        RECT 169.950 322.950 172.050 323.400 ;
        RECT 97.950 321.600 100.050 322.050 ;
        RECT 169.950 321.600 172.050 321.900 ;
        RECT 97.950 320.400 172.050 321.600 ;
        RECT 97.950 319.950 100.050 320.400 ;
        RECT 169.950 319.800 172.050 320.400 ;
        RECT 211.950 321.600 214.050 322.050 ;
        RECT 232.950 321.600 235.050 322.050 ;
        RECT 211.950 320.400 235.050 321.600 ;
        RECT 211.950 319.950 214.050 320.400 ;
        RECT 232.950 319.950 235.050 320.400 ;
        RECT 133.950 318.600 136.050 319.050 ;
        RECT 199.950 318.600 202.050 319.050 ;
        RECT 250.950 318.600 253.050 319.050 ;
        RECT 133.950 317.400 159.600 318.600 ;
        RECT 133.950 316.950 136.050 317.400 ;
        RECT 158.400 315.600 159.600 317.400 ;
        RECT 199.950 317.400 253.050 318.600 ;
        RECT 199.950 316.950 202.050 317.400 ;
        RECT 250.950 316.950 253.050 317.400 ;
        RECT 193.950 315.600 196.050 316.050 ;
        RECT 214.950 315.600 217.050 316.050 ;
        RECT 158.400 314.400 217.050 315.600 ;
        RECT 193.950 313.950 196.050 314.400 ;
        RECT 214.950 313.950 217.050 314.400 ;
        RECT 262.950 315.600 265.050 316.050 ;
        RECT 310.950 315.600 313.050 316.050 ;
        RECT 337.950 315.600 340.050 316.050 ;
        RECT 262.950 314.400 340.050 315.600 ;
        RECT 262.950 313.950 265.050 314.400 ;
        RECT 310.950 313.950 313.050 314.400 ;
        RECT 337.950 313.950 340.050 314.400 ;
        RECT 139.950 312.600 142.050 313.050 ;
        RECT 154.950 312.600 157.050 313.050 ;
        RECT 190.950 312.600 193.050 313.050 ;
        RECT 139.950 311.400 193.050 312.600 ;
        RECT 139.950 310.950 142.050 311.400 ;
        RECT 154.950 310.950 157.050 311.400 ;
        RECT 190.950 310.950 193.050 311.400 ;
        RECT 94.950 309.600 97.050 310.050 ;
        RECT 115.950 309.600 118.050 310.050 ;
        RECT 94.950 308.400 118.050 309.600 ;
        RECT 94.950 307.950 97.050 308.400 ;
        RECT 115.950 307.950 118.050 308.400 ;
        RECT 163.950 309.600 166.050 310.050 ;
        RECT 205.950 309.600 208.050 310.050 ;
        RECT 163.950 308.400 208.050 309.600 ;
        RECT 163.950 307.950 166.050 308.400 ;
        RECT 205.950 307.950 208.050 308.400 ;
        RECT 70.950 306.600 73.050 307.050 ;
        RECT 91.950 306.600 94.050 307.050 ;
        RECT 118.950 306.600 121.050 307.050 ;
        RECT 70.950 305.400 121.050 306.600 ;
        RECT 70.950 304.950 73.050 305.400 ;
        RECT 91.950 304.950 94.050 305.400 ;
        RECT 118.950 304.950 121.050 305.400 ;
        RECT 235.950 306.600 238.050 307.050 ;
        RECT 253.950 306.600 256.050 307.050 ;
        RECT 235.950 305.400 256.050 306.600 ;
        RECT 235.950 304.950 238.050 305.400 ;
        RECT 253.950 304.950 256.050 305.400 ;
        RECT 112.950 303.600 115.050 304.050 ;
        RECT 133.950 303.600 136.050 304.050 ;
        RECT 112.950 302.400 136.050 303.600 ;
        RECT 112.950 301.950 115.050 302.400 ;
        RECT 133.950 301.950 136.050 302.400 ;
        RECT 217.950 303.600 220.050 304.050 ;
        RECT 223.950 303.600 226.050 304.050 ;
        RECT 217.950 302.400 226.050 303.600 ;
        RECT 217.950 301.950 220.050 302.400 ;
        RECT 223.950 301.950 226.050 302.400 ;
        RECT 229.950 303.600 232.050 304.050 ;
        RECT 256.950 303.600 259.050 304.050 ;
        RECT 229.950 302.400 259.050 303.600 ;
        RECT 229.950 301.950 232.050 302.400 ;
        RECT 256.950 301.950 259.050 302.400 ;
        RECT 265.950 303.600 268.050 304.050 ;
        RECT 280.950 303.600 283.050 304.050 ;
        RECT 331.950 303.600 334.050 304.050 ;
        RECT 265.950 302.400 334.050 303.600 ;
        RECT 265.950 301.950 268.050 302.400 ;
        RECT 280.950 301.950 283.050 302.400 ;
        RECT 331.950 301.950 334.050 302.400 ;
        RECT 28.950 300.600 31.050 301.050 ;
        RECT 67.950 300.600 70.050 301.050 ;
        RECT 28.950 299.400 70.050 300.600 ;
        RECT 28.950 298.950 31.050 299.400 ;
        RECT 67.950 298.950 70.050 299.400 ;
        RECT 79.950 300.600 82.050 301.050 ;
        RECT 94.950 300.600 97.050 301.050 ;
        RECT 79.950 299.400 97.050 300.600 ;
        RECT 79.950 298.950 82.050 299.400 ;
        RECT 94.950 298.950 97.050 299.400 ;
        RECT 136.950 300.600 139.050 301.050 ;
        RECT 187.950 300.600 190.050 301.050 ;
        RECT 208.950 300.600 211.050 301.050 ;
        RECT 136.950 299.400 211.050 300.600 ;
        RECT 136.950 298.950 139.050 299.400 ;
        RECT 187.950 298.950 190.050 299.400 ;
        RECT 208.950 298.950 211.050 299.400 ;
        RECT 52.950 297.600 55.050 298.050 ;
        RECT 85.950 297.600 88.050 298.050 ;
        RECT 163.950 297.600 166.050 298.050 ;
        RECT 52.950 296.400 69.600 297.600 ;
        RECT 52.950 295.950 55.050 296.400 ;
        RECT 68.400 294.600 69.600 296.400 ;
        RECT 85.950 296.400 111.600 297.600 ;
        RECT 85.950 295.950 88.050 296.400 ;
        RECT 68.400 293.400 75.600 294.600 ;
        RECT 64.950 291.450 67.050 291.900 ;
        RECT 70.950 291.450 73.050 291.900 ;
        RECT 64.950 290.250 73.050 291.450 ;
        RECT 64.950 289.800 67.050 290.250 ;
        RECT 70.950 289.800 73.050 290.250 ;
        RECT 74.400 285.600 75.600 293.400 ;
        RECT 97.950 293.100 100.050 295.200 ;
        RECT 82.950 288.600 85.050 288.900 ;
        RECT 94.950 288.600 97.050 288.900 ;
        RECT 82.950 287.400 97.050 288.600 ;
        RECT 82.950 286.800 85.050 287.400 ;
        RECT 94.950 286.800 97.050 287.400 ;
        RECT 98.400 286.050 99.600 293.100 ;
        RECT 110.400 288.900 111.600 296.400 ;
        RECT 155.400 296.400 166.050 297.600 ;
        RECT 115.950 292.950 118.050 295.050 ;
        RECT 121.950 294.600 124.050 295.200 ;
        RECT 130.950 294.600 133.050 295.200 ;
        RECT 121.950 293.400 133.050 294.600 ;
        RECT 121.950 293.100 124.050 293.400 ;
        RECT 130.950 293.100 133.050 293.400 ;
        RECT 148.950 293.100 151.050 295.200 ;
        RECT 109.950 286.800 112.050 288.900 ;
        RECT 79.950 285.600 82.050 286.050 ;
        RECT 74.400 284.400 82.050 285.600 ;
        RECT 79.950 283.950 82.050 284.400 ;
        RECT 97.950 285.600 100.050 286.050 ;
        RECT 112.950 285.600 115.050 286.050 ;
        RECT 97.950 284.400 115.050 285.600 ;
        RECT 116.400 285.600 117.600 292.950 ;
        RECT 133.950 288.600 136.050 288.900 ;
        RECT 149.400 288.600 150.600 293.100 ;
        RECT 155.400 291.600 156.600 296.400 ;
        RECT 163.950 295.950 166.050 296.400 ;
        RECT 184.950 297.600 187.050 298.050 ;
        RECT 199.950 297.600 202.050 298.050 ;
        RECT 184.950 296.400 202.050 297.600 ;
        RECT 184.950 295.950 187.050 296.400 ;
        RECT 199.950 295.950 202.050 296.400 ;
        RECT 217.950 295.950 220.050 298.050 ;
        RECT 232.950 297.600 237.000 298.050 ;
        RECT 253.950 297.600 258.000 298.050 ;
        RECT 232.950 295.950 237.600 297.600 ;
        RECT 253.950 295.950 258.600 297.600 ;
        RECT 157.950 294.600 162.000 295.050 ;
        RECT 157.950 292.950 162.600 294.600 ;
        RECT 169.950 292.950 172.050 295.050 ;
        RECT 175.950 293.100 178.050 295.200 ;
        RECT 181.950 293.100 184.050 295.200 ;
        RECT 152.400 290.400 156.600 291.600 ;
        RECT 152.400 288.900 153.600 290.400 ;
        RECT 161.400 289.050 162.600 292.950 ;
        RECT 133.950 287.400 150.600 288.600 ;
        RECT 133.950 286.800 136.050 287.400 ;
        RECT 151.950 286.800 154.050 288.900 ;
        RECT 160.950 286.950 163.050 289.050 ;
        RECT 170.400 288.600 171.600 292.950 ;
        RECT 172.950 288.600 175.050 288.900 ;
        RECT 170.400 287.400 175.050 288.600 ;
        RECT 172.950 286.800 175.050 287.400 ;
        RECT 176.400 286.050 177.600 293.100 ;
        RECT 182.400 291.600 183.600 293.100 ;
        RECT 193.950 291.600 196.050 295.050 ;
        RECT 205.800 293.100 207.900 295.200 ;
        RECT 182.400 291.000 186.600 291.600 ;
        RECT 193.950 291.000 198.600 291.600 ;
        RECT 182.400 290.400 187.050 291.000 ;
        RECT 194.400 290.400 198.600 291.000 ;
        RECT 184.950 286.950 187.050 290.400 ;
        RECT 197.400 288.900 198.600 290.400 ;
        RECT 196.950 286.800 199.050 288.900 ;
        RECT 206.250 286.050 207.450 293.100 ;
        RECT 208.950 292.950 211.050 295.050 ;
        RECT 209.400 289.050 210.600 292.950 ;
        RECT 208.950 286.950 211.050 289.050 ;
        RECT 218.400 286.050 219.600 295.950 ;
        RECT 229.950 293.100 232.050 295.200 ;
        RECT 230.400 286.050 231.600 293.100 ;
        RECT 236.400 286.050 237.600 295.950 ;
        RECT 250.950 293.100 253.050 295.200 ;
        RECT 257.400 294.600 258.600 295.950 ;
        RECT 265.950 294.600 268.050 295.200 ;
        RECT 257.400 293.400 268.050 294.600 ;
        RECT 265.950 293.100 268.050 293.400 ;
        RECT 251.400 288.600 252.600 293.100 ;
        RECT 307.800 291.600 309.900 292.050 ;
        RECT 293.400 290.400 309.900 291.600 ;
        RECT 256.950 288.600 259.050 288.900 ;
        RECT 251.400 287.400 259.050 288.600 ;
        RECT 256.950 286.800 259.050 287.400 ;
        RECT 262.950 288.600 265.050 288.900 ;
        RECT 293.400 288.600 294.600 290.400 ;
        RECT 307.800 289.950 309.900 290.400 ;
        RECT 310.950 291.750 313.050 292.200 ;
        RECT 334.950 291.750 337.050 292.200 ;
        RECT 310.950 290.550 337.050 291.750 ;
        RECT 310.950 290.100 313.050 290.550 ;
        RECT 334.950 290.100 337.050 290.550 ;
        RECT 262.950 287.400 294.600 288.600 ;
        RECT 262.950 286.800 265.050 287.400 ;
        RECT 145.950 285.600 148.050 286.050 ;
        RECT 116.400 284.400 148.050 285.600 ;
        RECT 97.950 283.950 100.050 284.400 ;
        RECT 112.950 283.950 115.050 284.400 ;
        RECT 145.950 283.950 148.050 284.400 ;
        RECT 175.950 283.950 178.050 286.050 ;
        RECT 205.800 283.950 207.900 286.050 ;
        RECT 214.950 284.400 219.600 286.050 ;
        RECT 214.950 283.950 219.000 284.400 ;
        RECT 229.950 283.950 232.050 286.050 ;
        RECT 235.950 283.950 238.050 286.050 ;
        RECT 67.950 282.600 70.050 283.050 ;
        RECT 76.950 282.600 79.050 283.050 ;
        RECT 67.950 281.400 79.050 282.600 ;
        RECT 67.950 280.950 70.050 281.400 ;
        RECT 76.950 280.950 79.050 281.400 ;
        RECT 157.950 282.600 160.050 283.050 ;
        RECT 166.950 282.600 169.050 283.050 ;
        RECT 157.950 281.400 169.050 282.600 ;
        RECT 157.950 280.950 160.050 281.400 ;
        RECT 166.950 280.950 169.050 281.400 ;
        RECT 178.950 282.600 181.050 283.050 ;
        RECT 208.950 282.600 211.050 283.050 ;
        RECT 178.950 281.400 211.050 282.600 ;
        RECT 178.950 280.950 181.050 281.400 ;
        RECT 208.950 280.950 211.050 281.400 ;
        RECT 73.950 279.600 76.050 280.050 ;
        RECT 139.950 279.600 142.050 280.050 ;
        RECT 175.950 279.600 178.050 280.050 ;
        RECT 73.950 278.400 178.050 279.600 ;
        RECT 73.950 277.950 76.050 278.400 ;
        RECT 139.950 277.950 142.050 278.400 ;
        RECT 175.950 277.950 178.050 278.400 ;
        RECT 184.950 279.600 187.050 280.050 ;
        RECT 202.950 279.600 205.050 280.050 ;
        RECT 184.950 278.400 205.050 279.600 ;
        RECT 184.950 277.950 187.050 278.400 ;
        RECT 202.950 277.950 205.050 278.400 ;
        RECT 217.950 279.600 220.050 280.050 ;
        RECT 244.950 279.600 247.050 280.050 ;
        RECT 217.950 278.400 247.050 279.600 ;
        RECT 217.950 277.950 220.050 278.400 ;
        RECT 244.950 277.950 247.050 278.400 ;
        RECT 79.950 276.600 82.050 277.050 ;
        RECT 106.950 276.600 109.050 277.050 ;
        RECT 79.950 275.400 109.050 276.600 ;
        RECT 79.950 274.950 82.050 275.400 ;
        RECT 106.950 274.950 109.050 275.400 ;
        RECT 205.950 276.600 208.050 277.050 ;
        RECT 232.950 276.600 235.050 277.050 ;
        RECT 205.950 275.400 235.050 276.600 ;
        RECT 205.950 274.950 208.050 275.400 ;
        RECT 232.950 274.950 235.050 275.400 ;
        RECT 58.950 273.600 61.050 274.050 ;
        RECT 73.950 273.600 76.050 274.050 ;
        RECT 58.950 272.400 76.050 273.600 ;
        RECT 58.950 271.950 61.050 272.400 ;
        RECT 73.950 271.950 76.050 272.400 ;
        RECT 169.950 270.600 172.050 271.050 ;
        RECT 181.950 270.600 184.050 271.050 ;
        RECT 190.950 270.600 193.050 271.050 ;
        RECT 169.950 269.400 193.050 270.600 ;
        RECT 169.950 268.950 172.050 269.400 ;
        RECT 181.950 268.950 184.050 269.400 ;
        RECT 190.950 268.950 193.050 269.400 ;
        RECT 199.950 270.600 202.050 271.050 ;
        RECT 205.950 270.600 208.050 271.050 ;
        RECT 199.950 269.400 208.050 270.600 ;
        RECT 199.950 268.950 202.050 269.400 ;
        RECT 205.950 268.950 208.050 269.400 ;
        RECT 268.950 270.600 271.050 271.050 ;
        RECT 310.950 270.600 313.050 271.050 ;
        RECT 268.950 269.400 313.050 270.600 ;
        RECT 268.950 268.950 271.050 269.400 ;
        RECT 310.950 268.950 313.050 269.400 ;
        RECT 70.950 267.600 73.050 268.050 ;
        RECT 118.950 267.600 121.050 268.050 ;
        RECT 70.950 266.400 121.050 267.600 ;
        RECT 70.950 265.950 73.050 266.400 ;
        RECT 118.950 265.950 121.050 266.400 ;
        RECT 166.950 267.600 171.000 268.050 ;
        RECT 175.950 267.600 178.050 268.050 ;
        RECT 196.950 267.600 199.050 268.050 ;
        RECT 166.950 265.950 171.600 267.600 ;
        RECT 175.950 266.400 199.050 267.600 ;
        RECT 175.950 265.950 178.050 266.400 ;
        RECT 196.950 265.950 199.050 266.400 ;
        RECT 256.950 267.600 259.050 268.050 ;
        RECT 331.950 267.600 334.050 268.050 ;
        RECT 346.950 267.600 349.050 268.050 ;
        RECT 256.950 266.400 349.050 267.600 ;
        RECT 256.950 265.950 259.050 266.400 ;
        RECT 170.400 264.600 171.600 265.950 ;
        RECT 170.400 263.400 177.600 264.600 ;
        RECT 1.950 261.750 4.050 262.200 ;
        RECT 13.950 261.750 16.050 262.200 ;
        RECT 1.950 260.550 16.050 261.750 ;
        RECT 91.950 261.600 94.050 262.200 ;
        RECT 96.000 261.600 99.900 262.050 ;
        RECT 1.950 260.100 4.050 260.550 ;
        RECT 13.950 260.100 16.050 260.550 ;
        RECT 86.400 260.400 94.050 261.600 ;
        RECT 86.400 256.050 87.600 260.400 ;
        RECT 91.950 260.100 94.050 260.400 ;
        RECT 95.400 259.950 99.900 261.600 ;
        RECT 112.950 261.600 115.050 262.200 ;
        RECT 121.950 261.600 124.050 262.200 ;
        RECT 112.950 260.400 124.050 261.600 ;
        RECT 112.950 260.100 115.050 260.400 ;
        RECT 121.950 260.100 124.050 260.400 ;
        RECT 145.950 259.950 148.050 262.050 ;
        RECT 151.950 260.100 154.050 262.200 ;
        RECT 85.950 253.950 88.050 256.050 ;
        RECT 95.400 255.900 96.600 259.950 ;
        RECT 94.950 253.800 97.050 255.900 ;
        RECT 139.950 255.600 142.050 255.900 ;
        RECT 146.400 255.600 147.600 259.950 ;
        RECT 139.950 254.400 147.600 255.600 ;
        RECT 139.950 253.800 142.050 254.400 ;
        RECT 148.950 253.800 151.050 255.900 ;
        RECT 152.400 255.600 153.600 260.100 ;
        RECT 166.950 259.950 169.050 262.050 ;
        RECT 160.800 255.600 162.900 256.050 ;
        RECT 167.400 255.600 168.600 259.950 ;
        RECT 176.400 255.900 177.600 263.400 ;
        RECT 187.950 262.950 193.050 265.050 ;
        RECT 213.000 264.600 217.050 265.050 ;
        RECT 212.400 262.950 217.050 264.600 ;
        RECT 181.950 261.600 184.050 262.050 ;
        RECT 195.000 261.600 199.050 262.050 ;
        RECT 181.950 260.400 189.600 261.600 ;
        RECT 181.950 259.950 184.050 260.400 ;
        RECT 188.400 255.900 189.600 260.400 ;
        RECT 194.400 259.950 199.050 261.600 ;
        RECT 202.950 260.100 205.050 262.200 ;
        RECT 194.400 255.900 195.600 259.950 ;
        RECT 203.400 256.050 204.600 260.100 ;
        RECT 152.400 254.400 162.900 255.600 ;
        RECT 160.800 253.950 162.900 254.400 ;
        RECT 164.400 254.400 168.600 255.600 ;
        RECT 149.400 253.050 150.600 253.800 ;
        RECT 164.400 253.050 165.600 254.400 ;
        RECT 175.950 253.800 178.050 255.900 ;
        RECT 187.950 253.800 190.050 255.900 ;
        RECT 193.950 253.800 196.050 255.900 ;
        RECT 203.400 254.400 208.050 256.050 ;
        RECT 212.400 255.900 213.600 262.950 ;
        RECT 217.950 260.100 220.050 262.200 ;
        RECT 204.000 253.950 208.050 254.400 ;
        RECT 211.950 253.800 214.050 255.900 ;
        RECT 218.400 255.600 219.600 260.100 ;
        RECT 235.950 259.950 238.050 262.050 ;
        RECT 268.950 259.950 271.050 262.050 ;
        RECT 274.950 261.600 277.050 262.200 ;
        RECT 274.950 260.400 282.450 261.600 ;
        RECT 274.950 260.100 277.050 260.400 ;
        RECT 236.400 256.050 237.600 259.950 ;
        RECT 269.400 256.050 270.600 259.950 ;
        RECT 281.250 256.050 282.450 260.400 ;
        RECT 289.950 260.100 292.050 262.200 ;
        RECT 290.400 258.600 291.600 260.100 ;
        RECT 284.400 258.000 291.600 258.600 ;
        RECT 283.950 257.400 291.600 258.000 ;
        RECT 226.950 255.600 229.050 255.900 ;
        RECT 218.400 254.400 229.050 255.600 ;
        RECT 226.950 253.800 229.050 254.400 ;
        RECT 235.950 253.950 238.050 256.050 ;
        RECT 256.950 255.600 259.050 255.900 ;
        RECT 268.950 255.600 271.050 256.050 ;
        RECT 256.950 254.400 271.050 255.600 ;
        RECT 256.950 253.800 259.050 254.400 ;
        RECT 268.950 253.950 271.050 254.400 ;
        RECT 280.800 253.950 282.900 256.050 ;
        RECT 283.950 253.950 286.050 257.400 ;
        RECT 296.400 255.900 297.600 266.400 ;
        RECT 331.950 265.950 334.050 266.400 ;
        RECT 346.950 265.950 349.050 266.400 ;
        RECT 352.950 265.050 355.050 265.200 ;
        RECT 352.950 264.600 357.000 265.050 ;
        RECT 352.950 263.100 357.600 264.600 ;
        RECT 354.000 262.950 357.600 263.100 ;
        RECT 304.950 261.600 307.050 262.200 ;
        RECT 316.950 261.600 319.050 262.200 ;
        RECT 304.950 260.400 309.600 261.600 ;
        RECT 304.950 260.100 307.050 260.400 ;
        RECT 292.950 255.600 295.050 255.900 ;
        RECT 295.950 255.600 298.050 255.900 ;
        RECT 292.950 254.400 298.050 255.600 ;
        RECT 308.400 255.600 309.600 260.400 ;
        RECT 316.950 260.400 330.600 261.600 ;
        RECT 316.950 260.100 319.050 260.400 ;
        RECT 325.800 255.600 327.900 256.050 ;
        RECT 329.400 255.900 330.600 260.400 ;
        RECT 331.950 260.100 334.050 262.200 ;
        RECT 308.400 254.400 327.900 255.600 ;
        RECT 109.950 252.600 112.050 253.050 ;
        RECT 121.950 252.600 124.050 253.050 ;
        RECT 109.950 251.400 124.050 252.600 ;
        RECT 109.950 250.950 112.050 251.400 ;
        RECT 121.950 250.950 124.050 251.400 ;
        RECT 145.950 252.600 150.600 253.050 ;
        RECT 163.950 252.600 166.050 253.050 ;
        RECT 145.950 251.400 166.050 252.600 ;
        RECT 145.950 250.950 150.000 251.400 ;
        RECT 163.950 250.950 166.050 251.400 ;
        RECT 259.950 252.600 262.050 253.050 ;
        RECT 281.400 252.600 282.600 253.950 ;
        RECT 292.950 253.800 295.050 254.400 ;
        RECT 295.950 253.800 298.050 254.400 ;
        RECT 325.800 253.950 327.900 254.400 ;
        RECT 328.950 253.800 331.050 255.900 ;
        RECT 332.400 255.600 333.600 260.100 ;
        RECT 343.950 259.950 346.050 262.050 ;
        RECT 352.950 259.950 355.050 262.050 ;
        RECT 344.400 256.050 345.600 259.950 ;
        RECT 340.800 255.600 342.900 256.050 ;
        RECT 332.400 254.400 342.900 255.600 ;
        RECT 340.800 253.950 342.900 254.400 ;
        RECT 343.950 253.950 346.050 256.050 ;
        RECT 353.400 253.050 354.600 259.950 ;
        RECT 356.400 255.600 357.600 262.950 ;
        RECT 356.400 255.000 360.600 255.600 ;
        RECT 356.400 254.400 361.050 255.000 ;
        RECT 259.950 251.400 282.600 252.600 ;
        RECT 259.950 250.950 262.050 251.400 ;
        RECT 352.950 250.950 355.050 253.050 ;
        RECT 358.950 250.950 361.050 254.400 ;
        RECT 85.950 249.600 88.050 250.050 ;
        RECT 103.950 249.600 106.050 250.050 ;
        RECT 85.950 248.400 106.050 249.600 ;
        RECT 85.950 247.950 88.050 248.400 ;
        RECT 103.950 247.950 106.050 248.400 ;
        RECT 235.950 249.600 238.050 250.050 ;
        RECT 265.950 249.600 268.050 250.050 ;
        RECT 235.950 248.400 268.050 249.600 ;
        RECT 235.950 247.950 238.050 248.400 ;
        RECT 265.950 247.950 268.050 248.400 ;
        RECT 325.950 249.600 328.050 250.050 ;
        RECT 355.950 249.600 358.050 250.050 ;
        RECT 325.950 248.400 358.050 249.600 ;
        RECT 325.950 247.950 328.050 248.400 ;
        RECT 355.950 247.950 358.050 248.400 ;
        RECT 124.950 246.600 127.050 247.050 ;
        RECT 199.950 246.600 202.050 247.050 ;
        RECT 124.950 245.400 202.050 246.600 ;
        RECT 124.950 244.950 127.050 245.400 ;
        RECT 199.950 244.950 202.050 245.400 ;
        RECT 334.950 246.600 337.050 247.050 ;
        RECT 352.950 246.600 355.050 247.050 ;
        RECT 334.950 245.400 355.050 246.600 ;
        RECT 334.950 244.950 337.050 245.400 ;
        RECT 352.950 244.950 355.050 245.400 ;
        RECT 130.950 243.600 133.050 244.050 ;
        RECT 151.950 243.600 154.050 244.050 ;
        RECT 160.800 243.600 162.900 244.050 ;
        RECT 130.950 242.400 162.900 243.600 ;
        RECT 130.950 241.950 133.050 242.400 ;
        RECT 151.950 241.950 154.050 242.400 ;
        RECT 160.800 241.950 162.900 242.400 ;
        RECT 163.950 243.600 166.050 244.050 ;
        RECT 205.950 243.600 208.050 244.050 ;
        RECT 163.950 242.400 208.050 243.600 ;
        RECT 163.950 241.950 166.050 242.400 ;
        RECT 205.950 241.950 208.050 242.400 ;
        RECT 283.950 243.600 286.050 244.050 ;
        RECT 319.950 243.600 322.050 244.050 ;
        RECT 283.950 242.400 322.050 243.600 ;
        RECT 283.950 241.950 286.050 242.400 ;
        RECT 319.950 241.950 322.050 242.400 ;
        RECT 1.950 240.600 4.050 241.050 ;
        RECT 82.950 240.600 85.050 241.050 ;
        RECT 94.950 240.600 97.050 241.050 ;
        RECT 1.950 239.400 97.050 240.600 ;
        RECT 1.950 238.950 4.050 239.400 ;
        RECT 82.950 238.950 85.050 239.400 ;
        RECT 94.950 238.950 97.050 239.400 ;
        RECT 169.950 240.600 172.050 241.050 ;
        RECT 190.950 240.600 193.050 241.050 ;
        RECT 271.950 240.600 274.050 241.050 ;
        RECT 169.950 239.400 274.050 240.600 ;
        RECT 169.950 238.950 172.050 239.400 ;
        RECT 190.950 238.950 193.050 239.400 ;
        RECT 271.950 238.950 274.050 239.400 ;
        RECT 34.950 237.600 37.050 238.050 ;
        RECT 43.950 237.600 46.050 238.050 ;
        RECT 34.950 236.400 46.050 237.600 ;
        RECT 34.950 235.950 37.050 236.400 ;
        RECT 43.950 235.950 46.050 236.400 ;
        RECT 73.950 237.600 76.050 238.050 ;
        RECT 88.950 237.600 91.050 238.050 ;
        RECT 73.950 236.400 91.050 237.600 ;
        RECT 73.950 235.950 76.050 236.400 ;
        RECT 88.950 235.950 91.050 236.400 ;
        RECT 103.950 237.600 106.050 238.050 ;
        RECT 142.950 237.600 145.050 238.050 ;
        RECT 103.950 236.400 145.050 237.600 ;
        RECT 103.950 235.950 106.050 236.400 ;
        RECT 142.950 235.950 145.050 236.400 ;
        RECT 160.950 237.600 163.050 238.050 ;
        RECT 226.950 237.600 229.050 238.050 ;
        RECT 160.950 236.400 229.050 237.600 ;
        RECT 160.950 235.950 163.050 236.400 ;
        RECT 226.950 235.950 229.050 236.400 ;
        RECT 313.950 234.600 316.050 235.050 ;
        RECT 358.950 234.600 361.050 235.050 ;
        RECT 313.950 233.400 361.050 234.600 ;
        RECT 313.950 232.950 316.050 233.400 ;
        RECT 358.950 232.950 361.050 233.400 ;
        RECT 55.950 231.600 58.050 232.050 ;
        RECT 76.950 231.600 79.050 232.050 ;
        RECT 55.950 230.400 79.050 231.600 ;
        RECT 55.950 229.950 58.050 230.400 ;
        RECT 76.950 229.950 79.050 230.400 ;
        RECT 130.950 231.600 133.050 232.050 ;
        RECT 139.950 231.600 142.050 232.050 ;
        RECT 130.950 230.400 142.050 231.600 ;
        RECT 130.950 229.950 133.050 230.400 ;
        RECT 139.950 229.950 142.050 230.400 ;
        RECT 307.950 231.600 310.050 232.050 ;
        RECT 325.950 231.600 328.050 232.050 ;
        RECT 307.950 230.400 328.050 231.600 ;
        RECT 307.950 229.950 310.050 230.400 ;
        RECT 325.950 229.950 328.050 230.400 ;
        RECT 43.950 228.600 46.050 229.050 ;
        RECT 82.950 228.600 85.050 229.050 ;
        RECT 43.950 227.400 85.050 228.600 ;
        RECT 43.950 226.950 46.050 227.400 ;
        RECT 82.950 226.950 85.050 227.400 ;
        RECT 100.950 228.600 103.050 229.050 ;
        RECT 148.950 228.600 151.050 229.050 ;
        RECT 100.950 227.400 151.050 228.600 ;
        RECT 100.950 226.950 103.050 227.400 ;
        RECT 148.950 226.950 151.050 227.400 ;
        RECT 205.950 228.600 208.050 229.050 ;
        RECT 238.950 228.600 241.050 229.050 ;
        RECT 205.950 227.400 241.050 228.600 ;
        RECT 205.950 226.950 208.050 227.400 ;
        RECT 238.950 226.950 241.050 227.400 ;
        RECT 271.950 228.600 274.050 229.050 ;
        RECT 295.950 228.600 298.050 229.050 ;
        RECT 271.950 227.400 298.050 228.600 ;
        RECT 271.950 226.950 274.050 227.400 ;
        RECT 295.950 226.950 298.050 227.400 ;
        RECT 73.950 225.600 76.050 226.050 ;
        RECT 103.950 225.600 106.050 226.050 ;
        RECT 73.950 224.400 106.050 225.600 ;
        RECT 73.950 223.950 76.050 224.400 ;
        RECT 103.950 223.950 106.050 224.400 ;
        RECT 328.950 225.600 331.050 226.050 ;
        RECT 340.950 225.600 343.050 226.050 ;
        RECT 328.950 224.400 343.050 225.600 ;
        RECT 328.950 223.950 331.050 224.400 ;
        RECT 340.950 223.950 343.050 224.400 ;
        RECT 37.950 222.600 40.050 223.050 ;
        RECT 106.950 222.600 109.050 223.050 ;
        RECT 112.950 222.600 115.050 223.050 ;
        RECT 145.950 222.600 148.050 223.050 ;
        RECT 37.950 221.400 60.600 222.600 ;
        RECT 37.950 220.950 40.050 221.400 ;
        RECT 16.950 219.600 19.050 220.050 ;
        RECT 16.950 218.400 27.600 219.600 ;
        RECT 16.950 217.950 19.050 218.400 ;
        RECT 7.950 216.600 10.050 217.200 ;
        RECT 5.400 215.400 10.050 216.600 ;
        RECT 5.400 211.050 6.600 215.400 ;
        RECT 7.950 215.100 10.050 215.400 ;
        RECT 4.950 208.950 7.050 211.050 ;
        RECT 26.400 210.600 27.600 218.400 ;
        RECT 55.950 215.100 58.050 217.200 ;
        RECT 28.950 213.600 31.050 214.050 ;
        RECT 56.400 213.600 57.600 215.100 ;
        RECT 28.950 212.400 57.600 213.600 ;
        RECT 28.950 211.950 31.050 212.400 ;
        RECT 34.950 210.600 37.050 210.900 ;
        RECT 26.400 209.400 37.050 210.600 ;
        RECT 34.950 208.800 37.050 209.400 ;
        RECT 49.950 210.600 52.050 211.050 ;
        RECT 56.400 210.600 57.600 212.400 ;
        RECT 59.400 210.900 60.600 221.400 ;
        RECT 106.950 221.400 148.050 222.600 ;
        RECT 106.950 220.950 109.050 221.400 ;
        RECT 112.950 220.950 115.050 221.400 ;
        RECT 145.950 220.950 148.050 221.400 ;
        RECT 226.950 222.600 229.050 223.050 ;
        RECT 262.950 222.600 265.050 223.050 ;
        RECT 226.950 221.400 265.050 222.600 ;
        RECT 226.950 220.950 229.050 221.400 ;
        RECT 262.950 220.950 265.050 221.400 ;
        RECT 277.950 222.600 280.050 223.050 ;
        RECT 301.950 222.600 304.050 223.050 ;
        RECT 352.950 222.600 355.050 223.050 ;
        RECT 277.950 221.400 304.050 222.600 ;
        RECT 277.950 220.950 280.050 221.400 ;
        RECT 75.000 219.600 79.050 220.050 ;
        RECT 74.400 217.950 79.050 219.600 ;
        RECT 64.950 214.800 67.050 216.900 ;
        RECT 49.950 209.400 57.600 210.600 ;
        RECT 49.950 208.950 52.050 209.400 ;
        RECT 58.950 208.800 61.050 210.900 ;
        RECT 65.400 208.050 66.600 214.800 ;
        RECT 61.950 206.400 66.600 208.050 ;
        RECT 74.400 208.050 75.600 217.950 ;
        RECT 91.800 215.100 93.900 217.200 ;
        RECT 94.950 216.600 97.050 217.050 ;
        RECT 127.950 216.750 130.050 217.200 ;
        RECT 133.950 216.750 136.050 217.200 ;
        RECT 94.950 215.400 105.600 216.600 ;
        RECT 92.400 210.600 93.600 215.100 ;
        RECT 94.950 214.950 97.050 215.400 ;
        RECT 104.400 210.900 105.600 215.400 ;
        RECT 127.950 215.550 136.050 216.750 ;
        RECT 148.950 216.600 151.050 220.050 ;
        RECT 187.950 219.600 190.050 220.050 ;
        RECT 199.950 219.600 202.050 220.050 ;
        RECT 187.950 218.400 202.050 219.600 ;
        RECT 187.950 217.950 190.050 218.400 ;
        RECT 199.950 217.950 202.050 218.400 ;
        RECT 241.950 219.600 244.050 220.050 ;
        RECT 259.950 219.600 262.050 220.050 ;
        RECT 241.950 218.400 262.050 219.600 ;
        RECT 241.950 217.950 244.050 218.400 ;
        RECT 259.950 217.950 262.050 218.400 ;
        RECT 166.950 216.600 169.050 217.050 ;
        RECT 178.950 216.600 181.050 217.200 ;
        RECT 208.950 216.600 211.050 217.200 ;
        RECT 148.950 216.000 153.600 216.600 ;
        RECT 127.950 215.100 130.050 215.550 ;
        RECT 133.950 215.100 136.050 215.550 ;
        RECT 149.400 215.400 153.600 216.000 ;
        RECT 152.400 213.600 153.600 215.400 ;
        RECT 166.950 215.400 181.050 216.600 ;
        RECT 166.950 214.950 169.050 215.400 ;
        RECT 178.950 215.100 181.050 215.400 ;
        RECT 200.400 215.400 211.050 216.600 ;
        RECT 140.400 212.400 153.600 213.600 ;
        RECT 97.950 210.600 100.050 210.900 ;
        RECT 92.400 209.400 100.050 210.600 ;
        RECT 97.950 208.800 100.050 209.400 ;
        RECT 103.950 208.800 106.050 210.900 ;
        RECT 140.400 208.050 141.600 212.400 ;
        RECT 74.400 206.400 79.050 208.050 ;
        RECT 61.950 205.950 66.000 206.400 ;
        RECT 75.000 205.950 79.050 206.400 ;
        RECT 127.950 207.600 130.050 208.050 ;
        RECT 133.950 207.600 136.050 208.050 ;
        RECT 127.950 206.400 136.050 207.600 ;
        RECT 127.950 205.950 130.050 206.400 ;
        RECT 133.950 205.950 136.050 206.400 ;
        RECT 139.950 205.950 142.050 208.050 ;
        RECT 152.400 207.600 153.600 212.400 ;
        RECT 181.950 210.600 184.050 210.900 ;
        RECT 196.950 210.600 199.050 210.900 ;
        RECT 200.400 210.600 201.600 215.400 ;
        RECT 208.950 215.100 211.050 215.400 ;
        RECT 214.950 214.950 217.050 217.050 ;
        RECT 220.950 214.950 223.050 217.050 ;
        RECT 253.950 215.100 256.050 217.200 ;
        RECT 215.400 211.050 216.600 214.950 ;
        RECT 205.950 210.600 208.050 211.050 ;
        RECT 181.950 209.400 208.050 210.600 ;
        RECT 181.950 208.800 184.050 209.400 ;
        RECT 196.950 208.800 199.050 209.400 ;
        RECT 205.950 208.950 208.050 209.400 ;
        RECT 214.950 208.950 217.050 211.050 ;
        RECT 221.400 210.600 222.600 214.950 ;
        RECT 229.950 210.600 232.050 211.050 ;
        RECT 221.400 209.400 232.050 210.600 ;
        RECT 229.950 208.950 232.050 209.400 ;
        RECT 244.950 210.600 247.050 210.900 ;
        RECT 254.400 210.600 255.600 215.100 ;
        RECT 265.950 214.950 268.050 217.050 ;
        RECT 289.950 216.600 292.050 217.200 ;
        RECT 284.400 215.400 292.050 216.600 ;
        RECT 266.400 211.050 267.600 214.950 ;
        RECT 284.400 211.050 285.600 215.400 ;
        RECT 289.950 215.100 292.050 215.400 ;
        RECT 244.950 209.400 255.600 210.600 ;
        RECT 244.950 208.800 247.050 209.400 ;
        RECT 265.950 208.950 268.050 211.050 ;
        RECT 283.950 208.950 286.050 211.050 ;
        RECT 293.400 210.900 294.600 221.400 ;
        RECT 301.950 220.950 304.050 221.400 ;
        RECT 314.400 221.400 355.050 222.600 ;
        RECT 295.950 215.100 298.050 217.200 ;
        RECT 306.000 216.600 310.050 217.050 ;
        RECT 292.950 208.800 295.050 210.900 ;
        RECT 157.950 207.600 160.050 208.050 ;
        RECT 152.400 206.400 160.050 207.600 ;
        RECT 157.950 205.950 160.050 206.400 ;
        RECT 211.950 207.600 214.050 208.050 ;
        RECT 238.950 207.600 241.050 208.050 ;
        RECT 256.950 207.600 259.050 208.050 ;
        RECT 280.950 207.600 283.050 208.050 ;
        RECT 211.950 206.400 283.050 207.600 ;
        RECT 296.400 207.600 297.600 215.100 ;
        RECT 305.400 214.950 310.050 216.600 ;
        RECT 305.400 210.900 306.600 214.950 ;
        RECT 314.400 210.900 315.600 221.400 ;
        RECT 352.950 220.950 355.050 221.400 ;
        RECT 358.950 219.600 361.050 220.050 ;
        RECT 329.400 218.400 361.050 219.600 ;
        RECT 304.950 208.800 307.050 210.900 ;
        RECT 313.950 208.800 316.050 210.900 ;
        RECT 329.400 208.050 330.600 218.400 ;
        RECT 358.950 217.950 361.050 218.400 ;
        RECT 346.950 214.950 349.050 217.050 ;
        RECT 343.950 210.600 346.050 210.900 ;
        RECT 347.400 210.600 348.600 214.950 ;
        RECT 355.950 210.600 358.050 210.900 ;
        RECT 343.950 209.400 358.050 210.600 ;
        RECT 343.950 208.800 346.050 209.400 ;
        RECT 355.950 208.800 358.050 209.400 ;
        RECT 301.950 207.600 304.050 208.050 ;
        RECT 296.400 206.400 304.050 207.600 ;
        RECT 211.950 205.950 214.050 206.400 ;
        RECT 238.950 205.950 241.050 206.400 ;
        RECT 256.950 205.950 259.050 206.400 ;
        RECT 280.950 205.950 283.050 206.400 ;
        RECT 301.950 205.950 304.050 206.400 ;
        RECT 328.950 205.950 331.050 208.050 ;
        RECT 4.950 204.600 7.050 205.050 ;
        RECT 19.950 204.600 22.050 205.050 ;
        RECT 52.950 204.600 55.050 205.050 ;
        RECT 88.950 204.600 91.050 205.050 ;
        RECT 148.950 204.600 151.050 205.050 ;
        RECT 154.950 204.600 157.050 205.050 ;
        RECT 4.950 203.400 60.600 204.600 ;
        RECT 4.950 202.950 7.050 203.400 ;
        RECT 19.950 202.950 22.050 203.400 ;
        RECT 52.950 202.950 55.050 203.400 ;
        RECT 28.950 201.600 31.050 202.050 ;
        RECT 40.950 201.600 43.050 202.050 ;
        RECT 28.950 200.400 43.050 201.600 ;
        RECT 59.400 201.600 60.600 203.400 ;
        RECT 88.950 203.400 126.600 204.600 ;
        RECT 88.950 202.950 91.050 203.400 ;
        RECT 64.950 201.600 67.050 202.050 ;
        RECT 59.400 200.400 67.050 201.600 ;
        RECT 125.400 201.600 126.600 203.400 ;
        RECT 148.950 203.400 157.050 204.600 ;
        RECT 148.950 202.950 151.050 203.400 ;
        RECT 154.950 202.950 157.050 203.400 ;
        RECT 187.950 204.600 190.050 205.050 ;
        RECT 217.950 204.600 220.050 205.050 ;
        RECT 187.950 203.400 220.050 204.600 ;
        RECT 187.950 202.950 190.050 203.400 ;
        RECT 217.950 202.950 220.050 203.400 ;
        RECT 136.950 201.600 139.050 202.050 ;
        RECT 125.400 200.400 139.050 201.600 ;
        RECT 28.950 199.950 31.050 200.400 ;
        RECT 40.950 199.950 43.050 200.400 ;
        RECT 64.950 199.950 67.050 200.400 ;
        RECT 136.950 199.950 139.050 200.400 ;
        RECT 157.950 201.600 160.050 202.050 ;
        RECT 187.950 201.600 190.050 201.900 ;
        RECT 157.950 200.400 190.050 201.600 ;
        RECT 157.950 199.950 160.050 200.400 ;
        RECT 187.950 199.800 190.050 200.400 ;
        RECT 199.950 201.600 202.050 202.050 ;
        RECT 214.950 201.600 217.050 202.050 ;
        RECT 199.950 200.400 217.050 201.600 ;
        RECT 199.950 199.950 202.050 200.400 ;
        RECT 214.950 199.950 217.050 200.400 ;
        RECT 229.950 201.600 232.050 202.050 ;
        RECT 274.950 201.600 277.050 202.050 ;
        RECT 229.950 200.400 277.050 201.600 ;
        RECT 229.950 199.950 232.050 200.400 ;
        RECT 274.950 199.950 277.050 200.400 ;
        RECT 280.950 201.600 283.050 202.050 ;
        RECT 304.950 201.600 307.050 202.050 ;
        RECT 280.950 200.400 307.050 201.600 ;
        RECT 280.950 199.950 283.050 200.400 ;
        RECT 304.950 199.950 307.050 200.400 ;
        RECT 313.950 201.600 316.050 202.050 ;
        RECT 346.950 201.600 349.050 202.050 ;
        RECT 313.950 200.400 349.050 201.600 ;
        RECT 313.950 199.950 316.050 200.400 ;
        RECT 346.950 199.950 349.050 200.400 ;
        RECT 1.950 198.600 4.050 199.050 ;
        RECT 10.950 198.600 13.050 199.050 ;
        RECT 1.950 197.400 13.050 198.600 ;
        RECT 1.950 196.950 4.050 197.400 ;
        RECT 10.950 196.950 13.050 197.400 ;
        RECT 205.950 198.600 208.050 199.050 ;
        RECT 268.950 198.600 271.050 199.050 ;
        RECT 205.950 197.400 271.050 198.600 ;
        RECT 205.950 196.950 208.050 197.400 ;
        RECT 268.950 196.950 271.050 197.400 ;
        RECT 283.950 198.600 286.050 199.050 ;
        RECT 325.950 198.600 328.050 199.050 ;
        RECT 283.950 197.400 328.050 198.600 ;
        RECT 283.950 196.950 286.050 197.400 ;
        RECT 325.950 196.950 328.050 197.400 ;
        RECT 205.950 195.600 208.050 195.900 ;
        RECT 223.950 195.600 226.050 196.050 ;
        RECT 205.950 194.400 226.050 195.600 ;
        RECT 205.950 193.800 208.050 194.400 ;
        RECT 223.950 193.950 226.050 194.400 ;
        RECT 292.950 195.600 295.050 196.050 ;
        RECT 331.950 195.600 334.050 196.050 ;
        RECT 292.950 194.400 334.050 195.600 ;
        RECT 292.950 193.950 295.050 194.400 ;
        RECT 331.950 193.950 334.050 194.400 ;
        RECT 52.950 192.600 55.050 193.050 ;
        RECT 94.950 192.600 97.050 193.050 ;
        RECT 52.950 191.400 97.050 192.600 ;
        RECT 52.950 190.950 55.050 191.400 ;
        RECT 94.950 190.950 97.050 191.400 ;
        RECT 103.950 192.600 106.050 193.050 ;
        RECT 118.950 192.600 121.050 193.050 ;
        RECT 103.950 191.400 121.050 192.600 ;
        RECT 103.950 190.950 106.050 191.400 ;
        RECT 118.950 190.950 121.050 191.400 ;
        RECT 130.950 192.600 133.050 193.050 ;
        RECT 139.950 192.600 142.050 193.050 ;
        RECT 130.950 191.400 142.050 192.600 ;
        RECT 130.950 190.950 133.050 191.400 ;
        RECT 139.950 190.950 142.050 191.400 ;
        RECT 154.950 192.600 157.050 193.050 ;
        RECT 172.950 192.600 175.050 193.050 ;
        RECT 154.950 191.400 175.050 192.600 ;
        RECT 154.950 190.950 157.050 191.400 ;
        RECT 172.950 190.950 175.050 191.400 ;
        RECT 301.950 192.600 304.050 193.050 ;
        RECT 349.950 192.600 352.050 193.050 ;
        RECT 301.950 191.400 352.050 192.600 ;
        RECT 301.950 190.950 304.050 191.400 ;
        RECT 349.950 190.950 352.050 191.400 ;
        RECT 1.950 189.600 4.050 190.050 ;
        RECT 49.950 189.600 52.050 190.050 ;
        RECT 1.950 188.400 52.050 189.600 ;
        RECT 1.950 187.950 4.050 188.400 ;
        RECT 49.950 187.950 52.050 188.400 ;
        RECT 61.950 189.600 64.050 190.050 ;
        RECT 67.950 189.600 70.050 190.050 ;
        RECT 61.950 188.400 70.050 189.600 ;
        RECT 61.950 187.950 64.050 188.400 ;
        RECT 67.950 187.950 70.050 188.400 ;
        RECT 109.950 189.600 112.050 190.050 ;
        RECT 115.950 189.600 118.050 190.050 ;
        RECT 109.950 188.400 118.050 189.600 ;
        RECT 109.950 187.950 112.050 188.400 ;
        RECT 115.950 187.950 118.050 188.400 ;
        RECT 139.950 189.600 142.050 189.900 ;
        RECT 166.950 189.600 169.050 190.050 ;
        RECT 139.950 188.400 169.050 189.600 ;
        RECT 139.950 187.800 142.050 188.400 ;
        RECT 166.950 187.950 169.050 188.400 ;
        RECT 265.950 189.600 268.050 190.050 ;
        RECT 277.950 189.600 280.050 190.050 ;
        RECT 265.950 188.400 280.050 189.600 ;
        RECT 265.950 187.950 268.050 188.400 ;
        RECT 277.950 187.950 280.050 188.400 ;
        RECT 304.950 189.600 307.050 190.050 ;
        RECT 340.950 189.600 343.050 190.050 ;
        RECT 304.950 188.400 343.050 189.600 ;
        RECT 304.950 187.950 307.050 188.400 ;
        RECT 340.950 187.950 343.050 188.400 ;
        RECT 103.800 184.950 105.900 187.050 ;
        RECT 118.950 186.600 121.050 187.050 ;
        RECT 127.950 186.600 130.050 187.050 ;
        RECT 118.950 185.400 130.050 186.600 ;
        RECT 118.950 184.950 121.050 185.400 ;
        RECT 127.950 184.950 130.050 185.400 ;
        RECT 205.950 186.600 208.050 187.050 ;
        RECT 262.950 186.600 265.050 187.050 ;
        RECT 268.950 186.600 271.050 187.050 ;
        RECT 205.950 185.400 222.600 186.600 ;
        RECT 205.950 184.950 208.050 185.400 ;
        RECT 67.950 183.750 70.050 184.200 ;
        RECT 79.950 183.750 82.050 184.200 ;
        RECT 67.950 182.550 82.050 183.750 ;
        RECT 67.950 182.100 70.050 182.550 ;
        RECT 79.950 182.100 82.050 182.550 ;
        RECT 85.950 183.600 88.050 184.200 ;
        RECT 85.950 182.400 93.600 183.600 ;
        RECT 85.950 182.100 88.050 182.400 ;
        RECT 1.950 178.950 4.050 181.050 ;
        RECT 28.950 180.450 31.050 180.900 ;
        RECT 52.800 180.450 54.900 180.900 ;
        RECT 28.950 179.250 54.900 180.450 ;
        RECT 2.400 175.050 3.600 178.950 ;
        RECT 28.950 178.800 31.050 179.250 ;
        RECT 52.800 178.800 54.900 179.250 ;
        RECT 64.950 179.100 67.050 181.200 ;
        RECT 49.950 177.600 52.050 178.050 ;
        RECT 65.400 177.600 66.600 179.100 ;
        RECT 88.950 177.600 91.050 178.050 ;
        RECT 49.950 176.400 91.050 177.600 ;
        RECT 92.400 177.600 93.600 182.400 ;
        RECT 104.250 177.900 105.450 184.950 ;
        RECT 121.950 181.950 124.050 184.050 ;
        RECT 133.950 181.950 136.050 184.050 ;
        RECT 139.950 183.600 142.050 184.200 ;
        RECT 137.400 182.400 142.050 183.600 ;
        RECT 122.400 178.050 123.600 181.950 ;
        RECT 97.950 177.600 100.050 177.900 ;
        RECT 92.400 176.400 100.050 177.600 ;
        RECT 49.950 175.950 52.050 176.400 ;
        RECT 88.950 175.950 91.050 176.400 ;
        RECT 97.950 175.800 100.050 176.400 ;
        RECT 103.800 175.800 105.900 177.900 ;
        RECT 121.950 175.950 124.050 178.050 ;
        RECT 1.950 172.950 4.050 175.050 ;
        RECT 73.950 174.600 76.050 175.050 ;
        RECT 91.950 174.600 94.050 175.050 ;
        RECT 73.950 173.400 94.050 174.600 ;
        RECT 73.950 172.950 76.050 173.400 ;
        RECT 91.950 172.950 94.050 173.400 ;
        RECT 127.950 174.600 130.050 175.050 ;
        RECT 134.400 174.600 135.600 181.950 ;
        RECT 137.400 175.050 138.600 182.400 ;
        RECT 139.950 182.100 142.050 182.400 ;
        RECT 148.950 182.100 151.050 184.200 ;
        RECT 172.950 183.600 175.050 184.200 ;
        RECT 161.400 182.400 175.050 183.600 ;
        RECT 149.400 175.050 150.600 182.100 ;
        RECT 161.400 180.600 162.600 182.400 ;
        RECT 172.950 182.100 175.050 182.400 ;
        RECT 199.950 180.600 202.050 181.050 ;
        RECT 221.400 180.900 222.600 185.400 ;
        RECT 262.950 185.400 271.050 186.600 ;
        RECT 262.950 184.950 265.050 185.400 ;
        RECT 268.950 184.950 271.050 185.400 ;
        RECT 296.400 185.400 303.600 186.600 ;
        RECT 286.950 181.950 289.050 184.050 ;
        RECT 158.400 179.400 162.600 180.600 ;
        RECT 188.400 179.400 202.050 180.600 ;
        RECT 158.400 177.900 159.600 179.400 ;
        RECT 157.950 175.800 160.050 177.900 ;
        RECT 188.400 175.050 189.600 179.400 ;
        RECT 199.950 178.950 202.050 179.400 ;
        RECT 220.950 178.800 223.050 180.900 ;
        RECT 287.400 178.050 288.600 181.950 ;
        RECT 271.950 177.450 274.050 177.900 ;
        RECT 277.950 177.450 280.050 177.900 ;
        RECT 271.950 176.250 280.050 177.450 ;
        RECT 271.950 175.800 274.050 176.250 ;
        RECT 277.950 175.800 280.050 176.250 ;
        RECT 286.950 175.950 289.050 178.050 ;
        RECT 127.950 173.400 135.600 174.600 ;
        RECT 127.950 172.950 130.050 173.400 ;
        RECT 136.950 172.950 139.050 175.050 ;
        RECT 145.950 173.400 150.600 175.050 ;
        RECT 145.950 172.950 150.000 173.400 ;
        RECT 187.950 172.950 190.050 175.050 ;
        RECT 296.400 174.600 297.600 185.400 ;
        RECT 298.950 182.100 301.050 184.200 ;
        RECT 302.400 183.600 303.600 185.400 ;
        RECT 331.950 184.950 334.050 187.050 ;
        RECT 304.950 183.600 307.050 184.200 ;
        RECT 319.950 183.600 322.050 184.200 ;
        RECT 328.950 183.600 331.050 184.200 ;
        RECT 302.400 182.400 307.050 183.600 ;
        RECT 304.950 182.100 307.050 182.400 ;
        RECT 308.400 182.400 322.050 183.600 ;
        RECT 299.400 177.600 300.600 182.100 ;
        RECT 308.400 177.900 309.600 182.400 ;
        RECT 319.950 182.100 322.050 182.400 ;
        RECT 323.400 182.400 331.050 183.600 ;
        RECT 323.400 177.900 324.600 182.400 ;
        RECT 328.950 182.100 331.050 182.400 ;
        RECT 332.400 177.900 333.600 184.950 ;
        RECT 299.400 176.400 303.600 177.600 ;
        RECT 296.400 174.000 300.600 174.600 ;
        RECT 296.400 173.400 301.050 174.000 ;
        RECT 118.950 171.600 121.050 172.050 ;
        RECT 65.400 170.400 121.050 171.600 ;
        RECT 28.950 168.600 31.050 169.050 ;
        RECT 65.400 168.600 66.600 170.400 ;
        RECT 118.950 169.950 121.050 170.400 ;
        RECT 157.950 171.600 160.050 172.050 ;
        RECT 184.950 171.600 187.050 172.050 ;
        RECT 157.950 170.400 187.050 171.600 ;
        RECT 157.950 169.950 160.050 170.400 ;
        RECT 184.950 169.950 187.050 170.400 ;
        RECT 298.950 169.950 301.050 173.400 ;
        RECT 302.400 171.600 303.600 176.400 ;
        RECT 307.950 175.800 310.050 177.900 ;
        RECT 322.950 175.800 325.050 177.900 ;
        RECT 331.950 175.800 334.050 177.900 ;
        RECT 316.950 171.600 319.050 172.050 ;
        RECT 302.400 170.400 319.050 171.600 ;
        RECT 316.950 169.950 319.050 170.400 ;
        RECT 28.950 167.400 66.600 168.600 ;
        RECT 88.950 168.600 91.050 169.050 ;
        RECT 109.950 168.600 112.050 169.050 ;
        RECT 88.950 167.400 112.050 168.600 ;
        RECT 28.950 166.950 31.050 167.400 ;
        RECT 88.950 166.950 91.050 167.400 ;
        RECT 109.950 166.950 112.050 167.400 ;
        RECT 271.950 168.600 274.050 169.050 ;
        RECT 295.950 168.600 298.050 169.050 ;
        RECT 271.950 167.400 298.050 168.600 ;
        RECT 271.950 166.950 274.050 167.400 ;
        RECT 295.950 166.950 298.050 167.400 ;
        RECT 127.950 165.600 130.050 166.050 ;
        RECT 154.950 165.600 157.050 166.050 ;
        RECT 127.950 164.400 157.050 165.600 ;
        RECT 127.950 163.950 130.050 164.400 ;
        RECT 154.950 163.950 157.050 164.400 ;
        RECT 265.950 162.600 268.050 163.050 ;
        RECT 316.950 162.600 319.050 163.050 ;
        RECT 265.950 161.400 319.050 162.600 ;
        RECT 265.950 160.950 268.050 161.400 ;
        RECT 316.950 160.950 319.050 161.400 ;
        RECT 1.950 156.600 4.050 157.050 ;
        RECT 13.950 156.600 16.050 157.050 ;
        RECT 1.950 155.400 16.050 156.600 ;
        RECT 1.950 154.950 4.050 155.400 ;
        RECT 13.950 154.950 16.050 155.400 ;
        RECT 118.950 156.600 121.050 157.050 ;
        RECT 127.950 156.600 130.050 157.050 ;
        RECT 118.950 155.400 130.050 156.600 ;
        RECT 118.950 154.950 121.050 155.400 ;
        RECT 127.950 154.950 130.050 155.400 ;
        RECT 139.950 156.600 142.050 157.050 ;
        RECT 160.950 156.600 163.050 157.050 ;
        RECT 175.950 156.600 178.050 157.050 ;
        RECT 223.950 156.600 226.050 157.050 ;
        RECT 139.950 155.400 226.050 156.600 ;
        RECT 139.950 154.950 142.050 155.400 ;
        RECT 160.950 154.950 163.050 155.400 ;
        RECT 175.950 154.950 178.050 155.400 ;
        RECT 223.950 154.950 226.050 155.400 ;
        RECT 232.950 156.600 235.050 157.050 ;
        RECT 277.950 156.600 280.050 157.050 ;
        RECT 232.950 155.400 280.050 156.600 ;
        RECT 232.950 154.950 235.050 155.400 ;
        RECT 277.950 154.950 280.050 155.400 ;
        RECT 322.950 156.600 325.050 157.050 ;
        RECT 346.950 156.600 349.050 157.050 ;
        RECT 322.950 155.400 349.050 156.600 ;
        RECT 322.950 154.950 325.050 155.400 ;
        RECT 346.950 154.950 349.050 155.400 ;
        RECT 91.950 153.600 94.050 154.050 ;
        RECT 130.950 153.600 133.050 154.050 ;
        RECT 91.950 152.400 133.050 153.600 ;
        RECT 224.400 153.600 225.600 154.950 ;
        RECT 241.950 153.600 244.050 154.050 ;
        RECT 224.400 152.400 244.050 153.600 ;
        RECT 91.950 151.950 94.050 152.400 ;
        RECT 130.950 151.950 133.050 152.400 ;
        RECT 241.950 151.950 244.050 152.400 ;
        RECT 13.950 147.600 16.050 148.050 ;
        RECT 73.950 147.600 76.050 148.050 ;
        RECT 13.950 146.400 76.050 147.600 ;
        RECT 13.950 145.950 16.050 146.400 ;
        RECT 73.950 145.950 76.050 146.400 ;
        RECT 97.950 147.600 100.050 148.050 ;
        RECT 118.950 147.600 121.050 148.050 ;
        RECT 97.950 146.400 121.050 147.600 ;
        RECT 97.950 145.950 100.050 146.400 ;
        RECT 118.950 145.950 121.050 146.400 ;
        RECT 241.950 147.600 244.050 148.050 ;
        RECT 280.950 147.600 283.050 148.050 ;
        RECT 241.950 146.400 283.050 147.600 ;
        RECT 241.950 145.950 244.050 146.400 ;
        RECT 280.950 145.950 283.050 146.400 ;
        RECT 106.950 144.600 109.050 145.050 ;
        RECT 130.950 144.600 133.050 145.050 ;
        RECT 139.950 144.600 142.050 145.050 ;
        RECT 106.950 143.400 117.600 144.600 ;
        RECT 106.950 142.950 109.050 143.400 ;
        RECT 79.950 141.600 82.050 142.050 ;
        RECT 112.950 141.600 115.050 142.050 ;
        RECT 79.950 140.400 115.050 141.600 ;
        RECT 116.400 141.600 117.600 143.400 ;
        RECT 130.950 143.400 142.050 144.600 ;
        RECT 130.950 142.950 133.050 143.400 ;
        RECT 139.950 142.950 142.050 143.400 ;
        RECT 175.950 144.600 178.050 145.050 ;
        RECT 202.950 144.600 205.050 145.050 ;
        RECT 208.950 144.600 211.050 145.050 ;
        RECT 175.950 143.400 211.050 144.600 ;
        RECT 175.950 142.950 178.050 143.400 ;
        RECT 202.950 142.950 205.050 143.400 ;
        RECT 208.950 142.950 211.050 143.400 ;
        RECT 253.950 144.600 256.050 145.050 ;
        RECT 274.950 144.600 277.050 145.050 ;
        RECT 253.950 143.400 277.050 144.600 ;
        RECT 253.950 142.950 256.050 143.400 ;
        RECT 274.950 142.950 277.050 143.400 ;
        RECT 295.950 144.600 300.000 145.050 ;
        RECT 295.950 142.950 300.600 144.600 ;
        RECT 127.950 141.600 130.050 142.050 ;
        RECT 145.950 141.600 148.050 142.050 ;
        RECT 116.400 140.400 126.600 141.600 ;
        RECT 79.950 139.950 82.050 140.400 ;
        RECT 112.950 139.950 115.050 140.400 ;
        RECT 28.950 138.600 31.050 139.050 ;
        RECT 28.950 138.000 54.600 138.600 ;
        RECT 28.950 137.400 55.050 138.000 ;
        RECT 28.950 136.950 31.050 137.400 ;
        RECT 25.950 133.950 28.050 136.050 ;
        RECT 52.950 133.950 55.050 137.400 ;
        RECT 73.950 137.100 76.050 139.200 ;
        RECT 79.950 137.100 82.050 139.200 ;
        RECT 91.950 137.100 94.050 139.200 ;
        RECT 117.000 138.600 121.050 139.050 ;
        RECT 64.950 135.600 67.050 135.900 ;
        RECT 74.400 135.600 75.600 137.100 ;
        RECT 64.950 134.400 75.600 135.600 ;
        RECT 26.400 126.600 27.600 133.950 ;
        RECT 64.950 133.800 67.050 134.400 ;
        RECT 80.400 132.600 81.600 137.100 ;
        RECT 85.950 132.600 88.050 133.050 ;
        RECT 80.400 131.400 88.050 132.600 ;
        RECT 92.400 132.600 93.600 137.100 ;
        RECT 116.400 136.950 121.050 138.600 ;
        RECT 109.950 132.600 112.050 132.900 ;
        RECT 116.400 132.600 117.600 136.950 ;
        RECT 125.400 132.900 126.600 140.400 ;
        RECT 127.950 140.400 148.050 141.600 ;
        RECT 299.400 141.600 300.600 142.950 ;
        RECT 349.950 141.600 352.050 142.050 ;
        RECT 355.950 141.600 358.050 142.050 ;
        RECT 299.400 140.400 358.050 141.600 ;
        RECT 127.950 139.950 130.050 140.400 ;
        RECT 145.950 139.950 148.050 140.400 ;
        RECT 349.950 139.950 352.050 140.400 ;
        RECT 355.950 139.950 358.050 140.400 ;
        RECT 154.950 138.600 157.050 139.200 ;
        RECT 159.000 138.600 163.050 139.050 ;
        RECT 131.400 137.400 157.050 138.600 ;
        RECT 92.400 132.000 99.600 132.600 ;
        RECT 92.400 131.400 100.050 132.000 ;
        RECT 85.950 130.950 88.050 131.400 ;
        RECT 70.950 129.600 73.050 130.050 ;
        RECT 91.950 129.600 94.050 130.050 ;
        RECT 70.950 128.400 94.050 129.600 ;
        RECT 70.950 127.950 73.050 128.400 ;
        RECT 91.950 127.950 94.050 128.400 ;
        RECT 97.950 127.950 100.050 131.400 ;
        RECT 109.950 131.400 117.600 132.600 ;
        RECT 109.950 130.800 112.050 131.400 ;
        RECT 124.950 130.800 127.050 132.900 ;
        RECT 115.950 129.600 118.050 130.050 ;
        RECT 131.400 129.600 132.600 137.400 ;
        RECT 154.950 137.100 157.050 137.400 ;
        RECT 158.400 136.950 163.050 138.600 ;
        RECT 169.950 138.600 172.050 139.200 ;
        RECT 175.950 138.600 178.050 139.200 ;
        RECT 190.950 138.600 193.050 139.200 ;
        RECT 169.950 137.400 178.050 138.600 ;
        RECT 169.950 137.100 172.050 137.400 ;
        RECT 175.950 137.100 178.050 137.400 ;
        RECT 179.400 137.400 193.050 138.600 ;
        RECT 158.400 132.900 159.600 136.950 ;
        RECT 179.400 135.600 180.600 137.400 ;
        RECT 190.950 137.100 193.050 137.400 ;
        RECT 199.950 137.100 202.050 139.200 ;
        RECT 164.400 135.000 180.600 135.600 ;
        RECT 163.950 134.400 180.600 135.000 ;
        RECT 157.950 130.800 160.050 132.900 ;
        RECT 163.950 130.950 166.050 134.400 ;
        RECT 200.400 132.600 201.600 137.100 ;
        RECT 232.950 136.950 235.050 139.050 ;
        RECT 241.950 138.600 244.050 139.200 ;
        RECT 253.950 138.600 256.050 139.200 ;
        RECT 241.950 137.400 256.050 138.600 ;
        RECT 241.950 137.100 244.050 137.400 ;
        RECT 253.950 137.100 256.050 137.400 ;
        RECT 265.950 137.100 268.050 139.200 ;
        RECT 205.950 132.600 208.050 133.050 ;
        RECT 200.400 131.400 208.050 132.600 ;
        RECT 233.400 132.600 234.600 136.950 ;
        RECT 238.950 132.600 241.050 132.900 ;
        RECT 233.400 131.400 241.050 132.600 ;
        RECT 205.950 130.950 208.050 131.400 ;
        RECT 238.950 130.800 241.050 131.400 ;
        RECT 256.950 132.600 259.050 132.900 ;
        RECT 266.400 132.600 267.600 137.100 ;
        RECT 316.950 134.100 319.050 136.200 ;
        RECT 256.950 131.400 267.600 132.600 ;
        RECT 268.950 132.600 271.050 132.900 ;
        RECT 280.950 132.600 283.050 132.900 ;
        RECT 268.950 131.400 283.050 132.600 ;
        RECT 256.950 130.800 259.050 131.400 ;
        RECT 268.950 130.800 271.050 131.400 ;
        RECT 280.950 130.800 283.050 131.400 ;
        RECT 286.950 132.600 289.050 132.900 ;
        RECT 317.400 132.600 318.600 134.100 ;
        RECT 286.950 131.400 318.600 132.600 ;
        RECT 286.950 130.800 289.050 131.400 ;
        RECT 115.950 128.400 132.600 129.600 ;
        RECT 157.950 129.600 160.050 130.050 ;
        RECT 166.950 129.600 169.050 130.050 ;
        RECT 157.950 128.400 169.050 129.600 ;
        RECT 115.950 127.950 118.050 128.400 ;
        RECT 157.950 127.950 160.050 128.400 ;
        RECT 166.950 127.950 169.050 128.400 ;
        RECT 88.950 126.600 91.050 127.050 ;
        RECT 26.400 125.400 91.050 126.600 ;
        RECT 88.950 124.950 91.050 125.400 ;
        RECT 145.950 126.600 148.050 127.050 ;
        RECT 158.400 126.600 159.600 127.950 ;
        RECT 145.950 125.400 159.600 126.600 ;
        RECT 178.950 126.600 181.050 127.050 ;
        RECT 193.950 126.600 196.050 127.050 ;
        RECT 178.950 125.400 196.050 126.600 ;
        RECT 145.950 124.950 148.050 125.400 ;
        RECT 178.950 124.950 181.050 125.400 ;
        RECT 193.950 124.950 196.050 125.400 ;
        RECT 52.950 123.600 55.050 124.050 ;
        RECT 17.400 122.400 55.050 123.600 ;
        RECT 4.950 120.600 7.050 121.050 ;
        RECT 17.400 120.600 18.600 122.400 ;
        RECT 52.950 121.950 55.050 122.400 ;
        RECT 58.950 123.600 61.050 124.050 ;
        RECT 64.950 123.600 67.050 124.050 ;
        RECT 58.950 122.400 67.050 123.600 ;
        RECT 58.950 121.950 61.050 122.400 ;
        RECT 64.950 121.950 67.050 122.400 ;
        RECT 97.950 123.600 100.050 124.050 ;
        RECT 103.950 123.600 106.050 124.050 ;
        RECT 97.950 122.400 106.050 123.600 ;
        RECT 97.950 121.950 100.050 122.400 ;
        RECT 103.950 121.950 106.050 122.400 ;
        RECT 121.950 123.600 124.050 124.050 ;
        RECT 139.950 123.600 142.050 124.050 ;
        RECT 121.950 122.400 142.050 123.600 ;
        RECT 121.950 121.950 124.050 122.400 ;
        RECT 139.950 121.950 142.050 122.400 ;
        RECT 4.950 119.400 18.600 120.600 ;
        RECT 112.950 120.600 115.050 121.050 ;
        RECT 133.950 120.600 136.050 121.050 ;
        RECT 112.950 119.400 136.050 120.600 ;
        RECT 4.950 118.950 7.050 119.400 ;
        RECT 112.950 118.950 115.050 119.400 ;
        RECT 133.950 118.950 136.050 119.400 ;
        RECT 157.950 120.600 160.050 121.050 ;
        RECT 184.950 120.600 187.050 121.050 ;
        RECT 157.950 119.400 187.050 120.600 ;
        RECT 157.950 118.950 160.050 119.400 ;
        RECT 184.950 118.950 187.050 119.400 ;
        RECT 25.950 117.600 28.050 118.050 ;
        RECT 49.950 117.600 52.050 118.050 ;
        RECT 25.950 116.400 52.050 117.600 ;
        RECT 25.950 115.950 28.050 116.400 ;
        RECT 49.950 115.950 52.050 116.400 ;
        RECT 76.950 117.600 79.050 118.050 ;
        RECT 97.950 117.600 100.050 118.050 ;
        RECT 76.950 116.400 100.050 117.600 ;
        RECT 76.950 115.950 79.050 116.400 ;
        RECT 97.950 115.950 100.050 116.400 ;
        RECT 301.950 117.600 304.050 118.050 ;
        RECT 310.950 117.600 313.050 118.050 ;
        RECT 301.950 116.400 313.050 117.600 ;
        RECT 301.950 115.950 304.050 116.400 ;
        RECT 310.950 115.950 313.050 116.400 ;
        RECT 13.950 114.600 16.050 115.050 ;
        RECT 37.950 114.600 40.050 115.050 ;
        RECT 58.950 114.600 61.050 115.050 ;
        RECT 85.950 114.600 88.050 115.050 ;
        RECT 13.950 113.400 61.050 114.600 ;
        RECT 13.950 112.950 16.050 113.400 ;
        RECT 37.950 112.950 40.050 113.400 ;
        RECT 58.950 112.950 61.050 113.400 ;
        RECT 65.400 113.400 88.050 114.600 ;
        RECT 16.950 111.600 19.050 112.050 ;
        RECT 31.950 111.600 34.050 112.050 ;
        RECT 16.950 110.400 34.050 111.600 ;
        RECT 16.950 109.950 19.050 110.400 ;
        RECT 31.950 109.950 34.050 110.400 ;
        RECT 46.950 111.600 49.050 112.050 ;
        RECT 65.400 111.600 66.600 113.400 ;
        RECT 85.950 112.950 88.050 113.400 ;
        RECT 154.950 114.600 157.050 115.050 ;
        RECT 169.950 114.600 172.050 115.050 ;
        RECT 154.950 113.400 172.050 114.600 ;
        RECT 154.950 112.950 157.050 113.400 ;
        RECT 169.950 112.950 172.050 113.400 ;
        RECT 325.950 114.600 328.050 115.050 ;
        RECT 337.950 114.600 340.050 115.050 ;
        RECT 346.950 114.600 349.050 115.050 ;
        RECT 325.950 113.400 349.050 114.600 ;
        RECT 325.950 112.950 328.050 113.400 ;
        RECT 337.950 112.950 340.050 113.400 ;
        RECT 346.950 112.950 349.050 113.400 ;
        RECT 46.950 110.400 66.600 111.600 ;
        RECT 103.950 111.600 106.050 112.050 ;
        RECT 115.950 111.600 118.050 112.050 ;
        RECT 103.950 110.400 118.050 111.600 ;
        RECT 46.950 109.950 49.050 110.400 ;
        RECT 103.950 109.950 106.050 110.400 ;
        RECT 115.950 109.950 118.050 110.400 ;
        RECT 172.950 111.600 175.050 112.050 ;
        RECT 202.950 111.600 205.050 112.050 ;
        RECT 250.950 111.600 253.050 112.050 ;
        RECT 172.950 110.400 253.050 111.600 ;
        RECT 172.950 109.950 175.050 110.400 ;
        RECT 202.950 109.950 205.050 110.400 ;
        RECT 250.950 109.950 253.050 110.400 ;
        RECT 70.950 106.950 73.050 109.050 ;
        RECT 97.950 108.600 100.050 109.050 ;
        RECT 112.950 108.600 115.050 109.050 ;
        RECT 97.950 107.400 115.050 108.600 ;
        RECT 97.950 106.950 100.050 107.400 ;
        RECT 112.950 106.950 115.050 107.400 ;
        RECT 169.950 108.600 172.050 109.050 ;
        RECT 199.950 108.600 202.050 109.050 ;
        RECT 210.000 108.600 214.050 109.050 ;
        RECT 169.950 107.400 202.050 108.600 ;
        RECT 169.950 106.950 172.050 107.400 ;
        RECT 199.950 106.950 202.050 107.400 ;
        RECT 209.400 106.950 214.050 108.600 ;
        RECT 25.950 104.100 28.050 106.200 ;
        RECT 45.000 105.600 49.050 106.050 ;
        RECT 26.400 99.600 27.600 104.100 ;
        RECT 44.400 103.950 49.050 105.600 ;
        RECT 34.950 99.600 37.050 99.900 ;
        RECT 26.400 98.400 37.050 99.600 ;
        RECT 34.950 97.800 37.050 98.400 ;
        RECT 40.950 99.600 43.050 99.900 ;
        RECT 44.400 99.600 45.600 103.950 ;
        RECT 71.400 99.900 72.600 106.950 ;
        RECT 73.950 105.600 76.050 106.200 ;
        RECT 91.950 105.600 94.050 106.200 ;
        RECT 73.950 104.400 94.050 105.600 ;
        RECT 73.950 104.100 76.050 104.400 ;
        RECT 91.950 104.100 94.050 104.400 ;
        RECT 163.950 105.600 166.050 106.050 ;
        RECT 190.950 105.600 195.000 106.050 ;
        RECT 163.950 104.400 189.600 105.600 ;
        RECT 92.400 102.600 93.600 104.100 ;
        RECT 163.950 103.950 166.050 104.400 ;
        RECT 89.400 101.400 93.600 102.600 ;
        RECT 133.950 102.450 136.050 102.900 ;
        RECT 157.950 102.450 160.050 102.900 ;
        RECT 40.950 98.400 45.600 99.600 ;
        RECT 61.950 99.600 64.050 99.900 ;
        RECT 70.950 99.600 73.050 99.900 ;
        RECT 61.950 98.400 73.050 99.600 ;
        RECT 40.950 97.800 43.050 98.400 ;
        RECT 61.950 97.800 64.050 98.400 ;
        RECT 70.950 97.800 73.050 98.400 ;
        RECT 82.950 99.600 85.050 99.900 ;
        RECT 89.400 99.600 90.600 101.400 ;
        RECT 133.950 101.250 160.050 102.450 ;
        RECT 133.950 100.800 136.050 101.250 ;
        RECT 157.950 100.800 160.050 101.250 ;
        RECT 163.950 102.750 166.050 102.900 ;
        RECT 169.950 102.750 172.050 103.200 ;
        RECT 163.950 101.550 172.050 102.750 ;
        RECT 163.950 100.800 166.050 101.550 ;
        RECT 169.950 101.100 172.050 101.550 ;
        RECT 188.400 99.900 189.600 104.400 ;
        RECT 190.950 103.950 195.600 105.600 ;
        RECT 194.400 100.050 195.600 103.950 ;
        RECT 209.400 100.050 210.600 106.950 ;
        RECT 214.950 104.100 217.050 106.200 ;
        RECT 229.950 105.600 232.050 106.200 ;
        RECT 256.950 105.600 259.050 106.200 ;
        RECT 229.950 104.400 237.600 105.600 ;
        RECT 229.950 104.100 232.050 104.400 ;
        RECT 82.950 98.400 90.600 99.600 ;
        RECT 82.950 97.800 85.050 98.400 ;
        RECT 187.950 97.800 190.050 99.900 ;
        RECT 193.950 97.950 196.050 100.050 ;
        RECT 208.950 97.950 211.050 100.050 ;
        RECT 215.400 99.600 216.600 104.100 ;
        RECT 236.400 100.050 237.600 104.400 ;
        RECT 248.400 104.400 259.050 105.600 ;
        RECT 248.400 100.050 249.600 104.400 ;
        RECT 256.950 104.100 259.050 104.400 ;
        RECT 289.950 102.450 292.050 102.900 ;
        RECT 310.950 102.450 313.050 102.900 ;
        RECT 289.950 101.250 313.050 102.450 ;
        RECT 289.950 100.800 292.050 101.250 ;
        RECT 310.950 100.800 313.050 101.250 ;
        RECT 226.950 99.600 229.050 99.900 ;
        RECT 212.400 98.400 229.050 99.600 ;
        RECT 202.950 96.600 205.050 97.050 ;
        RECT 212.400 96.600 213.600 98.400 ;
        RECT 226.950 97.800 229.050 98.400 ;
        RECT 235.950 97.950 238.050 100.050 ;
        RECT 247.950 97.950 250.050 100.050 ;
        RECT 202.950 95.400 213.600 96.600 ;
        RECT 202.950 94.950 205.050 95.400 ;
        RECT 52.950 93.600 55.050 94.050 ;
        RECT 64.950 93.600 67.050 94.050 ;
        RECT 52.950 92.400 67.050 93.600 ;
        RECT 52.950 91.950 55.050 92.400 ;
        RECT 64.950 91.950 67.050 92.400 ;
        RECT 175.950 93.600 178.050 94.050 ;
        RECT 193.950 93.600 196.050 94.050 ;
        RECT 217.950 93.600 220.050 94.050 ;
        RECT 229.950 93.600 232.050 94.050 ;
        RECT 175.950 92.400 232.050 93.600 ;
        RECT 175.950 91.950 178.050 92.400 ;
        RECT 193.950 91.950 196.050 92.400 ;
        RECT 217.950 91.950 220.050 92.400 ;
        RECT 229.950 91.950 232.050 92.400 ;
        RECT 235.950 93.600 238.050 94.050 ;
        RECT 259.950 93.600 262.050 94.050 ;
        RECT 235.950 92.400 262.050 93.600 ;
        RECT 235.950 91.950 238.050 92.400 ;
        RECT 259.950 91.950 262.050 92.400 ;
        RECT 253.950 90.600 256.050 91.050 ;
        RECT 259.950 90.600 262.050 90.900 ;
        RECT 253.950 89.400 262.050 90.600 ;
        RECT 253.950 88.950 256.050 89.400 ;
        RECT 259.950 88.800 262.050 89.400 ;
        RECT 25.950 87.600 28.050 88.050 ;
        RECT 94.950 87.600 97.050 88.050 ;
        RECT 25.950 86.400 97.050 87.600 ;
        RECT 25.950 85.950 28.050 86.400 ;
        RECT 94.950 85.950 97.050 86.400 ;
        RECT 103.950 87.600 106.050 88.050 ;
        RECT 196.950 87.600 199.050 88.050 ;
        RECT 103.950 86.400 199.050 87.600 ;
        RECT 103.950 85.950 106.050 86.400 ;
        RECT 196.950 85.950 199.050 86.400 ;
        RECT 232.950 87.600 235.050 88.050 ;
        RECT 238.950 87.600 241.050 88.050 ;
        RECT 232.950 86.400 241.050 87.600 ;
        RECT 232.950 85.950 235.050 86.400 ;
        RECT 238.950 85.950 241.050 86.400 ;
        RECT 145.950 81.600 148.050 82.050 ;
        RECT 154.950 81.600 157.050 82.050 ;
        RECT 145.950 80.400 157.050 81.600 ;
        RECT 145.950 79.950 148.050 80.400 ;
        RECT 154.950 79.950 157.050 80.400 ;
        RECT 148.950 78.600 151.050 79.050 ;
        RECT 181.950 78.600 184.050 79.050 ;
        RECT 148.950 77.400 184.050 78.600 ;
        RECT 148.950 76.950 151.050 77.400 ;
        RECT 181.950 76.950 184.050 77.400 ;
        RECT 196.950 78.600 199.050 79.050 ;
        RECT 232.950 78.600 235.050 79.050 ;
        RECT 196.950 77.400 235.050 78.600 ;
        RECT 196.950 76.950 199.050 77.400 ;
        RECT 232.950 76.950 235.050 77.400 ;
        RECT 1.950 75.600 4.050 76.050 ;
        RECT 40.950 75.600 43.050 76.050 ;
        RECT 1.950 74.400 43.050 75.600 ;
        RECT 1.950 73.950 4.050 74.400 ;
        RECT 40.950 73.950 43.050 74.400 ;
        RECT 16.950 72.600 19.050 73.050 ;
        RECT 2.400 71.400 19.050 72.600 ;
        RECT 2.400 54.600 3.600 71.400 ;
        RECT 16.950 70.950 19.050 71.400 ;
        RECT 121.950 72.600 124.050 73.050 ;
        RECT 157.950 72.600 160.050 73.050 ;
        RECT 259.950 72.600 262.050 73.050 ;
        RECT 121.950 71.400 262.050 72.600 ;
        RECT 121.950 70.950 124.050 71.400 ;
        RECT 157.950 70.950 160.050 71.400 ;
        RECT 259.950 70.950 262.050 71.400 ;
        RECT 97.950 69.600 100.050 70.050 ;
        RECT 127.950 69.600 130.050 70.050 ;
        RECT 178.950 69.600 181.050 70.050 ;
        RECT 97.950 68.400 181.050 69.600 ;
        RECT 97.950 67.950 100.050 68.400 ;
        RECT 127.950 67.950 130.050 68.400 ;
        RECT 178.950 67.950 181.050 68.400 ;
        RECT 184.950 69.600 187.050 70.050 ;
        RECT 205.950 69.600 208.050 70.050 ;
        RECT 184.950 68.400 208.050 69.600 ;
        RECT 184.950 67.950 187.050 68.400 ;
        RECT 205.950 67.950 208.050 68.400 ;
        RECT 220.950 69.600 223.050 70.050 ;
        RECT 244.950 69.600 247.050 70.050 ;
        RECT 220.950 68.400 247.050 69.600 ;
        RECT 220.950 67.950 223.050 68.400 ;
        RECT 244.950 67.950 247.050 68.400 ;
        RECT 4.950 66.600 7.050 67.050 ;
        RECT 10.950 66.600 13.050 67.050 ;
        RECT 103.800 66.600 105.900 67.050 ;
        RECT 4.950 65.400 13.050 66.600 ;
        RECT 4.950 64.950 7.050 65.400 ;
        RECT 10.950 64.950 13.050 65.400 ;
        RECT 83.400 65.400 105.900 66.600 ;
        RECT 58.950 63.600 61.050 64.050 ;
        RECT 79.950 63.600 82.050 64.050 ;
        RECT 58.950 62.400 82.050 63.600 ;
        RECT 58.950 61.950 61.050 62.400 ;
        RECT 79.950 61.950 82.050 62.400 ;
        RECT 4.950 60.600 7.050 61.200 ;
        RECT 13.950 60.600 16.050 61.050 ;
        RECT 4.950 59.400 12.600 60.600 ;
        RECT 4.950 59.100 7.050 59.400 ;
        RECT 7.950 54.600 10.050 54.900 ;
        RECT 2.400 53.400 10.050 54.600 ;
        RECT 7.950 52.800 10.050 53.400 ;
        RECT 11.400 52.050 12.600 59.400 ;
        RECT 13.950 59.400 33.600 60.600 ;
        RECT 13.950 58.950 16.050 59.400 ;
        RECT 32.400 55.050 33.600 59.400 ;
        RECT 83.400 58.050 84.600 65.400 ;
        RECT 103.800 64.950 105.900 65.400 ;
        RECT 106.950 66.600 109.050 67.050 ;
        RECT 115.950 66.600 118.050 67.050 ;
        RECT 106.950 65.400 118.050 66.600 ;
        RECT 106.950 64.950 109.050 65.400 ;
        RECT 115.950 64.950 118.050 65.400 ;
        RECT 160.950 66.600 163.050 67.050 ;
        RECT 187.950 66.600 190.050 67.050 ;
        RECT 217.950 66.600 220.050 67.050 ;
        RECT 160.950 65.400 220.050 66.600 ;
        RECT 160.950 64.950 163.050 65.400 ;
        RECT 187.950 64.950 190.050 65.400 ;
        RECT 217.950 64.950 220.050 65.400 ;
        RECT 247.950 66.600 250.050 67.050 ;
        RECT 271.950 66.600 274.050 67.050 ;
        RECT 247.950 65.400 274.050 66.600 ;
        RECT 247.950 64.950 250.050 65.400 ;
        RECT 271.950 64.950 274.050 65.400 ;
        RECT 157.950 61.950 160.050 64.050 ;
        RECT 229.950 63.600 232.050 64.050 ;
        RECT 277.950 63.600 280.050 64.050 ;
        RECT 185.400 62.400 201.600 63.600 ;
        RECT 109.950 59.100 112.050 61.200 ;
        RECT 115.950 60.600 120.000 61.050 ;
        RECT 147.000 60.600 151.050 61.050 ;
        RECT 154.950 60.600 157.050 61.200 ;
        RECT 82.950 55.950 85.050 58.050 ;
        RECT 110.400 57.600 111.600 59.100 ;
        RECT 115.950 58.950 120.600 60.600 ;
        RECT 119.400 57.600 120.600 58.950 ;
        RECT 146.400 58.950 151.050 60.600 ;
        RECT 152.400 59.400 157.050 60.600 ;
        RECT 110.400 57.000 117.600 57.600 ;
        RECT 110.400 56.400 118.050 57.000 ;
        RECT 119.400 56.400 123.600 57.600 ;
        RECT 31.950 52.950 34.050 55.050 ;
        RECT 97.950 54.450 100.050 54.900 ;
        RECT 112.800 54.450 114.900 54.900 ;
        RECT 97.950 53.250 114.900 54.450 ;
        RECT 97.950 52.800 100.050 53.250 ;
        RECT 112.800 52.800 114.900 53.250 ;
        RECT 115.950 52.950 118.050 56.400 ;
        RECT 122.400 54.600 123.600 56.400 ;
        RECT 124.950 54.600 127.050 54.900 ;
        RECT 122.400 53.400 127.050 54.600 ;
        RECT 124.950 52.800 127.050 53.400 ;
        RECT 130.950 54.600 133.050 55.050 ;
        RECT 146.400 54.600 147.600 58.950 ;
        RECT 152.400 57.600 153.600 59.400 ;
        RECT 154.950 59.100 157.050 59.400 ;
        RECT 158.400 57.600 159.600 61.950 ;
        RECT 163.950 58.950 166.050 61.050 ;
        RECT 178.950 59.100 181.050 61.200 ;
        RECT 149.400 57.000 153.600 57.600 ;
        RECT 130.950 53.400 147.600 54.600 ;
        RECT 148.950 56.400 153.600 57.000 ;
        RECT 155.400 56.400 159.600 57.600 ;
        RECT 130.950 52.950 133.050 53.400 ;
        RECT 148.950 52.950 151.050 56.400 ;
        RECT 155.400 54.600 156.600 56.400 ;
        RECT 164.400 55.050 165.600 58.950 ;
        RECT 152.400 53.400 156.600 54.600 ;
        RECT 10.950 49.950 13.050 52.050 ;
        RECT 127.950 51.600 130.050 52.050 ;
        RECT 152.400 51.600 153.600 53.400 ;
        RECT 163.800 52.950 165.900 55.050 ;
        RECT 166.950 54.600 169.050 54.900 ;
        RECT 179.400 54.600 180.600 59.100 ;
        RECT 166.950 53.400 180.600 54.600 ;
        RECT 166.950 52.800 169.050 53.400 ;
        RECT 185.400 52.050 186.600 62.400 ;
        RECT 200.400 61.200 201.600 62.400 ;
        RECT 224.400 62.400 232.050 63.600 ;
        RECT 187.950 58.950 190.050 61.050 ;
        RECT 193.950 59.100 196.050 61.200 ;
        RECT 199.950 59.100 202.050 61.200 ;
        RECT 127.950 50.400 153.600 51.600 ;
        RECT 127.950 49.950 130.050 50.400 ;
        RECT 184.950 49.950 187.050 52.050 ;
        RECT 188.400 51.600 189.600 58.950 ;
        RECT 194.400 55.050 195.600 59.100 ;
        RECT 205.950 58.950 208.050 61.050 ;
        RECT 214.950 59.100 217.050 61.200 ;
        RECT 206.400 55.050 207.600 58.950 ;
        RECT 190.950 53.400 195.600 55.050 ;
        RECT 190.950 52.950 195.000 53.400 ;
        RECT 205.950 52.950 208.050 55.050 ;
        RECT 196.950 51.600 199.050 52.050 ;
        RECT 188.400 50.400 199.050 51.600 ;
        RECT 196.950 49.950 199.050 50.400 ;
        RECT 202.950 51.600 205.050 52.050 ;
        RECT 215.400 51.600 216.600 59.100 ;
        RECT 220.950 58.950 223.050 61.050 ;
        RECT 221.400 55.050 222.600 58.950 ;
        RECT 224.400 55.050 225.600 62.400 ;
        RECT 229.950 61.950 232.050 62.400 ;
        RECT 257.400 62.400 280.050 63.600 ;
        RECT 232.950 60.600 235.050 61.050 ;
        RECT 232.950 59.400 240.600 60.600 ;
        RECT 232.950 58.950 235.050 59.400 ;
        RECT 220.800 52.950 222.900 55.050 ;
        RECT 223.950 52.950 226.050 55.050 ;
        RECT 239.400 54.900 240.600 59.400 ;
        RECT 257.400 57.600 258.600 62.400 ;
        RECT 277.950 61.950 280.050 62.400 ;
        RECT 259.950 59.100 262.050 61.200 ;
        RECT 265.950 59.100 268.050 61.200 ;
        RECT 245.400 56.400 258.600 57.600 ;
        RECT 245.400 54.900 246.600 56.400 ;
        RECT 238.950 52.800 241.050 54.900 ;
        RECT 244.950 52.800 247.050 54.900 ;
        RECT 202.950 50.400 216.600 51.600 ;
        RECT 247.950 51.600 250.050 52.050 ;
        RECT 260.400 51.600 261.600 59.100 ;
        RECT 266.400 55.050 267.600 59.100 ;
        RECT 266.400 53.400 271.050 55.050 ;
        RECT 267.000 52.950 271.050 53.400 ;
        RECT 280.950 54.600 283.050 54.900 ;
        RECT 307.950 54.600 310.050 58.050 ;
        RECT 280.950 54.000 310.050 54.600 ;
        RECT 280.950 53.400 309.600 54.000 ;
        RECT 280.950 52.800 283.050 53.400 ;
        RECT 247.950 50.400 261.600 51.600 ;
        RECT 202.950 49.950 205.050 50.400 ;
        RECT 247.950 49.950 250.050 50.400 ;
        RECT 133.950 48.600 136.050 49.050 ;
        RECT 148.950 48.600 151.050 49.050 ;
        RECT 160.950 48.600 163.050 49.050 ;
        RECT 133.950 47.400 163.050 48.600 ;
        RECT 133.950 46.950 136.050 47.400 ;
        RECT 148.950 46.950 151.050 47.400 ;
        RECT 160.950 46.950 163.050 47.400 ;
        RECT 220.950 48.600 223.050 49.050 ;
        RECT 229.950 48.600 232.050 49.050 ;
        RECT 220.950 47.400 232.050 48.600 ;
        RECT 220.950 46.950 223.050 47.400 ;
        RECT 229.950 46.950 232.050 47.400 ;
        RECT 178.950 45.600 181.050 46.050 ;
        RECT 190.950 45.600 193.050 46.050 ;
        RECT 235.950 45.600 238.050 46.050 ;
        RECT 178.950 44.400 238.050 45.600 ;
        RECT 178.950 43.950 181.050 44.400 ;
        RECT 190.950 43.950 193.050 44.400 ;
        RECT 235.950 43.950 238.050 44.400 ;
        RECT 265.950 45.600 268.050 46.050 ;
        RECT 274.950 45.600 277.050 46.050 ;
        RECT 265.950 44.400 277.050 45.600 ;
        RECT 265.950 43.950 268.050 44.400 ;
        RECT 274.950 43.950 277.050 44.400 ;
        RECT 142.950 42.600 145.050 43.050 ;
        RECT 151.950 42.600 154.050 43.050 ;
        RECT 142.950 41.400 154.050 42.600 ;
        RECT 142.950 40.950 145.050 41.400 ;
        RECT 151.950 40.950 154.050 41.400 ;
        RECT 181.950 42.600 184.050 43.050 ;
        RECT 211.950 42.600 214.050 43.050 ;
        RECT 181.950 41.400 214.050 42.600 ;
        RECT 181.950 40.950 184.050 41.400 ;
        RECT 211.950 40.950 214.050 41.400 ;
        RECT 79.950 39.600 82.050 40.050 ;
        RECT 106.950 39.600 109.050 40.050 ;
        RECT 79.950 38.400 109.050 39.600 ;
        RECT 79.950 37.950 82.050 38.400 ;
        RECT 106.950 37.950 109.050 38.400 ;
        RECT 130.950 39.600 133.050 40.050 ;
        RECT 157.950 39.600 160.050 40.050 ;
        RECT 130.950 38.400 160.050 39.600 ;
        RECT 130.950 37.950 133.050 38.400 ;
        RECT 157.950 37.950 160.050 38.400 ;
        RECT 184.950 39.600 187.050 40.050 ;
        RECT 199.950 39.600 202.050 40.050 ;
        RECT 184.950 38.400 202.050 39.600 ;
        RECT 184.950 37.950 187.050 38.400 ;
        RECT 199.950 37.950 202.050 38.400 ;
        RECT 109.950 36.600 112.050 37.050 ;
        RECT 127.950 36.600 130.050 37.050 ;
        RECT 109.950 35.400 130.050 36.600 ;
        RECT 109.950 34.950 112.050 35.400 ;
        RECT 127.950 34.950 130.050 35.400 ;
        RECT 160.950 36.600 163.050 37.050 ;
        RECT 178.950 36.600 181.050 37.050 ;
        RECT 160.950 35.400 181.050 36.600 ;
        RECT 160.950 34.950 163.050 35.400 ;
        RECT 178.950 34.950 181.050 35.400 ;
        RECT 205.950 36.600 208.050 37.050 ;
        RECT 214.950 36.600 217.050 37.050 ;
        RECT 232.950 36.600 235.050 37.050 ;
        RECT 253.800 36.600 255.900 37.050 ;
        RECT 268.950 36.600 271.050 37.050 ;
        RECT 346.950 36.600 349.050 37.050 ;
        RECT 205.950 35.400 255.900 36.600 ;
        RECT 205.950 34.950 208.050 35.400 ;
        RECT 214.950 34.950 217.050 35.400 ;
        RECT 232.950 34.950 235.050 35.400 ;
        RECT 253.800 34.950 255.900 35.400 ;
        RECT 257.400 35.400 349.050 36.600 ;
        RECT 257.400 34.050 258.600 35.400 ;
        RECT 268.950 34.950 271.050 35.400 ;
        RECT 346.950 34.950 349.050 35.400 ;
        RECT 115.950 33.600 118.050 34.050 ;
        RECT 130.950 33.600 133.050 34.050 ;
        RECT 115.950 32.400 133.050 33.600 ;
        RECT 115.950 31.950 118.050 32.400 ;
        RECT 130.950 31.950 133.050 32.400 ;
        RECT 172.950 33.600 175.050 34.050 ;
        RECT 223.950 33.600 226.050 34.050 ;
        RECT 172.950 32.400 226.050 33.600 ;
        RECT 172.950 31.950 175.050 32.400 ;
        RECT 223.950 31.950 226.050 32.400 ;
        RECT 241.950 33.600 244.050 34.050 ;
        RECT 256.950 33.600 259.050 34.050 ;
        RECT 334.950 33.600 337.050 34.050 ;
        RECT 241.950 32.400 259.050 33.600 ;
        RECT 241.950 31.950 244.050 32.400 ;
        RECT 256.950 31.950 259.050 32.400 ;
        RECT 323.400 32.400 337.050 33.600 ;
        RECT 323.400 31.050 324.600 32.400 ;
        RECT 334.950 31.950 337.050 32.400 ;
        RECT 142.950 30.600 145.050 31.050 ;
        RECT 163.950 30.600 166.050 31.050 ;
        RECT 238.950 30.600 241.050 31.050 ;
        RECT 142.950 29.400 166.050 30.600 ;
        RECT 142.950 28.950 145.050 29.400 ;
        RECT 163.950 28.950 166.050 29.400 ;
        RECT 224.400 29.400 241.050 30.600 ;
        RECT 10.950 27.600 13.050 28.200 ;
        RECT 76.950 27.600 79.050 28.050 ;
        RECT 10.950 26.400 79.050 27.600 ;
        RECT 10.950 26.100 13.050 26.400 ;
        RECT 76.950 25.950 79.050 26.400 ;
        RECT 94.950 27.750 97.050 28.200 ;
        RECT 109.950 27.750 112.050 28.200 ;
        RECT 94.950 26.550 112.050 27.750 ;
        RECT 94.950 26.100 97.050 26.550 ;
        RECT 109.950 26.100 112.050 26.550 ;
        RECT 115.950 26.100 118.050 28.200 ;
        RECT 133.950 27.600 136.050 28.200 ;
        RECT 142.950 27.600 145.050 28.200 ;
        RECT 133.950 26.400 145.050 27.600 ;
        RECT 133.950 26.100 136.050 26.400 ;
        RECT 142.950 26.100 145.050 26.400 ;
        RECT 154.950 26.100 157.050 28.200 ;
        RECT 181.950 27.600 184.050 28.200 ;
        RECT 176.400 26.400 184.050 27.600 ;
        RECT 25.950 24.450 28.050 25.050 ;
        RECT 40.950 24.450 43.050 24.900 ;
        RECT 25.950 23.250 43.050 24.450 ;
        RECT 25.950 22.950 28.050 23.250 ;
        RECT 40.950 22.800 43.050 23.250 ;
        RECT 116.400 21.600 117.600 26.100 ;
        RECT 121.950 21.600 124.050 21.900 ;
        RECT 116.400 20.400 124.050 21.600 ;
        RECT 121.950 19.800 124.050 20.400 ;
        RECT 145.950 21.600 148.050 21.900 ;
        RECT 155.400 21.600 156.600 26.100 ;
        RECT 176.400 21.900 177.600 26.400 ;
        RECT 181.950 26.100 184.050 26.400 ;
        RECT 193.950 26.100 196.050 28.200 ;
        RECT 178.950 24.600 181.050 25.050 ;
        RECT 194.400 24.600 195.600 26.100 ;
        RECT 217.950 25.950 220.050 28.050 ;
        RECT 178.950 23.400 195.600 24.600 ;
        RECT 178.950 22.950 181.050 23.400 ;
        RECT 218.400 22.050 219.600 25.950 ;
        RECT 145.950 20.400 156.600 21.600 ;
        RECT 157.950 21.600 160.050 21.900 ;
        RECT 166.950 21.600 169.050 21.900 ;
        RECT 157.950 20.400 169.050 21.600 ;
        RECT 145.950 19.800 148.050 20.400 ;
        RECT 157.950 19.800 160.050 20.400 ;
        RECT 166.950 19.800 169.050 20.400 ;
        RECT 175.950 19.800 178.050 21.900 ;
        RECT 202.950 21.600 205.050 21.900 ;
        RECT 211.950 21.600 214.050 21.900 ;
        RECT 202.950 20.400 214.050 21.600 ;
        RECT 202.950 19.800 205.050 20.400 ;
        RECT 211.950 19.800 214.050 20.400 ;
        RECT 217.950 19.950 220.050 22.050 ;
        RECT 224.400 19.050 225.600 29.400 ;
        RECT 238.950 28.950 241.050 29.400 ;
        RECT 253.950 30.600 256.050 31.050 ;
        RECT 322.950 30.600 325.050 31.050 ;
        RECT 253.950 29.400 325.050 30.600 ;
        RECT 253.950 28.950 256.050 29.400 ;
        RECT 322.950 28.950 325.050 29.400 ;
        RECT 232.950 25.950 235.050 28.050 ;
        RECT 247.950 25.950 250.050 28.050 ;
        RECT 264.000 27.600 268.050 28.050 ;
        RECT 263.400 25.950 268.050 27.600 ;
        RECT 233.400 21.600 234.600 25.950 ;
        RECT 238.950 21.600 241.050 21.900 ;
        RECT 233.400 20.400 241.050 21.600 ;
        RECT 238.950 19.800 241.050 20.400 ;
        RECT 244.950 21.600 247.050 21.900 ;
        RECT 248.400 21.600 249.600 25.950 ;
        RECT 244.950 20.400 249.600 21.600 ;
        RECT 253.950 21.600 256.050 21.900 ;
        RECT 263.400 21.600 264.600 25.950 ;
        RECT 253.950 20.400 264.600 21.600 ;
        RECT 244.950 19.800 247.050 20.400 ;
        RECT 253.950 19.800 256.050 20.400 ;
        RECT 82.950 18.600 85.050 19.050 ;
        RECT 103.950 18.600 106.050 19.050 ;
        RECT 82.950 17.400 106.050 18.600 ;
        RECT 82.950 16.950 85.050 17.400 ;
        RECT 103.950 16.950 106.050 17.400 ;
        RECT 220.950 17.400 225.600 19.050 ;
        RECT 220.950 16.950 225.000 17.400 ;
        RECT 121.950 15.600 124.050 16.050 ;
        RECT 178.950 15.600 181.050 16.050 ;
        RECT 121.950 14.400 181.050 15.600 ;
        RECT 121.950 13.950 124.050 14.400 ;
        RECT 178.950 13.950 181.050 14.400 ;
        RECT 112.950 12.600 115.050 13.050 ;
        RECT 136.950 12.600 139.050 13.050 ;
        RECT 112.950 11.400 139.050 12.600 ;
        RECT 112.950 10.950 115.050 11.400 ;
        RECT 136.950 10.950 139.050 11.400 ;
        RECT 217.950 12.600 220.050 13.050 ;
        RECT 286.950 12.600 289.050 13.050 ;
        RECT 217.950 11.400 289.050 12.600 ;
        RECT 217.950 10.950 220.050 11.400 ;
        RECT 286.950 10.950 289.050 11.400 ;
        RECT 196.950 3.600 199.050 4.050 ;
        RECT 253.950 3.600 256.050 4.050 ;
        RECT 196.950 2.400 256.050 3.600 ;
        RECT 196.950 1.950 199.050 2.400 ;
        RECT 253.950 1.950 256.050 2.400 ;
  END
END counter16
END LIBRARY

