magic
tech scmos
magscale 1 30
timestamp 1749790639
<< checkpaint >>
rect 9150 9150 180850 180850
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI
timestamp 1725930584
transform 0 -1 171100 -1 0 75646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_1
timestamp 1725930584
transform 0 -1 171098 -1 0 62146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_2
timestamp 1725930584
transform 0 -1 171100 -1 0 102646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_3
timestamp 1725930584
transform 0 -1 171100 -1 0 89146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_4
timestamp 1725930584
transform 0 -1 171102 -1 0 129646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_5
timestamp 1725930584
transform 0 -1 171100 -1 0 116146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_6
timestamp 1725930584
transform 1 0 73845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_7
timestamp 1725930584
transform 1 0 60345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_8
timestamp 1725930584
transform 1 0 100845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_9
timestamp 1725930584
transform 1 0 87345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_10
timestamp 1725930584
transform 1 0 127845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_11
timestamp 1725930584
transform 1 0 114345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_12
timestamp 1725930584
transform 0 1 18899 -1 0 75655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_13
timestamp 1725930584
transform 0 1 18899 -1 0 62155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_14
timestamp 1725930584
transform 0 1 18900 -1 0 102655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_15
timestamp 1725930584
transform 0 1 18900 -1 0 89155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_16
timestamp 1725930584
transform 1 0 73845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_17
timestamp 1725930584
transform 0 1 18897 -1 0 116155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_18
timestamp 1725930584
transform 0 1 18900 -1 0 129655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_19
timestamp 1725930584
transform 1 0 60345 0 -1 171101
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_20
timestamp 1725930584
transform 1 0 100845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_21
timestamp 1725930584
transform 1 0 87344 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_22
timestamp 1725930584
transform 1 0 127845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_23
timestamp 1725930584
transform 1 0 114345 0 -1 171100
box -60 0 1860 25060
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 43621 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1569139307
transform 1 0 141360 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1569139307
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1569139307
transform 1 0 43638 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1569139307
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1569139307
transform 0 1 18900 -1 0 146379
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1569139307
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1569139307
transform 0 -1 171100 -1 0 146346
box -35 0 5035 25060
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1569139307
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1569139307
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1569139307
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use PIC  clk ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use PIC  down
timestamp 1569139307
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use PIC  enable
timestamp 1569139307
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use PIC  INV_IN
timestamp 1569139307
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use PIC  NAND_IN
timestamp 1569139307
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
use PIC  reset
timestamp 1569139307
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use PIC  up
timestamp 1569139307
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use POB8  hsync ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use POB8  INV_OUT1
timestamp 1569139307
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use POB8  INV_OUT8
timestamp 1569139307
transform 0 -1 171100 1 0 102500
box -100 -9150 12100 25300
use POB8  NAND_OUT1
timestamp 1569139307
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use POB8  NAND_OUT8
timestamp 1569139307
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use POB8  p_tick
timestamp 1569139307
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use POB8  rgb
timestamp 1569139307
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use POB8  vsync
timestamp 1569139307
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use PANA  INV_INA ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 0 1 18900 -1 0 87500
box -100 -9150 12095 25300
use PANA  INV_OUT1A
timestamp 1569139307
transform 0 1 18900 -1 0 74000
box -100 -9150 12095 25300
use PANA  INV_OUT8A
timestamp 1569139307
transform 0 1 18900 -1 0 60500
box -100 -9150 12095 25300
use PANA  NAND_OUT1A
timestamp 1569139307
transform 0 1 18900 -1 0 128000
box -100 -9150 12095 25300
use PANA  NAND_OUT8A
timestamp 1569139307
transform 0 1 18900 -1 0 114500
box -100 -9150 12095 25300
use PANA  PANA_0
timestamp 1569139307
transform 0 1 18900 -1 0 141500
box -100 -9150 12095 25300
use PVSS  GND ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 62000 0 1 18900
box 0 -9150 12000 25300
use PVSS  PVSS_0
timestamp 1569139307
transform 1 0 129500 0 1 18900
box 0 -9150 12000 25300
use PVSS  PVSS_1
timestamp 1569139307
transform 1 0 129500 0 -1 171100
box 0 -9150 12000 25300
use PVSS  PVSS_2
timestamp 1569139307
transform 0 1 18900 -1 0 101000
box 0 -9150 12000 25300
use PVDD  PVDD_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 48500 0 1 18900
box 0 -9150 12000 25300
use PVDD  PVDD_1
timestamp 1569139307
transform 0 -1 171100 1 0 89000
box 0 -9150 12000 25300
use PVDD  VCC
timestamp 1569139307
transform 1 0 48500 0 -1 171100
box 0 -9150 12000 25300
<< end >>