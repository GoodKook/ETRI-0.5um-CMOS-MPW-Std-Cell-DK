magic
tech scmos
magscale 1 2
timestamp 1727166839
<< metal1 >>
rect -63 5738 -3 5998
rect 5950 5982 6043 5998
rect 4727 5917 4813 5923
rect 3967 5903 3980 5907
rect 3967 5893 3983 5903
rect 3627 5877 3694 5883
rect 3977 5867 3983 5893
rect 1177 5857 1213 5863
rect 2827 5857 2873 5863
rect 3967 5857 3983 5867
rect 3967 5853 3980 5857
rect 2967 5837 3113 5843
rect 4087 5837 4153 5843
rect 4727 5837 4793 5843
rect 5067 5837 5173 5843
rect 3007 5817 3033 5823
rect 4873 5823 4887 5833
rect 4873 5820 4933 5823
rect 4877 5817 4933 5820
rect -63 5722 30 5738
rect -63 5218 -3 5722
rect 1707 5617 1753 5623
rect 2427 5617 2493 5623
rect 2507 5617 2533 5623
rect 4447 5617 4493 5623
rect 4967 5617 5033 5623
rect 5787 5617 5853 5623
rect 5867 5617 5913 5623
rect 5027 5603 5040 5607
rect 5027 5593 5043 5603
rect 5167 5603 5180 5607
rect 5167 5593 5183 5603
rect 3940 5583 3953 5587
rect 3787 5577 3834 5583
rect 3937 5577 3953 5583
rect 3940 5573 3953 5577
rect 5037 5567 5043 5593
rect 2957 5560 3013 5563
rect 2953 5557 3013 5560
rect 2953 5547 2967 5557
rect 5027 5557 5043 5567
rect 5027 5553 5040 5557
rect 2447 5537 2473 5543
rect 3413 5543 3427 5553
rect 3413 5540 3473 5543
rect 3417 5537 3473 5540
rect 5177 5546 5183 5593
rect 5983 5478 6043 5982
rect 5950 5462 6043 5478
rect 147 5377 183 5383
rect 177 5347 183 5377
rect 4287 5377 4323 5383
rect 4317 5347 4323 5377
rect 177 5337 193 5347
rect 180 5333 193 5337
rect 1527 5337 1573 5343
rect 4317 5337 4333 5347
rect 4320 5333 4333 5337
rect 287 5317 353 5323
rect 1467 5317 1533 5323
rect 1907 5317 2053 5323
rect 2547 5317 2633 5323
rect 4227 5317 4293 5323
rect 4387 5317 4493 5323
rect 5407 5317 5453 5323
rect 5827 5317 5873 5323
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 3307 5117 3373 5123
rect 4747 5117 4773 5123
rect 1907 5097 2013 5103
rect 2227 5097 2273 5103
rect 2787 5097 2893 5103
rect 3347 5097 3413 5103
rect 5687 5097 5773 5103
rect 300 5083 313 5087
rect 297 5073 313 5083
rect 2700 5083 2713 5087
rect 2697 5073 2713 5083
rect 3800 5083 3813 5087
rect 3797 5073 3813 5083
rect 4047 5083 4060 5087
rect 4047 5073 4063 5083
rect 4467 5083 4480 5087
rect 4467 5073 4483 5083
rect 5067 5083 5080 5087
rect 5067 5073 5083 5083
rect 5547 5077 5613 5083
rect 5700 5083 5713 5087
rect 5697 5073 5713 5083
rect 297 5047 303 5073
rect 2697 5047 2703 5073
rect 297 5037 313 5047
rect 300 5033 313 5037
rect 2697 5037 2713 5047
rect 2700 5033 2713 5037
rect 3797 5043 3803 5073
rect 4057 5047 4063 5073
rect 3747 5037 3803 5043
rect 4047 5037 4063 5047
rect 4477 5047 4483 5073
rect 4477 5037 4493 5047
rect 4047 5033 4060 5037
rect 4480 5033 4493 5037
rect 5077 5043 5083 5073
rect 5697 5047 5703 5073
rect 5077 5037 5133 5043
rect 5687 5037 5703 5047
rect 5687 5033 5700 5037
rect 4807 5017 4873 5023
rect 5983 4958 6043 5462
rect 5950 4942 6043 4958
rect 3807 4863 3820 4867
rect 3807 4853 3823 4863
rect 5667 4863 5680 4867
rect 5700 4863 5713 4867
rect 5667 4853 5683 4863
rect 3817 4827 3823 4853
rect 287 4817 333 4823
rect 3807 4817 3823 4827
rect 3807 4813 3820 4817
rect 2067 4797 2133 4803
rect 5327 4797 5433 4803
rect 5677 4803 5683 4853
rect 5697 4853 5713 4863
rect 5697 4827 5703 4853
rect 5697 4817 5713 4827
rect 5700 4813 5713 4817
rect 5827 4817 5933 4823
rect 5677 4797 5733 4803
rect 4287 4777 4353 4783
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 3607 4657 3633 4663
rect 2787 4637 2813 4643
rect 167 4577 203 4583
rect 197 4527 203 4577
rect 1327 4577 1383 4583
rect 327 4557 373 4563
rect 1377 4563 1383 4577
rect 4347 4577 4453 4583
rect 5667 4577 5713 4583
rect 5727 4577 5773 4583
rect 2820 4563 2833 4567
rect 1377 4557 1403 4563
rect 1397 4527 1403 4557
rect 197 4517 213 4527
rect 200 4513 213 4517
rect 1387 4517 1403 4527
rect 2817 4553 2833 4563
rect 3287 4563 3300 4567
rect 3780 4563 3793 4567
rect 3287 4553 3303 4563
rect 2817 4527 2823 4553
rect 3297 4543 3303 4553
rect 3777 4553 3793 4563
rect 3907 4563 3920 4567
rect 4600 4563 4613 4567
rect 3907 4553 3923 4563
rect 3297 4537 3333 4543
rect 3777 4527 3783 4553
rect 3917 4527 3923 4553
rect 4597 4553 4613 4563
rect 5827 4563 5840 4567
rect 5827 4553 5843 4563
rect 2817 4517 2833 4527
rect 1387 4513 1400 4517
rect 2820 4513 2833 4517
rect 3127 4517 3173 4523
rect 3777 4517 3793 4527
rect 3780 4513 3793 4517
rect 3907 4517 3923 4527
rect 3907 4513 3920 4517
rect 4597 4523 4603 4553
rect 5837 4527 5843 4553
rect 4567 4517 4603 4523
rect 5347 4517 5373 4523
rect 5827 4523 5843 4527
rect 5827 4517 5873 4523
rect 5827 4513 5840 4517
rect 2807 4477 2833 4483
rect 807 4457 853 4463
rect 2327 4457 2353 4463
rect 5983 4438 6043 4942
rect 5950 4422 6043 4438
rect 5647 4397 5673 4403
rect 67 4377 93 4383
rect 447 4377 513 4383
rect 2067 4377 2113 4383
rect 567 4357 593 4363
rect 1387 4357 1433 4363
rect 3647 4357 3713 4363
rect 4547 4357 4613 4363
rect 5007 4357 5073 4363
rect 180 4343 193 4347
rect 177 4333 193 4343
rect 2787 4343 2800 4347
rect 3820 4343 3833 4347
rect 2787 4333 2803 4343
rect 177 4307 183 4333
rect 2797 4307 2803 4333
rect 177 4297 193 4307
rect 180 4293 193 4297
rect 2787 4297 2803 4307
rect 3817 4333 3833 4343
rect 4387 4343 4400 4347
rect 4693 4343 4707 4353
rect 4387 4333 4403 4343
rect 4693 4340 4723 4343
rect 4697 4337 4723 4340
rect 3817 4307 3823 4333
rect 4397 4307 4403 4333
rect 4513 4307 4527 4313
rect 3817 4297 3833 4307
rect 2787 4293 2800 4297
rect 3820 4293 3833 4297
rect 4387 4297 4403 4307
rect 4387 4293 4400 4297
rect 4507 4300 4527 4307
rect 4717 4307 4723 4337
rect 4867 4343 4880 4347
rect 5520 4343 5533 4347
rect 4867 4333 4883 4343
rect 4877 4307 4883 4333
rect 4507 4297 4523 4300
rect 4717 4297 4733 4307
rect 4507 4293 4520 4297
rect 4720 4293 4733 4297
rect 4867 4297 4883 4307
rect 5517 4333 5533 4343
rect 5827 4343 5840 4347
rect 5827 4333 5843 4343
rect 5517 4307 5523 4333
rect 5837 4307 5843 4333
rect 5517 4297 5533 4307
rect 4867 4293 4880 4297
rect 5520 4293 5533 4297
rect 5827 4297 5843 4307
rect 5827 4293 5840 4297
rect 2907 4277 2973 4283
rect 4227 4277 4293 4283
rect 4487 4277 4513 4283
rect 4987 4277 5093 4283
rect 5767 4277 5873 4283
rect 5047 4257 5113 4263
rect 2767 4237 2853 4243
rect 27 4197 53 4203
rect 4887 4197 4913 4203
rect -63 4162 30 4178
rect -63 3658 -3 4162
rect 587 4117 623 4123
rect 617 4067 623 4117
rect 5087 4117 5113 4123
rect 167 4057 243 4063
rect 617 4057 633 4067
rect 237 4043 243 4057
rect 620 4053 633 4057
rect 2447 4057 2493 4063
rect 2507 4057 2553 4063
rect 3897 4057 3973 4063
rect 237 4037 263 4043
rect 1857 4037 1913 4043
rect 387 4017 454 4023
rect 3487 3997 3553 4003
rect 3897 3987 3903 4057
rect 4087 4057 4113 4063
rect 4807 4057 4833 4063
rect 4947 4057 5013 4063
rect 5313 4063 5327 4073
rect 5287 4060 5327 4063
rect 5287 4057 5323 4060
rect 5807 4057 5913 4063
rect 4057 4037 4093 4043
rect 4057 4007 4063 4037
rect 4193 4043 4207 4053
rect 4193 4040 4223 4043
rect 4197 4037 4223 4040
rect 4217 4007 4223 4037
rect 4047 3997 4063 4007
rect 4047 3993 4060 3997
rect 4207 3997 4223 4007
rect 4207 3993 4220 3997
rect 4237 3987 4243 4053
rect 4357 4007 4363 4053
rect 4660 4043 4673 4047
rect 4347 3997 4363 4007
rect 4657 4033 4673 4043
rect 4907 4043 4920 4047
rect 4940 4043 4953 4047
rect 4907 4033 4923 4043
rect 4657 4007 4663 4033
rect 4657 3997 4673 4007
rect 4347 3993 4360 3997
rect 4660 3993 4673 3997
rect 4917 4003 4923 4033
rect 4897 4000 4923 4003
rect 4893 3997 4923 4000
rect 4937 4033 4953 4043
rect 5067 4037 5103 4043
rect 4937 4007 4943 4033
rect 5097 4007 5103 4037
rect 5247 4037 5273 4043
rect 5560 4043 5573 4047
rect 5557 4033 5573 4043
rect 5557 4007 5563 4033
rect 4937 3997 4953 4007
rect 4893 3987 4907 3997
rect 4940 3993 4953 3997
rect 5097 3997 5113 4007
rect 5100 3993 5113 3997
rect 5547 3997 5563 4007
rect 5547 3993 5560 3997
rect 2167 3977 2193 3983
rect 5707 3977 5733 3983
rect 5247 3957 5313 3963
rect 5983 3918 6043 4422
rect 5950 3902 6043 3918
rect 3327 3837 3393 3843
rect 4913 3843 4927 3853
rect 4847 3840 4927 3843
rect 4847 3837 4923 3840
rect 5367 3843 5380 3847
rect 5367 3833 5383 3843
rect 167 3823 180 3827
rect 4440 3823 4453 3827
rect 167 3813 183 3823
rect 177 3783 183 3813
rect 4437 3813 4453 3823
rect 4577 3817 4613 3823
rect 4437 3787 4443 3813
rect 4577 3787 4583 3817
rect 5020 3823 5033 3827
rect 5017 3813 5033 3823
rect 5200 3823 5213 3827
rect 5197 3813 5213 3823
rect 5347 3823 5360 3827
rect 5347 3813 5363 3823
rect 4717 3787 4723 3813
rect 5017 3787 5023 3813
rect 177 3777 213 3783
rect 3887 3777 3913 3783
rect 4437 3777 4453 3787
rect 4440 3773 4453 3777
rect 4567 3777 4583 3787
rect 4567 3773 4580 3777
rect 5007 3777 5023 3787
rect 5197 3787 5203 3813
rect 5357 3787 5363 3813
rect 5377 3807 5383 3833
rect 5377 3806 5400 3807
rect 5377 3797 5393 3806
rect 5380 3793 5393 3797
rect 5197 3777 5213 3787
rect 5007 3773 5020 3777
rect 5200 3773 5213 3777
rect 5347 3777 5363 3787
rect 5537 3783 5543 3873
rect 5537 3777 5563 3783
rect 5347 3773 5360 3777
rect 5557 3767 5563 3777
rect 327 3757 393 3763
rect 1047 3757 1113 3763
rect 1227 3757 1253 3763
rect 5147 3757 5253 3763
rect 5557 3757 5573 3767
rect 5560 3753 5573 3757
rect 307 3677 353 3683
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 3047 3557 3093 3563
rect 4027 3557 4073 3563
rect 887 3537 913 3543
rect 2027 3537 2073 3543
rect 3307 3537 3393 3543
rect 4587 3537 4613 3543
rect 3327 3523 3340 3527
rect 3327 3513 3343 3523
rect 3867 3517 3933 3523
rect 367 3503 380 3507
rect 367 3497 394 3503
rect 367 3493 380 3497
rect 3337 3487 3343 3513
rect 3327 3477 3343 3487
rect 3917 3487 3923 3517
rect 5120 3523 5133 3527
rect 5117 3513 5133 3523
rect 5227 3523 5240 3527
rect 5227 3513 5243 3523
rect 5117 3503 5123 3513
rect 5097 3497 5123 3503
rect 3917 3477 3933 3487
rect 3327 3473 3340 3477
rect 3920 3473 3933 3477
rect 5097 3483 5103 3497
rect 5237 3487 5243 3513
rect 5067 3477 5103 3483
rect 5227 3477 5243 3487
rect 5227 3473 5240 3477
rect 1887 3457 1933 3463
rect 2507 3457 2553 3463
rect 5393 3463 5407 3473
rect 5347 3460 5407 3463
rect 5347 3457 5403 3460
rect 5627 3457 5693 3463
rect 3173 3423 3187 3433
rect 3173 3420 3213 3423
rect 3177 3417 3213 3420
rect 5983 3398 6043 3902
rect 5950 3382 6043 3398
rect 4647 3360 4703 3363
rect 4647 3357 4707 3360
rect 4693 3347 4707 3357
rect 2227 3337 2253 3343
rect 1333 3303 1347 3313
rect 1413 3303 1427 3313
rect 1333 3300 1427 3303
rect 4527 3317 4553 3323
rect 4847 3317 4913 3323
rect 5287 3317 5373 3323
rect 3873 3303 3887 3313
rect 3873 3300 3923 3303
rect 1337 3297 1423 3300
rect 3877 3297 3923 3300
rect 3917 3267 3923 3297
rect 4047 3303 4060 3307
rect 5780 3303 5793 3307
rect 4047 3293 4063 3303
rect 4057 3267 4063 3293
rect 5777 3293 5793 3303
rect 5907 3303 5920 3307
rect 5907 3293 5923 3303
rect 5777 3267 5783 3293
rect 5917 3267 5923 3293
rect 1207 3257 1253 3263
rect 3917 3257 3933 3267
rect 3920 3253 3933 3257
rect 4057 3257 4073 3267
rect 4060 3253 4073 3257
rect 5777 3257 5793 3267
rect 5780 3253 5793 3257
rect 5907 3257 5923 3267
rect 5907 3253 5920 3257
rect 3927 3237 3953 3243
rect 4167 3237 4253 3243
rect 4647 3237 4713 3243
rect 5127 3237 5213 3243
rect 5467 3237 5513 3243
rect 2747 3217 2833 3223
rect 3907 3217 3933 3223
rect 5127 3217 5153 3223
rect -63 3122 30 3138
rect -63 2618 -3 3122
rect 5687 3057 5713 3063
rect 3987 3017 4053 3023
rect 4907 3017 5013 3023
rect 5240 3023 5253 3027
rect 5237 3013 5253 3023
rect 5837 3017 5893 3023
rect 717 2997 753 3003
rect 807 2983 820 2987
rect 807 2977 834 2983
rect 807 2973 820 2977
rect 5237 2963 5243 3013
rect 5567 2997 5613 3003
rect 5707 3003 5720 3007
rect 5707 2993 5723 3003
rect 5267 2983 5280 2987
rect 5267 2977 5294 2983
rect 5267 2973 5280 2977
rect 5217 2957 5243 2963
rect 5397 2957 5433 2963
rect 5217 2947 5223 2957
rect 5717 2963 5723 2993
rect 5837 2963 5843 3017
rect 5717 2957 5743 2963
rect 5837 2957 5863 2963
rect 5207 2937 5223 2947
rect 5737 2947 5743 2957
rect 5737 2937 5753 2947
rect 5207 2933 5220 2937
rect 5740 2933 5753 2937
rect 5857 2943 5863 2957
rect 5857 2937 5913 2943
rect 5983 2878 6043 3382
rect 5950 2862 6043 2878
rect 727 2797 793 2803
rect 280 2783 293 2787
rect 277 2773 293 2783
rect 613 2783 627 2793
rect 597 2780 627 2783
rect 3687 2797 3713 2803
rect 4233 2803 4247 2813
rect 4233 2800 4263 2803
rect 4237 2797 4263 2800
rect 3353 2783 3367 2792
rect 3560 2783 3573 2787
rect 3353 2780 3423 2783
rect 597 2777 623 2780
rect 3357 2777 3423 2780
rect 277 2726 283 2773
rect 597 2706 603 2777
rect 3417 2747 3423 2777
rect 3557 2773 3573 2783
rect 3827 2777 3853 2783
rect 4127 2783 4140 2787
rect 4160 2783 4173 2787
rect 4127 2780 4143 2783
rect 4127 2773 4147 2780
rect 3557 2747 3563 2773
rect 4133 2766 4147 2773
rect 4157 2773 4173 2783
rect 4257 2783 4263 2797
rect 4287 2797 4333 2803
rect 4437 2797 4513 2803
rect 4257 2777 4283 2783
rect 4157 2747 4163 2773
rect 2547 2737 2573 2743
rect 3417 2737 3433 2747
rect 3420 2733 3433 2737
rect 3557 2737 3573 2747
rect 3560 2733 3573 2737
rect 4157 2737 4173 2747
rect 4160 2733 4173 2737
rect 4277 2743 4283 2777
rect 4257 2737 4283 2743
rect 4437 2747 4443 2797
rect 5097 2797 5133 2803
rect 4927 2777 4963 2783
rect 4957 2747 4963 2777
rect 5097 2747 5103 2797
rect 5420 2783 5433 2787
rect 5417 2773 5433 2783
rect 5827 2783 5840 2787
rect 5827 2773 5843 2783
rect 5417 2747 5423 2773
rect 4437 2737 4453 2747
rect 4257 2707 4263 2737
rect 4440 2733 4453 2737
rect 4957 2737 4973 2747
rect 4960 2733 4973 2737
rect 5097 2737 5113 2747
rect 5100 2733 5113 2737
rect 5417 2737 5433 2747
rect 5420 2733 5433 2737
rect 4287 2717 4333 2723
rect 4427 2717 4473 2723
rect 5387 2717 5453 2723
rect 5837 2723 5843 2773
rect 5837 2717 5893 2723
rect -63 2602 30 2618
rect -63 2098 -3 2602
rect 1747 2517 1853 2523
rect 4107 2517 4133 2523
rect 3727 2497 3773 2503
rect 5007 2497 5083 2503
rect 460 2483 473 2487
rect 457 2473 473 2483
rect 4133 2483 4147 2492
rect 4700 2483 4713 2487
rect 4097 2480 4147 2483
rect 4097 2477 4143 2480
rect 4697 2477 4713 2483
rect 457 2426 463 2473
rect 4097 2447 4103 2477
rect 4700 2473 4713 2477
rect 4907 2483 4920 2487
rect 4907 2473 4923 2483
rect 5027 2483 5040 2487
rect 5027 2473 5043 2483
rect 4547 2457 4603 2463
rect 4917 2447 4923 2473
rect 5037 2447 5043 2473
rect 5077 2463 5083 2497
rect 5407 2497 5453 2503
rect 5667 2497 5793 2503
rect 5397 2483 5403 2493
rect 5397 2477 5423 2483
rect 5077 2457 5103 2463
rect 5206 2457 5253 2463
rect 4087 2437 4103 2447
rect 4087 2433 4100 2437
rect 4907 2437 4923 2447
rect 4907 2433 4920 2437
rect 5027 2437 5043 2447
rect 5417 2447 5423 2477
rect 5417 2437 5433 2447
rect 5027 2433 5040 2437
rect 5420 2433 5433 2437
rect 5983 2358 6043 2862
rect 5950 2342 6043 2358
rect 3227 2277 3273 2283
rect 5227 2277 5293 2283
rect 767 2257 813 2263
rect 3420 2263 3433 2267
rect 3417 2253 3433 2263
rect 3707 2263 3720 2267
rect 3707 2253 3723 2263
rect 3867 2257 3943 2263
rect 4407 2263 4420 2267
rect 4407 2253 4423 2263
rect 4567 2257 4613 2263
rect 4727 2263 4740 2267
rect 4727 2253 4743 2263
rect 4867 2263 4880 2267
rect 5080 2263 5093 2267
rect 4867 2253 4883 2263
rect 3417 2227 3423 2253
rect 3417 2217 3433 2227
rect 3420 2213 3433 2217
rect 1087 2197 1133 2203
rect 3527 2197 3613 2203
rect 3717 2206 3723 2253
rect 4060 2243 4073 2247
rect 4046 2237 4073 2243
rect 4060 2233 4073 2237
rect 4417 2223 4423 2253
rect 4737 2227 4743 2253
rect 4877 2227 4883 2253
rect 4417 2217 4443 2223
rect 4387 2197 4413 2203
rect 4437 2187 4443 2217
rect 4727 2217 4743 2227
rect 4727 2213 4740 2217
rect 4867 2217 4883 2227
rect 5077 2253 5093 2263
rect 5207 2263 5220 2267
rect 5207 2253 5223 2263
rect 5077 2227 5083 2253
rect 5217 2227 5223 2253
rect 5077 2217 5093 2227
rect 4867 2213 4880 2217
rect 5080 2213 5093 2217
rect 5207 2217 5223 2227
rect 5207 2213 5220 2217
rect 5667 2197 5733 2203
rect 3567 2186 3580 2187
rect 4420 2186 4443 2187
rect 3567 2173 3573 2186
rect 4427 2177 4443 2186
rect 4427 2173 4440 2177
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 2867 1977 2913 1983
rect 3127 1977 3233 1983
rect 4867 1977 4893 1983
rect 5067 1977 5113 1983
rect 5527 1977 5573 1983
rect 5767 1977 5853 1983
rect 320 1963 333 1967
rect 317 1953 333 1963
rect 317 1926 323 1953
rect 477 1923 483 1973
rect 500 1963 513 1967
rect 457 1917 483 1923
rect 497 1953 513 1963
rect 2027 1957 2073 1963
rect 4267 1957 4313 1963
rect 4847 1957 4873 1963
rect 5467 1957 5503 1963
rect 497 1927 503 1953
rect 5497 1927 5503 1957
rect 5647 1957 5693 1963
rect 5807 1963 5820 1967
rect 5807 1953 5823 1963
rect 497 1917 513 1927
rect 457 1887 463 1917
rect 500 1913 513 1917
rect 4687 1917 4733 1923
rect 5497 1917 5513 1927
rect 5500 1913 5513 1917
rect 5817 1923 5823 1953
rect 5797 1917 5823 1923
rect 487 1897 553 1903
rect 2987 1897 3073 1903
rect 4107 1897 4193 1903
rect 5797 1887 5803 1917
rect 5827 1897 5873 1903
rect 5983 1838 6043 2342
rect 5950 1822 6043 1838
rect 3947 1797 3973 1803
rect 5667 1797 5693 1803
rect 727 1737 753 1743
rect 2960 1743 2973 1747
rect 2957 1733 2973 1743
rect 4587 1743 4600 1747
rect 4587 1733 4603 1743
rect 4887 1737 4933 1743
rect 5357 1737 5413 1743
rect 2957 1707 2963 1733
rect 4597 1707 4603 1733
rect 5357 1707 5363 1737
rect 5540 1743 5553 1747
rect 5537 1733 5553 1743
rect 2957 1697 2973 1707
rect 2960 1693 2973 1697
rect 4227 1697 4323 1703
rect 4587 1697 4603 1707
rect 4587 1693 4600 1697
rect 5347 1697 5363 1707
rect 5537 1703 5543 1733
rect 5537 1697 5563 1703
rect 5347 1693 5360 1697
rect 4687 1677 4753 1683
rect 4767 1677 4833 1683
rect 5067 1677 5133 1683
rect 5227 1677 5293 1683
rect 5557 1683 5563 1697
rect 5557 1677 5593 1683
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 2767 1457 2793 1463
rect 4087 1457 4113 1463
rect 5087 1457 5153 1463
rect 1133 1443 1147 1453
rect 1133 1440 1163 1443
rect 1137 1437 1163 1440
rect 447 1377 473 1383
rect 1157 1383 1163 1437
rect 3387 1443 3400 1447
rect 3387 1433 3403 1443
rect 4587 1437 4623 1443
rect 3397 1403 3403 1433
rect 4617 1423 4623 1437
rect 5267 1443 5280 1447
rect 5760 1443 5773 1447
rect 5267 1433 5283 1443
rect 4760 1423 4772 1427
rect 4617 1417 4643 1423
rect 4746 1417 4772 1423
rect 4760 1413 4772 1417
rect 4807 1417 4854 1423
rect 5277 1407 5283 1433
rect 5757 1433 5773 1443
rect 5757 1407 5763 1433
rect 3397 1397 3433 1403
rect 4957 1397 5033 1403
rect 5277 1397 5293 1407
rect 5280 1393 5293 1397
rect 5757 1397 5773 1407
rect 5760 1393 5773 1397
rect 1157 1377 1193 1383
rect 3247 1377 3273 1383
rect 5087 1377 5133 1383
rect 4247 1337 4293 1343
rect 5983 1318 6043 1822
rect 5950 1302 6043 1318
rect 5197 1237 5233 1243
rect 1200 1223 1213 1227
rect 1197 1213 1213 1223
rect 2337 1217 2373 1223
rect 5147 1223 5160 1227
rect 5197 1223 5203 1237
rect 5347 1237 5373 1243
rect 5447 1237 5473 1243
rect 5600 1243 5613 1247
rect 5597 1233 5613 1243
rect 5147 1213 5163 1223
rect 1197 1183 1203 1213
rect 2187 1197 2234 1203
rect 5157 1187 5163 1213
rect 1177 1180 1203 1183
rect 1173 1177 1203 1180
rect 1173 1167 1187 1177
rect 5147 1177 5163 1187
rect 5177 1217 5203 1223
rect 5177 1187 5183 1217
rect 5307 1223 5320 1227
rect 5307 1213 5323 1223
rect 5317 1187 5323 1213
rect 5597 1187 5603 1233
rect 5727 1217 5763 1223
rect 5177 1177 5193 1187
rect 5147 1173 5160 1177
rect 5180 1173 5193 1177
rect 5307 1177 5323 1187
rect 5307 1173 5320 1177
rect 5587 1177 5603 1187
rect 5757 1183 5763 1217
rect 5757 1177 5783 1183
rect 5587 1173 5600 1177
rect 5777 1167 5783 1177
rect 887 1157 913 1163
rect 1347 1157 1393 1163
rect 1847 1157 1893 1163
rect 1967 1157 2053 1163
rect 4307 1157 4333 1163
rect 5187 1157 5213 1163
rect 5777 1157 5793 1167
rect 5780 1153 5793 1157
rect 5147 1117 5173 1123
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 533 943 547 953
rect 533 940 563 943
rect 537 937 563 940
rect 557 923 563 937
rect 587 937 613 943
rect 707 937 813 943
rect 1847 937 1873 943
rect 4847 937 4903 943
rect 557 917 583 923
rect 577 863 583 917
rect 3967 917 3993 923
rect 4897 887 4903 937
rect 5327 937 5413 943
rect 5747 937 5853 943
rect 5220 923 5233 927
rect 5027 917 5083 923
rect 5077 887 5083 917
rect 5217 913 5233 923
rect 5520 923 5533 927
rect 5517 913 5533 923
rect 5217 887 5223 913
rect 5517 887 5523 913
rect 4897 877 4913 887
rect 4900 873 4913 877
rect 5077 877 5093 887
rect 5080 873 5093 877
rect 5207 873 5233 887
rect 5517 877 5533 887
rect 5520 873 5533 877
rect 5647 877 5673 883
rect 5907 877 5933 883
rect 547 857 583 863
rect 3467 857 3493 863
rect 3667 857 3793 863
rect 5983 798 6043 1302
rect 5950 782 6043 798
rect 3947 753 3953 767
rect 5247 737 5283 743
rect 4887 703 4900 707
rect 4887 693 4903 703
rect 200 683 213 687
rect 47 677 94 683
rect 197 677 213 683
rect 200 673 213 677
rect 4897 667 4903 693
rect 5097 697 5133 703
rect 5097 683 5103 697
rect 5066 677 5103 683
rect 3387 657 3413 663
rect 4887 657 4903 667
rect 5277 663 5283 737
rect 5467 737 5493 743
rect 5547 717 5583 723
rect 5577 663 5583 717
rect 5707 717 5753 723
rect 5860 703 5873 707
rect 5857 693 5873 703
rect 5277 657 5303 663
rect 5577 657 5603 663
rect 4887 653 4900 657
rect 5107 637 5193 643
rect 5247 637 5273 643
rect 5297 643 5303 657
rect 5597 647 5603 657
rect 5297 637 5333 643
rect 5597 637 5613 647
rect 5600 633 5613 637
rect 5857 643 5863 693
rect 5857 637 5893 643
rect -63 522 30 538
rect -63 18 -3 522
rect 3767 417 3873 423
rect 4667 417 4693 423
rect 5667 417 5713 423
rect 2587 397 2613 403
rect 5787 403 5800 407
rect 5787 393 5803 403
rect 5797 367 5803 393
rect 5237 360 5293 363
rect 5233 357 5293 360
rect 5233 347 5247 357
rect 5787 357 5803 367
rect 5787 353 5800 357
rect 1847 337 1893 343
rect 5983 278 6043 782
rect 5950 262 6043 278
rect 4947 237 4973 243
rect 1107 197 1153 203
rect 4107 197 4143 203
rect 4137 147 4143 197
rect 4137 137 4153 147
rect 4140 133 4153 137
rect 1807 117 1833 123
rect 4707 117 4733 123
rect -63 2 30 18
rect 5983 2 6043 262
<< m2contact >>
rect 4713 5914 4727 5928
rect 4813 5913 4827 5927
rect 3953 5893 3967 5907
rect 3613 5873 3627 5887
rect 1213 5853 1227 5867
rect 2813 5853 2827 5867
rect 2873 5853 2887 5867
rect 3953 5853 3967 5867
rect 2953 5833 2967 5847
rect 3113 5833 3127 5847
rect 4073 5833 4087 5847
rect 4153 5833 4167 5847
rect 4713 5833 4727 5847
rect 4793 5833 4807 5847
rect 4873 5833 4887 5847
rect 5053 5833 5067 5847
rect 5173 5833 5187 5847
rect 2993 5813 3007 5827
rect 3033 5813 3047 5827
rect 4933 5813 4947 5827
rect 1693 5613 1707 5627
rect 1753 5613 1767 5627
rect 2413 5613 2427 5627
rect 2493 5613 2507 5627
rect 2533 5613 2547 5627
rect 4433 5613 4447 5627
rect 4493 5613 4507 5627
rect 4953 5613 4967 5627
rect 5033 5613 5047 5627
rect 5773 5613 5787 5627
rect 5853 5613 5867 5627
rect 5913 5613 5927 5627
rect 5013 5593 5027 5607
rect 5153 5593 5167 5607
rect 3773 5573 3787 5587
rect 3953 5573 3967 5587
rect 3013 5553 3027 5567
rect 3413 5553 3427 5567
rect 5013 5553 5027 5567
rect 2433 5533 2447 5547
rect 2473 5533 2487 5547
rect 2953 5533 2967 5547
rect 3473 5533 3487 5547
rect 5173 5532 5187 5546
rect 133 5373 147 5387
rect 4273 5373 4287 5387
rect 193 5333 207 5347
rect 1513 5333 1527 5347
rect 1573 5333 1587 5347
rect 4333 5333 4347 5347
rect 273 5312 287 5326
rect 353 5313 367 5327
rect 1453 5313 1467 5327
rect 1533 5313 1547 5327
rect 1893 5313 1907 5327
rect 2053 5313 2067 5327
rect 2533 5313 2547 5327
rect 2633 5313 2647 5327
rect 4213 5313 4227 5327
rect 4293 5312 4307 5326
rect 4373 5313 4387 5327
rect 4493 5313 4507 5327
rect 5393 5313 5407 5327
rect 5453 5313 5467 5327
rect 5813 5313 5827 5327
rect 5873 5313 5887 5327
rect 3293 5113 3307 5127
rect 3373 5113 3387 5127
rect 4733 5113 4747 5127
rect 4773 5113 4787 5127
rect 1893 5093 1907 5107
rect 2013 5093 2027 5107
rect 2213 5093 2227 5107
rect 2273 5093 2287 5107
rect 2773 5093 2787 5107
rect 2893 5093 2907 5107
rect 3333 5093 3347 5107
rect 3413 5093 3427 5107
rect 5673 5093 5687 5107
rect 5773 5093 5787 5107
rect 313 5073 327 5087
rect 2713 5073 2727 5087
rect 3813 5073 3827 5087
rect 4033 5073 4047 5087
rect 4453 5073 4467 5087
rect 5053 5073 5067 5087
rect 5533 5073 5547 5087
rect 5613 5073 5627 5087
rect 5713 5073 5727 5087
rect 313 5033 327 5047
rect 2713 5033 2727 5047
rect 3733 5033 3747 5047
rect 4033 5033 4047 5047
rect 4493 5033 4507 5047
rect 5133 5033 5147 5047
rect 5673 5033 5687 5047
rect 4793 5013 4807 5027
rect 4873 5013 4887 5027
rect 3793 4853 3807 4867
rect 5653 4853 5667 4867
rect 273 4813 287 4827
rect 333 4813 347 4827
rect 3793 4813 3807 4827
rect 2053 4793 2067 4807
rect 2133 4793 2147 4807
rect 5313 4793 5327 4807
rect 5433 4793 5447 4807
rect 5713 4853 5727 4867
rect 5713 4813 5727 4827
rect 5813 4813 5827 4827
rect 5933 4813 5947 4827
rect 5733 4793 5747 4807
rect 4273 4773 4287 4787
rect 4353 4773 4367 4787
rect 3593 4653 3607 4667
rect 3633 4653 3647 4667
rect 2773 4633 2787 4647
rect 2813 4633 2827 4647
rect 153 4573 167 4587
rect 1313 4573 1327 4587
rect 313 4553 327 4567
rect 373 4553 387 4567
rect 4333 4573 4347 4587
rect 4453 4573 4467 4587
rect 5653 4573 5667 4587
rect 5713 4573 5727 4587
rect 5773 4573 5787 4587
rect 213 4513 227 4527
rect 1373 4513 1387 4527
rect 2833 4553 2847 4567
rect 3273 4553 3287 4567
rect 3793 4553 3807 4567
rect 3893 4553 3907 4567
rect 3333 4532 3347 4546
rect 4613 4553 4627 4567
rect 5813 4553 5827 4567
rect 2833 4513 2847 4527
rect 3113 4513 3127 4527
rect 3173 4513 3187 4527
rect 3793 4513 3807 4527
rect 3893 4513 3907 4527
rect 4553 4513 4567 4527
rect 5333 4513 5347 4527
rect 5373 4513 5387 4527
rect 5813 4513 5827 4527
rect 5873 4513 5887 4527
rect 2793 4472 2807 4486
rect 2833 4473 2847 4487
rect 793 4453 807 4467
rect 853 4453 867 4467
rect 2313 4453 2327 4467
rect 2353 4453 2367 4467
rect 5633 4393 5647 4407
rect 5673 4393 5687 4407
rect 53 4373 67 4387
rect 93 4373 107 4387
rect 433 4373 447 4387
rect 513 4373 527 4387
rect 2053 4373 2067 4387
rect 2113 4373 2127 4387
rect 553 4354 567 4368
rect 593 4353 607 4367
rect 1373 4353 1387 4367
rect 1433 4353 1447 4367
rect 3633 4353 3647 4367
rect 3713 4353 3727 4367
rect 4533 4353 4547 4367
rect 4613 4354 4627 4368
rect 4693 4353 4707 4367
rect 4993 4354 5007 4368
rect 5073 4353 5087 4367
rect 193 4333 207 4347
rect 2773 4333 2787 4347
rect 193 4293 207 4307
rect 2773 4293 2787 4307
rect 3833 4333 3847 4347
rect 4373 4333 4387 4347
rect 4513 4313 4527 4327
rect 3833 4293 3847 4307
rect 4373 4293 4387 4307
rect 4493 4293 4507 4307
rect 4853 4333 4867 4347
rect 4733 4293 4747 4307
rect 4853 4293 4867 4307
rect 5533 4333 5547 4347
rect 5813 4333 5827 4347
rect 5533 4293 5547 4307
rect 5813 4293 5827 4307
rect 2893 4273 2907 4287
rect 2973 4273 2987 4287
rect 4213 4273 4227 4287
rect 4293 4273 4307 4287
rect 4473 4273 4487 4287
rect 4513 4273 4527 4287
rect 4973 4273 4987 4287
rect 5093 4273 5107 4287
rect 5753 4273 5767 4287
rect 5873 4273 5887 4287
rect 5033 4253 5047 4267
rect 5113 4253 5127 4267
rect 2753 4233 2767 4247
rect 2853 4233 2867 4247
rect 13 4193 27 4207
rect 53 4193 67 4207
rect 4873 4193 4887 4207
rect 4913 4193 4927 4207
rect 573 4113 587 4127
rect 5073 4113 5087 4127
rect 5113 4113 5127 4127
rect 5313 4073 5327 4087
rect 153 4053 167 4067
rect 633 4053 647 4067
rect 2433 4053 2447 4067
rect 2493 4053 2507 4067
rect 2553 4053 2567 4067
rect 1913 4033 1927 4047
rect 373 4013 387 4027
rect 3473 3993 3487 4007
rect 3553 3993 3567 4007
rect 3973 4053 3987 4067
rect 4073 4053 4087 4067
rect 4113 4053 4127 4067
rect 4193 4053 4207 4067
rect 4233 4053 4247 4067
rect 4353 4053 4367 4067
rect 4793 4053 4807 4067
rect 4833 4053 4847 4067
rect 4933 4053 4947 4067
rect 5013 4053 5027 4067
rect 5273 4053 5287 4067
rect 5793 4053 5807 4067
rect 5913 4053 5927 4067
rect 4093 4033 4107 4047
rect 4033 3993 4047 4007
rect 4193 3993 4207 4007
rect 4333 3993 4347 4007
rect 4673 4033 4687 4047
rect 4893 4033 4907 4047
rect 4673 3993 4687 4007
rect 4953 4033 4967 4047
rect 5053 4033 5067 4047
rect 5233 4033 5247 4047
rect 5273 4032 5287 4046
rect 5573 4033 5587 4047
rect 4953 3993 4967 4007
rect 5113 3993 5127 4007
rect 5533 3993 5547 4007
rect 2153 3973 2167 3987
rect 2193 3973 2207 3987
rect 3893 3973 3907 3987
rect 4233 3973 4247 3987
rect 4893 3973 4907 3987
rect 5693 3972 5707 3986
rect 5733 3973 5747 3987
rect 5233 3953 5247 3967
rect 5313 3953 5327 3967
rect 5533 3873 5547 3887
rect 4913 3853 4927 3867
rect 3313 3833 3327 3847
rect 3393 3833 3407 3847
rect 4833 3833 4847 3847
rect 5353 3833 5367 3847
rect 153 3813 167 3827
rect 4453 3813 4467 3827
rect 4613 3813 4627 3827
rect 4713 3813 4727 3827
rect 5033 3813 5047 3827
rect 5213 3813 5227 3827
rect 5333 3813 5347 3827
rect 213 3773 227 3787
rect 3873 3773 3887 3787
rect 3913 3773 3927 3787
rect 4453 3773 4467 3787
rect 4553 3773 4567 3787
rect 4713 3773 4727 3787
rect 4993 3773 5007 3787
rect 5393 3792 5407 3806
rect 5213 3773 5227 3787
rect 5333 3773 5347 3787
rect 313 3753 327 3767
rect 393 3753 407 3767
rect 1033 3753 1047 3767
rect 1113 3753 1127 3767
rect 1213 3753 1227 3767
rect 1253 3753 1267 3767
rect 5133 3753 5147 3767
rect 5253 3753 5267 3767
rect 5573 3753 5587 3767
rect 293 3673 307 3687
rect 353 3673 367 3687
rect 3033 3553 3047 3567
rect 3093 3553 3107 3567
rect 4013 3553 4027 3567
rect 4073 3553 4087 3567
rect 873 3533 887 3547
rect 913 3533 927 3547
rect 2013 3533 2027 3547
rect 2073 3533 2087 3547
rect 3293 3534 3307 3548
rect 3393 3533 3407 3547
rect 4573 3533 4587 3547
rect 4613 3533 4627 3547
rect 3313 3513 3327 3527
rect 3853 3513 3867 3527
rect 353 3493 367 3507
rect 3313 3473 3327 3487
rect 3933 3513 3947 3527
rect 5133 3513 5147 3527
rect 5213 3513 5227 3527
rect 3933 3473 3947 3487
rect 5053 3473 5067 3487
rect 5213 3473 5227 3487
rect 5393 3473 5407 3487
rect 1873 3453 1887 3467
rect 1933 3453 1947 3467
rect 2493 3453 2507 3467
rect 2553 3453 2567 3467
rect 5333 3453 5347 3467
rect 5613 3453 5627 3467
rect 5693 3453 5707 3467
rect 3173 3433 3187 3447
rect 3213 3413 3227 3427
rect 4633 3353 4647 3367
rect 2213 3333 2227 3347
rect 2253 3333 2267 3347
rect 4693 3333 4707 3347
rect 1333 3313 1347 3327
rect 1413 3313 1427 3327
rect 3873 3313 3887 3327
rect 4513 3313 4527 3327
rect 4553 3313 4567 3327
rect 4833 3313 4847 3327
rect 4913 3313 4927 3327
rect 5273 3313 5287 3327
rect 5373 3313 5387 3327
rect 4033 3293 4047 3307
rect 5793 3293 5807 3307
rect 5893 3293 5907 3307
rect 1193 3253 1207 3267
rect 1253 3253 1267 3267
rect 3933 3253 3947 3267
rect 4073 3253 4087 3267
rect 5793 3253 5807 3267
rect 5893 3253 5907 3267
rect 3913 3233 3927 3247
rect 3953 3233 3967 3247
rect 4153 3233 4167 3247
rect 4253 3231 4267 3245
rect 4633 3233 4647 3247
rect 4713 3233 4727 3247
rect 5113 3233 5127 3247
rect 5213 3233 5227 3247
rect 5453 3233 5467 3247
rect 5513 3233 5527 3247
rect 2733 3213 2747 3227
rect 2833 3213 2847 3227
rect 3893 3213 3907 3227
rect 3933 3213 3947 3227
rect 5113 3212 5127 3226
rect 5153 3213 5167 3227
rect 5673 3053 5687 3067
rect 5713 3053 5727 3067
rect 3973 3014 3987 3028
rect 4053 3012 4067 3026
rect 4893 3013 4907 3027
rect 5013 3013 5027 3027
rect 5253 3013 5267 3027
rect 753 2993 767 3007
rect 793 2973 807 2987
rect 5553 2993 5567 3007
rect 5613 2993 5627 3007
rect 5693 2993 5707 3007
rect 5253 2973 5267 2987
rect 5433 2953 5447 2967
rect 5893 3013 5907 3027
rect 5193 2933 5207 2947
rect 5753 2933 5767 2947
rect 5913 2933 5927 2947
rect 4233 2813 4247 2827
rect 613 2793 627 2807
rect 713 2793 727 2807
rect 793 2793 807 2807
rect 293 2773 307 2787
rect 3353 2792 3367 2806
rect 3673 2793 3687 2807
rect 3713 2793 3727 2807
rect 273 2712 287 2726
rect 3573 2773 3587 2787
rect 3813 2773 3827 2787
rect 3853 2773 3867 2787
rect 4113 2773 4127 2787
rect 4133 2752 4147 2766
rect 4173 2773 4187 2787
rect 4273 2793 4287 2807
rect 4333 2793 4347 2807
rect 2533 2733 2547 2747
rect 2573 2733 2587 2747
rect 3433 2733 3447 2747
rect 3573 2733 3587 2747
rect 4173 2733 4187 2747
rect 4513 2793 4527 2807
rect 4913 2773 4927 2787
rect 5133 2793 5147 2807
rect 5433 2773 5447 2787
rect 5813 2773 5827 2787
rect 4453 2733 4467 2747
rect 4973 2733 4987 2747
rect 5113 2733 5127 2747
rect 5433 2733 5447 2747
rect 4273 2713 4287 2727
rect 4333 2713 4347 2727
rect 4413 2713 4427 2727
rect 4473 2713 4487 2727
rect 5373 2713 5387 2727
rect 5453 2713 5467 2727
rect 5893 2711 5907 2725
rect 593 2692 607 2706
rect 4253 2693 4267 2707
rect 1733 2513 1747 2527
rect 1853 2513 1867 2527
rect 4093 2513 4107 2527
rect 4133 2513 4147 2527
rect 3713 2493 3727 2507
rect 3773 2493 3787 2507
rect 4133 2492 4147 2506
rect 4993 2493 5007 2507
rect 473 2473 487 2487
rect 4713 2473 4727 2487
rect 4893 2473 4907 2487
rect 5013 2473 5027 2487
rect 4533 2453 4547 2467
rect 5393 2493 5407 2507
rect 5453 2493 5467 2507
rect 5653 2493 5667 2507
rect 5793 2493 5807 2507
rect 5253 2453 5267 2467
rect 4073 2433 4087 2447
rect 4893 2433 4907 2447
rect 5013 2433 5027 2447
rect 5433 2433 5447 2447
rect 453 2412 467 2426
rect 3213 2273 3227 2287
rect 3273 2273 3287 2287
rect 5213 2273 5227 2287
rect 5293 2274 5307 2288
rect 753 2253 767 2267
rect 813 2253 827 2267
rect 3433 2253 3447 2267
rect 3693 2253 3707 2267
rect 3853 2253 3867 2267
rect 4393 2253 4407 2267
rect 4553 2253 4567 2267
rect 4613 2253 4627 2267
rect 4713 2253 4727 2267
rect 4853 2253 4867 2267
rect 3433 2213 3447 2227
rect 1073 2193 1087 2207
rect 1133 2193 1147 2207
rect 3513 2193 3527 2207
rect 3613 2193 3627 2207
rect 4073 2233 4087 2247
rect 3713 2192 3727 2206
rect 4373 2193 4387 2207
rect 4413 2193 4427 2207
rect 4713 2213 4727 2227
rect 4853 2213 4867 2227
rect 5093 2253 5107 2267
rect 5193 2253 5207 2267
rect 5093 2213 5107 2227
rect 5193 2213 5207 2227
rect 5653 2193 5667 2207
rect 5733 2193 5747 2207
rect 3553 2173 3567 2187
rect 3573 2172 3587 2186
rect 4413 2172 4427 2186
rect 3993 2113 4007 2127
rect 473 1973 487 1987
rect 2853 1973 2867 1987
rect 2913 1973 2927 1987
rect 3113 1973 3127 1987
rect 3233 1973 3247 1987
rect 4853 1973 4867 1987
rect 4893 1973 4907 1987
rect 5053 1973 5067 1987
rect 5113 1973 5127 1987
rect 5513 1973 5527 1987
rect 5573 1973 5587 1987
rect 5753 1973 5767 1987
rect 5853 1973 5867 1987
rect 333 1953 347 1967
rect 313 1912 327 1926
rect 513 1953 527 1967
rect 2013 1953 2027 1967
rect 2073 1953 2087 1967
rect 4253 1953 4267 1967
rect 4313 1953 4327 1967
rect 4833 1953 4847 1967
rect 4873 1953 4887 1967
rect 5453 1953 5467 1967
rect 5633 1953 5647 1967
rect 5693 1953 5707 1967
rect 5793 1953 5807 1967
rect 513 1913 527 1927
rect 4673 1913 4687 1927
rect 4733 1913 4747 1927
rect 5513 1913 5527 1927
rect 473 1893 487 1907
rect 553 1893 567 1907
rect 2973 1893 2987 1907
rect 3073 1893 3087 1907
rect 4093 1893 4107 1907
rect 4193 1893 4207 1907
rect 5813 1893 5827 1907
rect 5873 1893 5887 1907
rect 453 1873 467 1887
rect 5793 1873 5807 1887
rect 3933 1793 3947 1807
rect 3973 1793 3987 1807
rect 5653 1793 5667 1807
rect 5693 1793 5707 1807
rect 713 1733 727 1747
rect 753 1733 767 1747
rect 2973 1733 2987 1747
rect 4573 1733 4587 1747
rect 4873 1733 4887 1747
rect 4933 1733 4947 1747
rect 5413 1733 5427 1747
rect 5553 1733 5567 1747
rect 2973 1693 2987 1707
rect 4213 1693 4227 1707
rect 4573 1693 4587 1707
rect 5333 1693 5347 1707
rect 4673 1673 4687 1687
rect 4753 1673 4767 1687
rect 4833 1673 4847 1687
rect 5053 1673 5067 1687
rect 5133 1671 5147 1685
rect 5213 1673 5227 1687
rect 5293 1673 5307 1687
rect 5593 1673 5607 1687
rect 1133 1453 1147 1467
rect 2753 1453 2767 1467
rect 2793 1454 2807 1468
rect 4073 1453 4087 1467
rect 4113 1453 4127 1467
rect 5073 1454 5087 1468
rect 5153 1453 5167 1467
rect 433 1373 447 1387
rect 473 1373 487 1387
rect 3373 1433 3387 1447
rect 4573 1433 4587 1447
rect 5253 1433 5267 1447
rect 4772 1413 4786 1427
rect 4793 1413 4807 1427
rect 5773 1433 5787 1447
rect 3433 1393 3447 1407
rect 5033 1393 5047 1407
rect 5293 1393 5307 1407
rect 5773 1393 5787 1407
rect 1193 1371 1207 1385
rect 3233 1372 3247 1386
rect 3273 1373 3287 1387
rect 5073 1373 5087 1387
rect 5133 1373 5147 1387
rect 4233 1333 4247 1347
rect 4293 1333 4307 1347
rect 1213 1213 1227 1227
rect 2373 1213 2387 1227
rect 5133 1213 5147 1227
rect 5233 1233 5247 1247
rect 5333 1233 5347 1247
rect 5373 1233 5387 1247
rect 5433 1234 5447 1248
rect 5473 1233 5487 1247
rect 5613 1233 5627 1247
rect 2173 1193 2187 1207
rect 5133 1173 5147 1187
rect 5293 1213 5307 1227
rect 5713 1213 5727 1227
rect 5193 1173 5207 1187
rect 5293 1173 5307 1187
rect 5573 1173 5587 1187
rect 873 1153 887 1167
rect 913 1153 927 1167
rect 1173 1153 1187 1167
rect 1333 1153 1347 1167
rect 1393 1153 1407 1167
rect 1833 1153 1847 1167
rect 1893 1153 1907 1167
rect 1953 1153 1967 1167
rect 2053 1153 2067 1167
rect 4293 1153 4307 1167
rect 4333 1153 4347 1167
rect 5173 1153 5187 1167
rect 5213 1151 5227 1165
rect 5793 1153 5807 1167
rect 5133 1113 5147 1127
rect 5173 1113 5187 1127
rect 2273 1073 2287 1087
rect 533 953 547 967
rect 573 933 587 947
rect 613 934 627 948
rect 693 933 707 947
rect 813 933 827 947
rect 1833 933 1847 947
rect 1873 933 1887 947
rect 4833 933 4847 947
rect 533 853 547 867
rect 3953 913 3967 927
rect 3993 913 4007 927
rect 5313 932 5327 946
rect 5413 933 5427 947
rect 5733 933 5747 947
rect 5853 933 5867 947
rect 5013 913 5027 927
rect 5233 913 5247 927
rect 5533 913 5547 927
rect 4913 873 4927 887
rect 5093 873 5107 887
rect 5193 873 5207 887
rect 5233 873 5247 887
rect 5533 873 5547 887
rect 5633 873 5647 887
rect 5673 873 5687 887
rect 5893 873 5907 887
rect 5933 873 5947 887
rect 3453 853 3467 867
rect 3493 853 3507 867
rect 3653 853 3667 867
rect 3793 853 3807 867
rect 3933 753 3947 767
rect 3953 753 3967 767
rect 5233 733 5247 747
rect 4873 693 4887 707
rect 33 673 47 687
rect 213 673 227 687
rect 5133 693 5147 707
rect 3373 653 3387 667
rect 3413 653 3427 667
rect 4873 653 4887 667
rect 5453 733 5467 747
rect 5493 733 5507 747
rect 5533 714 5547 728
rect 5693 713 5707 727
rect 5753 713 5767 727
rect 5873 693 5887 707
rect 5093 633 5107 647
rect 5193 633 5207 647
rect 5233 633 5247 647
rect 5273 633 5287 647
rect 5333 633 5347 647
rect 5613 633 5627 647
rect 5893 633 5907 647
rect 5013 553 5027 567
rect 3753 413 3767 427
rect 3873 413 3887 427
rect 4653 413 4667 427
rect 4693 413 4707 427
rect 5653 413 5667 427
rect 5713 413 5727 427
rect 2573 393 2587 407
rect 2613 393 2627 407
rect 5773 393 5787 407
rect 5293 353 5307 367
rect 5773 353 5787 367
rect 1833 333 1847 347
rect 1893 333 1907 347
rect 5233 333 5247 347
rect 4933 233 4947 247
rect 4973 232 4987 246
rect 1093 193 1107 207
rect 1153 193 1167 207
rect 4093 193 4107 207
rect 4153 133 4167 147
rect 1793 113 1807 127
rect 1833 113 1847 127
rect 4693 113 4707 127
rect 4733 113 4747 127
<< metal2 >>
rect 816 6007 824 6044
rect 2936 6007 2944 6044
rect 3536 6007 3544 6044
rect 4696 6007 4704 6044
rect 4716 6036 4744 6044
rect 156 5607 164 5913
rect 213 5900 227 5913
rect 216 5896 224 5900
rect 376 5867 384 5896
rect 720 5864 733 5867
rect 56 5507 64 5553
rect 96 5527 104 5553
rect 96 5376 104 5492
rect 136 5387 144 5513
rect 16 4207 24 5113
rect 36 4467 44 5374
rect 76 5340 84 5344
rect 73 5327 87 5340
rect 116 5207 124 5344
rect 56 4867 64 5073
rect 96 4856 104 4993
rect 56 4816 73 4824
rect 16 3827 24 4172
rect 16 3727 24 3773
rect 36 3627 44 4413
rect 56 4387 64 4816
rect 96 4556 104 4613
rect 136 4556 144 4653
rect 156 4587 164 5553
rect 176 5327 184 5852
rect 196 5566 204 5593
rect 236 5467 244 5564
rect 316 5560 324 5564
rect 256 5387 264 5533
rect 276 5347 284 5493
rect 196 5088 204 5333
rect 236 5127 244 5332
rect 213 4860 227 4873
rect 216 4856 224 4860
rect 276 4827 284 5312
rect 296 5207 304 5553
rect 313 5547 327 5560
rect 376 5467 384 5853
rect 416 5604 424 5864
rect 476 5860 484 5864
rect 473 5847 487 5860
rect 516 5627 524 5833
rect 656 5747 664 5864
rect 716 5860 733 5864
rect 713 5853 733 5860
rect 836 5860 844 5864
rect 713 5847 727 5853
rect 833 5847 847 5860
rect 916 5847 924 5993
rect 2447 5956 2473 5964
rect 1116 5896 1124 5933
rect 1316 5896 1324 5933
rect 1216 5867 1224 5893
rect 1516 5866 1524 5933
rect 1636 5896 1644 5933
rect 396 5596 424 5604
rect 516 5604 524 5613
rect 496 5596 524 5604
rect 396 5404 404 5596
rect 376 5396 404 5404
rect 376 5376 384 5396
rect 356 5340 364 5344
rect 396 5340 404 5344
rect 456 5340 464 5344
rect 353 5327 367 5340
rect 393 5327 407 5340
rect 453 5327 467 5340
rect 316 5087 324 5313
rect 516 5287 524 5344
rect 556 5327 564 5613
rect 656 5596 664 5693
rect 716 5566 724 5733
rect 833 5600 847 5613
rect 836 5596 844 5600
rect 596 5507 604 5564
rect 676 5560 684 5564
rect 673 5547 687 5560
rect 736 5427 744 5594
rect 776 5544 784 5564
rect 776 5536 804 5544
rect 576 5388 584 5413
rect 696 5344 704 5374
rect 696 5336 724 5344
rect 296 5047 304 5074
rect 356 5076 364 5193
rect 556 5127 564 5313
rect 533 5080 547 5093
rect 536 5076 544 5080
rect 327 5044 340 5047
rect 327 5036 344 5044
rect 327 5033 340 5036
rect 376 4868 384 5044
rect 436 4887 444 5053
rect 516 4907 524 5044
rect 576 5007 584 5093
rect 296 4587 304 4653
rect 316 4567 324 4613
rect 300 4564 313 4567
rect 296 4556 313 4564
rect 196 4527 204 4554
rect 300 4553 313 4556
rect 116 4387 124 4524
rect 227 4524 240 4527
rect 227 4516 244 4524
rect 227 4513 240 4516
rect 96 4336 104 4373
rect 156 4347 164 4512
rect 116 4267 124 4304
rect 56 3747 64 4193
rect 96 4036 104 4133
rect 156 4067 164 4193
rect 156 4036 164 4053
rect 176 4047 184 4373
rect 196 4347 204 4453
rect 216 4336 224 4373
rect 96 3828 104 3973
rect 116 3947 124 4004
rect 136 3816 144 3933
rect 156 3827 164 3853
rect 116 3547 124 3784
rect 176 3607 184 3993
rect 196 3967 204 4293
rect 216 4007 224 4233
rect 276 4167 284 4524
rect 296 4306 304 4493
rect 336 4467 344 4813
rect 356 4667 364 4824
rect 416 4604 424 4853
rect 436 4627 444 4873
rect 493 4860 507 4873
rect 496 4856 504 4860
rect 536 4856 544 4933
rect 476 4820 484 4824
rect 473 4807 487 4820
rect 516 4804 524 4824
rect 516 4796 544 4804
rect 396 4596 424 4604
rect 356 4387 364 4573
rect 396 4567 404 4596
rect 413 4560 427 4573
rect 480 4564 493 4567
rect 416 4556 424 4560
rect 476 4556 493 4564
rect 480 4553 493 4556
rect 376 4487 384 4553
rect 376 4336 384 4413
rect 396 4387 404 4513
rect 436 4487 444 4524
rect 436 4306 444 4373
rect 396 4296 424 4304
rect 296 3867 304 3964
rect 116 3304 124 3484
rect 176 3447 184 3514
rect 196 3387 204 3853
rect 316 3827 324 4004
rect 376 3967 384 4013
rect 216 3647 224 3773
rect 316 3767 324 3792
rect 336 3786 344 3933
rect 396 3907 404 4273
rect 416 4067 424 4296
rect 456 4247 464 4513
rect 476 4287 484 4453
rect 516 4387 524 4613
rect 536 4527 544 4796
rect 576 4564 584 4893
rect 596 4607 604 5073
rect 716 5047 724 5336
rect 796 5207 804 5536
rect 856 5487 864 5564
rect 896 5507 904 5613
rect 916 5467 924 5833
rect 996 5596 1004 5653
rect 1016 5647 1024 5693
rect 1136 5687 1144 5844
rect 1296 5787 1304 5864
rect 1336 5827 1344 5864
rect 976 5560 984 5564
rect 973 5547 987 5560
rect 856 5388 864 5413
rect 636 4947 644 5032
rect 676 4927 684 5044
rect 736 4944 744 5113
rect 816 5007 824 5044
rect 856 4987 864 5293
rect 876 5047 884 5332
rect 916 5307 924 5344
rect 956 5287 964 5374
rect 976 5307 984 5453
rect 996 5347 1004 5513
rect 1053 5380 1067 5393
rect 1076 5384 1084 5673
rect 1156 5596 1164 5773
rect 1336 5608 1344 5813
rect 1476 5707 1484 5864
rect 1536 5827 1544 5893
rect 1576 5787 1584 5864
rect 1616 5827 1624 5864
rect 1496 5647 1504 5673
rect 1136 5507 1144 5564
rect 1236 5527 1244 5573
rect 1276 5487 1284 5564
rect 1376 5527 1384 5573
rect 1516 5567 1524 5773
rect 1656 5707 1664 5864
rect 1536 5564 1544 5594
rect 1536 5556 1564 5564
rect 1596 5560 1604 5564
rect 1436 5527 1444 5552
rect 1056 5376 1064 5380
rect 1076 5376 1104 5384
rect 1096 5127 1104 5376
rect 1116 5147 1124 5373
rect 736 4936 764 4944
rect 656 4856 664 4913
rect 636 4820 644 4824
rect 633 4807 647 4820
rect 756 4787 764 4936
rect 776 4827 784 4893
rect 876 4787 884 4824
rect 556 4556 584 4564
rect 556 4368 564 4556
rect 636 4520 644 4524
rect 633 4507 647 4520
rect 696 4367 704 4593
rect 756 4487 764 4524
rect 796 4467 804 4513
rect 513 4340 527 4352
rect 516 4336 524 4340
rect 536 4107 544 4304
rect 576 4127 584 4153
rect 416 3848 424 4053
rect 496 3960 504 3964
rect 493 3947 507 3960
rect 316 3707 324 3753
rect 256 3516 264 3693
rect 356 3687 364 3833
rect 536 3816 544 3913
rect 556 3887 564 4021
rect 576 3927 584 4092
rect 576 3816 584 3853
rect 596 3847 604 4353
rect 716 4336 724 4393
rect 616 4147 624 4334
rect 656 4267 664 4304
rect 616 4047 624 4133
rect 636 4127 644 4193
rect 633 4040 647 4053
rect 636 4036 644 4040
rect 396 3780 404 3784
rect 376 3747 384 3772
rect 393 3767 407 3780
rect 636 3784 644 3833
rect 376 3687 384 3712
rect 296 3516 304 3673
rect 356 3507 364 3652
rect 556 3627 564 3784
rect 516 3527 524 3593
rect 596 3587 604 3784
rect 616 3776 644 3784
rect 616 3567 624 3776
rect 636 3527 644 3753
rect 656 3627 664 3853
rect 676 3767 684 3873
rect 696 3827 704 3953
rect 736 3947 744 4034
rect 716 3816 724 3873
rect 756 3824 764 4353
rect 776 4147 784 4393
rect 816 4347 824 4773
rect 916 4727 924 4856
rect 876 4568 884 4713
rect 836 4507 844 4554
rect 856 4367 864 4453
rect 856 4336 864 4353
rect 893 4340 907 4353
rect 896 4336 904 4340
rect 836 4247 844 4304
rect 956 4207 964 4973
rect 976 4867 984 4933
rect 996 4927 1004 5073
rect 1016 4947 1024 5113
rect 1116 5047 1124 5074
rect 1056 5007 1064 5044
rect 1136 5044 1144 5293
rect 1156 5267 1164 5344
rect 1196 5088 1204 5332
rect 1236 5267 1244 5393
rect 1296 5307 1304 5344
rect 1236 5076 1244 5133
rect 1136 5036 1164 5044
rect 1067 4996 1084 5004
rect 993 4884 1007 4892
rect 993 4880 1024 4884
rect 996 4876 1024 4880
rect 1016 4856 1024 4876
rect 1076 4864 1084 4996
rect 1076 4856 1104 4864
rect 996 4527 1004 4824
rect 1036 4556 1044 4753
rect 1056 4567 1064 4793
rect 1156 4724 1164 5036
rect 1176 4767 1184 4993
rect 1216 4887 1224 5044
rect 1256 4967 1264 5044
rect 1296 5024 1304 5113
rect 1316 5047 1324 5253
rect 1396 5088 1404 5373
rect 1500 5344 1513 5347
rect 1456 5327 1464 5344
rect 1496 5336 1513 5344
rect 1500 5333 1513 5336
rect 1536 5327 1544 5533
rect 1556 5427 1564 5556
rect 1593 5547 1607 5560
rect 1676 5564 1684 5594
rect 1696 5567 1704 5613
rect 1656 5556 1684 5564
rect 1556 5344 1564 5413
rect 1556 5336 1573 5344
rect 1587 5344 1600 5347
rect 1587 5336 1604 5344
rect 1587 5333 1600 5336
rect 1456 5224 1464 5313
rect 1656 5307 1664 5556
rect 1716 5564 1724 5953
rect 1796 5896 1804 5953
rect 2076 5896 2084 5953
rect 2116 5907 2124 5933
rect 1776 5747 1784 5864
rect 1916 5647 1924 5864
rect 1753 5600 1767 5613
rect 1756 5596 1764 5600
rect 1796 5596 1804 5633
rect 1936 5596 1944 5633
rect 1976 5608 1984 5852
rect 1716 5556 1744 5564
rect 1736 5376 1744 5556
rect 1776 5527 1784 5564
rect 1876 5376 1884 5594
rect 2016 5566 2024 5773
rect 2096 5647 2104 5852
rect 2156 5787 2164 5953
rect 2213 5900 2227 5913
rect 2236 5907 2244 5953
rect 2216 5896 2224 5900
rect 2093 5600 2107 5612
rect 2136 5607 2144 5633
rect 2096 5596 2104 5600
rect 2116 5507 2124 5564
rect 1916 5376 1924 5473
rect 1716 5267 1724 5344
rect 1756 5307 1764 5332
rect 1456 5216 1484 5224
rect 1436 5076 1444 5113
rect 1296 5016 1324 5024
rect 1276 4787 1284 4824
rect 1316 4787 1324 5016
rect 1336 4868 1344 5073
rect 1416 4987 1424 5044
rect 1396 4856 1404 4953
rect 1476 4927 1484 5216
rect 1796 5127 1804 5374
rect 1976 5346 1984 5473
rect 2033 5388 2047 5393
rect 2156 5387 2164 5613
rect 2176 5567 2184 5733
rect 2256 5624 2264 5913
rect 2456 5896 2464 5933
rect 2276 5827 2284 5893
rect 2336 5687 2344 5864
rect 2247 5616 2264 5624
rect 2233 5600 2247 5613
rect 2236 5596 2244 5600
rect 2336 5544 2344 5613
rect 2356 5567 2364 5793
rect 2396 5747 2404 5894
rect 2636 5896 2644 5953
rect 2596 5866 2604 5893
rect 2476 5807 2484 5864
rect 2516 5787 2524 5864
rect 2656 5860 2664 5864
rect 2653 5847 2667 5860
rect 2696 5807 2704 5864
rect 2716 5787 2724 5833
rect 2736 5807 2744 5894
rect 2800 5864 2813 5867
rect 2796 5856 2813 5864
rect 2800 5853 2813 5856
rect 2413 5600 2427 5613
rect 2416 5596 2424 5600
rect 2456 5596 2464 5633
rect 2436 5560 2444 5564
rect 2316 5536 2344 5544
rect 2433 5547 2447 5560
rect 2193 5380 2207 5393
rect 2296 5388 2304 5433
rect 2196 5376 2204 5380
rect 2296 5347 2304 5374
rect 1896 5340 1904 5344
rect 1893 5327 1907 5340
rect 2056 5327 2064 5344
rect 1596 5076 1604 5113
rect 1536 4987 1544 5044
rect 1636 4987 1644 5074
rect 1496 4824 1504 4973
rect 1576 4856 1584 4913
rect 1416 4787 1424 4824
rect 1456 4816 1504 4824
rect 1136 4716 1164 4724
rect 1116 4527 1124 4554
rect 1076 4427 1084 4524
rect 976 4307 984 4373
rect 1116 4304 1124 4334
rect 1096 4296 1124 4304
rect 1076 4267 1084 4290
rect 836 4036 844 4133
rect 856 4107 864 4173
rect 916 4004 924 4193
rect 1096 4147 1104 4296
rect 1136 4187 1144 4716
rect 1416 4624 1424 4773
rect 1556 4764 1564 4824
rect 1656 4787 1664 5053
rect 1756 5007 1764 5044
rect 1796 4987 1804 5033
rect 1736 4856 1744 4973
rect 1716 4804 1724 4812
rect 1716 4796 1744 4804
rect 1573 4764 1587 4773
rect 1556 4760 1587 4764
rect 1556 4756 1584 4760
rect 1396 4616 1424 4624
rect 1313 4560 1327 4573
rect 1316 4556 1324 4560
rect 1356 4556 1364 4593
rect 1196 4467 1204 4524
rect 1256 4507 1264 4553
rect 1216 4336 1224 4373
rect 1196 4284 1204 4304
rect 1236 4284 1244 4304
rect 1176 4276 1204 4284
rect 1216 4276 1244 4284
rect 1176 4247 1184 4276
rect 1216 4264 1224 4276
rect 1196 4256 1224 4264
rect 976 4036 984 4113
rect 1036 4006 1044 4073
rect 916 3996 944 4004
rect 756 3816 784 3824
rect 856 3816 864 3853
rect 896 3824 904 3993
rect 896 3816 924 3824
rect 736 3587 744 3772
rect 776 3667 784 3816
rect 836 3780 844 3784
rect 833 3767 847 3780
rect 607 3524 620 3527
rect 607 3513 624 3524
rect 660 3524 673 3527
rect 656 3516 673 3524
rect 660 3513 673 3516
rect 736 3524 744 3552
rect 716 3516 744 3524
rect 116 3296 144 3304
rect 136 3264 144 3296
rect 16 3260 44 3264
rect 16 3256 47 3260
rect 16 3044 24 3256
rect 33 3247 47 3256
rect 16 3036 33 3044
rect 36 2996 44 3033
rect 96 3024 104 3193
rect 76 3020 104 3024
rect 73 3016 104 3020
rect 73 3007 87 3016
rect 86 3000 87 3007
rect 136 2907 144 2996
rect 136 2744 144 2813
rect 36 2707 44 2744
rect 156 2707 164 3033
rect 256 2707 264 3373
rect 336 3296 344 3433
rect 276 3267 284 3296
rect 296 3256 313 3264
rect 276 2747 284 2950
rect 296 2787 304 3256
rect 373 3000 387 3013
rect 416 3004 424 3413
rect 436 3027 444 3444
rect 476 3404 484 3433
rect 496 3427 504 3452
rect 476 3396 504 3404
rect 496 3296 504 3396
rect 616 3287 624 3513
rect 756 3307 764 3613
rect 916 3587 924 3816
rect 836 3516 844 3573
rect 873 3520 887 3533
rect 876 3516 884 3520
rect 776 3447 784 3513
rect 916 3487 924 3533
rect 856 3447 864 3484
rect 936 3447 944 3996
rect 956 3827 964 4004
rect 976 3816 984 3853
rect 1016 3816 1024 3933
rect 1056 3827 1064 4113
rect 1096 4067 1104 4133
rect 1096 4036 1104 4053
rect 1176 4007 1184 4193
rect 996 3780 1004 3784
rect 1036 3780 1044 3784
rect 993 3767 1007 3780
rect 1033 3767 1047 3780
rect 1076 3767 1084 3993
rect 1096 3667 1104 3813
rect 1116 3767 1124 3833
rect 1173 3820 1187 3833
rect 1196 3827 1204 4256
rect 1236 4127 1244 4253
rect 1276 4207 1284 4413
rect 1296 4267 1304 4524
rect 1336 4520 1344 4524
rect 1333 4507 1347 4520
rect 1376 4427 1384 4513
rect 1373 4340 1387 4353
rect 1396 4347 1404 4616
rect 1376 4336 1384 4340
rect 1236 4067 1244 4113
rect 1256 4036 1264 4073
rect 1313 4040 1327 4053
rect 1316 4036 1324 4040
rect 1176 3816 1184 3820
rect 1216 3767 1224 3873
rect 1236 3827 1244 4004
rect 1276 3887 1284 4004
rect 1396 3964 1404 3992
rect 1416 3987 1424 4513
rect 1456 4447 1464 4524
rect 1436 4367 1444 4393
rect 1476 4387 1484 4493
rect 1536 4447 1544 4593
rect 1556 4344 1564 4613
rect 1576 4527 1584 4756
rect 1656 4556 1664 4633
rect 1676 4467 1684 4524
rect 1716 4447 1724 4554
rect 1736 4507 1744 4796
rect 1756 4567 1764 4812
rect 1796 4556 1804 4893
rect 1816 4827 1824 5074
rect 1836 5047 1844 5253
rect 2056 5167 2064 5313
rect 2216 5307 2224 5344
rect 1893 5088 1907 5093
rect 1936 5076 1973 5084
rect 2013 5080 2027 5093
rect 2016 5076 2024 5080
rect 2096 5087 2104 5293
rect 1916 4987 1924 5032
rect 1976 5007 1984 5074
rect 1836 4627 1844 4933
rect 2036 4856 2044 5032
rect 2116 4987 2124 5153
rect 1896 4820 1904 4824
rect 1893 4807 1907 4820
rect 2053 4807 2067 4812
rect 2093 4807 2107 4812
rect 2136 4807 2144 5093
rect 2176 5076 2184 5233
rect 2256 5207 2264 5344
rect 2316 5287 2324 5536
rect 2473 5547 2487 5552
rect 2276 5107 2284 5213
rect 2213 5080 2227 5093
rect 2256 5096 2273 5104
rect 2216 5076 2224 5080
rect 2196 4907 2204 5044
rect 2196 4884 2204 4893
rect 2176 4876 2204 4884
rect 2176 4856 2184 4876
rect 1936 4556 1944 4713
rect 2056 4604 2064 4793
rect 2236 4787 2244 4893
rect 2256 4727 2264 5096
rect 2296 4884 2304 5073
rect 2396 5046 2404 5133
rect 2296 4876 2324 4884
rect 2316 4868 2324 4876
rect 2356 4856 2364 4973
rect 2396 4868 2404 5032
rect 2036 4596 2064 4604
rect 1776 4520 1784 4524
rect 1773 4507 1787 4520
rect 1876 4407 1884 4512
rect 1556 4336 1584 4344
rect 1436 4087 1444 4332
rect 1476 4147 1484 4304
rect 1436 4007 1444 4036
rect 1496 3996 1524 4004
rect 1516 3967 1524 3996
rect 1396 3956 1424 3964
rect 1273 3820 1287 3833
rect 1336 3824 1344 3873
rect 1276 3816 1284 3820
rect 1336 3816 1364 3824
rect 1256 3780 1264 3784
rect 1253 3767 1267 3780
rect 1176 3627 1184 3753
rect 1256 3667 1264 3753
rect 1416 3707 1424 3956
rect 1536 3927 1544 4073
rect 976 3528 984 3593
rect 1196 3567 1204 3653
rect 1056 3476 1084 3484
rect 1056 3347 1064 3476
rect 1136 3387 1144 3514
rect 1256 3516 1264 3553
rect 1156 3367 1164 3513
rect 636 3264 644 3293
rect 476 3244 484 3252
rect 476 3236 504 3244
rect 496 3008 504 3236
rect 516 3027 524 3252
rect 736 3260 744 3264
rect 733 3247 747 3260
rect 376 2996 384 3000
rect 416 2996 444 3004
rect 336 2776 344 2933
rect 356 2907 364 2964
rect 396 2746 404 2952
rect 436 2784 444 2996
rect 456 2966 464 2993
rect 536 2960 544 2964
rect 416 2776 444 2784
rect 456 2776 464 2952
rect 533 2947 547 2960
rect 496 2776 504 2813
rect 416 2746 424 2776
rect 556 2746 564 2813
rect 296 2736 313 2744
rect 156 2507 164 2693
rect 33 2480 47 2493
rect 36 2476 44 2480
rect 136 2387 144 2476
rect 156 2227 164 2493
rect 216 2440 224 2444
rect 213 2427 227 2440
rect 256 2424 264 2633
rect 236 2416 264 2424
rect 236 2264 244 2416
rect 216 2256 244 2264
rect 36 2204 44 2210
rect 16 2196 44 2204
rect 16 2047 24 2196
rect 96 2187 104 2224
rect 256 2207 264 2393
rect 276 2287 284 2712
rect 296 2264 304 2736
rect 376 2476 384 2693
rect 396 2687 404 2732
rect 276 2256 304 2264
rect 336 2256 344 2413
rect 356 2387 364 2444
rect 276 2144 284 2256
rect 396 2226 404 2432
rect 436 2387 444 2693
rect 576 2587 584 3013
rect 776 3004 784 3313
rect 767 2996 784 3004
rect 656 2887 664 2964
rect 756 2927 764 2993
rect 796 2987 804 3333
rect 893 3300 907 3313
rect 896 3296 904 3300
rect 1136 3296 1144 3333
rect 916 3067 924 3264
rect 956 3008 964 3293
rect 1076 3266 1084 3293
rect 1196 3267 1204 3433
rect 1296 3427 1304 3573
rect 1316 3486 1324 3653
rect 1376 3516 1384 3553
rect 1416 3447 1424 3613
rect 933 2966 947 2981
rect 676 2847 684 2924
rect 976 2887 984 3053
rect 1036 3008 1044 3033
rect 1176 2996 1184 3133
rect 713 2807 727 2813
rect 596 2727 604 2793
rect 613 2787 627 2793
rect 693 2780 707 2793
rect 696 2776 704 2780
rect 736 2746 744 2833
rect 807 2804 820 2807
rect 807 2793 824 2804
rect 816 2776 824 2793
rect 616 2736 644 2744
rect 616 2707 624 2736
rect 756 2727 764 2753
rect 996 2747 1004 2813
rect 1016 2790 1024 2953
rect 1136 2947 1144 2964
rect 796 2740 804 2744
rect 793 2727 807 2740
rect 596 2607 604 2692
rect 456 2447 464 2513
rect 476 2487 484 2573
rect 536 2476 544 2513
rect 636 2487 644 2713
rect 316 2207 324 2224
rect 276 2136 304 2144
rect 96 1956 104 2033
rect 96 1527 104 1704
rect 196 1706 204 2033
rect 236 1956 244 2033
rect 96 1487 104 1513
rect 36 1436 44 1473
rect 56 967 64 1313
rect 116 1216 124 1393
rect 136 1327 144 1693
rect 156 1287 164 1533
rect 236 1307 244 1353
rect 276 1327 284 2113
rect 296 1907 304 2136
rect 316 1947 324 2193
rect 336 1980 404 1984
rect 333 1976 404 1980
rect 333 1967 347 1976
rect 396 1956 404 1976
rect 436 1956 444 2153
rect 456 1964 464 2412
rect 516 2387 524 2444
rect 513 2260 527 2273
rect 516 2256 524 2260
rect 556 2256 564 2433
rect 656 2264 664 2533
rect 696 2476 704 2593
rect 753 2480 767 2493
rect 756 2476 764 2480
rect 636 2256 664 2264
rect 636 2226 644 2256
rect 496 2187 504 2212
rect 536 2204 544 2224
rect 516 2196 544 2204
rect 516 2147 524 2196
rect 473 1987 487 1993
rect 456 1956 484 1964
rect 416 1920 424 1924
rect 296 1404 304 1673
rect 316 1444 324 1912
rect 413 1907 427 1920
rect 476 1907 484 1956
rect 416 1736 424 1793
rect 336 1467 344 1693
rect 356 1587 364 1704
rect 396 1700 404 1704
rect 393 1687 407 1700
rect 316 1436 344 1444
rect 373 1440 387 1453
rect 376 1436 384 1440
rect 156 1216 164 1273
rect 136 947 144 1184
rect 36 607 44 673
rect 56 27 64 913
rect 196 887 204 1293
rect 296 1227 304 1390
rect 356 1367 364 1404
rect 436 1387 444 1573
rect 456 1487 464 1873
rect 496 1748 504 2093
rect 516 1967 524 2053
rect 536 1968 544 2173
rect 576 2167 584 2224
rect 556 2047 564 2113
rect 576 1956 584 1993
rect 616 1956 624 2153
rect 676 2067 684 2224
rect 556 1920 564 1924
rect 513 1907 527 1913
rect 553 1907 567 1920
rect 676 1736 684 1793
rect 716 1747 724 1953
rect 736 1748 744 2053
rect 756 1964 764 2253
rect 776 2226 784 2253
rect 796 2067 804 2713
rect 836 2687 844 2744
rect 896 2740 904 2744
rect 893 2727 907 2740
rect 816 2327 824 2473
rect 836 2407 844 2652
rect 856 2507 864 2713
rect 916 2436 944 2444
rect 936 2407 944 2436
rect 813 2267 827 2273
rect 896 2256 904 2313
rect 836 2067 844 2113
rect 936 2107 944 2393
rect 956 2027 964 2513
rect 976 2287 984 2473
rect 1016 2387 1024 2444
rect 1056 2440 1064 2444
rect 1053 2427 1067 2440
rect 996 2220 1004 2224
rect 993 2207 1007 2220
rect 856 1964 864 2013
rect 756 1956 784 1964
rect 836 1956 864 1964
rect 893 1960 907 1973
rect 896 1956 904 1960
rect 996 1867 1004 2153
rect 1036 2147 1044 2224
rect 1076 2207 1084 2273
rect 1096 2267 1104 2732
rect 1136 2667 1144 2933
rect 1216 2927 1224 3293
rect 1236 3227 1244 3353
rect 1296 3296 1304 3353
rect 1333 3307 1347 3313
rect 1156 2547 1164 2913
rect 1236 2907 1244 2994
rect 1256 2927 1264 3253
rect 1316 3187 1324 3264
rect 1356 3247 1364 3433
rect 1436 3347 1444 3913
rect 1556 3824 1564 4133
rect 1576 4067 1584 4336
rect 1596 4267 1604 4353
rect 1673 4340 1687 4353
rect 1793 4340 1807 4353
rect 1676 4336 1684 4340
rect 1796 4336 1804 4340
rect 1836 4336 1844 4393
rect 1656 4227 1664 4304
rect 1776 4227 1784 4304
rect 1576 4036 1624 4044
rect 1653 4040 1667 4053
rect 1656 4036 1664 4040
rect 1576 3927 1584 4036
rect 1676 4000 1684 4004
rect 1673 3987 1687 4000
rect 1556 3816 1584 3824
rect 1476 3547 1484 3784
rect 1536 3747 1544 3784
rect 1576 3767 1584 3816
rect 1596 3787 1604 3953
rect 1656 3816 1664 3913
rect 1576 3607 1584 3753
rect 1496 3516 1504 3553
rect 1533 3520 1547 3533
rect 1536 3516 1544 3520
rect 1476 3447 1484 3484
rect 1376 3187 1384 3313
rect 1396 3266 1404 3333
rect 1413 3307 1427 3313
rect 1456 3296 1464 3353
rect 1516 3307 1524 3353
rect 1436 3227 1444 3264
rect 1316 3147 1324 3173
rect 1336 2996 1344 3033
rect 1216 2776 1224 2873
rect 1316 2827 1324 2964
rect 1396 2867 1404 3053
rect 1433 3008 1447 3013
rect 1476 2996 1484 3053
rect 1516 3007 1524 3252
rect 1536 3107 1544 3413
rect 1576 3407 1584 3533
rect 1596 3447 1604 3513
rect 1616 3467 1624 3693
rect 1676 3667 1684 3784
rect 1716 3664 1724 3973
rect 1736 3707 1744 4173
rect 1896 4147 1904 4554
rect 1916 4306 1924 4353
rect 1936 4107 1944 4493
rect 1956 4467 1964 4524
rect 2016 4507 2024 4554
rect 2036 4527 2044 4596
rect 2076 4556 2084 4613
rect 1956 4347 1964 4453
rect 1993 4340 2007 4353
rect 1996 4336 2004 4340
rect 2036 4336 2044 4433
rect 2096 4407 2104 4453
rect 2156 4447 2164 4633
rect 2176 4427 2184 4613
rect 2196 4587 2204 4653
rect 2216 4556 2224 4613
rect 2376 4568 2384 4673
rect 2396 4604 2404 4854
rect 2416 4627 2424 5233
rect 2436 5087 2444 5453
rect 2476 5376 2484 5533
rect 2496 5467 2504 5613
rect 2516 5607 2524 5773
rect 2533 5600 2547 5613
rect 2536 5596 2544 5600
rect 2576 5596 2584 5633
rect 2636 5527 2644 5633
rect 2656 5547 2664 5613
rect 2753 5600 2767 5613
rect 2756 5596 2764 5600
rect 2516 5376 2524 5433
rect 2496 5307 2504 5344
rect 2536 5340 2544 5344
rect 2533 5327 2547 5340
rect 2496 5187 2504 5293
rect 2453 5080 2467 5093
rect 2456 5076 2464 5080
rect 2496 5076 2504 5133
rect 2496 4856 2504 4993
rect 2516 4907 2524 5044
rect 2476 4747 2484 4812
rect 2516 4787 2524 4824
rect 2556 4767 2564 5173
rect 2576 5147 2584 5374
rect 2596 5347 2604 5453
rect 2656 5376 2664 5473
rect 2676 5467 2684 5553
rect 2696 5388 2704 5564
rect 2716 5504 2724 5533
rect 2736 5527 2744 5564
rect 2716 5496 2744 5504
rect 2636 5327 2644 5344
rect 2596 4907 2604 5273
rect 2636 5076 2644 5313
rect 2676 5187 2684 5332
rect 2736 5207 2744 5496
rect 2796 5467 2804 5833
rect 2756 5287 2764 5453
rect 2776 5387 2784 5413
rect 2816 5376 2824 5793
rect 2876 5707 2884 5853
rect 2896 5847 2904 5993
rect 2953 5847 2967 5852
rect 3036 5827 3044 5894
rect 3276 5896 3284 5933
rect 3176 5866 3184 5893
rect 3116 5860 3124 5864
rect 2856 5607 2864 5693
rect 2896 5596 2904 5633
rect 2936 5596 2944 5693
rect 2953 5547 2967 5552
rect 2696 5047 2704 5193
rect 2776 5107 2784 5213
rect 2727 5084 2740 5087
rect 2727 5076 2744 5084
rect 2773 5080 2787 5093
rect 2776 5076 2784 5080
rect 2727 5073 2740 5076
rect 2576 4787 2584 4854
rect 2636 4804 2644 4824
rect 2616 4796 2644 4804
rect 2616 4747 2624 4796
rect 2396 4596 2424 4604
rect 2416 4556 2424 4596
rect 2496 4587 2504 4633
rect 2453 4560 2467 4573
rect 2456 4556 2464 4560
rect 2316 4467 2324 4533
rect 2053 4387 2067 4393
rect 2127 4373 2133 4387
rect 2016 4247 2024 4304
rect 1796 3967 1804 4004
rect 1796 3816 1804 3893
rect 1816 3847 1824 3964
rect 1896 3867 1904 4093
rect 1976 4036 1984 4213
rect 1916 3927 1924 4033
rect 1956 3967 1964 4004
rect 1996 3927 2004 4004
rect 2056 3927 2064 4293
rect 2076 4247 2084 4373
rect 2136 4247 2144 4304
rect 2196 4227 2204 4433
rect 2276 4336 2284 4393
rect 2153 4040 2167 4053
rect 2156 4036 2164 4040
rect 2256 4036 2264 4304
rect 2296 4300 2304 4304
rect 2293 4287 2307 4300
rect 2336 4167 2344 4553
rect 2356 4307 2364 4453
rect 2376 4187 2384 4453
rect 2396 4348 2404 4473
rect 2436 4467 2444 4524
rect 2496 4404 2504 4573
rect 2516 4526 2524 4593
rect 2556 4556 2564 4593
rect 2596 4556 2604 4633
rect 2636 4487 2644 4773
rect 2656 4527 2664 4653
rect 2716 4647 2724 5033
rect 2776 4868 2784 4973
rect 2816 4867 2824 5273
rect 2836 5207 2844 5344
rect 2836 5088 2844 5133
rect 2876 5084 2884 5453
rect 2936 5376 2944 5513
rect 2976 5507 2984 5594
rect 2996 5547 3004 5813
rect 3076 5684 3084 5852
rect 3113 5847 3127 5860
rect 3076 5676 3093 5684
rect 3096 5596 3104 5673
rect 3116 5608 3124 5833
rect 3196 5807 3204 5894
rect 3296 5860 3304 5864
rect 3293 5847 3307 5860
rect 3336 5847 3344 5893
rect 3476 5787 3484 5893
rect 3616 5887 3624 5933
rect 3756 5896 3764 5953
rect 3136 5567 3144 5633
rect 3236 5596 3244 5633
rect 3356 5596 3364 5633
rect 3027 5564 3040 5567
rect 3027 5556 3044 5564
rect 3076 5560 3084 5564
rect 3027 5553 3040 5556
rect 3073 5547 3087 5560
rect 3256 5527 3264 5564
rect 2896 5267 2904 5374
rect 3036 5346 3044 5393
rect 3096 5376 3104 5513
rect 3296 5487 3304 5594
rect 3436 5567 3444 5633
rect 3336 5527 3344 5564
rect 3376 5560 3384 5564
rect 3373 5547 3387 5560
rect 3413 5547 3427 5553
rect 3476 5547 3484 5773
rect 3516 5707 3524 5864
rect 3636 5847 3644 5893
rect 3676 5873 3693 5887
rect 3676 5787 3684 5873
rect 3816 5844 3824 5993
rect 4716 5984 4724 6036
rect 4687 5976 4724 5984
rect 3953 5907 3967 5913
rect 3836 5847 3844 5894
rect 3976 5866 3984 5893
rect 3736 5747 3744 5844
rect 3796 5836 3824 5844
rect 3736 5687 3744 5733
rect 3616 5608 3624 5633
rect 3556 5527 3564 5564
rect 3133 5380 3147 5393
rect 3136 5376 3144 5380
rect 3196 5346 3204 5413
rect 3436 5376 3444 5473
rect 3576 5467 3584 5493
rect 3596 5487 3604 5553
rect 3616 5504 3624 5594
rect 3636 5567 3644 5673
rect 3696 5596 3704 5633
rect 3773 5567 3787 5573
rect 3716 5527 3724 5564
rect 3616 5496 3644 5504
rect 3636 5467 3644 5496
rect 3756 5487 3764 5553
rect 3776 5507 3784 5532
rect 3516 5387 3524 5413
rect 3596 5376 3604 5413
rect 3696 5388 3704 5433
rect 3736 5376 3784 5384
rect 2956 5307 2964 5344
rect 3116 5267 3124 5344
rect 3196 5307 3204 5332
rect 3256 5267 3264 5344
rect 3316 5247 3324 5344
rect 3416 5247 3424 5344
rect 3456 5304 3464 5332
rect 3456 5296 3484 5304
rect 2896 5107 2904 5213
rect 2856 5076 2884 5084
rect 2756 4667 2764 4824
rect 2796 4816 2824 4824
rect 2776 4607 2784 4633
rect 2776 4567 2784 4593
rect 2756 4487 2764 4524
rect 2496 4396 2524 4404
rect 2453 4344 2467 4353
rect 2436 4340 2467 4344
rect 2436 4336 2464 4340
rect 2476 4267 2484 4304
rect 2516 4267 2524 4396
rect 2313 4040 2327 4053
rect 2396 4048 2404 4093
rect 2316 4036 2324 4040
rect 2433 4040 2447 4053
rect 2436 4036 2444 4040
rect 2136 3927 2144 4004
rect 2153 3967 2167 3973
rect 2176 3944 2184 3993
rect 2207 3973 2213 3987
rect 2276 3947 2284 4004
rect 2176 3936 2193 3944
rect 1776 3780 1784 3784
rect 1773 3767 1787 3780
rect 1716 3656 1733 3664
rect 1660 3484 1673 3487
rect 1656 3480 1673 3484
rect 1653 3473 1673 3480
rect 1653 3467 1667 3473
rect 1596 3347 1604 3433
rect 1676 3367 1684 3433
rect 1616 3187 1624 3264
rect 1596 2967 1604 3093
rect 1456 2927 1464 2964
rect 1527 2956 1544 2964
rect 1516 2788 1524 2953
rect 1256 2776 1304 2784
rect 1296 2707 1304 2776
rect 1316 2747 1324 2774
rect 1136 2387 1144 2444
rect 1176 2287 1184 2444
rect 1216 2347 1224 2433
rect 1236 2427 1244 2473
rect 1256 2387 1264 2613
rect 1276 2447 1284 2633
rect 1376 2627 1384 2744
rect 1436 2707 1444 2773
rect 1316 2407 1324 2444
rect 1356 2440 1364 2444
rect 1353 2427 1367 2440
rect 1396 2440 1404 2444
rect 1096 2207 1104 2253
rect 1136 2220 1144 2224
rect 1133 2207 1147 2220
rect 1176 2187 1184 2224
rect 1216 2147 1224 2273
rect 1256 2256 1264 2293
rect 1236 2067 1244 2113
rect 1276 2067 1284 2224
rect 1316 2067 1324 2333
rect 1336 2187 1344 2293
rect 1376 2256 1384 2433
rect 1393 2427 1407 2440
rect 1456 2407 1464 2773
rect 1556 2667 1564 2774
rect 1576 2744 1584 2853
rect 1616 2847 1624 3013
rect 1636 3004 1644 3253
rect 1656 3027 1664 3333
rect 1676 3267 1684 3332
rect 1696 3187 1704 3413
rect 1736 3327 1744 3653
rect 1856 3587 1864 3833
rect 2196 3816 2204 3933
rect 1936 3707 1944 3784
rect 1756 3427 1764 3573
rect 1836 3516 1844 3553
rect 1816 3407 1824 3484
rect 1876 3467 1884 3593
rect 1936 3480 1944 3484
rect 1873 3447 1887 3453
rect 1756 3296 1764 3333
rect 1793 3300 1807 3313
rect 1796 3296 1804 3300
rect 1756 3164 1764 3213
rect 1776 3187 1784 3264
rect 1796 3207 1804 3233
rect 1756 3156 1784 3164
rect 1736 3004 1744 3093
rect 1636 2996 1664 3004
rect 1716 2996 1764 3004
rect 1576 2736 1593 2744
rect 1596 2684 1604 2733
rect 1616 2707 1624 2744
rect 1596 2676 1624 2684
rect 1476 2427 1484 2653
rect 1596 2484 1604 2533
rect 1576 2476 1604 2484
rect 1596 2407 1604 2433
rect 1616 2367 1624 2676
rect 1636 2446 1644 2553
rect 1656 2488 1664 2693
rect 1736 2567 1744 2833
rect 1756 2744 1764 2996
rect 1776 2867 1784 3156
rect 1896 3087 1904 3473
rect 1933 3467 1947 3480
rect 1996 3447 2004 3772
rect 2076 3747 2084 3784
rect 2176 3747 2184 3784
rect 2216 3767 2224 3784
rect 2207 3756 2224 3767
rect 2207 3753 2220 3756
rect 2076 3567 2084 3733
rect 2016 3464 2024 3533
rect 2036 3484 2044 3553
rect 2073 3547 2087 3553
rect 2096 3516 2104 3593
rect 2276 3587 2284 3813
rect 2356 3727 2364 3784
rect 2396 3744 2404 3973
rect 2416 3967 2424 4004
rect 2476 3824 2484 4153
rect 2536 4067 2544 4433
rect 2576 4407 2584 4453
rect 2596 4336 2604 4373
rect 2676 4348 2684 4393
rect 2736 4336 2744 4473
rect 2776 4347 2784 4513
rect 2796 4507 2804 4753
rect 2816 4747 2824 4816
rect 2836 4807 2844 5074
rect 2856 4947 2864 5076
rect 3076 5076 3084 5173
rect 3116 5167 3124 5213
rect 2936 4947 2944 5044
rect 2976 4987 2984 5044
rect 2856 4784 2864 4854
rect 2836 4776 2864 4784
rect 2816 4647 2824 4733
rect 2553 4067 2567 4073
rect 2496 4006 2504 4053
rect 2536 4036 2544 4053
rect 2576 4036 2584 4213
rect 2616 4036 2624 4133
rect 2656 4007 2664 4173
rect 2596 3947 2604 4004
rect 2387 3736 2404 3744
rect 2456 3816 2484 3824
rect 2036 3476 2064 3484
rect 2016 3456 2044 3464
rect 1916 3310 1924 3433
rect 2036 3307 2044 3456
rect 1916 3127 1924 3296
rect 1956 3207 1964 3264
rect 1813 3000 1827 3013
rect 1816 2996 1824 3000
rect 1836 2907 1844 2964
rect 1916 2960 1924 2964
rect 1736 2527 1744 2553
rect 1756 2547 1764 2730
rect 1716 2407 1724 2444
rect 1416 2220 1424 2224
rect 1413 2207 1427 2220
rect 1416 2167 1424 2193
rect 1456 2167 1464 2293
rect 1536 2256 1544 2353
rect 1496 2207 1504 2254
rect 1133 1970 1147 1973
rect 1196 1956 1244 1964
rect 1436 1956 1444 2053
rect 1476 1956 1524 1964
rect 756 1706 764 1733
rect 916 1707 924 1734
rect 536 1667 544 1704
rect 536 1547 544 1653
rect 696 1627 704 1704
rect 707 1616 724 1624
rect 476 1400 484 1404
rect 473 1387 487 1400
rect 536 1367 544 1434
rect 616 1436 624 1473
rect 653 1440 667 1453
rect 656 1436 664 1440
rect 556 1406 564 1433
rect 716 1406 724 1616
rect 836 1487 844 1704
rect 936 1627 944 1833
rect 956 1747 964 1853
rect 1016 1847 1024 1956
rect 1076 1916 1104 1924
rect 1096 1887 1104 1916
rect 996 1736 1004 1773
rect 976 1667 984 1704
rect 1116 1527 1124 1913
rect 1236 1887 1244 1956
rect 1516 1927 1524 1956
rect 1316 1916 1344 1924
rect 276 1180 284 1184
rect 273 1167 287 1180
rect 316 1167 324 1273
rect 316 967 324 1153
rect 236 916 244 953
rect 140 884 153 887
rect 136 876 153 884
rect 140 873 153 876
rect 336 867 344 1214
rect 356 1186 364 1313
rect 456 1216 464 1353
rect 496 1167 504 1313
rect 536 1216 544 1332
rect 636 1327 644 1404
rect 676 1367 684 1404
rect 656 1307 664 1333
rect 836 1327 844 1452
rect 856 1227 864 1513
rect 1136 1484 1144 1833
rect 1336 1807 1344 1916
rect 1276 1704 1284 1733
rect 1236 1696 1264 1704
rect 1256 1527 1264 1696
rect 1296 1667 1304 1713
rect 1316 1706 1324 1773
rect 1456 1706 1464 1924
rect 1476 1747 1484 1873
rect 1536 1867 1544 2193
rect 1616 2087 1624 2313
rect 1716 2256 1724 2372
rect 1756 2268 1764 2333
rect 1656 2220 1664 2224
rect 1653 2207 1667 2220
rect 1756 2224 1764 2254
rect 1736 2216 1764 2224
rect 1576 1956 1584 2073
rect 1616 1956 1624 2033
rect 1716 1927 1724 2193
rect 1516 1736 1524 1833
rect 1556 1736 1564 1813
rect 1536 1667 1544 1704
rect 1136 1476 1164 1484
rect 1056 1436 1064 1473
rect 1133 1448 1147 1453
rect 536 967 544 1153
rect 496 916 504 953
rect 556 944 564 1172
rect 596 1147 604 1184
rect 536 936 564 944
rect 536 916 544 936
rect 627 936 693 944
rect 136 736 144 853
rect 296 696 304 733
rect 213 667 227 673
rect 116 487 124 593
rect 116 396 124 473
rect 356 396 364 473
rect 376 447 384 853
rect 416 704 424 913
rect 576 887 584 933
rect 656 880 664 884
rect 653 867 667 880
rect 396 696 424 704
rect 396 547 404 696
rect 416 627 424 653
rect 416 427 424 613
rect 436 587 444 664
rect 476 487 484 664
rect 176 364 184 393
rect 96 267 104 364
rect 136 356 184 364
rect 216 327 224 364
rect 96 207 104 253
rect 216 227 224 313
rect 156 146 164 213
rect 256 187 264 364
rect 316 267 324 293
rect 416 284 424 364
rect 436 307 444 353
rect 456 284 464 394
rect 476 287 484 433
rect 496 324 504 653
rect 516 647 524 733
rect 536 567 544 853
rect 576 696 584 753
rect 616 708 624 853
rect 656 827 664 853
rect 716 767 724 933
rect 596 660 604 664
rect 593 647 607 660
rect 573 400 587 413
rect 616 407 624 553
rect 576 396 584 400
rect 556 360 564 364
rect 553 347 567 360
rect 596 344 604 364
rect 576 336 604 344
rect 576 324 584 336
rect 496 316 584 324
rect 616 307 624 353
rect 636 347 644 493
rect 656 427 664 753
rect 756 408 764 953
rect 776 887 784 1184
rect 876 1167 884 1433
rect 916 1367 924 1404
rect 956 1367 964 1404
rect 956 1307 964 1353
rect 896 1147 904 1213
rect 1016 1186 1024 1353
rect 813 920 827 933
rect 816 916 824 920
rect 776 667 784 694
rect 776 587 784 653
rect 796 647 804 694
rect 916 567 924 1153
rect 976 1027 984 1184
rect 996 944 1004 1133
rect 1036 1047 1044 1392
rect 1076 1384 1084 1404
rect 1056 1376 1084 1384
rect 987 936 1004 944
rect 976 916 984 933
rect 956 827 964 884
rect 1056 747 1064 1376
rect 1156 1367 1164 1476
rect 1276 1427 1284 1613
rect 1200 1385 1220 1387
rect 1207 1373 1213 1385
rect 1116 1216 1124 1313
rect 1156 1307 1164 1353
rect 1236 1347 1244 1404
rect 1156 1216 1164 1293
rect 1136 1127 1144 1184
rect 1173 1167 1187 1172
rect 1196 1067 1204 1333
rect 1213 1227 1227 1233
rect 1276 1180 1284 1184
rect 1273 1167 1287 1180
rect 1316 1167 1324 1353
rect 1336 1167 1344 1653
rect 1376 1587 1384 1653
rect 1376 1436 1384 1573
rect 1596 1507 1604 1793
rect 1616 1627 1624 1713
rect 1636 1607 1644 1873
rect 1676 1736 1684 1833
rect 1716 1787 1724 1913
rect 1736 1887 1744 2216
rect 1776 2207 1784 2493
rect 1796 2387 1804 2744
rect 1856 2527 1864 2613
rect 1896 2567 1904 2953
rect 1913 2947 1927 2960
rect 1976 2887 1984 2994
rect 1996 2927 2004 3153
rect 2036 3147 2044 3193
rect 2056 3167 2064 3476
rect 2076 3187 2084 3484
rect 2116 3447 2124 3484
rect 2136 3476 2164 3484
rect 2116 3296 2124 3433
rect 2136 3387 2144 3476
rect 2153 3300 2167 3313
rect 2196 3307 2204 3373
rect 2216 3347 2224 3493
rect 2156 3296 2164 3300
rect 2180 3264 2193 3267
rect 2016 3047 2024 3113
rect 2116 3107 2124 3233
rect 2136 3187 2144 3264
rect 2176 3256 2193 3264
rect 2180 3253 2193 3256
rect 2216 3247 2224 3312
rect 2116 3004 2124 3093
rect 2096 2996 2124 3004
rect 2116 2884 2124 2953
rect 2136 2907 2144 3073
rect 2116 2876 2144 2884
rect 1976 2776 1984 2852
rect 2036 2746 2044 2813
rect 2136 2776 2144 2876
rect 2176 2784 2184 3173
rect 2216 2996 2224 3053
rect 2236 3027 2244 3573
rect 2336 3516 2344 3553
rect 2256 3407 2264 3473
rect 2256 3287 2264 3333
rect 2316 3296 2324 3393
rect 2356 3347 2364 3433
rect 2376 3324 2384 3733
rect 2396 3387 2404 3573
rect 2416 3487 2424 3713
rect 2456 3707 2464 3816
rect 2456 3516 2464 3633
rect 2496 3587 2504 3784
rect 2576 3747 2584 3893
rect 2596 3827 2604 3933
rect 2676 3784 2684 4334
rect 2696 3907 2704 4292
rect 2716 4267 2724 4304
rect 2716 4147 2724 4253
rect 2776 4247 2784 4293
rect 2736 4036 2744 4233
rect 2756 4167 2764 4233
rect 2796 3864 2804 4472
rect 2816 4447 2824 4612
rect 2836 4567 2844 4776
rect 2856 4556 2864 4653
rect 2896 4556 2904 4793
rect 2916 4747 2924 4824
rect 3016 4727 3024 5032
rect 3056 4987 3064 5044
rect 3076 4856 3084 4893
rect 3136 4864 3144 5113
rect 3156 4947 3164 5173
rect 3213 5080 3227 5093
rect 3216 5076 3224 5080
rect 3296 5047 3304 5113
rect 3196 5007 3204 5044
rect 3287 5036 3304 5047
rect 3287 5033 3300 5036
rect 3127 4856 3144 4864
rect 3056 4647 3064 4824
rect 3096 4767 3104 4824
rect 2836 4487 2844 4513
rect 2876 4504 2884 4524
rect 2976 4524 2984 4554
rect 2996 4527 3004 4633
rect 3053 4560 3067 4573
rect 3056 4556 3064 4560
rect 2956 4516 2984 4524
rect 2876 4496 2904 4504
rect 2853 4484 2867 4493
rect 2853 4480 2884 4484
rect 2856 4476 2884 4480
rect 2816 4306 2824 4353
rect 2836 4347 2844 4452
rect 2876 4336 2884 4476
rect 2896 4367 2904 4496
rect 2896 4300 2904 4304
rect 2816 4087 2824 4292
rect 2893 4287 2907 4300
rect 2936 4264 2944 4493
rect 2956 4287 2964 4516
rect 3036 4520 3044 4524
rect 3033 4507 3047 4520
rect 3136 4524 3144 4812
rect 3156 4767 3164 4893
rect 3176 4787 3184 4953
rect 3196 4868 3204 4933
rect 3156 4647 3164 4713
rect 3276 4707 3284 4854
rect 3296 4824 3304 4993
rect 3316 4887 3324 5074
rect 3336 5044 3344 5093
rect 3376 5076 3384 5113
rect 3413 5080 3427 5093
rect 3416 5076 3424 5080
rect 3476 5047 3484 5296
rect 3676 5267 3684 5344
rect 3336 5036 3364 5044
rect 3356 4856 3364 5036
rect 3396 5007 3404 5044
rect 3496 5007 3504 5073
rect 3476 4856 3484 4933
rect 3516 4867 3524 5213
rect 3676 5144 3684 5173
rect 3696 5167 3704 5293
rect 3716 5227 3724 5253
rect 3776 5247 3784 5376
rect 3676 5136 3713 5144
rect 3696 5076 3704 5113
rect 3736 5087 3744 5233
rect 3296 4816 3324 4824
rect 3127 4516 3144 4524
rect 3116 4487 3124 4513
rect 3156 4507 3164 4633
rect 3213 4560 3227 4573
rect 3216 4556 3224 4560
rect 3273 4567 3287 4573
rect 3296 4527 3304 4773
rect 3187 4524 3200 4527
rect 3187 4516 3204 4524
rect 3187 4513 3200 4516
rect 2976 4287 2984 4373
rect 3036 4336 3044 4413
rect 3056 4367 3064 4453
rect 3073 4340 3087 4353
rect 3096 4347 3104 4413
rect 3076 4336 3084 4340
rect 2936 4256 2964 4264
rect 2836 4147 2844 4193
rect 2856 4187 2864 4233
rect 2916 4167 2924 4193
rect 2896 4107 2904 4133
rect 2787 3856 2804 3864
rect 2616 3747 2624 3784
rect 2656 3776 2684 3784
rect 2596 3607 2604 3653
rect 2616 3627 2624 3693
rect 2476 3467 2484 3484
rect 2536 3467 2544 3514
rect 2556 3467 2564 3533
rect 2616 3516 2624 3613
rect 2656 3507 2664 3776
rect 2676 3687 2684 3733
rect 2696 3727 2704 3853
rect 2776 3816 2784 3853
rect 2836 3828 2844 4093
rect 2876 4036 2884 4073
rect 2956 4004 2964 4256
rect 3096 4247 3104 4292
rect 3116 4267 3124 4473
rect 3136 4427 3144 4492
rect 3196 4336 3204 4493
rect 3236 4347 3244 4453
rect 2916 4000 2924 4004
rect 2913 3987 2927 4000
rect 2936 3996 2964 4004
rect 2836 3707 2844 3814
rect 2936 3784 2944 3996
rect 2976 3987 2984 4093
rect 3016 4048 3024 4113
rect 3096 4004 3104 4233
rect 3136 4187 3144 4333
rect 3176 4127 3184 4292
rect 3216 4287 3224 4304
rect 3196 4036 3204 4253
rect 3216 4227 3224 4273
rect 3256 4207 3264 4473
rect 3316 4367 3324 4816
rect 3336 4567 3344 4824
rect 3376 4687 3384 4824
rect 3416 4567 3424 4853
rect 3456 4767 3464 4824
rect 3436 4556 3444 4613
rect 3336 4487 3344 4532
rect 3396 4516 3413 4524
rect 3476 4524 3484 4733
rect 3496 4567 3504 4824
rect 3536 4584 3544 5033
rect 3576 5007 3584 5044
rect 3616 5007 3624 5074
rect 3756 5047 3764 5113
rect 3676 4967 3684 5044
rect 3556 4747 3564 4913
rect 3613 4860 3627 4873
rect 3616 4856 3624 4860
rect 3596 4727 3604 4824
rect 3676 4707 3684 4893
rect 3606 4672 3607 4680
rect 3593 4667 3607 4672
rect 3536 4576 3584 4584
rect 3576 4556 3584 4576
rect 3616 4526 3624 4673
rect 3636 4667 3644 4693
rect 3696 4687 3704 4933
rect 3736 4907 3744 5033
rect 3756 4856 3764 4993
rect 3776 4987 3784 5074
rect 3796 4867 3804 5836
rect 3836 5747 3844 5833
rect 3956 5587 3964 5853
rect 3976 5667 3984 5852
rect 4016 5827 4024 5933
rect 4096 5896 4104 5933
rect 4276 5896 4284 5933
rect 4456 5907 4464 5933
rect 4076 5860 4084 5864
rect 4073 5847 4087 5860
rect 4156 5847 4164 5893
rect 4336 5866 4344 5893
rect 4476 5866 4484 5913
rect 4536 5896 4544 5953
rect 3976 5608 3984 5653
rect 4016 5596 4024 5813
rect 4216 5747 4224 5864
rect 4236 5787 4244 5833
rect 4256 5807 4264 5864
rect 4396 5860 4404 5864
rect 4056 5596 4064 5673
rect 4036 5560 4044 5564
rect 4033 5547 4047 5560
rect 4076 5507 4084 5564
rect 4116 5547 4124 5693
rect 3816 5267 3824 5493
rect 3876 5376 3884 5453
rect 4036 5376 4044 5433
rect 3856 5267 3864 5344
rect 3816 5087 3824 5193
rect 3856 5147 3864 5253
rect 4016 5227 4024 5332
rect 3827 5084 3840 5087
rect 3827 5076 3844 5084
rect 3827 5073 3840 5076
rect 3896 5007 3904 5044
rect 3636 4568 3644 4613
rect 3716 4556 3724 4813
rect 3736 4767 3744 4824
rect 3756 4568 3764 4793
rect 3476 4516 3504 4524
rect 3516 4520 3524 4524
rect 3376 4347 3384 4373
rect 3296 4227 3304 4304
rect 3356 4247 3364 4292
rect 3396 4267 3404 4493
rect 3416 4487 3424 4513
rect 3416 4307 3424 4433
rect 3476 4427 3484 4493
rect 3476 4336 3484 4413
rect 3496 4407 3504 4516
rect 3513 4507 3527 4520
rect 3636 4507 3644 4554
rect 3526 4500 3527 4507
rect 3536 4467 3544 4493
rect 3236 4044 3244 4113
rect 3236 4036 3264 4044
rect 3056 4000 3064 4004
rect 3053 3987 3067 4000
rect 3076 3996 3104 4004
rect 2927 3776 2944 3784
rect 2676 3487 2684 3573
rect 2713 3520 2727 3533
rect 2716 3516 2724 3520
rect 2816 3516 2824 3553
rect 2876 3516 2884 3573
rect 2476 3456 2493 3467
rect 2480 3453 2493 3456
rect 2596 3407 2604 3484
rect 2376 3316 2404 3324
rect 2396 3296 2404 3316
rect 2296 3260 2304 3264
rect 2293 3247 2307 3260
rect 2476 3264 2484 3373
rect 2256 2996 2264 3173
rect 2316 2967 2324 3133
rect 2336 3047 2344 3252
rect 2376 3107 2384 3253
rect 2416 3047 2424 3133
rect 2456 3127 2464 3213
rect 2476 3167 2484 3250
rect 2516 3227 2524 3264
rect 2616 3227 2624 3353
rect 2636 3107 2644 3473
rect 2656 3347 2664 3453
rect 2656 3207 2664 3333
rect 2736 3327 2744 3353
rect 2776 3347 2784 3484
rect 2796 3407 2804 3473
rect 2916 3464 2924 3772
rect 2956 3667 2964 3753
rect 2976 3727 2984 3784
rect 2976 3687 2984 3713
rect 3076 3647 3084 3996
rect 3356 4004 3364 4053
rect 3156 3816 3164 3973
rect 2936 3484 2944 3613
rect 3036 3567 3044 3633
rect 3096 3627 3104 3813
rect 3216 3787 3224 4004
rect 3336 3996 3364 4004
rect 3136 3747 3144 3784
rect 3116 3607 3124 3693
rect 2916 3456 2944 3464
rect 2696 3227 2704 3264
rect 2736 3227 2744 3264
rect 2696 3127 2704 3213
rect 2733 3207 2747 3213
rect 2776 3107 2784 3333
rect 2796 3187 2804 3393
rect 2896 3347 2904 3393
rect 2853 3300 2867 3313
rect 2856 3296 2864 3300
rect 2896 3296 2904 3333
rect 2936 3267 2944 3456
rect 2956 3227 2964 3333
rect 3016 3296 3024 3333
rect 3036 3327 3044 3532
rect 3056 3487 3064 3573
rect 3096 3516 3104 3553
rect 3136 3547 3144 3613
rect 3156 3527 3164 3753
rect 3136 3516 3153 3524
rect 3056 3296 3064 3353
rect 3156 3327 3164 3473
rect 3176 3447 3184 3553
rect 3196 3310 3204 3693
rect 3236 3627 3244 3953
rect 3313 3847 3327 3853
rect 3336 3847 3344 3996
rect 3376 3984 3384 4213
rect 3456 4047 3464 4292
rect 3476 4007 3484 4253
rect 3356 3976 3384 3984
rect 3293 3820 3307 3833
rect 3296 3816 3304 3820
rect 3276 3687 3284 3784
rect 3316 3764 3324 3772
rect 3316 3756 3344 3764
rect 3216 3528 3224 3593
rect 3296 3548 3304 3573
rect 3316 3527 3324 3613
rect 3336 3527 3344 3756
rect 3356 3727 3364 3976
rect 3396 3847 3404 3873
rect 3396 3747 3404 3784
rect 3436 3780 3444 3784
rect 3433 3767 3447 3780
rect 2196 2807 2204 2953
rect 2276 2960 2284 2964
rect 2273 2947 2287 2960
rect 2176 2776 2204 2784
rect 1956 2627 1964 2744
rect 1996 2687 2004 2744
rect 1856 2476 1864 2513
rect 1896 2476 1944 2484
rect 1993 2480 2007 2493
rect 1996 2476 2004 2480
rect 1816 2447 1824 2474
rect 1936 2387 1944 2476
rect 2016 2440 2024 2444
rect 2013 2427 2027 2440
rect 2056 2347 2064 2774
rect 2196 2727 2204 2776
rect 2207 2716 2224 2724
rect 1856 2256 1864 2313
rect 2116 2264 2124 2553
rect 2176 2407 2184 2444
rect 2216 2427 2224 2716
rect 2236 2507 2244 2793
rect 2256 2747 2264 2913
rect 2336 2827 2344 3033
rect 2416 2996 2424 3033
rect 2436 2956 2464 2964
rect 2336 2740 2344 2744
rect 2333 2727 2347 2740
rect 2396 2667 2404 2893
rect 2436 2827 2444 2933
rect 2456 2927 2464 2956
rect 2476 2947 2484 3093
rect 2496 2887 2504 2953
rect 2436 2776 2444 2813
rect 2536 2807 2544 2931
rect 2576 2867 2584 2964
rect 2676 2884 2684 3013
rect 2656 2876 2684 2884
rect 2576 2827 2584 2853
rect 2536 2747 2544 2793
rect 2613 2780 2627 2793
rect 2616 2776 2624 2780
rect 2656 2776 2664 2876
rect 2456 2740 2464 2744
rect 2453 2727 2467 2740
rect 2496 2687 2504 2744
rect 2556 2707 2564 2773
rect 2427 2676 2453 2684
rect 2276 2476 2284 2553
rect 2313 2480 2327 2493
rect 2316 2476 2324 2480
rect 2376 2440 2384 2444
rect 2256 2327 2264 2432
rect 2373 2427 2387 2440
rect 2116 2256 2144 2264
rect 1836 2167 1844 2224
rect 1776 1956 1784 1993
rect 1876 1970 1884 2210
rect 1956 2007 1964 2033
rect 1876 1847 1884 1956
rect 1896 1867 1904 1993
rect 1956 1956 1964 1993
rect 1976 1987 1984 2224
rect 2036 2226 2044 2253
rect 1996 2007 2004 2213
rect 2000 1964 2013 1967
rect 1996 1956 2013 1964
rect 2000 1953 2013 1956
rect 1936 1920 1944 1924
rect 1933 1907 1947 1920
rect 1716 1736 1724 1773
rect 1696 1667 1704 1704
rect 1816 1627 1824 1813
rect 1536 1404 1544 1433
rect 1396 1400 1404 1404
rect 1393 1387 1407 1400
rect 1436 1307 1444 1404
rect 1416 1216 1424 1253
rect 1396 1180 1404 1184
rect 1393 1167 1407 1180
rect 1436 1127 1444 1172
rect 1456 916 1464 953
rect 956 696 964 733
rect 416 276 464 284
rect 396 176 404 273
rect 536 176 544 293
rect 656 190 664 353
rect 776 184 784 533
rect 996 467 1004 664
rect 1076 527 1084 913
rect 1236 887 1244 914
rect 1156 807 1164 873
rect 1176 847 1184 884
rect 1156 696 1164 793
rect 1296 696 1304 872
rect 1136 660 1144 664
rect 1133 647 1147 660
rect 1016 424 1024 513
rect 1036 427 1044 453
rect 996 416 1024 424
rect 776 176 804 184
rect 796 144 804 176
rect 836 167 844 364
rect 916 360 924 364
rect 913 347 927 360
rect 876 176 884 313
rect 96 -24 104 13
rect 356 -24 364 144
rect 496 -24 504 144
rect 756 136 804 144
rect 956 -16 964 273
rect 976 247 984 394
rect 996 327 1004 416
rect 1027 404 1040 407
rect 1116 404 1124 533
rect 1156 447 1164 553
rect 1027 396 1044 404
rect 1096 396 1124 404
rect 1027 393 1040 396
rect 1156 366 1164 433
rect 996 188 1004 313
rect 1016 204 1024 353
rect 1053 344 1067 353
rect 1036 340 1067 344
rect 1036 336 1064 340
rect 1036 287 1044 336
rect 1196 207 1204 364
rect 1316 287 1324 613
rect 1436 507 1444 573
rect 1536 547 1544 873
rect 1556 847 1564 1493
rect 1616 1444 1624 1473
rect 1676 1444 1684 1513
rect 1596 1436 1624 1444
rect 1656 1436 1704 1444
rect 1696 1184 1704 1436
rect 1676 916 1684 993
rect 1616 880 1624 884
rect 1596 807 1604 873
rect 1613 867 1627 880
rect 1556 667 1564 694
rect 1696 666 1704 853
rect 1596 627 1604 664
rect 1656 656 1684 664
rect 1676 547 1684 656
rect 1016 196 1044 204
rect 1036 176 1044 196
rect 1167 204 1180 207
rect 1167 193 1184 204
rect 1096 144 1104 193
rect 1176 176 1184 193
rect 1253 190 1267 193
rect 1356 184 1364 364
rect 1336 176 1364 184
rect 1456 184 1464 533
rect 1536 447 1544 473
rect 1496 307 1504 352
rect 1456 176 1484 184
rect 1116 146 1124 173
rect 1056 136 1104 144
rect 1336 144 1344 176
rect 1476 144 1484 176
rect 1516 47 1524 333
rect 1536 287 1544 364
rect 1596 356 1624 364
rect 1576 176 1584 353
rect 1596 287 1604 356
rect 1676 307 1684 393
rect 1636 147 1644 273
rect 1696 247 1704 453
rect 1716 407 1724 1593
rect 1796 1448 1804 1573
rect 1836 1527 1844 1833
rect 1976 1704 1984 1773
rect 2016 1748 2024 1893
rect 2036 1787 2044 2093
rect 2136 2007 2144 2256
rect 2336 2147 2344 2212
rect 2056 1748 2064 1954
rect 2076 1927 2084 1953
rect 2016 1704 2024 1734
rect 2136 1706 2144 1773
rect 2216 1748 2224 1993
rect 2276 1956 2284 2013
rect 2296 1867 2304 1924
rect 2416 1907 2424 2353
rect 2436 2287 2444 2653
rect 2456 2267 2464 2613
rect 2556 2476 2564 2513
rect 2576 2487 2584 2733
rect 2596 2627 2604 2732
rect 2596 2436 2624 2444
rect 2476 2367 2484 2433
rect 2596 2387 2604 2436
rect 2476 2067 2484 2224
rect 2536 2067 2544 2313
rect 2556 2226 2564 2333
rect 2596 2256 2604 2373
rect 2536 1987 2544 2053
rect 2536 1964 2544 1973
rect 2516 1956 2544 1964
rect 2336 1736 2344 1773
rect 1936 1696 1964 1704
rect 1956 1527 1964 1696
rect 2016 1696 2044 1704
rect 1736 1186 1744 1253
rect 1836 1228 1844 1433
rect 1856 1347 1864 1473
rect 2036 1448 2044 1696
rect 2113 1440 2127 1453
rect 2116 1436 2124 1440
rect 1876 1407 1884 1434
rect 2016 1407 2024 1434
rect 1796 1107 1804 1153
rect 1736 886 1744 953
rect 1796 928 1804 1093
rect 1816 1087 1824 1184
rect 1876 1167 1884 1372
rect 1936 1347 1944 1404
rect 1896 1167 1904 1213
rect 1956 1180 1964 1184
rect 1996 1180 2004 1184
rect 1953 1167 1967 1180
rect 1993 1167 2007 1180
rect 1833 1147 1847 1153
rect 2036 1147 2044 1434
rect 2176 1406 2184 1733
rect 2236 1467 2244 1704
rect 2376 1587 2384 1704
rect 2496 1667 2504 1704
rect 2536 1607 2544 1893
rect 2136 1307 2144 1404
rect 2056 1167 2064 1273
rect 2096 1216 2104 1293
rect 2196 1247 2204 1453
rect 2336 1307 2344 1433
rect 2436 1406 2444 1433
rect 2456 1407 2464 1593
rect 2556 1587 2564 2212
rect 2676 2147 2684 2553
rect 2696 2347 2704 3092
rect 2816 3047 2824 3153
rect 2733 3000 2747 3013
rect 2816 3004 2824 3033
rect 2736 2996 2744 3000
rect 2796 2996 2824 3004
rect 2716 2746 2724 2953
rect 2836 2867 2844 3213
rect 2836 2776 2844 2832
rect 2856 2787 2864 3133
rect 2876 2907 2884 3213
rect 3036 3104 3044 3252
rect 3096 3244 3104 3264
rect 3076 3236 3104 3244
rect 3036 3096 3064 3104
rect 2916 2996 2924 3093
rect 2956 2956 2984 2964
rect 2936 2827 2944 2950
rect 2956 2787 2964 2833
rect 2976 2807 2984 2956
rect 3056 2867 3064 3096
rect 3076 3047 3084 3236
rect 3156 3227 3164 3264
rect 3216 3047 3224 3413
rect 3276 3387 3284 3484
rect 3296 3127 3304 3173
rect 3316 3087 3324 3473
rect 3336 3427 3344 3513
rect 3336 3227 3344 3373
rect 3356 3307 3364 3673
rect 3376 3527 3384 3573
rect 3393 3520 3407 3533
rect 3396 3516 3404 3520
rect 3436 3516 3444 3753
rect 3476 3687 3484 3972
rect 3496 3687 3504 4292
rect 3536 4267 3544 4334
rect 3556 4307 3564 4473
rect 3633 4344 3647 4353
rect 3627 4340 3647 4344
rect 3627 4336 3644 4340
rect 3516 3987 3524 4193
rect 3536 3967 3544 4232
rect 3596 4207 3604 4292
rect 3656 4287 3664 4353
rect 3676 4307 3684 4493
rect 3696 4467 3704 4512
rect 3756 4507 3764 4554
rect 3573 4040 3587 4053
rect 3576 4036 3584 4040
rect 3616 4036 3624 4273
rect 3676 4167 3684 4293
rect 3696 4147 3704 4393
rect 3716 4367 3724 4493
rect 3776 4407 3784 4753
rect 3796 4567 3804 4813
rect 3816 4807 3824 4973
rect 3816 4667 3824 4753
rect 3836 4627 3844 4973
rect 3856 4827 3864 4953
rect 3936 4947 3944 5153
rect 3973 5080 3987 5093
rect 4036 5087 4044 5273
rect 4096 5207 4104 5374
rect 4116 5307 4124 5453
rect 4136 5287 4144 5713
rect 4233 5600 4247 5613
rect 4236 5596 4244 5600
rect 4167 5564 4180 5567
rect 4167 5553 4184 5564
rect 4176 5507 4184 5553
rect 4156 5287 4164 5393
rect 4196 5376 4204 5513
rect 4216 5407 4224 5564
rect 4276 5387 4284 5613
rect 4296 5347 4304 5374
rect 4213 5327 4227 5332
rect 4256 5307 4264 5344
rect 4020 5084 4033 5087
rect 3976 5076 3984 5080
rect 4016 5076 4033 5084
rect 4020 5073 4033 5076
rect 3916 4856 3924 4893
rect 3976 4867 3984 4893
rect 3896 4707 3904 4824
rect 3936 4816 3964 4824
rect 3936 4727 3944 4816
rect 3996 4727 4004 4993
rect 4036 4967 4044 5033
rect 4056 4987 4064 5133
rect 4076 5007 4084 5093
rect 4036 4856 4044 4913
rect 4076 4856 4084 4913
rect 4136 4824 4144 5044
rect 4176 5007 4184 5044
rect 4116 4816 4144 4824
rect 3896 4567 3904 4613
rect 3733 4340 3747 4353
rect 3736 4336 3744 4340
rect 3756 4204 3764 4292
rect 3756 4196 3784 4204
rect 3656 4044 3664 4113
rect 3656 4036 3673 4044
rect 3736 4036 3744 4073
rect 3776 4027 3784 4196
rect 3796 4107 3804 4513
rect 3816 4427 3824 4524
rect 3856 4487 3864 4524
rect 3816 4306 3824 4353
rect 3836 4347 3844 4373
rect 3876 4336 3884 4493
rect 3896 4487 3904 4513
rect 3916 4507 3924 4673
rect 3936 4447 3944 4713
rect 4016 4707 4024 4812
rect 4056 4627 4064 4753
rect 3973 4584 3987 4593
rect 3973 4580 4004 4584
rect 3976 4576 4004 4580
rect 3996 4556 4004 4576
rect 3947 4436 3964 4444
rect 3836 4207 3844 4293
rect 3896 4247 3904 4304
rect 3556 3907 3564 3993
rect 3636 3927 3644 4004
rect 3616 3816 3624 3853
rect 3736 3827 3744 3973
rect 3516 3786 3524 3813
rect 3596 3747 3604 3784
rect 3656 3747 3664 3784
rect 3707 3784 3720 3787
rect 3707 3776 3724 3784
rect 3707 3773 3720 3776
rect 3736 3747 3744 3773
rect 3556 3607 3564 3713
rect 3473 3567 3487 3573
rect 3473 3560 3493 3567
rect 3476 3556 3493 3560
rect 3480 3553 3493 3556
rect 3453 3544 3467 3553
rect 3453 3540 3484 3544
rect 3456 3536 3484 3540
rect 3476 3524 3484 3536
rect 3476 3516 3493 3524
rect 3556 3516 3564 3553
rect 3596 3507 3604 3712
rect 3376 3296 3384 3413
rect 3416 3296 3424 3373
rect 3356 3167 3364 3253
rect 3436 3227 3444 3264
rect 3176 2996 3184 3033
rect 3316 2996 3324 3033
rect 3216 2847 3224 2993
rect 2736 2667 2744 2773
rect 2776 2707 2784 2744
rect 2876 2740 2884 2744
rect 2873 2727 2887 2740
rect 2836 2547 2844 2713
rect 2936 2667 2944 2744
rect 2976 2647 2984 2793
rect 2956 2636 2973 2644
rect 2736 2256 2744 2413
rect 2816 2327 2824 2433
rect 2956 2264 2964 2636
rect 2996 2624 3004 2773
rect 3096 2687 3104 2776
rect 3136 2747 3144 2833
rect 3213 2780 3227 2793
rect 3236 2787 3244 2893
rect 3216 2776 3224 2780
rect 2936 2256 2964 2264
rect 2976 2616 3004 2624
rect 2696 2127 2704 2254
rect 2796 2127 2804 2224
rect 2836 2167 2844 2254
rect 2896 2127 2904 2224
rect 2976 2167 2984 2616
rect 3256 2547 3264 2913
rect 3276 2807 3284 2964
rect 3356 2827 3364 3053
rect 3353 2787 3367 2792
rect 3336 2740 3344 2744
rect 3333 2727 3347 2740
rect 3076 2407 3084 2476
rect 3296 2476 3304 2533
rect 3376 2487 3384 3073
rect 3436 2960 3444 2964
rect 3433 2947 3447 2960
rect 3416 2936 3433 2944
rect 3396 2746 3404 2853
rect 3120 2444 3140 2447
rect 3127 2433 3144 2444
rect 3013 2260 3027 2273
rect 3016 2256 3024 2260
rect 2656 1956 2664 2013
rect 2696 1968 2704 2113
rect 2916 1987 2924 2133
rect 2576 1867 2584 1953
rect 2676 1607 2684 1924
rect 2776 1787 2784 1924
rect 2856 1827 2864 1973
rect 2916 1956 2924 1973
rect 2956 1956 2964 2013
rect 2796 1767 2804 1793
rect 2856 1764 2864 1813
rect 2836 1756 2864 1764
rect 2936 1764 2944 1924
rect 2936 1756 2964 1764
rect 2516 1347 2524 1404
rect 2396 1316 2444 1324
rect 2396 1287 2404 1316
rect 2176 1207 2184 1214
rect 2176 1147 2184 1193
rect 2356 1186 2364 1233
rect 2387 1213 2393 1227
rect 2416 1216 2424 1293
rect 2436 1287 2444 1316
rect 2516 1186 2524 1333
rect 1836 947 1844 1033
rect 1833 920 1847 933
rect 1836 916 1844 920
rect 1876 807 1884 933
rect 1976 916 1984 953
rect 1896 847 1904 913
rect 1916 787 1924 853
rect 1996 847 2004 884
rect 2016 876 2044 884
rect 2016 807 2024 876
rect 2096 807 2104 1013
rect 1816 660 1824 664
rect 1813 647 1827 660
rect 1836 624 1844 653
rect 1856 647 1864 753
rect 1956 696 2004 704
rect 2056 666 2064 793
rect 2116 787 2124 1133
rect 2536 1087 2544 1393
rect 2596 1387 2604 1573
rect 2287 1073 2293 1087
rect 2556 1067 2564 1373
rect 2596 1147 2604 1184
rect 2656 1147 2664 1214
rect 2456 1007 2464 1053
rect 2276 887 2284 973
rect 2216 707 2224 733
rect 2236 667 2244 873
rect 2276 696 2284 793
rect 2296 787 2304 913
rect 2376 847 2384 884
rect 2296 727 2304 773
rect 2316 696 2324 733
rect 2176 656 2193 664
rect 1807 616 1844 624
rect 1736 396 1744 593
rect 1816 404 1824 533
rect 1796 396 1824 404
rect 1896 360 1904 364
rect 1893 347 1907 360
rect 1556 47 1564 144
rect 1776 146 1784 253
rect 1836 207 1844 333
rect 1896 267 1904 312
rect 1856 176 1864 213
rect 1896 176 1904 253
rect 1916 187 1924 253
rect 1996 207 2004 533
rect 2076 396 2084 433
rect 2056 360 2064 364
rect 2053 347 2067 360
rect 2116 347 2124 613
rect 2196 547 2204 653
rect 2336 396 2344 664
rect 2396 567 2404 694
rect 2416 627 2424 953
rect 2616 916 2624 1053
rect 2473 708 2487 713
rect 2536 704 2544 914
rect 2676 847 2684 1233
rect 2736 1216 2744 1273
rect 2756 1247 2764 1453
rect 2776 1444 2784 1734
rect 2796 1468 2804 1753
rect 2836 1736 2844 1756
rect 2936 1667 2944 1734
rect 2956 1706 2964 1756
rect 2976 1747 2984 1893
rect 2996 1767 3004 2213
rect 3056 2147 3064 2224
rect 3096 2007 3104 2333
rect 3116 2227 3124 2273
rect 3136 2027 3144 2433
rect 3176 2347 3184 2432
rect 3356 2407 3364 2444
rect 3196 2284 3204 2353
rect 3273 2287 3287 2293
rect 3176 2276 3204 2284
rect 3176 2256 3184 2276
rect 3213 2260 3227 2273
rect 3216 2256 3224 2260
rect 3316 2256 3324 2313
rect 3376 2264 3384 2433
rect 3396 2327 3404 2653
rect 3416 2607 3424 2936
rect 3476 2907 3484 3353
rect 3496 3347 3504 3373
rect 3496 3127 3504 3312
rect 3556 3308 3564 3373
rect 3536 3260 3544 3264
rect 3476 2776 3484 2833
rect 3496 2827 3504 3113
rect 3516 2788 3524 3253
rect 3533 3247 3547 3260
rect 3536 3067 3544 3233
rect 3596 3087 3604 3472
rect 3616 3227 3624 3673
rect 3756 3524 3764 3893
rect 3776 3747 3784 4013
rect 3796 3927 3804 4033
rect 3896 4004 3904 4153
rect 3876 3996 3904 4004
rect 3876 3787 3884 3996
rect 3896 3887 3904 3973
rect 3916 3844 3924 4113
rect 3936 4004 3944 4233
rect 3956 4044 3964 4436
rect 3976 4267 3984 4524
rect 4036 4387 4044 4493
rect 4076 4347 4084 4713
rect 4047 4344 4060 4347
rect 4047 4336 4064 4344
rect 4047 4333 4060 4336
rect 3996 4127 4004 4293
rect 4016 4267 4024 4304
rect 4036 4087 4044 4293
rect 3973 4067 3987 4073
rect 3956 4036 3984 4044
rect 3936 3996 3964 4004
rect 3936 3947 3944 3996
rect 3956 3927 3964 3996
rect 3907 3836 3924 3844
rect 3896 3786 3904 3833
rect 4036 3824 4044 3993
rect 4056 3847 4064 4173
rect 4076 4084 4084 4293
rect 4096 4167 4104 4693
rect 4116 4527 4124 4816
rect 4156 4727 4164 4933
rect 4216 4927 4224 5074
rect 4236 4868 4244 5173
rect 4256 4947 4264 5272
rect 4296 5076 4304 5312
rect 4316 5187 4324 5673
rect 4336 5604 4344 5852
rect 4393 5847 4407 5860
rect 4556 5827 4564 5852
rect 4596 5807 4604 5953
rect 4336 5596 4364 5604
rect 4396 5596 4404 5733
rect 4576 5627 4584 5733
rect 4616 5687 4624 5933
rect 4636 5687 4644 5973
rect 4707 5914 4713 5927
rect 4707 5913 4720 5914
rect 4696 5860 4704 5864
rect 4693 5847 4707 5860
rect 4436 5587 4444 5613
rect 4456 5567 4464 5613
rect 4493 5600 4507 5613
rect 4496 5596 4504 5600
rect 4576 5567 4584 5613
rect 4613 5600 4627 5613
rect 4616 5596 4624 5600
rect 4596 5467 4604 5513
rect 4636 5507 4644 5564
rect 4356 5388 4364 5413
rect 4336 5284 4344 5333
rect 4416 5340 4424 5344
rect 4373 5327 4387 5332
rect 4413 5327 4427 5340
rect 4336 5276 4364 5284
rect 4336 5087 4344 5253
rect 4276 4967 4284 5033
rect 4356 4887 4364 5276
rect 4416 5267 4424 5313
rect 4456 5307 4464 5373
rect 4596 5346 4604 5373
rect 4496 5340 4504 5344
rect 4536 5340 4544 5344
rect 4493 5327 4507 5340
rect 4476 5316 4493 5324
rect 4456 5087 4464 5213
rect 4376 5007 4384 5073
rect 4396 4884 4404 5033
rect 4436 4967 4444 5044
rect 4376 4876 4404 4884
rect 4276 4787 4284 4824
rect 4156 4568 4164 4692
rect 4216 4627 4224 4713
rect 4216 4556 4224 4613
rect 4176 4520 4184 4524
rect 4173 4507 4187 4520
rect 4116 4327 4124 4353
rect 4156 4336 4164 4413
rect 4193 4340 4207 4353
rect 4236 4347 4244 4513
rect 4256 4507 4264 4773
rect 4276 4567 4284 4633
rect 4316 4607 4324 4873
rect 4376 4856 4384 4876
rect 4356 4664 4364 4773
rect 4376 4684 4384 4713
rect 4396 4707 4404 4824
rect 4413 4684 4427 4693
rect 4376 4680 4427 4684
rect 4376 4676 4424 4680
rect 4356 4656 4384 4664
rect 4320 4584 4333 4587
rect 4316 4573 4333 4584
rect 4316 4556 4324 4573
rect 4356 4567 4364 4593
rect 4336 4487 4344 4524
rect 4196 4336 4204 4340
rect 4256 4327 4264 4353
rect 4216 4300 4224 4304
rect 4213 4287 4227 4300
rect 4216 4187 4224 4273
rect 4256 4267 4264 4313
rect 4276 4207 4284 4453
rect 4336 4336 4344 4473
rect 4356 4407 4364 4513
rect 4376 4347 4384 4656
rect 4293 4287 4307 4293
rect 4316 4267 4324 4304
rect 4316 4167 4324 4253
rect 4076 4076 4104 4084
rect 4076 4007 4084 4053
rect 4096 4047 4104 4076
rect 4113 4040 4127 4053
rect 4116 4036 4124 4040
rect 4156 4036 4164 4113
rect 4193 4048 4207 4053
rect 4016 3816 4044 3824
rect 3856 3607 3864 3753
rect 3856 3544 3864 3593
rect 3856 3536 3884 3544
rect 3747 3516 3764 3524
rect 3840 3524 3853 3527
rect 3836 3516 3853 3524
rect 3840 3513 3853 3516
rect 3656 3296 3664 3333
rect 3716 3307 3724 3470
rect 3696 3167 3704 3264
rect 3616 3004 3624 3053
rect 3636 3027 3644 3153
rect 3596 2996 3624 3004
rect 3576 2787 3584 2964
rect 3636 2947 3644 3013
rect 3596 2788 3604 2893
rect 3636 2776 3644 2833
rect 3676 2807 3684 3093
rect 3716 3067 3724 3133
rect 3736 3107 3744 3513
rect 3756 3247 3764 3413
rect 3776 3387 3784 3484
rect 3876 3427 3884 3536
rect 3776 3067 3784 3333
rect 3896 3324 3904 3772
rect 3916 3607 3924 3773
rect 3916 3347 3924 3593
rect 4016 3567 4024 3816
rect 4056 3764 4064 3784
rect 4056 3756 4084 3764
rect 3947 3524 3960 3527
rect 3947 3516 3964 3524
rect 4013 3520 4027 3532
rect 4016 3516 4024 3520
rect 3947 3513 3960 3516
rect 3936 3387 3944 3473
rect 3976 3407 3984 3484
rect 3940 3366 3960 3367
rect 3947 3363 3960 3366
rect 3947 3360 3964 3363
rect 3947 3353 3967 3360
rect 3953 3347 3967 3353
rect 3896 3316 3924 3324
rect 3873 3307 3887 3313
rect 3816 3227 3824 3264
rect 3856 3260 3864 3264
rect 3853 3247 3867 3260
rect 3896 3227 3904 3273
rect 3916 3247 3924 3316
rect 3976 3296 3984 3353
rect 4036 3307 4044 3353
rect 3947 3264 3960 3267
rect 3947 3256 3964 3264
rect 3947 3253 3960 3256
rect 3967 3244 3980 3247
rect 3967 3233 3984 3244
rect 3816 3127 3824 3213
rect 3716 2960 3724 2964
rect 3713 2947 3727 2960
rect 3796 2947 3804 3073
rect 3856 2996 3864 3053
rect 3447 2744 3460 2747
rect 3447 2736 3464 2744
rect 3447 2733 3460 2736
rect 3556 2724 3564 2773
rect 3536 2716 3564 2724
rect 3376 2256 3404 2264
rect 3396 2226 3404 2256
rect 3196 2220 3204 2224
rect 3296 2220 3304 2224
rect 3193 2207 3207 2220
rect 3293 2207 3307 2220
rect 3100 1984 3113 1987
rect 3096 1973 3113 1984
rect 2996 1736 3004 1753
rect 3016 1747 3024 1973
rect 3096 1956 3104 1973
rect 3036 1787 3044 1953
rect 3076 1920 3084 1924
rect 3116 1920 3124 1924
rect 3073 1907 3087 1920
rect 3113 1907 3127 1920
rect 3073 1887 3087 1893
rect 3156 1887 3164 1993
rect 3196 1968 3204 2153
rect 3233 1960 3247 1973
rect 3313 1960 3327 1973
rect 3236 1956 3244 1960
rect 3316 1956 3324 1960
rect 3176 1747 3184 1913
rect 3216 1887 3224 1924
rect 3416 1887 3424 2533
rect 3536 2507 3544 2716
rect 3576 2707 3584 2733
rect 3656 2707 3664 2744
rect 3556 2696 3573 2704
rect 3436 2387 3444 2473
rect 3456 2327 3464 2493
rect 3556 2476 3564 2696
rect 3456 2307 3464 2313
rect 3447 2296 3464 2307
rect 3447 2293 3460 2296
rect 3436 2280 3504 2284
rect 3433 2276 3504 2280
rect 3433 2267 3447 2276
rect 3496 2256 3504 2276
rect 3556 2267 3564 2413
rect 3596 2367 3604 2553
rect 3616 2427 3624 2493
rect 3676 2476 3684 2593
rect 3696 2507 3704 2773
rect 3716 2746 3724 2793
rect 3756 2776 3764 2933
rect 3836 2867 3844 2964
rect 3896 2907 3904 3113
rect 3916 3027 3924 3212
rect 3936 3127 3944 3213
rect 3936 3008 3944 3113
rect 3976 3028 3984 3233
rect 3996 3227 4004 3264
rect 3996 3004 4004 3093
rect 3987 2996 4004 3004
rect 3816 2787 3824 2833
rect 3836 2788 3844 2853
rect 3956 2807 3964 2964
rect 3776 2507 3784 2744
rect 3836 2567 3844 2774
rect 3976 2776 3984 2933
rect 3856 2667 3864 2773
rect 3713 2480 3727 2493
rect 3756 2496 3773 2504
rect 3716 2476 3724 2480
rect 3656 2440 3664 2444
rect 3653 2427 3667 2440
rect 3596 2264 3604 2353
rect 3576 2256 3604 2264
rect 3616 2256 3624 2313
rect 3476 2220 3484 2224
rect 3516 2220 3524 2224
rect 2973 1687 2987 1693
rect 2896 1567 2904 1613
rect 2776 1436 2793 1444
rect 2893 1440 2907 1453
rect 2896 1436 2904 1440
rect 2956 1436 2964 1493
rect 2976 1444 2984 1593
rect 2996 1467 3004 1653
rect 2976 1436 3004 1444
rect 2996 1404 3004 1436
rect 2816 1347 2824 1404
rect 2976 1396 3004 1404
rect 2776 1216 2784 1333
rect 2716 1067 2724 1184
rect 2716 787 2724 913
rect 2527 696 2544 704
rect 2436 487 2444 694
rect 2616 647 2624 733
rect 2636 667 2644 693
rect 2776 664 2784 773
rect 2676 660 2684 664
rect 2673 647 2687 660
rect 1796 127 1804 173
rect 2036 147 2044 213
rect 2216 188 2224 364
rect 2276 347 2284 373
rect 2276 227 2284 253
rect 1836 140 1844 144
rect 1833 127 1847 140
rect 2276 144 2284 213
rect 2316 188 2324 352
rect 2353 347 2367 352
rect 2396 227 2404 393
rect 2416 367 2424 433
rect 2536 247 2544 364
rect 2576 347 2584 393
rect 2596 267 2604 413
rect 2627 404 2640 407
rect 2627 396 2644 404
rect 2627 393 2640 396
rect 2656 287 2664 352
rect 2696 347 2704 553
rect 2776 427 2784 650
rect 2796 647 2804 1073
rect 2816 727 2824 1273
rect 2836 1186 2844 1233
rect 2873 1220 2887 1233
rect 2876 1216 2884 1220
rect 2896 1147 2904 1184
rect 2876 916 2884 1093
rect 2956 1067 2964 1253
rect 2916 916 2924 973
rect 2956 827 2964 933
rect 2856 696 2864 733
rect 2893 700 2907 713
rect 2896 696 2904 700
rect 2816 666 2824 692
rect 2916 647 2924 664
rect 2476 146 2484 233
rect 2236 136 2284 144
rect 2636 144 2644 253
rect 2656 146 2664 233
rect 2696 176 2704 312
rect 2736 247 2744 364
rect 2776 360 2784 364
rect 2773 347 2787 360
rect 2836 327 2844 394
rect 2796 146 2804 213
rect 2836 187 2844 313
rect 2856 267 2864 453
rect 2916 408 2924 633
rect 2956 587 2964 694
rect 2956 467 2964 573
rect 2976 567 2984 1396
rect 3016 1287 3024 1693
rect 3036 1547 3044 1704
rect 3096 1667 3104 1690
rect 3156 1667 3164 1704
rect 3176 1607 3184 1693
rect 3196 1667 3204 1793
rect 3016 1216 3024 1252
rect 3096 1187 3104 1353
rect 3116 1167 3124 1593
rect 3136 1287 3144 1533
rect 3216 1487 3224 1813
rect 3273 1740 3287 1753
rect 3276 1736 3284 1740
rect 3316 1647 3324 1753
rect 3376 1748 3384 1873
rect 3436 1867 3444 2213
rect 3473 2207 3487 2220
rect 3513 2207 3527 2220
rect 3556 2187 3564 2232
rect 3576 2226 3584 2256
rect 3696 2267 3704 2444
rect 3716 2227 3724 2353
rect 3756 2284 3764 2496
rect 3876 2476 3884 2773
rect 3916 2587 3924 2744
rect 3956 2740 3964 2744
rect 3953 2727 3967 2740
rect 3736 2276 3764 2284
rect 3627 2196 3653 2204
rect 3580 2186 3593 2187
rect 3587 2173 3593 2186
rect 3676 1956 3684 1993
rect 3496 1920 3504 1924
rect 3493 1907 3507 1920
rect 3507 1896 3524 1904
rect 3416 1736 3424 1793
rect 3336 1587 3344 1734
rect 3516 1744 3524 1896
rect 3636 1867 3644 1924
rect 3696 1787 3704 1913
rect 3716 1807 3724 2192
rect 3736 1926 3744 2276
rect 3776 2264 3784 2472
rect 3756 2256 3784 2264
rect 3816 2256 3824 2333
rect 3856 2267 3864 2444
rect 3756 2207 3764 2256
rect 3796 2167 3804 2212
rect 3836 2187 3844 2224
rect 3896 2087 3904 2393
rect 3916 2107 3924 2313
rect 3936 2239 3944 2533
rect 3996 2488 4004 2733
rect 4016 2507 4024 2993
rect 4036 2787 4044 3253
rect 4056 3047 4064 3713
rect 4076 3687 4084 3756
rect 4116 3727 4124 3953
rect 4136 3947 4144 4004
rect 4176 3967 4184 3992
rect 4193 3987 4207 3993
rect 4216 3947 4224 4113
rect 4236 4067 4244 4133
rect 4256 4044 4264 4073
rect 4276 4048 4284 4073
rect 4356 4067 4364 4193
rect 4376 4087 4384 4293
rect 4396 4267 4404 4676
rect 4436 4664 4444 4854
rect 4456 4787 4464 4913
rect 4476 4887 4484 5316
rect 4533 5327 4547 5340
rect 4516 5076 4524 5133
rect 4556 5088 4564 5113
rect 4493 5024 4507 5033
rect 4493 5020 4524 5024
rect 4496 5016 4524 5020
rect 4516 4856 4524 5016
rect 4536 5007 4544 5044
rect 4576 4987 4584 5044
rect 4596 4967 4604 5013
rect 4616 4927 4624 5433
rect 4656 5376 4664 5473
rect 4676 5447 4684 5553
rect 4696 5467 4704 5833
rect 4716 5727 4724 5833
rect 4776 5747 4784 5993
rect 4796 5847 4804 5973
rect 4836 5947 4844 6044
rect 4876 5987 4884 6044
rect 4827 5924 4840 5927
rect 4827 5913 4844 5924
rect 4836 5896 4844 5913
rect 5196 5896 5204 5953
rect 4896 5860 4904 5864
rect 4856 5787 4864 5852
rect 4893 5847 4907 5860
rect 4873 5827 4887 5833
rect 4886 5820 4887 5827
rect 4716 5567 4724 5673
rect 4716 5447 4724 5532
rect 4736 5527 4744 5733
rect 4856 5724 4864 5773
rect 4856 5716 4884 5724
rect 4776 5596 4784 5693
rect 4836 5608 4844 5633
rect 4876 5564 4884 5716
rect 4916 5704 4924 5853
rect 4936 5827 4944 5893
rect 5056 5860 5064 5864
rect 4907 5696 4924 5704
rect 4896 5567 4904 5693
rect 4953 5600 4967 5613
rect 4956 5596 4964 5600
rect 5016 5607 5024 5852
rect 5053 5847 5067 5860
rect 5096 5807 5104 5894
rect 5173 5847 5187 5852
rect 5033 5608 5047 5613
rect 5156 5607 5164 5793
rect 4696 5376 4704 5413
rect 4636 5046 4644 5293
rect 4756 5167 4764 5453
rect 4776 5287 4784 5513
rect 4796 5447 4804 5564
rect 4856 5556 4884 5564
rect 4856 5376 4864 5556
rect 4976 5427 4984 5564
rect 4996 5467 5004 5513
rect 5016 5504 5024 5553
rect 5036 5527 5044 5594
rect 5176 5567 5184 5833
rect 5276 5827 5284 5894
rect 5376 5707 5384 5894
rect 5296 5596 5304 5693
rect 5336 5567 5344 5633
rect 5476 5608 5484 5933
rect 5496 5787 5504 5894
rect 5536 5827 5544 5864
rect 5636 5667 5644 5893
rect 5656 5864 5664 5913
rect 5693 5900 5707 5913
rect 5696 5896 5704 5900
rect 5916 5896 5924 5933
rect 5656 5856 5684 5864
rect 5576 5596 5584 5653
rect 5096 5544 5104 5552
rect 5076 5536 5104 5544
rect 5016 5496 5044 5504
rect 4996 5376 5004 5453
rect 5036 5376 5044 5496
rect 5076 5346 5084 5536
rect 5116 5427 5124 5533
rect 4836 5307 4844 5344
rect 4836 5247 4844 5293
rect 4876 5247 4884 5344
rect 5016 5307 5024 5344
rect 5116 5344 5124 5413
rect 5176 5376 5184 5532
rect 5416 5487 5424 5564
rect 5316 5376 5324 5453
rect 5456 5447 5464 5564
rect 5116 5336 5164 5344
rect 4773 5127 4787 5133
rect 4727 5113 4733 5127
rect 4753 5080 4767 5093
rect 4756 5076 4764 5080
rect 4656 5007 4664 5074
rect 4736 4947 4744 5032
rect 4796 5027 4804 5173
rect 4873 5088 4887 5093
rect 4996 5076 5004 5133
rect 5056 5087 5064 5273
rect 4856 5040 4864 5044
rect 4853 5027 4867 5040
rect 4896 5027 4904 5044
rect 4887 5016 4904 5027
rect 4887 5013 4900 5016
rect 4713 4860 4727 4873
rect 4716 4856 4724 4860
rect 4536 4787 4544 4824
rect 4576 4820 4584 4824
rect 4573 4807 4587 4820
rect 4587 4796 4604 4804
rect 4416 4656 4444 4664
rect 4416 4467 4424 4656
rect 4436 4526 4444 4593
rect 4453 4568 4467 4573
rect 4536 4556 4544 4773
rect 4576 4526 4584 4673
rect 4556 4427 4564 4513
rect 4453 4340 4467 4353
rect 4456 4336 4464 4340
rect 4516 4327 4524 4393
rect 4416 4064 4424 4273
rect 4436 4227 4444 4304
rect 4476 4300 4484 4304
rect 4473 4287 4487 4300
rect 4493 4287 4507 4293
rect 4376 4056 4424 4064
rect 4236 4036 4264 4044
rect 4236 4004 4244 4036
rect 4376 4044 4384 4056
rect 4356 4036 4384 4044
rect 4236 4000 4264 4004
rect 4236 3996 4267 4000
rect 4253 3987 4267 3996
rect 4233 3967 4247 3973
rect 4296 3967 4304 4004
rect 4136 3727 4144 3853
rect 4156 3667 4164 3814
rect 4316 3816 4324 3973
rect 4336 3827 4344 3993
rect 4356 3847 4364 4036
rect 4456 4036 4464 4133
rect 4387 4004 4400 4007
rect 4387 3993 4404 4004
rect 4436 4000 4444 4004
rect 4396 3904 4404 3993
rect 4433 3987 4447 4000
rect 4476 3967 4484 3993
rect 4396 3896 4424 3904
rect 4196 3607 4204 3784
rect 4236 3747 4244 3784
rect 4076 3367 4084 3553
rect 4176 3528 4184 3553
rect 4116 3447 4124 3484
rect 4156 3464 4164 3484
rect 4136 3456 4164 3464
rect 4136 3296 4144 3456
rect 4176 3307 4184 3393
rect 4076 3067 4084 3253
rect 4116 3227 4124 3264
rect 4156 3260 4164 3264
rect 4153 3247 4167 3260
rect 4176 3107 4184 3253
rect 4056 2947 4064 3012
rect 4196 3004 4204 3353
rect 4216 3187 4224 3673
rect 4276 3567 4284 3813
rect 4236 3307 4244 3373
rect 4276 3296 4284 3353
rect 4296 3327 4304 3473
rect 4316 3308 4324 3513
rect 4336 3427 4344 3773
rect 4356 3747 4364 3784
rect 4336 3266 4344 3353
rect 4260 3245 4280 3247
rect 4236 3207 4244 3233
rect 4267 3244 4280 3245
rect 4296 3244 4304 3264
rect 4356 3264 4364 3693
rect 4376 3527 4384 3773
rect 4396 3547 4404 3873
rect 4416 3544 4424 3896
rect 4436 3667 4444 3893
rect 4456 3827 4464 3933
rect 4476 3907 4484 3953
rect 4496 3887 4504 4252
rect 4516 3947 4524 4273
rect 4536 4247 4544 4353
rect 4576 4344 4584 4413
rect 4596 4367 4604 4796
rect 4616 4687 4624 4854
rect 4656 4787 4664 4824
rect 4693 4807 4707 4812
rect 4616 4567 4624 4633
rect 4616 4487 4624 4513
rect 4636 4464 4644 4524
rect 4676 4487 4684 4524
rect 4636 4456 4693 4464
rect 4616 4368 4624 4393
rect 4696 4367 4704 4432
rect 4693 4348 4707 4353
rect 4556 4336 4584 4344
rect 4536 4047 4544 4193
rect 4556 4067 4564 4336
rect 4716 4307 4724 4513
rect 4736 4407 4744 4653
rect 4756 4467 4764 5013
rect 4916 4967 4924 5013
rect 4936 4987 4944 5053
rect 4776 4647 4784 4933
rect 4956 4867 4964 5074
rect 4796 4556 4804 4633
rect 4816 4587 4824 4753
rect 4836 4627 4844 4673
rect 4876 4667 4884 4824
rect 4916 4687 4924 4813
rect 4916 4647 4924 4673
rect 4976 4627 4984 4824
rect 5016 4807 5024 4824
rect 5016 4664 5024 4793
rect 5016 4656 5044 4664
rect 4996 4568 5004 4593
rect 4776 4336 4784 4373
rect 4813 4340 4827 4353
rect 4853 4347 4867 4353
rect 4816 4336 4824 4340
rect 4596 4267 4604 4292
rect 4636 4247 4644 4304
rect 4596 4036 4604 4073
rect 4556 4000 4564 4004
rect 4553 3987 4567 4000
rect 4536 3907 4544 3953
rect 4467 3784 4480 3787
rect 4467 3776 4484 3784
rect 4467 3773 4480 3776
rect 4536 3727 4544 3784
rect 4416 3536 4444 3544
rect 4393 3520 4407 3533
rect 4436 3528 4444 3536
rect 4396 3516 4404 3520
rect 4416 3427 4424 3484
rect 4436 3367 4444 3453
rect 4476 3347 4484 3653
rect 4496 3527 4504 3713
rect 4536 3516 4544 3653
rect 4556 3547 4564 3773
rect 4576 3747 4584 3814
rect 4576 3607 4584 3733
rect 4596 3567 4604 3873
rect 4616 3827 4624 3993
rect 4636 3987 4644 4113
rect 4656 4006 4664 4093
rect 4676 4047 4684 4292
rect 4696 4127 4704 4253
rect 4716 4167 4724 4233
rect 4736 4048 4744 4293
rect 4756 4147 4764 4292
rect 4796 4067 4804 4133
rect 4816 4044 4824 4253
rect 4836 4147 4844 4304
rect 4856 4267 4864 4293
rect 4876 4224 4884 4453
rect 4896 4307 4904 4554
rect 4856 4220 4884 4224
rect 4853 4216 4884 4220
rect 4853 4207 4867 4216
rect 4916 4207 4924 4373
rect 4936 4364 4944 4512
rect 5036 4387 5044 4656
rect 5056 4527 5064 4993
rect 5076 4847 5084 5332
rect 5196 5287 5204 5344
rect 5276 5327 5284 5374
rect 5196 5247 5204 5273
rect 5096 5047 5104 5153
rect 5336 5088 5344 5332
rect 5376 5247 5384 5344
rect 5116 5027 5124 5074
rect 5136 4987 5144 5033
rect 5156 4864 5164 4933
rect 5176 4927 5184 5044
rect 5236 5027 5244 5073
rect 5156 4856 5184 4864
rect 5136 4787 5144 4824
rect 5176 4667 5184 4856
rect 5196 4807 5204 4973
rect 5376 4967 5384 5153
rect 5396 5044 5404 5313
rect 5416 5247 5424 5393
rect 5473 5380 5487 5393
rect 5476 5376 5484 5380
rect 5636 5376 5644 5564
rect 5676 5427 5684 5856
rect 5716 5844 5724 5864
rect 5696 5836 5724 5844
rect 5696 5507 5704 5836
rect 5756 5827 5764 5864
rect 5716 5424 5724 5813
rect 5816 5628 5824 5893
rect 5856 5627 5864 5864
rect 5773 5600 5787 5613
rect 5896 5607 5904 5864
rect 5776 5596 5784 5600
rect 5716 5416 5744 5424
rect 5456 5340 5464 5344
rect 5453 5327 5467 5340
rect 5656 5327 5664 5344
rect 5736 5344 5744 5416
rect 5796 5376 5804 5473
rect 5716 5336 5744 5344
rect 5527 5074 5533 5087
rect 5520 5073 5533 5074
rect 5556 5047 5564 5073
rect 5396 5036 5413 5044
rect 5416 5007 5424 5032
rect 5076 4484 5084 4653
rect 5176 4568 5184 4613
rect 5056 4476 5084 4484
rect 4936 4356 4964 4364
rect 4956 4336 4964 4356
rect 4987 4354 4993 4367
rect 4987 4353 5000 4354
rect 4976 4300 4984 4304
rect 4973 4287 4987 4300
rect 4796 4036 4824 4044
rect 4833 4040 4847 4053
rect 4876 4048 4884 4193
rect 4933 4184 4947 4193
rect 4916 4180 4947 4184
rect 4916 4176 4944 4180
rect 4836 4036 4844 4040
rect 4656 3887 4664 3992
rect 4676 3867 4684 3993
rect 4716 3967 4724 3993
rect 4716 3827 4724 3953
rect 4756 3816 4764 3893
rect 4796 3816 4804 4036
rect 4896 4047 4904 4093
rect 4893 3987 4907 3992
rect 4816 3887 4824 3933
rect 4836 3847 4844 3953
rect 4700 3786 4713 3787
rect 4676 3727 4684 3784
rect 4707 3773 4713 3786
rect 4776 3747 4784 3784
rect 4856 3744 4864 3913
rect 4896 3827 4904 3952
rect 4916 3907 4924 4176
rect 4956 4147 4964 4213
rect 4976 4187 4984 4252
rect 4996 4247 5004 4273
rect 4976 4087 4984 4152
rect 4996 4067 5004 4233
rect 5036 4227 5044 4253
rect 5056 4207 5064 4476
rect 5116 4467 5124 4524
rect 5156 4520 5164 4524
rect 5153 4507 5167 4520
rect 5216 4467 5224 4893
rect 5296 4856 5304 4893
rect 5416 4856 5424 4893
rect 5456 4856 5464 4993
rect 5496 4827 5504 4893
rect 5276 4767 5284 4824
rect 5316 4820 5324 4824
rect 5313 4807 5327 4820
rect 5253 4560 5267 4573
rect 5256 4556 5264 4560
rect 5296 4556 5304 4673
rect 5356 4587 5364 4793
rect 5320 4524 5333 4527
rect 5316 4516 5333 4524
rect 5320 4513 5333 4516
rect 5076 4407 5084 4453
rect 5276 4447 5284 4512
rect 5356 4507 5364 4573
rect 5376 4527 5384 4773
rect 5396 4747 5404 4824
rect 5433 4807 5447 4812
rect 5516 4687 5524 4854
rect 5416 4520 5424 4524
rect 5413 4507 5427 4520
rect 5093 4367 5107 4373
rect 5087 4360 5107 4367
rect 5087 4356 5104 4360
rect 5087 4353 5100 4356
rect 5156 4336 5164 4433
rect 5216 4307 5224 4373
rect 5316 4336 5324 4493
rect 5096 4300 5104 4304
rect 5056 4104 5064 4172
rect 5076 4127 5084 4293
rect 5093 4287 5107 4300
rect 5096 4107 5104 4273
rect 5116 4207 5124 4253
rect 5136 4247 5144 4304
rect 5236 4296 5253 4304
rect 5056 4096 5084 4104
rect 4936 3967 4944 4053
rect 4967 4044 4980 4047
rect 4967 4036 4984 4044
rect 5013 4040 5027 4053
rect 5053 4047 5067 4053
rect 5016 4036 5024 4040
rect 4967 4033 4980 4036
rect 4953 3987 4967 3993
rect 4996 3947 5004 4004
rect 5076 3947 5084 4096
rect 5116 4047 5124 4113
rect 5136 4036 5144 4133
rect 5176 4036 5184 4073
rect 5236 4047 5244 4296
rect 5296 4207 5304 4304
rect 5096 3907 5104 4033
rect 4913 3847 4927 3853
rect 4980 3784 4993 3787
rect 4936 3747 4944 3784
rect 4976 3776 4993 3784
rect 4980 3773 4993 3776
rect 4847 3736 4864 3744
rect 4676 3587 4684 3713
rect 4573 3520 4587 3533
rect 4576 3516 4584 3520
rect 4356 3256 4384 3264
rect 4267 3236 4304 3244
rect 4267 3233 4284 3236
rect 4236 3004 4244 3193
rect 4276 3008 4284 3233
rect 4176 2996 4204 3004
rect 4216 2996 4244 3004
rect 4096 2867 4104 2964
rect 4136 2960 4144 2964
rect 4133 2947 4147 2960
rect 4073 2780 4087 2793
rect 4113 2787 4127 2793
rect 4136 2787 4144 2853
rect 4076 2776 4084 2780
rect 4036 2647 4044 2733
rect 4056 2707 4064 2744
rect 4116 2647 4124 2673
rect 4036 2476 4044 2533
rect 4136 2527 4144 2752
rect 4156 2587 4164 2853
rect 4176 2787 4184 2996
rect 4236 2827 4244 2953
rect 4296 2907 4304 2953
rect 4316 2947 4324 3093
rect 4196 2776 4204 2813
rect 4176 2607 4184 2733
rect 4156 2527 4164 2573
rect 4216 2567 4224 2744
rect 4276 2727 4284 2793
rect 4296 2746 4304 2893
rect 4336 2807 4344 3173
rect 4376 3007 4384 3256
rect 4396 3067 4404 3264
rect 4436 2996 4444 3033
rect 4476 2996 4484 3193
rect 4496 3147 4504 3473
rect 4516 3367 4524 3484
rect 4616 3407 4624 3533
rect 4636 3486 4644 3553
rect 4756 3427 4764 3633
rect 4776 3424 4784 3653
rect 4836 3516 4844 3733
rect 4976 3707 4984 3753
rect 4996 3687 5004 3713
rect 4876 3516 4884 3613
rect 4796 3447 4804 3473
rect 4816 3424 4824 3484
rect 4776 3416 4824 3424
rect 4556 3327 4564 3373
rect 4636 3367 4644 3413
rect 4496 3008 4504 3133
rect 4516 3087 4524 3313
rect 4576 3296 4584 3353
rect 4636 3266 4644 3293
rect 4633 3247 4647 3252
rect 4656 3207 4664 3353
rect 4676 3267 4684 3413
rect 4776 3387 4784 3416
rect 4693 3347 4707 3353
rect 4716 3296 4724 3333
rect 4716 3187 4724 3233
rect 4356 2827 4364 2993
rect 4456 2960 4464 2964
rect 4453 2947 4467 2960
rect 4436 2936 4453 2944
rect 4376 2804 4384 2853
rect 4356 2796 4384 2804
rect 4356 2776 4364 2796
rect 4307 2736 4324 2744
rect 4336 2740 4344 2744
rect 4273 2707 4287 2713
rect 4096 2467 4104 2513
rect 4060 2444 4073 2447
rect 4016 2327 4024 2444
rect 4056 2436 4073 2444
rect 4060 2433 4073 2436
rect 4076 2247 4084 2273
rect 3936 1968 3944 1993
rect 3836 1847 3844 1953
rect 3896 1920 3904 1924
rect 3893 1907 3907 1920
rect 3976 1807 3984 2053
rect 3996 1827 4004 2113
rect 4096 1907 4104 2373
rect 4116 2226 4124 2513
rect 4133 2487 4147 2492
rect 4216 2446 4224 2493
rect 4156 2287 4164 2432
rect 4216 2256 4224 2393
rect 4236 2387 4244 2673
rect 4256 2444 4264 2693
rect 4296 2476 4304 2653
rect 4316 2507 4324 2736
rect 4333 2727 4347 2740
rect 4416 2727 4424 2813
rect 4436 2807 4444 2936
rect 4436 2746 4444 2793
rect 4496 2776 4504 2813
rect 4516 2807 4524 3033
rect 4576 2996 4584 3033
rect 4616 2996 4624 3173
rect 4676 3087 4684 3113
rect 4536 2847 4544 2993
rect 4656 2966 4664 3073
rect 4736 3024 4744 3252
rect 4776 3227 4784 3264
rect 4716 3016 4744 3024
rect 4716 2996 4724 3016
rect 4596 2907 4604 2952
rect 4736 2927 4744 2964
rect 4596 2788 4604 2813
rect 4336 2547 4344 2713
rect 4456 2707 4464 2733
rect 4473 2727 4487 2732
rect 4516 2707 4524 2744
rect 4336 2476 4344 2512
rect 4256 2436 4284 2444
rect 4116 1907 4124 2212
rect 4156 2187 4164 2224
rect 4256 2107 4264 2253
rect 4276 2224 4284 2436
rect 4296 2347 4304 2413
rect 4316 2367 4324 2444
rect 4356 2407 4364 2444
rect 4356 2256 4364 2353
rect 4396 2267 4404 2593
rect 4436 2476 4444 2513
rect 4473 2480 4487 2493
rect 4476 2476 4484 2480
rect 4536 2467 4544 2613
rect 4456 2407 4464 2444
rect 4556 2364 4564 2713
rect 4576 2627 4584 2773
rect 4596 2707 4604 2774
rect 4756 2744 4764 2774
rect 4676 2647 4684 2744
rect 4716 2627 4724 2744
rect 4736 2736 4764 2744
rect 4736 2564 4744 2736
rect 4776 2727 4784 2853
rect 4796 2746 4804 2833
rect 4816 2787 4824 3333
rect 4836 3147 4844 3313
rect 4856 3308 4864 3484
rect 4916 3327 4924 3613
rect 4936 3427 4944 3533
rect 4956 3527 4964 3653
rect 4996 3524 5004 3673
rect 5016 3547 5024 3893
rect 5036 3827 5044 3873
rect 5116 3816 5124 3993
rect 5156 3984 5164 4004
rect 5136 3976 5164 3984
rect 5136 3827 5144 3976
rect 5036 3687 5044 3733
rect 5036 3627 5044 3673
rect 4976 3516 5004 3524
rect 5036 3516 5044 3613
rect 5056 3587 5064 3784
rect 5096 3747 5104 3784
rect 5133 3767 5147 3773
rect 5116 3687 5124 3753
rect 4936 3296 4944 3373
rect 4956 3304 4964 3473
rect 5016 3447 5024 3484
rect 5027 3436 5044 3444
rect 4956 3296 4984 3304
rect 4916 3247 4924 3264
rect 4856 2996 4864 3073
rect 4916 3067 4924 3233
rect 4976 3164 4984 3296
rect 4956 3156 4984 3164
rect 4956 3084 4964 3156
rect 4936 3076 4964 3084
rect 4893 3027 4907 3033
rect 4893 3000 4907 3013
rect 4896 2996 4904 3000
rect 4836 2847 4844 2953
rect 4876 2807 4884 2964
rect 4866 2793 4867 2800
rect 4853 2780 4867 2793
rect 4916 2787 4924 2913
rect 4936 2867 4944 3076
rect 4956 2967 4964 3053
rect 4976 2867 4984 3133
rect 4996 3107 5004 3413
rect 5016 3027 5024 3313
rect 5036 3307 5044 3436
rect 5056 3327 5064 3473
rect 5076 3296 5084 3593
rect 5096 3347 5104 3633
rect 5116 3587 5124 3652
rect 5136 3527 5144 3693
rect 5156 3647 5164 3953
rect 5196 3947 5204 4004
rect 5236 3967 5244 3993
rect 5256 3967 5264 4133
rect 5296 4127 5304 4193
rect 5273 4067 5287 4073
rect 5296 4047 5304 4092
rect 5313 4067 5327 4073
rect 5356 4047 5364 4333
rect 5376 4227 5384 4433
rect 5416 4336 5424 4393
rect 5456 4367 5464 4524
rect 5496 4267 5504 4493
rect 5516 4487 5524 4554
rect 5536 4447 5544 4953
rect 5556 4947 5564 5033
rect 5576 5007 5584 5273
rect 5656 5167 5664 5313
rect 5673 5087 5687 5093
rect 5716 5087 5724 5336
rect 5856 5340 5864 5344
rect 5813 5327 5827 5332
rect 5853 5327 5867 5340
rect 5627 5084 5640 5087
rect 5627 5076 5644 5084
rect 5627 5073 5640 5076
rect 5773 5080 5787 5093
rect 5776 5076 5784 5080
rect 5656 5024 5664 5044
rect 5636 5016 5664 5024
rect 5636 4868 5644 5016
rect 5676 4944 5684 5033
rect 5667 4936 5684 4944
rect 5656 4867 5664 4933
rect 5556 4507 5564 4713
rect 5576 4627 5584 4824
rect 5616 4820 5624 4824
rect 5613 4807 5627 4820
rect 5613 4560 5627 4573
rect 5653 4560 5667 4573
rect 5676 4567 5684 4873
rect 5616 4556 5624 4560
rect 5656 4556 5664 4560
rect 5616 4447 5624 4473
rect 5636 4467 5644 4524
rect 5516 4307 5524 4393
rect 5556 4387 5564 4413
rect 5676 4407 5684 4513
rect 5696 4467 5704 5053
rect 5756 5040 5764 5044
rect 5753 5027 5767 5040
rect 5716 4867 5724 5013
rect 5736 4856 5744 4893
rect 5776 4856 5784 4933
rect 5836 4867 5844 5233
rect 5716 4587 5724 4813
rect 5736 4587 5744 4793
rect 5756 4787 5764 4824
rect 5736 4556 5744 4573
rect 5773 4568 5787 4573
rect 5816 4567 5824 4813
rect 5620 4404 5633 4407
rect 5616 4393 5633 4404
rect 5533 4347 5547 4353
rect 5616 4336 5624 4393
rect 5336 4036 5353 4044
rect 5176 3807 5184 3833
rect 5176 3684 5184 3713
rect 5196 3707 5204 3893
rect 5216 3827 5224 3873
rect 5236 3847 5244 3893
rect 5276 3867 5284 4032
rect 5316 3847 5324 3953
rect 5336 3827 5344 3853
rect 5356 3847 5364 3993
rect 5376 3907 5384 4113
rect 5373 3824 5387 3833
rect 5396 3827 5404 4033
rect 5416 3987 5424 4093
rect 5436 4047 5444 4253
rect 5456 4036 5464 4113
rect 5493 4040 5507 4053
rect 5536 4044 5544 4293
rect 5556 4267 5564 4304
rect 5576 4047 5584 4273
rect 5596 4048 5604 4304
rect 5636 4048 5644 4253
rect 5496 4036 5504 4040
rect 5536 4036 5564 4044
rect 5476 3947 5484 4004
rect 5536 3947 5544 3993
rect 5526 3933 5527 3940
rect 5513 3924 5527 3933
rect 5556 3927 5564 4036
rect 5676 4047 5684 4393
rect 5696 4007 5704 4453
rect 5716 4387 5724 4413
rect 5736 4336 5744 4493
rect 5756 4467 5764 4524
rect 5796 4447 5804 4524
rect 5816 4347 5824 4513
rect 5836 4507 5844 4554
rect 5856 4447 5864 5213
rect 5876 4567 5884 5313
rect 5896 5227 5904 5374
rect 5916 4727 5924 5613
rect 5936 4827 5944 5413
rect 5956 5047 5964 5593
rect 5976 4887 5984 5493
rect 5873 4507 5887 4513
rect 5896 4427 5904 4524
rect 5936 4336 5944 4493
rect 5956 4347 5964 4513
rect 5756 4287 5764 4304
rect 5513 3920 5544 3924
rect 5516 3916 5544 3920
rect 5356 3820 5387 3824
rect 5356 3816 5384 3820
rect 5227 3784 5240 3787
rect 5227 3776 5244 3784
rect 5227 3773 5240 3776
rect 5320 3784 5333 3787
rect 5316 3776 5333 3784
rect 5320 3773 5333 3776
rect 5176 3676 5204 3684
rect 5116 3367 5124 3514
rect 5156 3516 5164 3593
rect 5196 3527 5204 3676
rect 5216 3647 5224 3752
rect 5196 3516 5213 3527
rect 5200 3513 5213 3516
rect 5236 3487 5244 3733
rect 5256 3687 5264 3753
rect 5356 3727 5364 3816
rect 5456 3816 5464 3873
rect 5496 3816 5504 3853
rect 5516 3827 5524 3893
rect 5536 3887 5544 3916
rect 5547 3856 5564 3864
rect 5136 3307 5144 3393
rect 5036 3167 5044 3253
rect 5056 3227 5064 3264
rect 5096 3256 5124 3264
rect 5096 3227 5104 3256
rect 5127 3233 5133 3247
rect 5156 3227 5164 3313
rect 5176 3307 5184 3413
rect 5196 3324 5204 3433
rect 5216 3427 5224 3473
rect 5196 3316 5224 3324
rect 5216 3296 5224 3316
rect 5256 3296 5264 3593
rect 5276 3587 5284 3613
rect 5296 3528 5304 3553
rect 5276 3327 5284 3472
rect 5316 3467 5324 3484
rect 5316 3456 5333 3467
rect 5320 3453 5333 3456
rect 5356 3407 5364 3473
rect 5376 3387 5384 3753
rect 5396 3687 5404 3792
rect 5476 3780 5484 3784
rect 5473 3767 5487 3780
rect 5536 3764 5544 3852
rect 5556 3824 5564 3856
rect 5576 3847 5584 3993
rect 5616 3984 5624 4004
rect 5616 3976 5644 3984
rect 5596 3867 5604 3913
rect 5556 3816 5584 3824
rect 5616 3816 5624 3953
rect 5636 3947 5644 3976
rect 5636 3847 5644 3933
rect 5596 3780 5604 3784
rect 5516 3756 5544 3764
rect 5396 3527 5404 3633
rect 5416 3627 5424 3713
rect 5416 3516 5424 3553
rect 5476 3516 5484 3633
rect 5496 3527 5504 3593
rect 5393 3467 5407 3473
rect 5187 3264 5200 3267
rect 5187 3256 5204 3264
rect 5187 3253 5200 3256
rect 5056 3067 5064 3213
rect 5016 2996 5024 3013
rect 5096 2884 5104 3153
rect 5116 2947 5124 3212
rect 5176 3187 5184 3232
rect 5196 3167 5204 3213
rect 5216 3187 5224 3233
rect 5156 2996 5164 3153
rect 5196 3087 5204 3153
rect 5196 2996 5204 3073
rect 5216 3007 5224 3093
rect 5176 2960 5184 2964
rect 5096 2876 5124 2884
rect 4856 2776 4864 2780
rect 4727 2556 4744 2564
rect 4716 2487 4724 2553
rect 4736 2427 4744 2474
rect 4656 2400 4664 2404
rect 4653 2387 4667 2400
rect 4556 2356 4584 2364
rect 4513 2260 4527 2273
rect 4516 2256 4524 2260
rect 4276 2216 4304 2224
rect 3496 1736 3524 1744
rect 3476 1706 3484 1733
rect 3396 1687 3404 1704
rect 3396 1567 3404 1673
rect 3227 1476 3244 1484
rect 3236 1407 3244 1476
rect 3176 1327 3184 1392
rect 3227 1386 3240 1387
rect 3227 1373 3233 1386
rect 3256 1347 3264 1493
rect 3360 1444 3373 1447
rect 3356 1436 3373 1444
rect 3360 1433 3373 1436
rect 3273 1367 3287 1373
rect 3336 1347 3344 1404
rect 3376 1367 3384 1393
rect 3396 1347 3404 1553
rect 3456 1487 3464 1593
rect 3416 1227 3424 1453
rect 3456 1436 3464 1473
rect 3496 1436 3504 1736
rect 3536 1667 3544 1704
rect 3576 1700 3584 1704
rect 3573 1687 3587 1700
rect 3656 1527 3664 1773
rect 3876 1736 3884 1793
rect 3696 1667 3704 1704
rect 3736 1607 3744 1704
rect 3636 1516 3653 1524
rect 3476 1400 3484 1404
rect 3433 1387 3447 1393
rect 3473 1387 3487 1400
rect 3176 1216 3224 1224
rect 3156 1047 3164 1172
rect 3053 920 3067 933
rect 3096 927 3104 973
rect 3056 916 3064 920
rect 3176 887 3184 1153
rect 3336 987 3344 1184
rect 3393 1167 3407 1170
rect 3036 847 3044 884
rect 3076 824 3084 884
rect 3196 847 3204 916
rect 3076 816 3104 824
rect 3056 696 3064 733
rect 3096 667 3104 816
rect 3176 696 3184 813
rect 3336 807 3344 916
rect 3156 627 3164 664
rect 3196 607 3204 664
rect 3036 396 3044 473
rect 2976 366 2984 393
rect 2876 176 2884 213
rect 2896 207 2904 364
rect 2596 136 2644 144
rect 1896 -16 1904 113
rect 2936 -16 2944 193
rect 3016 176 3024 313
rect 3056 227 3064 364
rect 3096 327 3104 353
rect 3136 264 3144 413
rect 3156 366 3164 453
rect 3196 396 3204 593
rect 3256 427 3264 793
rect 3287 756 3313 764
rect 3296 696 3304 733
rect 3356 487 3364 1053
rect 3396 916 3404 1033
rect 3416 947 3424 1093
rect 3436 1067 3444 1333
rect 3456 1187 3464 1233
rect 3496 1216 3504 1313
rect 3576 1027 3584 1273
rect 3596 1186 3604 1313
rect 3636 1287 3644 1516
rect 3676 1436 3684 1473
rect 3733 1440 3747 1453
rect 3736 1436 3744 1440
rect 3776 1307 3784 1733
rect 3836 1507 3844 1704
rect 3796 1404 3804 1433
rect 3816 1407 3824 1473
rect 3896 1436 3904 1513
rect 3936 1464 3944 1793
rect 3956 1706 3964 1773
rect 4036 1647 4044 1704
rect 3936 1456 3964 1464
rect 3876 1367 3884 1404
rect 3936 1367 3944 1434
rect 3656 1216 3664 1253
rect 3736 1180 3744 1184
rect 3733 1167 3747 1180
rect 3796 1147 3804 1184
rect 3836 1047 3844 1273
rect 3856 1186 3864 1293
rect 3436 916 3444 973
rect 3376 667 3384 873
rect 3456 880 3464 884
rect 3453 867 3467 880
rect 3476 696 3484 853
rect 3493 847 3507 853
rect 3376 396 3384 453
rect 3316 287 3324 364
rect 3136 256 3164 264
rect 3156 187 3164 256
rect 2956 147 2964 176
rect 3176 144 3184 213
rect 3416 187 3424 653
rect 3036 107 3044 144
rect 3036 47 3044 93
rect 3356 27 3364 133
rect 3436 127 3444 473
rect 3456 366 3464 664
rect 3516 627 3524 1013
rect 3836 928 3844 1033
rect 3636 880 3644 884
rect 3633 867 3647 880
rect 3653 844 3667 853
rect 3627 840 3667 844
rect 3627 836 3664 840
rect 3696 707 3704 914
rect 3956 927 3964 1456
rect 3976 1247 3984 1593
rect 4076 1467 4084 1753
rect 4116 1736 4124 1833
rect 4136 1807 4144 2093
rect 4176 1956 4184 2073
rect 4256 1967 4264 2093
rect 4196 1920 4204 1924
rect 4193 1907 4207 1920
rect 4153 1740 4167 1753
rect 4156 1736 4164 1740
rect 4216 1707 4224 1793
rect 4136 1667 4144 1704
rect 4216 1647 4224 1693
rect 4076 1327 4084 1404
rect 4076 1287 4084 1313
rect 4096 1307 4104 1393
rect 4116 1387 4124 1453
rect 4156 1436 4164 1493
rect 4236 1444 4244 1924
rect 4256 1707 4264 1913
rect 4276 1847 4284 1954
rect 4296 1867 4304 2216
rect 4336 2167 4344 2224
rect 4376 2207 4384 2224
rect 4416 2207 4424 2233
rect 4356 2067 4364 2193
rect 4373 2187 4387 2193
rect 4356 1956 4364 2013
rect 4316 1926 4324 1953
rect 4376 1887 4384 1912
rect 4416 1907 4424 2172
rect 4456 2167 4464 2224
rect 4456 1867 4464 1924
rect 4376 1736 4384 1773
rect 4256 1667 4264 1693
rect 4356 1547 4364 1684
rect 4436 1567 4444 1853
rect 4516 1847 4524 2173
rect 4556 1964 4564 2253
rect 4576 2087 4584 2356
rect 4596 2226 4604 2353
rect 4627 2264 4640 2267
rect 4627 2256 4644 2264
rect 4627 2253 4640 2256
rect 4716 2267 4724 2293
rect 4756 2264 4764 2633
rect 4776 2307 4784 2573
rect 4796 2527 4804 2732
rect 4836 2707 4844 2744
rect 4936 2727 4944 2793
rect 5016 2776 5024 2813
rect 5053 2780 5067 2793
rect 5076 2787 5084 2873
rect 5056 2776 5064 2780
rect 4896 2487 4904 2633
rect 4916 2547 4924 2673
rect 4936 2488 4944 2713
rect 4956 2507 4964 2773
rect 4987 2744 5000 2747
rect 4987 2736 5004 2744
rect 5036 2740 5044 2744
rect 4987 2733 5000 2736
rect 5033 2727 5047 2740
rect 4996 2507 5004 2613
rect 4916 2476 4933 2484
rect 4836 2327 4844 2444
rect 4876 2440 4884 2444
rect 4873 2427 4887 2440
rect 4916 2446 4924 2476
rect 5016 2487 5024 2613
rect 4796 2268 4804 2313
rect 4736 2256 4764 2264
rect 4656 2167 4664 2224
rect 4696 2107 4704 2212
rect 4536 1956 4564 1964
rect 4536 1926 4544 1956
rect 4676 1927 4684 1954
rect 4236 1436 4264 1444
rect 4196 1400 4204 1404
rect 4193 1387 4207 1400
rect 4216 1327 4224 1353
rect 4236 1307 4244 1333
rect 4256 1287 4264 1436
rect 4316 1436 4324 1493
rect 4276 1347 4284 1433
rect 4336 1396 4364 1404
rect 4293 1327 4307 1333
rect 4093 1220 4107 1233
rect 4096 1216 4104 1220
rect 3996 1087 4004 1214
rect 4076 1164 4084 1184
rect 4056 1156 4084 1164
rect 4056 928 4064 1156
rect 4136 1147 4144 1253
rect 4336 1247 4344 1396
rect 4356 1216 4364 1253
rect 4396 1247 4404 1353
rect 4396 1216 4404 1233
rect 4416 1224 4424 1353
rect 4436 1307 4444 1433
rect 4416 1216 4444 1224
rect 4216 1047 4224 1184
rect 4296 1167 4304 1213
rect 4436 1186 4444 1216
rect 4336 1180 4344 1184
rect 4333 1167 4347 1180
rect 4236 916 4244 1073
rect 3776 880 3784 884
rect 3773 867 3787 880
rect 3816 867 3824 884
rect 3807 856 3824 867
rect 3807 853 3820 856
rect 3856 707 3864 872
rect 3876 867 3884 913
rect 3927 753 3933 767
rect 3967 753 3973 767
rect 3996 744 4004 913
rect 4076 880 4084 884
rect 4073 867 4087 880
rect 4116 880 4124 884
rect 3976 736 4004 744
rect 3756 696 3804 704
rect 3576 607 3584 664
rect 3796 607 3804 696
rect 3873 700 3887 713
rect 3876 696 3884 700
rect 3936 667 3944 732
rect 3807 596 3824 604
rect 3496 396 3504 553
rect 3753 400 3767 413
rect 3793 400 3807 413
rect 3816 407 3824 596
rect 3856 427 3864 653
rect 3976 464 3984 736
rect 3996 720 4044 724
rect 3993 716 4044 720
rect 3993 707 4007 716
rect 4036 696 4044 716
rect 4096 704 4104 873
rect 4113 867 4127 880
rect 4196 807 4204 893
rect 4096 696 4113 704
rect 4193 704 4207 713
rect 4216 704 4224 773
rect 4193 700 4224 704
rect 4196 696 4224 700
rect 4116 667 4124 694
rect 3976 456 4004 464
rect 3756 396 3764 400
rect 3796 396 3804 400
rect 3873 404 3887 413
rect 3867 400 3887 404
rect 3913 400 3927 413
rect 3867 396 3884 400
rect 3916 396 3924 400
rect 3856 366 3864 392
rect 3976 366 3984 433
rect 3516 227 3524 364
rect 3456 27 3464 213
rect 3596 146 3604 213
rect 3696 176 3704 213
rect 3516 140 3524 144
rect 3513 127 3527 140
rect 3636 87 3644 173
rect 3856 167 3864 213
rect 3676 140 3684 144
rect 3673 127 3687 140
rect 3716 107 3724 144
rect 3816 87 3824 144
rect 3876 107 3884 176
rect 3707 76 3733 84
rect 3996 47 4004 456
rect 4080 204 4093 207
rect 4076 193 4093 204
rect 4076 176 4084 193
rect 4116 188 4124 613
rect 4176 607 4184 664
rect 4236 427 4244 853
rect 4336 747 4344 913
rect 4356 867 4364 1153
rect 4456 1047 4464 1832
rect 4576 1747 4584 1893
rect 4476 1607 4484 1733
rect 4516 1700 4524 1704
rect 4496 1464 4504 1693
rect 4513 1687 4527 1700
rect 4596 1706 4604 1912
rect 4636 1744 4644 1924
rect 4616 1736 4644 1744
rect 4656 1736 4664 1813
rect 4676 1804 4684 1873
rect 4696 1867 4704 1973
rect 4716 1926 4724 2213
rect 4736 1987 4744 2256
rect 4833 2260 4847 2273
rect 4856 2267 4864 2293
rect 4836 2256 4844 2260
rect 4876 2226 4884 2253
rect 4776 1968 4784 2013
rect 4816 1956 4824 2212
rect 4856 2004 4864 2213
rect 4836 1996 4864 2004
rect 4836 1967 4844 1996
rect 4896 1987 4904 2433
rect 5000 2444 5013 2447
rect 4996 2440 5013 2444
rect 4993 2433 5013 2440
rect 4993 2427 5007 2433
rect 5036 2367 5044 2473
rect 4916 2007 4924 2273
rect 4996 2256 5004 2313
rect 4976 2187 4984 2224
rect 4736 1887 4744 1913
rect 4796 1887 4804 1924
rect 4676 1796 4704 1804
rect 4696 1748 4704 1796
rect 4496 1456 4524 1464
rect 4516 1436 4524 1456
rect 4576 1447 4584 1693
rect 4616 1687 4624 1736
rect 4676 1700 4684 1704
rect 4673 1687 4687 1700
rect 4756 1687 4764 1793
rect 4856 1787 4864 1973
rect 4976 1956 4984 2152
rect 4876 1747 4884 1953
rect 4896 1706 4904 1773
rect 4956 1747 4964 1773
rect 4976 1736 4984 1833
rect 5016 1787 5024 2053
rect 5056 2027 5064 2493
rect 5076 2344 5084 2733
rect 5096 2627 5104 2853
rect 5116 2787 5124 2876
rect 5136 2807 5144 2953
rect 5173 2947 5187 2960
rect 5176 2807 5184 2933
rect 5196 2887 5204 2933
rect 5166 2793 5167 2800
rect 5153 2780 5167 2793
rect 5156 2776 5164 2780
rect 5116 2587 5124 2733
rect 5136 2687 5144 2744
rect 5216 2587 5224 2953
rect 5096 2387 5104 2412
rect 5076 2336 5104 2344
rect 5076 2226 5084 2313
rect 5096 2267 5104 2336
rect 5156 2287 5164 2404
rect 5136 2276 5153 2284
rect 5136 2268 5144 2276
rect 5176 2256 5184 2353
rect 5196 2267 5204 2373
rect 5096 2147 5104 2213
rect 5216 2226 5224 2273
rect 5196 2187 5204 2213
rect 5036 1926 5044 1993
rect 5053 1967 5067 1973
rect 5073 1960 5087 1973
rect 5113 1960 5127 1973
rect 5076 1956 5084 1960
rect 5116 1956 5124 1960
rect 5136 1867 5144 1924
rect 4836 1700 4844 1704
rect 4833 1687 4847 1700
rect 4496 1244 4504 1404
rect 4536 1347 4544 1404
rect 4476 1240 4504 1244
rect 4473 1236 4504 1240
rect 4473 1227 4487 1236
rect 4513 1220 4527 1233
rect 4516 1216 4524 1220
rect 4556 1216 4564 1293
rect 4596 1224 4604 1553
rect 4616 1244 4624 1533
rect 4633 1427 4647 1433
rect 4796 1427 4804 1553
rect 4636 1267 4644 1421
rect 4616 1236 4644 1244
rect 4596 1216 4624 1224
rect 4496 1180 4504 1184
rect 4493 1167 4507 1180
rect 4536 1144 4544 1184
rect 4536 1136 4564 1144
rect 4376 787 4384 913
rect 4436 876 4484 884
rect 4536 867 4544 1113
rect 4556 787 4564 1136
rect 4616 1127 4624 1216
rect 4636 1087 4644 1236
rect 4676 1216 4684 1333
rect 4696 1327 4704 1364
rect 4716 1216 4724 1313
rect 4776 1307 4784 1413
rect 4816 1364 4824 1593
rect 4916 1527 4924 1733
rect 4936 1587 4944 1733
rect 4996 1567 5004 1704
rect 4816 1356 4844 1364
rect 4596 916 4604 953
rect 4653 920 4667 933
rect 4656 916 4664 920
rect 4476 707 4484 773
rect 4136 367 4144 394
rect 4236 387 4244 413
rect 4296 396 4304 433
rect 4316 427 4324 664
rect 4356 366 4364 653
rect 4567 656 4584 664
rect 4496 396 4504 613
rect 4576 404 4584 656
rect 4596 527 4604 853
rect 4696 827 4704 1184
rect 4776 1147 4784 1253
rect 4816 1216 4824 1333
rect 4836 1247 4844 1356
rect 4976 1327 4984 1413
rect 4996 1347 5004 1513
rect 4716 847 4724 953
rect 4836 947 4844 1184
rect 4773 928 4787 933
rect 4616 664 4624 733
rect 4676 696 4684 753
rect 4696 587 4704 664
rect 4736 627 4744 664
rect 4776 627 4784 853
rect 4796 847 4804 884
rect 4836 827 4844 884
rect 4856 827 4864 873
rect 4876 707 4884 1233
rect 4933 1220 4947 1233
rect 4936 1216 4944 1220
rect 4976 1216 4984 1313
rect 5016 1224 5024 1673
rect 5036 1547 5044 1704
rect 5053 1687 5067 1693
rect 5076 1468 5084 1813
rect 5136 1787 5144 1853
rect 5176 1827 5184 2013
rect 5096 1706 5104 1773
rect 5153 1740 5167 1753
rect 5196 1747 5204 2093
rect 5236 1987 5244 3193
rect 5256 3027 5264 3233
rect 5276 3167 5284 3264
rect 5316 3247 5324 3333
rect 5336 3127 5344 3373
rect 5413 3347 5427 3353
rect 5407 3340 5427 3347
rect 5407 3336 5424 3340
rect 5407 3333 5420 3336
rect 5373 3300 5387 3313
rect 5376 3296 5384 3300
rect 5436 3304 5444 3473
rect 5456 3407 5464 3484
rect 5436 3296 5464 3304
rect 5376 3067 5384 3213
rect 5396 3087 5404 3264
rect 5256 2904 5264 2973
rect 5256 2896 5273 2904
rect 5276 2804 5284 2893
rect 5336 2867 5344 2924
rect 5276 2796 5304 2804
rect 5296 2776 5304 2796
rect 5256 2467 5264 2553
rect 5316 2488 5324 2733
rect 5336 2647 5344 2744
rect 5376 2727 5384 2853
rect 5396 2607 5404 2813
rect 5416 2727 5424 3113
rect 5436 3008 5444 3253
rect 5456 3247 5464 3296
rect 5456 3027 5464 3073
rect 5476 3047 5484 3373
rect 5496 3307 5504 3473
rect 5516 3447 5524 3756
rect 5536 3308 5544 3553
rect 5556 3467 5564 3773
rect 5593 3767 5607 3780
rect 5576 3707 5584 3753
rect 5636 3707 5644 3784
rect 5656 3727 5664 3773
rect 5576 3527 5584 3693
rect 5676 3667 5684 3853
rect 5696 3647 5704 3972
rect 5716 3827 5724 4033
rect 5736 3987 5744 4093
rect 5756 4047 5764 4273
rect 5796 4207 5804 4304
rect 5816 4147 5824 4293
rect 5836 4207 5844 4334
rect 5976 4327 5984 4373
rect 5876 4300 5884 4304
rect 5873 4287 5887 4300
rect 5793 4040 5807 4053
rect 5796 4036 5804 4040
rect 5836 4036 5844 4093
rect 5856 4047 5864 4213
rect 5776 3984 5784 4004
rect 5776 3976 5804 3984
rect 5756 3816 5764 3893
rect 5776 3887 5784 3953
rect 5796 3907 5804 3976
rect 5816 3967 5824 3992
rect 5793 3820 5807 3833
rect 5796 3816 5804 3820
rect 5736 3780 5744 3784
rect 5733 3767 5747 3780
rect 5776 3727 5784 3784
rect 5656 3516 5664 3553
rect 5756 3516 5764 3553
rect 5576 3387 5584 3473
rect 5596 3447 5604 3484
rect 5556 3327 5564 3353
rect 5516 3260 5524 3264
rect 5496 3067 5504 3253
rect 5513 3247 5527 3260
rect 5556 3227 5564 3264
rect 5536 3107 5544 3173
rect 5556 3147 5564 3192
rect 5496 3008 5504 3032
rect 5556 3007 5564 3053
rect 5433 2947 5447 2953
rect 5476 2907 5484 2964
rect 5516 2847 5524 2964
rect 5556 2907 5564 2953
rect 5576 2907 5584 3253
rect 5596 3187 5604 3293
rect 5596 3008 5604 3173
rect 5616 3147 5624 3453
rect 5636 3227 5644 3484
rect 5696 3467 5704 3514
rect 5836 3484 5844 3713
rect 5856 3607 5864 3993
rect 5876 3987 5884 4193
rect 5896 3947 5904 4253
rect 5916 4107 5924 4292
rect 5956 4267 5964 4293
rect 5927 4064 5940 4067
rect 5927 4053 5944 4064
rect 5936 4036 5944 4053
rect 5976 4047 5984 4153
rect 5956 3996 5984 4004
rect 5976 3987 5984 3996
rect 5736 3480 5744 3484
rect 5733 3467 5747 3480
rect 5746 3460 5747 3467
rect 5656 3307 5664 3373
rect 5696 3327 5704 3353
rect 5696 3296 5704 3313
rect 5756 3307 5764 3453
rect 5776 3344 5784 3484
rect 5816 3476 5844 3484
rect 5816 3367 5824 3476
rect 5856 3387 5864 3553
rect 5776 3336 5804 3344
rect 5676 3107 5684 3264
rect 5636 3007 5644 3093
rect 5656 2996 5664 3073
rect 5676 3027 5684 3053
rect 5696 3047 5704 3233
rect 5716 3067 5724 3264
rect 5776 3227 5784 3313
rect 5796 3307 5804 3336
rect 5833 3300 5847 3313
rect 5876 3308 5884 3753
rect 5836 3296 5844 3300
rect 5896 3307 5904 3653
rect 5696 3007 5704 3033
rect 5716 3027 5724 3053
rect 5436 2787 5444 2813
rect 5513 2780 5527 2793
rect 5516 2776 5524 2780
rect 5596 2776 5604 2833
rect 5616 2827 5624 2993
rect 5636 2776 5644 2853
rect 5456 2740 5464 2744
rect 5496 2740 5504 2744
rect 5396 2507 5404 2593
rect 5256 2267 5264 2313
rect 5296 2288 5304 2433
rect 5336 2304 5344 2444
rect 5376 2440 5384 2444
rect 5373 2427 5387 2440
rect 5336 2296 5364 2304
rect 5333 2260 5347 2273
rect 5356 2267 5364 2296
rect 5336 2256 5344 2260
rect 5356 2167 5364 2213
rect 5236 1956 5244 1973
rect 5276 1956 5284 2013
rect 5256 1767 5264 1912
rect 5276 1787 5284 1893
rect 5296 1887 5304 1924
rect 5336 1907 5344 2133
rect 5376 2027 5384 2293
rect 5396 2007 5404 2433
rect 5416 2107 5424 2673
rect 5436 2507 5444 2733
rect 5453 2727 5467 2740
rect 5493 2727 5507 2740
rect 5453 2480 5467 2493
rect 5456 2476 5464 2480
rect 5496 2476 5504 2633
rect 5436 2267 5444 2433
rect 5476 2327 5484 2444
rect 5536 2364 5544 2573
rect 5556 2547 5564 2773
rect 5616 2527 5624 2744
rect 5556 2427 5564 2512
rect 5653 2488 5667 2493
rect 5666 2480 5667 2488
rect 5676 2487 5684 2813
rect 5696 2687 5704 2853
rect 5716 2807 5724 3013
rect 5736 3007 5744 3113
rect 5776 3008 5784 3213
rect 5796 3004 5804 3253
rect 5816 3087 5824 3252
rect 5856 3244 5864 3264
rect 5836 3236 5864 3244
rect 5836 3187 5844 3236
rect 5796 2996 5824 3004
rect 5756 2960 5764 2964
rect 5736 2827 5744 2953
rect 5753 2947 5767 2960
rect 5816 2924 5824 2996
rect 5836 2944 5844 3093
rect 5876 2996 5884 3073
rect 5896 3027 5904 3253
rect 5916 3127 5924 3293
rect 5936 3107 5944 3893
rect 5913 3000 5927 3013
rect 5956 3007 5964 3933
rect 5976 3527 5984 3973
rect 5976 3207 5984 3253
rect 5916 2996 5924 3000
rect 5836 2936 5864 2944
rect 5796 2916 5824 2924
rect 5796 2807 5804 2916
rect 5716 2784 5724 2793
rect 5716 2776 5744 2784
rect 5816 2787 5824 2893
rect 5756 2740 5764 2744
rect 5753 2727 5767 2740
rect 5796 2627 5804 2744
rect 5836 2707 5844 2913
rect 5756 2476 5764 2533
rect 5793 2480 5807 2493
rect 5796 2476 5804 2480
rect 5596 2440 5604 2444
rect 5576 2387 5584 2433
rect 5593 2427 5607 2440
rect 5536 2356 5564 2364
rect 5476 2256 5484 2292
rect 5513 2260 5527 2273
rect 5516 2256 5524 2260
rect 5456 2127 5464 2224
rect 5296 1764 5304 1873
rect 5276 1756 5304 1764
rect 5156 1736 5164 1740
rect 5176 1700 5184 1704
rect 5173 1687 5187 1700
rect 5116 1507 5124 1573
rect 5136 1487 5144 1671
rect 5196 1664 5204 1693
rect 5216 1687 5224 1753
rect 5276 1736 5284 1756
rect 5316 1736 5324 1793
rect 5336 1787 5344 1853
rect 5296 1700 5304 1704
rect 5293 1687 5307 1700
rect 5176 1656 5204 1664
rect 5113 1440 5127 1453
rect 5136 1447 5144 1473
rect 5116 1436 5124 1440
rect 5047 1404 5060 1407
rect 5047 1396 5064 1404
rect 5047 1393 5060 1396
rect 5133 1387 5147 1393
rect 5067 1373 5073 1387
rect 5016 1216 5044 1224
rect 4816 607 4824 664
rect 4556 396 4584 404
rect 4616 396 4624 573
rect 4653 400 4667 413
rect 4693 407 4707 413
rect 4656 396 4664 400
rect 4536 367 4544 394
rect 4136 146 4144 353
rect 4276 184 4284 352
rect 4436 267 4444 364
rect 4476 307 4484 364
rect 4556 227 4564 396
rect 4756 396 4764 433
rect 4276 176 4304 184
rect 4356 147 4364 174
rect 4556 167 4564 213
rect 4616 176 4624 293
rect 4056 107 4064 144
rect 4156 107 4164 133
rect 4236 107 4244 144
rect 4676 146 4684 353
rect 4696 127 4704 393
rect 4796 366 4804 533
rect 4876 467 4884 653
rect 4896 507 4904 1033
rect 4916 927 4924 1173
rect 4996 1107 5004 1184
rect 4993 920 5007 933
rect 5016 927 5024 1073
rect 4996 916 5004 920
rect 4927 884 4940 887
rect 4927 876 4944 884
rect 4927 873 4940 876
rect 4916 666 4924 852
rect 4916 427 4924 652
rect 4936 607 4944 853
rect 4976 827 4984 884
rect 5036 807 5044 1216
rect 5136 1227 5144 1333
rect 5056 1127 5064 1214
rect 5056 847 5064 1113
rect 5076 724 5084 993
rect 5116 947 5124 1184
rect 5136 1127 5144 1173
rect 5136 916 5144 1053
rect 5156 1007 5164 1453
rect 5176 1167 5184 1656
rect 5296 1587 5304 1652
rect 5316 1607 5324 1673
rect 5256 1447 5264 1493
rect 5236 1367 5244 1392
rect 5276 1248 5284 1493
rect 5316 1448 5324 1533
rect 5336 1487 5344 1693
rect 5356 1507 5364 1973
rect 5456 1967 5464 1993
rect 5376 1707 5384 1953
rect 5416 1847 5424 1924
rect 5456 1827 5464 1912
rect 5376 1527 5384 1573
rect 5336 1464 5344 1473
rect 5336 1456 5364 1464
rect 5356 1436 5364 1456
rect 5233 1220 5247 1233
rect 5296 1227 5304 1393
rect 5336 1307 5344 1404
rect 5396 1324 5404 1813
rect 5476 1767 5484 2193
rect 5507 1973 5513 1987
rect 5536 1956 5544 2033
rect 5556 2027 5564 2356
rect 5576 2267 5584 2313
rect 5636 2307 5644 2444
rect 5593 2260 5607 2273
rect 5596 2256 5604 2260
rect 5656 2220 5664 2224
rect 5653 2207 5667 2220
rect 5696 2047 5704 2253
rect 5573 1960 5587 1973
rect 5576 1956 5584 1960
rect 5413 1747 5427 1753
rect 5496 1736 5504 1913
rect 5516 1824 5524 1913
rect 5556 1827 5564 1924
rect 5516 1816 5544 1824
rect 5536 1804 5544 1816
rect 5536 1796 5564 1804
rect 5516 1747 5524 1793
rect 5427 1704 5440 1707
rect 5427 1696 5444 1704
rect 5427 1693 5440 1696
rect 5376 1316 5404 1324
rect 5236 1216 5244 1220
rect 5193 1167 5207 1173
rect 5176 987 5184 1113
rect 5173 920 5187 933
rect 5196 927 5204 1013
rect 5176 916 5184 920
rect 5096 767 5104 873
rect 5076 716 5104 724
rect 5096 647 5104 716
rect 5116 666 5124 793
rect 5196 724 5204 873
rect 5216 807 5224 1151
rect 5256 1027 5264 1184
rect 5296 1007 5304 1173
rect 5236 927 5244 973
rect 5316 967 5324 1273
rect 5376 1247 5384 1316
rect 5276 916 5284 953
rect 5313 920 5327 932
rect 5336 927 5344 1233
rect 5316 916 5324 920
rect 5236 747 5244 873
rect 5133 707 5147 713
rect 5176 716 5204 724
rect 5176 696 5184 716
rect 5213 708 5227 713
rect 5196 660 5204 664
rect 4816 347 4824 394
rect 4916 307 4924 364
rect 4896 188 4904 253
rect 4936 247 4944 353
rect 4736 140 4744 144
rect 4733 127 4747 140
rect 4776 107 4784 144
rect 4856 140 4884 144
rect 4853 136 4884 140
rect 4853 127 4867 136
rect 4956 107 4964 413
rect 4976 267 4984 593
rect 5013 547 5027 553
rect 4976 147 4984 232
rect 4996 188 5004 453
rect 5076 396 5084 453
rect 5096 407 5104 633
rect 5056 360 5064 364
rect 5053 347 5067 360
rect 5116 207 5124 652
rect 5156 396 5164 652
rect 5193 647 5207 660
rect 5236 587 5244 633
rect 5193 400 5207 413
rect 5196 396 5204 400
rect 5136 147 5144 353
rect 5216 176 5224 364
rect 5233 347 5247 352
rect 5256 307 5264 833
rect 5296 704 5304 884
rect 5356 767 5364 1233
rect 5396 1216 5404 1293
rect 5416 1247 5424 1593
rect 5436 1248 5444 1673
rect 5476 1607 5484 1704
rect 5476 1436 5484 1553
rect 5516 1447 5524 1693
rect 5536 1467 5544 1773
rect 5556 1747 5564 1796
rect 5596 1736 5604 1873
rect 5636 1847 5644 1953
rect 5656 1807 5664 2013
rect 5556 1547 5564 1693
rect 5576 1667 5584 1704
rect 5596 1587 5604 1673
rect 5616 1627 5624 1704
rect 5656 1667 5664 1693
rect 5527 1436 5544 1444
rect 5496 1307 5504 1404
rect 5576 1406 5584 1453
rect 5596 1444 5604 1513
rect 5676 1487 5684 1973
rect 5696 1967 5704 2012
rect 5716 1987 5724 2473
rect 5736 2267 5744 2293
rect 5776 2268 5784 2353
rect 5816 2327 5824 2444
rect 5796 2220 5804 2224
rect 5736 2087 5744 2193
rect 5736 1956 5744 2073
rect 5756 1987 5764 2212
rect 5793 2207 5807 2220
rect 5856 2207 5864 2936
rect 5876 2787 5884 2873
rect 5916 2827 5924 2933
rect 5936 2807 5944 2964
rect 5956 2927 5964 2953
rect 5976 2867 5984 3133
rect 5776 1987 5784 2193
rect 5796 2127 5804 2193
rect 5876 2087 5884 2713
rect 5776 1956 5784 1973
rect 5796 1967 5804 2033
rect 5876 1984 5884 2073
rect 5896 2007 5904 2711
rect 5916 2027 5924 2673
rect 5936 2647 5944 2732
rect 5936 2307 5944 2633
rect 5876 1976 5904 1984
rect 5716 1807 5724 1924
rect 5816 1907 5824 1973
rect 5853 1968 5867 1973
rect 5896 1956 5904 1976
rect 5936 1967 5944 2253
rect 5876 1920 5884 1924
rect 5873 1907 5887 1920
rect 5696 1604 5704 1793
rect 5716 1727 5724 1793
rect 5736 1747 5744 1853
rect 5756 1736 5764 1773
rect 5796 1748 5804 1873
rect 5696 1596 5724 1604
rect 5596 1436 5624 1444
rect 5653 1440 5667 1453
rect 5696 1447 5704 1573
rect 5656 1436 5664 1440
rect 5416 1180 5424 1184
rect 5376 847 5384 1173
rect 5413 1167 5427 1180
rect 5456 1147 5464 1173
rect 5456 967 5464 1112
rect 5427 944 5440 947
rect 5427 933 5444 944
rect 5436 916 5444 933
rect 5476 927 5484 1233
rect 5496 1227 5504 1293
rect 5516 1247 5524 1393
rect 5536 1216 5544 1253
rect 5576 1227 5584 1353
rect 5576 1147 5584 1173
rect 5496 947 5504 1093
rect 5316 724 5324 753
rect 5376 744 5384 773
rect 5336 736 5384 744
rect 5396 744 5404 913
rect 5456 880 5464 884
rect 5453 867 5467 880
rect 5476 747 5484 873
rect 5496 747 5504 933
rect 5516 887 5524 1053
rect 5536 927 5544 993
rect 5596 987 5604 1333
rect 5676 1307 5684 1404
rect 5613 1247 5627 1253
rect 5696 1247 5704 1393
rect 5716 1347 5724 1596
rect 5756 1504 5764 1653
rect 5776 1547 5784 1704
rect 5756 1496 5784 1504
rect 5716 1227 5724 1293
rect 5616 1147 5624 1212
rect 5616 1136 5633 1147
rect 5620 1133 5633 1136
rect 5573 944 5587 953
rect 5573 940 5604 944
rect 5576 936 5604 940
rect 5553 920 5567 933
rect 5556 916 5564 920
rect 5596 916 5604 936
rect 5396 736 5424 744
rect 5336 724 5344 736
rect 5316 716 5344 724
rect 5276 696 5304 704
rect 5336 696 5344 716
rect 5276 647 5284 696
rect 5276 287 5284 612
rect 5316 607 5324 652
rect 5356 644 5364 664
rect 5356 636 5384 644
rect 5333 627 5347 633
rect 5333 400 5347 413
rect 5336 396 5344 400
rect 5296 327 5304 353
rect 5316 184 5324 352
rect 5376 347 5384 636
rect 5396 227 5404 413
rect 5416 407 5424 736
rect 5456 667 5464 733
rect 5536 728 5544 873
rect 5620 884 5633 887
rect 5616 876 5633 884
rect 5620 873 5633 876
rect 5453 400 5467 413
rect 5456 396 5464 400
rect 5436 327 5444 364
rect 5496 327 5504 613
rect 5556 587 5564 653
rect 5576 647 5584 793
rect 5596 707 5604 833
rect 5616 787 5624 813
rect 5616 696 5624 733
rect 5636 724 5644 852
rect 5656 787 5664 973
rect 5676 887 5684 1153
rect 5696 1087 5704 1184
rect 5716 916 5724 1013
rect 5736 947 5744 1453
rect 5756 924 5764 1473
rect 5776 1447 5784 1496
rect 5796 1436 5804 1673
rect 5816 1467 5824 1692
rect 5836 1436 5844 1493
rect 5856 1467 5864 1873
rect 5876 1667 5884 1793
rect 5896 1607 5904 1773
rect 5876 1444 5884 1533
rect 5916 1507 5924 1924
rect 5936 1706 5944 1913
rect 5876 1436 5904 1444
rect 5776 1227 5784 1393
rect 5896 1404 5904 1436
rect 5856 1304 5864 1404
rect 5876 1396 5904 1404
rect 5876 1304 5884 1396
rect 5856 1296 5884 1304
rect 5816 1216 5824 1253
rect 5796 1180 5804 1184
rect 5776 947 5784 1173
rect 5793 1167 5807 1180
rect 5836 1147 5844 1184
rect 5816 928 5824 1113
rect 5856 987 5864 1173
rect 5876 1127 5884 1296
rect 5756 916 5784 924
rect 5776 727 5784 916
rect 5853 920 5867 933
rect 5896 927 5904 1373
rect 5916 1087 5924 1253
rect 5856 916 5864 920
rect 5880 884 5893 887
rect 5836 827 5844 884
rect 5876 876 5893 884
rect 5880 873 5893 876
rect 5636 716 5664 724
rect 5656 696 5664 716
rect 5516 227 5524 433
rect 5576 424 5584 453
rect 5596 447 5604 653
rect 5616 427 5624 633
rect 5636 507 5644 664
rect 5676 587 5684 653
rect 5696 607 5704 713
rect 5716 427 5724 713
rect 5753 700 5767 713
rect 5756 696 5764 700
rect 5796 696 5804 813
rect 5576 416 5604 424
rect 5596 396 5604 416
rect 5556 287 5564 364
rect 5636 247 5644 393
rect 5656 366 5664 413
rect 5736 396 5744 433
rect 5776 407 5784 613
rect 5760 364 5773 367
rect 5756 356 5773 364
rect 5760 353 5773 356
rect 5316 176 5344 184
rect 5296 146 5304 173
rect 5436 167 5444 213
rect 5493 180 5507 193
rect 5496 176 5504 180
rect 5576 146 5584 213
rect 5656 204 5664 352
rect 5636 196 5664 204
rect 5636 176 5644 196
rect 5676 176 5684 293
rect 5796 207 5804 393
rect 5816 366 5824 653
rect 5836 427 5844 773
rect 5856 667 5864 853
rect 5876 707 5884 853
rect 5896 696 5904 753
rect 5916 727 5924 973
rect 5936 887 5944 1613
rect 5876 396 5884 493
rect 5896 407 5904 633
rect 5716 146 5724 193
rect 5816 176 5824 313
rect 5896 307 5904 353
rect 5856 176 5864 233
rect 5916 146 5924 413
rect 5956 327 5964 2693
rect 5976 2446 5984 2773
rect 5976 1807 5984 2293
rect 5976 827 5984 1733
rect 5976 407 5984 453
rect 5836 47 5844 144
rect 956 -24 984 -16
rect 1896 -24 1924 -16
rect 2916 -24 2944 -16
rect 3396 -24 3404 13
rect 3496 -24 3504 13
<< m3contact >>
rect 813 5993 827 6007
rect 913 5993 927 6007
rect 2893 5993 2907 6007
rect 2933 5993 2947 6007
rect 3533 5993 3547 6007
rect 3813 5993 3827 6007
rect 4693 5993 4707 6007
rect 153 5913 167 5927
rect 213 5913 227 5927
rect 113 5894 127 5908
rect 93 5852 107 5866
rect 73 5594 87 5608
rect 132 5594 146 5608
rect 293 5896 307 5910
rect 373 5896 387 5910
rect 533 5896 547 5910
rect 172 5852 186 5866
rect 193 5852 207 5866
rect 233 5852 247 5866
rect 373 5853 387 5867
rect 153 5593 167 5607
rect 53 5553 67 5567
rect 92 5553 106 5567
rect 113 5552 127 5566
rect 153 5553 167 5567
rect 93 5513 107 5527
rect 133 5513 147 5527
rect 53 5493 67 5507
rect 93 5492 107 5506
rect 33 5374 47 5388
rect 13 5113 27 5127
rect 73 5313 87 5327
rect 113 5193 127 5207
rect 53 5073 67 5087
rect 93 5074 107 5088
rect 113 5032 127 5046
rect 93 4993 107 5007
rect 53 4853 67 4867
rect 33 4453 47 4467
rect 33 4413 47 4427
rect 13 4172 27 4186
rect 13 3813 27 3827
rect 13 3773 27 3787
rect 13 3713 27 3727
rect 73 4812 87 4826
rect 113 4812 127 4826
rect 133 4653 147 4667
rect 93 4613 107 4627
rect 193 5593 207 5607
rect 253 5594 267 5608
rect 193 5552 207 5566
rect 293 5553 307 5567
rect 253 5533 267 5547
rect 233 5453 247 5467
rect 213 5374 227 5388
rect 273 5493 287 5507
rect 253 5373 267 5387
rect 173 5313 187 5327
rect 233 5332 247 5346
rect 273 5333 287 5347
rect 233 5113 247 5127
rect 193 5074 207 5088
rect 233 5074 247 5088
rect 213 5032 227 5046
rect 213 4873 227 4887
rect 313 5533 327 5547
rect 473 5833 487 5847
rect 513 5833 527 5847
rect 733 5853 747 5867
rect 713 5833 727 5847
rect 1713 5953 1727 5967
rect 1793 5953 1807 5967
rect 2073 5953 2087 5967
rect 2153 5953 2167 5967
rect 2233 5953 2247 5967
rect 2433 5953 2447 5967
rect 2473 5953 2487 5967
rect 2633 5953 2647 5967
rect 1113 5933 1127 5947
rect 1313 5933 1327 5947
rect 1513 5933 1527 5947
rect 1633 5933 1647 5947
rect 1213 5893 1227 5907
rect 1453 5894 1467 5908
rect 973 5852 987 5866
rect 1533 5893 1547 5907
rect 1593 5894 1607 5908
rect 833 5833 847 5847
rect 913 5833 927 5847
rect 653 5733 667 5747
rect 713 5733 727 5747
rect 653 5693 667 5707
rect 513 5613 527 5627
rect 553 5613 567 5627
rect 433 5596 447 5610
rect 373 5453 387 5467
rect 413 5374 427 5388
rect 313 5313 327 5327
rect 393 5313 407 5327
rect 453 5313 467 5327
rect 293 5193 307 5207
rect 293 5074 307 5088
rect 613 5594 627 5608
rect 833 5613 847 5627
rect 893 5613 907 5627
rect 733 5594 747 5608
rect 793 5594 807 5608
rect 633 5552 647 5566
rect 713 5552 727 5566
rect 673 5533 687 5547
rect 593 5493 607 5507
rect 813 5552 827 5566
rect 573 5413 587 5427
rect 733 5413 747 5427
rect 573 5374 587 5388
rect 633 5376 647 5390
rect 693 5374 707 5388
rect 733 5374 747 5388
rect 553 5313 567 5327
rect 513 5273 527 5287
rect 353 5193 367 5207
rect 553 5113 567 5127
rect 533 5093 547 5107
rect 573 5093 587 5107
rect 393 5074 407 5088
rect 493 5074 507 5088
rect 433 5053 447 5067
rect 293 5033 307 5047
rect 593 5073 607 5087
rect 653 5074 667 5088
rect 573 4993 587 5007
rect 533 4933 547 4947
rect 513 4893 527 4907
rect 433 4873 447 4887
rect 493 4873 507 4887
rect 373 4854 387 4868
rect 413 4853 427 4867
rect 233 4812 247 4826
rect 293 4653 307 4667
rect 313 4613 327 4627
rect 293 4573 307 4587
rect 193 4554 207 4568
rect 253 4554 267 4568
rect 153 4512 167 4526
rect 193 4513 207 4527
rect 113 4373 127 4387
rect 133 4334 147 4348
rect 193 4453 207 4467
rect 173 4373 187 4387
rect 153 4333 167 4347
rect 113 4253 127 4267
rect 153 4193 167 4207
rect 93 4133 107 4147
rect 213 4373 227 4387
rect 173 4033 187 4047
rect 93 3973 107 3987
rect 173 3993 187 4007
rect 113 3933 127 3947
rect 133 3933 147 3947
rect 93 3814 107 3828
rect 153 3853 167 3867
rect 53 3733 67 3747
rect 33 3613 47 3627
rect 233 4292 247 4306
rect 213 4233 227 4247
rect 293 4493 307 4507
rect 353 4653 367 4667
rect 573 4893 587 4907
rect 473 4793 487 4807
rect 433 4613 447 4627
rect 513 4613 527 4627
rect 353 4573 367 4587
rect 333 4453 347 4467
rect 413 4573 427 4587
rect 393 4553 407 4567
rect 493 4553 507 4567
rect 393 4513 407 4527
rect 373 4473 387 4487
rect 373 4413 387 4427
rect 353 4373 367 4387
rect 333 4334 347 4348
rect 453 4513 467 4527
rect 433 4473 447 4487
rect 393 4373 407 4387
rect 293 4292 307 4306
rect 353 4292 367 4306
rect 393 4273 407 4287
rect 273 4153 287 4167
rect 213 3993 227 4007
rect 193 3953 207 3967
rect 193 3853 207 3867
rect 293 3853 307 3867
rect 173 3593 187 3607
rect 113 3533 127 3547
rect 93 3514 107 3528
rect 133 3514 147 3528
rect 173 3514 187 3528
rect 73 3472 87 3486
rect 173 3433 187 3447
rect 253 3814 267 3828
rect 373 3953 387 3967
rect 333 3933 347 3947
rect 313 3813 327 3827
rect 313 3792 327 3806
rect 233 3772 247 3786
rect 273 3772 287 3786
rect 433 4292 447 4306
rect 473 4453 487 4467
rect 753 5332 767 5346
rect 893 5493 907 5507
rect 853 5473 867 5487
rect 1013 5693 1027 5707
rect 993 5653 1007 5667
rect 953 5594 967 5608
rect 1433 5852 1447 5866
rect 1333 5813 1347 5827
rect 1153 5773 1167 5787
rect 1293 5773 1307 5787
rect 1073 5673 1087 5687
rect 1133 5673 1147 5687
rect 1013 5633 1027 5647
rect 973 5533 987 5547
rect 993 5513 1007 5527
rect 913 5453 927 5467
rect 973 5453 987 5467
rect 853 5413 867 5427
rect 853 5374 867 5388
rect 893 5374 907 5388
rect 953 5374 967 5388
rect 873 5332 887 5346
rect 853 5293 867 5307
rect 793 5193 807 5207
rect 733 5113 747 5127
rect 633 5032 647 5046
rect 633 4933 647 4947
rect 713 5033 727 5047
rect 793 5074 807 5088
rect 773 5032 787 5046
rect 813 4993 827 5007
rect 913 5293 927 5307
rect 1053 5393 1067 5407
rect 1113 5594 1127 5608
rect 1513 5852 1527 5866
rect 1533 5813 1547 5827
rect 1613 5813 1627 5827
rect 1513 5773 1527 5787
rect 1573 5773 1587 5787
rect 1473 5693 1487 5707
rect 1493 5673 1507 5687
rect 1493 5633 1507 5647
rect 1293 5594 1307 5608
rect 1333 5594 1347 5608
rect 1413 5594 1427 5608
rect 1453 5594 1467 5608
rect 1233 5573 1247 5587
rect 1373 5573 1387 5587
rect 1233 5513 1247 5527
rect 1133 5493 1147 5507
rect 1313 5552 1327 5566
rect 1653 5693 1667 5707
rect 1533 5594 1547 5608
rect 1573 5594 1587 5608
rect 1613 5594 1627 5608
rect 1673 5594 1687 5608
rect 1433 5552 1447 5566
rect 1473 5552 1487 5566
rect 1513 5553 1527 5567
rect 1533 5533 1547 5547
rect 1373 5513 1387 5527
rect 1433 5513 1447 5527
rect 1273 5473 1287 5487
rect 1233 5393 1247 5407
rect 993 5333 1007 5347
rect 1033 5332 1047 5346
rect 973 5293 987 5307
rect 953 5273 967 5287
rect 1113 5373 1127 5387
rect 1173 5374 1187 5388
rect 1133 5293 1147 5307
rect 1113 5133 1127 5147
rect 1013 5113 1027 5127
rect 1093 5113 1107 5127
rect 933 5074 947 5088
rect 993 5073 1007 5087
rect 873 5033 887 5047
rect 913 5032 927 5046
rect 953 5032 967 5046
rect 853 4973 867 4987
rect 953 4973 967 4987
rect 653 4913 667 4927
rect 673 4913 687 4927
rect 693 4856 707 4870
rect 633 4793 647 4807
rect 773 4893 787 4907
rect 913 4856 927 4870
rect 773 4813 787 4827
rect 813 4810 827 4824
rect 753 4773 767 4787
rect 813 4773 827 4787
rect 873 4773 887 4787
rect 593 4593 607 4607
rect 693 4593 707 4607
rect 533 4513 547 4527
rect 593 4554 607 4568
rect 653 4554 667 4568
rect 633 4493 647 4507
rect 513 4352 527 4366
rect 733 4554 747 4568
rect 773 4554 787 4568
rect 793 4513 807 4527
rect 753 4473 767 4487
rect 713 4393 727 4407
rect 773 4393 787 4407
rect 693 4353 707 4367
rect 553 4333 567 4347
rect 473 4273 487 4287
rect 453 4233 467 4247
rect 573 4153 587 4167
rect 533 4093 547 4107
rect 573 4092 587 4106
rect 413 4053 427 4067
rect 393 3893 407 3907
rect 493 3933 507 3947
rect 533 3913 547 3927
rect 353 3833 367 3847
rect 413 3834 427 3848
rect 333 3772 347 3786
rect 253 3693 267 3707
rect 313 3693 327 3707
rect 213 3633 227 3647
rect 413 3813 427 3827
rect 453 3814 467 3828
rect 573 3913 587 3927
rect 553 3873 567 3887
rect 573 3853 587 3867
rect 613 4334 627 4348
rect 673 4334 687 4348
rect 753 4353 767 4367
rect 693 4292 707 4306
rect 653 4253 667 4267
rect 633 4193 647 4207
rect 613 4133 627 4147
rect 633 4113 647 4127
rect 613 4033 627 4047
rect 673 4034 687 4048
rect 733 4034 747 4048
rect 653 3992 667 4006
rect 693 3992 707 4006
rect 693 3953 707 3967
rect 673 3873 687 3887
rect 653 3853 667 3867
rect 593 3833 607 3847
rect 633 3833 647 3847
rect 373 3772 387 3786
rect 433 3772 447 3786
rect 373 3733 387 3747
rect 373 3712 387 3726
rect 373 3673 387 3687
rect 353 3652 367 3666
rect 553 3613 567 3627
rect 513 3593 527 3607
rect 593 3573 607 3587
rect 633 3753 647 3767
rect 613 3553 627 3567
rect 733 3933 747 3947
rect 713 3873 727 3887
rect 693 3813 707 3827
rect 873 4713 887 4727
rect 913 4713 927 4727
rect 833 4554 847 4568
rect 873 4554 887 4568
rect 913 4554 927 4568
rect 893 4512 907 4526
rect 833 4493 847 4507
rect 853 4353 867 4367
rect 893 4353 907 4367
rect 813 4333 827 4347
rect 833 4233 847 4247
rect 973 4933 987 4947
rect 1073 5074 1087 5088
rect 1113 5074 1127 5088
rect 1113 5033 1127 5047
rect 1193 5332 1207 5346
rect 1153 5253 1167 5267
rect 1313 5374 1327 5388
rect 1393 5373 1407 5387
rect 1433 5374 1447 5388
rect 1473 5374 1487 5388
rect 1293 5293 1307 5307
rect 1233 5253 1247 5267
rect 1313 5253 1327 5267
rect 1233 5133 1247 5147
rect 1193 5074 1207 5088
rect 1293 5113 1307 5127
rect 1053 4993 1067 5007
rect 1013 4933 1027 4947
rect 993 4913 1007 4927
rect 993 4892 1007 4906
rect 973 4853 987 4867
rect 1053 4854 1067 4868
rect 1033 4812 1047 4826
rect 1053 4793 1067 4807
rect 1033 4753 1047 4767
rect 1173 5032 1187 5046
rect 1173 4993 1187 5007
rect 1633 5552 1647 5566
rect 1593 5533 1607 5547
rect 1553 5413 1567 5427
rect 1613 5374 1627 5388
rect 1693 5553 1707 5567
rect 1753 5894 1767 5908
rect 1933 5894 1947 5908
rect 2033 5894 2047 5908
rect 2113 5933 2127 5947
rect 2113 5893 2127 5907
rect 1813 5852 1827 5866
rect 1773 5733 1787 5747
rect 1973 5852 1987 5866
rect 2053 5852 2067 5866
rect 2093 5852 2107 5866
rect 1793 5633 1807 5647
rect 1912 5633 1926 5647
rect 1933 5633 1947 5647
rect 1873 5594 1887 5608
rect 2013 5773 2027 5787
rect 1973 5594 1987 5608
rect 1693 5374 1707 5388
rect 1813 5552 1827 5566
rect 1773 5513 1787 5527
rect 1793 5374 1807 5388
rect 2213 5913 2227 5927
rect 2453 5933 2467 5947
rect 2253 5913 2267 5927
rect 2233 5893 2247 5907
rect 2193 5852 2207 5866
rect 2153 5773 2167 5787
rect 2173 5733 2187 5747
rect 2093 5633 2107 5647
rect 2133 5633 2147 5647
rect 2093 5612 2107 5626
rect 2053 5594 2067 5608
rect 2153 5613 2167 5627
rect 2133 5593 2147 5607
rect 1913 5552 1927 5566
rect 1953 5552 1967 5566
rect 2013 5552 2027 5566
rect 2073 5552 2087 5566
rect 2113 5493 2127 5507
rect 1913 5473 1927 5487
rect 1973 5473 1987 5487
rect 1653 5293 1667 5307
rect 1753 5332 1767 5346
rect 1753 5293 1767 5307
rect 1713 5253 1727 5267
rect 1433 5113 1447 5127
rect 1333 5073 1347 5087
rect 1393 5074 1407 5088
rect 1313 5033 1327 5047
rect 1253 4953 1267 4967
rect 1213 4873 1227 4887
rect 1213 4810 1227 4824
rect 1373 5032 1387 5046
rect 1413 4973 1427 4987
rect 1393 4953 1407 4967
rect 1333 4854 1347 4868
rect 2033 5393 2047 5407
rect 2033 5374 2047 5388
rect 2073 5374 2087 5388
rect 2233 5613 2247 5627
rect 2273 5893 2287 5907
rect 2313 5894 2327 5908
rect 2353 5894 2367 5908
rect 2393 5894 2407 5908
rect 2493 5894 2507 5908
rect 2273 5813 2287 5827
rect 2353 5793 2367 5807
rect 2333 5673 2347 5687
rect 2333 5613 2347 5627
rect 2273 5594 2287 5608
rect 2173 5553 2187 5567
rect 2253 5552 2267 5566
rect 2293 5552 2307 5566
rect 2593 5893 2607 5907
rect 2673 5894 2687 5908
rect 2733 5894 2747 5908
rect 2773 5894 2787 5908
rect 2473 5793 2487 5807
rect 2593 5852 2607 5866
rect 2653 5833 2667 5847
rect 2713 5833 2727 5847
rect 2693 5793 2707 5807
rect 2793 5833 2807 5847
rect 2733 5793 2747 5807
rect 2513 5773 2527 5787
rect 2713 5773 2727 5787
rect 2393 5733 2407 5747
rect 2453 5633 2467 5647
rect 2353 5553 2367 5567
rect 2393 5552 2407 5566
rect 2293 5433 2307 5447
rect 2193 5393 2207 5407
rect 2153 5373 2167 5387
rect 2233 5374 2247 5388
rect 2293 5374 2307 5388
rect 1933 5332 1947 5346
rect 1973 5332 1987 5346
rect 2013 5332 2027 5346
rect 1833 5253 1847 5267
rect 1593 5113 1607 5127
rect 1793 5113 1807 5127
rect 1553 5074 1567 5088
rect 1633 5074 1647 5088
rect 1733 5074 1747 5088
rect 1773 5074 1787 5088
rect 1813 5074 1827 5088
rect 1573 5032 1587 5046
rect 1653 5053 1667 5067
rect 1493 4973 1507 4987
rect 1533 4973 1547 4987
rect 1633 4973 1647 4987
rect 1473 4913 1487 4927
rect 1433 4854 1447 4868
rect 1573 4913 1587 4927
rect 1613 4854 1627 4868
rect 1273 4773 1287 4787
rect 1313 4773 1327 4787
rect 1413 4773 1427 4787
rect 1173 4753 1187 4767
rect 1053 4553 1067 4567
rect 1113 4554 1127 4568
rect 993 4513 1007 4527
rect 1113 4513 1127 4527
rect 1073 4413 1087 4427
rect 973 4373 987 4387
rect 1113 4334 1127 4348
rect 973 4293 987 4307
rect 1013 4290 1027 4304
rect 1073 4290 1087 4304
rect 1073 4253 1087 4267
rect 913 4193 927 4207
rect 953 4193 967 4207
rect 853 4173 867 4187
rect 773 4133 787 4147
rect 833 4133 847 4147
rect 793 4034 807 4048
rect 853 4093 867 4107
rect 813 3992 827 4006
rect 893 3993 907 4007
rect 1593 4812 1607 4826
rect 1713 5032 1727 5046
rect 1793 5033 1807 5047
rect 1753 4993 1767 5007
rect 1733 4973 1747 4987
rect 1793 4973 1807 4987
rect 1693 4854 1707 4868
rect 1793 4893 1807 4907
rect 1713 4812 1727 4826
rect 1753 4812 1767 4826
rect 1573 4773 1587 4787
rect 1653 4773 1667 4787
rect 1353 4593 1367 4607
rect 1173 4554 1187 4568
rect 1253 4553 1267 4567
rect 1253 4493 1267 4507
rect 1193 4453 1207 4467
rect 1273 4413 1287 4427
rect 1213 4373 1227 4387
rect 1173 4334 1187 4348
rect 1173 4233 1187 4247
rect 1173 4193 1187 4207
rect 1133 4173 1147 4187
rect 1093 4133 1107 4147
rect 973 4113 987 4127
rect 1053 4113 1067 4127
rect 1033 4073 1047 4087
rect 853 3853 867 3867
rect 733 3772 747 3786
rect 673 3753 687 3767
rect 653 3613 667 3627
rect 873 3772 887 3786
rect 833 3753 847 3767
rect 773 3653 787 3667
rect 753 3613 767 3627
rect 733 3573 747 3587
rect 733 3552 747 3566
rect 513 3513 527 3527
rect 593 3513 607 3527
rect 633 3513 647 3527
rect 673 3513 687 3527
rect 493 3492 507 3506
rect 273 3472 287 3486
rect 533 3470 547 3484
rect 493 3452 507 3466
rect 333 3433 347 3447
rect 193 3373 207 3387
rect 253 3373 267 3387
rect 213 3296 227 3310
rect 93 3250 107 3264
rect 133 3250 147 3264
rect 33 3233 47 3247
rect 93 3193 107 3207
rect 33 3033 47 3047
rect 153 3033 167 3047
rect 72 2993 86 3007
rect 93 2996 107 3010
rect 133 2996 147 3010
rect 133 2893 147 2907
rect 133 2813 147 2827
rect 93 2730 107 2744
rect 133 2730 147 2744
rect 213 2950 227 2964
rect 213 2776 227 2790
rect 273 3296 287 3310
rect 413 3413 427 3427
rect 273 3253 287 3267
rect 273 2950 287 2964
rect 313 3252 327 3266
rect 353 3252 367 3266
rect 373 3013 387 3027
rect 333 2994 347 3008
rect 473 3433 487 3447
rect 493 3413 507 3427
rect 553 3296 567 3310
rect 833 3573 847 3587
rect 913 3573 927 3587
rect 773 3513 787 3527
rect 813 3472 827 3486
rect 913 3473 927 3487
rect 993 3992 1007 4006
rect 1033 3992 1047 4006
rect 1013 3933 1027 3947
rect 973 3853 987 3867
rect 953 3813 967 3827
rect 1093 4053 1107 4067
rect 1073 3993 1087 4007
rect 1053 3813 1067 3827
rect 993 3753 1007 3767
rect 1133 3992 1147 4006
rect 1173 3993 1187 4007
rect 1113 3833 1127 3847
rect 1173 3833 1187 3847
rect 1093 3813 1107 3827
rect 1073 3753 1087 3767
rect 1233 4253 1247 4267
rect 1333 4493 1347 4507
rect 1373 4413 1387 4427
rect 1553 4613 1567 4627
rect 1533 4593 1547 4607
rect 1433 4554 1447 4568
rect 1473 4554 1487 4568
rect 1413 4513 1427 4527
rect 1393 4333 1407 4347
rect 1353 4292 1367 4306
rect 1293 4253 1307 4267
rect 1273 4193 1287 4207
rect 1233 4113 1247 4127
rect 1253 4073 1267 4087
rect 1233 4053 1247 4067
rect 1313 4053 1327 4067
rect 1373 4036 1387 4050
rect 1213 3873 1227 3887
rect 1193 3813 1207 3827
rect 1153 3772 1167 3786
rect 1393 3992 1407 4006
rect 1493 4512 1507 4526
rect 1473 4493 1487 4507
rect 1453 4433 1467 4447
rect 1433 4393 1447 4407
rect 1533 4433 1547 4447
rect 1473 4373 1487 4387
rect 1433 4332 1447 4346
rect 1493 4334 1507 4348
rect 1533 4334 1547 4348
rect 1653 4633 1667 4647
rect 1613 4554 1627 4568
rect 1713 4554 1727 4568
rect 1573 4513 1587 4527
rect 1633 4512 1647 4526
rect 1673 4453 1687 4467
rect 1753 4553 1767 4567
rect 2093 5293 2107 5307
rect 2213 5293 2227 5307
rect 2053 5153 2067 5167
rect 1893 5074 1907 5088
rect 1973 5074 1987 5088
rect 2053 5074 2067 5088
rect 2173 5233 2187 5247
rect 2113 5153 2127 5167
rect 1833 5033 1847 5047
rect 1873 5032 1887 5046
rect 1913 5032 1927 5046
rect 2093 5073 2107 5087
rect 2033 5032 2047 5046
rect 2073 5032 2087 5046
rect 1973 4993 1987 5007
rect 1913 4973 1927 4987
rect 1833 4933 1847 4947
rect 1813 4813 1827 4827
rect 1873 4854 1887 4868
rect 1913 4854 1927 4868
rect 2133 5093 2147 5107
rect 2113 4973 2127 4987
rect 2073 4854 2087 4868
rect 1933 4812 1947 4826
rect 2053 4812 2067 4826
rect 1893 4793 1907 4807
rect 2093 4812 2107 4826
rect 2293 5333 2307 5347
rect 2473 5552 2487 5566
rect 2433 5453 2447 5467
rect 2373 5374 2387 5388
rect 2353 5332 2367 5346
rect 2313 5273 2327 5287
rect 2413 5233 2427 5247
rect 2273 5213 2287 5227
rect 2253 5193 2267 5207
rect 2393 5133 2407 5147
rect 2193 4893 2207 4907
rect 2233 4893 2247 4907
rect 2193 4812 2207 4826
rect 2093 4793 2107 4807
rect 1933 4713 1947 4727
rect 1833 4613 1847 4627
rect 1833 4554 1847 4568
rect 1893 4554 1907 4568
rect 2233 4773 2247 4787
rect 2293 5073 2307 5087
rect 2333 5074 2347 5088
rect 2353 5032 2367 5046
rect 2393 5032 2407 5046
rect 2353 4973 2367 4987
rect 2313 4854 2327 4868
rect 2393 4854 2407 4868
rect 2293 4812 2307 4826
rect 2333 4812 2347 4826
rect 2253 4713 2267 4727
rect 2373 4673 2387 4687
rect 2193 4653 2207 4667
rect 2153 4633 2167 4647
rect 2073 4613 2087 4627
rect 1973 4554 1987 4568
rect 2013 4554 2027 4568
rect 1813 4512 1827 4526
rect 1873 4512 1887 4526
rect 1733 4493 1747 4507
rect 1773 4493 1787 4507
rect 1713 4433 1727 4447
rect 1833 4393 1847 4407
rect 1873 4393 1887 4407
rect 1593 4353 1607 4367
rect 1673 4353 1687 4367
rect 1513 4292 1527 4306
rect 1473 4133 1487 4147
rect 1553 4133 1567 4147
rect 1433 4073 1447 4087
rect 1533 4073 1547 4087
rect 1433 4036 1447 4050
rect 1433 3993 1447 4007
rect 1413 3973 1427 3987
rect 1273 3873 1287 3887
rect 1333 3873 1347 3887
rect 1273 3833 1287 3847
rect 1233 3813 1247 3827
rect 1293 3772 1307 3786
rect 1173 3753 1187 3767
rect 1093 3653 1107 3667
rect 1513 3953 1527 3967
rect 1433 3913 1447 3927
rect 1533 3913 1547 3927
rect 1413 3693 1427 3707
rect 1193 3653 1207 3667
rect 1253 3653 1267 3667
rect 1313 3653 1327 3667
rect 1173 3613 1187 3627
rect 973 3593 987 3607
rect 1293 3573 1307 3587
rect 1193 3553 1207 3567
rect 1253 3553 1267 3567
rect 973 3514 987 3528
rect 1013 3514 1027 3528
rect 1132 3514 1146 3528
rect 993 3472 1007 3486
rect 773 3433 787 3447
rect 853 3433 867 3447
rect 933 3433 947 3447
rect 1153 3513 1167 3527
rect 1193 3516 1207 3530
rect 1133 3373 1147 3387
rect 1193 3433 1207 3447
rect 1153 3353 1167 3367
rect 793 3333 807 3347
rect 1053 3333 1067 3347
rect 1133 3333 1147 3347
rect 773 3313 787 3327
rect 633 3293 647 3307
rect 753 3293 767 3307
rect 613 3273 627 3287
rect 473 3252 487 3266
rect 513 3252 527 3266
rect 433 3013 447 3027
rect 633 3250 647 3264
rect 673 3250 687 3264
rect 733 3233 747 3247
rect 513 3013 527 3027
rect 573 3013 587 3027
rect 333 2933 347 2947
rect 393 2952 407 2966
rect 353 2893 367 2907
rect 273 2733 287 2747
rect 453 2993 467 3007
rect 493 2994 507 3008
rect 453 2952 467 2966
rect 533 2933 547 2947
rect 493 2813 507 2827
rect 553 2813 567 2827
rect 33 2693 47 2707
rect 153 2693 167 2707
rect 253 2693 267 2707
rect 253 2633 267 2647
rect 33 2493 47 2507
rect 153 2493 167 2507
rect 93 2476 107 2490
rect 133 2476 147 2490
rect 133 2373 147 2387
rect 213 2413 227 2427
rect 253 2393 267 2407
rect 33 2210 47 2224
rect 153 2213 167 2227
rect 273 2273 287 2287
rect 313 2732 327 2746
rect 353 2732 367 2746
rect 392 2732 406 2746
rect 413 2732 427 2746
rect 473 2732 487 2746
rect 513 2732 527 2746
rect 553 2732 567 2746
rect 373 2693 387 2707
rect 333 2474 347 2488
rect 433 2693 447 2707
rect 393 2673 407 2687
rect 333 2413 347 2427
rect 393 2432 407 2446
rect 353 2373 367 2387
rect 253 2193 267 2207
rect 93 2173 107 2187
rect 893 3313 907 3327
rect 853 3294 867 3308
rect 953 3293 967 3307
rect 993 3294 1007 3308
rect 1033 3294 1047 3308
rect 1073 3293 1087 3307
rect 873 3252 887 3266
rect 913 3053 927 3067
rect 1413 3613 1427 3627
rect 1373 3553 1387 3567
rect 1313 3472 1327 3486
rect 1353 3472 1367 3486
rect 1353 3433 1367 3447
rect 1413 3433 1427 3447
rect 1293 3413 1307 3427
rect 1233 3353 1247 3367
rect 1293 3353 1307 3367
rect 1213 3293 1227 3307
rect 1013 3252 1027 3266
rect 1073 3252 1087 3266
rect 1153 3252 1167 3266
rect 1173 3133 1187 3147
rect 973 3053 987 3067
rect 953 2994 967 3008
rect 933 2952 947 2966
rect 653 2873 667 2887
rect 753 2913 767 2927
rect 873 2912 887 2926
rect 1033 3033 1047 3047
rect 1033 2994 1047 3008
rect 1013 2953 1027 2967
rect 973 2873 987 2887
rect 673 2833 687 2847
rect 733 2833 747 2847
rect 713 2813 727 2827
rect 593 2793 607 2807
rect 693 2793 707 2807
rect 613 2773 627 2787
rect 653 2774 667 2788
rect 993 2813 1007 2827
rect 753 2753 767 2767
rect 593 2713 607 2727
rect 673 2732 687 2746
rect 733 2732 747 2746
rect 1053 2952 1067 2966
rect 1133 2933 1147 2947
rect 1013 2776 1027 2790
rect 1073 2776 1087 2790
rect 633 2713 647 2727
rect 753 2713 767 2727
rect 793 2713 807 2727
rect 613 2693 627 2707
rect 593 2593 607 2607
rect 473 2573 487 2587
rect 573 2573 587 2587
rect 453 2513 467 2527
rect 533 2513 547 2527
rect 493 2474 507 2488
rect 693 2593 707 2607
rect 653 2533 667 2547
rect 633 2473 647 2487
rect 453 2433 467 2447
rect 433 2373 447 2387
rect 353 2212 367 2226
rect 393 2212 407 2226
rect 313 2193 327 2207
rect 273 2113 287 2127
rect 13 2033 27 2047
rect 93 2033 107 2047
rect 193 2033 207 2047
rect 233 2033 247 2047
rect 133 1693 147 1707
rect 93 1513 107 1527
rect 33 1473 47 1487
rect 93 1473 107 1487
rect 93 1436 107 1450
rect 113 1393 127 1407
rect 53 1313 67 1327
rect 193 1692 207 1706
rect 233 1692 247 1706
rect 153 1533 167 1547
rect 133 1313 147 1327
rect 213 1390 227 1404
rect 233 1353 247 1367
rect 433 2153 447 2167
rect 353 1954 367 1968
rect 553 2433 567 2447
rect 513 2373 527 2387
rect 513 2273 527 2287
rect 573 2430 587 2444
rect 753 2493 767 2507
rect 693 2254 707 2268
rect 773 2253 787 2267
rect 493 2212 507 2226
rect 493 2173 507 2187
rect 533 2173 547 2187
rect 513 2133 527 2147
rect 493 2093 507 2107
rect 473 1993 487 2007
rect 313 1933 327 1947
rect 373 1912 387 1926
rect 293 1893 307 1907
rect 293 1673 307 1687
rect 413 1893 427 1907
rect 413 1793 427 1807
rect 373 1734 387 1748
rect 333 1693 347 1707
rect 393 1673 407 1687
rect 353 1573 367 1587
rect 433 1573 447 1587
rect 333 1453 347 1467
rect 373 1453 387 1467
rect 293 1390 307 1404
rect 273 1313 287 1327
rect 193 1293 207 1307
rect 233 1293 247 1307
rect 153 1273 167 1287
rect 93 1172 107 1186
rect 53 953 67 967
rect 133 933 147 947
rect 53 913 67 927
rect 93 914 107 928
rect 33 593 47 607
rect 253 1214 267 1228
rect 393 1392 407 1406
rect 513 2053 527 2067
rect 633 2212 647 2226
rect 573 2153 587 2167
rect 613 2153 627 2167
rect 553 2113 567 2127
rect 553 2033 567 2047
rect 573 1993 587 2007
rect 533 1954 547 1968
rect 713 2212 727 2226
rect 673 2053 687 2067
rect 733 2053 747 2067
rect 713 1953 727 1967
rect 513 1893 527 1907
rect 593 1912 607 1926
rect 653 1910 667 1924
rect 673 1793 687 1807
rect 493 1734 507 1748
rect 573 1734 587 1748
rect 773 2212 787 2226
rect 953 2730 967 2744
rect 993 2733 1007 2747
rect 1093 2732 1107 2746
rect 853 2713 867 2727
rect 893 2713 907 2727
rect 833 2673 847 2687
rect 833 2652 847 2666
rect 813 2473 827 2487
rect 953 2513 967 2527
rect 853 2493 867 2507
rect 873 2474 887 2488
rect 833 2393 847 2407
rect 933 2393 947 2407
rect 813 2313 827 2327
rect 893 2313 907 2327
rect 813 2273 827 2287
rect 853 2254 867 2268
rect 833 2212 847 2226
rect 873 2212 887 2226
rect 833 2113 847 2127
rect 933 2093 947 2107
rect 793 2053 807 2067
rect 833 2053 847 2067
rect 973 2473 987 2487
rect 1033 2474 1047 2488
rect 1053 2413 1067 2427
rect 1013 2373 1027 2387
rect 973 2273 987 2287
rect 1073 2273 1087 2287
rect 1013 2254 1027 2268
rect 993 2193 1007 2207
rect 993 2153 1007 2167
rect 853 2013 867 2027
rect 953 2013 967 2027
rect 893 1973 907 1987
rect 953 1956 967 1970
rect 1333 3293 1347 3307
rect 1233 3213 1247 3227
rect 1233 2994 1247 3008
rect 1153 2913 1167 2927
rect 1213 2913 1227 2927
rect 1133 2653 1147 2667
rect 1273 3252 1287 3266
rect 1633 4334 1647 4348
rect 1793 4353 1807 4367
rect 1593 4253 1607 4267
rect 1693 4292 1707 4306
rect 1813 4292 1827 4306
rect 1653 4213 1667 4227
rect 1773 4213 1787 4227
rect 1733 4173 1747 4187
rect 1573 4053 1587 4067
rect 1653 4053 1667 4067
rect 1633 3992 1647 4006
rect 1673 3973 1687 3987
rect 1713 3973 1727 3987
rect 1593 3953 1607 3967
rect 1573 3913 1587 3927
rect 1653 3913 1667 3927
rect 1593 3773 1607 3787
rect 1633 3772 1647 3786
rect 1573 3753 1587 3767
rect 1533 3733 1547 3747
rect 1613 3693 1627 3707
rect 1573 3593 1587 3607
rect 1493 3553 1507 3567
rect 1473 3533 1487 3547
rect 1533 3533 1547 3547
rect 1573 3533 1587 3547
rect 1513 3472 1527 3486
rect 1473 3433 1487 3447
rect 1533 3413 1547 3427
rect 1453 3353 1467 3367
rect 1513 3353 1527 3367
rect 1393 3333 1407 3347
rect 1433 3333 1447 3347
rect 1373 3313 1387 3327
rect 1353 3233 1367 3247
rect 1413 3293 1427 3307
rect 1513 3293 1527 3307
rect 1393 3252 1407 3266
rect 1492 3252 1506 3266
rect 1513 3252 1527 3266
rect 1433 3213 1447 3227
rect 1313 3173 1327 3187
rect 1373 3173 1387 3187
rect 1313 3133 1327 3147
rect 1393 3053 1407 3067
rect 1473 3053 1487 3067
rect 1333 3033 1347 3047
rect 1293 2994 1307 3008
rect 1253 2913 1267 2927
rect 1233 2893 1247 2907
rect 1213 2873 1227 2887
rect 1353 2952 1367 2966
rect 1433 3013 1447 3027
rect 1433 2994 1447 3008
rect 1593 3513 1607 3527
rect 1673 3653 1687 3667
rect 1933 4493 1947 4507
rect 1913 4353 1927 4367
rect 1913 4292 1927 4306
rect 1893 4133 1907 4147
rect 2113 4554 2127 4568
rect 2033 4513 2047 4527
rect 2093 4512 2107 4526
rect 2013 4493 2027 4507
rect 1953 4453 1967 4467
rect 2093 4453 2107 4467
rect 2033 4433 2047 4447
rect 1993 4353 2007 4367
rect 1953 4333 1967 4347
rect 2173 4613 2187 4627
rect 2153 4433 2167 4447
rect 2213 4613 2227 4627
rect 2193 4573 2207 4587
rect 2573 5633 2587 5647
rect 2633 5633 2647 5647
rect 2513 5593 2527 5607
rect 2553 5552 2567 5566
rect 2593 5552 2607 5566
rect 2653 5613 2667 5627
rect 2753 5613 2767 5627
rect 2713 5594 2727 5608
rect 2673 5553 2687 5567
rect 2653 5533 2667 5547
rect 2633 5513 2647 5527
rect 2653 5473 2667 5487
rect 2493 5453 2507 5467
rect 2593 5453 2607 5467
rect 2513 5433 2527 5447
rect 2573 5374 2587 5388
rect 2493 5293 2507 5307
rect 2493 5173 2507 5187
rect 2553 5173 2567 5187
rect 2493 5133 2507 5147
rect 2453 5093 2467 5107
rect 2433 5073 2447 5087
rect 2473 5032 2487 5046
rect 2493 4993 2507 5007
rect 2453 4854 2467 4868
rect 2513 4893 2527 4907
rect 2473 4812 2487 4826
rect 2513 4773 2527 4787
rect 2673 5453 2687 5467
rect 2713 5533 2727 5547
rect 2733 5513 2747 5527
rect 2693 5374 2707 5388
rect 2593 5333 2607 5347
rect 2673 5332 2687 5346
rect 2593 5273 2607 5287
rect 2573 5133 2587 5147
rect 2813 5793 2827 5807
rect 2753 5453 2767 5467
rect 2793 5453 2807 5467
rect 2773 5413 2787 5427
rect 2773 5373 2787 5387
rect 3753 5953 3767 5967
rect 3273 5933 3287 5947
rect 3613 5933 3627 5947
rect 2933 5894 2947 5908
rect 2973 5894 2987 5908
rect 3033 5894 3047 5908
rect 3093 5894 3107 5908
rect 3133 5894 3147 5908
rect 2953 5852 2967 5866
rect 2993 5852 3007 5866
rect 2893 5833 2907 5847
rect 3172 5893 3186 5907
rect 3193 5894 3207 5908
rect 3233 5894 3247 5908
rect 3073 5852 3087 5866
rect 2852 5693 2866 5707
rect 2873 5693 2887 5707
rect 2933 5693 2947 5707
rect 2893 5633 2907 5647
rect 2853 5593 2867 5607
rect 2973 5594 2987 5608
rect 2873 5552 2887 5566
rect 2913 5552 2927 5566
rect 2953 5552 2967 5566
rect 2933 5513 2947 5527
rect 2873 5453 2887 5467
rect 2793 5332 2807 5346
rect 2753 5273 2767 5287
rect 2813 5273 2827 5287
rect 2773 5213 2787 5227
rect 2693 5193 2707 5207
rect 2733 5193 2747 5207
rect 2673 5173 2687 5187
rect 2653 5032 2667 5046
rect 2693 5033 2707 5047
rect 2593 4893 2607 4907
rect 2573 4854 2587 4868
rect 2613 4854 2627 4868
rect 2653 4854 2667 4868
rect 2573 4773 2587 4787
rect 2553 4753 2567 4767
rect 2633 4773 2647 4787
rect 2473 4733 2487 4747
rect 2613 4733 2627 4747
rect 2493 4633 2507 4647
rect 2593 4633 2607 4647
rect 2413 4613 2427 4627
rect 2273 4554 2287 4568
rect 2333 4553 2347 4567
rect 2373 4554 2387 4568
rect 2513 4593 2527 4607
rect 2553 4593 2567 4607
rect 2453 4573 2467 4587
rect 2493 4573 2507 4587
rect 2313 4533 2327 4547
rect 2233 4512 2247 4526
rect 2193 4433 2207 4447
rect 2173 4413 2187 4427
rect 2053 4393 2067 4407
rect 2093 4393 2107 4407
rect 2073 4373 2087 4387
rect 2133 4373 2147 4387
rect 1973 4292 1987 4306
rect 2053 4293 2067 4307
rect 2013 4233 2027 4247
rect 1973 4213 1987 4227
rect 1893 4093 1907 4107
rect 1933 4093 1947 4107
rect 1793 3953 1807 3967
rect 1793 3893 1807 3907
rect 1953 3953 1967 3967
rect 2113 4334 2127 4348
rect 2153 4334 2167 4348
rect 2073 4233 2087 4247
rect 2133 4233 2147 4247
rect 2273 4393 2287 4407
rect 2193 4213 2207 4227
rect 2153 4053 2167 4067
rect 2113 4034 2127 4048
rect 2293 4273 2307 4287
rect 2393 4512 2407 4526
rect 2393 4473 2407 4487
rect 2373 4453 2387 4467
rect 2353 4293 2367 4307
rect 2433 4453 2447 4467
rect 2513 4512 2527 4526
rect 2573 4512 2587 4526
rect 2653 4653 2667 4667
rect 2753 5032 2767 5046
rect 2773 4973 2787 4987
rect 2773 4854 2787 4868
rect 2833 5193 2847 5207
rect 2833 5133 2847 5147
rect 2833 5074 2847 5088
rect 2893 5374 2907 5388
rect 3173 5852 3187 5866
rect 3093 5673 3107 5687
rect 3053 5594 3067 5608
rect 3333 5893 3347 5907
rect 3393 5894 3407 5908
rect 3473 5893 3487 5907
rect 3533 5894 3547 5908
rect 3573 5894 3587 5908
rect 3253 5852 3267 5866
rect 3413 5852 3427 5866
rect 3293 5833 3307 5847
rect 3333 5833 3347 5847
rect 3193 5793 3207 5807
rect 3633 5893 3647 5907
rect 3473 5773 3487 5787
rect 3133 5633 3147 5647
rect 3233 5633 3247 5647
rect 3353 5633 3367 5647
rect 3433 5633 3447 5647
rect 3113 5594 3127 5608
rect 3193 5594 3207 5608
rect 3293 5594 3307 5608
rect 3393 5594 3407 5608
rect 3133 5553 3147 5567
rect 3213 5552 3227 5566
rect 2993 5533 3007 5547
rect 3073 5533 3087 5547
rect 3093 5513 3107 5527
rect 3253 5513 3267 5527
rect 2973 5493 2987 5507
rect 3033 5393 3047 5407
rect 2973 5374 2987 5388
rect 3373 5533 3387 5547
rect 3433 5553 3447 5567
rect 3553 5852 3567 5866
rect 3633 5833 3647 5847
rect 3793 5852 3807 5866
rect 4633 5973 4647 5987
rect 4673 5973 4687 5987
rect 4773 5993 4787 6007
rect 4533 5953 4547 5967
rect 4593 5953 4607 5967
rect 4013 5933 4027 5947
rect 4093 5933 4107 5947
rect 4273 5933 4287 5947
rect 4453 5933 4467 5947
rect 3953 5913 3967 5927
rect 3833 5894 3847 5908
rect 3873 5894 3887 5908
rect 3913 5894 3927 5908
rect 3973 5893 3987 5907
rect 3893 5852 3907 5866
rect 3933 5852 3947 5866
rect 3673 5773 3687 5787
rect 3733 5733 3747 5747
rect 3513 5693 3527 5707
rect 3633 5673 3647 5687
rect 3733 5673 3747 5687
rect 3613 5633 3627 5647
rect 3533 5594 3547 5608
rect 3573 5594 3587 5608
rect 3613 5594 3627 5608
rect 3513 5552 3527 5566
rect 3413 5533 3427 5547
rect 3593 5553 3607 5567
rect 3333 5513 3347 5527
rect 3553 5513 3567 5527
rect 3573 5493 3587 5507
rect 3293 5473 3307 5487
rect 3433 5473 3447 5487
rect 3193 5413 3207 5427
rect 3133 5393 3147 5407
rect 3273 5374 3287 5388
rect 3693 5633 3707 5647
rect 3733 5594 3747 5608
rect 3633 5553 3647 5567
rect 3673 5552 3687 5566
rect 3752 5553 3766 5567
rect 3773 5553 3787 5567
rect 3713 5513 3727 5527
rect 3593 5473 3607 5487
rect 3773 5532 3787 5546
rect 3773 5493 3787 5507
rect 3753 5473 3767 5487
rect 3573 5453 3587 5467
rect 3633 5453 3647 5467
rect 3693 5433 3707 5447
rect 3513 5413 3527 5427
rect 3593 5413 3607 5427
rect 3513 5373 3527 5387
rect 3693 5374 3707 5388
rect 2993 5332 3007 5346
rect 3033 5332 3047 5346
rect 2953 5293 2967 5307
rect 3153 5332 3167 5346
rect 3193 5332 3207 5346
rect 3193 5293 3207 5307
rect 2893 5253 2907 5267
rect 3113 5253 3127 5267
rect 3253 5253 3267 5267
rect 3453 5332 3467 5346
rect 3573 5332 3587 5346
rect 3313 5233 3327 5247
rect 3413 5233 3427 5247
rect 2893 5213 2907 5227
rect 3113 5213 3127 5227
rect 3073 5173 3087 5187
rect 2813 4853 2827 4867
rect 2793 4753 2807 4767
rect 2753 4653 2767 4667
rect 2713 4633 2727 4647
rect 2773 4593 2787 4607
rect 2693 4554 2707 4568
rect 2733 4554 2747 4568
rect 2773 4553 2787 4567
rect 2653 4513 2667 4527
rect 2713 4512 2727 4526
rect 2773 4513 2787 4527
rect 2633 4473 2647 4487
rect 2732 4473 2746 4487
rect 2753 4473 2767 4487
rect 2573 4453 2587 4467
rect 2533 4433 2547 4447
rect 2453 4353 2467 4367
rect 2393 4334 2407 4348
rect 2413 4292 2427 4306
rect 2473 4253 2487 4267
rect 2513 4253 2527 4267
rect 2373 4173 2387 4187
rect 2333 4153 2347 4167
rect 2473 4153 2487 4167
rect 2393 4093 2407 4107
rect 2313 4053 2327 4067
rect 2393 4034 2407 4048
rect 2173 3993 2187 4007
rect 2153 3953 2167 3967
rect 2213 3973 2227 3987
rect 2393 3973 2407 3987
rect 2193 3933 2207 3947
rect 2273 3933 2287 3947
rect 1913 3913 1927 3927
rect 1993 3913 2007 3927
rect 2053 3913 2067 3927
rect 2133 3913 2147 3927
rect 1893 3853 1907 3867
rect 1813 3833 1827 3847
rect 1853 3833 1867 3847
rect 1813 3772 1827 3786
rect 1773 3753 1787 3767
rect 1733 3693 1747 3707
rect 1733 3653 1747 3667
rect 1693 3514 1707 3528
rect 1673 3473 1687 3487
rect 1613 3453 1627 3467
rect 1653 3453 1667 3467
rect 1593 3433 1607 3447
rect 1673 3433 1687 3447
rect 1573 3393 1587 3407
rect 1693 3413 1707 3427
rect 1673 3353 1687 3367
rect 1593 3333 1607 3347
rect 1652 3333 1666 3347
rect 1593 3294 1607 3308
rect 1573 3252 1587 3266
rect 1633 3253 1647 3267
rect 1613 3173 1627 3187
rect 1533 3093 1547 3107
rect 1593 3093 1607 3107
rect 1513 2993 1527 3007
rect 1613 3013 1627 3027
rect 1513 2953 1527 2967
rect 1593 2953 1607 2967
rect 1453 2913 1467 2927
rect 1393 2853 1407 2867
rect 1313 2813 1327 2827
rect 1573 2853 1587 2867
rect 1193 2732 1207 2746
rect 1233 2732 1247 2746
rect 1313 2774 1327 2788
rect 1353 2774 1367 2788
rect 1393 2774 1407 2788
rect 1432 2773 1446 2787
rect 1453 2773 1467 2787
rect 1513 2774 1527 2788
rect 1553 2774 1567 2788
rect 1313 2733 1327 2747
rect 1293 2693 1307 2707
rect 1273 2633 1287 2647
rect 1253 2613 1267 2627
rect 1153 2533 1167 2547
rect 1153 2474 1167 2488
rect 1193 2474 1207 2488
rect 1233 2473 1247 2487
rect 1133 2373 1147 2387
rect 1213 2433 1227 2447
rect 1233 2413 1247 2427
rect 1433 2693 1447 2707
rect 1373 2613 1387 2627
rect 1333 2474 1347 2488
rect 1273 2433 1287 2447
rect 1373 2433 1387 2447
rect 1353 2413 1367 2427
rect 1313 2393 1327 2407
rect 1253 2373 1267 2387
rect 1213 2333 1227 2347
rect 1313 2333 1327 2347
rect 1253 2293 1267 2307
rect 1173 2273 1187 2287
rect 1213 2273 1227 2287
rect 1093 2253 1107 2267
rect 1153 2254 1167 2268
rect 1093 2193 1107 2207
rect 1173 2173 1187 2187
rect 1033 2133 1047 2147
rect 1213 2133 1227 2147
rect 1233 2113 1247 2127
rect 1333 2293 1347 2307
rect 1393 2413 1407 2427
rect 1493 2732 1507 2746
rect 1673 3332 1687 3346
rect 1673 3253 1687 3267
rect 2233 3814 2247 3828
rect 2273 3813 2287 3827
rect 1993 3772 2007 3786
rect 1933 3693 1947 3707
rect 1873 3593 1887 3607
rect 1753 3573 1767 3587
rect 1853 3573 1867 3587
rect 1833 3553 1847 3567
rect 1793 3514 1807 3528
rect 1753 3413 1767 3427
rect 1953 3514 1967 3528
rect 1893 3473 1907 3487
rect 1873 3433 1887 3447
rect 1813 3393 1827 3407
rect 1753 3333 1767 3347
rect 1733 3313 1747 3327
rect 1793 3313 1807 3327
rect 1833 3296 1847 3310
rect 1733 3252 1747 3266
rect 1753 3213 1767 3227
rect 1693 3173 1707 3187
rect 1793 3233 1807 3247
rect 1793 3193 1807 3207
rect 1773 3173 1787 3187
rect 1733 3093 1747 3107
rect 1653 3013 1667 3027
rect 1613 2833 1627 2847
rect 1733 2833 1747 2847
rect 1633 2774 1647 2788
rect 1673 2776 1687 2790
rect 1593 2733 1607 2747
rect 1613 2693 1627 2707
rect 1653 2693 1667 2707
rect 1473 2653 1487 2667
rect 1553 2653 1567 2667
rect 1593 2533 1607 2547
rect 1513 2476 1527 2490
rect 1593 2433 1607 2447
rect 1473 2413 1487 2427
rect 1453 2393 1467 2407
rect 1593 2393 1607 2407
rect 1633 2553 1647 2567
rect 2193 3753 2207 3767
rect 2073 3733 2087 3747
rect 2173 3733 2187 3747
rect 2093 3593 2107 3607
rect 2033 3553 2047 3567
rect 2073 3553 2087 3567
rect 2373 3733 2387 3747
rect 2413 3953 2427 3967
rect 2573 4393 2587 4407
rect 2673 4393 2687 4407
rect 2593 4373 2607 4387
rect 2633 4334 2647 4348
rect 2673 4334 2687 4348
rect 2913 5074 2927 5088
rect 2953 5074 2967 5088
rect 3153 5173 3167 5187
rect 3113 5153 3127 5167
rect 3133 5113 3147 5127
rect 2893 5032 2907 5046
rect 3013 5032 3027 5046
rect 2973 4973 2987 4987
rect 2853 4933 2867 4947
rect 2933 4933 2947 4947
rect 2853 4854 2867 4868
rect 2953 4854 2967 4868
rect 2833 4793 2847 4807
rect 2893 4793 2907 4807
rect 2813 4733 2827 4747
rect 2813 4612 2827 4626
rect 2793 4493 2807 4507
rect 2573 4292 2587 4306
rect 2613 4292 2627 4306
rect 2573 4213 2587 4227
rect 2553 4073 2567 4087
rect 2533 4053 2547 4067
rect 2653 4173 2667 4187
rect 2613 4133 2627 4147
rect 2493 3992 2507 4006
rect 2553 3992 2567 4006
rect 2653 3993 2667 4007
rect 2593 3933 2607 3947
rect 2573 3893 2587 3907
rect 2353 3713 2367 3727
rect 2233 3573 2247 3587
rect 2273 3573 2287 3587
rect 2213 3493 2227 3507
rect 1913 3433 1927 3447
rect 1993 3433 2007 3447
rect 1913 3296 1927 3310
rect 2033 3293 2047 3307
rect 2013 3250 2027 3264
rect 1953 3193 1967 3207
rect 2033 3193 2047 3207
rect 1993 3153 2007 3167
rect 1913 3113 1927 3127
rect 1893 3073 1907 3087
rect 1813 3013 1827 3027
rect 1853 2994 1867 3008
rect 1973 2994 1987 3008
rect 1893 2953 1907 2967
rect 1833 2893 1847 2907
rect 1773 2853 1787 2867
rect 1753 2730 1767 2744
rect 1733 2553 1747 2567
rect 1753 2533 1767 2547
rect 1773 2493 1787 2507
rect 1653 2474 1667 2488
rect 1693 2474 1707 2488
rect 1733 2474 1747 2488
rect 1633 2432 1647 2446
rect 1673 2432 1687 2446
rect 1713 2393 1727 2407
rect 1713 2372 1727 2386
rect 1533 2353 1547 2367
rect 1613 2353 1627 2367
rect 1453 2293 1467 2307
rect 1413 2193 1427 2207
rect 1333 2173 1347 2187
rect 1493 2254 1507 2268
rect 1613 2313 1627 2327
rect 1573 2254 1587 2268
rect 1553 2212 1567 2226
rect 1493 2193 1507 2207
rect 1533 2193 1547 2207
rect 1413 2153 1427 2167
rect 1453 2153 1467 2167
rect 1233 2053 1247 2067
rect 1273 2053 1287 2067
rect 1313 2053 1327 2067
rect 1433 2053 1447 2067
rect 1133 1973 1147 1987
rect 1013 1956 1027 1970
rect 1133 1956 1147 1970
rect 953 1853 967 1867
rect 993 1853 1007 1867
rect 933 1833 947 1847
rect 733 1734 747 1748
rect 813 1734 827 1748
rect 853 1734 867 1748
rect 913 1734 927 1748
rect 533 1653 547 1667
rect 753 1692 767 1706
rect 793 1692 807 1706
rect 693 1613 707 1627
rect 533 1533 547 1547
rect 453 1473 467 1487
rect 613 1473 627 1487
rect 493 1434 507 1448
rect 532 1434 546 1448
rect 553 1433 567 1447
rect 653 1453 667 1467
rect 873 1692 887 1706
rect 913 1693 927 1707
rect 1113 1913 1127 1927
rect 1093 1873 1107 1887
rect 1013 1833 1027 1847
rect 993 1773 1007 1787
rect 953 1733 967 1747
rect 1053 1736 1067 1750
rect 1013 1692 1027 1706
rect 973 1653 987 1667
rect 933 1613 947 1627
rect 1233 1873 1247 1887
rect 1133 1833 1147 1847
rect 853 1513 867 1527
rect 1113 1513 1127 1527
rect 833 1473 847 1487
rect 833 1452 847 1466
rect 773 1434 787 1448
rect 553 1392 567 1406
rect 353 1353 367 1367
rect 453 1353 467 1367
rect 533 1353 547 1367
rect 353 1313 367 1327
rect 313 1273 327 1287
rect 293 1213 307 1227
rect 233 1172 247 1186
rect 333 1214 347 1228
rect 273 1153 287 1167
rect 313 1153 327 1167
rect 233 953 247 967
rect 313 953 327 967
rect 153 873 167 887
rect 193 873 207 887
rect 413 1214 427 1228
rect 533 1332 547 1346
rect 493 1313 507 1327
rect 353 1172 367 1186
rect 393 1172 407 1186
rect 433 1172 447 1186
rect 713 1392 727 1406
rect 753 1392 767 1406
rect 793 1392 807 1406
rect 673 1353 687 1367
rect 653 1333 667 1347
rect 633 1313 647 1327
rect 833 1313 847 1327
rect 653 1293 667 1307
rect 573 1214 587 1228
rect 653 1216 667 1230
rect 1053 1473 1067 1487
rect 1333 1793 1347 1807
rect 1313 1773 1327 1787
rect 1273 1733 1287 1747
rect 1293 1713 1307 1727
rect 1173 1690 1187 1704
rect 1273 1690 1287 1704
rect 1373 1734 1387 1748
rect 1413 1734 1427 1748
rect 1513 1913 1527 1927
rect 1473 1873 1487 1887
rect 1673 2254 1687 2268
rect 1753 2333 1767 2347
rect 1753 2254 1767 2268
rect 1693 2212 1707 2226
rect 1653 2193 1667 2207
rect 1713 2193 1727 2207
rect 1573 2073 1587 2087
rect 1613 2073 1627 2087
rect 1613 2033 1627 2047
rect 1593 1912 1607 1926
rect 1653 1910 1667 1924
rect 1713 1913 1727 1927
rect 1633 1873 1647 1887
rect 1533 1853 1547 1867
rect 1513 1833 1527 1847
rect 1473 1733 1487 1747
rect 1553 1813 1567 1827
rect 1593 1793 1607 1807
rect 1313 1692 1327 1706
rect 1353 1692 1367 1706
rect 1393 1692 1407 1706
rect 1453 1692 1467 1706
rect 1493 1692 1507 1706
rect 1293 1653 1307 1667
rect 1333 1653 1347 1667
rect 1373 1653 1387 1667
rect 1533 1653 1547 1667
rect 1273 1613 1287 1627
rect 1253 1513 1267 1527
rect 873 1433 887 1447
rect 933 1434 947 1448
rect 1093 1434 1107 1448
rect 1133 1434 1147 1448
rect 853 1213 867 1227
rect 553 1172 567 1186
rect 493 1153 507 1167
rect 533 1153 547 1167
rect 493 953 507 967
rect 373 914 387 928
rect 413 913 427 927
rect 593 1133 607 1147
rect 753 953 767 967
rect 713 933 727 947
rect 133 853 147 867
rect 333 853 347 867
rect 373 853 387 867
rect 293 733 307 747
rect 333 694 347 708
rect 213 653 227 667
rect 313 652 327 666
rect 113 593 127 607
rect 113 473 127 487
rect 353 473 367 487
rect 173 393 187 407
rect 233 394 247 408
rect 613 913 627 927
rect 673 914 687 928
rect 513 872 527 886
rect 573 873 587 887
rect 613 853 627 867
rect 653 853 667 867
rect 513 733 527 747
rect 453 694 467 708
rect 413 653 427 667
rect 413 613 427 627
rect 393 533 407 547
rect 373 433 387 447
rect 433 573 447 587
rect 493 653 507 667
rect 473 473 487 487
rect 473 433 487 447
rect 413 413 427 427
rect 393 394 407 408
rect 453 394 467 408
rect 213 313 227 327
rect 93 253 107 267
rect 153 213 167 227
rect 213 213 227 227
rect 93 193 107 207
rect 113 174 127 188
rect 213 174 227 188
rect 373 352 387 366
rect 313 293 327 307
rect 393 273 407 287
rect 433 353 447 367
rect 433 293 447 307
rect 513 633 527 647
rect 573 753 587 767
rect 653 813 667 827
rect 653 753 667 767
rect 713 753 727 767
rect 613 694 627 708
rect 593 633 607 647
rect 533 553 547 567
rect 613 553 627 567
rect 573 413 587 427
rect 533 394 547 408
rect 633 493 647 507
rect 613 393 627 407
rect 553 333 567 347
rect 613 353 627 367
rect 693 694 707 708
rect 713 652 727 666
rect 653 413 667 427
rect 833 1170 847 1184
rect 1033 1392 1047 1406
rect 913 1353 927 1367
rect 953 1353 967 1367
rect 1013 1353 1027 1367
rect 953 1293 967 1307
rect 893 1213 907 1227
rect 953 1214 967 1228
rect 933 1172 947 1186
rect 893 1133 907 1147
rect 853 914 867 928
rect 773 873 787 887
rect 833 872 847 886
rect 873 872 887 886
rect 772 694 786 708
rect 793 694 807 708
rect 833 694 847 708
rect 873 694 887 708
rect 773 653 787 667
rect 853 652 867 666
rect 793 633 807 647
rect 773 573 787 587
rect 1013 1172 1027 1186
rect 993 1133 1007 1147
rect 973 1013 987 1027
rect 973 933 987 947
rect 1113 1392 1127 1406
rect 1033 1033 1047 1047
rect 1013 914 1027 928
rect 993 872 1007 886
rect 953 813 967 827
rect 1213 1434 1227 1448
rect 1273 1413 1287 1427
rect 1193 1392 1207 1406
rect 1213 1371 1227 1385
rect 1153 1353 1167 1367
rect 1113 1313 1127 1327
rect 1313 1353 1327 1367
rect 1193 1333 1207 1347
rect 1233 1333 1247 1347
rect 1153 1293 1167 1307
rect 1093 1172 1107 1186
rect 1173 1172 1187 1186
rect 1133 1113 1147 1127
rect 1213 1233 1227 1247
rect 1253 1214 1267 1228
rect 1233 1172 1247 1186
rect 1373 1573 1387 1587
rect 1613 1713 1627 1727
rect 1613 1613 1627 1627
rect 1673 1833 1687 1847
rect 1853 2730 1867 2744
rect 1853 2613 1867 2627
rect 1913 2933 1927 2947
rect 2113 3433 2127 3447
rect 2133 3373 2147 3387
rect 2193 3373 2207 3387
rect 2153 3313 2167 3327
rect 2213 3312 2227 3326
rect 2193 3293 2207 3307
rect 2113 3233 2127 3247
rect 2073 3173 2087 3187
rect 2053 3153 2067 3167
rect 2033 3133 2047 3147
rect 2013 3113 2027 3127
rect 2193 3253 2207 3267
rect 2213 3233 2227 3247
rect 2133 3173 2147 3187
rect 2173 3173 2187 3187
rect 2113 3093 2127 3107
rect 2013 3033 2027 3047
rect 2033 2996 2047 3010
rect 2133 3073 2147 3087
rect 2113 2953 2127 2967
rect 1993 2913 2007 2927
rect 1973 2873 1987 2887
rect 2133 2893 2147 2907
rect 1973 2852 1987 2866
rect 2033 2813 2047 2827
rect 2053 2774 2067 2788
rect 2093 2774 2107 2788
rect 2213 3053 2227 3067
rect 2333 3553 2347 3567
rect 2273 3516 2287 3530
rect 2253 3473 2267 3487
rect 2353 3433 2367 3447
rect 2253 3393 2267 3407
rect 2313 3393 2327 3407
rect 2353 3333 2367 3347
rect 2413 3713 2427 3727
rect 2393 3573 2407 3587
rect 2453 3693 2467 3707
rect 2453 3633 2467 3647
rect 2593 3813 2607 3827
rect 2633 3814 2647 3828
rect 2693 4292 2707 4306
rect 2753 4292 2767 4306
rect 2713 4253 2727 4267
rect 2733 4233 2747 4247
rect 2773 4233 2787 4247
rect 2713 4133 2727 4147
rect 2753 4153 2767 4167
rect 2753 3992 2767 4006
rect 2693 3893 2707 3907
rect 2693 3853 2707 3867
rect 2773 3853 2787 3867
rect 2853 4653 2867 4667
rect 2913 4733 2927 4747
rect 3093 5032 3107 5046
rect 3053 4973 3067 4987
rect 3073 4893 3087 4907
rect 3113 4854 3127 4868
rect 3213 5093 3227 5107
rect 3253 5074 3267 5088
rect 3313 5074 3327 5088
rect 3233 5032 3247 5046
rect 3273 5033 3287 5047
rect 3193 4993 3207 5007
rect 3293 4993 3307 5007
rect 3173 4953 3187 4967
rect 3153 4933 3167 4947
rect 3153 4893 3167 4907
rect 3013 4713 3027 4727
rect 3133 4812 3147 4826
rect 3093 4753 3107 4767
rect 2993 4633 3007 4647
rect 3053 4633 3067 4647
rect 2933 4554 2947 4568
rect 2973 4554 2987 4568
rect 2853 4493 2867 4507
rect 2913 4512 2927 4526
rect 3053 4573 3067 4587
rect 3093 4554 3107 4568
rect 2833 4452 2847 4466
rect 2813 4433 2827 4447
rect 2813 4353 2827 4367
rect 2833 4333 2847 4347
rect 2933 4493 2947 4507
rect 2893 4353 2907 4367
rect 2813 4292 2827 4306
rect 2853 4292 2867 4306
rect 2993 4513 3007 4527
rect 3073 4512 3087 4526
rect 3193 4933 3207 4947
rect 3193 4854 3207 4868
rect 3233 4854 3247 4868
rect 3273 4854 3287 4868
rect 3213 4812 3227 4826
rect 3173 4773 3187 4787
rect 3153 4753 3167 4767
rect 3153 4713 3167 4727
rect 3713 5332 3727 5346
rect 3693 5293 3707 5307
rect 3673 5253 3687 5267
rect 3513 5213 3527 5227
rect 3493 5073 3507 5087
rect 3313 4873 3327 4887
rect 3433 5032 3447 5046
rect 3473 5033 3487 5047
rect 3393 4993 3407 5007
rect 3493 4993 3507 5007
rect 3473 4933 3487 4947
rect 3413 4853 3427 4867
rect 3673 5173 3687 5187
rect 3713 5253 3727 5267
rect 3733 5233 3747 5247
rect 3773 5233 3787 5247
rect 3713 5213 3727 5227
rect 3693 5153 3707 5167
rect 3713 5133 3727 5147
rect 3693 5113 3707 5127
rect 3553 5074 3567 5088
rect 3613 5074 3627 5088
rect 3653 5074 3667 5088
rect 3753 5113 3767 5127
rect 3533 5033 3547 5047
rect 3513 4853 3527 4867
rect 3293 4773 3307 4787
rect 3273 4693 3287 4707
rect 3153 4633 3167 4647
rect 3033 4493 3047 4507
rect 3213 4573 3227 4587
rect 3273 4573 3287 4587
rect 3253 4554 3267 4568
rect 3233 4512 3247 4526
rect 3293 4513 3307 4527
rect 3132 4492 3146 4506
rect 3153 4493 3167 4507
rect 3193 4493 3207 4507
rect 3113 4473 3127 4487
rect 3053 4453 3067 4467
rect 3033 4413 3047 4427
rect 2973 4373 2987 4387
rect 3093 4413 3107 4427
rect 3052 4353 3066 4367
rect 3073 4353 3087 4367
rect 3093 4333 3107 4347
rect 3013 4292 3027 4306
rect 3053 4292 3067 4306
rect 3093 4292 3107 4306
rect 2953 4273 2967 4287
rect 2833 4193 2847 4207
rect 2913 4193 2927 4207
rect 2853 4173 2867 4187
rect 2913 4153 2927 4167
rect 2833 4133 2847 4147
rect 2893 4133 2907 4147
rect 2833 4093 2847 4107
rect 2893 4093 2907 4107
rect 2813 4073 2827 4087
rect 2573 3733 2587 3747
rect 2613 3733 2627 3747
rect 2613 3693 2627 3707
rect 2593 3653 2607 3667
rect 2613 3613 2627 3627
rect 2593 3593 2607 3607
rect 2493 3573 2507 3587
rect 2553 3533 2567 3547
rect 2493 3514 2507 3528
rect 2533 3514 2547 3528
rect 2413 3473 2427 3487
rect 2673 3733 2687 3747
rect 2873 4073 2887 4087
rect 3133 4413 3147 4427
rect 3133 4333 3147 4347
rect 3253 4473 3267 4487
rect 3233 4453 3247 4467
rect 3233 4333 3247 4347
rect 3113 4253 3127 4267
rect 3093 4233 3107 4247
rect 3013 4113 3027 4127
rect 2973 4093 2987 4107
rect 2913 3973 2927 3987
rect 2833 3814 2847 3828
rect 2893 3814 2907 3828
rect 2733 3772 2747 3786
rect 2693 3713 2707 3727
rect 2873 3772 2887 3786
rect 2913 3772 2927 3786
rect 3013 4034 3027 4048
rect 3173 4292 3187 4306
rect 3133 4173 3147 4187
rect 3213 4273 3227 4287
rect 3193 4253 3207 4267
rect 3173 4113 3187 4127
rect 3153 4034 3167 4048
rect 3213 4213 3227 4227
rect 3373 4673 3387 4687
rect 3333 4553 3347 4567
rect 3373 4554 3387 4568
rect 3453 4753 3467 4767
rect 3473 4733 3487 4747
rect 3433 4613 3447 4627
rect 3413 4553 3427 4567
rect 3413 4513 3427 4527
rect 3733 5073 3747 5087
rect 3773 5074 3787 5088
rect 3573 4993 3587 5007
rect 3613 4993 3627 5007
rect 3713 5032 3727 5046
rect 3753 5033 3767 5047
rect 3673 4953 3687 4967
rect 3693 4933 3707 4947
rect 3553 4913 3567 4927
rect 3673 4893 3687 4907
rect 3613 4873 3627 4887
rect 3553 4733 3567 4747
rect 3633 4812 3647 4826
rect 3593 4713 3607 4727
rect 3633 4693 3647 4707
rect 3673 4693 3687 4707
rect 3592 4672 3606 4686
rect 3613 4673 3627 4687
rect 3493 4553 3507 4567
rect 3533 4554 3547 4568
rect 3753 4993 3767 5007
rect 3733 4893 3747 4907
rect 3773 4973 3787 4987
rect 3833 5833 3847 5847
rect 3833 5733 3847 5747
rect 3973 5852 3987 5866
rect 4053 5894 4067 5908
rect 4153 5893 4167 5907
rect 4233 5894 4247 5908
rect 4333 5893 4347 5907
rect 4373 5894 4387 5908
rect 4413 5894 4427 5908
rect 4473 5913 4487 5927
rect 4453 5893 4467 5907
rect 4113 5852 4127 5866
rect 4013 5813 4027 5827
rect 3973 5653 3987 5667
rect 3973 5594 3987 5608
rect 4233 5833 4247 5847
rect 4333 5852 4347 5866
rect 4253 5793 4267 5807
rect 4233 5773 4247 5787
rect 4213 5733 4227 5747
rect 4133 5713 4147 5727
rect 4113 5693 4127 5707
rect 4053 5673 4067 5687
rect 3873 5533 3887 5547
rect 4033 5533 4047 5547
rect 4113 5533 4127 5547
rect 3813 5493 3827 5507
rect 4073 5493 4087 5507
rect 3873 5453 3887 5467
rect 4113 5453 4127 5467
rect 4033 5433 4047 5447
rect 3913 5374 3927 5388
rect 3993 5374 4007 5388
rect 4093 5374 4107 5388
rect 3893 5332 3907 5346
rect 4013 5332 4027 5346
rect 4053 5332 4067 5346
rect 3813 5253 3827 5267
rect 3853 5253 3867 5267
rect 3813 5193 3827 5207
rect 4033 5273 4047 5287
rect 4013 5213 4027 5227
rect 3933 5153 3947 5167
rect 3853 5133 3867 5147
rect 3873 5074 3887 5088
rect 3853 5032 3867 5046
rect 3893 4993 3907 5007
rect 3812 4973 3826 4987
rect 3833 4973 3847 4987
rect 3713 4813 3727 4827
rect 3693 4673 3707 4687
rect 3633 4613 3647 4627
rect 3633 4554 3647 4568
rect 3673 4554 3687 4568
rect 3773 4812 3787 4826
rect 3753 4793 3767 4807
rect 3733 4753 3747 4767
rect 3773 4753 3787 4767
rect 3753 4554 3767 4568
rect 3393 4493 3407 4507
rect 3333 4473 3347 4487
rect 3373 4373 3387 4387
rect 3313 4353 3327 4367
rect 3333 4334 3347 4348
rect 3373 4333 3387 4347
rect 3353 4292 3367 4306
rect 3473 4493 3487 4507
rect 3413 4473 3427 4487
rect 3413 4433 3427 4447
rect 3473 4413 3487 4427
rect 3553 4512 3567 4526
rect 3613 4512 3627 4526
rect 3693 4512 3707 4526
rect 3512 4493 3526 4507
rect 3533 4493 3547 4507
rect 3633 4493 3647 4507
rect 3673 4493 3687 4507
rect 3553 4473 3567 4487
rect 3533 4453 3547 4467
rect 3493 4393 3507 4407
rect 3533 4334 3547 4348
rect 3413 4293 3427 4307
rect 3453 4292 3467 4306
rect 3493 4292 3507 4306
rect 3393 4253 3407 4267
rect 3353 4233 3367 4247
rect 3293 4213 3307 4227
rect 3373 4213 3387 4227
rect 3253 4193 3267 4207
rect 3233 4113 3247 4127
rect 3353 4053 3367 4067
rect 3313 4036 3327 4050
rect 2973 3973 2987 3987
rect 3053 3973 3067 3987
rect 2993 3814 3007 3828
rect 2833 3693 2847 3707
rect 2673 3673 2687 3687
rect 2673 3573 2687 3587
rect 2873 3573 2887 3587
rect 2653 3493 2667 3507
rect 2813 3553 2827 3567
rect 2713 3533 2727 3547
rect 2753 3514 2767 3528
rect 2533 3453 2547 3467
rect 2633 3473 2647 3487
rect 2673 3473 2687 3487
rect 2593 3393 2607 3407
rect 2393 3373 2407 3387
rect 2473 3373 2487 3387
rect 2353 3294 2367 3308
rect 2253 3273 2267 3287
rect 2333 3252 2347 3266
rect 2373 3253 2387 3267
rect 2613 3353 2627 3367
rect 2293 3233 2307 3247
rect 2253 3173 2267 3187
rect 2233 3013 2247 3027
rect 2313 3133 2327 3147
rect 2473 3250 2487 3264
rect 2453 3213 2467 3227
rect 2413 3133 2427 3147
rect 2373 3093 2387 3107
rect 2573 3250 2587 3264
rect 2513 3213 2527 3227
rect 2613 3213 2627 3227
rect 2473 3153 2487 3167
rect 2453 3113 2467 3127
rect 2733 3472 2747 3486
rect 2653 3453 2667 3467
rect 2733 3353 2747 3367
rect 2653 3333 2667 3347
rect 2793 3473 2807 3487
rect 2953 3753 2967 3767
rect 3013 3772 3027 3786
rect 2973 3713 2987 3727
rect 2973 3673 2987 3687
rect 2953 3653 2967 3667
rect 3173 3992 3187 4006
rect 3153 3973 3167 3987
rect 3093 3813 3107 3827
rect 3033 3633 3047 3647
rect 3073 3633 3087 3647
rect 2933 3613 2947 3627
rect 3233 3953 3247 3967
rect 3173 3772 3187 3786
rect 3213 3773 3227 3787
rect 3153 3753 3167 3767
rect 3133 3733 3147 3747
rect 3113 3693 3127 3707
rect 3093 3613 3107 3627
rect 3133 3613 3147 3627
rect 3113 3593 3127 3607
rect 3053 3573 3067 3587
rect 3033 3532 3047 3546
rect 2933 3470 2947 3484
rect 2993 3470 3007 3484
rect 2793 3393 2807 3407
rect 2893 3393 2907 3407
rect 2773 3333 2787 3347
rect 2733 3313 2747 3327
rect 2713 3294 2727 3308
rect 2693 3213 2707 3227
rect 2653 3193 2667 3207
rect 2733 3193 2747 3207
rect 2693 3113 2707 3127
rect 2893 3333 2907 3347
rect 2853 3313 2867 3327
rect 2953 3333 2967 3347
rect 3013 3333 3027 3347
rect 2833 3252 2847 3266
rect 2873 3252 2887 3266
rect 2933 3253 2947 3267
rect 3133 3533 3147 3547
rect 3193 3693 3207 3707
rect 3173 3553 3187 3567
rect 3153 3513 3167 3527
rect 3053 3473 3067 3487
rect 3113 3472 3127 3486
rect 3153 3473 3167 3487
rect 3053 3353 3067 3367
rect 3033 3313 3047 3327
rect 3153 3313 3167 3327
rect 3313 3853 3327 3867
rect 3473 4253 3487 4267
rect 3453 4033 3467 4047
rect 3433 3990 3447 4004
rect 3293 3833 3307 3847
rect 3333 3833 3347 3847
rect 3313 3772 3327 3786
rect 3273 3673 3287 3687
rect 3233 3613 3247 3627
rect 3313 3613 3327 3627
rect 3213 3593 3227 3607
rect 3293 3573 3307 3587
rect 3213 3514 3227 3528
rect 3253 3514 3267 3528
rect 3473 3972 3487 3986
rect 3393 3873 3407 3887
rect 3413 3814 3427 3828
rect 3433 3753 3447 3767
rect 3393 3733 3407 3747
rect 3353 3713 3367 3727
rect 3353 3673 3367 3687
rect 3293 3513 3307 3527
rect 3333 3513 3347 3527
rect 3193 3296 3207 3310
rect 2993 3252 3007 3266
rect 3033 3252 3047 3266
rect 2873 3213 2887 3227
rect 2953 3213 2967 3227
rect 2793 3173 2807 3187
rect 2813 3153 2827 3167
rect 2473 3093 2487 3107
rect 2633 3093 2647 3107
rect 2333 3033 2347 3047
rect 2413 3033 2427 3047
rect 2193 2953 2207 2967
rect 2233 2952 2247 2966
rect 2313 2953 2327 2967
rect 2273 2933 2287 2947
rect 2253 2913 2267 2927
rect 2193 2793 2207 2807
rect 2233 2793 2247 2807
rect 2033 2732 2047 2746
rect 1993 2673 2007 2687
rect 1953 2613 1967 2627
rect 1893 2553 1907 2567
rect 1813 2474 1827 2488
rect 1993 2493 2007 2507
rect 1813 2433 1827 2447
rect 1873 2432 1887 2446
rect 2013 2413 2027 2427
rect 1793 2373 1807 2387
rect 1933 2373 1947 2387
rect 2113 2732 2127 2746
rect 2153 2732 2167 2746
rect 2193 2713 2207 2727
rect 2113 2553 2127 2567
rect 2053 2333 2067 2347
rect 1853 2313 1867 2327
rect 1813 2254 1827 2268
rect 2033 2253 2047 2267
rect 2093 2256 2107 2270
rect 2153 2474 2167 2488
rect 2373 2994 2387 3008
rect 2393 2952 2407 2966
rect 2433 2933 2447 2947
rect 2393 2893 2407 2907
rect 2333 2813 2347 2827
rect 2313 2774 2327 2788
rect 2353 2774 2367 2788
rect 2253 2733 2267 2747
rect 2293 2732 2307 2746
rect 2333 2713 2347 2727
rect 2693 3092 2707 3106
rect 2773 3093 2787 3107
rect 2673 3013 2687 3027
rect 2553 2994 2567 3008
rect 2493 2953 2507 2967
rect 2473 2933 2487 2947
rect 2453 2913 2467 2927
rect 2533 2952 2547 2966
rect 2533 2931 2547 2945
rect 2493 2873 2507 2887
rect 2433 2813 2447 2827
rect 2613 2950 2627 2964
rect 2573 2853 2587 2867
rect 2573 2813 2587 2827
rect 2533 2793 2547 2807
rect 2613 2793 2627 2807
rect 2473 2774 2487 2788
rect 2553 2773 2567 2787
rect 2453 2713 2467 2727
rect 2553 2693 2567 2707
rect 2413 2673 2427 2687
rect 2453 2673 2467 2687
rect 2493 2673 2507 2687
rect 2393 2653 2407 2667
rect 2433 2653 2447 2667
rect 2273 2553 2287 2567
rect 2233 2493 2247 2507
rect 2313 2493 2327 2507
rect 2253 2432 2267 2446
rect 2293 2432 2307 2446
rect 2213 2413 2227 2427
rect 2173 2393 2187 2407
rect 2373 2413 2387 2427
rect 2413 2353 2427 2367
rect 2253 2313 2267 2327
rect 1773 2193 1787 2207
rect 1873 2210 1887 2224
rect 1913 2210 1927 2224
rect 1833 2153 1847 2167
rect 1773 1993 1787 2007
rect 1953 2033 1967 2047
rect 1893 1993 1907 2007
rect 1953 1993 1967 2007
rect 1833 1956 1847 1970
rect 1873 1956 1887 1970
rect 1733 1873 1747 1887
rect 1993 2213 2007 2227
rect 2033 2212 2047 2226
rect 2033 2093 2047 2107
rect 1993 1993 2007 2007
rect 1973 1973 1987 1987
rect 1973 1912 1987 1926
rect 1933 1893 1947 1907
rect 2013 1893 2027 1907
rect 1893 1853 1907 1867
rect 1833 1833 1847 1847
rect 1873 1833 1887 1847
rect 1813 1813 1827 1827
rect 1713 1773 1727 1787
rect 1753 1736 1767 1750
rect 1693 1653 1707 1667
rect 1813 1613 1827 1627
rect 1633 1593 1647 1607
rect 1713 1593 1727 1607
rect 1673 1513 1687 1527
rect 1553 1493 1567 1507
rect 1593 1493 1607 1507
rect 1413 1434 1427 1448
rect 1533 1433 1547 1447
rect 1393 1373 1407 1387
rect 1473 1390 1487 1404
rect 1533 1390 1547 1404
rect 1433 1293 1447 1307
rect 1413 1253 1427 1267
rect 1473 1216 1487 1230
rect 1433 1172 1447 1186
rect 1273 1153 1287 1167
rect 1313 1153 1327 1167
rect 1433 1113 1447 1127
rect 1193 1053 1207 1067
rect 1453 953 1467 967
rect 1073 913 1087 927
rect 1133 914 1147 928
rect 1233 914 1247 928
rect 1273 914 1287 928
rect 1513 916 1527 930
rect 953 733 967 747
rect 1053 733 1067 747
rect 913 553 927 567
rect 773 533 787 547
rect 673 394 687 408
rect 713 394 727 408
rect 753 394 767 408
rect 653 353 667 367
rect 633 333 647 347
rect 533 293 547 307
rect 613 293 627 307
rect 473 273 487 287
rect 313 253 327 267
rect 253 173 267 187
rect 693 352 707 366
rect 573 176 587 190
rect 653 176 667 190
rect 1153 873 1167 887
rect 1233 873 1247 887
rect 1293 872 1307 886
rect 1173 833 1187 847
rect 1153 793 1167 807
rect 1113 694 1127 708
rect 1253 694 1267 708
rect 1333 870 1347 884
rect 1533 873 1547 887
rect 1433 694 1447 708
rect 1473 696 1487 710
rect 1273 652 1287 666
rect 1413 652 1427 666
rect 1133 633 1147 647
rect 1313 613 1327 627
rect 1153 553 1167 567
rect 1113 533 1127 547
rect 1013 513 1027 527
rect 1073 513 1087 527
rect 993 453 1007 467
rect 1033 453 1047 467
rect 813 394 827 408
rect 853 394 867 408
rect 973 394 987 408
rect 93 132 107 146
rect 153 132 167 146
rect 193 132 207 146
rect 233 132 247 146
rect 913 333 927 347
rect 873 313 887 327
rect 953 273 967 287
rect 833 153 847 167
rect 53 13 67 27
rect 93 13 107 27
rect 693 130 707 144
rect 893 132 907 146
rect 1033 413 1047 427
rect 1013 393 1027 407
rect 1153 433 1167 447
rect 1013 353 1027 367
rect 1053 353 1067 367
rect 1213 394 1227 408
rect 993 313 1007 327
rect 973 233 987 247
rect 1153 352 1167 366
rect 1033 273 1047 287
rect 1233 352 1247 366
rect 1433 573 1447 587
rect 1613 1473 1627 1487
rect 1593 1170 1607 1184
rect 1653 1170 1667 1184
rect 1693 1170 1707 1184
rect 1673 993 1687 1007
rect 1633 914 1647 928
rect 1593 873 1607 887
rect 1553 833 1567 847
rect 1653 872 1667 886
rect 1613 853 1627 867
rect 1693 853 1707 867
rect 1593 793 1607 807
rect 1553 694 1567 708
rect 1553 653 1567 667
rect 1593 613 1607 627
rect 1693 652 1707 666
rect 1453 533 1467 547
rect 1533 533 1547 547
rect 1673 533 1687 547
rect 1433 493 1447 507
rect 1373 394 1387 408
rect 1413 394 1427 408
rect 1313 273 1327 287
rect 993 174 1007 188
rect 1193 193 1207 207
rect 1253 193 1267 207
rect 1013 132 1027 146
rect 1113 173 1127 187
rect 1253 176 1267 190
rect 1393 352 1407 366
rect 1533 473 1547 487
rect 1693 453 1707 467
rect 1533 433 1547 447
rect 1513 394 1527 408
rect 1553 394 1567 408
rect 1673 393 1687 407
rect 1493 352 1507 366
rect 1513 333 1527 347
rect 1493 293 1507 307
rect 1113 132 1127 146
rect 1153 132 1167 146
rect 1193 132 1207 146
rect 1333 130 1347 144
rect 1373 130 1387 144
rect 1433 130 1447 144
rect 1473 130 1487 144
rect 1573 353 1587 367
rect 1533 273 1547 287
rect 1673 293 1687 307
rect 1593 273 1607 287
rect 1633 273 1647 287
rect 1793 1573 1807 1587
rect 1973 1773 1987 1787
rect 2193 2254 2207 2268
rect 2213 2212 2227 2226
rect 2333 2212 2347 2226
rect 2333 2133 2347 2147
rect 2273 2013 2287 2027
rect 2133 1993 2147 2007
rect 2213 1993 2227 2007
rect 2053 1954 2067 1968
rect 2033 1773 2047 1787
rect 2113 1954 2127 1968
rect 2153 1954 2167 1968
rect 2073 1913 2087 1927
rect 2133 1912 2147 1926
rect 2133 1773 2147 1787
rect 2013 1734 2027 1748
rect 2053 1734 2067 1748
rect 2253 1912 2267 1926
rect 2333 1910 2347 1924
rect 2453 2613 2467 2627
rect 2433 2273 2447 2287
rect 2553 2513 2567 2527
rect 2493 2476 2507 2490
rect 2593 2732 2607 2746
rect 2633 2732 2647 2746
rect 2593 2613 2607 2627
rect 2673 2553 2687 2567
rect 2573 2473 2587 2487
rect 2473 2433 2487 2447
rect 2593 2373 2607 2387
rect 2473 2353 2487 2367
rect 2553 2333 2567 2347
rect 2533 2313 2547 2327
rect 2453 2253 2467 2267
rect 2633 2254 2647 2268
rect 2553 2212 2567 2226
rect 2613 2212 2627 2226
rect 2473 2053 2487 2067
rect 2533 2053 2547 2067
rect 2533 1973 2547 1987
rect 2453 1956 2467 1970
rect 2413 1893 2427 1907
rect 2533 1893 2547 1907
rect 2293 1853 2307 1867
rect 2333 1773 2347 1787
rect 2173 1733 2187 1747
rect 2213 1734 2227 1748
rect 1873 1690 1887 1704
rect 1973 1690 1987 1704
rect 1833 1513 1847 1527
rect 1953 1513 1967 1527
rect 1853 1473 1867 1487
rect 1753 1434 1767 1448
rect 1793 1434 1807 1448
rect 1833 1433 1847 1447
rect 1773 1392 1787 1406
rect 1733 1253 1747 1267
rect 2093 1692 2107 1706
rect 2133 1692 2147 1706
rect 2113 1453 2127 1467
rect 1873 1434 1887 1448
rect 1913 1434 1927 1448
rect 1953 1434 1967 1448
rect 2012 1434 2026 1448
rect 2033 1434 2047 1448
rect 2073 1434 2087 1448
rect 1873 1393 1887 1407
rect 1873 1372 1887 1386
rect 1853 1333 1867 1347
rect 1793 1214 1807 1228
rect 1833 1214 1847 1228
rect 1733 1172 1747 1186
rect 1773 1172 1787 1186
rect 1793 1153 1807 1167
rect 1793 1093 1807 1107
rect 1733 953 1747 967
rect 1973 1392 1987 1406
rect 2013 1393 2027 1407
rect 1933 1333 1947 1347
rect 1893 1213 1907 1227
rect 1933 1214 1947 1228
rect 1973 1214 1987 1228
rect 1873 1153 1887 1167
rect 1993 1153 2007 1167
rect 2433 1690 2447 1704
rect 2493 1653 2507 1667
rect 2453 1593 2467 1607
rect 2533 1593 2547 1607
rect 2373 1573 2387 1587
rect 2193 1453 2207 1467
rect 2233 1453 2247 1467
rect 2093 1392 2107 1406
rect 2173 1392 2187 1406
rect 2093 1293 2107 1307
rect 2133 1293 2147 1307
rect 2053 1273 2067 1287
rect 2253 1434 2267 1448
rect 2333 1433 2347 1447
rect 2373 1434 2387 1448
rect 2433 1433 2447 1447
rect 2233 1392 2247 1406
rect 2273 1392 2287 1406
rect 2813 3033 2827 3047
rect 2733 3013 2747 3027
rect 2713 2953 2727 2967
rect 2853 3133 2867 3147
rect 2833 2853 2847 2867
rect 2833 2832 2847 2846
rect 2733 2773 2747 2787
rect 2793 2774 2807 2788
rect 2913 3093 2927 3107
rect 2933 2950 2947 2964
rect 2873 2893 2887 2907
rect 2953 2833 2967 2847
rect 2933 2813 2947 2827
rect 2993 2950 3007 2964
rect 3153 3213 3167 3227
rect 3273 3373 3287 3387
rect 3273 3296 3287 3310
rect 3293 3173 3307 3187
rect 3293 3113 3307 3127
rect 3333 3413 3347 3427
rect 3333 3373 3347 3387
rect 3373 3573 3387 3587
rect 3373 3513 3387 3527
rect 3653 4353 3667 4367
rect 3613 4334 3627 4348
rect 3553 4293 3567 4307
rect 3593 4292 3607 4306
rect 3533 4253 3547 4267
rect 3533 4232 3547 4246
rect 3513 4193 3527 4207
rect 3513 3973 3527 3987
rect 3713 4493 3727 4507
rect 3753 4493 3767 4507
rect 3693 4453 3707 4467
rect 3693 4393 3707 4407
rect 3673 4293 3687 4307
rect 3613 4273 3627 4287
rect 3653 4273 3667 4287
rect 3593 4193 3607 4207
rect 3573 4053 3587 4067
rect 3673 4153 3687 4167
rect 3813 4793 3827 4807
rect 3813 4753 3827 4767
rect 3813 4653 3827 4667
rect 3853 4953 3867 4967
rect 3973 5093 3987 5107
rect 4113 5293 4127 5307
rect 4313 5673 4327 5687
rect 4233 5613 4247 5627
rect 4273 5613 4287 5627
rect 4193 5594 4207 5608
rect 4153 5553 4167 5567
rect 4193 5513 4207 5527
rect 4173 5493 4187 5507
rect 4153 5393 4167 5407
rect 4213 5393 4227 5407
rect 4233 5374 4247 5388
rect 4293 5374 4307 5388
rect 4213 5332 4227 5346
rect 4293 5333 4307 5347
rect 4253 5293 4267 5307
rect 4132 5273 4146 5287
rect 4153 5273 4167 5287
rect 4253 5272 4267 5286
rect 4093 5193 4107 5207
rect 4233 5173 4247 5187
rect 4053 5133 4067 5147
rect 3993 5032 4007 5046
rect 3993 4993 4007 5007
rect 3933 4933 3947 4947
rect 3913 4893 3927 4907
rect 3973 4893 3987 4907
rect 3973 4853 3987 4867
rect 3853 4813 3867 4827
rect 4073 5093 4087 5107
rect 4113 5074 4127 5088
rect 4153 5074 4167 5088
rect 4213 5074 4227 5088
rect 4073 4993 4087 5007
rect 4053 4973 4067 4987
rect 4033 4953 4047 4967
rect 4033 4913 4047 4927
rect 4073 4913 4087 4927
rect 4013 4812 4027 4826
rect 4053 4812 4067 4826
rect 4093 4812 4107 4826
rect 4173 4993 4187 5007
rect 4153 4933 4167 4947
rect 3933 4713 3947 4727
rect 3993 4713 4007 4727
rect 3893 4693 3907 4707
rect 3913 4673 3927 4687
rect 3833 4613 3847 4627
rect 3893 4613 3907 4627
rect 3833 4554 3847 4568
rect 3873 4554 3887 4568
rect 3773 4393 3787 4407
rect 3733 4353 3747 4367
rect 3753 4292 3767 4306
rect 3693 4133 3707 4147
rect 3653 4113 3667 4127
rect 3733 4073 3747 4087
rect 3673 4036 3687 4050
rect 3873 4493 3887 4507
rect 3853 4473 3867 4487
rect 3813 4413 3827 4427
rect 3833 4373 3847 4387
rect 3813 4353 3827 4367
rect 3913 4493 3927 4507
rect 3893 4473 3907 4487
rect 4053 4753 4067 4767
rect 4013 4693 4027 4707
rect 4073 4713 4087 4727
rect 4053 4613 4067 4627
rect 3973 4593 3987 4607
rect 4033 4554 4047 4568
rect 3933 4433 3947 4447
rect 3913 4334 3927 4348
rect 3813 4292 3827 4306
rect 3853 4292 3867 4306
rect 3893 4233 3907 4247
rect 3933 4233 3947 4247
rect 3833 4193 3847 4207
rect 3893 4153 3907 4167
rect 3793 4093 3807 4107
rect 3793 4033 3807 4047
rect 3773 4013 3787 4027
rect 3533 3953 3547 3967
rect 3593 3992 3607 4006
rect 3733 3973 3747 3987
rect 3633 3913 3647 3927
rect 3553 3893 3567 3907
rect 3613 3853 3627 3867
rect 3513 3813 3527 3827
rect 3573 3814 3587 3828
rect 3753 3893 3767 3907
rect 3733 3813 3747 3827
rect 3513 3772 3527 3786
rect 3553 3772 3567 3786
rect 3693 3773 3707 3787
rect 3733 3773 3747 3787
rect 3593 3733 3607 3747
rect 3653 3733 3667 3747
rect 3733 3733 3747 3747
rect 3553 3713 3567 3727
rect 3472 3673 3486 3687
rect 3493 3673 3507 3687
rect 3593 3712 3607 3726
rect 3553 3593 3567 3607
rect 3473 3573 3487 3587
rect 3453 3553 3467 3567
rect 3493 3553 3507 3567
rect 3553 3553 3567 3567
rect 3493 3516 3507 3530
rect 3613 3673 3627 3687
rect 3593 3493 3607 3507
rect 3413 3472 3427 3486
rect 3453 3472 3467 3486
rect 3593 3472 3607 3486
rect 3373 3413 3387 3427
rect 3353 3293 3367 3307
rect 3413 3373 3427 3387
rect 3493 3373 3507 3387
rect 3553 3373 3567 3387
rect 3473 3353 3487 3367
rect 3353 3253 3367 3267
rect 3333 3213 3347 3227
rect 3393 3252 3407 3266
rect 3433 3213 3447 3227
rect 3353 3153 3367 3167
rect 3313 3073 3327 3087
rect 3373 3073 3387 3087
rect 3353 3053 3367 3067
rect 3073 3033 3087 3047
rect 3173 3033 3187 3047
rect 3213 3033 3227 3047
rect 3313 3033 3327 3047
rect 3113 2996 3127 3010
rect 3213 2993 3227 3007
rect 3053 2853 3067 2867
rect 3253 2913 3267 2927
rect 3233 2893 3247 2907
rect 3133 2833 3147 2847
rect 3213 2833 3227 2847
rect 2973 2793 2987 2807
rect 2853 2773 2867 2787
rect 2953 2773 2967 2787
rect 2713 2732 2727 2746
rect 2813 2732 2827 2746
rect 2833 2713 2847 2727
rect 2873 2713 2887 2727
rect 2773 2693 2787 2707
rect 2733 2653 2747 2667
rect 2933 2653 2947 2667
rect 2993 2773 3007 2787
rect 3053 2776 3067 2790
rect 3093 2776 3107 2790
rect 2833 2533 2847 2547
rect 2733 2476 2747 2490
rect 2793 2476 2807 2490
rect 2853 2476 2867 2490
rect 2913 2476 2927 2490
rect 2813 2433 2827 2447
rect 2733 2413 2747 2427
rect 2693 2333 2707 2347
rect 2693 2254 2707 2268
rect 2813 2313 2827 2327
rect 2773 2254 2787 2268
rect 2833 2254 2847 2268
rect 2973 2633 2987 2647
rect 3213 2793 3227 2807
rect 3233 2773 3247 2787
rect 3133 2733 3147 2747
rect 3173 2732 3187 2746
rect 3093 2673 3107 2687
rect 2673 2133 2687 2147
rect 2753 2212 2767 2226
rect 2833 2153 2847 2167
rect 3353 2813 3367 2827
rect 3273 2793 3287 2807
rect 3313 2774 3327 2788
rect 3353 2773 3367 2787
rect 3293 2732 3307 2746
rect 3333 2713 3347 2727
rect 3253 2533 3267 2547
rect 3293 2533 3307 2547
rect 3073 2476 3087 2490
rect 3033 2430 3047 2444
rect 3153 2474 3167 2488
rect 3333 2474 3347 2488
rect 3413 2994 3427 3008
rect 3393 2853 3407 2867
rect 3393 2732 3407 2746
rect 3393 2653 3407 2667
rect 3373 2473 3387 2487
rect 3113 2430 3127 2444
rect 3073 2393 3087 2407
rect 3093 2333 3107 2347
rect 3013 2273 3027 2287
rect 2993 2213 3007 2227
rect 2973 2153 2987 2167
rect 2913 2133 2927 2147
rect 2693 2113 2707 2127
rect 2793 2113 2807 2127
rect 2893 2113 2907 2127
rect 2653 2013 2667 2027
rect 2573 1953 2587 1967
rect 2953 2013 2967 2027
rect 2693 1954 2707 1968
rect 2813 1954 2827 1968
rect 2633 1912 2647 1926
rect 2573 1853 2587 1867
rect 2613 1736 2627 1750
rect 2853 1813 2867 1827
rect 2793 1793 2807 1807
rect 2773 1773 2787 1787
rect 2793 1753 2807 1767
rect 2713 1734 2727 1748
rect 2773 1734 2787 1748
rect 2733 1692 2747 1706
rect 2673 1593 2687 1607
rect 2553 1573 2567 1587
rect 2593 1573 2607 1587
rect 2493 1434 2507 1448
rect 2553 1434 2567 1448
rect 2393 1392 2407 1406
rect 2432 1392 2446 1406
rect 2453 1393 2467 1407
rect 2533 1393 2547 1407
rect 2513 1333 2527 1347
rect 2333 1293 2347 1307
rect 2413 1293 2427 1307
rect 2393 1273 2407 1287
rect 2193 1233 2207 1247
rect 2353 1233 2367 1247
rect 2133 1214 2147 1228
rect 2173 1214 2187 1228
rect 2113 1172 2127 1186
rect 2393 1213 2407 1227
rect 2433 1273 2447 1287
rect 2453 1214 2467 1228
rect 2353 1172 2367 1186
rect 2433 1172 2447 1186
rect 2473 1172 2487 1186
rect 2513 1172 2527 1186
rect 1833 1133 1847 1147
rect 2033 1133 2047 1147
rect 2113 1133 2127 1147
rect 2173 1133 2187 1147
rect 1813 1073 1827 1087
rect 1833 1033 1847 1047
rect 2093 1013 2107 1027
rect 1973 953 1987 967
rect 1793 914 1807 928
rect 1733 872 1747 886
rect 1813 872 1827 886
rect 1893 913 1907 927
rect 1933 914 1947 928
rect 1953 872 1967 886
rect 1913 853 1927 867
rect 1893 833 1907 847
rect 1873 793 1887 807
rect 1993 833 2007 847
rect 2013 793 2027 807
rect 2053 793 2067 807
rect 2093 793 2107 807
rect 1913 773 1927 787
rect 1853 753 1867 767
rect 1753 694 1767 708
rect 1793 694 1807 708
rect 1773 652 1787 666
rect 1833 653 1847 667
rect 1813 633 1827 647
rect 1793 613 1807 627
rect 2653 1434 2667 1448
rect 2713 1434 2727 1448
rect 2693 1392 2707 1406
rect 2553 1373 2567 1387
rect 2593 1373 2607 1387
rect 2293 1073 2307 1087
rect 2533 1073 2547 1087
rect 2733 1273 2747 1287
rect 2673 1233 2687 1247
rect 2613 1214 2627 1228
rect 2653 1214 2667 1228
rect 2593 1133 2607 1147
rect 2653 1133 2667 1147
rect 2453 1053 2467 1067
rect 2553 1053 2567 1067
rect 2613 1053 2627 1067
rect 2453 993 2467 1007
rect 2273 973 2287 987
rect 2153 916 2167 930
rect 2213 916 2227 930
rect 2413 953 2427 967
rect 2293 913 2307 927
rect 2333 914 2347 928
rect 2233 873 2247 887
rect 2273 873 2287 887
rect 2113 773 2127 787
rect 2213 733 2227 747
rect 2213 693 2227 707
rect 2273 793 2287 807
rect 2373 833 2387 847
rect 2293 773 2307 787
rect 2313 733 2327 747
rect 2293 713 2307 727
rect 2353 694 2367 708
rect 2393 694 2407 708
rect 1933 652 1947 666
rect 2053 652 2067 666
rect 2113 650 2127 664
rect 2193 653 2207 667
rect 2233 653 2247 667
rect 1853 633 1867 647
rect 2113 613 2127 627
rect 1733 593 1747 607
rect 1713 393 1727 407
rect 1813 533 1827 547
rect 1993 533 2007 547
rect 1913 394 1927 408
rect 1773 253 1787 267
rect 1693 233 1707 247
rect 1713 174 1727 188
rect 1593 132 1607 146
rect 1633 133 1647 147
rect 1893 312 1907 326
rect 1892 253 1906 267
rect 1913 253 1927 267
rect 1853 213 1867 227
rect 1833 193 1847 207
rect 1793 173 1807 187
rect 2073 433 2087 447
rect 2033 394 2047 408
rect 2293 652 2307 666
rect 2193 533 2207 547
rect 2193 394 2207 408
rect 2233 394 2247 408
rect 2453 914 2467 928
rect 2493 914 2507 928
rect 2533 914 2547 928
rect 2473 872 2487 886
rect 2473 713 2487 727
rect 2433 694 2447 708
rect 2473 694 2487 708
rect 2513 694 2527 708
rect 2873 1734 2887 1748
rect 2933 1734 2947 1748
rect 2853 1692 2867 1706
rect 2893 1692 2907 1706
rect 3053 2133 3067 2147
rect 3113 2273 3127 2287
rect 3113 2213 3127 2227
rect 3173 2432 3187 2446
rect 3313 2432 3327 2446
rect 3373 2433 3387 2447
rect 3353 2393 3367 2407
rect 3193 2353 3207 2367
rect 3173 2333 3187 2347
rect 3313 2313 3327 2327
rect 3273 2293 3287 2307
rect 3353 2254 3367 2268
rect 3433 2933 3447 2947
rect 3493 3333 3507 3347
rect 3493 3312 3507 3326
rect 3553 3294 3567 3308
rect 3513 3253 3527 3267
rect 3493 3113 3507 3127
rect 3473 2893 3487 2907
rect 3473 2833 3487 2847
rect 3493 2813 3507 2827
rect 3533 3233 3547 3247
rect 3733 3513 3747 3527
rect 3913 4113 3927 4127
rect 3853 3990 3867 4004
rect 3793 3913 3807 3927
rect 3833 3816 3847 3830
rect 3893 3873 3907 3887
rect 3893 3833 3907 3847
rect 4013 4512 4027 4526
rect 4033 4493 4047 4507
rect 4033 4373 4047 4387
rect 4093 4693 4107 4707
rect 4033 4333 4047 4347
rect 4073 4333 4087 4347
rect 3993 4293 4007 4307
rect 3973 4253 3987 4267
rect 4033 4293 4047 4307
rect 4073 4293 4087 4307
rect 4013 4253 4027 4267
rect 3993 4113 4007 4127
rect 4053 4173 4067 4187
rect 3973 4073 3987 4087
rect 4033 4073 4047 4087
rect 4013 4034 4027 4048
rect 3933 3933 3947 3947
rect 3993 3992 4007 4006
rect 3953 3913 3967 3927
rect 3933 3814 3947 3828
rect 4213 4913 4227 4927
rect 4433 5852 4447 5866
rect 4473 5852 4487 5866
rect 4513 5852 4527 5866
rect 4553 5852 4567 5866
rect 4393 5833 4407 5847
rect 4553 5813 4567 5827
rect 4613 5933 4627 5947
rect 4593 5793 4607 5807
rect 4393 5733 4407 5747
rect 4573 5733 4587 5747
rect 4693 5913 4707 5927
rect 4673 5894 4687 5908
rect 4713 5893 4727 5907
rect 4733 5852 4747 5866
rect 4693 5833 4707 5847
rect 4612 5673 4626 5687
rect 4633 5673 4647 5687
rect 4453 5613 4467 5627
rect 4573 5613 4587 5627
rect 4613 5613 4627 5627
rect 4433 5573 4447 5587
rect 4533 5594 4547 5608
rect 4653 5594 4667 5608
rect 4373 5552 4387 5566
rect 4453 5553 4467 5567
rect 4513 5552 4527 5566
rect 4573 5553 4587 5567
rect 4593 5513 4607 5527
rect 4673 5553 4687 5567
rect 4633 5493 4647 5507
rect 4653 5473 4667 5487
rect 4593 5453 4607 5467
rect 4613 5433 4627 5447
rect 4353 5413 4367 5427
rect 4353 5374 4367 5388
rect 4393 5374 4407 5388
rect 4453 5373 4467 5387
rect 4513 5374 4527 5388
rect 4553 5374 4567 5388
rect 4593 5373 4607 5387
rect 4373 5332 4387 5346
rect 4413 5313 4427 5327
rect 4333 5253 4347 5267
rect 4313 5173 4327 5187
rect 4333 5073 4347 5087
rect 4273 5033 4287 5047
rect 4313 5032 4327 5046
rect 4273 4953 4287 4967
rect 4253 4933 4267 4947
rect 4453 5293 4467 5307
rect 4413 5253 4427 5267
rect 4453 5213 4467 5227
rect 4373 5073 4387 5087
rect 4413 5074 4427 5088
rect 4393 5033 4407 5047
rect 4373 4993 4387 5007
rect 4313 4873 4327 4887
rect 4353 4873 4367 4887
rect 4433 4953 4447 4967
rect 4453 4913 4467 4927
rect 4233 4854 4247 4868
rect 4213 4812 4227 4826
rect 4253 4773 4267 4787
rect 4153 4713 4167 4727
rect 4213 4713 4227 4727
rect 4153 4692 4167 4706
rect 4213 4613 4227 4627
rect 4153 4554 4167 4568
rect 4113 4513 4127 4527
rect 4233 4513 4247 4527
rect 4173 4493 4187 4507
rect 4153 4413 4167 4427
rect 4113 4353 4127 4367
rect 4193 4353 4207 4367
rect 4273 4633 4287 4647
rect 4433 4854 4447 4868
rect 4353 4812 4367 4826
rect 4373 4713 4387 4727
rect 4392 4693 4406 4707
rect 4413 4693 4427 4707
rect 4313 4593 4327 4607
rect 4353 4593 4367 4607
rect 4273 4553 4287 4567
rect 4353 4553 4367 4567
rect 4293 4512 4307 4526
rect 4253 4493 4267 4507
rect 4353 4513 4367 4527
rect 4333 4473 4347 4487
rect 4273 4453 4287 4467
rect 4253 4353 4267 4367
rect 4233 4333 4247 4347
rect 4113 4313 4127 4327
rect 4253 4313 4267 4327
rect 4173 4292 4187 4306
rect 4253 4253 4267 4267
rect 4353 4393 4367 4407
rect 4293 4293 4307 4307
rect 4353 4292 4367 4306
rect 4313 4253 4327 4267
rect 4273 4193 4287 4207
rect 4213 4173 4227 4187
rect 4353 4193 4367 4207
rect 4093 4153 4107 4167
rect 4313 4153 4327 4167
rect 4233 4133 4247 4147
rect 4153 4113 4167 4127
rect 4213 4113 4227 4127
rect 4193 4034 4207 4048
rect 4073 3993 4087 4007
rect 4113 3953 4127 3967
rect 4053 3833 4067 3847
rect 3893 3772 3907 3786
rect 3853 3753 3867 3767
rect 3773 3733 3787 3747
rect 3853 3593 3867 3607
rect 3793 3514 3807 3528
rect 3673 3470 3687 3484
rect 3713 3470 3727 3484
rect 3653 3333 3667 3347
rect 3713 3293 3727 3307
rect 3613 3213 3627 3227
rect 3633 3153 3647 3167
rect 3693 3153 3707 3167
rect 3593 3073 3607 3087
rect 3533 3053 3547 3067
rect 3613 3053 3627 3067
rect 3553 2994 3567 3008
rect 3713 3133 3727 3147
rect 3673 3093 3687 3107
rect 3633 3013 3647 3027
rect 3513 2774 3527 2788
rect 3633 2933 3647 2947
rect 3593 2893 3607 2907
rect 3633 2833 3647 2847
rect 3553 2773 3567 2787
rect 3593 2774 3607 2788
rect 3753 3413 3767 3427
rect 3813 3472 3827 3486
rect 3873 3413 3887 3427
rect 3773 3373 3787 3387
rect 3773 3333 3787 3347
rect 3753 3233 3767 3247
rect 3733 3093 3747 3107
rect 3953 3772 3967 3786
rect 3913 3593 3927 3607
rect 4073 3814 4087 3828
rect 4053 3713 4067 3727
rect 4013 3532 4027 3546
rect 3973 3393 3987 3407
rect 3933 3373 3947 3387
rect 3933 3352 3947 3366
rect 3973 3353 3987 3367
rect 4033 3353 4047 3367
rect 3913 3333 3927 3347
rect 3953 3333 3967 3347
rect 3833 3294 3847 3308
rect 3873 3293 3887 3307
rect 3893 3273 3907 3287
rect 3853 3233 3867 3247
rect 4013 3294 4027 3308
rect 3813 3213 3827 3227
rect 3913 3212 3927 3226
rect 3813 3113 3827 3127
rect 3893 3113 3907 3127
rect 3793 3073 3807 3087
rect 3713 3053 3727 3067
rect 3773 3053 3787 3067
rect 3733 2994 3747 3008
rect 3853 3053 3867 3067
rect 3713 2933 3727 2947
rect 3753 2933 3767 2947
rect 3793 2933 3807 2947
rect 3693 2773 3707 2787
rect 3493 2732 3507 2746
rect 3413 2593 3427 2607
rect 3413 2533 3427 2547
rect 3393 2313 3407 2327
rect 3193 2193 3207 2207
rect 3333 2212 3347 2226
rect 3393 2212 3407 2226
rect 3293 2193 3307 2207
rect 3193 2153 3207 2167
rect 3133 2013 3147 2027
rect 3093 1993 3107 2007
rect 3153 1993 3167 2007
rect 3013 1973 3027 1987
rect 2993 1753 3007 1767
rect 3033 1953 3047 1967
rect 3113 1893 3127 1907
rect 3193 1954 3207 1968
rect 3313 1973 3327 1987
rect 3373 1956 3387 1970
rect 3173 1913 3187 1927
rect 3073 1873 3087 1887
rect 3153 1873 3167 1887
rect 3033 1773 3047 1787
rect 3253 1912 3267 1926
rect 3613 2732 3627 2746
rect 3453 2493 3467 2507
rect 3533 2493 3547 2507
rect 3433 2473 3447 2487
rect 3433 2373 3447 2387
rect 3493 2474 3507 2488
rect 3573 2693 3587 2707
rect 3653 2693 3667 2707
rect 3673 2593 3687 2607
rect 3593 2553 3607 2567
rect 3533 2432 3547 2446
rect 3553 2413 3567 2427
rect 3453 2313 3467 2327
rect 3433 2293 3447 2307
rect 3453 2254 3467 2268
rect 3613 2493 3627 2507
rect 3933 3113 3947 3127
rect 3913 3013 3927 3027
rect 4033 3253 4047 3267
rect 3993 3213 4007 3227
rect 3993 3093 4007 3107
rect 3933 2994 3947 3008
rect 3973 2993 3987 3007
rect 4013 2993 4027 3007
rect 3893 2893 3907 2907
rect 3833 2853 3847 2867
rect 3813 2833 3827 2847
rect 3793 2774 3807 2788
rect 3973 2933 3987 2947
rect 3953 2793 3967 2807
rect 3833 2774 3847 2788
rect 3713 2732 3727 2746
rect 3873 2773 3887 2787
rect 3933 2774 3947 2788
rect 3853 2653 3867 2667
rect 3833 2553 3847 2567
rect 3693 2493 3707 2507
rect 3613 2413 3627 2427
rect 3653 2413 3667 2427
rect 3593 2353 3607 2367
rect 3553 2253 3567 2267
rect 3613 2313 3627 2327
rect 3553 2232 3567 2246
rect 3213 1873 3227 1887
rect 3373 1873 3387 1887
rect 3413 1873 3427 1887
rect 3213 1813 3227 1827
rect 3193 1793 3207 1807
rect 3013 1733 3027 1747
rect 3173 1733 3187 1747
rect 2952 1692 2966 1706
rect 3013 1693 3027 1707
rect 2973 1673 2987 1687
rect 2933 1653 2947 1667
rect 2993 1653 3007 1667
rect 2893 1613 2907 1627
rect 2973 1593 2987 1607
rect 2893 1553 2907 1567
rect 2953 1493 2967 1507
rect 2893 1453 2907 1467
rect 2793 1433 2807 1447
rect 2833 1434 2847 1448
rect 2993 1453 3007 1467
rect 2773 1333 2787 1347
rect 2813 1333 2827 1347
rect 2753 1233 2767 1247
rect 2813 1273 2827 1287
rect 2753 1172 2767 1186
rect 2793 1073 2807 1087
rect 2713 1053 2727 1067
rect 2713 913 2727 927
rect 2753 914 2767 928
rect 2673 833 2687 847
rect 2713 773 2727 787
rect 2773 773 2787 787
rect 2613 733 2627 747
rect 2553 696 2567 710
rect 2413 613 2427 627
rect 2393 553 2407 567
rect 2493 652 2507 666
rect 2633 693 2647 707
rect 2633 653 2647 667
rect 2733 650 2747 664
rect 2773 650 2787 664
rect 2613 633 2627 647
rect 2673 633 2687 647
rect 2693 553 2707 567
rect 2433 473 2447 487
rect 2413 433 2427 447
rect 2393 393 2407 407
rect 2273 373 2287 387
rect 2173 352 2187 366
rect 2053 333 2067 347
rect 2113 333 2127 347
rect 2033 213 2047 227
rect 1993 193 2007 207
rect 1913 173 1927 187
rect 1693 132 1707 146
rect 1733 132 1747 146
rect 1773 132 1787 146
rect 2113 176 2127 190
rect 2313 352 2327 366
rect 2353 352 2367 366
rect 2273 333 2287 347
rect 2273 253 2287 267
rect 2273 213 2287 227
rect 2213 174 2227 188
rect 1873 132 1887 146
rect 1933 130 1947 144
rect 1993 130 2007 144
rect 2033 133 2047 147
rect 2353 333 2367 347
rect 2593 413 2607 427
rect 2473 394 2487 408
rect 2513 394 2527 408
rect 2413 353 2427 367
rect 2493 352 2507 366
rect 2573 333 2587 347
rect 2653 352 2667 366
rect 2953 1253 2967 1267
rect 2833 1233 2847 1247
rect 2873 1233 2887 1247
rect 2913 1214 2927 1228
rect 2833 1172 2847 1186
rect 2893 1133 2907 1147
rect 2873 1093 2887 1107
rect 2953 1053 2967 1067
rect 2913 973 2927 987
rect 2953 933 2967 947
rect 2893 872 2907 886
rect 2953 813 2967 827
rect 2853 733 2867 747
rect 2813 713 2827 727
rect 2813 692 2827 706
rect 2893 713 2907 727
rect 2953 694 2967 708
rect 2813 652 2827 666
rect 2873 652 2887 666
rect 2793 633 2807 647
rect 2913 633 2927 647
rect 2853 453 2867 467
rect 2773 413 2787 427
rect 2753 394 2767 408
rect 2793 394 2807 408
rect 2833 394 2847 408
rect 2693 333 2707 347
rect 2693 312 2707 326
rect 2653 273 2667 287
rect 2593 253 2607 267
rect 2633 253 2647 267
rect 2473 233 2487 247
rect 2533 233 2547 247
rect 2393 213 2407 227
rect 2313 174 2327 188
rect 2373 174 2387 188
rect 2413 176 2427 190
rect 2353 132 2367 146
rect 2473 132 2487 146
rect 2653 233 2667 247
rect 2773 333 2787 347
rect 2833 313 2847 327
rect 2733 233 2747 247
rect 2793 213 2807 227
rect 2733 174 2747 188
rect 2953 573 2967 587
rect 3093 1690 3107 1704
rect 3173 1693 3187 1707
rect 3093 1653 3107 1667
rect 3153 1653 3167 1667
rect 3193 1653 3207 1667
rect 3113 1593 3127 1607
rect 3173 1593 3187 1607
rect 3033 1533 3047 1547
rect 3073 1390 3087 1404
rect 3093 1353 3107 1367
rect 3013 1273 3027 1287
rect 3013 1252 3027 1266
rect 3033 1172 3047 1186
rect 3093 1173 3107 1187
rect 3133 1533 3147 1547
rect 3273 1753 3287 1767
rect 3313 1753 3327 1767
rect 3473 2193 3487 2207
rect 3653 2254 3667 2268
rect 3713 2353 3727 2367
rect 3773 2472 3787 2486
rect 3833 2474 3847 2488
rect 3993 2733 4007 2747
rect 3953 2713 3967 2727
rect 3913 2573 3927 2587
rect 3933 2533 3947 2547
rect 3573 2212 3587 2226
rect 3633 2212 3647 2226
rect 3673 2212 3687 2226
rect 3713 2213 3727 2227
rect 3653 2193 3667 2207
rect 3593 2173 3607 2187
rect 3673 1993 3687 2007
rect 3613 1954 3627 1968
rect 3493 1893 3507 1907
rect 3433 1853 3447 1867
rect 3413 1793 3427 1807
rect 3333 1734 3347 1748
rect 3373 1734 3387 1748
rect 3313 1633 3327 1647
rect 3473 1733 3487 1747
rect 3693 1913 3707 1927
rect 3633 1853 3647 1867
rect 3813 2432 3827 2446
rect 3813 2333 3827 2347
rect 3893 2393 3907 2407
rect 3793 2212 3807 2226
rect 3753 2193 3767 2207
rect 3833 2173 3847 2187
rect 3793 2153 3807 2167
rect 3913 2313 3927 2327
rect 4173 3992 4187 4006
rect 4193 3973 4207 3987
rect 4173 3953 4187 3967
rect 4252 4073 4266 4087
rect 4273 4073 4287 4087
rect 4593 5332 4607 5346
rect 4533 5313 4547 5327
rect 4513 5133 4527 5147
rect 4553 5113 4567 5127
rect 4553 5074 4567 5088
rect 4473 4873 4487 4887
rect 4533 4993 4547 5007
rect 4593 5013 4607 5027
rect 4573 4973 4587 4987
rect 4593 4953 4607 4967
rect 4793 5973 4807 5987
rect 4873 5973 4887 5987
rect 5193 5953 5207 5967
rect 4833 5933 4847 5947
rect 4873 5894 4887 5908
rect 4933 5893 4947 5907
rect 4993 5894 5007 5908
rect 5033 5894 5047 5908
rect 5093 5894 5107 5908
rect 5153 5894 5167 5908
rect 5473 5933 5487 5947
rect 5913 5933 5927 5947
rect 5273 5894 5287 5908
rect 5333 5894 5347 5908
rect 5373 5894 5387 5908
rect 5413 5894 5427 5908
rect 4853 5852 4867 5866
rect 4913 5853 4927 5867
rect 4893 5833 4907 5847
rect 4872 5813 4886 5827
rect 4853 5773 4867 5787
rect 4733 5733 4747 5747
rect 4773 5733 4787 5747
rect 4713 5713 4727 5727
rect 4713 5673 4727 5687
rect 4713 5553 4727 5567
rect 4713 5532 4727 5546
rect 4693 5453 4707 5467
rect 4773 5693 4787 5707
rect 4833 5633 4847 5647
rect 4833 5594 4847 5608
rect 4893 5693 4907 5707
rect 5013 5852 5027 5866
rect 4993 5594 5007 5608
rect 5133 5852 5147 5866
rect 5173 5852 5187 5866
rect 5093 5793 5107 5807
rect 5153 5793 5167 5807
rect 5033 5594 5047 5608
rect 5073 5594 5087 5608
rect 5113 5594 5127 5608
rect 4733 5513 4747 5527
rect 4773 5513 4787 5527
rect 4753 5453 4767 5467
rect 4673 5433 4687 5447
rect 4713 5433 4727 5447
rect 4693 5413 4707 5427
rect 4673 5332 4687 5346
rect 4713 5332 4727 5346
rect 4633 5293 4647 5307
rect 4793 5433 4807 5447
rect 4893 5553 4907 5567
rect 4933 5552 4947 5566
rect 4993 5513 5007 5527
rect 5313 5852 5327 5866
rect 5273 5813 5287 5827
rect 5433 5852 5447 5866
rect 5293 5693 5307 5707
rect 5373 5693 5387 5707
rect 5253 5594 5267 5608
rect 5333 5633 5347 5647
rect 5653 5913 5667 5927
rect 5693 5913 5707 5927
rect 5493 5894 5507 5908
rect 5553 5894 5567 5908
rect 5593 5894 5607 5908
rect 5633 5893 5647 5907
rect 5573 5852 5587 5866
rect 5533 5813 5547 5827
rect 5493 5773 5507 5787
rect 5733 5894 5747 5908
rect 5813 5893 5827 5907
rect 5873 5894 5887 5908
rect 5573 5653 5587 5667
rect 5633 5653 5647 5667
rect 5393 5594 5407 5608
rect 5433 5594 5447 5608
rect 5473 5594 5487 5608
rect 5613 5594 5627 5608
rect 5093 5552 5107 5566
rect 5133 5552 5147 5566
rect 5173 5553 5187 5567
rect 5233 5552 5247 5566
rect 5273 5552 5287 5566
rect 5333 5553 5347 5567
rect 5033 5513 5047 5527
rect 4993 5453 5007 5467
rect 4973 5413 4987 5427
rect 4893 5374 4907 5388
rect 5113 5533 5127 5547
rect 5113 5413 5127 5427
rect 4833 5293 4847 5307
rect 4773 5273 4787 5287
rect 4973 5332 4987 5346
rect 5073 5332 5087 5346
rect 5413 5473 5427 5487
rect 5313 5453 5327 5467
rect 5213 5374 5227 5388
rect 5273 5374 5287 5388
rect 5593 5552 5607 5566
rect 5453 5433 5467 5447
rect 5413 5393 5427 5407
rect 5473 5393 5487 5407
rect 5353 5374 5367 5388
rect 5013 5293 5027 5307
rect 5053 5273 5067 5287
rect 4833 5233 4847 5247
rect 4873 5233 4887 5247
rect 4793 5173 4807 5187
rect 4753 5153 4767 5167
rect 4773 5133 4787 5147
rect 4713 5113 4727 5127
rect 4753 5093 4767 5107
rect 4653 5074 4667 5088
rect 4713 5074 4727 5088
rect 4633 5032 4647 5046
rect 4693 5032 4707 5046
rect 4733 5032 4747 5046
rect 4653 4993 4667 5007
rect 4993 5133 5007 5147
rect 4873 5093 4887 5107
rect 4833 5074 4847 5088
rect 4873 5074 4887 5088
rect 4953 5074 4967 5088
rect 5033 5074 5047 5088
rect 4933 5053 4947 5067
rect 4753 5013 4767 5027
rect 4853 5013 4867 5027
rect 4913 5013 4927 5027
rect 4733 4933 4747 4947
rect 4613 4913 4627 4927
rect 4713 4873 4727 4887
rect 4553 4854 4567 4868
rect 4613 4854 4627 4868
rect 4673 4854 4687 4868
rect 4573 4793 4587 4807
rect 4453 4773 4467 4787
rect 4533 4773 4547 4787
rect 4433 4593 4447 4607
rect 4453 4554 4467 4568
rect 4493 4554 4507 4568
rect 4573 4673 4587 4687
rect 4433 4512 4447 4526
rect 4473 4512 4487 4526
rect 4513 4512 4527 4526
rect 4413 4453 4427 4467
rect 4573 4512 4587 4526
rect 4552 4413 4566 4427
rect 4573 4413 4587 4427
rect 4513 4393 4527 4407
rect 4453 4353 4467 4367
rect 4413 4273 4427 4287
rect 4393 4253 4407 4267
rect 4373 4073 4387 4087
rect 4493 4273 4507 4287
rect 4493 4252 4507 4266
rect 4433 4213 4447 4227
rect 4453 4133 4467 4147
rect 4273 4034 4287 4048
rect 4313 4034 4327 4048
rect 4253 3973 4267 3987
rect 4313 3973 4327 3987
rect 4233 3953 4247 3967
rect 4293 3953 4307 3967
rect 4133 3933 4147 3947
rect 4213 3933 4227 3947
rect 4133 3853 4147 3867
rect 4153 3814 4167 3828
rect 4213 3814 4227 3828
rect 4112 3713 4126 3727
rect 4133 3713 4147 3727
rect 4073 3673 4087 3687
rect 4273 3813 4287 3827
rect 4413 4034 4427 4048
rect 4373 3993 4387 4007
rect 4473 3993 4487 4007
rect 4433 3973 4447 3987
rect 4473 3953 4487 3967
rect 4453 3933 4467 3947
rect 4393 3873 4407 3887
rect 4353 3833 4367 3847
rect 4333 3813 4347 3827
rect 4153 3653 4167 3667
rect 4233 3733 4247 3747
rect 4213 3673 4227 3687
rect 4193 3593 4207 3607
rect 4173 3553 4187 3567
rect 4133 3514 4147 3528
rect 4173 3514 4187 3528
rect 4113 3433 4127 3447
rect 4073 3353 4087 3367
rect 4093 3294 4107 3308
rect 4173 3393 4187 3407
rect 4193 3353 4207 3367
rect 4173 3293 4187 3307
rect 4173 3253 4187 3267
rect 4113 3213 4127 3227
rect 4173 3093 4187 3107
rect 4073 3053 4087 3067
rect 4053 3033 4067 3047
rect 4113 2994 4127 3008
rect 4333 3773 4347 3787
rect 4273 3553 4287 3567
rect 4273 3514 4287 3528
rect 4313 3513 4327 3527
rect 4253 3472 4267 3486
rect 4293 3473 4307 3487
rect 4233 3373 4247 3387
rect 4273 3353 4287 3367
rect 4233 3293 4247 3307
rect 4293 3313 4307 3327
rect 4373 3773 4387 3787
rect 4353 3733 4367 3747
rect 4353 3693 4367 3707
rect 4333 3413 4347 3427
rect 4333 3353 4347 3367
rect 4313 3294 4327 3308
rect 4253 3252 4267 3266
rect 4233 3233 4247 3247
rect 4333 3252 4347 3266
rect 4393 3533 4407 3547
rect 4433 3893 4447 3907
rect 4473 3893 4487 3907
rect 4693 4812 4707 4826
rect 4693 4793 4707 4807
rect 4653 4773 4667 4787
rect 4613 4673 4627 4687
rect 4733 4653 4747 4667
rect 4613 4633 4627 4647
rect 4653 4554 4667 4568
rect 4693 4554 4707 4568
rect 4613 4513 4627 4527
rect 4613 4473 4627 4487
rect 4713 4513 4727 4527
rect 4673 4473 4687 4487
rect 4693 4453 4707 4467
rect 4693 4432 4707 4446
rect 4613 4393 4627 4407
rect 4593 4353 4607 4367
rect 4533 4233 4547 4247
rect 4533 4193 4547 4207
rect 4613 4333 4627 4347
rect 4653 4334 4667 4348
rect 4693 4334 4707 4348
rect 4933 4973 4947 4987
rect 4913 4953 4927 4967
rect 4773 4933 4787 4947
rect 4853 4854 4867 4868
rect 4893 4854 4907 4868
rect 5013 5032 5027 5046
rect 5053 4993 5067 5007
rect 4953 4853 4967 4867
rect 4993 4854 5007 4868
rect 4833 4812 4847 4826
rect 4813 4753 4827 4767
rect 4772 4633 4786 4647
rect 4793 4633 4807 4647
rect 4833 4673 4847 4687
rect 4913 4813 4927 4827
rect 4913 4673 4927 4687
rect 4873 4653 4887 4667
rect 4913 4633 4927 4647
rect 5013 4793 5027 4807
rect 4833 4613 4847 4627
rect 4973 4613 4987 4627
rect 4993 4593 5007 4607
rect 4813 4573 4827 4587
rect 4833 4554 4847 4568
rect 4893 4554 4907 4568
rect 4953 4554 4967 4568
rect 4993 4554 5007 4568
rect 4813 4512 4827 4526
rect 4853 4512 4867 4526
rect 4753 4453 4767 4467
rect 4873 4453 4887 4467
rect 4733 4393 4747 4407
rect 4773 4373 4787 4387
rect 4813 4353 4827 4367
rect 4853 4353 4867 4367
rect 4593 4292 4607 4306
rect 4593 4253 4607 4267
rect 4673 4292 4687 4306
rect 4713 4293 4727 4307
rect 4633 4233 4647 4247
rect 4633 4113 4647 4127
rect 4593 4073 4607 4087
rect 4553 4053 4567 4067
rect 4533 4033 4547 4047
rect 4613 3993 4627 4007
rect 4553 3973 4567 3987
rect 4533 3953 4547 3967
rect 4513 3933 4527 3947
rect 4533 3893 4547 3907
rect 4493 3873 4507 3887
rect 4593 3873 4607 3887
rect 4493 3814 4507 3828
rect 4573 3814 4587 3828
rect 4493 3713 4507 3727
rect 4533 3713 4547 3727
rect 4433 3653 4447 3667
rect 4473 3653 4487 3667
rect 4373 3513 4387 3527
rect 4433 3514 4447 3528
rect 4433 3453 4447 3467
rect 4413 3413 4427 3427
rect 4433 3353 4447 3367
rect 4533 3653 4547 3667
rect 4493 3513 4507 3527
rect 4573 3733 4587 3747
rect 4573 3593 4587 3607
rect 4653 4093 4667 4107
rect 4693 4253 4707 4267
rect 4713 4233 4727 4247
rect 4713 4153 4727 4167
rect 4693 4113 4707 4127
rect 4753 4292 4767 4306
rect 4793 4292 4807 4306
rect 4813 4253 4827 4267
rect 4753 4133 4767 4147
rect 4793 4133 4807 4147
rect 4733 4034 4747 4048
rect 4853 4253 4867 4267
rect 4933 4512 4947 4526
rect 4973 4512 4987 4526
rect 4913 4373 4927 4387
rect 4893 4293 4907 4307
rect 5333 5332 5347 5346
rect 5273 5313 5287 5327
rect 5193 5273 5207 5287
rect 5193 5233 5207 5247
rect 5093 5153 5107 5167
rect 5393 5313 5407 5327
rect 5373 5233 5387 5247
rect 5373 5153 5387 5167
rect 5113 5074 5127 5088
rect 5153 5074 5167 5088
rect 5193 5074 5207 5088
rect 5093 5033 5107 5047
rect 5233 5073 5247 5087
rect 5273 5074 5287 5088
rect 5333 5074 5347 5088
rect 5113 5013 5127 5027
rect 5133 4973 5147 4987
rect 5153 4933 5167 4947
rect 5113 4854 5127 4868
rect 5313 5032 5327 5046
rect 5233 5013 5247 5027
rect 5193 4973 5207 4987
rect 5173 4913 5187 4927
rect 5073 4833 5087 4847
rect 5133 4773 5147 4787
rect 5513 5374 5527 5388
rect 5713 5813 5727 5827
rect 5753 5813 5767 5827
rect 5693 5493 5707 5507
rect 5673 5413 5687 5427
rect 5813 5614 5827 5628
rect 5813 5593 5827 5607
rect 5893 5593 5907 5607
rect 5753 5552 5767 5566
rect 5793 5552 5807 5566
rect 5793 5473 5807 5487
rect 5673 5374 5687 5388
rect 5493 5332 5507 5346
rect 5693 5332 5707 5346
rect 5833 5374 5847 5388
rect 5893 5374 5907 5388
rect 5653 5313 5667 5327
rect 5573 5273 5587 5287
rect 5413 5233 5427 5247
rect 5433 5074 5447 5088
rect 5473 5074 5487 5088
rect 5513 5074 5527 5088
rect 5553 5073 5567 5087
rect 5413 5032 5427 5046
rect 5453 5032 5467 5046
rect 5493 5032 5507 5046
rect 5553 5033 5567 5047
rect 5413 4993 5427 5007
rect 5453 4993 5467 5007
rect 5373 4953 5387 4967
rect 5213 4893 5227 4907
rect 5293 4893 5307 4907
rect 5413 4893 5427 4907
rect 5193 4793 5207 4807
rect 5073 4653 5087 4667
rect 5173 4653 5187 4667
rect 5053 4513 5067 4527
rect 5173 4613 5187 4627
rect 5133 4554 5147 4568
rect 5173 4554 5187 4568
rect 5033 4373 5047 4387
rect 4973 4353 4987 4367
rect 4993 4333 5007 4347
rect 5013 4292 5027 4306
rect 4993 4273 5007 4287
rect 4973 4252 4987 4266
rect 4953 4213 4967 4227
rect 4853 4193 4867 4207
rect 4933 4193 4947 4207
rect 4833 4133 4847 4147
rect 4893 4093 4907 4107
rect 4653 3992 4667 4006
rect 4633 3973 4647 3987
rect 4653 3873 4667 3887
rect 4692 3992 4706 4006
rect 4713 3993 4727 4007
rect 4713 3953 4727 3967
rect 4673 3853 4687 3867
rect 4653 3814 4667 3828
rect 4753 3893 4767 3907
rect 4873 4034 4887 4048
rect 4853 3992 4867 4006
rect 4893 3992 4907 4006
rect 4833 3953 4847 3967
rect 4813 3933 4827 3947
rect 4813 3873 4827 3887
rect 4893 3952 4907 3966
rect 4853 3913 4867 3927
rect 4633 3772 4647 3786
rect 4693 3772 4707 3786
rect 4813 3772 4827 3786
rect 4773 3733 4787 3747
rect 4833 3733 4847 3747
rect 4993 4233 5007 4247
rect 4973 4173 4987 4187
rect 4973 4152 4987 4166
rect 4953 4133 4967 4147
rect 4973 4073 4987 4087
rect 5033 4213 5047 4227
rect 5153 4493 5167 4507
rect 5253 4854 5267 4868
rect 5533 4953 5547 4967
rect 5493 4893 5507 4907
rect 5513 4854 5527 4868
rect 5353 4793 5367 4807
rect 5273 4753 5287 4767
rect 5293 4673 5307 4687
rect 5253 4573 5267 4587
rect 5373 4773 5387 4787
rect 5353 4573 5367 4587
rect 5273 4512 5287 4526
rect 5073 4453 5087 4467
rect 5113 4453 5127 4467
rect 5213 4453 5227 4467
rect 5433 4812 5447 4826
rect 5493 4813 5507 4827
rect 5393 4733 5407 4747
rect 5513 4673 5527 4687
rect 5433 4554 5447 4568
rect 5473 4554 5487 4568
rect 5513 4554 5527 4568
rect 5313 4493 5327 4507
rect 5353 4493 5367 4507
rect 5413 4493 5427 4507
rect 5153 4433 5167 4447
rect 5273 4433 5287 4447
rect 5073 4393 5087 4407
rect 5093 4373 5107 4387
rect 5113 4334 5127 4348
rect 5213 4373 5227 4387
rect 5273 4334 5287 4348
rect 5373 4433 5387 4447
rect 5353 4333 5367 4347
rect 5073 4293 5087 4307
rect 5053 4193 5067 4207
rect 5053 4172 5067 4186
rect 5213 4293 5227 4307
rect 5133 4233 5147 4247
rect 5113 4193 5127 4207
rect 5133 4133 5147 4147
rect 4993 4053 5007 4067
rect 5053 4053 5067 4067
rect 4953 3973 4967 3987
rect 4933 3953 4947 3967
rect 5033 3992 5047 4006
rect 5093 4093 5107 4107
rect 5092 4033 5106 4047
rect 5113 4033 5127 4047
rect 5173 4073 5187 4087
rect 5213 4034 5227 4048
rect 5253 4292 5267 4306
rect 5293 4193 5307 4207
rect 5253 4133 5267 4147
rect 4993 3933 5007 3947
rect 5073 3933 5087 3947
rect 4913 3893 4927 3907
rect 5013 3893 5027 3907
rect 5093 3893 5107 3907
rect 4913 3833 4927 3847
rect 4893 3813 4907 3827
rect 4953 3814 4967 3828
rect 4973 3753 4987 3767
rect 4933 3733 4947 3747
rect 4673 3713 4687 3727
rect 4773 3653 4787 3667
rect 4753 3633 4767 3647
rect 4673 3573 4687 3587
rect 4593 3553 4607 3567
rect 4633 3553 4647 3567
rect 4553 3533 4567 3547
rect 4493 3473 4507 3487
rect 4473 3333 4487 3347
rect 4413 3294 4427 3308
rect 4453 3294 4467 3308
rect 4233 3193 4247 3207
rect 4213 3173 4227 3187
rect 4333 3173 4347 3187
rect 4313 3093 4327 3107
rect 4053 2933 4067 2947
rect 4133 2933 4147 2947
rect 4093 2853 4107 2867
rect 4132 2853 4146 2867
rect 4153 2853 4167 2867
rect 4073 2793 4087 2807
rect 4033 2773 4047 2787
rect 4113 2793 4127 2807
rect 4133 2773 4147 2787
rect 4033 2733 4047 2747
rect 4093 2732 4107 2746
rect 4053 2693 4067 2707
rect 4113 2673 4127 2687
rect 4033 2633 4047 2647
rect 4113 2633 4127 2647
rect 4033 2533 4047 2547
rect 4013 2493 4027 2507
rect 3993 2474 4007 2488
rect 4273 2994 4287 3008
rect 4232 2953 4246 2967
rect 4253 2952 4267 2966
rect 4293 2953 4307 2967
rect 4313 2933 4327 2947
rect 4293 2893 4307 2907
rect 4193 2813 4207 2827
rect 4233 2774 4247 2788
rect 4173 2593 4187 2607
rect 4153 2573 4167 2587
rect 4433 3252 4447 3266
rect 4473 3193 4487 3207
rect 4393 3053 4407 3067
rect 4433 3033 4447 3047
rect 4352 2993 4366 3007
rect 4372 2993 4386 3007
rect 4393 2994 4407 3008
rect 4553 3472 4567 3486
rect 4713 3514 4727 3528
rect 4633 3472 4647 3486
rect 4673 3472 4687 3486
rect 4633 3413 4647 3427
rect 4673 3413 4687 3427
rect 4753 3413 4767 3427
rect 4993 3713 5007 3727
rect 4973 3693 4987 3707
rect 4993 3673 5007 3687
rect 4953 3653 4967 3667
rect 4873 3613 4887 3627
rect 4913 3613 4927 3627
rect 4793 3473 4807 3487
rect 4793 3433 4807 3447
rect 4613 3393 4627 3407
rect 4553 3373 4567 3387
rect 4513 3353 4527 3367
rect 4573 3353 4587 3367
rect 4653 3353 4667 3367
rect 4493 3133 4507 3147
rect 4633 3293 4647 3307
rect 4553 3252 4567 3266
rect 4593 3252 4607 3266
rect 4633 3252 4647 3266
rect 4773 3373 4787 3387
rect 4693 3353 4707 3367
rect 4713 3333 4727 3347
rect 4813 3333 4827 3347
rect 4753 3294 4767 3308
rect 4673 3253 4687 3267
rect 4733 3252 4747 3266
rect 4653 3193 4667 3207
rect 4613 3173 4627 3187
rect 4713 3173 4727 3187
rect 4513 3073 4527 3087
rect 4513 3033 4527 3047
rect 4573 3033 4587 3047
rect 4493 2994 4507 3008
rect 4413 2952 4427 2966
rect 4373 2853 4387 2867
rect 4353 2813 4367 2827
rect 4413 2813 4427 2827
rect 4293 2732 4307 2746
rect 4273 2693 4287 2707
rect 4233 2673 4247 2687
rect 4213 2553 4227 2567
rect 4113 2513 4127 2527
rect 4153 2513 4167 2527
rect 4093 2453 4107 2467
rect 3973 2432 3987 2446
rect 4093 2373 4107 2387
rect 4013 2313 4027 2327
rect 4073 2273 4087 2287
rect 3913 2093 3927 2107
rect 3893 2073 3907 2087
rect 3973 2053 3987 2067
rect 3933 1993 3947 2007
rect 3773 1954 3787 1968
rect 3833 1953 3847 1967
rect 3873 1954 3887 1968
rect 3933 1954 3947 1968
rect 3733 1912 3747 1926
rect 3793 1912 3807 1926
rect 3893 1893 3907 1907
rect 3833 1833 3847 1847
rect 4053 1954 4067 1968
rect 4033 1912 4047 1926
rect 4213 2493 4227 2507
rect 4133 2473 4147 2487
rect 4173 2474 4187 2488
rect 4153 2432 4167 2446
rect 4213 2432 4227 2446
rect 4213 2393 4227 2407
rect 4153 2273 4167 2287
rect 4173 2254 4187 2268
rect 4293 2653 4307 2667
rect 4373 2732 4387 2746
rect 4453 2933 4467 2947
rect 4493 2813 4507 2827
rect 4433 2793 4447 2807
rect 4533 2993 4547 3007
rect 4673 3113 4687 3127
rect 4652 3073 4666 3087
rect 4673 3073 4687 3087
rect 4773 3213 4787 3227
rect 4753 2994 4767 3008
rect 4593 2952 4607 2966
rect 4653 2952 4667 2966
rect 4693 2952 4707 2966
rect 4733 2913 4747 2927
rect 4593 2893 4607 2907
rect 4773 2853 4787 2867
rect 4533 2833 4547 2847
rect 4593 2813 4607 2827
rect 4533 2774 4547 2788
rect 4572 2773 4586 2787
rect 4593 2774 4607 2788
rect 4653 2774 4667 2788
rect 4693 2774 4707 2788
rect 4753 2774 4767 2788
rect 4433 2732 4447 2746
rect 4473 2732 4487 2746
rect 4553 2713 4567 2727
rect 4453 2693 4467 2707
rect 4513 2693 4527 2707
rect 4533 2613 4547 2627
rect 4393 2593 4407 2607
rect 4333 2533 4347 2547
rect 4333 2512 4347 2526
rect 4313 2493 4327 2507
rect 4233 2373 4247 2387
rect 4253 2253 4267 2267
rect 4113 2212 4127 2226
rect 4193 2212 4207 2226
rect 4153 2173 4167 2187
rect 4293 2413 4307 2427
rect 4353 2393 4367 2407
rect 4313 2353 4327 2367
rect 4353 2353 4367 2367
rect 4293 2333 4307 2347
rect 4313 2254 4327 2268
rect 4433 2513 4447 2527
rect 4473 2493 4487 2507
rect 4453 2393 4467 2407
rect 4633 2732 4647 2746
rect 4593 2693 4607 2707
rect 4673 2633 4687 2647
rect 4573 2613 4587 2627
rect 4713 2613 4727 2627
rect 4713 2553 4727 2567
rect 4793 2833 4807 2847
rect 4933 3533 4947 3547
rect 4953 3513 4967 3527
rect 5033 3873 5047 3887
rect 5073 3814 5087 3828
rect 5153 3953 5167 3967
rect 5133 3813 5147 3827
rect 5033 3733 5047 3747
rect 5033 3673 5047 3687
rect 5033 3613 5047 3627
rect 5013 3533 5027 3547
rect 5133 3773 5147 3787
rect 5113 3753 5127 3767
rect 5093 3733 5107 3747
rect 5133 3693 5147 3707
rect 5113 3673 5127 3687
rect 5113 3652 5127 3666
rect 5093 3633 5107 3647
rect 5073 3593 5087 3607
rect 5053 3573 5067 3587
rect 4953 3473 4967 3487
rect 4933 3413 4947 3427
rect 4933 3373 4947 3387
rect 4853 3294 4867 3308
rect 4893 3294 4907 3308
rect 5013 3433 5027 3447
rect 4993 3413 5007 3427
rect 4873 3252 4887 3266
rect 4913 3233 4927 3247
rect 4833 3133 4847 3147
rect 4853 3073 4867 3087
rect 4973 3133 4987 3147
rect 4913 3053 4927 3067
rect 4893 3033 4907 3047
rect 4833 2953 4847 2967
rect 4833 2833 4847 2847
rect 4913 2913 4927 2927
rect 4852 2793 4866 2807
rect 4873 2793 4887 2807
rect 4813 2773 4827 2787
rect 4953 3053 4967 3067
rect 4953 2953 4967 2967
rect 5013 3313 5027 3327
rect 4993 3093 5007 3107
rect 5053 3313 5067 3327
rect 5033 3293 5047 3307
rect 5113 3573 5127 3587
rect 5113 3514 5127 3528
rect 5233 3993 5247 4007
rect 5293 4113 5307 4127
rect 5293 4092 5307 4106
rect 5273 4073 5287 4087
rect 5313 4053 5327 4067
rect 5413 4393 5427 4407
rect 5493 4493 5507 4507
rect 5453 4353 5467 4367
rect 5453 4292 5467 4306
rect 5513 4473 5527 4487
rect 5653 5153 5667 5167
rect 5813 5332 5827 5346
rect 5853 5313 5867 5327
rect 5833 5233 5847 5247
rect 5673 5073 5687 5087
rect 5733 5074 5747 5088
rect 5693 5053 5707 5067
rect 5573 4993 5587 5007
rect 5553 4933 5567 4947
rect 5653 4933 5667 4947
rect 5593 4854 5607 4868
rect 5633 4854 5647 4868
rect 5673 4873 5687 4887
rect 5553 4713 5567 4727
rect 5613 4793 5627 4807
rect 5573 4613 5587 4627
rect 5613 4573 5627 4587
rect 5673 4553 5687 4567
rect 5593 4512 5607 4526
rect 5553 4493 5567 4507
rect 5613 4473 5627 4487
rect 5673 4513 5687 4527
rect 5633 4453 5647 4467
rect 5533 4433 5547 4447
rect 5613 4433 5627 4447
rect 5553 4413 5567 4427
rect 5513 4393 5527 4407
rect 5793 5032 5807 5046
rect 5713 5013 5727 5027
rect 5753 5013 5767 5027
rect 5773 4933 5787 4947
rect 5733 4893 5747 4907
rect 5853 5213 5867 5227
rect 5833 4853 5847 4867
rect 5793 4812 5807 4826
rect 5753 4773 5767 4787
rect 5733 4573 5747 4587
rect 5773 4554 5787 4568
rect 5833 4554 5847 4568
rect 5733 4493 5747 4507
rect 5693 4453 5707 4467
rect 5553 4373 5567 4387
rect 5533 4353 5547 4367
rect 5573 4334 5587 4348
rect 5513 4293 5527 4307
rect 5433 4253 5447 4267
rect 5493 4253 5507 4267
rect 5373 4213 5387 4227
rect 5373 4113 5387 4127
rect 5293 4033 5307 4047
rect 5353 4033 5367 4047
rect 5253 3953 5267 3967
rect 5193 3933 5207 3947
rect 5193 3893 5207 3907
rect 5233 3893 5247 3907
rect 5173 3833 5187 3847
rect 5173 3793 5187 3807
rect 5173 3713 5187 3727
rect 5213 3873 5227 3887
rect 5313 3992 5327 4006
rect 5353 3993 5367 4007
rect 5273 3853 5287 3867
rect 5333 3853 5347 3867
rect 5233 3833 5247 3847
rect 5313 3833 5327 3847
rect 5253 3814 5267 3828
rect 5293 3814 5307 3828
rect 5413 4093 5427 4107
rect 5393 4033 5407 4047
rect 5373 3893 5387 3907
rect 5373 3833 5387 3847
rect 5453 4113 5467 4127
rect 5433 4033 5447 4047
rect 5493 4053 5507 4067
rect 5573 4273 5587 4287
rect 5553 4253 5567 4267
rect 5633 4253 5647 4267
rect 5413 3973 5427 3987
rect 5513 3992 5527 4006
rect 5473 3933 5487 3947
rect 5512 3933 5526 3947
rect 5533 3933 5547 3947
rect 5593 4034 5607 4048
rect 5633 4034 5647 4048
rect 5673 4033 5687 4047
rect 5713 4413 5727 4427
rect 5713 4373 5727 4387
rect 5753 4453 5767 4467
rect 5793 4433 5807 4447
rect 5773 4334 5787 4348
rect 5833 4493 5847 4507
rect 5893 5213 5907 5227
rect 5953 5593 5967 5607
rect 5933 5413 5947 5427
rect 5973 5493 5987 5507
rect 5953 5033 5967 5047
rect 5973 4873 5987 4887
rect 5913 4713 5927 4727
rect 5873 4553 5887 4567
rect 5933 4554 5947 4568
rect 5873 4493 5887 4507
rect 5853 4433 5867 4447
rect 5953 4513 5967 4527
rect 5933 4493 5947 4507
rect 5893 4413 5907 4427
rect 5833 4334 5847 4348
rect 5893 4334 5907 4348
rect 5973 4373 5987 4387
rect 5733 4093 5747 4107
rect 5713 4033 5727 4047
rect 5573 3993 5587 4007
rect 5513 3893 5527 3907
rect 5453 3873 5467 3887
rect 5273 3772 5287 3786
rect 5213 3752 5227 3766
rect 5193 3693 5207 3707
rect 5153 3633 5167 3647
rect 5153 3593 5167 3607
rect 5233 3733 5247 3747
rect 5213 3633 5227 3647
rect 5393 3813 5407 3827
rect 5493 3853 5507 3867
rect 5553 3913 5567 3927
rect 5533 3852 5547 3866
rect 5513 3813 5527 3827
rect 5373 3753 5387 3767
rect 5353 3713 5367 3727
rect 5253 3673 5267 3687
rect 5273 3613 5287 3627
rect 5253 3593 5267 3607
rect 5173 3472 5187 3486
rect 5233 3473 5247 3487
rect 5193 3433 5207 3447
rect 5173 3413 5187 3427
rect 5133 3393 5147 3407
rect 5113 3353 5127 3367
rect 5093 3333 5107 3347
rect 5153 3313 5167 3327
rect 5133 3293 5147 3307
rect 5033 3253 5047 3267
rect 5133 3233 5147 3247
rect 5213 3413 5227 3427
rect 5173 3293 5187 3307
rect 5273 3573 5287 3587
rect 5293 3553 5307 3567
rect 5293 3514 5307 3528
rect 5333 3514 5347 3528
rect 5273 3472 5287 3486
rect 5353 3473 5367 3487
rect 5353 3393 5367 3407
rect 5433 3772 5447 3786
rect 5473 3753 5487 3767
rect 5653 3992 5667 4006
rect 5693 3993 5707 4007
rect 5613 3953 5627 3967
rect 5593 3913 5607 3927
rect 5593 3853 5607 3867
rect 5573 3833 5587 3847
rect 5633 3933 5647 3947
rect 5673 3853 5687 3867
rect 5633 3833 5647 3847
rect 5553 3773 5567 3787
rect 5413 3713 5427 3727
rect 5393 3673 5407 3687
rect 5393 3633 5407 3647
rect 5473 3633 5487 3647
rect 5413 3613 5427 3627
rect 5413 3553 5427 3567
rect 5393 3513 5407 3527
rect 5493 3593 5507 3607
rect 5493 3513 5507 3527
rect 5433 3473 5447 3487
rect 5393 3453 5407 3467
rect 5333 3373 5347 3387
rect 5373 3373 5387 3387
rect 5313 3333 5327 3347
rect 5173 3253 5187 3267
rect 5233 3252 5247 3266
rect 5173 3232 5187 3246
rect 5253 3233 5267 3247
rect 5053 3213 5067 3227
rect 5093 3213 5107 3227
rect 5033 3153 5047 3167
rect 5093 3153 5107 3167
rect 5053 3053 5067 3067
rect 5053 2994 5067 3008
rect 5033 2952 5047 2966
rect 5073 2873 5087 2887
rect 5193 3213 5207 3227
rect 5173 3173 5187 3187
rect 5233 3193 5247 3207
rect 5213 3173 5227 3187
rect 5153 3153 5167 3167
rect 5193 3153 5207 3167
rect 5213 3093 5227 3107
rect 5193 3073 5207 3087
rect 5213 2993 5227 3007
rect 5133 2953 5147 2967
rect 5113 2933 5127 2947
rect 4933 2853 4947 2867
rect 4973 2853 4987 2867
rect 5013 2813 5027 2827
rect 4933 2793 4947 2807
rect 4793 2732 4807 2746
rect 4773 2713 4787 2727
rect 4753 2633 4767 2647
rect 4733 2474 4747 2488
rect 4733 2413 4747 2427
rect 4653 2373 4667 2387
rect 4513 2273 4527 2287
rect 4473 2254 4487 2268
rect 4413 2233 4427 2247
rect 4133 2093 4147 2107
rect 4253 2093 4267 2107
rect 4113 1893 4127 1907
rect 4113 1833 4127 1847
rect 3993 1813 4007 1827
rect 3713 1793 3727 1807
rect 3873 1793 3887 1807
rect 3653 1773 3667 1787
rect 3693 1773 3707 1787
rect 3433 1692 3447 1706
rect 3473 1692 3487 1706
rect 3393 1673 3407 1687
rect 3333 1573 3347 1587
rect 3453 1593 3467 1607
rect 3393 1553 3407 1567
rect 3253 1493 3267 1507
rect 3213 1473 3227 1487
rect 3193 1434 3207 1448
rect 3173 1392 3187 1406
rect 3233 1393 3247 1407
rect 3213 1373 3227 1387
rect 3313 1434 3327 1448
rect 3293 1392 3307 1406
rect 3273 1353 3287 1367
rect 3373 1393 3387 1407
rect 3373 1353 3387 1367
rect 3453 1473 3467 1487
rect 3413 1453 3427 1467
rect 3253 1333 3267 1347
rect 3333 1333 3347 1347
rect 3393 1333 3407 1347
rect 3173 1313 3187 1327
rect 3133 1273 3147 1287
rect 3553 1734 3567 1748
rect 3573 1673 3587 1687
rect 3533 1653 3547 1667
rect 3713 1734 3727 1748
rect 3773 1733 3787 1747
rect 3693 1653 3707 1667
rect 3733 1593 3747 1607
rect 3433 1373 3447 1387
rect 3553 1390 3567 1404
rect 3473 1373 3487 1387
rect 3433 1333 3447 1347
rect 3413 1213 3427 1227
rect 3153 1172 3167 1186
rect 3113 1153 3127 1167
rect 3173 1153 3187 1167
rect 3153 1033 3167 1047
rect 3093 973 3107 987
rect 3053 933 3067 947
rect 3013 914 3027 928
rect 3093 913 3107 927
rect 3393 1170 3407 1184
rect 3393 1153 3407 1167
rect 3413 1093 3427 1107
rect 3353 1053 3367 1067
rect 3333 973 3347 987
rect 3193 916 3207 930
rect 3233 916 3247 930
rect 3293 916 3307 930
rect 3333 916 3347 930
rect 3033 833 3047 847
rect 3113 870 3127 884
rect 3173 873 3187 887
rect 3193 833 3207 847
rect 3053 733 3067 747
rect 3013 694 3027 708
rect 3173 813 3187 827
rect 3253 793 3267 807
rect 3333 793 3347 807
rect 3213 694 3227 708
rect 3033 652 3047 666
rect 3093 653 3107 667
rect 3153 613 3167 627
rect 3193 593 3207 607
rect 2973 553 2987 567
rect 3033 473 3047 487
rect 2953 453 2967 467
rect 2913 394 2927 408
rect 2973 393 2987 407
rect 3153 453 3167 467
rect 3133 413 3147 427
rect 3073 394 3087 408
rect 2853 253 2867 267
rect 2873 213 2887 227
rect 2833 173 2847 187
rect 2973 352 2987 366
rect 3013 352 3027 366
rect 3013 313 3027 327
rect 2893 193 2907 207
rect 2933 193 2947 207
rect 2533 130 2547 144
rect 2653 132 2667 146
rect 2713 132 2727 146
rect 2753 132 2767 146
rect 2793 132 2807 146
rect 2853 132 2867 146
rect 2893 132 2907 146
rect 1893 113 1907 127
rect 1513 33 1527 47
rect 1553 33 1567 47
rect 2953 176 2967 190
rect 3093 353 3107 367
rect 3093 313 3107 327
rect 3273 753 3287 767
rect 3313 753 3327 767
rect 3293 733 3307 747
rect 3313 652 3327 666
rect 3393 1033 3407 1047
rect 3493 1313 3507 1327
rect 3593 1313 3607 1327
rect 3453 1233 3467 1247
rect 3573 1273 3587 1287
rect 3533 1214 3547 1228
rect 3453 1173 3467 1187
rect 3513 1172 3527 1186
rect 3433 1053 3447 1067
rect 3653 1513 3667 1527
rect 3673 1473 3687 1487
rect 3733 1453 3747 1467
rect 3893 1692 3907 1706
rect 3893 1513 3907 1527
rect 3833 1493 3847 1507
rect 3813 1473 3827 1487
rect 3793 1433 3807 1447
rect 3853 1434 3867 1448
rect 3953 1773 3967 1787
rect 4073 1753 4087 1767
rect 4013 1734 4027 1748
rect 3953 1692 3967 1706
rect 3993 1692 4007 1706
rect 4033 1633 4047 1647
rect 3973 1593 3987 1607
rect 3933 1434 3947 1448
rect 3792 1390 3806 1404
rect 3813 1393 3827 1407
rect 3873 1353 3887 1367
rect 3933 1353 3947 1367
rect 3773 1293 3787 1307
rect 3853 1293 3867 1307
rect 3633 1273 3647 1287
rect 3833 1273 3847 1287
rect 3653 1253 3667 1267
rect 3593 1172 3607 1186
rect 3633 1172 3647 1186
rect 3673 1172 3687 1186
rect 3733 1153 3747 1167
rect 3793 1133 3807 1147
rect 3913 1216 3927 1230
rect 3853 1172 3867 1186
rect 3833 1033 3847 1047
rect 3513 1013 3527 1027
rect 3573 1013 3587 1027
rect 3433 973 3447 987
rect 3413 933 3427 947
rect 3473 914 3487 928
rect 3373 873 3387 887
rect 3413 872 3427 886
rect 3473 853 3487 867
rect 3433 694 3447 708
rect 3493 833 3507 847
rect 3353 473 3367 487
rect 3373 453 3387 467
rect 3253 413 3267 427
rect 3333 394 3347 408
rect 3153 352 3167 366
rect 3213 352 3227 366
rect 3353 352 3367 366
rect 3313 273 3327 287
rect 3053 213 3067 227
rect 3093 176 3107 190
rect 3173 213 3187 227
rect 3153 173 3167 187
rect 2953 133 2967 147
rect 2993 132 3007 146
rect 3373 174 3387 188
rect 3433 473 3447 487
rect 3413 173 3427 187
rect 3173 130 3187 144
rect 3213 130 3227 144
rect 3273 130 3287 144
rect 3353 133 3367 147
rect 3033 93 3047 107
rect 3033 33 3047 47
rect 3393 132 3407 146
rect 3593 914 3607 928
rect 3653 914 3667 928
rect 3693 914 3707 928
rect 3753 914 3767 928
rect 3793 914 3807 928
rect 3833 914 3847 928
rect 3633 853 3647 867
rect 3613 833 3627 847
rect 3553 694 3567 708
rect 3593 694 3607 708
rect 3873 913 3887 927
rect 3933 914 3947 928
rect 4173 2073 4187 2087
rect 4213 1954 4227 1968
rect 4273 1954 4287 1968
rect 4133 1793 4147 1807
rect 4213 1793 4227 1807
rect 4153 1753 4167 1767
rect 4173 1692 4187 1706
rect 4133 1653 4147 1667
rect 4213 1633 4227 1647
rect 4153 1493 4167 1507
rect 4013 1434 4027 1448
rect 4053 1434 4067 1448
rect 4033 1392 4047 1406
rect 4093 1393 4107 1407
rect 4073 1313 4087 1327
rect 4213 1434 4227 1448
rect 4253 1913 4267 1927
rect 4353 2193 4367 2207
rect 4333 2153 4347 2167
rect 4373 2173 4387 2187
rect 4353 2053 4367 2067
rect 4353 2013 4367 2027
rect 4313 1912 4327 1926
rect 4373 1912 4387 1926
rect 4493 2212 4507 2226
rect 4513 2173 4527 2187
rect 4453 2153 4467 2167
rect 4473 1954 4487 1968
rect 4413 1893 4427 1907
rect 4373 1873 4387 1887
rect 4293 1853 4307 1867
rect 4432 1853 4446 1867
rect 4453 1853 4467 1867
rect 4273 1833 4287 1847
rect 4373 1773 4387 1787
rect 4253 1693 4267 1707
rect 4253 1653 4267 1667
rect 4593 2353 4607 2367
rect 4713 2293 4727 2307
rect 4673 2254 4687 2268
rect 4773 2573 4787 2587
rect 4893 2732 4907 2746
rect 4953 2773 4967 2787
rect 5053 2793 5067 2807
rect 5093 2853 5107 2867
rect 5073 2773 5087 2787
rect 4933 2713 4947 2727
rect 4833 2693 4847 2707
rect 4913 2673 4927 2687
rect 4893 2633 4907 2647
rect 4793 2513 4807 2527
rect 4813 2474 4827 2488
rect 4853 2474 4867 2488
rect 4913 2533 4927 2547
rect 5073 2733 5087 2747
rect 5033 2713 5047 2727
rect 4992 2613 5006 2627
rect 5013 2613 5027 2627
rect 4953 2493 4967 2507
rect 4933 2474 4947 2488
rect 4973 2474 4987 2488
rect 5053 2493 5067 2507
rect 5033 2473 5047 2487
rect 4873 2413 4887 2427
rect 4793 2313 4807 2327
rect 4833 2313 4847 2327
rect 4773 2293 4787 2307
rect 4853 2293 4867 2307
rect 4833 2273 4847 2287
rect 4593 2212 4607 2226
rect 4693 2212 4707 2226
rect 4653 2153 4667 2167
rect 4693 2093 4707 2107
rect 4573 2073 4587 2087
rect 4693 1973 4707 1987
rect 4573 1954 4587 1968
rect 4613 1954 4627 1968
rect 4673 1954 4687 1968
rect 4533 1912 4547 1926
rect 4593 1912 4607 1926
rect 4573 1893 4587 1907
rect 4453 1832 4467 1846
rect 4513 1833 4527 1847
rect 4433 1553 4447 1567
rect 4353 1533 4367 1547
rect 4313 1493 4327 1507
rect 4113 1373 4127 1387
rect 4193 1373 4207 1387
rect 4213 1353 4227 1367
rect 4213 1313 4227 1327
rect 4093 1293 4107 1307
rect 4233 1293 4247 1307
rect 4273 1433 4287 1447
rect 4373 1434 4387 1448
rect 4433 1433 4447 1447
rect 4273 1333 4287 1347
rect 4293 1313 4307 1327
rect 4073 1273 4087 1287
rect 4253 1273 4267 1287
rect 4133 1253 4147 1267
rect 3973 1233 3987 1247
rect 4093 1233 4107 1247
rect 3993 1214 4007 1228
rect 4053 1214 4067 1228
rect 4033 1172 4047 1186
rect 3993 1073 4007 1087
rect 4392 1353 4406 1367
rect 4413 1353 4427 1367
rect 4353 1253 4367 1267
rect 4333 1233 4347 1247
rect 4193 1214 4207 1228
rect 4293 1213 4307 1227
rect 4393 1233 4407 1247
rect 4433 1293 4447 1307
rect 4173 1172 4187 1186
rect 4133 1133 4147 1147
rect 4373 1172 4387 1186
rect 4433 1172 4447 1186
rect 4353 1153 4367 1167
rect 4233 1073 4247 1087
rect 4213 1033 4227 1047
rect 4053 914 4067 928
rect 4293 916 4307 930
rect 4333 913 4347 927
rect 3853 872 3867 886
rect 3773 853 3787 867
rect 3913 872 3927 886
rect 3873 853 3887 867
rect 3913 753 3927 767
rect 3973 753 3987 767
rect 3933 732 3947 746
rect 4193 893 4207 907
rect 4093 873 4107 887
rect 4073 853 4087 867
rect 3873 713 3887 727
rect 3693 693 3707 707
rect 3513 613 3527 627
rect 3613 652 3627 666
rect 3733 652 3747 666
rect 3853 693 3867 707
rect 3832 652 3846 666
rect 3853 653 3867 667
rect 3573 593 3587 607
rect 3793 593 3807 607
rect 3493 553 3507 567
rect 3613 394 3627 408
rect 3793 413 3807 427
rect 3893 652 3907 666
rect 3933 653 3947 667
rect 3993 693 4007 707
rect 4113 853 4127 867
rect 4233 853 4247 867
rect 4193 793 4207 807
rect 4213 773 4227 787
rect 4193 713 4207 727
rect 4113 694 4127 708
rect 4153 694 4167 708
rect 4013 652 4027 666
rect 4053 652 4067 666
rect 4113 653 4127 667
rect 4113 613 4127 627
rect 3973 433 3987 447
rect 3853 413 3867 427
rect 3813 393 3827 407
rect 3853 392 3867 406
rect 3913 413 3927 427
rect 3453 352 3467 366
rect 3633 352 3647 366
rect 3733 352 3747 366
rect 3773 352 3787 366
rect 3853 352 3867 366
rect 3893 352 3907 366
rect 3933 352 3947 366
rect 3973 352 3987 366
rect 3453 213 3467 227
rect 3513 213 3527 227
rect 3593 213 3607 227
rect 3693 213 3707 227
rect 3853 213 3867 227
rect 3433 113 3447 127
rect 3493 174 3507 188
rect 3533 174 3547 188
rect 3633 173 3647 187
rect 3553 132 3567 146
rect 3593 132 3607 146
rect 3513 113 3527 127
rect 3873 176 3887 190
rect 3933 176 3947 190
rect 3853 153 3867 167
rect 3673 113 3687 127
rect 3753 130 3767 144
rect 3713 93 3727 107
rect 3873 93 3887 107
rect 3633 73 3647 87
rect 3693 73 3707 87
rect 3733 73 3747 87
rect 3813 73 3827 87
rect 4053 394 4067 408
rect 4033 352 4047 366
rect 4073 352 4087 366
rect 4173 593 4187 607
rect 4473 1733 4487 1747
rect 4533 1734 4547 1748
rect 4493 1693 4507 1707
rect 4473 1593 4487 1607
rect 4553 1692 4567 1706
rect 4673 1873 4687 1887
rect 4653 1813 4667 1827
rect 4793 2254 4807 2268
rect 4873 2253 4887 2267
rect 4773 2212 4787 2226
rect 4813 2212 4827 2226
rect 4773 2013 4787 2027
rect 4733 1973 4747 1987
rect 4773 1954 4787 1968
rect 4873 2212 4887 2226
rect 4913 2432 4927 2446
rect 4953 2432 4967 2446
rect 4993 2413 5007 2427
rect 5033 2353 5047 2367
rect 4993 2313 5007 2327
rect 4913 2273 4927 2287
rect 4953 2254 4967 2268
rect 5013 2212 5027 2226
rect 4973 2173 4987 2187
rect 4973 2152 4987 2166
rect 4913 1993 4927 2007
rect 4713 1912 4727 1926
rect 4753 1912 4767 1926
rect 4733 1873 4747 1887
rect 4793 1873 4807 1887
rect 4693 1853 4707 1867
rect 4753 1793 4767 1807
rect 4513 1673 4527 1687
rect 4553 1434 4567 1448
rect 4593 1692 4607 1706
rect 4693 1734 4707 1748
rect 4713 1692 4727 1706
rect 4933 1954 4947 1968
rect 5013 2053 5027 2067
rect 4853 1773 4867 1787
rect 4813 1734 4827 1748
rect 4853 1734 4867 1748
rect 4913 1912 4927 1926
rect 4953 1912 4967 1926
rect 4973 1833 4987 1847
rect 4893 1773 4907 1787
rect 4953 1773 4967 1787
rect 4913 1733 4927 1747
rect 4953 1733 4967 1747
rect 5213 2953 5227 2967
rect 5173 2933 5187 2947
rect 5193 2873 5207 2887
rect 5152 2793 5166 2807
rect 5173 2793 5187 2807
rect 5113 2773 5127 2787
rect 5093 2613 5107 2627
rect 5173 2732 5187 2746
rect 5133 2673 5147 2687
rect 5113 2573 5127 2587
rect 5213 2573 5227 2587
rect 5093 2412 5107 2426
rect 5093 2373 5107 2387
rect 5073 2313 5087 2327
rect 5193 2373 5207 2387
rect 5173 2353 5187 2367
rect 5153 2273 5167 2287
rect 5133 2254 5147 2268
rect 5073 2212 5087 2226
rect 5113 2212 5127 2226
rect 5153 2212 5167 2226
rect 5213 2212 5227 2226
rect 5193 2173 5207 2187
rect 5093 2133 5107 2147
rect 5193 2093 5207 2107
rect 5053 2013 5067 2027
rect 5173 2013 5187 2027
rect 5033 1993 5047 2007
rect 5053 1953 5067 1967
rect 5073 1973 5087 1987
rect 5033 1912 5047 1926
rect 5093 1912 5107 1926
rect 5133 1853 5147 1867
rect 5073 1813 5087 1827
rect 5013 1773 5027 1787
rect 5013 1734 5027 1748
rect 4793 1692 4807 1706
rect 4893 1692 4907 1706
rect 4613 1673 4627 1687
rect 4813 1593 4827 1607
rect 4593 1553 4607 1567
rect 4793 1553 4807 1567
rect 4533 1333 4547 1347
rect 4553 1293 4567 1307
rect 4473 1213 4487 1227
rect 4513 1233 4527 1247
rect 4613 1533 4627 1547
rect 4633 1433 4647 1447
rect 4673 1333 4687 1347
rect 4633 1253 4647 1267
rect 4493 1153 4507 1167
rect 4573 1172 4587 1186
rect 4533 1113 4547 1127
rect 4453 1033 4467 1047
rect 4373 913 4387 927
rect 4413 914 4427 928
rect 4353 853 4367 867
rect 4533 853 4547 867
rect 4613 1113 4627 1127
rect 4692 1313 4706 1327
rect 4713 1313 4727 1327
rect 4933 1573 4947 1587
rect 5013 1673 5027 1687
rect 4993 1553 5007 1567
rect 4913 1513 4927 1527
rect 4993 1513 5007 1527
rect 4973 1413 4987 1427
rect 4813 1333 4827 1347
rect 4773 1293 4787 1307
rect 4773 1253 4787 1267
rect 4633 1073 4647 1087
rect 4593 953 4607 967
rect 4653 933 4667 947
rect 4593 853 4607 867
rect 4373 773 4387 787
rect 4473 773 4487 787
rect 4553 773 4567 787
rect 4333 733 4347 747
rect 4333 694 4347 708
rect 4373 696 4387 710
rect 4473 693 4487 707
rect 4293 433 4307 447
rect 4233 413 4247 427
rect 4133 394 4147 408
rect 4173 394 4187 408
rect 4353 653 4367 667
rect 4313 413 4327 427
rect 4233 373 4247 387
rect 4133 353 4147 367
rect 4493 650 4507 664
rect 4553 650 4567 664
rect 4493 613 4507 627
rect 4453 394 4467 408
rect 4533 394 4547 408
rect 4893 1352 4907 1366
rect 4993 1333 5007 1347
rect 4973 1313 4987 1327
rect 4833 1233 4847 1247
rect 4873 1233 4887 1247
rect 4933 1233 4947 1247
rect 4773 1133 4787 1147
rect 4713 953 4727 967
rect 4773 933 4787 947
rect 4773 914 4787 928
rect 4813 914 4827 928
rect 4753 872 4767 886
rect 4773 853 4787 867
rect 4713 833 4727 847
rect 4693 813 4707 827
rect 4673 753 4687 767
rect 4613 733 4627 747
rect 4713 694 4727 708
rect 4613 650 4627 664
rect 4793 833 4807 847
rect 4853 873 4867 887
rect 4832 813 4846 827
rect 4853 813 4867 827
rect 4833 694 4847 708
rect 5053 1693 5067 1707
rect 5033 1533 5047 1547
rect 5173 1813 5187 1827
rect 5093 1773 5107 1787
rect 5133 1773 5147 1787
rect 5153 1753 5167 1767
rect 5313 3233 5327 3247
rect 5273 3153 5287 3167
rect 5413 3353 5427 3367
rect 5393 3333 5407 3347
rect 5413 3294 5427 3308
rect 5493 3473 5507 3487
rect 5453 3393 5467 3407
rect 5473 3373 5487 3387
rect 5373 3213 5387 3227
rect 5333 3113 5347 3127
rect 5433 3253 5447 3267
rect 5413 3113 5427 3127
rect 5393 3073 5407 3087
rect 5373 3053 5387 3067
rect 5273 2893 5287 2907
rect 5333 2853 5347 2867
rect 5373 2853 5387 2867
rect 5273 2732 5287 2746
rect 5313 2733 5327 2747
rect 5253 2553 5267 2567
rect 5393 2813 5407 2827
rect 5333 2633 5347 2647
rect 5453 3073 5467 3087
rect 5533 3553 5547 3567
rect 5513 3433 5527 3447
rect 5593 3753 5607 3767
rect 5653 3773 5667 3787
rect 5653 3713 5667 3727
rect 5573 3693 5587 3707
rect 5633 3693 5647 3707
rect 5673 3653 5687 3667
rect 5793 4193 5807 4207
rect 5953 4333 5967 4347
rect 5973 4313 5987 4327
rect 5913 4292 5927 4306
rect 5953 4293 5967 4307
rect 5893 4253 5907 4267
rect 5853 4213 5867 4227
rect 5833 4193 5847 4207
rect 5813 4133 5827 4147
rect 5833 4093 5847 4107
rect 5753 4033 5767 4047
rect 5873 4193 5887 4207
rect 5853 4033 5867 4047
rect 5813 3992 5827 4006
rect 5853 3993 5867 4007
rect 5773 3953 5787 3967
rect 5753 3893 5767 3907
rect 5713 3813 5727 3827
rect 5813 3953 5827 3967
rect 5793 3893 5807 3907
rect 5773 3873 5787 3887
rect 5793 3833 5807 3847
rect 5733 3753 5747 3767
rect 5773 3713 5787 3727
rect 5833 3713 5847 3727
rect 5693 3633 5707 3647
rect 5653 3553 5667 3567
rect 5753 3553 5767 3567
rect 5573 3513 5587 3527
rect 5613 3514 5627 3528
rect 5693 3514 5707 3528
rect 5793 3514 5807 3528
rect 5573 3473 5587 3487
rect 5553 3453 5567 3467
rect 5593 3433 5607 3447
rect 5573 3373 5587 3387
rect 5553 3353 5567 3367
rect 5553 3313 5567 3327
rect 5493 3293 5507 3307
rect 5533 3294 5547 3308
rect 5593 3293 5607 3307
rect 5493 3253 5507 3267
rect 5573 3253 5587 3267
rect 5553 3213 5567 3227
rect 5553 3192 5567 3206
rect 5533 3173 5547 3187
rect 5553 3133 5567 3147
rect 5533 3093 5547 3107
rect 5493 3053 5507 3067
rect 5553 3053 5567 3067
rect 5472 3033 5486 3047
rect 5493 3032 5507 3046
rect 5453 3013 5467 3027
rect 5433 2994 5447 3008
rect 5493 2994 5507 3008
rect 5533 2994 5547 3008
rect 5433 2933 5447 2947
rect 5473 2893 5487 2907
rect 5553 2953 5567 2967
rect 5593 3173 5607 3187
rect 5873 3973 5887 3987
rect 5953 4253 5967 4267
rect 5973 4153 5987 4167
rect 5913 4093 5927 4107
rect 5973 4033 5987 4047
rect 5973 3973 5987 3987
rect 5893 3933 5907 3947
rect 5953 3933 5967 3947
rect 5933 3893 5947 3907
rect 5873 3753 5887 3767
rect 5853 3593 5867 3607
rect 5853 3553 5867 3567
rect 5732 3453 5746 3467
rect 5753 3453 5767 3467
rect 5653 3373 5667 3387
rect 5693 3353 5707 3367
rect 5693 3313 5707 3327
rect 5653 3293 5667 3307
rect 5732 3294 5746 3308
rect 5853 3373 5867 3387
rect 5813 3353 5827 3367
rect 5773 3313 5787 3327
rect 5753 3293 5767 3307
rect 5633 3213 5647 3227
rect 5613 3133 5627 3147
rect 5693 3233 5707 3247
rect 5633 3093 5647 3107
rect 5673 3093 5687 3107
rect 5593 2994 5607 3008
rect 5653 3073 5667 3087
rect 5633 2993 5647 3007
rect 5833 3313 5847 3327
rect 5893 3653 5907 3667
rect 5873 3294 5887 3308
rect 5913 3293 5927 3307
rect 5773 3213 5787 3227
rect 5733 3113 5747 3127
rect 5693 3033 5707 3047
rect 5673 3013 5687 3027
rect 5713 3013 5727 3027
rect 5552 2893 5566 2907
rect 5573 2893 5587 2907
rect 5513 2833 5527 2847
rect 5593 2833 5607 2847
rect 5433 2813 5447 2827
rect 5513 2793 5527 2807
rect 5473 2774 5487 2788
rect 5553 2773 5567 2787
rect 5673 2952 5687 2966
rect 5633 2853 5647 2867
rect 5693 2853 5707 2867
rect 5613 2813 5627 2827
rect 5673 2813 5687 2827
rect 5413 2713 5427 2727
rect 5413 2673 5427 2687
rect 5393 2593 5407 2607
rect 5313 2474 5327 2488
rect 5353 2474 5367 2488
rect 5293 2433 5307 2447
rect 5253 2313 5267 2327
rect 5393 2433 5407 2447
rect 5373 2413 5387 2427
rect 5333 2273 5347 2287
rect 5253 2253 5267 2267
rect 5293 2253 5307 2267
rect 5373 2293 5387 2307
rect 5353 2253 5367 2267
rect 5273 2212 5287 2226
rect 5313 2212 5327 2226
rect 5353 2213 5367 2227
rect 5353 2153 5367 2167
rect 5333 2133 5347 2147
rect 5273 2013 5287 2027
rect 5233 1973 5247 1987
rect 5253 1912 5267 1926
rect 5273 1893 5287 1907
rect 5373 2013 5387 2027
rect 5493 2713 5507 2727
rect 5493 2633 5507 2647
rect 5433 2493 5447 2507
rect 5533 2573 5547 2587
rect 5553 2533 5567 2547
rect 5553 2512 5567 2526
rect 5613 2513 5627 2527
rect 5613 2474 5627 2488
rect 5652 2474 5666 2488
rect 5733 2993 5747 3007
rect 5773 2994 5787 3008
rect 5813 3252 5827 3266
rect 5833 3173 5847 3187
rect 5833 3093 5847 3107
rect 5813 3073 5827 3087
rect 5733 2953 5747 2967
rect 5873 3073 5887 3087
rect 5913 3113 5927 3127
rect 5933 3093 5947 3107
rect 5913 3013 5927 3027
rect 5973 3513 5987 3527
rect 5973 3253 5987 3267
rect 5973 3193 5987 3207
rect 5973 3133 5987 3147
rect 5953 2993 5967 3007
rect 5893 2952 5907 2966
rect 5733 2813 5747 2827
rect 5833 2913 5847 2927
rect 5813 2893 5827 2907
rect 5713 2793 5727 2807
rect 5793 2793 5807 2807
rect 5773 2774 5787 2788
rect 5753 2713 5767 2727
rect 5693 2673 5707 2687
rect 5833 2693 5847 2707
rect 5793 2613 5807 2627
rect 5753 2533 5767 2547
rect 5673 2473 5687 2487
rect 5713 2473 5727 2487
rect 5573 2433 5587 2447
rect 5553 2413 5567 2427
rect 5593 2413 5607 2427
rect 5573 2373 5587 2387
rect 5473 2313 5487 2327
rect 5473 2292 5487 2306
rect 5433 2253 5447 2267
rect 5513 2273 5527 2287
rect 5493 2212 5507 2226
rect 5473 2193 5487 2207
rect 5453 2113 5467 2127
rect 5413 2093 5427 2107
rect 5393 1993 5407 2007
rect 5453 1993 5467 2007
rect 5353 1973 5367 1987
rect 5333 1893 5347 1907
rect 5293 1873 5307 1887
rect 5273 1773 5287 1787
rect 5213 1753 5227 1767
rect 5253 1753 5267 1767
rect 5333 1853 5347 1867
rect 5313 1793 5327 1807
rect 5193 1733 5207 1747
rect 5093 1692 5107 1706
rect 5133 1692 5147 1706
rect 5193 1693 5207 1707
rect 5173 1673 5187 1687
rect 5113 1573 5127 1587
rect 5113 1493 5127 1507
rect 5333 1773 5347 1787
rect 5253 1692 5267 1706
rect 5313 1673 5327 1687
rect 5133 1473 5147 1487
rect 5113 1453 5127 1467
rect 5073 1433 5087 1447
rect 5133 1433 5147 1447
rect 5093 1392 5107 1406
rect 5133 1393 5147 1407
rect 5053 1373 5067 1387
rect 5133 1333 5147 1347
rect 4913 1173 4927 1187
rect 4893 1033 4907 1047
rect 4733 613 4747 627
rect 4773 613 4787 627
rect 4853 652 4867 666
rect 4813 593 4827 607
rect 4613 573 4627 587
rect 4693 573 4707 587
rect 4593 513 4607 527
rect 4793 533 4807 547
rect 4753 433 4767 447
rect 4113 174 4127 188
rect 4193 352 4207 366
rect 4273 352 4287 366
rect 4313 352 4327 366
rect 4353 352 4367 366
rect 4173 174 4187 188
rect 4213 174 4227 188
rect 4533 353 4547 367
rect 4473 293 4487 307
rect 4433 253 4447 267
rect 4693 393 4707 407
rect 4593 352 4607 366
rect 4633 352 4647 366
rect 4673 353 4687 367
rect 4613 293 4627 307
rect 4553 213 4567 227
rect 4353 174 4367 188
rect 4553 153 4567 167
rect 4093 132 4107 146
rect 4133 132 4147 146
rect 4193 132 4207 146
rect 4353 133 4367 147
rect 4413 130 4427 144
rect 4473 130 4487 144
rect 4593 132 4607 146
rect 4633 132 4647 146
rect 4673 132 4687 146
rect 4953 1172 4967 1186
rect 4993 1093 5007 1107
rect 5013 1073 5027 1087
rect 4993 933 5007 947
rect 4913 913 4927 927
rect 4953 914 4967 928
rect 4912 852 4926 866
rect 4933 853 4947 867
rect 4913 652 4927 666
rect 4893 493 4907 507
rect 4873 453 4887 467
rect 4973 813 4987 827
rect 5053 1214 5067 1228
rect 5093 1214 5107 1228
rect 5053 1113 5067 1127
rect 5073 993 5087 1007
rect 5053 833 5067 847
rect 5033 793 5047 807
rect 5133 1053 5147 1067
rect 5113 933 5127 947
rect 5293 1652 5307 1666
rect 5313 1593 5327 1607
rect 5293 1573 5307 1587
rect 5313 1533 5327 1547
rect 5252 1493 5266 1507
rect 5273 1493 5287 1507
rect 5213 1434 5227 1448
rect 5233 1392 5247 1406
rect 5233 1353 5247 1367
rect 5373 1953 5387 1967
rect 5433 1954 5447 1968
rect 5453 1912 5467 1926
rect 5413 1833 5427 1847
rect 5393 1813 5407 1827
rect 5453 1813 5467 1827
rect 5373 1693 5387 1707
rect 5373 1573 5387 1587
rect 5373 1513 5387 1527
rect 5353 1493 5367 1507
rect 5333 1473 5347 1487
rect 5313 1434 5327 1448
rect 5273 1234 5287 1248
rect 5533 2033 5547 2047
rect 5493 1973 5507 1987
rect 5573 2313 5587 2327
rect 5633 2293 5647 2307
rect 5593 2273 5607 2287
rect 5573 2253 5587 2267
rect 5633 2254 5647 2268
rect 5693 2253 5707 2267
rect 5613 2212 5627 2226
rect 5693 2033 5707 2047
rect 5553 2013 5567 2027
rect 5653 2013 5667 2027
rect 5493 1913 5507 1927
rect 5413 1753 5427 1767
rect 5473 1753 5487 1767
rect 5453 1734 5467 1748
rect 5593 1912 5607 1926
rect 5593 1873 5607 1887
rect 5513 1793 5527 1807
rect 5553 1813 5567 1827
rect 5533 1773 5547 1787
rect 5513 1733 5527 1747
rect 5413 1693 5427 1707
rect 5433 1673 5447 1687
rect 5413 1593 5427 1607
rect 5333 1293 5347 1307
rect 5313 1273 5327 1287
rect 5273 1213 5287 1227
rect 5213 1172 5227 1186
rect 5193 1153 5207 1167
rect 5153 993 5167 1007
rect 5193 1013 5207 1027
rect 5173 973 5187 987
rect 5173 933 5187 947
rect 5193 913 5207 927
rect 5113 872 5127 886
rect 5153 872 5167 886
rect 5113 793 5127 807
rect 5093 753 5107 767
rect 4953 672 4967 686
rect 5133 713 5147 727
rect 5253 1013 5267 1027
rect 5293 993 5307 1007
rect 5233 973 5247 987
rect 5393 1293 5407 1307
rect 5353 1233 5367 1247
rect 5273 953 5287 967
rect 5313 953 5327 967
rect 5333 913 5347 927
rect 5213 793 5227 807
rect 5253 872 5267 886
rect 5253 833 5267 847
rect 5213 713 5227 727
rect 5213 694 5227 708
rect 5113 652 5127 666
rect 5153 652 5167 666
rect 4933 593 4947 607
rect 4973 593 4987 607
rect 4913 413 4927 427
rect 4953 413 4967 427
rect 4813 394 4827 408
rect 4853 394 4867 408
rect 4893 394 4907 408
rect 4733 352 4747 366
rect 4793 352 4807 366
rect 4873 352 4887 366
rect 4813 333 4827 347
rect 4933 353 4947 367
rect 4913 293 4927 307
rect 4893 253 4907 267
rect 4753 174 4767 188
rect 4793 174 4807 188
rect 4893 174 4907 188
rect 4733 113 4747 127
rect 4913 132 4927 146
rect 4853 113 4867 127
rect 5013 533 5027 547
rect 4993 453 5007 467
rect 5073 453 5087 467
rect 4973 253 4987 267
rect 5033 394 5047 408
rect 5093 393 5107 407
rect 5053 333 5067 347
rect 5233 573 5247 587
rect 5193 413 5207 427
rect 5133 353 5147 367
rect 5113 193 5127 207
rect 4993 174 5007 188
rect 5073 174 5087 188
rect 5173 352 5187 366
rect 5233 352 5247 366
rect 5513 1693 5527 1707
rect 5473 1593 5487 1607
rect 5473 1553 5487 1567
rect 5633 1833 5647 1847
rect 5693 2012 5707 2026
rect 5673 1973 5687 1987
rect 5633 1734 5647 1748
rect 5553 1693 5567 1707
rect 5573 1653 5587 1667
rect 5653 1693 5667 1707
rect 5653 1653 5667 1667
rect 5613 1613 5627 1627
rect 5593 1573 5607 1587
rect 5553 1533 5567 1547
rect 5593 1513 5607 1527
rect 5533 1453 5547 1467
rect 5573 1453 5587 1467
rect 5513 1433 5527 1447
rect 5513 1393 5527 1407
rect 5773 2432 5787 2446
rect 5773 2353 5787 2367
rect 5733 2293 5747 2307
rect 5813 2313 5827 2327
rect 5733 2253 5747 2267
rect 5772 2254 5786 2268
rect 5813 2254 5827 2268
rect 5753 2212 5767 2226
rect 5733 2073 5747 2087
rect 5713 1973 5727 1987
rect 5873 2873 5887 2887
rect 5913 2813 5927 2827
rect 5953 2953 5967 2967
rect 5953 2913 5967 2927
rect 5973 2853 5987 2867
rect 5933 2793 5947 2807
rect 5873 2773 5887 2787
rect 5913 2774 5927 2788
rect 5973 2773 5987 2787
rect 5893 2732 5907 2746
rect 5933 2732 5947 2746
rect 5873 2713 5887 2727
rect 5772 2193 5786 2207
rect 5793 2193 5807 2207
rect 5853 2193 5867 2207
rect 5793 2113 5807 2127
rect 5873 2073 5887 2087
rect 5793 2033 5807 2047
rect 5773 1973 5787 1987
rect 5813 1973 5827 1987
rect 5913 2673 5927 2687
rect 5953 2693 5967 2707
rect 5933 2633 5947 2647
rect 5933 2293 5947 2307
rect 5933 2253 5947 2267
rect 5913 2013 5927 2027
rect 5893 1993 5907 2007
rect 5753 1912 5767 1926
rect 5853 1954 5867 1968
rect 5933 1953 5947 1967
rect 5853 1873 5867 1887
rect 5733 1853 5747 1867
rect 5713 1793 5727 1807
rect 5753 1773 5767 1787
rect 5733 1733 5747 1747
rect 5793 1734 5807 1748
rect 5713 1713 5727 1727
rect 5753 1653 5767 1667
rect 5693 1573 5707 1587
rect 5673 1473 5687 1487
rect 5653 1453 5667 1467
rect 5693 1433 5707 1447
rect 5493 1293 5507 1307
rect 5413 1233 5427 1247
rect 5433 1213 5447 1227
rect 5373 1173 5387 1187
rect 5453 1173 5467 1187
rect 5413 1153 5427 1167
rect 5453 1133 5467 1147
rect 5453 1112 5467 1126
rect 5453 953 5467 967
rect 5393 913 5407 927
rect 5573 1392 5587 1406
rect 5633 1392 5647 1406
rect 5573 1353 5587 1367
rect 5533 1253 5547 1267
rect 5513 1233 5527 1247
rect 5493 1213 5507 1227
rect 5593 1333 5607 1347
rect 5573 1213 5587 1227
rect 5513 1172 5527 1186
rect 5553 1172 5567 1186
rect 5573 1133 5587 1147
rect 5493 1093 5507 1107
rect 5513 1053 5527 1067
rect 5493 933 5507 947
rect 5473 913 5487 927
rect 5373 833 5387 847
rect 5373 773 5387 787
rect 5313 753 5327 767
rect 5353 753 5367 767
rect 5473 873 5487 887
rect 5453 853 5467 867
rect 5533 993 5547 1007
rect 5693 1393 5707 1407
rect 5673 1293 5687 1307
rect 5613 1253 5627 1267
rect 5813 1692 5827 1706
rect 5793 1673 5807 1687
rect 5773 1533 5787 1547
rect 5753 1473 5767 1487
rect 5733 1453 5747 1467
rect 5713 1333 5727 1347
rect 5713 1293 5727 1307
rect 5693 1233 5707 1247
rect 5613 1212 5627 1226
rect 5673 1214 5687 1228
rect 5653 1172 5667 1186
rect 5673 1153 5687 1167
rect 5633 1133 5647 1147
rect 5593 973 5607 987
rect 5653 973 5667 987
rect 5573 953 5587 967
rect 5553 933 5567 947
rect 5513 873 5527 887
rect 5373 694 5387 708
rect 5313 652 5327 666
rect 5273 612 5287 626
rect 5253 293 5267 307
rect 5333 613 5347 627
rect 5313 593 5327 607
rect 5333 413 5347 427
rect 5313 352 5327 366
rect 5293 313 5307 327
rect 5273 273 5287 287
rect 5293 173 5307 187
rect 5393 413 5407 427
rect 5373 333 5387 347
rect 5473 733 5487 747
rect 5573 872 5587 886
rect 5633 852 5647 866
rect 5593 833 5607 847
rect 5573 793 5587 807
rect 5493 694 5507 708
rect 5533 693 5547 707
rect 5453 653 5467 667
rect 5513 652 5527 666
rect 5553 653 5567 667
rect 5493 613 5507 627
rect 5453 413 5467 427
rect 5413 393 5427 407
rect 5613 813 5627 827
rect 5613 773 5627 787
rect 5613 733 5627 747
rect 5593 693 5607 707
rect 5693 1073 5707 1087
rect 5713 1013 5727 1027
rect 5833 1493 5847 1507
rect 5813 1453 5827 1467
rect 5873 1793 5887 1807
rect 5893 1773 5907 1787
rect 5873 1653 5887 1667
rect 5893 1593 5907 1607
rect 5873 1533 5887 1547
rect 5853 1453 5867 1467
rect 5933 1913 5947 1927
rect 5933 1692 5947 1706
rect 5933 1613 5947 1627
rect 5913 1493 5927 1507
rect 5813 1392 5827 1406
rect 5893 1373 5907 1387
rect 5813 1253 5827 1267
rect 5773 1213 5787 1227
rect 5773 1173 5787 1187
rect 5853 1173 5867 1187
rect 5833 1133 5847 1147
rect 5813 1113 5827 1127
rect 5773 933 5787 947
rect 5873 1113 5887 1127
rect 5853 973 5867 987
rect 5673 873 5687 886
rect 5673 872 5687 873
rect 5733 872 5747 886
rect 5653 773 5667 787
rect 5813 914 5827 928
rect 5913 1253 5927 1267
rect 5913 1073 5927 1087
rect 5913 973 5927 987
rect 5893 913 5907 927
rect 5852 853 5866 867
rect 5873 853 5887 867
rect 5793 813 5807 827
rect 5833 813 5847 827
rect 5713 713 5727 727
rect 5773 713 5787 727
rect 5593 653 5607 667
rect 5573 633 5587 647
rect 5553 573 5567 587
rect 5573 453 5587 467
rect 5513 433 5527 447
rect 5433 313 5447 327
rect 5493 313 5507 327
rect 5593 433 5607 447
rect 5673 653 5687 667
rect 5693 593 5707 607
rect 5673 573 5687 587
rect 5633 493 5647 507
rect 5833 773 5847 787
rect 5773 652 5787 666
rect 5813 653 5827 667
rect 5773 613 5787 627
rect 5733 433 5747 447
rect 5613 413 5627 427
rect 5633 393 5647 407
rect 5553 273 5567 287
rect 5693 394 5707 408
rect 5793 393 5807 407
rect 5653 352 5667 366
rect 5713 352 5727 366
rect 5633 233 5647 247
rect 5393 213 5407 227
rect 5433 213 5447 227
rect 5513 213 5527 227
rect 5573 213 5587 227
rect 5373 174 5387 188
rect 4973 133 4987 147
rect 5033 132 5047 146
rect 5093 132 5107 146
rect 5133 133 5147 147
rect 5493 193 5507 207
rect 5433 153 5447 167
rect 5673 293 5687 307
rect 5893 753 5907 767
rect 5913 713 5927 727
rect 5853 653 5867 667
rect 5913 652 5927 666
rect 5873 493 5887 507
rect 5833 413 5847 427
rect 5913 413 5927 427
rect 5893 393 5907 407
rect 5813 352 5827 366
rect 5853 352 5867 366
rect 5893 353 5907 367
rect 5813 313 5827 327
rect 5713 193 5727 207
rect 5793 193 5807 207
rect 5893 293 5907 307
rect 5853 233 5867 247
rect 5973 2432 5987 2446
rect 5973 2293 5987 2307
rect 5973 1793 5987 1807
rect 5973 1733 5987 1747
rect 5973 813 5987 827
rect 5973 453 5987 467
rect 5973 393 5987 407
rect 5953 313 5967 327
rect 5193 132 5207 146
rect 5253 132 5267 146
rect 5293 132 5307 146
rect 5353 132 5367 146
rect 5393 132 5407 146
rect 5513 132 5527 146
rect 5573 132 5587 146
rect 5613 132 5627 146
rect 5653 132 5667 146
rect 5713 132 5727 146
rect 5793 132 5807 146
rect 4053 93 4067 107
rect 4153 93 4167 107
rect 4233 93 4247 107
rect 4773 93 4787 107
rect 4953 93 4967 107
rect 5913 132 5927 146
rect 3993 33 4007 47
rect 5833 33 5847 47
rect 3353 13 3367 27
rect 3393 13 3407 27
rect 3453 13 3467 27
rect 3493 13 3507 27
<< metal3 >>
rect 827 5996 913 6004
rect 2907 5996 2933 6004
rect 3547 5996 3813 6004
rect 4707 5996 4773 6004
rect 4647 5976 4673 5984
rect 4807 5976 4873 5984
rect 1727 5956 1793 5964
rect 2087 5956 2153 5964
rect 2247 5956 2433 5964
rect 2487 5956 2633 5964
rect 3767 5956 4533 5964
rect 4607 5956 5193 5964
rect 1127 5936 1313 5944
rect 1527 5936 1633 5944
rect 1647 5936 2113 5944
rect 2256 5936 2453 5944
rect 2256 5927 2264 5936
rect 3287 5936 3613 5944
rect 4027 5936 4093 5944
rect 4287 5936 4453 5944
rect 4627 5936 4833 5944
rect 5487 5936 5913 5944
rect 167 5916 213 5924
rect 2227 5916 2253 5924
rect 4487 5916 4693 5924
rect 5667 5916 5693 5924
rect 127 5896 293 5904
rect 387 5899 533 5907
rect 116 5884 124 5894
rect 1227 5896 1453 5904
rect 1547 5896 1593 5904
rect 1607 5896 1753 5904
rect 1816 5896 1933 5904
rect 116 5876 204 5884
rect 196 5866 204 5876
rect 107 5855 172 5863
rect 247 5856 373 5864
rect 1816 5866 1824 5896
rect 1947 5896 2033 5904
rect 2127 5896 2233 5904
rect 2287 5896 2313 5904
rect 2367 5897 2393 5905
rect 2507 5896 2593 5904
rect 2747 5897 2773 5905
rect 2987 5896 3033 5904
rect 3047 5897 3093 5905
rect 3147 5896 3172 5904
rect 2676 5884 2684 5894
rect 2936 5884 2944 5894
rect 3207 5897 3233 5905
rect 3347 5896 3393 5904
rect 3487 5896 3533 5904
rect 3587 5896 3633 5904
rect 3847 5897 3873 5905
rect 3953 5904 3967 5913
rect 3927 5900 3967 5904
rect 3927 5896 3964 5900
rect 3987 5896 4053 5904
rect 4167 5896 4233 5904
rect 4347 5896 4373 5904
rect 3336 5884 3344 5893
rect 2676 5876 3344 5884
rect 4416 5884 4424 5894
rect 4467 5896 4673 5904
rect 4716 5884 4724 5893
rect 4876 5884 4884 5894
rect 4947 5896 4993 5904
rect 5047 5896 5093 5904
rect 5107 5897 5153 5905
rect 5287 5897 5333 5905
rect 5387 5897 5413 5905
rect 5507 5897 5553 5905
rect 5607 5896 5633 5904
rect 5747 5896 5813 5904
rect 5827 5896 5873 5904
rect 4416 5876 4544 5884
rect 4716 5876 4884 5884
rect 747 5856 973 5864
rect 1447 5855 1513 5863
rect 1987 5855 2053 5863
rect 2107 5856 2193 5864
rect 2607 5855 2953 5863
rect 3007 5856 3073 5864
rect 3187 5855 3253 5863
rect 3427 5856 3553 5864
rect 3807 5855 3893 5863
rect 3947 5855 3973 5863
rect 4127 5855 4333 5863
rect 4447 5856 4473 5864
rect 4487 5855 4513 5863
rect 4536 5864 4544 5876
rect 4536 5856 4553 5864
rect 4747 5856 4853 5864
rect 4876 5864 4884 5876
rect 4876 5856 4913 5864
rect 5027 5856 5133 5864
rect 5187 5856 5313 5864
rect 5447 5856 5573 5864
rect 487 5836 513 5844
rect 527 5836 713 5844
rect 847 5836 913 5844
rect 2667 5836 2713 5844
rect 2807 5836 2893 5844
rect 3307 5836 3333 5844
rect 3647 5836 3833 5844
rect 4247 5836 4393 5844
rect 4707 5836 4893 5844
rect 1347 5816 1533 5824
rect 1627 5816 2273 5824
rect 2287 5816 4013 5824
rect 4567 5816 4872 5824
rect 4896 5824 4904 5833
rect 4896 5816 5273 5824
rect 5287 5816 5533 5824
rect 5727 5816 5753 5824
rect 2367 5796 2473 5804
rect 2707 5796 2733 5804
rect 2747 5796 2813 5804
rect 2827 5796 3193 5804
rect 4267 5796 4593 5804
rect 5107 5796 5153 5804
rect 1167 5776 1293 5784
rect 1307 5776 1513 5784
rect 1527 5776 1573 5784
rect 2027 5776 2153 5784
rect 2167 5776 2513 5784
rect 2727 5776 3473 5784
rect 3687 5776 4233 5784
rect 4867 5776 5493 5784
rect 667 5736 713 5744
rect 1787 5736 2173 5744
rect 2407 5736 3733 5744
rect 3847 5736 4213 5744
rect 4407 5736 4573 5744
rect 4747 5736 4773 5744
rect 4147 5716 4713 5724
rect 667 5696 1013 5704
rect 1487 5696 1653 5704
rect 1667 5696 2852 5704
rect 2887 5696 2933 5704
rect 2947 5696 3513 5704
rect 4127 5696 4773 5704
rect 4907 5696 5293 5704
rect 5307 5696 5373 5704
rect 1087 5676 1133 5684
rect 1507 5676 2333 5684
rect 3107 5676 3633 5684
rect 3747 5676 4053 5684
rect 4327 5676 4612 5684
rect 4647 5676 4713 5684
rect 1007 5656 3973 5664
rect 5587 5656 5633 5664
rect 1027 5636 1493 5644
rect 1807 5636 1912 5644
rect 1947 5636 2093 5644
rect 2107 5636 2133 5644
rect 2467 5636 2573 5644
rect 2587 5636 2633 5644
rect 2907 5636 3133 5644
rect 3247 5636 3353 5644
rect 3367 5636 3433 5644
rect 3627 5636 3693 5644
rect 4847 5636 5333 5644
rect 527 5616 553 5624
rect 847 5616 893 5624
rect 2107 5616 2153 5624
rect 2167 5616 2224 5624
rect 95 5596 132 5604
rect 76 5584 84 5594
rect 56 5580 84 5584
rect 53 5576 84 5580
rect 53 5567 67 5576
rect 95 5567 103 5596
rect 167 5596 193 5604
rect 127 5555 153 5563
rect 167 5555 193 5563
rect 256 5564 264 5594
rect 256 5556 293 5564
rect 436 5564 444 5596
rect 627 5596 733 5604
rect 747 5597 793 5605
rect 807 5596 953 5604
rect 967 5596 1113 5604
rect 1347 5596 1413 5604
rect 1547 5597 1573 5605
rect 1627 5597 1673 5605
rect 1887 5597 1973 5605
rect 1987 5596 2053 5604
rect 2076 5596 2133 5604
rect 1296 5584 1304 5594
rect 1247 5576 1304 5584
rect 1456 5584 1464 5594
rect 1387 5576 1464 5584
rect 436 5556 633 5564
rect 727 5555 813 5563
rect 1327 5556 1433 5564
rect 1487 5556 1513 5564
rect 1647 5556 1693 5564
rect 2076 5566 2084 5596
rect 2216 5604 2224 5616
rect 2247 5616 2333 5624
rect 2667 5616 2753 5624
rect 4247 5616 4273 5624
rect 4287 5616 4453 5624
rect 4587 5616 4613 5624
rect 5800 5624 5813 5627
rect 5796 5614 5813 5624
rect 5796 5613 5820 5614
rect 2216 5596 2273 5604
rect 2513 5584 2527 5593
rect 2513 5580 2584 5584
rect 2516 5576 2584 5580
rect 1827 5556 1913 5564
rect 1967 5555 2013 5563
rect 2187 5556 2253 5564
rect 2307 5556 2353 5564
rect 2367 5556 2393 5564
rect 2487 5555 2553 5563
rect 2576 5564 2584 5576
rect 2576 5556 2593 5564
rect 2716 5564 2724 5594
rect 2987 5597 3053 5605
rect 3127 5597 3193 5605
rect 3307 5597 3393 5605
rect 3587 5597 3613 5605
rect 3987 5597 4193 5605
rect 4547 5596 4653 5604
rect 4667 5596 4833 5604
rect 5047 5597 5073 5605
rect 5156 5596 5253 5604
rect 2687 5556 2724 5564
rect 2856 5564 2864 5593
rect 2856 5556 2873 5564
rect 2927 5555 2953 5563
rect 3147 5556 3213 5564
rect 3447 5556 3513 5564
rect 3536 5564 3544 5594
rect 3736 5567 3744 5594
rect 4376 5576 4433 5584
rect 3536 5556 3593 5564
rect 3647 5556 3673 5564
rect 3736 5556 3752 5567
rect 3740 5553 3752 5556
rect 3787 5556 4153 5564
rect 4376 5566 4384 5576
rect 4996 5584 5004 5594
rect 4996 5576 5024 5584
rect 4467 5556 4513 5564
rect 4587 5556 4624 5564
rect 267 5536 313 5544
rect 687 5536 973 5544
rect 1547 5536 1593 5544
rect 2667 5536 2713 5544
rect 3007 5544 3020 5547
rect 3007 5536 3073 5544
rect 3007 5533 3024 5536
rect 3387 5536 3413 5544
rect 107 5516 133 5524
rect 1007 5516 1233 5524
rect 1247 5516 1373 5524
rect 1447 5516 1773 5524
rect 2647 5516 2733 5524
rect 3016 5524 3024 5533
rect 3787 5536 3873 5544
rect 4047 5536 4113 5544
rect 4616 5544 4624 5556
rect 4687 5556 4713 5564
rect 4907 5556 4933 5564
rect 5016 5564 5024 5576
rect 5016 5556 5093 5564
rect 5116 5547 5124 5594
rect 5156 5584 5164 5596
rect 5447 5597 5473 5605
rect 5396 5584 5404 5594
rect 5136 5576 5164 5584
rect 5316 5576 5404 5584
rect 5136 5566 5144 5576
rect 5187 5555 5233 5563
rect 5316 5564 5324 5576
rect 5287 5556 5324 5564
rect 5347 5556 5593 5564
rect 5616 5564 5624 5594
rect 5796 5566 5804 5613
rect 5827 5596 5893 5604
rect 5907 5596 5953 5604
rect 5616 5556 5753 5564
rect 4616 5536 4713 5544
rect 2947 5516 3024 5524
rect 3107 5516 3253 5524
rect 3267 5516 3333 5524
rect 3567 5516 3713 5524
rect 3727 5516 4193 5524
rect 4607 5516 4733 5524
rect 4747 5516 4773 5524
rect 5007 5516 5033 5524
rect 67 5496 93 5504
rect 287 5496 593 5504
rect 907 5496 1133 5504
rect 2127 5496 2973 5504
rect 3587 5496 3773 5504
rect 3827 5496 4073 5504
rect 4187 5496 4633 5504
rect 5707 5496 5973 5504
rect 867 5476 1273 5484
rect 1927 5476 1973 5484
rect 1987 5476 2653 5484
rect 2976 5484 2984 5493
rect 2976 5476 3293 5484
rect 3447 5476 3593 5484
rect 3607 5476 3753 5484
rect 3767 5476 4653 5484
rect 5427 5476 5793 5484
rect 247 5456 373 5464
rect 927 5456 973 5464
rect 2447 5456 2493 5464
rect 2607 5456 2673 5464
rect 2767 5456 2793 5464
rect 2887 5456 3573 5464
rect 3647 5456 3873 5464
rect 4127 5456 4593 5464
rect 4707 5456 4753 5464
rect 5007 5456 5313 5464
rect 2307 5436 2513 5444
rect 3707 5436 4033 5444
rect 4627 5436 4673 5444
rect 4727 5436 4793 5444
rect 4807 5436 5453 5444
rect 587 5416 733 5424
rect 747 5416 853 5424
rect 1567 5416 2773 5424
rect 3207 5416 3513 5424
rect 3607 5416 4353 5424
rect 4707 5416 4973 5424
rect 4987 5416 5113 5424
rect 5687 5416 5933 5424
rect 1067 5396 1233 5404
rect 2047 5396 2193 5404
rect 3047 5396 3133 5404
rect 3596 5404 3604 5413
rect 3147 5396 3604 5404
rect 4167 5396 4213 5404
rect 5427 5396 5473 5404
rect 47 5377 213 5385
rect 227 5376 253 5384
rect 427 5377 573 5385
rect 647 5376 693 5384
rect 707 5377 733 5385
rect 907 5377 953 5385
rect 856 5364 864 5374
rect 1127 5376 1173 5384
rect 856 5356 1084 5364
rect 247 5335 273 5343
rect 767 5336 873 5344
rect 1007 5336 1033 5344
rect 1076 5344 1084 5356
rect 1076 5336 1193 5344
rect 1316 5344 1324 5374
rect 1407 5376 1433 5384
rect 1627 5376 1693 5384
rect 1707 5377 1793 5385
rect 1936 5376 2033 5384
rect 1476 5344 1484 5374
rect 1936 5346 1944 5376
rect 2087 5376 2153 5384
rect 2247 5377 2293 5385
rect 2387 5376 2573 5384
rect 2587 5377 2693 5385
rect 2787 5384 2800 5387
rect 2787 5373 2804 5384
rect 2907 5377 2973 5385
rect 1316 5336 1753 5344
rect 1987 5335 2013 5343
rect 2307 5336 2353 5344
rect 2796 5346 2804 5373
rect 2607 5336 2673 5344
rect 3007 5335 3033 5343
rect 3167 5335 3193 5343
rect 3276 5344 3284 5374
rect 3527 5376 3693 5384
rect 3927 5376 3993 5384
rect 4007 5377 4093 5385
rect 4247 5377 4293 5385
rect 4407 5376 4453 5384
rect 4356 5364 4364 5374
rect 4467 5376 4513 5384
rect 4567 5376 4593 5384
rect 4907 5376 5213 5384
rect 5287 5377 5353 5385
rect 5376 5376 5513 5384
rect 5216 5364 5224 5374
rect 5376 5364 5384 5376
rect 5687 5376 5833 5384
rect 5847 5377 5893 5385
rect 4356 5356 4704 5364
rect 5216 5356 5384 5364
rect 3276 5336 3453 5344
rect 3587 5336 3713 5344
rect 3907 5336 4013 5344
rect 4067 5336 4213 5344
rect 4307 5336 4373 5344
rect 4607 5335 4673 5343
rect 4696 5344 4704 5356
rect 4696 5336 4713 5344
rect 4987 5335 5073 5343
rect 5347 5336 5493 5344
rect 5707 5336 5813 5344
rect 87 5316 173 5324
rect 187 5316 313 5324
rect 327 5316 393 5324
rect 467 5316 553 5324
rect 4427 5316 4533 5324
rect 5287 5316 5393 5324
rect 5667 5316 5853 5324
rect 867 5296 913 5304
rect 987 5296 1133 5304
rect 1307 5296 1653 5304
rect 1767 5296 2093 5304
rect 2227 5296 2493 5304
rect 2967 5296 3193 5304
rect 3707 5296 4113 5304
rect 4267 5296 4453 5304
rect 4467 5296 4633 5304
rect 4847 5296 5013 5304
rect 527 5276 953 5284
rect 2327 5276 2593 5284
rect 2767 5276 2813 5284
rect 4047 5276 4132 5284
rect 4167 5276 4253 5284
rect 4787 5276 5053 5284
rect 5207 5276 5573 5284
rect 1167 5256 1233 5264
rect 1247 5256 1313 5264
rect 1727 5256 1833 5264
rect 2907 5256 3113 5264
rect 3127 5256 3253 5264
rect 3267 5256 3673 5264
rect 3727 5256 3813 5264
rect 3867 5256 4333 5264
rect 4347 5256 4413 5264
rect 2187 5236 2413 5244
rect 3327 5236 3413 5244
rect 3427 5236 3733 5244
rect 3787 5236 4833 5244
rect 4887 5236 5193 5244
rect 5387 5236 5413 5244
rect 5427 5236 5833 5244
rect 2287 5216 2773 5224
rect 2907 5216 3113 5224
rect 3527 5216 3713 5224
rect 4027 5216 4453 5224
rect 5867 5216 5893 5224
rect 127 5196 293 5204
rect 307 5196 353 5204
rect 367 5196 793 5204
rect 2267 5196 2693 5204
rect 2707 5196 2733 5204
rect 2847 5196 3813 5204
rect 4107 5196 4344 5204
rect 2507 5176 2553 5184
rect 2687 5176 3073 5184
rect 3167 5176 3673 5184
rect 4247 5176 4313 5184
rect 4336 5184 4344 5196
rect 4336 5176 4793 5184
rect 2067 5156 2113 5164
rect 3127 5156 3693 5164
rect 3947 5156 4753 5164
rect 5107 5156 5373 5164
rect 5387 5156 5653 5164
rect 1127 5136 1233 5144
rect 2407 5136 2493 5144
rect 2587 5136 2833 5144
rect 3727 5136 3853 5144
rect 4067 5136 4513 5144
rect 4787 5136 4993 5144
rect 27 5116 233 5124
rect 567 5116 733 5124
rect 1027 5116 1093 5124
rect 1307 5116 1433 5124
rect 1607 5116 1793 5124
rect 1807 5116 3133 5124
rect 3707 5116 3753 5124
rect 4567 5116 4713 5124
rect 547 5096 573 5104
rect 2147 5096 2453 5104
rect 3227 5096 3784 5104
rect 3776 5088 3784 5096
rect 3987 5096 4073 5104
rect 4767 5096 4873 5104
rect 67 5076 93 5084
rect 116 5076 193 5084
rect 116 5046 124 5076
rect 307 5077 393 5085
rect 407 5076 493 5084
rect 236 5064 244 5074
rect 607 5076 653 5084
rect 676 5076 793 5084
rect 236 5056 433 5064
rect 676 5064 684 5076
rect 947 5076 993 5084
rect 1087 5077 1113 5085
rect 636 5056 684 5064
rect 227 5036 293 5044
rect 636 5046 644 5056
rect 727 5036 773 5044
rect 887 5036 913 5044
rect 967 5036 1113 5044
rect 1127 5036 1173 5044
rect 1196 5007 1204 5074
rect 1347 5076 1393 5084
rect 1567 5077 1633 5085
rect 1716 5076 1733 5084
rect 1716 5064 1724 5076
rect 1827 5077 1893 5085
rect 1987 5077 2053 5085
rect 1667 5056 1724 5064
rect 1776 5047 1784 5074
rect 2307 5076 2333 5084
rect 2847 5077 2913 5085
rect 3267 5077 3313 5085
rect 1327 5036 1373 5044
rect 1587 5036 1713 5044
rect 1776 5036 1793 5047
rect 1780 5033 1793 5036
rect 1847 5036 1873 5044
rect 1927 5036 2033 5044
rect 2096 5044 2104 5073
rect 2087 5036 2104 5044
rect 2367 5035 2393 5043
rect 2436 5044 2444 5073
rect 2956 5064 2964 5074
rect 3507 5076 3553 5084
rect 3627 5077 3653 5085
rect 3787 5077 3873 5085
rect 4167 5077 4213 5085
rect 4320 5084 4333 5087
rect 2956 5056 3024 5064
rect 2436 5036 2473 5044
rect 2667 5036 2693 5044
rect 3016 5046 3024 5056
rect 2707 5036 2753 5044
rect 2767 5036 2893 5044
rect 3027 5035 3093 5043
rect 3247 5036 3273 5044
rect 3447 5036 3473 5044
rect 3487 5036 3533 5044
rect 3736 5044 3744 5073
rect 3727 5036 3744 5044
rect 3767 5036 3853 5044
rect 4116 5044 4124 5074
rect 4316 5073 4333 5084
rect 4387 5076 4413 5084
rect 4436 5076 4553 5084
rect 4007 5036 4273 5044
rect 4316 5046 4324 5073
rect 4436 5064 4444 5076
rect 4667 5077 4713 5085
rect 4887 5077 4953 5085
rect 5127 5077 5153 5085
rect 4396 5060 4444 5064
rect 4393 5056 4444 5060
rect 4393 5047 4407 5056
rect 4647 5035 4693 5043
rect 4836 5044 4844 5074
rect 5036 5064 5044 5074
rect 5196 5064 5204 5074
rect 5247 5076 5273 5084
rect 5347 5076 5433 5084
rect 5487 5077 5513 5085
rect 5567 5076 5673 5084
rect 4947 5056 5204 5064
rect 4747 5036 4844 5044
rect 5027 5036 5093 5044
rect 5196 5044 5204 5056
rect 5736 5064 5744 5074
rect 5707 5056 5744 5064
rect 5196 5036 5313 5044
rect 5427 5035 5453 5043
rect 5507 5036 5553 5044
rect 5807 5036 5953 5044
rect 3296 5016 3844 5024
rect 3296 5007 3304 5016
rect 107 4996 573 5004
rect 827 4996 1053 5004
rect 1187 4996 1204 5007
rect 1187 4993 1200 4996
rect 1767 4996 1973 5004
rect 1987 4996 2493 5004
rect 3207 4996 3293 5004
rect 3407 4996 3493 5004
rect 3587 4996 3613 5004
rect 3627 4996 3753 5004
rect 3836 5004 3844 5016
rect 4336 5016 4593 5024
rect 3836 4996 3893 5004
rect 4007 4996 4073 5004
rect 4336 5004 4344 5016
rect 4767 5016 4853 5024
rect 4927 5016 5113 5024
rect 5127 5016 5233 5024
rect 5727 5016 5753 5024
rect 4187 4996 4344 5004
rect 4387 4996 4533 5004
rect 4756 5004 4764 5013
rect 4667 4996 4764 5004
rect 5067 4996 5413 5004
rect 5467 4996 5573 5004
rect 867 4976 953 4984
rect 1427 4976 1493 4984
rect 1507 4976 1533 4984
rect 1647 4976 1733 4984
rect 1807 4976 1913 4984
rect 2127 4976 2353 4984
rect 2787 4976 2973 4984
rect 2987 4976 3053 4984
rect 3787 4976 3812 4984
rect 3847 4976 4053 4984
rect 4587 4976 4933 4984
rect 5147 4976 5193 4984
rect 1267 4956 1393 4964
rect 3187 4956 3673 4964
rect 3867 4956 4033 4964
rect 4287 4956 4433 4964
rect 4607 4956 4913 4964
rect 5387 4956 5533 4964
rect 547 4936 633 4944
rect 987 4936 1013 4944
rect 1847 4936 2853 4944
rect 2947 4936 3153 4944
rect 3207 4936 3473 4944
rect 3707 4936 3933 4944
rect 4167 4936 4253 4944
rect 4747 4936 4773 4944
rect 5167 4936 5553 4944
rect 5667 4936 5773 4944
rect 667 4916 673 4924
rect 687 4916 993 4924
rect 1487 4916 1573 4924
rect 3567 4916 4033 4924
rect 4087 4916 4213 4924
rect 4467 4916 4613 4924
rect 5187 4916 5504 4924
rect 5496 4907 5504 4916
rect 527 4896 573 4904
rect 787 4896 993 4904
rect 1807 4896 2193 4904
rect 2207 4896 2233 4904
rect 2247 4896 2513 4904
rect 2607 4896 3073 4904
rect 3167 4896 3304 4904
rect 227 4876 433 4884
rect 447 4876 493 4884
rect 3296 4884 3304 4896
rect 3687 4896 3733 4904
rect 3927 4896 3973 4904
rect 5227 4896 5293 4904
rect 5307 4896 5413 4904
rect 5507 4896 5733 4904
rect 3296 4876 3313 4884
rect 3327 4876 3613 4884
rect 4327 4876 4353 4884
rect 4487 4876 4713 4884
rect 5687 4876 5973 4884
rect 67 4864 80 4867
rect 67 4853 84 4864
rect 387 4856 413 4864
rect 707 4859 913 4867
rect 987 4856 1044 4864
rect 76 4826 84 4853
rect 127 4816 233 4824
rect 1036 4826 1044 4856
rect 787 4816 813 4824
rect 1056 4807 1064 4854
rect 1216 4824 1224 4873
rect 1347 4857 1433 4865
rect 1627 4856 1693 4864
rect 1707 4856 1873 4864
rect 1927 4856 2073 4864
rect 2087 4856 2313 4864
rect 2407 4857 2453 4865
rect 2587 4857 2613 4865
rect 2667 4856 2773 4864
rect 2827 4856 2853 4864
rect 2867 4857 2953 4865
rect 3127 4857 3193 4865
rect 3247 4857 3273 4865
rect 3427 4856 3513 4864
rect 3956 4856 3973 4864
rect 3956 4844 3964 4856
rect 3987 4856 4233 4864
rect 4247 4857 4433 4865
rect 4567 4856 4613 4864
rect 4627 4857 4673 4865
rect 4867 4856 4884 4864
rect 3676 4836 3964 4844
rect 1607 4816 1713 4824
rect 1767 4816 1813 4824
rect 1947 4816 2053 4824
rect 2107 4816 2193 4824
rect 2207 4816 2293 4824
rect 2347 4816 2473 4824
rect 3147 4815 3213 4823
rect 3676 4824 3684 4836
rect 3647 4816 3713 4824
rect 3787 4815 3853 4823
rect 3867 4815 4013 4823
rect 4107 4816 4213 4824
rect 4227 4816 4353 4824
rect 4707 4816 4833 4824
rect 4876 4824 4884 4856
rect 4907 4856 4953 4864
rect 4967 4856 4993 4864
rect 5007 4856 5113 4864
rect 5136 4856 5253 4864
rect 5136 4844 5144 4856
rect 5527 4857 5593 4865
rect 5647 4856 5833 4864
rect 5087 4836 5144 4844
rect 4876 4816 4913 4824
rect 5447 4816 5493 4824
rect 5796 4826 5804 4856
rect 487 4796 633 4804
rect 1907 4796 2093 4804
rect 2847 4796 2893 4804
rect 3767 4796 3813 4804
rect 4056 4804 4064 4812
rect 3827 4796 4064 4804
rect 4587 4796 4693 4804
rect 5027 4796 5193 4804
rect 5367 4796 5613 4804
rect 767 4776 813 4784
rect 827 4776 873 4784
rect 887 4776 1273 4784
rect 1327 4776 1413 4784
rect 1587 4776 1653 4784
rect 2247 4776 2513 4784
rect 2587 4776 2633 4784
rect 3187 4776 3293 4784
rect 4267 4776 4453 4784
rect 4547 4776 4653 4784
rect 4667 4776 5133 4784
rect 5387 4776 5753 4784
rect 1047 4756 1173 4764
rect 2567 4756 2793 4764
rect 3107 4756 3153 4764
rect 3467 4756 3733 4764
rect 3747 4756 3773 4764
rect 3827 4756 4053 4764
rect 4827 4756 5273 4764
rect 2487 4736 2613 4744
rect 2827 4736 2913 4744
rect 3487 4736 3553 4744
rect 5276 4744 5284 4753
rect 5276 4736 5393 4744
rect 887 4716 913 4724
rect 1947 4716 2253 4724
rect 3027 4716 3153 4724
rect 3607 4716 3933 4724
rect 3947 4716 3993 4724
rect 4087 4716 4153 4724
rect 4227 4716 4373 4724
rect 5567 4716 5913 4724
rect 3596 4704 3604 4713
rect 3287 4696 3604 4704
rect 3647 4696 3673 4704
rect 3687 4696 3893 4704
rect 4027 4696 4093 4704
rect 4167 4696 4392 4704
rect 4427 4696 4764 4704
rect 2387 4676 2764 4684
rect 2756 4667 2764 4676
rect 3387 4676 3592 4684
rect 3627 4676 3693 4684
rect 3927 4676 4573 4684
rect 4587 4676 4613 4684
rect 4756 4684 4764 4696
rect 4756 4676 4833 4684
rect 4927 4676 5293 4684
rect 5307 4676 5513 4684
rect 147 4656 293 4664
rect 307 4656 353 4664
rect 2207 4656 2653 4664
rect 2767 4656 2853 4664
rect 2867 4656 3813 4664
rect 4747 4656 4873 4664
rect 5087 4656 5173 4664
rect 1667 4636 2153 4644
rect 2507 4636 2593 4644
rect 2607 4636 2713 4644
rect 3007 4636 3053 4644
rect 3167 4636 4273 4644
rect 4627 4636 4772 4644
rect 4807 4636 4913 4644
rect 107 4616 313 4624
rect 447 4616 513 4624
rect 1567 4616 1833 4624
rect 2087 4616 2173 4624
rect 2187 4616 2213 4624
rect 2427 4616 2813 4624
rect 3447 4616 3633 4624
rect 3847 4616 3893 4624
rect 4067 4616 4213 4624
rect 4847 4616 4973 4624
rect 5187 4616 5573 4624
rect 607 4596 693 4604
rect 1367 4596 1533 4604
rect 1547 4596 2144 4604
rect 367 4576 413 4584
rect 2136 4584 2144 4596
rect 2527 4596 2553 4604
rect 2567 4596 2773 4604
rect 3276 4596 3973 4604
rect 3276 4587 3284 4596
rect 4327 4596 4353 4604
rect 4447 4596 4993 4604
rect 2136 4576 2193 4584
rect 2467 4576 2493 4584
rect 3067 4576 3213 4584
rect 3227 4576 3273 4584
rect 5267 4576 5353 4584
rect 5627 4576 5733 4584
rect 207 4557 253 4565
rect 167 4516 193 4524
rect 296 4507 304 4573
rect 507 4556 593 4564
rect 667 4556 733 4564
rect 747 4556 764 4564
rect 396 4527 404 4553
rect 756 4544 764 4556
rect 787 4556 833 4564
rect 847 4557 873 4565
rect 927 4557 1053 4565
rect 1067 4557 1113 4565
rect 1187 4556 1253 4564
rect 1267 4556 1433 4564
rect 1627 4557 1713 4565
rect 756 4540 804 4544
rect 756 4536 807 4540
rect 793 4527 807 4536
rect 467 4516 533 4524
rect 907 4516 993 4524
rect 1127 4516 1413 4524
rect 1476 4507 1484 4554
rect 1847 4557 1893 4565
rect 1987 4557 2013 4565
rect 2287 4556 2333 4564
rect 1507 4516 1573 4524
rect 1756 4524 1764 4553
rect 2116 4544 2124 4554
rect 2347 4556 2373 4564
rect 2116 4536 2313 4544
rect 2696 4544 2704 4554
rect 2636 4536 2704 4544
rect 1647 4516 1764 4524
rect 1827 4515 1873 4523
rect 2047 4516 2093 4524
rect 2247 4516 2393 4524
rect 2407 4515 2513 4523
rect 2636 4524 2644 4536
rect 2587 4516 2644 4524
rect 2667 4516 2713 4524
rect 2736 4524 2744 4554
rect 2787 4556 2884 4564
rect 2736 4516 2773 4524
rect 2876 4524 2884 4556
rect 2947 4557 2973 4565
rect 3267 4556 3333 4564
rect 2876 4516 2913 4524
rect 3007 4516 3073 4524
rect 647 4496 833 4504
rect 1267 4496 1333 4504
rect 1747 4496 1773 4504
rect 1947 4496 2013 4504
rect 2807 4496 2853 4504
rect 2947 4496 3033 4504
rect 3096 4504 3104 4554
rect 3347 4556 3373 4564
rect 3400 4564 3413 4567
rect 3396 4553 3413 4564
rect 3647 4557 3673 4565
rect 3767 4557 3833 4565
rect 4047 4556 4153 4564
rect 3247 4516 3293 4524
rect 3396 4507 3404 4553
rect 3496 4524 3504 4553
rect 3427 4516 3504 4524
rect 3536 4507 3544 4554
rect 3567 4515 3613 4523
rect 3876 4524 3884 4554
rect 4287 4564 4300 4567
rect 4287 4553 4304 4564
rect 4467 4557 4493 4565
rect 4296 4544 4304 4553
rect 4236 4540 4304 4544
rect 4233 4536 4304 4540
rect 4233 4527 4247 4536
rect 3707 4516 3884 4524
rect 4027 4516 4113 4524
rect 4296 4526 4304 4536
rect 4356 4527 4364 4553
rect 4447 4515 4473 4523
rect 4527 4515 4573 4523
rect 4656 4524 4664 4554
rect 4627 4516 4664 4524
rect 4696 4527 4704 4554
rect 4696 4516 4713 4527
rect 4700 4513 4713 4516
rect 4816 4526 4824 4573
rect 4847 4556 4893 4564
rect 4907 4557 4953 4565
rect 5007 4556 5133 4564
rect 5487 4557 5513 4565
rect 4867 4516 4933 4524
rect 4987 4516 5053 4524
rect 5176 4524 5184 4554
rect 5176 4516 5273 4524
rect 5436 4524 5444 4554
rect 5787 4557 5833 4565
rect 5947 4556 6024 4564
rect 5676 4527 5684 4553
rect 5873 4544 5887 4553
rect 5873 4540 5904 4544
rect 5876 4536 5904 4540
rect 5436 4516 5593 4524
rect 5896 4524 5904 4536
rect 5896 4516 5953 4524
rect 3096 4496 3132 4504
rect 3167 4496 3193 4504
rect 3487 4496 3512 4504
rect 3647 4496 3673 4504
rect 3727 4496 3753 4504
rect 3887 4496 3913 4504
rect 4047 4496 4173 4504
rect 4187 4496 4253 4504
rect 5167 4496 5313 4504
rect 5327 4496 5353 4504
rect 5427 4496 5493 4504
rect 5507 4496 5553 4504
rect 5747 4496 5833 4504
rect 5887 4496 5933 4504
rect 387 4476 433 4484
rect 447 4476 753 4484
rect 2407 4476 2633 4484
rect 2647 4476 2732 4484
rect 2767 4476 3113 4484
rect 3267 4476 3333 4484
rect 3427 4476 3553 4484
rect 3867 4476 3893 4484
rect 4347 4476 4613 4484
rect 5527 4476 5613 4484
rect 47 4456 193 4464
rect 347 4456 473 4464
rect 1207 4456 1673 4464
rect 1687 4456 1953 4464
rect 1976 4456 2093 4464
rect 1467 4436 1533 4444
rect 1976 4444 1984 4456
rect 2387 4456 2433 4464
rect 2587 4456 2833 4464
rect 3067 4456 3233 4464
rect 3547 4456 3693 4464
rect 4287 4456 4413 4464
rect 4676 4447 4684 4473
rect 4707 4456 4753 4464
rect 4887 4456 5073 4464
rect 5127 4456 5213 4464
rect 5647 4456 5693 4464
rect 5707 4456 5753 4464
rect 1727 4436 1984 4444
rect 2047 4436 2153 4444
rect 2167 4436 2193 4444
rect 2547 4436 2813 4444
rect 2827 4436 3413 4444
rect 3427 4436 3933 4444
rect 4676 4446 4700 4447
rect 4676 4436 4693 4446
rect 4680 4433 4693 4436
rect 47 4416 373 4424
rect 1087 4416 1273 4424
rect 1716 4424 1724 4433
rect 5167 4436 5273 4444
rect 5387 4436 5533 4444
rect 5627 4436 5793 4444
rect 5807 4436 5853 4444
rect 1387 4416 1724 4424
rect 2187 4416 2524 4424
rect 727 4396 773 4404
rect 1447 4396 1833 4404
rect 1887 4396 2053 4404
rect 2107 4396 2273 4404
rect 2516 4404 2524 4416
rect 3047 4416 3093 4424
rect 3147 4416 3473 4424
rect 3656 4416 3813 4424
rect 2516 4396 2573 4404
rect 2687 4396 3493 4404
rect 3656 4404 3664 4416
rect 4167 4416 4552 4424
rect 4587 4416 5553 4424
rect 5727 4416 5893 4424
rect 3507 4396 3664 4404
rect 3707 4396 3773 4404
rect 4367 4396 4513 4404
rect 4627 4396 4733 4404
rect 5087 4396 5413 4404
rect 5527 4396 5744 4404
rect 127 4376 173 4384
rect 227 4376 353 4384
rect 407 4380 524 4384
rect 407 4376 527 4380
rect 356 4364 364 4373
rect 513 4366 527 4376
rect 987 4376 1213 4384
rect 1487 4376 2073 4384
rect 2147 4376 2593 4384
rect 2987 4376 3373 4384
rect 3847 4376 4033 4384
rect 4787 4376 4913 4384
rect 4927 4376 5033 4384
rect 5107 4376 5213 4384
rect 5567 4376 5713 4384
rect 5736 4384 5744 4396
rect 5736 4376 5973 4384
rect 356 4356 504 4364
rect 147 4336 153 4344
rect 167 4336 333 4344
rect 496 4344 504 4356
rect 707 4356 753 4364
rect 867 4356 893 4364
rect 1607 4356 1673 4364
rect 1687 4356 1793 4364
rect 1927 4356 1993 4364
rect 2467 4356 2813 4364
rect 2907 4356 3052 4364
rect 3087 4356 3313 4364
rect 3327 4356 3653 4364
rect 3667 4356 3733 4364
rect 3827 4356 4113 4364
rect 4207 4356 4253 4364
rect 4467 4356 4593 4364
rect 4827 4356 4853 4364
rect 4867 4356 4973 4364
rect 5467 4356 5533 4364
rect 496 4336 553 4344
rect 336 4324 344 4334
rect 627 4337 673 4345
rect 827 4336 1064 4344
rect 276 4316 344 4324
rect 276 4304 284 4316
rect 247 4296 284 4304
rect 307 4295 353 4303
rect 447 4295 693 4303
rect 1056 4304 1064 4336
rect 1127 4337 1173 4345
rect 987 4296 1013 4304
rect 1056 4296 1073 4304
rect 1396 4304 1404 4333
rect 1447 4336 1493 4344
rect 1547 4336 1633 4344
rect 1967 4344 1980 4347
rect 1967 4333 1984 4344
rect 2167 4337 2393 4345
rect 2647 4337 2673 4345
rect 1976 4306 1984 4333
rect 1367 4296 1513 4304
rect 1707 4296 1813 4304
rect 1827 4295 1913 4303
rect 2116 4304 2124 4334
rect 2847 4344 2860 4347
rect 2847 4333 2864 4344
rect 3107 4336 3133 4344
rect 3247 4336 3333 4344
rect 2856 4324 2864 4333
rect 3336 4324 3344 4334
rect 3547 4337 3613 4345
rect 3927 4336 3944 4344
rect 2856 4316 3024 4324
rect 2067 4296 2124 4304
rect 2336 4296 2353 4304
rect 407 4276 473 4284
rect 2336 4284 2344 4296
rect 2856 4306 2864 4316
rect 3016 4306 3024 4316
rect 3196 4316 3344 4324
rect 2367 4296 2413 4304
rect 2427 4296 2573 4304
rect 2627 4295 2693 4303
rect 2767 4295 2813 4303
rect 3067 4295 3093 4303
rect 3196 4304 3204 4316
rect 3187 4296 3204 4304
rect 3376 4304 3384 4333
rect 3367 4296 3384 4304
rect 3427 4296 3453 4304
rect 3507 4296 3553 4304
rect 3567 4296 3593 4304
rect 3687 4296 3753 4304
rect 3827 4295 3853 4303
rect 3936 4304 3944 4336
rect 4220 4344 4233 4347
rect 4216 4333 4233 4344
rect 4667 4337 4693 4345
rect 5287 4336 5353 4344
rect 4036 4307 4044 4333
rect 4076 4307 4084 4333
rect 4216 4324 4224 4333
rect 4127 4316 4224 4324
rect 3936 4296 3993 4304
rect 4176 4306 4184 4316
rect 4616 4324 4624 4333
rect 4267 4316 4624 4324
rect 4307 4296 4353 4304
rect 4367 4296 4593 4304
rect 4687 4296 4713 4304
rect 4727 4296 4753 4304
rect 4807 4296 4893 4304
rect 4996 4287 5004 4333
rect 5027 4296 5073 4304
rect 5116 4304 5124 4334
rect 5847 4337 5893 4345
rect 5087 4296 5124 4304
rect 5227 4296 5253 4304
rect 5467 4296 5513 4304
rect 5576 4287 5584 4334
rect 5776 4304 5784 4334
rect 5956 4307 5964 4333
rect 5987 4316 6024 4324
rect 5776 4296 5913 4304
rect 6016 4296 6024 4316
rect 2307 4276 2344 4284
rect 2967 4276 3213 4284
rect 3627 4276 3653 4284
rect 4427 4276 4493 4284
rect 127 4256 653 4264
rect 1087 4256 1233 4264
rect 1307 4256 1593 4264
rect 2487 4256 2513 4264
rect 2527 4256 2713 4264
rect 3127 4256 3193 4264
rect 3407 4256 3464 4264
rect 227 4236 453 4244
rect 847 4236 1173 4244
rect 2027 4236 2073 4244
rect 2087 4236 2133 4244
rect 2747 4236 2773 4244
rect 2787 4236 3093 4244
rect 3456 4244 3464 4256
rect 3487 4256 3533 4264
rect 3656 4264 3664 4273
rect 3656 4256 3973 4264
rect 4027 4256 4253 4264
rect 4267 4256 4313 4264
rect 4407 4256 4493 4264
rect 4607 4256 4693 4264
rect 4827 4256 4853 4264
rect 4896 4256 4973 4264
rect 3367 4236 3424 4244
rect 3456 4236 3533 4244
rect 1667 4216 1773 4224
rect 1787 4216 1973 4224
rect 2207 4216 2573 4224
rect 3227 4216 3293 4224
rect 3307 4216 3373 4224
rect 3416 4224 3424 4236
rect 3907 4236 3933 4244
rect 4547 4236 4633 4244
rect 4896 4244 4904 4256
rect 5447 4256 5493 4264
rect 5567 4256 5633 4264
rect 5907 4256 5953 4264
rect 4727 4236 4904 4244
rect 5007 4236 5133 4244
rect 3416 4216 4433 4224
rect 4967 4216 5033 4224
rect 5387 4216 5853 4224
rect 167 4196 633 4204
rect 927 4196 953 4204
rect 1187 4196 1273 4204
rect 2847 4196 2913 4204
rect 3267 4196 3513 4204
rect 3607 4196 3833 4204
rect 4287 4196 4353 4204
rect 4547 4196 4853 4204
rect 4947 4196 5053 4204
rect 5127 4196 5293 4204
rect 5807 4196 5833 4204
rect 5847 4196 5873 4204
rect 27 4176 853 4184
rect 1147 4176 1733 4184
rect 2387 4176 2653 4184
rect 2867 4176 3133 4184
rect 4067 4176 4213 4184
rect 4987 4176 5053 4184
rect 287 4156 573 4164
rect 2347 4156 2473 4164
rect 2496 4156 2753 4164
rect 107 4136 613 4144
rect 787 4136 833 4144
rect 1107 4136 1473 4144
rect 1487 4136 1553 4144
rect 2496 4144 2504 4156
rect 2927 4156 3673 4164
rect 3907 4156 4093 4164
rect 4327 4156 4713 4164
rect 4987 4156 5973 4164
rect 1907 4136 2504 4144
rect 2627 4136 2713 4144
rect 2727 4136 2833 4144
rect 2907 4136 3693 4144
rect 4247 4136 4453 4144
rect 4767 4136 4793 4144
rect 4847 4136 4953 4144
rect 5016 4136 5133 4144
rect 647 4116 973 4124
rect 1067 4116 1233 4124
rect 3027 4116 3173 4124
rect 3247 4116 3653 4124
rect 3927 4116 3993 4124
rect 4007 4116 4153 4124
rect 4227 4116 4633 4124
rect 5016 4124 5024 4136
rect 5267 4136 5813 4144
rect 4707 4116 5024 4124
rect 5307 4116 5373 4124
rect 5387 4116 5453 4124
rect 547 4096 573 4104
rect 867 4096 1893 4104
rect 1947 4096 2393 4104
rect 2407 4096 2833 4104
rect 2847 4096 2893 4104
rect 2987 4096 3793 4104
rect 3807 4096 4653 4104
rect 4907 4096 5093 4104
rect 5107 4096 5293 4104
rect 5307 4096 5413 4104
rect 5747 4096 5833 4104
rect 5847 4096 5913 4104
rect 1047 4076 1253 4084
rect 1447 4076 1533 4084
rect 2567 4076 2813 4084
rect 2827 4076 2873 4084
rect 3656 4076 3733 4084
rect 427 4056 1093 4064
rect 1247 4056 1313 4064
rect 1587 4056 1653 4064
rect 2167 4056 2313 4064
rect 2327 4056 2533 4064
rect 3367 4056 3573 4064
rect 3656 4064 3664 4076
rect 3987 4076 4033 4084
rect 4047 4076 4252 4084
rect 4287 4076 4373 4084
rect 4607 4076 4973 4084
rect 5187 4076 5273 4084
rect 3636 4056 3664 4064
rect 96 4036 173 4044
rect 96 3987 104 4036
rect 627 4036 664 4044
rect 187 3996 213 4004
rect 656 4006 664 4036
rect 687 4037 733 4045
rect 1387 4039 1433 4047
rect 2936 4036 3013 4044
rect 796 4004 804 4034
rect 707 3996 804 4004
rect 827 3996 893 4004
rect 1007 3995 1033 4003
rect 1047 3996 1073 4004
rect 1147 3995 1173 4003
rect 1187 3995 1393 4003
rect 1447 3996 1633 4004
rect 2116 4004 2124 4034
rect 2116 3996 2173 4004
rect 2396 3987 2404 4034
rect 2936 4024 2944 4036
rect 2816 4016 2944 4024
rect 2507 3995 2553 4003
rect 2667 3996 2753 4004
rect 2816 4004 2824 4016
rect 2767 3996 2824 4004
rect 3156 3987 3164 4034
rect 3316 4004 3324 4036
rect 3456 4004 3464 4033
rect 3187 3996 3324 4004
rect 3447 3996 3464 4004
rect 3636 4004 3644 4056
rect 4567 4056 4624 4064
rect 3607 3996 3644 4004
rect 1427 3976 1673 3984
rect 1687 3976 1713 3984
rect 2227 3976 2304 3984
rect 207 3956 373 3964
rect 387 3956 693 3964
rect 1527 3956 1593 3964
rect 1807 3956 1953 3964
rect 1967 3956 2084 3964
rect 127 3936 133 3944
rect 147 3936 333 3944
rect 347 3936 493 3944
rect 747 3936 1013 3944
rect 2076 3944 2084 3956
rect 2116 3956 2153 3964
rect 2116 3944 2124 3956
rect 2296 3964 2304 3976
rect 2927 3976 2973 3984
rect 2987 3976 3053 3984
rect 3487 3976 3513 3984
rect 3676 3984 3684 4036
rect 3807 4036 4013 4044
rect 4027 4037 4193 4045
rect 4496 4036 4533 4044
rect 4276 4024 4284 4034
rect 3787 4016 4284 4024
rect 3856 4004 3864 4016
rect 4007 3996 4073 4004
rect 4316 4004 4324 4034
rect 4187 3996 4373 4004
rect 4193 3987 4207 3996
rect 4416 4004 4424 4034
rect 4416 3996 4473 4004
rect 3676 3976 3733 3984
rect 4267 3976 4313 3984
rect 4496 3984 4504 4036
rect 4616 4007 4624 4056
rect 5007 4056 5053 4064
rect 5327 4056 5493 4064
rect 4716 4036 4733 4044
rect 4716 4007 4724 4036
rect 4887 4036 5092 4044
rect 5113 4024 5127 4033
rect 5036 4020 5127 4024
rect 5216 4024 5224 4034
rect 5367 4036 5393 4044
rect 5293 4024 5307 4033
rect 5216 4020 5244 4024
rect 5293 4020 5324 4024
rect 5036 4016 5124 4020
rect 5216 4016 5247 4020
rect 5296 4016 5324 4020
rect 4667 3995 4692 4003
rect 5036 4006 5044 4016
rect 5233 4007 5247 4016
rect 4867 3995 4893 4003
rect 5316 4006 5324 4016
rect 4447 3976 4504 3984
rect 4567 3976 4633 3984
rect 5236 3984 5244 3993
rect 5436 4004 5444 4033
rect 5596 4007 5604 4034
rect 5367 3996 5444 4004
rect 5456 3996 5513 4004
rect 4967 3976 5024 3984
rect 2296 3956 2413 3964
rect 3247 3956 3533 3964
rect 4127 3956 4173 3964
rect 4247 3956 4293 3964
rect 4487 3956 4533 3964
rect 4727 3956 4833 3964
rect 4907 3956 4933 3964
rect 5016 3964 5024 3976
rect 5096 3976 5244 3984
rect 5096 3964 5104 3976
rect 5456 3984 5464 3996
rect 5587 3996 5604 4007
rect 5587 3993 5600 3996
rect 5427 3976 5464 3984
rect 5636 3967 5644 4034
rect 5687 4036 5713 4044
rect 5987 4036 6024 4044
rect 5667 3996 5693 4004
rect 5756 4004 5764 4033
rect 5856 4007 5864 4033
rect 5756 3996 5813 4004
rect 5887 3976 5973 3984
rect 5016 3956 5104 3964
rect 5167 3956 5253 3964
rect 5627 3956 5644 3967
rect 5627 3953 5640 3956
rect 5787 3956 5813 3964
rect 2076 3936 2124 3944
rect 2207 3936 2273 3944
rect 2287 3936 2593 3944
rect 3256 3936 3933 3944
rect 547 3916 573 3924
rect 1447 3916 1533 3924
rect 1587 3916 1653 3924
rect 1927 3916 1993 3924
rect 2007 3916 2053 3924
rect 2067 3916 2133 3924
rect 3256 3924 3264 3936
rect 4147 3936 4213 3944
rect 4467 3936 4513 3944
rect 4527 3936 4813 3944
rect 5007 3936 5073 3944
rect 5087 3936 5193 3944
rect 5487 3936 5512 3944
rect 5547 3936 5633 3944
rect 5907 3936 5953 3944
rect 2716 3916 3264 3924
rect 407 3896 1793 3904
rect 2587 3896 2693 3904
rect 2716 3904 2724 3916
rect 3647 3916 3793 3924
rect 3967 3916 4853 3924
rect 5567 3916 5593 3924
rect 2707 3896 2724 3904
rect 3567 3896 3753 3904
rect 4447 3896 4473 3904
rect 4547 3896 4753 3904
rect 4927 3896 5013 3904
rect 5107 3896 5193 3904
rect 5247 3896 5373 3904
rect 5527 3896 5753 3904
rect 5807 3896 5933 3904
rect 567 3876 673 3884
rect 687 3876 713 3884
rect 1227 3876 1273 3884
rect 1287 3876 1333 3884
rect 3407 3876 3893 3884
rect 4407 3876 4493 3884
rect 4607 3876 4653 3884
rect 4827 3876 5033 3884
rect 5047 3876 5213 3884
rect 5467 3876 5773 3884
rect -24 3856 153 3864
rect 207 3856 293 3864
rect 587 3856 653 3864
rect 867 3856 973 3864
rect 1907 3856 2693 3864
rect 2787 3856 3313 3864
rect 3627 3856 3864 3864
rect 367 3836 413 3844
rect 607 3836 633 3844
rect 1127 3836 1173 3844
rect 1187 3836 1273 3844
rect 1827 3836 1853 3844
rect 3307 3836 3333 3844
rect 3856 3844 3864 3856
rect 4056 3856 4133 3864
rect 4056 3847 4064 3856
rect 4596 3856 4673 3864
rect 3856 3836 3893 3844
rect 3956 3836 4053 3844
rect -24 3816 13 3824
rect 107 3816 244 3824
rect -24 3776 13 3784
rect 236 3786 244 3816
rect 267 3816 304 3824
rect 296 3807 304 3816
rect 327 3816 413 3824
rect 467 3816 624 3824
rect 296 3806 320 3807
rect 296 3796 313 3806
rect 300 3793 313 3796
rect 616 3804 624 3816
rect 707 3816 824 3824
rect 816 3804 824 3816
rect 1067 3816 1093 3824
rect 2247 3816 2273 3824
rect 2607 3816 2633 3824
rect 2847 3817 2893 3825
rect 3007 3816 3093 3824
rect 616 3796 744 3804
rect 816 3796 884 3804
rect 736 3786 744 3796
rect 876 3786 884 3796
rect 287 3775 333 3783
rect 387 3775 433 3783
rect 956 3784 964 3813
rect 956 3776 1153 3784
rect 1196 3767 1204 3813
rect 1236 3784 1244 3813
rect 1236 3776 1293 3784
rect 1307 3776 1593 3784
rect 1607 3776 1633 3784
rect 1827 3775 1993 3783
rect 2636 3784 2644 3814
rect 3427 3816 3513 3824
rect 3576 3804 3584 3814
rect 3847 3816 3933 3824
rect 3956 3824 3964 3836
rect 4367 3844 4380 3847
rect 4367 3833 4384 3844
rect 3947 3816 3964 3824
rect 4087 3817 4153 3825
rect 4227 3816 4273 3824
rect 3576 3796 3684 3804
rect 3676 3787 3684 3796
rect 3736 3787 3744 3813
rect 4336 3787 4344 3813
rect 4376 3787 4384 3833
rect 4507 3817 4573 3825
rect 4596 3804 4604 3856
rect 5287 3856 5333 3864
rect 5507 3856 5533 3864
rect 5607 3856 5673 3864
rect 4927 3836 5064 3844
rect 4667 3816 4893 3824
rect 4476 3796 4604 3804
rect 2636 3776 2733 3784
rect 2887 3775 2913 3783
rect 3187 3776 3213 3784
rect 3227 3776 3313 3784
rect 3527 3775 3553 3783
rect 3676 3776 3693 3787
rect 3680 3773 3693 3776
rect 3907 3775 3953 3783
rect 4476 3784 4484 3796
rect 4816 3786 4824 3816
rect 5056 3824 5064 3836
rect 5187 3836 5233 3844
rect 5327 3836 5373 3844
rect 5647 3836 5793 3844
rect 5056 3816 5073 3824
rect 5087 3816 5133 3824
rect 4956 3804 4964 3814
rect 5196 3816 5253 3824
rect 4956 3796 5173 3804
rect 4456 3776 4484 3784
rect 647 3756 673 3764
rect 687 3756 833 3764
rect 1007 3756 1073 3764
rect 1187 3756 1204 3767
rect 1187 3753 1200 3756
rect 1587 3756 1773 3764
rect 1787 3756 2193 3764
rect 3016 3764 3024 3772
rect 2967 3756 3153 3764
rect 3167 3756 3433 3764
rect 4456 3764 4464 3776
rect 4647 3775 4693 3783
rect 5076 3776 5133 3784
rect 3867 3756 4464 3764
rect 5076 3764 5084 3776
rect 5196 3767 5204 3816
rect 5307 3817 5393 3825
rect 5287 3776 5433 3784
rect 5516 3784 5524 3813
rect 5576 3804 5584 3833
rect 5556 3800 5584 3804
rect 5447 3776 5524 3784
rect 5553 3796 5584 3800
rect 5656 3816 5713 3824
rect 5553 3787 5567 3796
rect 5656 3787 5664 3816
rect 4987 3756 5084 3764
rect 5196 3766 5220 3767
rect 5196 3764 5213 3766
rect 5127 3756 5213 3764
rect 5200 3753 5213 3756
rect 67 3736 373 3744
rect 1547 3736 2073 3744
rect 2187 3736 2373 3744
rect 2587 3736 2613 3744
rect 2687 3736 3133 3744
rect 3147 3744 3160 3747
rect 3147 3733 3164 3744
rect 27 3716 373 3724
rect 2367 3716 2413 3724
rect 2707 3716 2973 3724
rect 3156 3724 3164 3733
rect 3336 3736 3393 3744
rect 3336 3724 3344 3736
rect 3436 3744 3444 3753
rect 5387 3756 5473 3764
rect 5487 3756 5593 3764
rect 5747 3756 5873 3764
rect 3436 3736 3593 3744
rect 3667 3736 3733 3744
rect 3787 3736 4233 3744
rect 4367 3736 4573 3744
rect 4787 3736 4833 3744
rect 4947 3736 5033 3744
rect 5107 3736 5233 3744
rect 3156 3716 3344 3724
rect 3367 3716 3553 3724
rect 267 3696 313 3704
rect 1427 3696 1613 3704
rect 1747 3696 1933 3704
rect 2356 3704 2364 3713
rect 3653 3724 3667 3733
rect 3607 3720 3667 3724
rect 3607 3716 3664 3720
rect 4067 3716 4112 3724
rect 4147 3716 4493 3724
rect 4507 3716 4533 3724
rect 4547 3716 4673 3724
rect 5007 3716 5173 3724
rect 5187 3716 5353 3724
rect 5427 3716 5653 3724
rect 5787 3716 5833 3724
rect 1947 3696 2364 3704
rect 2467 3696 2613 3704
rect 2847 3696 3113 3704
rect 3207 3696 4084 3704
rect 4076 3687 4084 3696
rect 4367 3696 4973 3704
rect 5147 3696 5193 3704
rect 5587 3696 5633 3704
rect 387 3676 2673 3684
rect 2987 3676 3273 3684
rect 3367 3676 3472 3684
rect 3507 3676 3613 3684
rect 4087 3676 4213 3684
rect 4227 3676 4993 3684
rect 5047 3676 5113 3684
rect 5267 3676 5393 3684
rect 367 3656 773 3664
rect 1107 3656 1193 3664
rect 1267 3656 1313 3664
rect 1687 3656 1733 3664
rect 2607 3656 2953 3664
rect 4167 3656 4433 3664
rect 4447 3656 4473 3664
rect 4547 3656 4773 3664
rect 4967 3656 5113 3664
rect 5687 3656 5893 3664
rect 227 3636 2453 3644
rect 2467 3636 3033 3644
rect 3087 3636 4753 3644
rect 5107 3636 5153 3644
rect 5227 3636 5393 3644
rect 5487 3636 5693 3644
rect 47 3616 553 3624
rect 667 3616 753 3624
rect 1187 3616 1413 3624
rect 2627 3616 2933 3624
rect 3107 3616 3133 3624
rect 3247 3616 3313 3624
rect 4887 3616 4913 3624
rect 4927 3616 5033 3624
rect 5287 3616 5413 3624
rect 187 3596 513 3604
rect 987 3596 1573 3604
rect 1887 3596 2093 3604
rect 2107 3596 2593 3604
rect 3127 3596 3213 3604
rect 3567 3596 3853 3604
rect 3927 3596 4193 3604
rect 4587 3596 5073 3604
rect 5087 3596 5153 3604
rect 5167 3596 5253 3604
rect 5507 3596 5853 3604
rect 456 3576 593 3584
rect 76 3536 113 3544
rect 76 3486 84 3536
rect 147 3517 173 3525
rect 96 3484 104 3514
rect 96 3476 273 3484
rect 456 3447 464 3576
rect 747 3576 833 3584
rect 927 3576 1293 3584
rect 1767 3576 1853 3584
rect 2247 3576 2273 3584
rect 2407 3576 2493 3584
rect 2507 3576 2584 3584
rect 476 3556 613 3564
rect 476 3467 484 3556
rect 747 3556 1193 3564
rect 1207 3556 1253 3564
rect 1387 3556 1493 3564
rect 1847 3556 2033 3564
rect 2087 3556 2333 3564
rect 2576 3564 2584 3576
rect 2687 3576 2873 3584
rect 3067 3576 3293 3584
rect 3387 3576 3473 3584
rect 4687 3576 5053 3584
rect 5127 3576 5273 3584
rect 2576 3556 2813 3564
rect 3187 3556 3453 3564
rect 3507 3556 3553 3564
rect 4187 3556 4273 3564
rect 4607 3556 4633 3564
rect 5307 3556 5413 3564
rect 5547 3556 5653 3564
rect 5767 3556 5853 3564
rect 1547 3536 1573 3544
rect 2567 3536 2713 3544
rect 496 3520 513 3524
rect 493 3516 513 3520
rect 493 3506 507 3516
rect 527 3516 593 3524
rect 620 3524 633 3527
rect 616 3513 633 3524
rect 687 3516 773 3524
rect 816 3516 973 3524
rect 616 3504 624 3513
rect 536 3496 624 3504
rect 536 3484 544 3496
rect 816 3486 824 3516
rect 1027 3517 1132 3525
rect 1167 3516 1193 3524
rect 1473 3524 1487 3533
rect 3047 3536 3133 3544
rect 4027 3536 4393 3544
rect 4947 3536 5013 3544
rect 1473 3520 1524 3524
rect 1476 3516 1524 3520
rect 1516 3486 1524 3516
rect 1607 3516 1693 3524
rect 1707 3516 1793 3524
rect 1967 3516 2204 3524
rect 2196 3507 2204 3516
rect 2196 3496 2213 3507
rect 2200 3493 2213 3496
rect 2276 3487 2284 3516
rect 2507 3517 2533 3525
rect 2756 3504 2764 3514
rect 3227 3517 3253 3525
rect 3307 3516 3333 3524
rect 3387 3516 3424 3524
rect 2667 3496 2764 3504
rect 927 3476 993 3484
rect 1327 3475 1353 3483
rect 1687 3476 1893 3484
rect 2267 3476 2284 3487
rect 2267 3473 2280 3476
rect 2427 3476 2633 3484
rect 2687 3476 2733 3484
rect 2756 3484 2764 3496
rect 3156 3487 3164 3513
rect 2756 3476 2793 3484
rect 2947 3473 2993 3481
rect 3067 3476 3113 3484
rect 3416 3486 3424 3516
rect 3496 3504 3504 3516
rect 3747 3516 3793 3524
rect 4187 3516 4264 3524
rect 3496 3496 3593 3504
rect 4136 3504 4144 3514
rect 3956 3496 4144 3504
rect 3467 3475 3593 3483
rect 3687 3473 3713 3481
rect 3956 3484 3964 3496
rect 4256 3486 4264 3516
rect 4287 3516 4313 3524
rect 4336 3516 4373 3524
rect 3827 3476 3964 3484
rect 4336 3484 4344 3516
rect 4307 3476 4344 3484
rect 4436 3467 4444 3514
rect 4496 3487 4504 3513
rect 4556 3486 4564 3533
rect 4727 3516 4784 3524
rect 4776 3487 4784 3516
rect 5127 3517 5293 3525
rect 4956 3487 4964 3513
rect 5336 3487 5344 3514
rect 5407 3516 5444 3524
rect 5436 3487 5444 3516
rect 5707 3517 5793 3525
rect 5807 3516 5973 3524
rect 5496 3487 5504 3513
rect 5576 3487 5584 3513
rect 5616 3504 5624 3514
rect 5616 3496 5784 3504
rect 4647 3475 4673 3483
rect 4776 3476 4793 3487
rect 4780 3473 4793 3476
rect 5187 3475 5233 3483
rect 5247 3475 5273 3483
rect 5336 3476 5353 3487
rect 5340 3473 5353 3476
rect 5776 3467 5784 3496
rect 476 3466 500 3467
rect 476 3456 493 3466
rect 480 3453 493 3456
rect 1627 3456 1653 3464
rect 2547 3456 2653 3464
rect 5407 3456 5553 3464
rect 5567 3456 5732 3464
rect 5767 3456 5784 3467
rect 5767 3453 5780 3456
rect 187 3436 333 3444
rect 456 3436 473 3447
rect 460 3433 473 3436
rect 787 3436 853 3444
rect 947 3436 1193 3444
rect 1367 3436 1413 3444
rect 1487 3436 1593 3444
rect 1687 3436 1873 3444
rect 1927 3436 1993 3444
rect 2127 3436 2353 3444
rect 4127 3436 4484 3444
rect 427 3416 493 3424
rect 1307 3416 1533 3424
rect 1707 3416 1753 3424
rect 3316 3416 3333 3424
rect 1587 3396 1813 3404
rect 2267 3396 2313 3404
rect 2607 3396 2793 3404
rect 3316 3404 3324 3416
rect 3347 3416 3373 3424
rect 3767 3416 3873 3424
rect 4176 3416 4333 3424
rect 4176 3407 4184 3416
rect 4427 3424 4440 3427
rect 4476 3424 4484 3436
rect 4807 3436 5013 3444
rect 5027 3436 5193 3444
rect 5527 3436 5593 3444
rect 4427 3413 4444 3424
rect 4476 3416 4633 3424
rect 4687 3416 4753 3424
rect 4947 3416 4993 3424
rect 5187 3416 5213 3424
rect 2907 3396 3324 3404
rect 3987 3396 4173 3404
rect 4436 3404 4444 3413
rect 4436 3396 4613 3404
rect 5147 3396 5353 3404
rect 5367 3396 5453 3404
rect 207 3376 253 3384
rect 1147 3376 2133 3384
rect 2147 3376 2193 3384
rect 2407 3376 2473 3384
rect 3287 3376 3333 3384
rect 3427 3376 3493 3384
rect 3567 3376 3773 3384
rect 3947 3376 4233 3384
rect 4567 3376 4773 3384
rect 4947 3376 5333 3384
rect 5347 3376 5373 3384
rect 5487 3376 5573 3384
rect 5667 3376 5853 3384
rect 1167 3356 1233 3364
rect 1307 3356 1453 3364
rect 1527 3356 1673 3364
rect 2627 3356 2733 3364
rect 3067 3356 3473 3364
rect 3487 3356 3933 3364
rect 3987 3356 4033 3364
rect 4087 3356 4193 3364
rect 4287 3356 4333 3364
rect 4447 3356 4513 3364
rect 4587 3356 4653 3364
rect 4707 3356 5113 3364
rect 5427 3356 5553 3364
rect 5707 3356 5813 3364
rect 807 3336 1053 3344
rect 1067 3336 1133 3344
rect 1407 3336 1433 3344
rect 1607 3336 1652 3344
rect 1687 3336 1753 3344
rect 2367 3336 2653 3344
rect 2787 3336 2893 3344
rect 2967 3336 3013 3344
rect 3507 3336 3653 3344
rect 3787 3336 3913 3344
rect 3967 3336 4473 3344
rect 4487 3336 4713 3344
rect 4827 3336 5093 3344
rect 5327 3336 5393 3344
rect 787 3316 893 3324
rect 1387 3316 1733 3324
rect 1747 3316 1793 3324
rect 2167 3316 2213 3324
rect 2747 3316 2853 3324
rect 2996 3316 3033 3324
rect 227 3299 273 3307
rect 107 3253 133 3261
rect 287 3256 313 3264
rect 367 3256 473 3264
rect 556 3264 564 3296
rect 647 3296 753 3304
rect 776 3296 853 3304
rect 776 3284 784 3296
rect 967 3296 993 3304
rect 1047 3296 1073 3304
rect 1227 3296 1333 3304
rect 1427 3296 1513 3304
rect 1607 3296 1744 3304
rect 1847 3299 1913 3307
rect 2020 3304 2033 3307
rect 627 3276 784 3284
rect 527 3256 564 3264
rect 647 3253 673 3261
rect 887 3256 1013 3264
rect 1087 3255 1153 3263
rect 1167 3256 1273 3264
rect 1407 3255 1492 3263
rect 1527 3255 1573 3263
rect 1647 3256 1673 3264
rect 1736 3266 1744 3296
rect 2016 3293 2033 3304
rect 2727 3296 2844 3304
rect 2016 3264 2024 3293
rect 2196 3267 2204 3293
rect 2267 3276 2344 3284
rect 2027 3260 2124 3264
rect 2027 3256 2127 3260
rect 2113 3247 2127 3256
rect 2336 3266 2344 3276
rect 2356 3267 2364 3294
rect 2356 3256 2373 3267
rect 2360 3253 2373 3256
rect 2836 3266 2844 3296
rect 2487 3253 2573 3261
rect 2887 3256 2933 3264
rect 2996 3266 3004 3316
rect 3076 3316 3153 3324
rect 3076 3304 3084 3316
rect 3507 3316 3924 3324
rect 3036 3296 3084 3304
rect 3207 3299 3273 3307
rect 3036 3266 3044 3296
rect 3396 3296 3553 3304
rect 3356 3267 3364 3293
rect 3396 3266 3404 3296
rect 3847 3296 3873 3304
rect 3916 3304 3924 3316
rect 4116 3316 4293 3324
rect 3916 3296 4013 3304
rect 4027 3296 4093 3304
rect 3713 3284 3727 3293
rect 3713 3280 3893 3284
rect 3716 3276 3893 3280
rect 4116 3284 4124 3316
rect 5027 3316 5053 3324
rect 5167 3316 5404 3324
rect 4247 3304 4260 3307
rect 4247 3293 4264 3304
rect 4327 3297 4413 3305
rect 4467 3296 4633 3304
rect 4767 3296 4844 3304
rect 4036 3280 4124 3284
rect 4033 3276 4124 3280
rect 4033 3267 4047 3276
rect 4176 3267 4184 3293
rect 3407 3256 3513 3264
rect 4256 3266 4264 3293
rect 4836 3284 4844 3296
rect 4867 3297 4893 3305
rect 5396 3304 5404 3316
rect 5567 3316 5693 3324
rect 5787 3316 5833 3324
rect 5396 3296 5413 3304
rect 5547 3296 5593 3304
rect 5696 3296 5732 3304
rect 4836 3276 4884 3284
rect 4347 3255 4433 3263
rect 4447 3256 4553 3264
rect 4607 3255 4633 3263
rect 4876 3266 4884 3276
rect 5036 3267 5044 3293
rect 4687 3256 4733 3264
rect 5136 3264 5144 3293
rect 5176 3267 5184 3293
rect 5496 3267 5504 3293
rect 5136 3256 5164 3264
rect 5156 3247 5164 3256
rect 5247 3256 5433 3264
rect 5656 3264 5664 3293
rect 5587 3256 5664 3264
rect 5696 3247 5704 3296
rect 5887 3296 5913 3304
rect 5756 3264 5764 3293
rect 5756 3256 5813 3264
rect 5987 3256 6024 3264
rect 47 3236 733 3244
rect 1367 3236 1464 3244
rect 1247 3216 1433 3224
rect 1456 3224 1464 3236
rect 1807 3236 2064 3244
rect 1456 3216 1753 3224
rect 2056 3224 2064 3236
rect 2227 3236 2293 3244
rect 3547 3236 3753 3244
rect 3767 3236 3853 3244
rect 3867 3236 4233 3244
rect 4927 3236 5133 3244
rect 5156 3246 5180 3247
rect 5156 3236 5173 3246
rect 5160 3233 5173 3236
rect 5267 3236 5313 3244
rect 2056 3216 2453 3224
rect 2527 3216 2613 3224
rect 2707 3216 2873 3224
rect 2967 3216 3153 3224
rect 3347 3216 3433 3224
rect 3627 3216 3813 3224
rect 3927 3216 3993 3224
rect 4007 3216 4113 3224
rect 4787 3216 5053 3224
rect 5107 3216 5193 3224
rect 5387 3216 5553 3224
rect 5647 3216 5773 3224
rect 107 3196 1793 3204
rect 1967 3196 2033 3204
rect 2667 3196 2733 3204
rect 4247 3196 4473 3204
rect 4667 3196 5233 3204
rect 5567 3196 5973 3204
rect 1327 3176 1373 3184
rect 1387 3176 1613 3184
rect 1707 3176 1773 3184
rect 2087 3176 2133 3184
rect 2147 3176 2173 3184
rect 2187 3176 2253 3184
rect 2807 3176 3293 3184
rect 4227 3176 4333 3184
rect 4347 3176 4613 3184
rect 4727 3176 5173 3184
rect 5227 3176 5533 3184
rect 5607 3176 5833 3184
rect 2007 3156 2053 3164
rect 2487 3156 2813 3164
rect 3367 3156 3633 3164
rect 3707 3156 5024 3164
rect 1187 3136 1313 3144
rect 2047 3136 2313 3144
rect 2427 3136 2853 3144
rect 3727 3136 4493 3144
rect 4847 3136 4973 3144
rect 5016 3144 5024 3156
rect 5047 3156 5093 3164
rect 5107 3156 5153 3164
rect 5207 3156 5273 3164
rect 5016 3136 5553 3144
rect 5627 3136 5973 3144
rect 1927 3116 2013 3124
rect 2467 3116 2693 3124
rect 3307 3116 3493 3124
rect 3827 3116 3893 3124
rect 3947 3116 4673 3124
rect 5347 3116 5413 3124
rect 5747 3116 5913 3124
rect 1547 3096 1593 3104
rect 1747 3096 2113 3104
rect 2387 3096 2473 3104
rect 2647 3096 2693 3104
rect 2787 3096 2913 3104
rect 3687 3096 3733 3104
rect 4007 3096 4173 3104
rect 4187 3096 4313 3104
rect 5007 3096 5213 3104
rect 5547 3096 5633 3104
rect 5647 3096 5673 3104
rect 5847 3096 5933 3104
rect 1907 3076 2133 3084
rect 3327 3076 3373 3084
rect 3607 3076 3793 3084
rect 3807 3076 4513 3084
rect 4527 3076 4652 3084
rect 4687 3076 4853 3084
rect 4867 3076 5193 3084
rect 5407 3076 5453 3084
rect 5667 3076 5813 3084
rect 5827 3076 5873 3084
rect 927 3056 973 3064
rect 1407 3056 1473 3064
rect 2156 3056 2213 3064
rect 47 3036 153 3044
rect 1047 3036 1333 3044
rect 2156 3044 2164 3056
rect 3367 3056 3533 3064
rect 3627 3056 3713 3064
rect 3787 3056 3853 3064
rect 4087 3056 4393 3064
rect 4927 3056 4953 3064
rect 5067 3056 5373 3064
rect 5507 3056 5553 3064
rect 2027 3036 2164 3044
rect 2347 3036 2413 3044
rect 2827 3036 3073 3044
rect 3087 3036 3173 3044
rect 3187 3036 3213 3044
rect 3327 3036 4053 3044
rect 4447 3036 4513 3044
rect 4587 3036 4893 3044
rect 5136 3036 5472 3044
rect 387 3016 433 3024
rect 527 3016 573 3024
rect 1447 3016 1613 3024
rect 1627 3016 1653 3024
rect 1667 3016 1813 3024
rect 2196 3016 2233 3024
rect -24 2996 72 3004
rect 107 2999 133 3007
rect 227 2953 273 2961
rect 336 2947 344 2994
rect 467 2996 493 3004
rect 967 2997 1033 3005
rect 1247 2997 1293 3005
rect 1356 2996 1433 3004
rect 407 2955 453 2963
rect 947 2955 1013 2963
rect 1356 2966 1364 2996
rect 1867 2997 1973 3005
rect 1516 2967 1524 2993
rect 1027 2955 1053 2963
rect 1607 2956 1893 2964
rect 2036 2964 2044 2996
rect 2196 2967 2204 3016
rect 2687 3016 2733 3024
rect 3647 3016 3913 3024
rect 2567 2996 2724 3004
rect 3127 2996 3213 3004
rect 2376 2984 2384 2994
rect 2296 2976 2384 2984
rect 2036 2956 2113 2964
rect 2296 2964 2304 2976
rect 2716 2967 2724 2996
rect 3427 2996 3553 3004
rect 3747 2996 3933 3004
rect 3956 2996 3973 3004
rect 3556 2984 3564 2994
rect 3956 2984 3964 2996
rect 4027 2996 4113 3004
rect 4287 2996 4352 3004
rect 4386 2993 4387 3000
rect 4407 2997 4493 3005
rect 4507 2996 4533 3004
rect 4636 2996 4753 3004
rect 4373 2984 4387 2993
rect 4636 2984 4644 2996
rect 4856 2996 4984 3004
rect 3556 2976 3964 2984
rect 4236 2980 4387 2984
rect 4233 2976 4383 2980
rect 4616 2976 4644 2984
rect 4233 2967 4247 2976
rect 2247 2956 2304 2964
rect 2327 2956 2393 2964
rect 2507 2956 2533 2964
rect 2547 2956 2613 2964
rect 2947 2953 2993 2961
rect 4246 2960 4247 2967
rect 4267 2956 4293 2964
rect 4307 2956 4413 2964
rect 4616 2964 4624 2976
rect 4856 2967 4864 2996
rect 4976 2984 4984 2996
rect 5016 2996 5053 3004
rect 5016 2984 5024 2996
rect 4976 2976 5024 2984
rect 5136 2967 5144 3036
rect 5507 3036 5693 3044
rect 5467 3016 5673 3024
rect 5727 3016 5913 3024
rect 5447 2997 5493 3005
rect 5547 2997 5593 3005
rect 5647 2996 5684 3004
rect 5216 2967 5224 2993
rect 4607 2956 4624 2964
rect 4667 2955 4693 2963
rect 4847 2956 4864 2967
rect 4847 2953 4860 2956
rect 4967 2956 5033 2964
rect 5676 2966 5684 2996
rect 5787 2996 5804 3004
rect 5736 2967 5744 2993
rect 5567 2956 5673 2964
rect 5796 2964 5804 2996
rect 5956 2967 5964 2993
rect 5796 2956 5893 2964
rect 547 2936 1133 2944
rect 2287 2936 2433 2944
rect 2487 2936 2533 2944
rect 767 2916 873 2924
rect 1167 2916 1213 2924
rect 1267 2916 1453 2924
rect 1913 2924 1927 2933
rect 3447 2936 3633 2944
rect 3727 2936 3753 2944
rect 3767 2936 3793 2944
rect 3807 2936 3973 2944
rect 4067 2936 4133 2944
rect 4327 2936 4453 2944
rect 5127 2936 5173 2944
rect 5187 2936 5433 2944
rect 1913 2920 1993 2924
rect 1916 2916 1993 2920
rect 2007 2916 2253 2924
rect 2467 2916 3253 2924
rect 4747 2916 4913 2924
rect 5847 2916 5953 2924
rect 147 2896 353 2904
rect 1247 2896 1833 2904
rect 2147 2896 2393 2904
rect 2887 2896 3233 2904
rect 3487 2896 3593 2904
rect 3907 2896 4293 2904
rect 4607 2896 5273 2904
rect 5487 2896 5552 2904
rect 5587 2896 5813 2904
rect 667 2876 973 2884
rect 987 2876 1213 2884
rect 1987 2876 2493 2884
rect 5087 2876 5193 2884
rect 5636 2876 5873 2884
rect 5636 2867 5644 2876
rect 1407 2856 1573 2864
rect 1787 2856 1973 2864
rect 2587 2856 2833 2864
rect 2847 2856 2984 2864
rect 687 2836 733 2844
rect 1627 2836 1733 2844
rect 2847 2836 2953 2844
rect 2976 2844 2984 2856
rect 3067 2856 3393 2864
rect 3847 2856 4093 2864
rect 4107 2856 4132 2864
rect 4167 2856 4373 2864
rect 4787 2856 4933 2864
rect 4987 2856 5093 2864
rect 5347 2856 5373 2864
rect 5387 2856 5633 2864
rect 5707 2856 5973 2864
rect 2976 2836 3133 2844
rect 3227 2836 3473 2844
rect 3647 2836 3813 2844
rect 4547 2836 4793 2844
rect 4807 2836 4833 2844
rect 5527 2836 5593 2844
rect 147 2816 493 2824
rect 567 2816 713 2824
rect 1007 2816 1313 2824
rect 2047 2816 2333 2824
rect 2447 2816 2573 2824
rect 2947 2816 3353 2824
rect 3507 2816 4193 2824
rect 4367 2816 4413 2824
rect 4507 2816 4593 2824
rect 5027 2816 5393 2824
rect 5447 2816 5613 2824
rect 5687 2816 5733 2824
rect 5927 2816 6004 2824
rect 607 2796 693 2804
rect 2207 2796 2233 2804
rect 2547 2796 2613 2804
rect 2987 2796 3213 2804
rect 3227 2796 3273 2804
rect 3967 2804 3980 2807
rect 3967 2793 3984 2804
rect 4087 2796 4113 2804
rect 4447 2796 4852 2804
rect 4887 2796 4933 2804
rect 5067 2796 5152 2804
rect 5187 2796 5264 2804
rect 216 2764 224 2776
rect 627 2776 653 2784
rect 1027 2779 1073 2787
rect 1327 2777 1353 2785
rect 1407 2776 1432 2784
rect 1467 2776 1513 2784
rect 1567 2777 1633 2785
rect 216 2756 753 2764
rect 107 2733 133 2741
rect 287 2736 313 2744
rect 367 2735 392 2743
rect 427 2735 473 2743
rect 527 2735 553 2743
rect 687 2735 733 2743
rect 967 2736 993 2744
rect 1107 2735 1193 2743
rect 1247 2736 1313 2744
rect 1327 2736 1493 2744
rect 1676 2744 1684 2776
rect 2067 2777 2093 2785
rect 2156 2776 2313 2784
rect 2156 2746 2164 2776
rect 2487 2776 2553 2784
rect 1607 2736 1684 2744
rect 1767 2733 1853 2741
rect 2047 2735 2113 2743
rect 2267 2736 2293 2744
rect 2356 2744 2364 2774
rect 2747 2776 2793 2784
rect 2816 2776 2853 2784
rect 2816 2746 2824 2776
rect 2967 2776 2993 2784
rect 3067 2779 3093 2787
rect 3247 2776 3284 2784
rect 3276 2764 3284 2776
rect 3327 2776 3353 2784
rect 3527 2776 3553 2784
rect 3607 2776 3693 2784
rect 3807 2777 3833 2785
rect 3887 2776 3933 2784
rect 3976 2764 3984 2793
rect 4147 2777 4233 2785
rect 4547 2776 4572 2784
rect 4607 2777 4653 2785
rect 4707 2777 4753 2785
rect 4827 2776 4953 2784
rect 5256 2784 5264 2796
rect 5527 2796 5713 2804
rect 5256 2776 5284 2784
rect 3276 2756 3304 2764
rect 3976 2760 4004 2764
rect 3976 2756 4007 2760
rect 2356 2736 2593 2744
rect 2647 2735 2713 2743
rect 3296 2746 3304 2756
rect 3993 2747 4007 2756
rect 4036 2747 4044 2773
rect 4536 2756 4644 2764
rect 3147 2736 3173 2744
rect 3407 2735 3493 2743
rect 3627 2735 3713 2743
rect 4107 2735 4293 2743
rect 4387 2735 4433 2743
rect 4536 2744 4544 2756
rect 4636 2746 4644 2756
rect 5076 2747 5084 2773
rect 5113 2764 5127 2773
rect 5113 2760 5184 2764
rect 5116 2756 5184 2760
rect 4487 2736 4544 2744
rect 4807 2735 4893 2743
rect 5176 2746 5184 2756
rect 5276 2746 5284 2776
rect 5316 2776 5473 2784
rect 5316 2747 5324 2776
rect 5567 2776 5773 2784
rect 5793 2784 5807 2793
rect 5896 2796 5933 2804
rect 5793 2780 5864 2784
rect 5796 2776 5864 2780
rect 607 2716 633 2724
rect 767 2716 793 2724
rect 867 2716 893 2724
rect 2207 2716 2333 2724
rect 2347 2716 2453 2724
rect 2847 2716 2873 2724
rect 3396 2724 3404 2732
rect 3347 2716 3404 2724
rect 3716 2724 3724 2732
rect 5856 2727 5864 2776
rect 5876 2744 5884 2773
rect 5896 2764 5904 2796
rect 5927 2776 5973 2784
rect 5996 2764 6004 2816
rect 5896 2756 5944 2764
rect 5936 2746 5944 2756
rect 5976 2756 6004 2764
rect 5876 2736 5893 2744
rect 3716 2716 3953 2724
rect 4567 2716 4773 2724
rect 4947 2716 5033 2724
rect 5427 2716 5493 2724
rect 5507 2716 5753 2724
rect 5856 2716 5873 2727
rect 5860 2713 5873 2716
rect 47 2696 153 2704
rect 267 2696 373 2704
rect 447 2696 613 2704
rect 1307 2696 1433 2704
rect 1447 2696 1613 2704
rect 1627 2696 1653 2704
rect 2567 2696 2773 2704
rect 3587 2696 3653 2704
rect 4067 2696 4273 2704
rect 4467 2696 4513 2704
rect 4607 2696 4833 2704
rect 5847 2696 5953 2704
rect 407 2676 833 2684
rect 2007 2676 2413 2684
rect 2467 2676 2493 2684
rect 2507 2676 3093 2684
rect 4127 2676 4233 2684
rect 4927 2676 5133 2684
rect 5427 2676 5693 2684
rect 5976 2684 5984 2756
rect 5927 2676 5984 2684
rect 847 2656 1133 2664
rect 1487 2656 1553 2664
rect 2407 2656 2433 2664
rect 2747 2656 2933 2664
rect 3407 2656 3853 2664
rect 3867 2656 4293 2664
rect 267 2636 1273 2644
rect 1287 2636 2973 2644
rect 4047 2636 4113 2644
rect 4687 2636 4753 2644
rect 4907 2636 5333 2644
rect 5507 2636 5933 2644
rect 1267 2616 1373 2624
rect 1867 2616 1953 2624
rect 2467 2616 2593 2624
rect 4547 2616 4573 2624
rect 4587 2616 4713 2624
rect 4727 2616 4992 2624
rect 5027 2616 5093 2624
rect 5516 2616 5793 2624
rect 607 2596 693 2604
rect 3427 2596 3673 2604
rect 4187 2596 4393 2604
rect 5516 2604 5524 2616
rect 5407 2596 5524 2604
rect 487 2576 573 2584
rect 3927 2576 4153 2584
rect 4787 2576 5113 2584
rect 5227 2576 5533 2584
rect 1647 2556 1733 2564
rect 1907 2556 2113 2564
rect 2287 2556 2673 2564
rect 3607 2556 3833 2564
rect 4227 2556 4713 2564
rect 4727 2556 5253 2564
rect 667 2536 1153 2544
rect 1607 2536 1753 2544
rect 1767 2536 2833 2544
rect 2553 2527 2567 2536
rect 3267 2536 3293 2544
rect 3307 2536 3413 2544
rect 3947 2536 4033 2544
rect 4347 2536 4913 2544
rect 5567 2536 5753 2544
rect 467 2516 533 2524
rect 856 2516 953 2524
rect 856 2507 864 2516
rect 4127 2516 4153 2524
rect 4167 2516 4333 2524
rect 4447 2516 4793 2524
rect 5567 2516 5613 2524
rect 47 2496 153 2504
rect 167 2496 753 2504
rect 767 2496 853 2504
rect 1787 2496 1993 2504
rect 2247 2496 2313 2504
rect 3467 2496 3533 2504
rect 3627 2496 3693 2504
rect 4027 2496 4213 2504
rect 4327 2496 4473 2504
rect 4967 2496 5053 2504
rect 5396 2496 5433 2504
rect 107 2479 133 2487
rect 507 2476 633 2484
rect 336 2427 344 2474
rect 496 2464 504 2474
rect 647 2476 813 2484
rect 827 2476 873 2484
rect 987 2476 1033 2484
rect 396 2456 504 2464
rect 396 2446 404 2456
rect 467 2433 553 2441
rect 567 2433 573 2441
rect 1156 2424 1164 2474
rect 1196 2447 1204 2474
rect 1247 2476 1333 2484
rect 1527 2476 1604 2484
rect 1596 2447 1604 2476
rect 1667 2477 1693 2485
rect 1747 2477 1813 2485
rect 2167 2476 2184 2484
rect 1196 2436 1213 2447
rect 1200 2433 1213 2436
rect 1287 2436 1373 2444
rect 1647 2435 1673 2443
rect 1827 2436 1873 2444
rect 2176 2444 2184 2476
rect 2296 2476 2493 2484
rect 2296 2446 2304 2476
rect 2807 2476 2853 2484
rect 2927 2479 3073 2487
rect 2176 2436 2253 2444
rect 2576 2444 2584 2473
rect 2487 2436 2584 2444
rect 2736 2427 2744 2476
rect 2796 2447 2804 2476
rect 3167 2476 3333 2484
rect 3387 2476 3433 2484
rect 3456 2476 3493 2484
rect 2796 2436 2813 2447
rect 2800 2433 2813 2436
rect 3047 2433 3113 2441
rect 3187 2436 3313 2444
rect 3456 2444 3464 2476
rect 3787 2476 3833 2484
rect 3847 2476 3993 2484
rect 4147 2476 4173 2484
rect 4747 2477 4813 2485
rect 4867 2477 4933 2485
rect 4987 2476 5033 2484
rect 5296 2476 5313 2484
rect 3536 2456 4093 2464
rect 3536 2446 3544 2456
rect 3816 2446 3824 2456
rect 3976 2446 3984 2456
rect 5296 2447 5304 2476
rect 3387 2436 3464 2444
rect 4167 2435 4213 2443
rect 4927 2435 4953 2443
rect 1067 2416 1233 2424
rect 1367 2416 1393 2424
rect 1407 2416 1473 2424
rect 2027 2416 2213 2424
rect 2316 2416 2373 2424
rect 213 2404 227 2413
rect 213 2400 253 2404
rect 216 2396 253 2400
rect 847 2396 933 2404
rect 1327 2396 1453 2404
rect 1607 2396 1713 2404
rect 2316 2404 2324 2416
rect 3567 2416 3613 2424
rect 3627 2416 3653 2424
rect 4307 2416 4733 2424
rect 4887 2416 4993 2424
rect 5356 2424 5364 2474
rect 5396 2447 5404 2496
rect 5616 2464 5624 2474
rect 5576 2460 5624 2464
rect 5573 2456 5624 2460
rect 5573 2447 5587 2456
rect 5107 2416 5364 2424
rect 2187 2396 2324 2404
rect 3087 2396 3353 2404
rect 3696 2396 3893 2404
rect 147 2376 353 2384
rect 447 2376 513 2384
rect 1027 2376 1133 2384
rect 1147 2376 1253 2384
rect 1727 2376 1793 2384
rect 1947 2376 2593 2384
rect 3696 2384 3704 2396
rect 4227 2396 4353 2404
rect 4367 2396 4453 2404
rect 5356 2404 5364 2416
rect 5387 2416 5553 2424
rect 5567 2416 5593 2424
rect 5656 2404 5664 2474
rect 5687 2476 5713 2484
rect 5787 2435 5973 2443
rect 5356 2396 5664 2404
rect 3447 2376 3704 2384
rect 4107 2376 4233 2384
rect 4667 2376 5093 2384
rect 5207 2376 5573 2384
rect 1547 2356 1613 2364
rect 2427 2356 2473 2364
rect 3207 2356 3593 2364
rect 3727 2356 4313 2364
rect 4367 2356 4593 2364
rect 4607 2356 5033 2364
rect 5187 2356 5773 2364
rect 1227 2336 1313 2344
rect 1767 2336 2053 2344
rect 2567 2336 2693 2344
rect 3107 2336 3173 2344
rect 3827 2336 4293 2344
rect 827 2316 893 2324
rect 1627 2316 1853 2324
rect 1867 2316 2253 2324
rect 2547 2316 2813 2324
rect 3327 2316 3393 2324
rect 3467 2316 3613 2324
rect 3927 2316 4013 2324
rect 4807 2316 4833 2324
rect 5007 2316 5073 2324
rect 5087 2316 5253 2324
rect 5267 2316 5473 2324
rect 5587 2316 5813 2324
rect 1267 2296 1333 2304
rect 1347 2296 1453 2304
rect 3287 2296 3433 2304
rect 4656 2296 4713 2304
rect 287 2276 513 2284
rect 987 2276 1073 2284
rect 1187 2276 1213 2284
rect 2447 2276 3013 2284
rect 3027 2276 3113 2284
rect 4087 2276 4153 2284
rect 4656 2284 4664 2296
rect 4787 2296 4853 2304
rect 5387 2296 5473 2304
rect 5647 2296 5733 2304
rect 5947 2296 5973 2304
rect 4527 2276 4664 2284
rect 4847 2276 4913 2284
rect 5167 2276 5324 2284
rect 707 2256 773 2264
rect 813 2264 827 2273
rect 813 2260 853 2264
rect 816 2256 853 2260
rect 876 2256 1013 2264
rect 396 2236 724 2244
rect -24 2204 -16 2224
rect 47 2216 153 2224
rect 396 2226 404 2236
rect 716 2226 724 2236
rect 876 2226 884 2256
rect 1107 2256 1153 2264
rect 1507 2257 1573 2265
rect 1687 2257 1753 2265
rect 1827 2256 2033 2264
rect 2107 2256 2193 2264
rect 2467 2256 2633 2264
rect 2647 2257 2693 2265
rect 2787 2257 2833 2265
rect 3367 2256 3444 2264
rect 3436 2244 3444 2256
rect 3467 2257 3553 2265
rect 3667 2256 3804 2264
rect 3436 2236 3553 2244
rect 367 2215 393 2223
rect 507 2215 633 2223
rect 787 2215 833 2223
rect 1567 2216 1693 2224
rect 1887 2213 1913 2221
rect 2007 2216 2033 2224
rect 2047 2215 2213 2223
rect 2347 2215 2553 2223
rect 2627 2216 2753 2224
rect 3007 2216 3113 2224
rect 3347 2215 3393 2223
rect 3587 2215 3633 2223
rect 3687 2215 3713 2223
rect 3796 2226 3804 2256
rect 4187 2256 4244 2264
rect 4236 2244 4244 2256
rect 4267 2256 4313 2264
rect 4687 2256 4793 2264
rect 4236 2236 4364 2244
rect 4127 2215 4193 2223
rect -24 2196 4 2204
rect -4 2184 4 2196
rect 267 2196 313 2204
rect 1007 2196 1093 2204
rect 1427 2196 1493 2204
rect 1507 2196 1533 2204
rect 1547 2196 1653 2204
rect 1727 2196 1773 2204
rect 3207 2196 3293 2204
rect 3576 2204 3584 2212
rect 4356 2207 4364 2236
rect 4476 2244 4484 2254
rect 4887 2256 4953 2264
rect 5016 2256 5133 2264
rect 4427 2236 4484 2244
rect 5016 2226 5024 2256
rect 5267 2256 5293 2264
rect 5316 2226 5324 2276
rect 5347 2276 5513 2284
rect 5527 2276 5593 2284
rect 5447 2256 5484 2264
rect 5356 2227 5364 2253
rect 4507 2215 4593 2223
rect 4707 2216 4773 2224
rect 4827 2215 4873 2223
rect 5087 2215 5113 2223
rect 5167 2216 5213 2224
rect 5227 2215 5273 2223
rect 5476 2207 5484 2256
rect 5647 2256 5693 2264
rect 5827 2256 5933 2264
rect 5573 2244 5587 2253
rect 5733 2244 5747 2253
rect 5573 2240 5604 2244
rect 5733 2240 5764 2244
rect 5576 2236 5604 2240
rect 5736 2236 5764 2240
rect 5596 2224 5604 2236
rect 5756 2226 5764 2236
rect 5507 2216 5613 2224
rect 5775 2207 5783 2254
rect 3487 2196 3584 2204
rect 3667 2196 3753 2204
rect 5807 2196 5853 2204
rect -4 2176 93 2184
rect 507 2176 533 2184
rect 1187 2176 1333 2184
rect 3607 2176 3833 2184
rect 3847 2176 4153 2184
rect 4167 2176 4373 2184
rect 4527 2176 4973 2184
rect 4987 2176 5193 2184
rect 447 2156 573 2164
rect 587 2156 613 2164
rect 627 2156 993 2164
rect 1007 2156 1413 2164
rect 1467 2156 1833 2164
rect 2847 2156 2973 2164
rect 2987 2156 3193 2164
rect 3807 2156 4333 2164
rect 4347 2156 4453 2164
rect 4667 2156 4973 2164
rect 4987 2156 5353 2164
rect 296 2136 513 2144
rect 296 2127 304 2136
rect 1047 2136 1213 2144
rect 1856 2136 2333 2144
rect 287 2116 304 2127
rect 287 2113 300 2116
rect 567 2116 833 2124
rect 1856 2124 1864 2136
rect 2687 2136 2913 2144
rect 2927 2136 3053 2144
rect 5107 2136 5333 2144
rect 1247 2116 1864 2124
rect 2707 2116 2793 2124
rect 2807 2116 2893 2124
rect 5467 2116 5793 2124
rect 507 2096 933 2104
rect 947 2096 2033 2104
rect 3927 2096 4133 2104
rect 4267 2096 4693 2104
rect 5207 2096 5413 2104
rect 1587 2076 1613 2084
rect 3907 2076 4173 2084
rect 4196 2076 4573 2084
rect 527 2056 673 2064
rect 747 2056 793 2064
rect 847 2056 1233 2064
rect 1287 2056 1313 2064
rect 1327 2056 1433 2064
rect 2487 2056 2533 2064
rect 4196 2064 4204 2076
rect 5747 2076 5873 2084
rect 3987 2056 4204 2064
rect 4367 2056 5013 2064
rect 27 2036 93 2044
rect 207 2036 233 2044
rect 247 2036 553 2044
rect 1627 2036 1953 2044
rect 5376 2036 5533 2044
rect 5376 2027 5384 2036
rect 5707 2036 5793 2044
rect 867 2016 953 2024
rect 2287 2016 2653 2024
rect 2967 2016 3133 2024
rect 4367 2016 4773 2024
rect 5067 2016 5173 2024
rect 5287 2016 5373 2024
rect 5567 2016 5653 2024
rect 5707 2016 5913 2024
rect 487 1996 573 2004
rect 1787 1996 1893 2004
rect 1967 1996 1993 2004
rect 2147 1996 2213 2004
rect 3107 1996 3153 2004
rect 3687 1996 3933 2004
rect 4927 1996 5033 2004
rect 5407 1996 5453 2004
rect 907 1976 1133 1984
rect 2547 1976 3013 1984
rect 3027 1976 3313 1984
rect 4707 1976 4733 1984
rect 4747 1976 5073 1984
rect 5247 1976 5353 1984
rect 5367 1976 5493 1984
rect 5687 1976 5713 1984
rect 5787 1976 5813 1984
rect 367 1956 533 1964
rect 547 1956 713 1964
rect 967 1959 1013 1967
rect 1847 1959 1873 1967
rect 327 1936 384 1944
rect 376 1926 384 1936
rect 1136 1927 1144 1956
rect 516 1920 593 1924
rect 513 1916 593 1920
rect 513 1907 527 1916
rect 607 1916 653 1924
rect 1127 1916 1144 1927
rect 1127 1913 1140 1916
rect 1527 1916 1593 1924
rect 1667 1916 1713 1924
rect 1976 1926 1984 1973
rect 2067 1957 2113 1965
rect 2087 1916 2133 1924
rect 2156 1924 2164 1954
rect 2156 1916 2253 1924
rect 2456 1924 2464 1956
rect 2587 1956 2693 1964
rect 2827 1956 3033 1964
rect 3196 1927 3204 1954
rect 2267 1916 2333 1924
rect 2456 1916 2633 1924
rect 3187 1916 3204 1927
rect 3187 1913 3200 1916
rect 3376 1924 3384 1956
rect 3627 1956 3704 1964
rect 3696 1927 3704 1956
rect 3787 1956 3833 1964
rect 3847 1956 3873 1964
rect 3947 1956 3984 1964
rect 3267 1916 3384 1924
rect 3747 1915 3793 1923
rect 3976 1924 3984 1956
rect 4067 1956 4204 1964
rect 4196 1944 4204 1956
rect 4227 1957 4273 1965
rect 4487 1956 4573 1964
rect 4627 1957 4673 1965
rect 4787 1956 4933 1964
rect 4976 1956 5053 1964
rect 4196 1940 4264 1944
rect 4196 1936 4267 1940
rect 4253 1927 4267 1936
rect 3976 1916 4033 1924
rect 4327 1915 4373 1923
rect 4547 1915 4593 1923
rect 4727 1915 4753 1923
rect 4767 1916 4913 1924
rect 4976 1924 4984 1956
rect 5387 1956 5433 1964
rect 5756 1956 5853 1964
rect 4967 1916 4984 1924
rect 5047 1915 5093 1923
rect 5267 1915 5453 1923
rect 5756 1926 5764 1956
rect 5507 1916 5593 1924
rect 307 1896 413 1904
rect 1947 1896 2013 1904
rect 2427 1896 2533 1904
rect 3127 1896 3493 1904
rect 3907 1896 4113 1904
rect 4427 1896 4573 1904
rect 5287 1896 5333 1904
rect 1107 1876 1233 1884
rect 1247 1876 1473 1884
rect 1647 1876 1733 1884
rect 3087 1876 3153 1884
rect 3167 1876 3213 1884
rect 3387 1876 3413 1884
rect 4387 1876 4673 1884
rect 4747 1876 4793 1884
rect 5307 1876 5593 1884
rect 5896 1884 5904 1993
rect 5936 1927 5944 1953
rect 5867 1876 5904 1884
rect 967 1856 993 1864
rect 1547 1860 1684 1864
rect 1547 1856 1687 1860
rect 1673 1847 1687 1856
rect 1907 1856 2293 1864
rect 2307 1856 2573 1864
rect 3447 1856 3633 1864
rect 4307 1856 4432 1864
rect 4467 1856 4693 1864
rect 5147 1856 5333 1864
rect 5636 1856 5733 1864
rect 5636 1847 5644 1856
rect 947 1836 1013 1844
rect 1147 1836 1513 1844
rect 1847 1836 1873 1844
rect 3847 1836 4113 1844
rect 4287 1836 4324 1844
rect 1136 1824 1144 1833
rect 956 1816 1144 1824
rect 427 1796 673 1804
rect 956 1804 964 1816
rect 1567 1816 1813 1824
rect 2867 1816 3213 1824
rect 4316 1824 4324 1836
rect 4467 1836 4513 1844
rect 4536 1836 4973 1844
rect 4536 1824 4544 1836
rect 5427 1836 5633 1844
rect 4007 1816 4304 1824
rect 4316 1816 4544 1824
rect 687 1796 964 1804
rect 1347 1796 1593 1804
rect 1607 1796 2793 1804
rect 3207 1796 3413 1804
rect 3727 1796 3873 1804
rect 4147 1796 4213 1804
rect 4296 1804 4304 1816
rect 4667 1816 5073 1824
rect 5187 1816 5393 1824
rect 5467 1816 5553 1824
rect 5567 1816 5704 1824
rect 5696 1807 5704 1816
rect 4296 1796 4753 1804
rect 5327 1796 5513 1804
rect 5696 1796 5713 1807
rect 5700 1793 5713 1796
rect 5887 1796 5973 1804
rect 1007 1776 1313 1784
rect 1727 1776 1973 1784
rect 2047 1776 2133 1784
rect 2147 1776 2333 1784
rect 2347 1776 2773 1784
rect 3047 1776 3653 1784
rect 3707 1776 3953 1784
rect 3967 1776 4373 1784
rect 4867 1776 4893 1784
rect 4967 1776 5013 1784
rect 5107 1776 5133 1784
rect 5287 1776 5324 1784
rect 2807 1756 2993 1764
rect 3287 1756 3313 1764
rect 4087 1756 4153 1764
rect 5167 1756 5213 1764
rect 336 1736 373 1744
rect 336 1707 344 1736
rect 507 1737 573 1745
rect 747 1737 813 1745
rect 867 1737 913 1745
rect 940 1744 953 1747
rect 936 1733 953 1744
rect 936 1724 944 1733
rect 876 1716 944 1724
rect 147 1696 193 1704
rect 207 1695 233 1703
rect 876 1706 884 1716
rect 767 1695 793 1703
rect 927 1696 1013 1704
rect 1056 1704 1064 1736
rect 1287 1736 1373 1744
rect 1416 1724 1424 1734
rect 1736 1736 1753 1744
rect 1307 1716 1424 1724
rect 1027 1696 1064 1704
rect 1187 1693 1273 1701
rect 1327 1695 1353 1703
rect 1407 1695 1453 1703
rect 1476 1704 1484 1733
rect 1736 1724 1744 1736
rect 2027 1737 2053 1745
rect 2187 1736 2213 1744
rect 2627 1736 2713 1744
rect 2727 1737 2773 1745
rect 2887 1737 2933 1745
rect 3027 1736 3064 1744
rect 3056 1724 3064 1736
rect 3347 1737 3373 1745
rect 3487 1736 3553 1744
rect 3727 1736 3773 1744
rect 3896 1736 4013 1744
rect 1627 1716 1744 1724
rect 2436 1716 3104 1724
rect 1476 1696 1493 1704
rect 1887 1693 1973 1701
rect 2107 1695 2133 1703
rect 2436 1704 2444 1716
rect 2747 1696 2853 1704
rect 2907 1695 2952 1703
rect 2976 1700 3013 1704
rect 2973 1696 3013 1700
rect 2973 1687 2987 1696
rect 3096 1704 3104 1716
rect 3176 1707 3184 1733
rect 3896 1706 3904 1736
rect 4027 1736 4184 1744
rect 4176 1706 4184 1736
rect 4487 1736 4533 1744
rect 4707 1736 4813 1744
rect 4867 1736 4913 1744
rect 4953 1724 4967 1733
rect 5016 1724 5024 1734
rect 4953 1720 5004 1724
rect 4956 1716 5004 1720
rect 5016 1720 5064 1724
rect 5016 1716 5067 1720
rect 3447 1695 3473 1703
rect 3967 1695 3993 1703
rect 4267 1696 4493 1704
rect 4567 1695 4593 1703
rect 4727 1696 4793 1704
rect 4807 1695 4893 1703
rect 4996 1704 5004 1716
rect 5053 1707 5067 1716
rect 5196 1707 5204 1733
rect 4996 1700 5024 1704
rect 4996 1696 5027 1700
rect 5013 1687 5027 1696
rect 5107 1695 5133 1703
rect 5256 1706 5264 1753
rect 5316 1687 5324 1776
rect 5347 1776 5533 1784
rect 5767 1776 5893 1784
rect 5413 1744 5427 1753
rect 5413 1740 5453 1744
rect 5416 1736 5453 1740
rect 5476 1724 5484 1753
rect 5556 1736 5633 1744
rect 5436 1716 5484 1724
rect 5387 1696 5413 1704
rect 5436 1687 5444 1716
rect 5516 1707 5524 1733
rect 5556 1707 5564 1736
rect 5656 1736 5733 1744
rect 5656 1707 5664 1736
rect 5807 1736 5973 1744
rect 307 1676 393 1684
rect 3407 1676 3573 1684
rect 4527 1676 4613 1684
rect 5716 1684 5724 1713
rect 5827 1695 5933 1703
rect 5716 1676 5793 1684
rect 547 1656 973 1664
rect 987 1656 1293 1664
rect 1307 1656 1333 1664
rect 1387 1656 1533 1664
rect 1547 1656 1693 1664
rect 2507 1656 2933 1664
rect 3007 1656 3093 1664
rect 3167 1656 3193 1664
rect 3547 1656 3693 1664
rect 4147 1656 4253 1664
rect 4616 1664 4624 1673
rect 5173 1664 5187 1673
rect 4616 1656 5293 1664
rect 3536 1644 3544 1653
rect 5587 1656 5653 1664
rect 5767 1656 5873 1664
rect 3327 1636 3544 1644
rect 4047 1636 4213 1644
rect 707 1616 933 1624
rect 947 1616 1273 1624
rect 1287 1616 1613 1624
rect 1827 1616 2893 1624
rect 5627 1616 5933 1624
rect 1647 1596 1713 1604
rect 2467 1596 2533 1604
rect 2687 1596 2973 1604
rect 3127 1596 3173 1604
rect 3467 1596 3733 1604
rect 3747 1596 3973 1604
rect 4487 1596 4813 1604
rect 5327 1596 5413 1604
rect 5487 1596 5893 1604
rect 367 1576 433 1584
rect 447 1576 1373 1584
rect 1807 1576 2373 1584
rect 2567 1576 2593 1584
rect 2976 1584 2984 1593
rect 2976 1576 3333 1584
rect 4947 1576 5113 1584
rect 5307 1576 5373 1584
rect 5607 1576 5693 1584
rect 2907 1556 3393 1564
rect 4447 1556 4593 1564
rect 4807 1556 4993 1564
rect 5007 1556 5473 1564
rect 167 1536 533 1544
rect 3047 1536 3133 1544
rect 4367 1536 4613 1544
rect 5047 1536 5313 1544
rect 5327 1536 5553 1544
rect 5787 1536 5873 1544
rect 107 1516 853 1524
rect 867 1516 1113 1524
rect 1127 1516 1253 1524
rect 1267 1516 1673 1524
rect 1687 1516 1833 1524
rect 1847 1516 1953 1524
rect 3667 1516 3893 1524
rect 4927 1516 4993 1524
rect 5387 1516 5593 1524
rect 1567 1496 1593 1504
rect 2967 1496 3253 1504
rect 3847 1496 4153 1504
rect 4167 1496 4313 1504
rect 5127 1496 5252 1504
rect 5287 1496 5353 1504
rect 5847 1496 5913 1504
rect 47 1476 93 1484
rect 467 1476 613 1484
rect 847 1476 1053 1484
rect 1627 1476 1853 1484
rect 3227 1476 3453 1484
rect 3687 1476 3813 1484
rect 5147 1476 5333 1484
rect 5687 1476 5753 1484
rect 347 1456 373 1464
rect 667 1456 833 1464
rect 2127 1456 2193 1464
rect 2207 1456 2233 1464
rect 2907 1456 2993 1464
rect 3007 1456 3413 1464
rect 3427 1456 3733 1464
rect 5056 1456 5113 1464
rect 96 1407 104 1436
rect 507 1437 532 1445
rect 567 1436 773 1444
rect 887 1436 933 1444
rect 1107 1437 1133 1445
rect 1156 1436 1213 1444
rect 1156 1424 1164 1436
rect 1427 1436 1533 1444
rect 1547 1436 1753 1444
rect 1807 1436 1833 1444
rect 1887 1437 1913 1445
rect 1967 1437 2012 1445
rect 2047 1437 2073 1445
rect 2096 1436 2253 1444
rect 1116 1416 1164 1424
rect 1196 1416 1273 1424
rect 96 1396 113 1407
rect 100 1393 113 1396
rect 1116 1406 1124 1416
rect 1196 1406 1204 1416
rect 2096 1424 2104 1436
rect 2347 1436 2373 1444
rect 2447 1436 2493 1444
rect 2567 1436 2653 1444
rect 2727 1436 2793 1444
rect 3207 1436 3313 1444
rect 1996 1416 2104 1424
rect 227 1393 293 1401
rect 407 1395 553 1403
rect 727 1395 753 1403
rect 807 1395 1033 1403
rect 1487 1393 1533 1401
rect 1787 1396 1873 1404
rect 1996 1404 2004 1416
rect 1987 1396 2004 1404
rect 2027 1396 2093 1404
rect 2187 1395 2233 1403
rect 2287 1396 2393 1404
rect 2407 1395 2432 1403
rect 2467 1396 2533 1404
rect 2836 1404 2844 1434
rect 3807 1436 3853 1444
rect 3947 1437 4013 1445
rect 4227 1436 4273 1444
rect 2707 1396 2844 1404
rect 1227 1376 1393 1384
rect 2176 1384 2184 1392
rect 1887 1376 2184 1384
rect 2567 1376 2593 1384
rect 2716 1384 2724 1396
rect 3087 1396 3173 1404
rect 3247 1395 3293 1403
rect 3387 1396 3553 1404
rect 3567 1393 3792 1401
rect 3827 1396 4033 1404
rect 4056 1404 4064 1434
rect 4387 1436 4433 1444
rect 4556 1424 4564 1434
rect 5056 1444 5064 1456
rect 5547 1456 5573 1464
rect 5667 1456 5724 1464
rect 4647 1436 5064 1444
rect 4556 1416 4973 1424
rect 4056 1396 4093 1404
rect 5076 1387 5084 1433
rect 5133 1424 5147 1433
rect 5096 1420 5147 1424
rect 5156 1436 5213 1444
rect 5096 1416 5144 1420
rect 5096 1406 5104 1416
rect 5156 1407 5164 1436
rect 5236 1436 5313 1444
rect 5147 1396 5164 1407
rect 5236 1406 5244 1436
rect 5516 1407 5524 1433
rect 5696 1407 5704 1433
rect 5716 1424 5724 1456
rect 5747 1456 5813 1464
rect 5716 1416 5744 1424
rect 5147 1393 5160 1396
rect 5587 1395 5633 1403
rect 5736 1404 5744 1416
rect 5736 1396 5813 1404
rect 2716 1376 3213 1384
rect 3447 1376 3473 1384
rect 4127 1376 4193 1384
rect 5067 1376 5084 1387
rect 5856 1384 5864 1453
rect 5856 1376 5893 1384
rect 5067 1373 5080 1376
rect 247 1356 353 1364
rect 467 1356 533 1364
rect 547 1356 673 1364
rect 687 1356 913 1364
rect 967 1356 1013 1364
rect 1027 1356 1153 1364
rect 1327 1356 3093 1364
rect 3287 1356 3373 1364
rect 3887 1356 3933 1364
rect 4227 1356 4392 1364
rect 4427 1356 4893 1364
rect 5247 1356 5573 1364
rect 547 1336 653 1344
rect 1207 1336 1233 1344
rect 1867 1336 1933 1344
rect 2527 1336 2773 1344
rect 2787 1336 2813 1344
rect 3267 1336 3333 1344
rect 3407 1336 3433 1344
rect 4287 1336 4533 1344
rect 4547 1336 4673 1344
rect 4687 1336 4813 1344
rect 5007 1336 5133 1344
rect 5607 1336 5713 1344
rect 67 1316 133 1324
rect 287 1316 353 1324
rect 507 1316 633 1324
rect 847 1316 1113 1324
rect 3187 1316 3493 1324
rect 3507 1316 3593 1324
rect 4087 1316 4213 1324
rect 4307 1316 4692 1324
rect 4727 1316 4973 1324
rect 207 1296 233 1304
rect 667 1296 953 1304
rect 1167 1296 1433 1304
rect 2107 1296 2133 1304
rect 2147 1296 2333 1304
rect 2347 1296 2413 1304
rect 3787 1296 3853 1304
rect 4107 1296 4233 1304
rect 4447 1296 4553 1304
rect 4787 1296 5333 1304
rect 5347 1296 5393 1304
rect 5507 1296 5673 1304
rect 5687 1296 5713 1304
rect 167 1276 313 1284
rect 2067 1276 2393 1284
rect 2447 1276 2733 1284
rect 2827 1276 3013 1284
rect 3147 1276 3573 1284
rect 3647 1276 3833 1284
rect 3847 1276 4073 1284
rect 4267 1276 5313 1284
rect 1427 1256 1733 1264
rect 2967 1256 3013 1264
rect 3027 1256 3653 1264
rect 4147 1256 4353 1264
rect 4647 1256 4773 1264
rect 5547 1256 5613 1264
rect 5827 1256 5913 1264
rect 2207 1236 2353 1244
rect 2687 1236 2753 1244
rect 2847 1236 2873 1244
rect 2887 1236 3453 1244
rect 3987 1236 4093 1244
rect 4107 1236 4333 1244
rect 4407 1236 4513 1244
rect 4847 1236 4873 1244
rect 4947 1236 5064 1244
rect 216 1216 253 1224
rect 216 1204 224 1216
rect 347 1217 413 1225
rect 436 1216 573 1224
rect 293 1204 307 1213
rect 96 1196 224 1204
rect 256 1200 307 1204
rect 256 1196 304 1200
rect 96 1186 104 1196
rect 256 1184 264 1196
rect 436 1186 444 1216
rect 840 1224 853 1227
rect 247 1176 264 1184
rect 367 1175 393 1183
rect 656 1184 664 1216
rect 836 1213 853 1224
rect 907 1216 953 1224
rect 1213 1224 1227 1233
rect 1213 1220 1253 1224
rect 1216 1216 1253 1220
rect 1456 1216 1473 1224
rect 1596 1216 1793 1224
rect 836 1184 844 1213
rect 1016 1196 1224 1204
rect 1016 1186 1024 1196
rect 567 1176 664 1184
rect 947 1175 1013 1183
rect 1107 1175 1173 1183
rect 1216 1184 1224 1196
rect 1216 1176 1233 1184
rect 1456 1184 1464 1216
rect 1596 1184 1604 1216
rect 1836 1204 1844 1214
rect 1907 1216 1933 1224
rect 2147 1217 2173 1225
rect 1816 1196 1844 1204
rect 1447 1176 1464 1184
rect 1667 1173 1693 1181
rect 1747 1175 1773 1183
rect 1816 1167 1824 1196
rect 1976 1184 1984 1214
rect 2407 1216 2453 1224
rect 2627 1217 2653 1225
rect 3400 1224 3413 1227
rect 1976 1176 2113 1184
rect 2367 1175 2433 1183
rect 2487 1175 2513 1183
rect 2767 1175 2833 1183
rect 2916 1184 2924 1214
rect 3396 1213 3413 1224
rect 3547 1216 3913 1224
rect 5056 1228 5064 1236
rect 5287 1236 5353 1244
rect 5376 1236 5413 1244
rect 2916 1176 3033 1184
rect 3107 1176 3153 1184
rect 3396 1184 3404 1213
rect 3676 1186 3684 1216
rect 3916 1204 3924 1216
rect 4007 1217 4053 1225
rect 4207 1216 4293 1224
rect 4487 1216 4584 1224
rect 3916 1196 4064 1204
rect 3467 1176 3513 1184
rect 3607 1175 3633 1183
rect 3867 1175 4033 1183
rect 4056 1184 4064 1196
rect 4576 1186 4584 1216
rect 5067 1217 5093 1225
rect 5116 1216 5273 1224
rect 5116 1204 5124 1216
rect 4976 1196 5124 1204
rect 4056 1176 4173 1184
rect 4387 1175 4433 1183
rect 4927 1176 4953 1184
rect 4976 1184 4984 1196
rect 5376 1187 5384 1236
rect 5707 1236 5864 1244
rect 5513 1224 5527 1233
rect 5513 1220 5564 1224
rect 5516 1216 5564 1220
rect 5436 1187 5444 1213
rect 5493 1204 5507 1213
rect 5493 1200 5524 1204
rect 5496 1196 5524 1200
rect 4967 1176 4984 1184
rect 5176 1176 5213 1184
rect 287 1156 313 1164
rect 507 1156 533 1164
rect 1287 1156 1313 1164
rect 1807 1156 1824 1167
rect 1807 1153 1820 1156
rect 1887 1156 1993 1164
rect 3127 1156 3173 1164
rect 3407 1156 3733 1164
rect 4367 1156 4493 1164
rect 607 1136 893 1144
rect 1007 1136 1833 1144
rect 2047 1136 2113 1144
rect 2187 1136 2593 1144
rect 2667 1136 2893 1144
rect 3807 1136 4133 1144
rect 5176 1144 5184 1176
rect 5436 1176 5453 1187
rect 5440 1173 5453 1176
rect 5516 1186 5524 1196
rect 5556 1186 5564 1216
rect 5587 1216 5613 1224
rect 5687 1216 5704 1224
rect 5567 1176 5653 1184
rect 5696 1167 5704 1216
rect 5776 1187 5784 1213
rect 5856 1187 5864 1236
rect 5207 1156 5413 1164
rect 5687 1156 5704 1167
rect 5687 1153 5700 1156
rect 4787 1136 5184 1144
rect 5467 1136 5573 1144
rect 5647 1136 5833 1144
rect 1147 1116 1433 1124
rect 4547 1116 4613 1124
rect 5067 1116 5453 1124
rect 5827 1116 5873 1124
rect 1807 1096 2873 1104
rect 2887 1096 3413 1104
rect 5007 1096 5493 1104
rect 1827 1076 2293 1084
rect 2547 1076 2793 1084
rect 4007 1076 4233 1084
rect 4647 1076 5013 1084
rect 5707 1076 5913 1084
rect 1207 1056 2453 1064
rect 2567 1056 2613 1064
rect 2727 1056 2953 1064
rect 3367 1056 3433 1064
rect 5147 1056 5513 1064
rect 1047 1036 1833 1044
rect 3167 1036 3393 1044
rect 3847 1036 4213 1044
rect 4467 1036 4893 1044
rect 987 1016 2093 1024
rect 3527 1016 3573 1024
rect 5207 1016 5253 1024
rect 5267 1016 5713 1024
rect 1687 996 2004 1004
rect 1996 984 2004 996
rect 2467 996 2924 1004
rect 2916 987 2924 996
rect 5087 996 5153 1004
rect 5307 996 5533 1004
rect 1996 976 2273 984
rect 2927 976 3093 984
rect 3347 976 3433 984
rect 5187 976 5233 984
rect 5607 976 5653 984
rect 5867 976 5913 984
rect 67 956 233 964
rect 327 956 493 964
rect 507 956 753 964
rect 1467 956 1733 964
rect 1987 956 2413 964
rect 4607 956 4713 964
rect 5287 956 5313 964
rect 5467 956 5573 964
rect 616 936 713 944
rect 67 916 93 924
rect 136 867 144 933
rect 616 927 624 936
rect 727 936 973 944
rect 2967 936 3053 944
rect 4356 936 4653 944
rect 387 916 413 924
rect 687 916 853 924
rect 1027 916 1073 924
rect 1087 916 1133 924
rect 1247 917 1273 925
rect 1516 904 1524 916
rect 1807 916 1893 924
rect 1636 904 1644 914
rect 2056 916 2153 924
rect 1516 900 1544 904
rect 1596 900 1644 904
rect 1516 896 1547 900
rect 1533 887 1547 896
rect 167 876 193 884
rect 527 876 573 884
rect 787 876 833 884
rect 887 876 993 884
rect 1167 876 1233 884
rect 1307 876 1333 884
rect 1593 896 1644 900
rect 1593 887 1607 896
rect 1667 875 1733 883
rect 1936 884 1944 914
rect 1827 876 1944 884
rect 2056 884 2064 916
rect 1967 876 2064 884
rect 2216 887 2224 916
rect 2307 916 2333 924
rect 2347 916 2453 924
rect 2507 917 2533 925
rect 2727 916 2753 924
rect 2216 876 2233 887
rect 2220 873 2233 876
rect 2287 876 2473 884
rect 3016 884 3024 914
rect 3107 924 3120 927
rect 3107 913 3124 924
rect 3207 919 3233 927
rect 3307 919 3333 927
rect 3116 884 3124 913
rect 2907 876 3024 884
rect 3187 876 3373 884
rect 3416 886 3424 933
rect 3487 916 3593 924
rect 3667 917 3693 925
rect 3707 916 3753 924
rect 3807 917 3833 925
rect 3887 916 3933 924
rect 4307 916 4333 924
rect 3867 875 3913 883
rect 4056 884 4064 914
rect 4296 904 4304 916
rect 4356 924 4364 936
rect 4787 936 4993 944
rect 5127 936 5164 944
rect 4347 916 4364 924
rect 4387 916 4413 924
rect 4427 916 4764 924
rect 4207 896 4304 904
rect 4056 876 4093 884
rect 4756 886 4764 916
rect 4776 867 4784 914
rect 4816 884 4824 914
rect 4816 876 4853 884
rect 347 856 373 864
rect 627 856 653 864
rect 1627 856 1693 864
rect 1707 856 1913 864
rect 3487 856 3633 864
rect 3647 856 3773 864
rect 3787 856 3873 864
rect 4087 856 4113 864
rect 4247 856 4353 864
rect 4547 856 4593 864
rect 4916 866 4924 913
rect 4956 884 4964 914
rect 5156 886 5164 936
rect 5276 944 5284 953
rect 5187 936 5284 944
rect 5507 936 5553 944
rect 5636 936 5773 944
rect 5207 916 5264 924
rect 5256 886 5264 916
rect 5347 916 5393 924
rect 5476 887 5484 913
rect 4956 876 5113 884
rect 5527 876 5573 884
rect 4947 856 5453 864
rect 5636 866 5644 936
rect 5687 875 5733 883
rect 5816 864 5824 914
rect 5896 867 5904 913
rect 5816 856 5852 864
rect 5887 856 5904 867
rect 5887 853 5900 856
rect 1187 836 1553 844
rect 1907 836 1993 844
rect 2387 836 2673 844
rect 3047 836 3193 844
rect 3507 836 3613 844
rect 4727 836 4793 844
rect 5067 836 5253 844
rect 5387 836 5593 844
rect 667 816 953 824
rect 2967 816 3173 824
rect 4707 816 4832 824
rect 4867 816 4973 824
rect 5627 816 5793 824
rect 5847 816 5973 824
rect 1167 796 1593 804
rect 1887 796 2013 804
rect 2067 796 2093 804
rect 2107 796 2273 804
rect 3267 796 3333 804
rect 3347 796 4193 804
rect 5047 796 5113 804
rect 5227 796 5573 804
rect 1927 776 2113 784
rect 2127 776 2293 784
rect 2727 776 2773 784
rect 4227 776 4373 784
rect 4487 776 4553 784
rect 5387 776 5613 784
rect 5667 776 5833 784
rect 587 756 653 764
rect 667 756 713 764
rect 1867 756 3273 764
rect 3327 756 3913 764
rect 3987 756 4673 764
rect 5107 756 5313 764
rect 5367 756 5893 764
rect 307 736 513 744
rect 967 736 1053 744
rect 2227 736 2313 744
rect 2627 736 2853 744
rect 3067 736 3293 744
rect 3307 736 3933 744
rect 4347 736 4613 744
rect 5096 744 5104 753
rect 5036 736 5104 744
rect 2487 716 2813 724
rect 2827 716 2893 724
rect 3887 724 3900 727
rect 3887 713 3904 724
rect 467 696 504 704
rect 227 656 313 664
rect 336 664 344 694
rect 496 667 504 696
rect 707 697 772 705
rect 807 697 833 705
rect 1267 696 1433 704
rect 1447 696 1473 704
rect 1567 697 1753 705
rect 1807 696 1844 704
rect 336 656 413 664
rect 616 664 624 694
rect 616 656 713 664
rect 787 656 853 664
rect 876 664 884 694
rect 1116 684 1124 694
rect 1116 676 1304 684
rect 876 656 1273 664
rect 1296 664 1304 676
rect 1836 667 1844 696
rect 2116 696 2213 704
rect 1296 656 1413 664
rect 1427 656 1553 664
rect 1707 655 1773 663
rect 1947 655 2053 663
rect 2116 664 2124 696
rect 2207 656 2233 664
rect 2296 666 2304 713
rect 2367 697 2393 705
rect 2447 697 2473 705
rect 2527 696 2553 704
rect 2647 696 2813 704
rect 2967 697 3013 705
rect 3227 696 3433 704
rect 3447 696 3553 704
rect 3607 696 3693 704
rect 2507 656 2633 664
rect 2747 653 2773 661
rect 2827 655 2873 663
rect 3047 656 3093 664
rect 3216 664 3224 694
rect 3896 704 3904 713
rect 4016 716 4193 724
rect 3896 696 3993 704
rect 3856 667 3864 693
rect 3216 656 3313 664
rect 3627 656 3733 664
rect 3747 656 3832 664
rect 3907 656 3933 664
rect 4016 666 4024 716
rect 4127 697 4153 705
rect 4347 696 4373 704
rect 4356 667 4364 696
rect 4487 704 4500 707
rect 4487 693 4504 704
rect 4727 696 4833 704
rect 5036 704 5044 736
rect 5487 736 5613 744
rect 5147 716 5213 724
rect 5727 716 5773 724
rect 5816 716 5913 724
rect 4956 700 5044 704
rect 4953 696 5044 700
rect 4067 656 4113 664
rect 4496 664 4504 693
rect 4953 686 4967 696
rect 5227 696 5324 704
rect 5316 666 5324 696
rect 5387 696 5493 704
rect 5536 667 5544 693
rect 5596 667 5604 693
rect 5816 667 5824 716
rect 4567 653 4613 661
rect 4867 655 4913 663
rect 5127 655 5153 663
rect 5467 656 5513 664
rect 5536 656 5553 667
rect 5540 653 5553 656
rect 5687 656 5773 664
rect 5867 656 5913 664
rect 527 636 593 644
rect 807 636 1133 644
rect 1827 636 1853 644
rect 2627 636 2673 644
rect 2807 636 2913 644
rect 5587 636 5684 644
rect 796 624 804 633
rect 427 616 804 624
rect 1327 616 1584 624
rect 47 596 113 604
rect 1576 604 1584 616
rect 1607 616 1793 624
rect 2127 616 2413 624
rect 3167 616 3513 624
rect 3527 616 4113 624
rect 4127 616 4493 624
rect 4507 616 4733 624
rect 4747 616 4773 624
rect 4787 616 5273 624
rect 5347 616 5493 624
rect 5676 624 5684 636
rect 5676 616 5773 624
rect 1576 596 1733 604
rect 3207 596 3573 604
rect 3807 596 4173 604
rect 4827 596 4933 604
rect 4947 596 4973 604
rect 5327 596 5693 604
rect 447 576 773 584
rect 1447 576 2953 584
rect 4627 576 4693 584
rect 4707 576 5233 584
rect 5567 576 5673 584
rect 547 556 613 564
rect 927 556 1153 564
rect 2407 556 2693 564
rect 2987 556 3493 564
rect 407 536 773 544
rect 787 536 1113 544
rect 1127 536 1453 544
rect 1467 536 1533 544
rect 1547 536 1673 544
rect 1687 536 1813 544
rect 1827 536 1993 544
rect 2007 536 2193 544
rect 4807 536 5013 544
rect 1027 516 1073 524
rect 4607 516 5664 524
rect 647 496 1433 504
rect 4907 496 5633 504
rect 5656 504 5664 516
rect 5656 496 5873 504
rect 127 476 353 484
rect 367 476 473 484
rect 1547 476 2433 484
rect 3047 476 3353 484
rect 3367 476 3433 484
rect 1007 456 1033 464
rect 1707 456 2853 464
rect 2967 456 3153 464
rect 3167 456 3373 464
rect 4887 456 4993 464
rect 5007 456 5073 464
rect 5587 456 5973 464
rect 387 436 473 444
rect 1167 436 1533 444
rect 2087 436 2413 444
rect 3987 436 4293 444
rect 4656 436 4753 444
rect 376 416 413 424
rect 187 396 233 404
rect 376 366 384 416
rect 587 416 653 424
rect 1047 424 1060 427
rect 1047 413 1064 424
rect 2607 416 2773 424
rect 2787 416 3133 424
rect 3147 416 3253 424
rect 3807 416 3853 424
rect 3867 416 3913 424
rect 4247 416 4313 424
rect 4656 424 4664 436
rect 5527 436 5593 444
rect 5607 436 5733 444
rect 4636 416 4664 424
rect 467 397 533 405
rect 396 364 404 394
rect 656 396 673 404
rect 616 367 624 393
rect 656 367 664 396
rect 727 397 753 405
rect 867 397 973 405
rect 396 356 433 364
rect 816 364 824 394
rect 1016 367 1024 393
rect 1056 367 1064 413
rect 1227 396 1373 404
rect 707 356 824 364
rect 1167 355 1233 363
rect 1247 356 1393 364
rect 1416 364 1424 394
rect 1416 356 1493 364
rect 1516 347 1524 394
rect 1556 367 1564 394
rect 1687 396 1713 404
rect 1727 396 1913 404
rect 1556 356 1573 367
rect 1560 353 1573 356
rect 2036 364 2044 394
rect 2036 356 2173 364
rect 567 336 633 344
rect 876 336 913 344
rect 876 327 884 336
rect 2067 336 2113 344
rect 2196 344 2204 394
rect 2236 364 2244 394
rect 2407 396 2473 404
rect 2527 396 2753 404
rect 2807 397 2833 405
rect 2927 396 2973 404
rect 2287 376 2344 384
rect 2236 356 2313 364
rect 2336 364 2344 376
rect 2336 356 2353 364
rect 2427 356 2493 364
rect 2756 364 2764 394
rect 3347 396 3613 404
rect 3776 396 3813 404
rect 3076 367 3084 394
rect 2667 356 2764 364
rect 2987 355 3013 363
rect 3076 356 3093 367
rect 3080 353 3093 356
rect 3776 366 3784 396
rect 3867 396 4053 404
rect 4147 397 4173 405
rect 4467 397 4533 405
rect 4036 376 4233 384
rect 4036 366 4044 376
rect 3167 355 3213 363
rect 3367 355 3453 363
rect 3647 356 3733 364
rect 3867 355 3893 363
rect 3947 355 3973 363
rect 4087 356 4133 364
rect 4207 356 4273 364
rect 4327 355 4353 363
rect 4636 366 4644 416
rect 4927 416 4953 424
rect 5207 416 5333 424
rect 5407 416 5453 424
rect 5627 416 5704 424
rect 5696 408 5704 416
rect 5847 416 5913 424
rect 4707 396 4813 404
rect 4827 397 4853 405
rect 4547 356 4593 364
rect 4687 356 4733 364
rect 4747 355 4793 363
rect 4807 356 4873 364
rect 4896 364 4904 394
rect 4896 356 4933 364
rect 5036 364 5044 394
rect 5107 396 5324 404
rect 5036 356 5133 364
rect 5316 366 5324 396
rect 5427 396 5633 404
rect 5707 396 5793 404
rect 5987 396 6024 404
rect 5896 367 5904 393
rect 5187 355 5233 363
rect 5667 355 5713 363
rect 5827 355 5853 363
rect 2196 336 2273 344
rect 2367 336 2573 344
rect 2707 336 2773 344
rect 4827 336 5053 344
rect 5067 336 5373 344
rect 227 316 873 324
rect 1007 316 1893 324
rect 1907 316 2693 324
rect 2707 316 2833 324
rect 3027 316 3093 324
rect 5307 316 5433 324
rect 5447 316 5493 324
rect 5827 316 5953 324
rect 327 296 433 304
rect 547 296 613 304
rect 1507 296 1673 304
rect 4487 296 4613 304
rect 4927 296 5253 304
rect 5687 296 5893 304
rect 407 276 473 284
rect 967 276 1033 284
rect 1327 276 1533 284
rect 1607 276 1633 284
rect 2667 276 3313 284
rect 5287 276 5553 284
rect 107 256 313 264
rect 1787 256 1892 264
rect 1927 256 2273 264
rect 2607 256 2633 264
rect 2867 256 4433 264
rect 4907 256 4973 264
rect 987 236 1693 244
rect 2487 236 2533 244
rect 2547 236 2653 244
rect 2667 236 2733 244
rect 5647 236 5853 244
rect 167 216 213 224
rect 1867 216 2033 224
rect 2287 216 2393 224
rect 2807 216 2873 224
rect 3067 216 3173 224
rect 3467 216 3513 224
rect 3607 216 3693 224
rect 3867 216 4553 224
rect 5407 216 5433 224
rect 5527 216 5573 224
rect 1207 196 1253 204
rect 1936 196 1993 204
rect 96 146 104 193
rect 127 176 213 184
rect 267 176 573 184
rect 587 179 653 187
rect 1007 176 1113 184
rect 1196 176 1253 184
rect 256 164 264 173
rect 236 156 264 164
rect 696 156 833 164
rect 236 146 244 156
rect 167 135 193 143
rect 696 144 704 156
rect 1196 146 1204 176
rect 1727 176 1793 184
rect 1836 164 1844 193
rect 1876 176 1913 184
rect 1836 156 1864 164
rect 907 136 1013 144
rect 1127 135 1153 143
rect 1347 133 1373 141
rect 1447 133 1473 141
rect 1607 136 1633 144
rect 1647 136 1693 144
rect 1747 135 1773 143
rect 1856 124 1864 156
rect 1876 146 1884 176
rect 1936 144 1944 196
rect 2907 196 2933 204
rect 5127 196 5493 204
rect 5727 196 5793 204
rect 2127 176 2213 184
rect 2327 177 2373 185
rect 2387 176 2413 184
rect 2636 176 2733 184
rect 2007 136 2033 144
rect 2367 135 2473 143
rect 2636 144 2644 176
rect 2847 184 2860 187
rect 2847 173 2864 184
rect 2967 179 3093 187
rect 3167 176 3284 184
rect 2856 146 2864 173
rect 2547 136 2644 144
rect 2667 135 2713 143
rect 2767 135 2793 143
rect 2907 136 2953 144
rect 2967 136 2993 144
rect 3276 144 3284 176
rect 3356 176 3373 184
rect 3356 147 3364 176
rect 3427 176 3493 184
rect 3547 176 3633 184
rect 3187 133 3213 141
rect 3496 144 3504 174
rect 3887 179 3933 187
rect 4096 176 4113 184
rect 3756 156 3853 164
rect 3407 136 3504 144
rect 3567 135 3593 143
rect 3756 144 3764 156
rect 4096 146 4104 176
rect 4127 177 4173 185
rect 4227 177 4353 185
rect 4596 176 4753 184
rect 4476 156 4553 164
rect 4147 135 4193 143
rect 4476 144 4484 156
rect 4596 146 4604 176
rect 4807 176 4893 184
rect 5007 177 5073 185
rect 5307 176 5373 184
rect 5356 156 5433 164
rect 4367 136 4413 144
rect 4647 135 4673 143
rect 4927 136 4973 144
rect 4987 136 5033 144
rect 5107 136 5133 144
rect 5356 146 5364 156
rect 5147 136 5193 144
rect 5267 135 5293 143
rect 5407 136 5513 144
rect 5587 135 5613 143
rect 5667 135 5713 143
rect 5807 135 5913 143
rect 1856 116 1893 124
rect 3447 116 3513 124
rect 3527 116 3673 124
rect 4747 116 4853 124
rect 3436 104 3444 113
rect 3047 96 3444 104
rect 3727 96 3873 104
rect 3887 96 4053 104
rect 4167 96 4233 104
rect 4787 96 4953 104
rect 3647 76 3693 84
rect 3747 76 3813 84
rect 1527 36 1553 44
rect 1567 36 3033 44
rect 4007 36 5833 44
rect 67 16 93 24
rect 3367 16 3393 24
rect 3467 16 3493 24
use NOR2X1  _723_
timestamp 0
transform 1 0 1190 0 1 1310
box -6 -8 86 268
use INVX2  _724_
timestamp 0
transform -1 0 710 0 -1 1830
box -6 -8 66 268
use NOR2X1  _725_
timestamp 0
transform -1 0 1730 0 -1 1830
box -6 -8 86 268
use OAI21X1  _726_
timestamp 0
transform -1 0 1450 0 1 1310
box -6 -8 106 268
use INVX2  _727_
timestamp 0
transform 1 0 1990 0 1 2350
box -6 -8 66 268
use NOR2X1  _728_
timestamp 0
transform -1 0 2130 0 1 3390
box -6 -8 86 268
use AOI22X1  _729_
timestamp 0
transform -1 0 890 0 -1 1830
box -6 -8 126 268
use OAI21X1  _730_
timestamp 0
transform -1 0 1130 0 1 1310
box -6 -8 106 268
use INVX1  _731_
timestamp 0
transform 1 0 470 0 1 1310
box -6 -8 66 268
use INVX1  _732_
timestamp 0
transform -1 0 3190 0 -1 1310
box -6 -8 66 268
use NAND2X1  _733_
timestamp 0
transform 1 0 1230 0 -1 1310
box -6 -8 86 268
use OAI21X1  _734_
timestamp 0
transform -1 0 1170 0 -1 1310
box -6 -8 106 268
use AOI22X1  _735_
timestamp 0
transform -1 0 630 0 1 1830
box -6 -8 126 268
use OAI21X1  _736_
timestamp 0
transform -1 0 690 0 1 1310
box -6 -8 106 268
use INVX1  _737_
timestamp 0
transform -1 0 1970 0 -1 790
box -6 -8 66 268
use NAND2X1  _738_
timestamp 0
transform 1 0 930 0 -1 1310
box -6 -8 86 268
use OAI21X1  _739_
timestamp 0
transform 1 0 530 0 -1 1310
box -6 -8 106 268
use AOI22X1  _740_
timestamp 0
transform -1 0 590 0 -1 2350
box -6 -8 126 268
use OAI21X1  _741_
timestamp 0
transform -1 0 470 0 -1 1310
box -6 -8 106 268
use NOR2X1  _742_
timestamp 0
transform 1 0 750 0 1 1310
box -6 -8 86 268
use OAI21X1  _743_
timestamp 0
transform -1 0 430 0 -1 1830
box -6 -8 106 268
use AOI22X1  _744_
timestamp 0
transform -1 0 450 0 1 1830
box -6 -8 126 268
use OAI21X1  _745_
timestamp 0
transform -1 0 410 0 1 1310
box -6 -8 106 268
use INVX2  _746_
timestamp 0
transform 1 0 3530 0 -1 3390
box -6 -8 66 268
use NAND2X1  _747_
timestamp 0
transform -1 0 3310 0 1 3390
box -6 -8 86 268
use OAI21X1  _748_
timestamp 0
transform 1 0 3370 0 -1 3390
box -6 -8 106 268
use INVX1  _749_
timestamp 0
transform 1 0 3930 0 -1 3910
box -6 -8 66 268
use NAND2X1  _750_
timestamp 0
transform -1 0 4030 0 1 3910
box -6 -8 86 268
use OAI21X1  _751_
timestamp 0
transform -1 0 4190 0 1 3910
box -6 -8 106 268
use INVX2  _752_
timestamp 0
transform 1 0 4050 0 -1 3910
box -6 -8 66 268
use NAND2X1  _753_
timestamp 0
transform -1 0 4330 0 1 3910
box -6 -8 86 268
use OAI21X1  _754_
timestamp 0
transform 1 0 4390 0 1 3910
box -6 -8 106 268
use INVX2  _755_
timestamp 0
transform -1 0 3750 0 1 2870
box -6 -8 66 268
use NAND2X1  _756_
timestamp 0
transform -1 0 4450 0 1 3390
box -6 -8 86 268
use OAI21X1  _757_
timestamp 0
transform 1 0 4510 0 1 3390
box -6 -8 106 268
use NAND2X1  _758_
timestamp 0
transform 1 0 3290 0 -1 2870
box -6 -8 86 268
use OAI21X1  _759_
timestamp 0
transform -1 0 3530 0 -1 2870
box -6 -8 106 268
use NAND2X1  _760_
timestamp 0
transform 1 0 3390 0 -1 3910
box -6 -8 86 268
use OAI21X1  _761_
timestamp 0
transform -1 0 3630 0 -1 3910
box -6 -8 106 268
use NAND2X1  _762_
timestamp 0
transform 1 0 2970 0 -1 3910
box -6 -8 86 268
use OAI21X1  _763_
timestamp 0
transform -1 0 3070 0 -1 3390
box -6 -8 106 268
use NAND2X1  _764_
timestamp 0
transform 1 0 3090 0 1 3390
box -6 -8 86 268
use OAI21X1  _765_
timestamp 0
transform -1 0 3470 0 1 3390
box -6 -8 106 268
use INVX1  _766_
timestamp 0
transform 1 0 2190 0 -1 2350
box -6 -8 66 268
use NAND2X1  _767_
timestamp 0
transform -1 0 2170 0 1 1830
box -6 -8 86 268
use OAI21X1  _768_
timestamp 0
transform 1 0 1930 0 1 1830
box -6 -8 106 268
use INVX1  _769_
timestamp 0
transform -1 0 1650 0 -1 2870
box -6 -8 66 268
use NAND2X1  _770_
timestamp 0
transform 1 0 1850 0 1 2350
box -6 -8 86 268
use OAI21X1  _771_
timestamp 0
transform 1 0 1670 0 1 2350
box -6 -8 106 268
use INVX1  _772_
timestamp 0
transform -1 0 1070 0 1 2870
box -6 -8 66 268
use NAND2X1  _773_
timestamp 0
transform 1 0 1810 0 1 2870
box -6 -8 86 268
use OAI21X1  _774_
timestamp 0
transform -1 0 1370 0 1 2870
box -6 -8 106 268
use INVX1  _775_
timestamp 0
transform 1 0 730 0 -1 5470
box -6 -8 66 268
use NAND2X1  _776_
timestamp 0
transform 1 0 1430 0 1 2870
box -6 -8 86 268
use OAI21X1  _777_
timestamp 0
transform 1 0 850 0 -1 5470
box -6 -8 106 268
use INVX1  _778_
timestamp 0
transform -1 0 130 0 -1 5990
box -6 -8 66 268
use NAND2X1  _779_
timestamp 0
transform 1 0 1770 0 -1 3910
box -6 -8 86 268
use OAI21X1  _780_
timestamp 0
transform -1 0 430 0 -1 5470
box -6 -8 106 268
use INVX1  _781_
timestamp 0
transform -1 0 870 0 -1 4430
box -6 -8 66 268
use NAND2X1  _782_
timestamp 0
transform 1 0 1950 0 -1 2870
box -6 -8 86 268
use OAI21X1  _783_
timestamp 0
transform 1 0 1170 0 -1 4430
box -6 -8 106 268
use INVX1  _784_
timestamp 0
transform 1 0 710 0 -1 3910
box -6 -8 66 268
use NAND2X1  _785_
timestamp 0
transform 1 0 970 0 1 3390
box -6 -8 86 268
use OAI21X1  _786_
timestamp 0
transform 1 0 810 0 1 3390
box -6 -8 106 268
use INVX1  _787_
timestamp 0
transform 1 0 1350 0 1 3390
box -6 -8 66 268
use NAND2X1  _788_
timestamp 0
transform 1 0 1790 0 1 3390
box -6 -8 86 268
use OAI21X1  _789_
timestamp 0
transform 1 0 1470 0 1 3390
box -6 -8 106 268
use INVX1  _790_
timestamp 0
transform 1 0 2710 0 -1 1830
box -6 -8 66 268
use NAND2X1  _791_
timestamp 0
transform 1 0 2910 0 1 1830
box -6 -8 86 268
use OAI21X1  _792_
timestamp 0
transform 1 0 2830 0 -1 1830
box -6 -8 106 268
use INVX1  _793_
timestamp 0
transform 1 0 3170 0 1 1310
box -6 -8 66 268
use NAND2X1  _794_
timestamp 0
transform 1 0 3450 0 1 1310
box -6 -8 86 268
use OAI21X1  _795_
timestamp 0
transform 1 0 3290 0 1 1310
box -6 -8 106 268
use INVX1  _796_
timestamp 0
transform -1 0 1310 0 1 790
box -6 -8 66 268
use NAND2X1  _797_
timestamp 0
transform 1 0 2450 0 1 790
box -6 -8 86 268
use OAI21X1  _798_
timestamp 0
transform 1 0 1610 0 1 790
box -6 -8 106 268
use INVX1  _799_
timestamp 0
transform 1 0 870 0 -1 270
box -6 -8 66 268
use NAND2X1  _800_
timestamp 0
transform 1 0 1150 0 -1 270
box -6 -8 86 268
use OAI21X1  _801_
timestamp 0
transform 1 0 990 0 -1 270
box -6 -8 106 268
use INVX1  _802_
timestamp 0
transform -1 0 4090 0 1 790
box -6 -8 66 268
use NAND2X1  _803_
timestamp 0
transform -1 0 3750 0 -1 1830
box -6 -8 86 268
use OAI21X1  _804_
timestamp 0
transform -1 0 4110 0 -1 1310
box -6 -8 106 268
use INVX1  _805_
timestamp 0
transform -1 0 4210 0 1 270
box -6 -8 66 268
use NAND2X1  _806_
timestamp 0
transform -1 0 4110 0 -1 270
box -6 -8 86 268
use OAI21X1  _807_
timestamp 0
transform 1 0 4170 0 -1 270
box -6 -8 106 268
use INVX1  _808_
timestamp 0
transform -1 0 2390 0 -1 270
box -6 -8 66 268
use NAND2X1  _809_
timestamp 0
transform 1 0 2850 0 -1 270
box -6 -8 86 268
use OAI21X1  _810_
timestamp 0
transform 1 0 2690 0 -1 270
box -6 -8 106 268
use INVX1  _811_
timestamp 0
transform 1 0 2210 0 -1 270
box -6 -8 66 268
use NAND2X1  _812_
timestamp 0
transform -1 0 1750 0 -1 270
box -6 -8 86 268
use OAI21X1  _813_
timestamp 0
transform -1 0 1910 0 -1 270
box -6 -8 106 268
use INVX1  _814_
timestamp 0
transform -1 0 2190 0 1 2350
box -6 -8 66 268
use NAND3X1  _815_
timestamp 0
transform 1 0 2170 0 -1 3910
box -6 -8 106 268
use OAI21X1  _816_
timestamp 0
transform 1 0 2250 0 1 2350
box -6 -8 106 268
use INVX8  _817_
timestamp 0
transform 1 0 2030 0 -1 1830
box -6 -8 126 268
use NAND2X1  _818_
timestamp 0
transform 1 0 2390 0 1 3910
box -6 -8 86 268
use NAND2X1  _819_
timestamp 0
transform -1 0 2170 0 1 3910
box -6 -8 86 268
use XNOR2X1  _820_
timestamp 0
transform 1 0 1750 0 1 3910
box -6 -8 146 268
use NAND2X1  _821_
timestamp 0
transform 1 0 1570 0 -1 3390
box -6 -8 86 268
use OAI21X1  _822_
timestamp 0
transform -1 0 1810 0 -1 3390
box -6 -8 106 268
use NOR2X1  _823_
timestamp 0
transform 1 0 1950 0 1 3910
box -6 -8 86 268
use NAND2X1  _824_
timestamp 0
transform -1 0 1990 0 1 4430
box -6 -8 86 268
use NAND2X1  _825_
timestamp 0
transform 1 0 2710 0 -1 4430
box -6 -8 86 268
use NOR2X1  _826_
timestamp 0
transform 1 0 2110 0 -1 4430
box -6 -8 86 268
use AOI22X1  _827_
timestamp 0
transform 1 0 2530 0 1 3910
box -6 -8 126 268
use OAI21X1  _828_
timestamp 0
transform -1 0 2050 0 -1 4430
box -6 -8 106 268
use INVX1  _829_
timestamp 0
transform -1 0 1210 0 1 4430
box -6 -8 66 268
use AND2X2  _830_
timestamp 0
transform -1 0 2330 0 1 3910
box -6 -8 106 268
use AND2X2  _831_
timestamp 0
transform -1 0 2490 0 -1 4430
box -6 -8 106 268
use NAND2X1  _832_
timestamp 0
transform 1 0 2250 0 -1 4430
box -6 -8 86 268
use INVX1  _833_
timestamp 0
transform -1 0 3250 0 -1 4950
box -6 -8 66 268
use INVX1  _834_
timestamp 0
transform -1 0 2770 0 1 3910
box -6 -8 66 268
use NAND2X1  _835_
timestamp 0
transform -1 0 2610 0 1 4430
box -6 -8 86 268
use OAI21X1  _836_
timestamp 0
transform -1 0 2770 0 1 4430
box -6 -8 106 268
use NAND3X1  _837_
timestamp 0
transform -1 0 1370 0 1 4430
box -6 -8 106 268
use NAND3X1  _838_
timestamp 0
transform 1 0 1770 0 -1 4430
box -6 -8 106 268
use INVX1  _839_
timestamp 0
transform -1 0 1390 0 -1 4430
box -6 -8 66 268
use AOI21X1  _840_
timestamp 0
transform -1 0 1710 0 -1 4430
box -6 -8 106 268
use OAI21X1  _841_
timestamp 0
transform -1 0 1550 0 -1 4430
box -6 -8 106 268
use INVX1  _842_
timestamp 0
transform 1 0 1130 0 -1 3390
box -6 -8 66 268
use NAND2X1  _843_
timestamp 0
transform 1 0 1270 0 -1 3390
box -6 -8 86 268
use AND2X2  _844_
timestamp 0
transform -1 0 1510 0 -1 3390
box -6 -8 106 268
use INVX1  _845_
timestamp 0
transform 1 0 1050 0 1 4950
box -6 -8 66 268
use NAND2X1  _846_
timestamp 0
transform 1 0 3450 0 -1 4950
box -6 -8 86 268
use AOI21X1  _847_
timestamp 0
transform 1 0 1430 0 1 4430
box -6 -8 106 268
use NAND2X1  _848_
timestamp 0
transform 1 0 2170 0 1 4950
box -6 -8 86 268
use NAND2X1  _849_
timestamp 0
transform 1 0 2750 0 -1 4950
box -6 -8 86 268
use NOR2X1  _850_
timestamp 0
transform 1 0 2610 0 -1 4950
box -6 -8 86 268
use AOI22X1  _851_
timestamp 0
transform -1 0 2470 0 1 4430
box -6 -8 126 268
use OAI21X1  _852_
timestamp 0
transform 1 0 2450 0 -1 4950
box -6 -8 106 268
use INVX1  _853_
timestamp 0
transform 1 0 2170 0 -1 4950
box -6 -8 66 268
use AND2X2  _854_
timestamp 0
transform -1 0 2290 0 1 4430
box -6 -8 106 268
use NAND2X1  _855_
timestamp 0
transform -1 0 2130 0 1 4430
box -6 -8 86 268
use INVX1  _856_
timestamp 0
transform -1 0 2370 0 1 4950
box -6 -8 66 268
use NAND3X1  _857_
timestamp 0
transform -1 0 2110 0 -1 4950
box -6 -8 106 268
use NAND3X1  _858_
timestamp 0
transform -1 0 1790 0 1 4950
box -6 -8 106 268
use OAI21X1  _859_
timestamp 0
transform -1 0 1690 0 1 4430
box -6 -8 106 268
use AOI21X1  _860_
timestamp 0
transform -1 0 1950 0 -1 4950
box -6 -8 106 268
use INVX2  _861_
timestamp 0
transform -1 0 3770 0 -1 4430
box -6 -8 66 268
use OAI21X1  _862_
timestamp 0
transform -1 0 3090 0 -1 4430
box -6 -8 106 268
use INVX2  _863_
timestamp 0
transform -1 0 2630 0 1 3390
box -6 -8 66 268
use INVX1  _864_
timestamp 0
transform -1 0 2650 0 -1 3910
box -6 -8 66 268
use OAI21X1  _865_
timestamp 0
transform -1 0 2650 0 -1 4430
box -6 -8 106 268
use AOI21X1  _866_
timestamp 0
transform -1 0 1850 0 1 4430
box -6 -8 106 268
use OAI21X1  _867_
timestamp 0
transform 1 0 1690 0 -1 4950
box -6 -8 106 268
use NAND3X1  _868_
timestamp 0
transform -1 0 1610 0 1 4950
box -6 -8 106 268
use INVX1  _869_
timestamp 0
transform -1 0 1630 0 -1 5470
box -6 -8 66 268
use NAND3X1  _870_
timestamp 0
transform 1 0 2010 0 1 4950
box -6 -8 106 268
use OAI21X1  _871_
timestamp 0
transform -1 0 1630 0 -1 4950
box -6 -8 106 268
use NAND3X1  _872_
timestamp 0
transform -1 0 1510 0 -1 5470
box -6 -8 106 268
use AOI21X1  _873_
timestamp 0
transform -1 0 1470 0 -1 4950
box -6 -8 106 268
use NAND3X1  _874_
timestamp 0
transform -1 0 1450 0 1 4950
box -6 -8 106 268
use NAND2X1  _875_
timestamp 0
transform -1 0 1210 0 -1 5470
box -6 -8 86 268
use OAI22X1  _876_
timestamp 0
transform 1 0 1170 0 1 4950
box -6 -8 126 268
use INVX1  _877_
timestamp 0
transform 1 0 230 0 1 5470
box -6 -8 66 268
use INVX1  _878_
timestamp 0
transform -1 0 1070 0 -1 5470
box -6 -8 66 268
use AOI21X1  _879_
timestamp 0
transform -1 0 1950 0 1 4950
box -6 -8 106 268
use OAI21X1  _880_
timestamp 0
transform 1 0 1690 0 -1 5470
box -6 -8 106 268
use OAI21X1  _881_
timestamp 0
transform -1 0 2530 0 1 4950
box -6 -8 106 268
use AND2X2  _882_
timestamp 0
transform 1 0 3290 0 -1 4430
box -6 -8 106 268
use NAND2X1  _883_
timestamp 0
transform 1 0 2850 0 -1 4430
box -6 -8 86 268
use AOI22X1  _884_
timestamp 0
transform -1 0 2950 0 1 4430
box -6 -8 126 268
use INVX1  _885_
timestamp 0
transform -1 0 2390 0 -1 5470
box -6 -8 66 268
use NAND2X1  _886_
timestamp 0
transform 1 0 2730 0 1 4950
box -6 -8 86 268
use INVX1  _887_
timestamp 0
transform -1 0 2670 0 1 4950
box -6 -8 66 268
use NAND3X1  _888_
timestamp 0
transform -1 0 2550 0 -1 5470
box -6 -8 106 268
use NAND2X1  _889_
timestamp 0
transform -1 0 3230 0 -1 4430
box -6 -8 86 268
use NOR2X1  _890_
timestamp 0
transform 1 0 3050 0 1 4950
box -6 -8 86 268
use OAI21X1  _891_
timestamp 0
transform 1 0 2690 0 1 5470
box -6 -8 106 268
use AOI21X1  _892_
timestamp 0
transform -1 0 2470 0 1 5470
box -6 -8 106 268
use AOI21X1  _893_
timestamp 0
transform 1 0 2290 0 -1 4950
box -6 -8 106 268
use NAND3X1  _894_
timestamp 0
transform -1 0 2270 0 -1 5470
box -6 -8 106 268
use OAI21X1  _895_
timestamp 0
transform -1 0 2710 0 -1 5470
box -6 -8 106 268
use AOI21X1  _896_
timestamp 0
transform 1 0 2010 0 -1 5470
box -6 -8 106 268
use NAND2X1  _897_
timestamp 0
transform 1 0 3590 0 -1 4950
box -6 -8 86 268
use INVX1  _898_
timestamp 0
transform -1 0 2910 0 -1 3910
box -6 -8 66 268
use INVX2  _899_
timestamp 0
transform 1 0 3410 0 1 2870
box -6 -8 66 268
use NAND2X1  _900_
timestamp 0
transform 1 0 3450 0 -1 4430
box -6 -8 86 268
use OAI21X1  _901_
timestamp 0
transform 1 0 3030 0 1 4430
box -6 -8 106 268
use OAI21X1  _902_
timestamp 0
transform -1 0 3130 0 -1 4950
box -6 -8 106 268
use OAI21X1  _903_
timestamp 0
transform -1 0 2310 0 1 5470
box -6 -8 106 268
use NAND3X1  _904_
timestamp 0
transform -1 0 1950 0 -1 5470
box -6 -8 106 268
use NAND3X1  _905_
timestamp 0
transform 1 0 2530 0 1 5470
box -6 -8 106 268
use INVX1  _906_
timestamp 0
transform -1 0 2230 0 -1 5990
box -6 -8 66 268
use NAND3X1  _907_
timestamp 0
transform -1 0 2110 0 -1 5990
box -6 -8 106 268
use NAND3X1  _908_
timestamp 0
transform -1 0 1830 0 -1 5990
box -6 -8 106 268
use INVX1  _909_
timestamp 0
transform -1 0 1330 0 -1 5470
box -6 -8 66 268
use AOI21X1  _910_
timestamp 0
transform 1 0 1570 0 1 5470
box -6 -8 106 268
use AOI21X1  _911_
timestamp 0
transform -1 0 1990 0 1 5470
box -6 -8 106 268
use INVX1  _912_
timestamp 0
transform -1 0 1950 0 -1 5990
box -6 -8 66 268
use OAI21X1  _913_
timestamp 0
transform -1 0 1830 0 1 5470
box -6 -8 106 268
use AOI21X1  _914_
timestamp 0
transform -1 0 1350 0 1 5470
box -6 -8 106 268
use NAND3X1  _915_
timestamp 0
transform 1 0 1410 0 1 5470
box -6 -8 106 268
use NAND2X1  _916_
timestamp 0
transform 1 0 1110 0 1 5470
box -6 -8 86 268
use OAI22X1  _917_
timestamp 0
transform 1 0 770 0 1 5470
box -6 -8 126 268
use AND2X2  _918_
timestamp 0
transform -1 0 3970 0 -1 4950
box -6 -8 106 268
use NAND2X1  _919_
timestamp 0
transform -1 0 2850 0 -1 5470
box -6 -8 86 268
use INVX1  _920_
timestamp 0
transform 1 0 2770 0 -1 5990
box -6 -8 66 268
use AOI21X1  _921_
timestamp 0
transform 1 0 2050 0 1 5470
box -6 -8 106 268
use NAND2X1  _922_
timestamp 0
transform 1 0 3730 0 -1 4950
box -6 -8 86 268
use AND2X2  _923_
timestamp 0
transform -1 0 3450 0 1 4430
box -6 -8 106 268
use OAI21X1  _924_
timestamp 0
transform 1 0 3190 0 1 4430
box -6 -8 106 268
use INVX2  _925_
timestamp 0
transform 1 0 3590 0 -1 4430
box -6 -8 66 268
use OAI21X1  _926_
timestamp 0
transform -1 0 3910 0 1 4950
box -6 -8 106 268
use NAND3X1  _927_
timestamp 0
transform 1 0 3650 0 1 4950
box -6 -8 106 268
use INVX1  _928_
timestamp 0
transform -1 0 3590 0 1 4950
box -6 -8 66 268
use NAND2X1  _929_
timestamp 0
transform -1 0 3390 0 -1 4950
box -6 -8 86 268
use OAI21X1  _930_
timestamp 0
transform 1 0 3190 0 1 4950
box -6 -8 106 268
use NAND3X1  _931_
timestamp 0
transform 1 0 3370 0 1 4950
box -6 -8 106 268
use NAND2X1  _932_
timestamp 0
transform -1 0 3470 0 -1 5470
box -6 -8 86 268
use OAI22X1  _933_
timestamp 0
transform -1 0 2990 0 1 4950
box -6 -8 126 268
use INVX1  _934_
timestamp 0
transform -1 0 4330 0 1 4950
box -6 -8 66 268
use NAND2X1  _935_
timestamp 0
transform 1 0 4970 0 -1 4950
box -6 -8 86 268
use NAND3X1  _936_
timestamp 0
transform -1 0 4230 0 -1 4430
box -6 -8 106 268
use NAND2X1  _937_
timestamp 0
transform -1 0 4370 0 -1 4430
box -6 -8 86 268
use NAND3X1  _938_
timestamp 0
transform -1 0 4710 0 1 4430
box -6 -8 106 268
use NAND3X1  _939_
timestamp 0
transform -1 0 4770 0 1 4950
box -6 -8 106 268
use INVX1  _940_
timestamp 0
transform 1 0 5110 0 -1 4950
box -6 -8 66 268
use AND2X2  _941_
timestamp 0
transform -1 0 4550 0 -1 3910
box -6 -8 106 268
use NAND2X1  _942_
timestamp 0
transform 1 0 4430 0 -1 4430
box -6 -8 86 268
use OAI21X1  _943_
timestamp 0
transform -1 0 3930 0 -1 4430
box -6 -8 106 268
use NAND3X1  _944_
timestamp 0
transform 1 0 4650 0 -1 4950
box -6 -8 106 268
use NAND3X1  _945_
timestamp 0
transform -1 0 4270 0 -1 5470
box -6 -8 106 268
use AOI21X1  _946_
timestamp 0
transform -1 0 4590 0 -1 4950
box -6 -8 106 268
use AOI21X1  _947_
timestamp 0
transform 1 0 4830 0 1 4950
box -6 -8 106 268
use OAI21X1  _948_
timestamp 0
transform -1 0 3930 0 -1 5470
box -6 -8 106 268
use NAND3X1  _949_
timestamp 0
transform -1 0 3750 0 1 5470
box -6 -8 106 268
use AND2X2  _950_
timestamp 0
transform -1 0 3330 0 -1 5470
box -6 -8 106 268
use NAND3X1  _951_
timestamp 0
transform -1 0 4430 0 -1 5470
box -6 -8 106 268
use OAI21X1  _952_
timestamp 0
transform 1 0 3990 0 -1 5470
box -6 -8 106 268
use NAND3X1  _953_
timestamp 0
transform -1 0 3010 0 -1 5470
box -6 -8 106 268
use NAND3X1  _954_
timestamp 0
transform -1 0 3110 0 1 5470
box -6 -8 106 268
use OAI21X1  _955_
timestamp 0
transform 1 0 2450 0 -1 5990
box -6 -8 106 268
use AOI21X1  _956_
timestamp 0
transform -1 0 3170 0 -1 5470
box -6 -8 106 268
use AOI21X1  _957_
timestamp 0
transform -1 0 3590 0 1 5470
box -6 -8 106 268
use OAI21X1  _958_
timestamp 0
transform -1 0 3270 0 1 5470
box -6 -8 106 268
use NAND3X1  _959_
timestamp 0
transform -1 0 2950 0 1 5470
box -6 -8 106 268
use NAND3X1  _960_
timestamp 0
transform -1 0 3010 0 -1 5990
box -6 -8 106 268
use OAI21X1  _961_
timestamp 0
transform 1 0 3330 0 1 5470
box -6 -8 106 268
use NAND3X1  _962_
timestamp 0
transform -1 0 2710 0 -1 5990
box -6 -8 106 268
use NAND2X1  _963_
timestamp 0
transform -1 0 1490 0 -1 5990
box -6 -8 86 268
use NAND2X1  _964_
timestamp 0
transform -1 0 1350 0 -1 5990
box -6 -8 86 268
use XNOR2X1  _965_
timestamp 0
transform 1 0 1070 0 -1 5990
box -6 -8 146 268
use NAND2X1  _966_
timestamp 0
transform 1 0 870 0 1 4430
box -6 -8 86 268
use OAI21X1  _967_
timestamp 0
transform -1 0 1070 0 -1 4950
box -6 -8 106 268
use INVX1  _968_
timestamp 0
transform 1 0 210 0 -1 5470
box -6 -8 66 268
use AOI22X1  _969_
timestamp 0
transform -1 0 1670 0 -1 5990
box -6 -8 126 268
use AOI21X1  _970_
timestamp 0
transform 1 0 3070 0 -1 5990
box -6 -8 106 268
use OAI21X1  _971_
timestamp 0
transform 1 0 3230 0 -1 5990
box -6 -8 106 268
use NAND2X1  _972_
timestamp 0
transform 1 0 3670 0 1 4430
box -6 -8 86 268
use OAI21X1  _973_
timestamp 0
transform 1 0 3510 0 1 4430
box -6 -8 106 268
use INVX1  _974_
timestamp 0
transform -1 0 5350 0 -1 5990
box -6 -8 66 268
use INVX1  _975_
timestamp 0
transform -1 0 3610 0 -1 5470
box -6 -8 66 268
use AOI21X1  _976_
timestamp 0
transform 1 0 3670 0 -1 5470
box -6 -8 106 268
use NAND2X1  _977_
timestamp 0
transform 1 0 3970 0 1 4950
box -6 -8 86 268
use AND2X2  _978_
timestamp 0
transform -1 0 4230 0 1 4430
box -6 -8 106 268
use OAI21X1  _979_
timestamp 0
transform 1 0 3970 0 1 4430
box -6 -8 106 268
use AND2X2  _980_
timestamp 0
transform -1 0 4290 0 -1 4950
box -6 -8 106 268
use OAI21X1  _981_
timestamp 0
transform 1 0 4030 0 -1 4950
box -6 -8 106 268
use NAND3X1  _982_
timestamp 0
transform 1 0 4110 0 1 4950
box -6 -8 106 268
use INVX1  _983_
timestamp 0
transform -1 0 4450 0 1 4950
box -6 -8 66 268
use NAND2X1  _984_
timestamp 0
transform 1 0 4350 0 -1 4950
box -6 -8 86 268
use OAI21X1  _985_
timestamp 0
transform 1 0 3810 0 1 4430
box -6 -8 106 268
use NAND3X1  _986_
timestamp 0
transform 1 0 4510 0 1 4950
box -6 -8 106 268
use NAND2X1  _987_
timestamp 0
transform -1 0 5210 0 1 4950
box -6 -8 86 268
use NOR2X1  _988_
timestamp 0
transform 1 0 4290 0 1 4430
box -6 -8 86 268
use AOI21X1  _989_
timestamp 0
transform -1 0 4550 0 1 4430
box -6 -8 106 268
use NAND2X1  _990_
timestamp 0
transform 1 0 4830 0 1 3910
box -6 -8 86 268
use NAND2X1  _991_
timestamp 0
transform -1 0 4690 0 -1 3910
box -6 -8 86 268
use NAND3X1  _992_
timestamp 0
transform 1 0 4970 0 1 3910
box -6 -8 106 268
use NAND2X1  _993_
timestamp 0
transform -1 0 5210 0 1 3390
box -6 -8 86 268
use NAND3X1  _994_
timestamp 0
transform 1 0 5050 0 -1 3910
box -6 -8 106 268
use NAND3X1  _995_
timestamp 0
transform 1 0 5090 0 -1 4430
box -6 -8 106 268
use INVX1  _996_
timestamp 0
transform 1 0 5310 0 1 3910
box -6 -8 66 268
use AND2X2  _997_
timestamp 0
transform 1 0 4970 0 1 3390
box -6 -8 106 268
use NAND2X1  _998_
timestamp 0
transform -1 0 4990 0 -1 3910
box -6 -8 86 268
use OAI21X1  _999_
timestamp 0
transform 1 0 4750 0 -1 3910
box -6 -8 106 268
use NAND3X1  _1000_
timestamp 0
transform 1 0 5250 0 -1 4430
box -6 -8 106 268
use NAND3X1  _1001_
timestamp 0
transform -1 0 5190 0 1 4430
box -6 -8 106 268
use AOI22X1  _1002_
timestamp 0
transform -1 0 4690 0 -1 4430
box -6 -8 126 268
use OAI21X1  _1003_
timestamp 0
transform -1 0 4910 0 -1 4950
box -6 -8 106 268
use AOI22X1  _1004_
timestamp 0
transform 1 0 4750 0 -1 4430
box -6 -8 126 268
use AOI21X1  _1005_
timestamp 0
transform -1 0 5030 0 -1 4430
box -6 -8 106 268
use OAI21X1  _1006_
timestamp 0
transform -1 0 4870 0 1 4430
box -6 -8 106 268
use NAND3X1  _1007_
timestamp 0
transform -1 0 5330 0 -1 4950
box -6 -8 106 268
use AND2X2  _1008_
timestamp 0
transform 1 0 5270 0 1 4950
box -6 -8 106 268
use NAND3X1  _1009_
timestamp 0
transform 1 0 5570 0 -1 4950
box -6 -8 106 268
use OAI21X1  _1010_
timestamp 0
transform 1 0 4930 0 1 4430
box -6 -8 106 268
use NAND3X1  _1011_
timestamp 0
transform -1 0 5390 0 -1 5470
box -6 -8 106 268
use NAND3X1  _1012_
timestamp 0
transform 1 0 4970 0 -1 5470
box -6 -8 106 268
use AOI21X1  _1013_
timestamp 0
transform 1 0 4490 0 -1 5470
box -6 -8 106 268
use OAI21X1  _1014_
timestamp 0
transform 1 0 4650 0 -1 5470
box -6 -8 106 268
use AOI21X1  _1015_
timestamp 0
transform 1 0 5450 0 -1 5470
box -6 -8 106 268
use AOI21X1  _1016_
timestamp 0
transform 1 0 5390 0 -1 4950
box -6 -8 106 268
use OAI21X1  _1017_
timestamp 0
transform -1 0 5230 0 -1 5470
box -6 -8 106 268
use NAND3X1  _1018_
timestamp 0
transform -1 0 5070 0 -1 5990
box -6 -8 106 268
use NAND3X1  _1019_
timestamp 0
transform -1 0 5010 0 1 5470
box -6 -8 106 268
use OAI21X1  _1020_
timestamp 0
transform -1 0 4910 0 -1 5470
box -6 -8 106 268
use NAND3X1  _1021_
timestamp 0
transform -1 0 4910 0 -1 5990
box -6 -8 106 268
use NAND2X1  _1022_
timestamp 0
transform 1 0 4510 0 -1 5990
box -6 -8 86 268
use XNOR2X1  _1023_
timestamp 0
transform -1 0 3810 0 -1 5990
box -6 -8 146 268
use NOR2X1  _1024_
timestamp 0
transform 1 0 2310 0 -1 5990
box -6 -8 86 268
use NAND3X1  _1025_
timestamp 0
transform -1 0 4450 0 -1 5990
box -6 -8 106 268
use INVX1  _1026_
timestamp 0
transform 1 0 3390 0 -1 5990
box -6 -8 66 268
use AOI21X1  _1027_
timestamp 0
transform 1 0 3510 0 -1 5990
box -6 -8 106 268
use AOI21X1  _1028_
timestamp 0
transform -1 0 4750 0 -1 5990
box -6 -8 106 268
use AOI21X1  _1029_
timestamp 0
transform 1 0 5130 0 -1 5990
box -6 -8 106 268
use OAI21X1  _1030_
timestamp 0
transform -1 0 4290 0 -1 5990
box -6 -8 106 268
use NAND3X1  _1031_
timestamp 0
transform -1 0 4130 0 -1 5990
box -6 -8 106 268
use NAND2X1  _1032_
timestamp 0
transform 1 0 950 0 1 5470
box -6 -8 86 268
use OAI22X1  _1033_
timestamp 0
transform 1 0 590 0 1 5470
box -6 -8 126 268
use OAI21X1  _1034_
timestamp 0
transform 1 0 3870 0 -1 5990
box -6 -8 106 268
use INVX1  _1035_
timestamp 0
transform 1 0 5410 0 -1 5990
box -6 -8 66 268
use AOI21X1  _1036_
timestamp 0
transform 1 0 5530 0 -1 5990
box -6 -8 106 268
use NAND2X1  _1037_
timestamp 0
transform 1 0 4990 0 1 4950
box -6 -8 86 268
use INVX1  _1038_
timestamp 0
transform 1 0 5850 0 1 270
box -6 -8 66 268
use INVX1  _1039_
timestamp 0
transform -1 0 5670 0 1 4950
box -6 -8 66 268
use AOI21X1  _1040_
timestamp 0
transform 1 0 5430 0 1 4950
box -6 -8 106 268
use NAND2X1  _1041_
timestamp 0
transform -1 0 4250 0 -1 3910
box -6 -8 86 268
use AND2X2  _1042_
timestamp 0
transform 1 0 4210 0 1 2870
box -6 -8 106 268
use OAI21X1  _1043_
timestamp 0
transform 1 0 4090 0 -1 3390
box -6 -8 106 268
use AND2X2  _1044_
timestamp 0
transform -1 0 4030 0 1 3390
box -6 -8 106 268
use OAI21X1  _1045_
timestamp 0
transform 1 0 3770 0 1 3390
box -6 -8 106 268
use NAND3X1  _1046_
timestamp 0
transform -1 0 4190 0 1 3390
box -6 -8 106 268
use INVX1  _1047_
timestamp 0
transform 1 0 4250 0 1 3390
box -6 -8 66 268
use NAND2X1  _1048_
timestamp 0
transform 1 0 4250 0 -1 3390
box -6 -8 86 268
use NAND2X1  _1049_
timestamp 0
transform -1 0 3870 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1050_
timestamp 0
transform -1 0 4030 0 -1 3390
box -6 -8 106 268
use NAND3X1  _1051_
timestamp 0
transform 1 0 4390 0 -1 3390
box -6 -8 106 268
use NAND2X1  _1052_
timestamp 0
transform -1 0 5350 0 1 3390
box -6 -8 86 268
use AOI22X1  _1053_
timestamp 0
transform 1 0 5230 0 -1 3910
box -6 -8 126 268
use NAND2X1  _1054_
timestamp 0
transform -1 0 5070 0 1 2870
box -6 -8 86 268
use NAND2X1  _1055_
timestamp 0
transform -1 0 5210 0 1 2870
box -6 -8 86 268
use NOR2X1  _1056_
timestamp 0
transform 1 0 5370 0 -1 3390
box -6 -8 86 268
use AOI22X1  _1057_
timestamp 0
transform 1 0 5190 0 -1 3390
box -6 -8 126 268
use OAI21X1  _1058_
timestamp 0
transform -1 0 5750 0 -1 3390
box -6 -8 106 268
use INVX1  _1059_
timestamp 0
transform -1 0 5690 0 1 2870
box -6 -8 66 268
use AND2X2  _1060_
timestamp 0
transform -1 0 5130 0 -1 3390
box -6 -8 106 268
use NAND2X1  _1061_
timestamp 0
transform 1 0 5510 0 -1 3390
box -6 -8 86 268
use INVX1  _1062_
timestamp 0
transform 1 0 5750 0 1 2870
box -6 -8 66 268
use NAND3X1  _1063_
timestamp 0
transform 1 0 5810 0 -1 3390
box -6 -8 106 268
use NAND3X1  _1064_
timestamp 0
transform 1 0 5730 0 -1 3910
box -6 -8 106 268
use AOI22X1  _1065_
timestamp 0
transform 1 0 5130 0 1 3910
box -6 -8 126 268
use OAI21X1  _1066_
timestamp 0
transform -1 0 5530 0 1 3910
box -6 -8 106 268
use AOI21X1  _1067_
timestamp 0
transform -1 0 5670 0 1 3390
box -6 -8 106 268
use OAI21X1  _1068_
timestamp 0
transform 1 0 4710 0 -1 3390
box -6 -8 106 268
use OAI21X1  _1069_
timestamp 0
transform 1 0 4810 0 1 3390
box -6 -8 106 268
use AOI21X1  _1070_
timestamp 0
transform 1 0 4870 0 -1 3390
box -6 -8 106 268
use OAI21X1  _1071_
timestamp 0
transform 1 0 5570 0 -1 3910
box -6 -8 106 268
use NAND3X1  _1072_
timestamp 0
transform 1 0 5590 0 1 3910
box -6 -8 106 268
use AND2X2  _1073_
timestamp 0
transform 1 0 5410 0 1 3390
box -6 -8 106 268
use NAND3X1  _1074_
timestamp 0
transform 1 0 5690 0 1 270
box -6 -8 106 268
use OAI21X1  _1075_
timestamp 0
transform -1 0 5510 0 -1 3910
box -6 -8 106 268
use NAND3X1  _1076_
timestamp 0
transform -1 0 5810 0 -1 4430
box -6 -8 106 268
use NAND3X1  _1077_
timestamp 0
transform 1 0 5730 0 1 4950
box -6 -8 106 268
use AOI21X1  _1078_
timestamp 0
transform 1 0 5250 0 1 4430
box -6 -8 106 268
use OAI21X1  _1079_
timestamp 0
transform 1 0 5730 0 -1 4950
box -6 -8 106 268
use AOI21X1  _1080_
timestamp 0
transform 1 0 5870 0 -1 4430
box -6 -8 106 268
use AOI21X1  _1081_
timestamp 0
transform 1 0 5550 0 -1 4430
box -6 -8 106 268
use OAI21X1  _1082_
timestamp 0
transform 1 0 5690 0 -1 5990
box -6 -8 106 268
use AOI21X1  _1083_
timestamp 0
transform -1 0 5830 0 1 5470
box -6 -8 106 268
use NAND3X1  _1084_
timestamp 0
transform 1 0 5730 0 1 4430
box -6 -8 106 268
use OAI21X1  _1085_
timestamp 0
transform -1 0 5870 0 -1 270
box -6 -8 106 268
use AOI21X1  _1086_
timestamp 0
transform -1 0 5710 0 -1 5470
box -6 -8 106 268
use OAI21X1  _1087_
timestamp 0
transform -1 0 5650 0 1 5470
box -6 -8 106 268
use AOI21X1  _1088_
timestamp 0
transform 1 0 5070 0 1 5470
box -6 -8 106 268
use OAI21X1  _1089_
timestamp 0
transform 1 0 5230 0 1 5470
box -6 -8 106 268
use NAND3X1  _1090_
timestamp 0
transform -1 0 5870 0 -1 5470
box -6 -8 106 268
use NAND3X1  _1091_
timestamp 0
transform 1 0 5850 0 -1 5990
box -6 -8 106 268
use NAND3X1  _1092_
timestamp 0
transform 1 0 5390 0 1 5470
box -6 -8 106 268
use NAND2X1  _1093_
timestamp 0
transform 1 0 4610 0 1 5470
box -6 -8 86 268
use XOR2X1  _1094_
timestamp 0
transform -1 0 3950 0 1 5470
box -6 -8 146 268
use NAND2X1  _1095_
timestamp 0
transform 1 0 1630 0 -1 3910
box -6 -8 86 268
use OAI21X1  _1096_
timestamp 0
transform -1 0 1690 0 1 3910
box -6 -8 106 268
use NAND2X1  _1097_
timestamp 0
transform 1 0 3850 0 1 1310
box -6 -8 86 268
use NAND2X1  _1098_
timestamp 0
transform -1 0 4410 0 1 5470
box -6 -8 86 268
use NAND2X1  _1099_
timestamp 0
transform -1 0 4550 0 1 5470
box -6 -8 86 268
use OAI21X1  _1100_
timestamp 0
transform 1 0 4170 0 1 5470
box -6 -8 106 268
use AOI21X1  _1101_
timestamp 0
transform -1 0 5670 0 1 4430
box -6 -8 106 268
use OAI21X1  _1102_
timestamp 0
transform 1 0 5410 0 1 4430
box -6 -8 106 268
use NAND2X1  _1103_
timestamp 0
transform 1 0 4550 0 -1 3390
box -6 -8 86 268
use INVX1  _1104_
timestamp 0
transform 1 0 5890 0 -1 790
box -6 -8 66 268
use INVX1  _1105_
timestamp 0
transform -1 0 5970 0 1 3910
box -6 -8 66 268
use AOI21X1  _1106_
timestamp 0
transform -1 0 5850 0 1 3910
box -6 -8 106 268
use INVX2  _1107_
timestamp 0
transform -1 0 3870 0 1 2870
box -6 -8 66 268
use NOR2X1  _1108_
timestamp 0
transform 1 0 4190 0 -1 2870
box -6 -8 86 268
use AND2X2  _1109_
timestamp 0
transform -1 0 4910 0 -1 2870
box -6 -8 106 268
use AOI22X1  _1110_
timestamp 0
transform -1 0 4490 0 1 2870
box -6 -8 126 268
use AOI21X1  _1111_
timestamp 0
transform 1 0 4470 0 -1 2870
box -6 -8 106 268
use XNOR2X1  _1112_
timestamp 0
transform 1 0 4590 0 1 2350
box -6 -8 146 268
use AOI21X1  _1113_
timestamp 0
transform 1 0 5870 0 1 2870
box -6 -8 106 268
use NAND2X1  _1114_
timestamp 0
transform 1 0 5130 0 -1 2870
box -6 -8 86 268
use NAND2X1  _1115_
timestamp 0
transform 1 0 4850 0 1 2870
box -6 -8 86 268
use NAND2X1  _1116_
timestamp 0
transform -1 0 4630 0 1 2870
box -6 -8 86 268
use OAI21X1  _1117_
timestamp 0
transform 1 0 4690 0 1 2870
box -6 -8 106 268
use OAI21X1  _1118_
timestamp 0
transform -1 0 5070 0 -1 2870
box -6 -8 106 268
use NOR2X1  _1119_
timestamp 0
transform 1 0 5610 0 -1 790
box -6 -8 86 268
use OAI21X1  _1120_
timestamp 0
transform 1 0 5470 0 1 2870
box -6 -8 106 268
use XOR2X1  _1121_
timestamp 0
transform -1 0 5410 0 1 2870
box -6 -8 146 268
use NOR2X1  _1122_
timestamp 0
transform 1 0 5590 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1123_
timestamp 0
transform 1 0 5590 0 1 2350
box -6 -8 106 268
use XOR2X1  _1124_
timestamp 0
transform 1 0 5090 0 1 2350
box -6 -8 146 268
use OAI21X1  _1125_
timestamp 0
transform -1 0 5530 0 -1 2870
box -6 -8 106 268
use NAND2X1  _1126_
timestamp 0
transform 1 0 5450 0 1 2350
box -6 -8 86 268
use NAND3X1  _1127_
timestamp 0
transform 1 0 5110 0 -1 2350
box -6 -8 106 268
use NAND3X1  _1128_
timestamp 0
transform 1 0 5750 0 -1 2350
box -6 -8 106 268
use AOI21X1  _1129_
timestamp 0
transform 1 0 5610 0 -1 270
box -6 -8 106 268
use OAI21X1  _1130_
timestamp 0
transform 1 0 5730 0 1 3390
box -6 -8 106 268
use AOI21X1  _1131_
timestamp 0
transform 1 0 5270 0 -1 2350
box -6 -8 106 268
use NAND2X1  _1132_
timestamp 0
transform 1 0 5890 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1133_
timestamp 0
transform 1 0 5730 0 -1 2870
box -6 -8 106 268
use AOI21X1  _1134_
timestamp 0
transform 1 0 5750 0 1 2350
box -6 -8 106 268
use OAI21X1  _1135_
timestamp 0
transform 1 0 5590 0 -1 2350
box -6 -8 106 268
use NAND3X1  _1136_
timestamp 0
transform 1 0 5810 0 1 790
box -6 -8 106 268
use NAND3X1  _1137_
timestamp 0
transform -1 0 5790 0 1 1830
box -6 -8 106 268
use OAI21X1  _1138_
timestamp 0
transform -1 0 5530 0 -1 2350
box -6 -8 106 268
use NAND3X1  _1139_
timestamp 0
transform 1 0 5230 0 1 1830
box -6 -8 106 268
use NAND3X1  _1140_
timestamp 0
transform 1 0 5570 0 -1 1830
box -6 -8 106 268
use INVX1  _1141_
timestamp 0
transform 1 0 5410 0 1 1830
box -6 -8 66 268
use AOI21X1  _1142_
timestamp 0
transform 1 0 5530 0 1 1830
box -6 -8 106 268
use AOI21X1  _1143_
timestamp 0
transform -1 0 5830 0 -1 1830
box -6 -8 106 268
use OAI21X1  _1144_
timestamp 0
transform -1 0 5510 0 -1 1830
box -6 -8 106 268
use NAND2X1  _1145_
timestamp 0
transform 1 0 5310 0 1 1310
box -6 -8 86 268
use XOR2X1  _1146_
timestamp 0
transform 1 0 4630 0 1 1310
box -6 -8 146 268
use OAI21X1  _1147_
timestamp 0
transform -1 0 4090 0 1 1310
box -6 -8 106 268
use INVX1  _1148_
timestamp 0
transform -1 0 5250 0 1 1310
box -6 -8 66 268
use AOI21X1  _1149_
timestamp 0
transform -1 0 5130 0 1 1310
box -6 -8 106 268
use AOI22X1  _1150_
timestamp 0
transform 1 0 4630 0 -1 2870
box -6 -8 126 268
use INVX1  _1151_
timestamp 0
transform 1 0 4450 0 1 1830
box -6 -8 66 268
use OAI21X1  _1152_
timestamp 0
transform -1 0 5390 0 1 2350
box -6 -8 106 268
use NOR2X1  _1153_
timestamp 0
transform -1 0 3230 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1154_
timestamp 0
transform -1 0 3610 0 1 2870
box -6 -8 86 268
use NAND2X1  _1155_
timestamp 0
transform 1 0 4050 0 -1 2870
box -6 -8 86 268
use OR2X2  _1156_
timestamp 0
transform -1 0 3570 0 1 2350
box -6 -8 106 268
use OAI21X1  _1157_
timestamp 0
transform 1 0 3590 0 -1 2870
box -6 -8 106 268
use NAND3X1  _1158_
timestamp 0
transform 1 0 3290 0 -1 2350
box -6 -8 106 268
use NAND2X1  _1159_
timestamp 0
transform 1 0 4430 0 1 2350
box -6 -8 86 268
use NAND2X1  _1160_
timestamp 0
transform 1 0 4330 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1161_
timestamp 0
transform -1 0 4370 0 1 2350
box -6 -8 106 268
use OAI21X1  _1162_
timestamp 0
transform 1 0 3610 0 -1 2350
box -6 -8 106 268
use NAND2X1  _1163_
timestamp 0
transform -1 0 3850 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1164_
timestamp 0
transform -1 0 4890 0 1 2350
box -6 -8 106 268
use NOR2X1  _1165_
timestamp 0
transform 1 0 4950 0 1 2350
box -6 -8 86 268
use NAND3X1  _1166_
timestamp 0
transform -1 0 4390 0 -1 2350
box -6 -8 106 268
use NAND3X1  _1167_
timestamp 0
transform -1 0 4710 0 -1 2350
box -6 -8 106 268
use AOI21X1  _1168_
timestamp 0
transform -1 0 5030 0 -1 2350
box -6 -8 106 268
use AOI21X1  _1169_
timestamp 0
transform 1 0 4450 0 -1 2350
box -6 -8 106 268
use INVX1  _1170_
timestamp 0
transform -1 0 4390 0 1 1830
box -6 -8 66 268
use OAI21X1  _1171_
timestamp 0
transform 1 0 4750 0 1 1830
box -6 -8 106 268
use NAND3X1  _1172_
timestamp 0
transform 1 0 4570 0 1 1830
box -6 -8 106 268
use NAND3X1  _1173_
timestamp 0
transform 1 0 4770 0 -1 2350
box -6 -8 106 268
use OAI21X1  _1174_
timestamp 0
transform 1 0 4910 0 1 1830
box -6 -8 106 268
use NAND3X1  _1175_
timestamp 0
transform 1 0 5070 0 1 1830
box -6 -8 106 268
use NAND2X1  _1176_
timestamp 0
transform -1 0 5190 0 -1 1830
box -6 -8 86 268
use NAND3X1  _1177_
timestamp 0
transform 1 0 5250 0 -1 1830
box -6 -8 106 268
use AOI21X1  _1178_
timestamp 0
transform 1 0 5850 0 1 1830
box -6 -8 106 268
use OAI21X1  _1179_
timestamp 0
transform -1 0 5870 0 1 1310
box -6 -8 106 268
use NAND3X1  _1180_
timestamp 0
transform 1 0 5610 0 1 1310
box -6 -8 106 268
use AND2X2  _1181_
timestamp 0
transform -1 0 5550 0 1 1310
box -6 -8 106 268
use XOR2X1  _1182_
timestamp 0
transform -1 0 4970 0 1 1310
box -6 -8 146 268
use NAND2X1  _1183_
timestamp 0
transform 1 0 4170 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1184_
timestamp 0
transform -1 0 4410 0 -1 1310
box -6 -8 106 268
use INVX1  _1185_
timestamp 0
transform -1 0 1450 0 -1 790
box -6 -8 66 268
use NAND2X1  _1186_
timestamp 0
transform 1 0 5510 0 -1 1310
box -6 -8 86 268
use NOR2X1  _1187_
timestamp 0
transform -1 0 5450 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1188_
timestamp 0
transform 1 0 5790 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1189_
timestamp 0
transform 1 0 5650 0 -1 1310
box -6 -8 86 268
use INVX1  _1190_
timestamp 0
transform -1 0 5750 0 1 790
box -6 -8 66 268
use AOI21X1  _1191_
timestamp 0
transform 1 0 5210 0 -1 1310
box -6 -8 106 268
use NAND2X1  _1192_
timestamp 0
transform -1 0 4570 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1193_
timestamp 0
transform -1 0 4230 0 -1 2350
box -6 -8 106 268
use INVX1  _1194_
timestamp 0
transform 1 0 5490 0 -1 270
box -6 -8 66 268
use OR2X2  _1195_
timestamp 0
transform 1 0 5270 0 -1 2870
box -6 -8 106 268
use NOR2X1  _1196_
timestamp 0
transform -1 0 4150 0 1 2870
box -6 -8 86 268
use OAI21X1  _1197_
timestamp 0
transform -1 0 3990 0 -1 2870
box -6 -8 106 268
use NAND2X1  _1198_
timestamp 0
transform 1 0 3930 0 1 2870
box -6 -8 86 268
use OAI21X1  _1199_
timestamp 0
transform 1 0 3810 0 1 2350
box -6 -8 106 268
use XOR2X1  _1200_
timestamp 0
transform 1 0 3930 0 -1 2350
box -6 -8 146 268
use AOI21X1  _1201_
timestamp 0
transform -1 0 4730 0 -1 1830
box -6 -8 106 268
use NAND3X1  _1202_
timestamp 0
transform 1 0 4790 0 -1 1830
box -6 -8 106 268
use INVX1  _1203_
timestamp 0
transform 1 0 5430 0 1 270
box -6 -8 66 268
use OAI21X1  _1204_
timestamp 0
transform 1 0 5330 0 -1 270
box -6 -8 106 268
use INVX1  _1205_
timestamp 0
transform 1 0 5310 0 1 270
box -6 -8 66 268
use NAND3X1  _1206_
timestamp 0
transform 1 0 5150 0 1 270
box -6 -8 106 268
use AND2X2  _1207_
timestamp 0
transform -1 0 5270 0 -1 270
box -6 -8 106 268
use NAND2X1  _1208_
timestamp 0
transform -1 0 5090 0 1 270
box -6 -8 86 268
use OR2X2  _1209_
timestamp 0
transform -1 0 5110 0 -1 270
box -6 -8 106 268
use NAND2X1  _1210_
timestamp 0
transform 1 0 4870 0 -1 270
box -6 -8 86 268
use NAND2X1  _1211_
timestamp 0
transform 1 0 4810 0 -1 790
box -6 -8 86 268
use AND2X2  _1212_
timestamp 0
transform -1 0 4850 0 1 5470
box -6 -8 106 268
use NAND3X1  _1213_
timestamp 0
transform 1 0 4010 0 1 5470
box -6 -8 106 268
use NAND3X1  _1214_
timestamp 0
transform -1 0 5050 0 -1 1830
box -6 -8 106 268
use AOI21X1  _1215_
timestamp 0
transform 1 0 4170 0 1 1830
box -6 -8 106 268
use INVX1  _1216_
timestamp 0
transform -1 0 5470 0 1 790
box -6 -8 66 268
use OAI21X1  _1217_
timestamp 0
transform 1 0 5250 0 1 790
box -6 -8 106 268
use NAND3X1  _1218_
timestamp 0
transform -1 0 4750 0 -1 790
box -6 -8 106 268
use OAI21X1  _1219_
timestamp 0
transform 1 0 1750 0 -1 790
box -6 -8 106 268
use NAND2X1  _1220_
timestamp 0
transform 1 0 670 0 1 270
box -6 -8 86 268
use AOI21X1  _1221_
timestamp 0
transform 1 0 5150 0 -1 790
box -6 -8 106 268
use INVX1  _1222_
timestamp 0
transform 1 0 4150 0 1 2350
box -6 -8 66 268
use OAI22X1  _1223_
timestamp 0
transform 1 0 3970 0 1 2350
box -6 -8 126 268
use OAI21X1  _1224_
timestamp 0
transform 1 0 3450 0 -1 2350
box -6 -8 106 268
use NOR2X1  _1225_
timestamp 0
transform 1 0 3750 0 -1 2870
box -6 -8 86 268
use INVX1  _1226_
timestamp 0
transform -1 0 3810 0 1 1830
box -6 -8 66 268
use OR2X2  _1227_
timestamp 0
transform 1 0 3870 0 1 1830
box -6 -8 106 268
use AND2X2  _1228_
timestamp 0
transform -1 0 3690 0 1 1830
box -6 -8 106 268
use XNOR2X1  _1229_
timestamp 0
transform -1 0 4430 0 -1 1830
box -6 -8 146 268
use XOR2X1  _1230_
timestamp 0
transform 1 0 4950 0 -1 790
box -6 -8 146 268
use INVX1  _1231_
timestamp 0
transform 1 0 4730 0 1 270
box -6 -8 66 268
use NAND3X1  _1232_
timestamp 0
transform -1 0 4670 0 1 270
box -6 -8 106 268
use OAI21X1  _1233_
timestamp 0
transform -1 0 4810 0 -1 270
box -6 -8 106 268
use NAND2X1  _1234_
timestamp 0
transform -1 0 4650 0 -1 270
box -6 -8 86 268
use NAND3X1  _1235_
timestamp 0
transform -1 0 4510 0 1 270
box -6 -8 106 268
use NAND2X1  _1236_
timestamp 0
transform 1 0 810 0 1 270
box -6 -8 86 268
use INVX1  _1237_
timestamp 0
transform -1 0 4450 0 1 790
box -6 -8 66 268
use NOR2X1  _1238_
timestamp 0
transform 1 0 5750 0 -1 790
box -6 -8 86 268
use AOI21X1  _1239_
timestamp 0
transform 1 0 5310 0 -1 790
box -6 -8 106 268
use NOR2X1  _1240_
timestamp 0
transform -1 0 5550 0 -1 790
box -6 -8 86 268
use NAND3X1  _1241_
timestamp 0
transform 1 0 4850 0 1 270
box -6 -8 106 268
use OAI21X1  _1242_
timestamp 0
transform 1 0 4930 0 -1 1310
box -6 -8 106 268
use NAND2X1  _1243_
timestamp 0
transform -1 0 4050 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1244_
timestamp 0
transform 1 0 3650 0 1 2350
box -6 -8 106 268
use OR2X2  _1245_
timestamp 0
transform -1 0 3910 0 -1 1830
box -6 -8 106 268
use INVX1  _1246_
timestamp 0
transform 1 0 4030 0 1 1830
box -6 -8 66 268
use OAI21X1  _1247_
timestamp 0
transform 1 0 4110 0 -1 1830
box -6 -8 106 268
use AND2X2  _1248_
timestamp 0
transform 1 0 4150 0 1 1310
box -6 -8 106 268
use NOR2X1  _1249_
timestamp 0
transform 1 0 4670 0 -1 1310
box -6 -8 86 268
use INVX1  _1250_
timestamp 0
transform 1 0 5090 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1251_
timestamp 0
transform -1 0 5630 0 1 790
box -6 -8 106 268
use AOI21X1  _1252_
timestamp 0
transform -1 0 5190 0 1 790
box -6 -8 106 268
use INVX1  _1253_
timestamp 0
transform 1 0 4810 0 -1 1310
box -6 -8 66 268
use OAI21X1  _1254_
timestamp 0
transform 1 0 4930 0 1 790
box -6 -8 106 268
use OAI22X1  _1255_
timestamp 0
transform 1 0 4750 0 1 790
box -6 -8 126 268
use INVX1  _1256_
timestamp 0
transform -1 0 4350 0 -1 790
box -6 -8 66 268
use AOI21X1  _1257_
timestamp 0
transform -1 0 4570 0 1 1310
box -6 -8 106 268
use AND2X2  _1258_
timestamp 0
transform 1 0 4310 0 1 1310
box -6 -8 106 268
use AOI22X1  _1259_
timestamp 0
transform 1 0 4490 0 -1 1310
box -6 -8 126 268
use NOR2X1  _1260_
timestamp 0
transform 1 0 1810 0 -1 2350
box -6 -8 86 268
use INVX1  _1261_
timestamp 0
transform 1 0 1250 0 -1 2350
box -6 -8 66 268
use NAND2X1  _1262_
timestamp 0
transform -1 0 1630 0 1 1830
box -6 -8 86 268
use NAND2X1  _1263_
timestamp 0
transform -1 0 1490 0 1 1830
box -6 -8 86 268
use NAND2X1  _1264_
timestamp 0
transform -1 0 1030 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1265_
timestamp 0
transform -1 0 1430 0 -1 1830
box -6 -8 106 268
use INVX1  _1266_
timestamp 0
transform -1 0 1530 0 -1 2870
box -6 -8 66 268
use NOR2X1  _1267_
timestamp 0
transform -1 0 1410 0 -1 2870
box -6 -8 86 268
use NOR2X1  _1268_
timestamp 0
transform -1 0 1370 0 1 2350
box -6 -8 86 268
use NOR2X1  _1269_
timestamp 0
transform -1 0 1070 0 1 2350
box -6 -8 86 268
use NAND2X1  _1270_
timestamp 0
transform -1 0 1190 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1271_
timestamp 0
transform 1 0 1130 0 1 2350
box -6 -8 106 268
use NAND2X1  _1272_
timestamp 0
transform -1 0 1050 0 -1 2350
box -6 -8 86 268
use NAND2X1  _1273_
timestamp 0
transform 1 0 670 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1274_
timestamp 0
transform -1 0 910 0 -1 2350
box -6 -8 106 268
use OAI21X1  _1275_
timestamp 0
transform -1 0 1270 0 -1 2870
box -6 -8 106 268
use XOR2X1  _1276_
timestamp 0
transform -1 0 950 0 1 2870
box -6 -8 146 268
use XNOR2X1  _1277_
timestamp 0
transform 1 0 610 0 1 2870
box -6 -8 146 268
use NAND2X1  _1278_
timestamp 0
transform -1 0 550 0 1 2350
box -6 -8 86 268
use OAI21X1  _1279_
timestamp 0
transform -1 0 710 0 -1 2870
box -6 -8 106 268
use NOR2X1  _1280_
timestamp 0
transform 1 0 990 0 -1 3390
box -6 -8 86 268
use AOI21X1  _1281_
timestamp 0
transform -1 0 930 0 -1 3390
box -6 -8 106 268
use NOR2X1  _1282_
timestamp 0
transform 1 0 770 0 1 4950
box -6 -8 86 268
use NOR2X1  _1283_
timestamp 0
transform 1 0 910 0 1 4950
box -6 -8 86 268
use NOR2X1  _1284_
timestamp 0
transform 1 0 630 0 1 4950
box -6 -8 86 268
use XOR2X1  _1285_
timestamp 0
transform -1 0 510 0 1 3390
box -6 -8 146 268
use NAND2X1  _1286_
timestamp 0
transform 1 0 310 0 -1 2870
box -6 -8 86 268
use OAI21X1  _1287_
timestamp 0
transform -1 0 410 0 1 2870
box -6 -8 106 268
use NAND2X1  _1288_
timestamp 0
transform 1 0 790 0 -1 2870
box -6 -8 86 268
use NAND2X1  _1289_
timestamp 0
transform 1 0 70 0 -1 5470
box -6 -8 86 268
use NAND2X1  _1290_
timestamp 0
transform 1 0 190 0 -1 5990
box -6 -8 86 268
use AND2X2  _1291_
timestamp 0
transform 1 0 70 0 1 5470
box -6 -8 106 268
use INVX1  _1292_
timestamp 0
transform -1 0 130 0 1 4950
box -6 -8 66 268
use INVX1  _1293_
timestamp 0
transform -1 0 670 0 -1 4950
box -6 -8 66 268
use OAI21X1  _1294_
timestamp 0
transform -1 0 550 0 -1 4950
box -6 -8 106 268
use INVX1  _1295_
timestamp 0
transform 1 0 210 0 -1 4950
box -6 -8 66 268
use NAND2X1  _1296_
timestamp 0
transform 1 0 70 0 -1 4950
box -6 -8 86 268
use NAND2X1  _1297_
timestamp 0
transform 1 0 190 0 1 4950
box -6 -8 86 268
use NAND2X1  _1298_
timestamp 0
transform 1 0 490 0 1 4950
box -6 -8 86 268
use OAI21X1  _1299_
timestamp 0
transform 1 0 450 0 -1 2870
box -6 -8 106 268
use NAND2X1  _1300_
timestamp 0
transform -1 0 530 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1301_
timestamp 0
transform 1 0 330 0 1 4950
box -6 -8 106 268
use OR2X2  _1302_
timestamp 0
transform -1 0 670 0 1 4430
box -6 -8 106 268
use NAND2X1  _1303_
timestamp 0
transform 1 0 730 0 1 4430
box -6 -8 86 268
use AND2X2  _1304_
timestamp 0
transform -1 0 490 0 1 4430
box -6 -8 106 268
use NOR2X1  _1305_
timestamp 0
transform -1 0 570 0 -1 4430
box -6 -8 86 268
use INVX1  _1306_
timestamp 0
transform -1 0 390 0 -1 4950
box -6 -8 66 268
use INVX1  _1307_
timestamp 0
transform 1 0 210 0 -1 4430
box -6 -8 66 268
use OAI21X1  _1308_
timestamp 0
transform 1 0 330 0 -1 4430
box -6 -8 106 268
use OAI21X1  _1309_
timestamp 0
transform 1 0 530 0 -1 3910
box -6 -8 106 268
use NAND2X1  _1310_
timestamp 0
transform 1 0 310 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1311_
timestamp 0
transform -1 0 170 0 1 4430
box -6 -8 106 268
use XOR2X1  _1312_
timestamp 0
transform -1 0 570 0 1 3910
box -6 -8 146 268
use NOR2X1  _1313_
timestamp 0
transform -1 0 150 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1314_
timestamp 0
transform -1 0 290 0 -1 3910
box -6 -8 86 268
use NAND2X1  _1315_
timestamp 0
transform -1 0 310 0 1 3390
box -6 -8 86 268
use OAI21X1  _1316_
timestamp 0
transform 1 0 70 0 1 3390
box -6 -8 106 268
use OAI21X1  _1317_
timestamp 0
transform -1 0 470 0 -1 3910
box -6 -8 106 268
use NOR2X1  _1318_
timestamp 0
transform -1 0 1290 0 1 3910
box -6 -8 86 268
use NAND2X1  _1319_
timestamp 0
transform 1 0 1250 0 -1 3910
box -6 -8 86 268
use INVX1  _1320_
timestamp 0
transform -1 0 1190 0 -1 3910
box -6 -8 66 268
use NOR2X1  _1321_
timestamp 0
transform -1 0 1010 0 1 3910
box -6 -8 86 268
use XNOR2X1  _1322_
timestamp 0
transform -1 0 370 0 1 3910
box -6 -8 146 268
use NAND2X1  _1323_
timestamp 0
transform 1 0 310 0 -1 2350
box -6 -8 86 268
use OAI21X1  _1324_
timestamp 0
transform -1 0 410 0 1 2350
box -6 -8 106 268
use NAND2X1  _1325_
timestamp 0
transform 1 0 1750 0 1 1310
box -6 -8 86 268
use OAI21X1  _1326_
timestamp 0
transform 1 0 230 0 1 4430
box -6 -8 106 268
use NAND2X1  _1327_
timestamp 0
transform 1 0 830 0 -1 3910
box -6 -8 86 268
use OAI21X1  _1328_
timestamp 0
transform 1 0 970 0 -1 3910
box -6 -8 106 268
use AND2X2  _1329_
timestamp 0
transform -1 0 170 0 1 3910
box -6 -8 106 268
use AOI21X1  _1330_
timestamp 0
transform 1 0 630 0 1 3910
box -6 -8 106 268
use NOR2X1  _1331_
timestamp 0
transform -1 0 150 0 -1 4430
box -6 -8 86 268
use NAND3X1  _1332_
timestamp 0
transform 1 0 650 0 -1 4430
box -6 -8 106 268
use NAND2X1  _1333_
timestamp 0
transform 1 0 790 0 1 3910
box -6 -8 86 268
use OR2X2  _1334_
timestamp 0
transform -1 0 2730 0 1 1310
box -6 -8 106 268
use NAND2X1  _1335_
timestamp 0
transform 1 0 2790 0 1 1310
box -6 -8 86 268
use AND2X2  _1336_
timestamp 0
transform -1 0 2570 0 1 1310
box -6 -8 106 268
use NOR2X1  _1337_
timestamp 0
transform -1 0 2290 0 1 1310
box -6 -8 86 268
use INVX1  _1338_
timestamp 0
transform 1 0 2210 0 -1 1830
box -6 -8 66 268
use INVX1  _1339_
timestamp 0
transform -1 0 2410 0 1 1310
box -6 -8 66 268
use OAI21X1  _1340_
timestamp 0
transform -1 0 2150 0 1 1310
box -6 -8 106 268
use OAI21X1  _1341_
timestamp 0
transform -1 0 1990 0 1 1310
box -6 -8 106 268
use OAI21X1  _1342_
timestamp 0
transform 1 0 2410 0 -1 1310
box -6 -8 106 268
use NOR2X1  _1343_
timestamp 0
transform 1 0 3490 0 -1 1310
box -6 -8 86 268
use NAND2X1  _1344_
timestamp 0
transform 1 0 3630 0 -1 1310
box -6 -8 86 268
use INVX1  _1345_
timestamp 0
transform 1 0 3010 0 -1 1310
box -6 -8 66 268
use NOR2X1  _1346_
timestamp 0
transform 1 0 2870 0 -1 1310
box -6 -8 86 268
use INVX1  _1347_
timestamp 0
transform -1 0 2630 0 -1 1310
box -6 -8 66 268
use XOR2X1  _1348_
timestamp 0
transform -1 0 2350 0 -1 1310
box -6 -8 146 268
use NAND2X1  _1349_
timestamp 0
transform -1 0 1450 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1350_
timestamp 0
transform -1 0 1850 0 -1 1310
box -6 -8 106 268
use NAND2X1  _1351_
timestamp 0
transform -1 0 550 0 1 790
box -6 -8 86 268
use NOR2X1  _1352_
timestamp 0
transform -1 0 2150 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1353_
timestamp 0
transform -1 0 2790 0 -1 1310
box -6 -8 106 268
use AOI21X1  _1354_
timestamp 0
transform -1 0 2010 0 -1 1310
box -6 -8 106 268
use NOR2X1  _1355_
timestamp 0
transform -1 0 1310 0 -1 790
box -6 -8 86 268
use NOR2X1  _1356_
timestamp 0
transform -1 0 1170 0 -1 790
box -6 -8 86 268
use NOR2X1  _1357_
timestamp 0
transform -1 0 890 0 -1 790
box -6 -8 86 268
use INVX1  _1358_
timestamp 0
transform 1 0 690 0 -1 790
box -6 -8 66 268
use AND2X2  _1359_
timestamp 0
transform 1 0 610 0 1 790
box -6 -8 106 268
use OAI21X1  _1360_
timestamp 0
transform 1 0 950 0 1 790
box -6 -8 106 268
use OAI21X1  _1361_
timestamp 0
transform -1 0 890 0 1 790
box -6 -8 106 268
use NOR2X1  _1362_
timestamp 0
transform -1 0 630 0 -1 790
box -6 -8 86 268
use NOR2X1  _1363_
timestamp 0
transform -1 0 350 0 -1 790
box -6 -8 86 268
use NOR2X1  _1364_
timestamp 0
transform 1 0 210 0 1 270
box -6 -8 86 268
use NAND2X1  _1365_
timestamp 0
transform 1 0 190 0 -1 270
box -6 -8 86 268
use INVX1  _1366_
timestamp 0
transform -1 0 130 0 -1 270
box -6 -8 66 268
use NOR2X1  _1367_
timestamp 0
transform -1 0 150 0 1 270
box -6 -8 86 268
use XOR2X1  _1368_
timestamp 0
transform -1 0 210 0 -1 790
box -6 -8 146 268
use NAND2X1  _1369_
timestamp 0
transform 1 0 230 0 -1 1310
box -6 -8 86 268
use OAI21X1  _1370_
timestamp 0
transform -1 0 170 0 -1 1310
box -6 -8 106 268
use NAND2X1  _1371_
timestamp 0
transform -1 0 2930 0 1 790
box -6 -8 86 268
use AOI21X1  _1372_
timestamp 0
transform 1 0 350 0 1 270
box -6 -8 106 268
use NAND2X1  _1373_
timestamp 0
transform -1 0 490 0 -1 790
box -6 -8 86 268
use OAI21X1  _1374_
timestamp 0
transform -1 0 610 0 1 270
box -6 -8 106 268
use NAND2X1  _1375_
timestamp 0
transform -1 0 4070 0 -1 790
box -6 -8 86 268
use NOR2X1  _1376_
timestamp 0
transform 1 0 4150 0 -1 790
box -6 -8 86 268
use INVX1  _1377_
timestamp 0
transform -1 0 3770 0 -1 790
box -6 -8 66 268
use AND2X2  _1378_
timestamp 0
transform 1 0 3830 0 -1 790
box -6 -8 106 268
use NOR2X1  _1379_
timestamp 0
transform -1 0 3070 0 -1 790
box -6 -8 86 268
use INVX1  _1380_
timestamp 0
transform -1 0 3230 0 1 270
box -6 -8 66 268
use INVX1  _1381_
timestamp 0
transform 1 0 3290 0 -1 790
box -6 -8 66 268
use OAI21X1  _1382_
timestamp 0
transform -1 0 3230 0 -1 790
box -6 -8 106 268
use OAI21X1  _1383_
timestamp 0
transform -1 0 3090 0 1 790
box -6 -8 106 268
use OAI21X1  _1384_
timestamp 0
transform 1 0 3550 0 -1 790
box -6 -8 106 268
use NOR2X1  _1385_
timestamp 0
transform 1 0 4270 0 1 270
box -6 -8 86 268
use NOR2X1  _1386_
timestamp 0
transform -1 0 4090 0 1 270
box -6 -8 86 268
use NOR2X1  _1387_
timestamp 0
transform -1 0 3950 0 1 270
box -6 -8 86 268
use INVX1  _1388_
timestamp 0
transform 1 0 3910 0 1 790
box -6 -8 66 268
use OR2X2  _1389_
timestamp 0
transform -1 0 3670 0 1 790
box -6 -8 106 268
use AOI21X1  _1390_
timestamp 0
transform 1 0 3750 0 1 790
box -6 -8 106 268
use AOI22X1  _1391_
timestamp 0
transform 1 0 3390 0 1 790
box -6 -8 126 268
use AOI21X1  _1392_
timestamp 0
transform -1 0 3810 0 1 270
box -6 -8 106 268
use INVX1  _1393_
timestamp 0
transform -1 0 3650 0 1 270
box -6 -8 66 268
use NOR2X1  _1394_
timestamp 0
transform -1 0 3490 0 -1 790
box -6 -8 86 268
use AOI21X1  _1395_
timestamp 0
transform -1 0 3390 0 1 270
box -6 -8 106 268
use INVX1  _1396_
timestamp 0
transform -1 0 2670 0 1 270
box -6 -8 66 268
use NOR2X1  _1397_
timestamp 0
transform 1 0 2310 0 1 270
box -6 -8 86 268
use OAI21X1  _1398_
timestamp 0
transform 1 0 2730 0 1 270
box -6 -8 106 268
use OAI22X1  _1399_
timestamp 0
transform 1 0 2270 0 -1 790
box -6 -8 126 268
use NAND2X1  _1400_
timestamp 0
transform -1 0 1850 0 1 790
box -6 -8 86 268
use NAND3X1  _1401_
timestamp 0
transform -1 0 2250 0 1 270
box -6 -8 106 268
use OAI21X1  _1402_
timestamp 0
transform -1 0 2550 0 1 270
box -6 -8 106 268
use NAND2X1  _1403_
timestamp 0
transform -1 0 2090 0 1 270
box -6 -8 86 268
use OAI21X1  _1404_
timestamp 0
transform -1 0 2010 0 1 790
box -6 -8 106 268
use INVX1  _1405_
timestamp 0
transform -1 0 3530 0 1 270
box -6 -8 66 268
use NAND3X1  _1406_
timestamp 0
transform 1 0 1490 0 -1 1830
box -6 -8 106 268
use NAND2X1  _1407_
timestamp 0
transform 1 0 3530 0 -1 1830
box -6 -8 86 268
use OAI21X1  _1408_
timestamp 0
transform 1 0 3370 0 -1 1830
box -6 -8 106 268
use INVX1  _1409_
timestamp 0
transform 1 0 3370 0 -1 270
box -6 -8 66 268
use NAND2X1  _1410_
timestamp 0
transform -1 0 3730 0 -1 270
box -6 -8 86 268
use OAI21X1  _1411_
timestamp 0
transform 1 0 3490 0 -1 270
box -6 -8 106 268
use INVX1  _1412_
timestamp 0
transform 1 0 2890 0 1 270
box -6 -8 66 268
use NAND2X1  _1413_
timestamp 0
transform 1 0 2990 0 -1 270
box -6 -8 86 268
use OAI21X1  _1414_
timestamp 0
transform 1 0 3010 0 1 270
box -6 -8 106 268
use INVX1  _1415_
timestamp 0
transform 1 0 1890 0 1 270
box -6 -8 66 268
use NAND2X1  _1416_
timestamp 0
transform -1 0 1610 0 -1 270
box -6 -8 86 268
use OAI21X1  _1417_
timestamp 0
transform 1 0 1490 0 1 270
box -6 -8 106 268
use NOR2X1  _1418_
timestamp 0
transform -1 0 970 0 1 1310
box -6 -8 86 268
use NOR2X1  _1419_
timestamp 0
transform 1 0 3130 0 1 2350
box -6 -8 86 268
use AOI21X1  _1420_
timestamp 0
transform 1 0 3290 0 1 2350
box -6 -8 106 268
use NOR2X1  _1421_
timestamp 0
transform -1 0 3130 0 1 1830
box -6 -8 86 268
use AOI21X1  _1422_
timestamp 0
transform 1 0 3190 0 1 1830
box -6 -8 106 268
use NOR2X1  _1423_
timestamp 0
transform -1 0 2530 0 -1 790
box -6 -8 86 268
use AOI21X1  _1424_
timestamp 0
transform -1 0 2930 0 -1 790
box -6 -8 106 268
use NOR2X1  _1425_
timestamp 0
transform 1 0 1190 0 1 270
box -6 -8 86 268
use AOI21X1  _1426_
timestamp 0
transform -1 0 1430 0 1 270
box -6 -8 106 268
use INVX1  _1427_
timestamp 0
transform 1 0 1930 0 1 3390
box -6 -8 66 268
use OAI21X1  _1428_
timestamp 0
transform -1 0 2290 0 1 2870
box -6 -8 106 268
use OAI21X1  _1429_
timestamp 0
transform -1 0 2450 0 1 2870
box -6 -8 106 268
use OAI21X1  _1430_
timestamp 0
transform 1 0 2430 0 -1 2870
box -6 -8 106 268
use OAI21X1  _1431_
timestamp 0
transform -1 0 2850 0 -1 2870
box -6 -8 106 268
use OAI21X1  _1432_
timestamp 0
transform 1 0 2110 0 -1 3390
box -6 -8 106 268
use OAI21X1  _1433_
timestamp 0
transform -1 0 2370 0 -1 3390
box -6 -8 106 268
use OAI21X1  _1434_
timestamp 0
transform -1 0 2370 0 -1 2870
box -6 -8 106 268
use OAI21X1  _1435_
timestamp 0
transform 1 0 2090 0 -1 2870
box -6 -8 106 268
use NOR2X1  _1436_
timestamp 0
transform -1 0 2310 0 1 1830
box -6 -8 86 268
use AOI21X1  _1437_
timestamp 0
transform -1 0 2710 0 1 1830
box -6 -8 106 268
use NOR2X1  _1438_
timestamp 0
transform -1 0 2650 0 -1 2350
box -6 -8 86 268
use AOI21X1  _1439_
timestamp 0
transform -1 0 2810 0 -1 2350
box -6 -8 106 268
use NOR2X1  _1440_
timestamp 0
transform -1 0 2590 0 1 2870
box -6 -8 86 268
use AOI21X1  _1441_
timestamp 0
transform 1 0 2590 0 -1 2870
box -6 -8 106 268
use NOR2X1  _1442_
timestamp 0
transform -1 0 1590 0 -1 2350
box -6 -8 86 268
use AOI21X1  _1443_
timestamp 0
transform 1 0 1650 0 -1 2350
box -6 -8 106 268
use NAND2X1  _1444_
timestamp 0
transform -1 0 2750 0 -1 3390
box -6 -8 86 268
use OAI21X1  _1445_
timestamp 0
transform -1 0 2910 0 -1 3390
box -6 -8 106 268
use NAND2X1  _1446_
timestamp 0
transform -1 0 3190 0 -1 3910
box -6 -8 86 268
use OAI21X1  _1447_
timestamp 0
transform -1 0 3230 0 1 3910
box -6 -8 106 268
use NAND2X1  _1448_
timestamp 0
transform -1 0 3330 0 -1 3910
box -6 -8 86 268
use OAI21X1  _1449_
timestamp 0
transform -1 0 3650 0 1 3910
box -6 -8 106 268
use NAND2X1  _1450_
timestamp 0
transform -1 0 2510 0 1 3390
box -6 -8 86 268
use OAI21X1  _1451_
timestamp 0
transform -1 0 2790 0 1 3390
box -6 -8 106 268
use DFFPOSX1  _1452_
timestamp 0
transform -1 0 3210 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1453_
timestamp 0
transform 1 0 3630 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1454_
timestamp 0
transform 1 0 3070 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1455_
timestamp 0
transform 1 0 3470 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1456_
timestamp 0
transform 1 0 1890 0 -1 2350
box -6 -8 246 268
use DFFPOSX1  _1457_
timestamp 0
transform -1 0 1610 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1458_
timestamp 0
transform 1 0 870 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1459_
timestamp 0
transform 1 0 430 0 -1 5470
box -6 -8 246 268
use DFFPOSX1  _1460_
timestamp 0
transform -1 0 510 0 -1 5990
box -6 -8 246 268
use DFFPOSX1  _1461_
timestamp 0
transform -1 0 1110 0 -1 4430
box -6 -8 246 268
use DFFPOSX1  _1462_
timestamp 0
transform -1 0 750 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1463_
timestamp 0
transform -1 0 1570 0 -1 3910
box -6 -8 246 268
use DFFPOSX1  _1464_
timestamp 0
transform 1 0 2410 0 -1 1830
box -6 -8 246 268
use DFFPOSX1  _1465_
timestamp 0
transform 1 0 2870 0 1 1310
box -6 -8 246 268
use DFFPOSX1  _1466_
timestamp 0
transform -1 0 1550 0 1 790
box -6 -8 246 268
use DFFPOSX1  _1467_
timestamp 0
transform -1 0 1130 0 1 270
box -6 -8 246 268
use DFFPOSX1  _1468_
timestamp 0
transform -1 0 4330 0 1 790
box -6 -8 246 268
use DFFPOSX1  _1469_
timestamp 0
transform -1 0 4510 0 -1 270
box -6 -8 246 268
use DFFPOSX1  _1470_
timestamp 0
transform -1 0 2630 0 -1 270
box -6 -8 246 268
use DFFPOSX1  _1471_
timestamp 0
transform 1 0 1910 0 -1 270
box -6 -8 246 268
use DFFPOSX1  _1472_
timestamp 0
transform -1 0 2590 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1473_
timestamp 0
transform -1 0 1750 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1474_
timestamp 0
transform -1 0 1290 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1475_
timestamp 0
transform -1 0 1310 0 -1 4950
box -6 -8 246 268
use DFFPOSX1  _1476_
timestamp 0
transform -1 0 750 0 -1 5990
box -6 -8 246 268
use DFFPOSX1  _1477_
timestamp 0
transform -1 0 910 0 -1 4950
box -6 -8 246 268
use DFFPOSX1  _1478_
timestamp 0
transform -1 0 530 0 1 5470
box -6 -8 246 268
use DFFPOSX1  _1479_
timestamp 0
transform 1 0 1290 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1480_
timestamp 0
transform -1 0 3770 0 1 1310
box -6 -8 246 268
use DFFPOSX1  _1481_
timestamp 0
transform 1 0 3710 0 -1 1310
box -6 -8 246 268
use DFFPOSX1  _1482_
timestamp 0
transform -1 0 1690 0 -1 790
box -6 -8 246 268
use DFFPOSX1  _1483_
timestamp 0
transform -1 0 790 0 -1 270
box -6 -8 246 268
use DFFPOSX1  _1484_
timestamp 0
transform -1 0 4690 0 1 790
box -6 -8 246 268
use DFFPOSX1  _1485_
timestamp 0
transform -1 0 4590 0 -1 790
box -6 -8 246 268
use DFFPOSX1  _1486_
timestamp 0
transform -1 0 1270 0 -1 1830
box -6 -8 246 268
use DFFPOSX1  _1487_
timestamp 0
transform -1 0 870 0 1 1830
box -6 -8 246 268
use DFFPOSX1  _1488_
timestamp 0
transform -1 0 790 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1489_
timestamp 0
transform 1 0 10 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1490_
timestamp 0
transform 1 0 10 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1491_
timestamp 0
transform -1 0 770 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1492_
timestamp 0
transform 1 0 10 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1493_
timestamp 0
transform 1 0 10 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1494_
timestamp 0
transform -1 0 1690 0 1 1310
box -6 -8 246 268
use DFFPOSX1  _1495_
timestamp 0
transform -1 0 1690 0 -1 1310
box -6 -8 246 268
use DFFPOSX1  _1496_
timestamp 0
transform -1 0 870 0 -1 1310
box -6 -8 246 268
use DFFPOSX1  _1497_
timestamp 0
transform 1 0 10 0 1 1310
box -6 -8 246 268
use DFFPOSX1  _1498_
timestamp 0
transform -1 0 3330 0 1 790
box -6 -8 246 268
use DFFPOSX1  _1499_
timestamp 0
transform -1 0 3430 0 -1 1310
box -6 -8 246 268
use DFFPOSX1  _1500_
timestamp 0
transform -1 0 2210 0 -1 790
box -6 -8 246 268
use DFFPOSX1  _1501_
timestamp 0
transform -1 0 2250 0 1 790
box -6 -8 246 268
use DFFPOSX1  _1502_
timestamp 0
transform 1 0 3070 0 -1 1830
box -6 -8 246 268
use DFFPOSX1  _1503_
timestamp 0
transform 1 0 3730 0 -1 270
box -6 -8 246 268
use DFFPOSX1  _1504_
timestamp 0
transform -1 0 3310 0 -1 270
box -6 -8 246 268
use DFFPOSX1  _1505_
timestamp 0
transform -1 0 1830 0 1 270
box -6 -8 246 268
use DFFPOSX1  _1506_
timestamp 0
transform 1 0 2830 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1507_
timestamp 0
transform 1 0 3290 0 1 1830
box -6 -8 246 268
use DFFPOSX1  _1508_
timestamp 0
transform -1 0 2770 0 -1 790
box -6 -8 246 268
use DFFPOSX1  _1509_
timestamp 0
transform -1 0 1470 0 -1 270
box -6 -8 246 268
use DFFPOSX1  _1510_
timestamp 0
transform -1 0 2050 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1511_
timestamp 0
transform 1 0 2850 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1512_
timestamp 0
transform -1 0 2370 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1513_
timestamp 0
transform -1 0 2130 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1514_
timestamp 0
transform -1 0 2550 0 1 1830
box -6 -8 246 268
use DFFPOSX1  _1515_
timestamp 0
transform -1 0 2830 0 1 2350
box -6 -8 246 268
use DFFPOSX1  _1516_
timestamp 0
transform -1 0 2830 0 1 2870
box -6 -8 246 268
use DFFPOSX1  _1517_
timestamp 0
transform -1 0 1890 0 -1 2870
box -6 -8 246 268
use DFFPOSX1  _1518_
timestamp 0
transform -1 0 2610 0 -1 3390
box -6 -8 246 268
use DFFPOSX1  _1519_
timestamp 0
transform 1 0 3230 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1520_
timestamp 0
transform 1 0 3650 0 1 3910
box -6 -8 246 268
use DFFPOSX1  _1521_
timestamp 0
transform 1 0 2790 0 1 3390
box -6 -8 246 268
use DFFPOSX1  _1522_
timestamp 0
transform 1 0 10 0 -1 2350
box -6 -8 246 268
use DFFPOSX1  _1523_
timestamp 0
transform -1 0 1870 0 1 1830
box -6 -8 246 268
use DFFPOSX1  _1524_
timestamp 0
transform -1 0 1970 0 -1 1830
box -6 -8 246 268
use DFFPOSX1  _1525_
timestamp 0
transform 1 0 870 0 1 1830
box -6 -8 246 268
use DFFPOSX1  _1526_
timestamp 0
transform 1 0 1110 0 1 1830
box -6 -8 246 268
use BUFX2  _1527_
timestamp 0
transform 1 0 5550 0 1 270
box -6 -8 86 268
use BUFX2  _1528_
timestamp 0
transform 1 0 3650 0 -1 3390
box -6 -8 86 268
use BUFX2  _1529_
timestamp 0
transform 1 0 4550 0 1 3910
box -6 -8 86 268
use BUFX2  _1530_
timestamp 0
transform 1 0 5410 0 -1 4430
box -6 -8 86 268
use BUFX2  _1531_
timestamp 0
transform 1 0 5890 0 1 4430
box -6 -8 86 268
use BUFX2  _1532_
timestamp 0
transform 1 0 950 0 -1 790
box -6 -8 86 268
use BUFX2  _1533_
timestamp 0
transform -1 0 550 0 -1 270
box -6 -8 86 268
use BUFX2  _1534_
timestamp 0
transform -1 0 410 0 -1 270
box -6 -8 86 268
use BUFX2  _1535_
timestamp 0
transform -1 0 150 0 1 790
box -6 -8 86 268
use BUFX2  BUFX2_insert0
timestamp 0
transform -1 0 1150 0 1 3910
box -6 -8 86 268
use BUFX2  BUFX2_insert1
timestamp 0
transform 1 0 3010 0 -1 2350
box -6 -8 86 268
use BUFX2  BUFX2_insert2
timestamp 0
transform -1 0 1190 0 1 790
box -6 -8 86 268
use BUFX2  BUFX2_insert3
timestamp 0
transform -1 0 1090 0 1 4430
box -6 -8 86 268
use BUFX2  BUFX2_insert4
timestamp 0
transform 1 0 1650 0 1 3390
box -6 -8 86 268
use BUFX2  BUFX2_insert5
timestamp 0
transform -1 0 2390 0 1 790
box -6 -8 86 268
use BUFX2  BUFX2_insert6
timestamp 0
transform 1 0 2990 0 -1 1830
box -6 -8 86 268
use BUFX2  BUFX2_insert15
timestamp 0
transform -1 0 2790 0 -1 3910
box -6 -8 86 268
use BUFX2  BUFX2_insert16
timestamp 0
transform -1 0 2970 0 -1 4950
box -6 -8 86 268
use BUFX2  BUFX2_insert17
timestamp 0
transform -1 0 4070 0 -1 4430
box -6 -8 86 268
use BUFX2  BUFX2_insert18
timestamp 0
transform 1 0 4310 0 -1 3910
box -6 -8 86 268
use BUFX2  BUFX2_insert19
timestamp 0
transform -1 0 590 0 -1 1830
box -6 -8 86 268
use BUFX2  BUFX2_insert20
timestamp 0
transform 1 0 1130 0 1 2870
box -6 -8 86 268
use BUFX2  BUFX2_insert21
timestamp 0
transform -1 0 550 0 1 2870
box -6 -8 86 268
use BUFX2  BUFX2_insert22
timestamp 0
transform -1 0 930 0 1 2350
box -6 -8 86 268
use BUFX2  BUFX2_insert23
timestamp 0
transform 1 0 2330 0 -1 1830
box -6 -8 86 268
use BUFX2  BUFX2_insert24
timestamp 0
transform 1 0 2770 0 1 1830
box -6 -8 86 268
use BUFX2  BUFX2_insert25
timestamp 0
transform 1 0 3270 0 1 2870
box -6 -8 86 268
use BUFX2  BUFX2_insert26
timestamp 0
transform -1 0 3230 0 -1 2870
box -6 -8 86 268
use BUFX2  BUFX2_insert27
timestamp 0
transform -1 0 2950 0 -1 2350
box -6 -8 86 268
use BUFX2  BUFX2_insert28
timestamp 0
transform -1 0 2970 0 1 2870
box -6 -8 86 268
use BUFX2  BUFX2_insert29
timestamp 0
transform 1 0 1370 0 -1 2350
box -6 -8 86 268
use BUFX2  BUFX2_insert30
timestamp 0
transform 1 0 4690 0 1 3910
box -6 -8 86 268
use BUFX2  BUFX2_insert31
timestamp 0
transform -1 0 3070 0 1 3910
box -6 -8 86 268
use BUFX2  BUFX2_insert32
timestamp 0
transform 1 0 4670 0 1 3390
box -6 -8 86 268
use BUFX2  BUFX2_insert33
timestamp 0
transform -1 0 2930 0 1 3910
box -6 -8 86 268
use CLKBUF1  CLKBUF1_insert7
timestamp 0
transform 1 0 810 0 -1 5990
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert8
timestamp 0
transform -1 0 270 0 -1 1830
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert9
timestamp 0
transform 1 0 2310 0 -1 2350
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert10
timestamp 0
transform -1 0 270 0 1 1830
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert11
timestamp 0
transform 1 0 210 0 1 790
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert12
timestamp 0
transform 1 0 2330 0 -1 3910
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert13
timestamp 0
transform 1 0 1910 0 -1 3910
box -6 -8 206 268
use CLKBUF1  CLKBUF1_insert14
timestamp 0
transform 1 0 2590 0 1 790
box -6 -8 206 268
use FILL  FILL87450x23550
timestamp 0
transform -1 0 5850 0 -1 1830
box -6 -8 26 268
use FILL  FILL87450x50850
timestamp 0
transform 1 0 5830 0 1 3390
box -6 -8 26 268
use FILL  FILL87450x54750
timestamp 0
transform -1 0 5850 0 -1 3910
box -6 -8 26 268
use FILL  FILL87450x70350
timestamp 0
transform -1 0 5850 0 -1 4950
box -6 -8 26 268
use FILL  FILL87450x74250
timestamp 0
transform 1 0 5830 0 1 4950
box -6 -8 26 268
use FILL  FILL87450x82050
timestamp 0
transform 1 0 5830 0 1 5470
box -6 -8 26 268
use FILL  FILL87750x23550
timestamp 0
transform -1 0 5870 0 -1 1830
box -6 -8 26 268
use FILL  FILL87750x31350
timestamp 0
transform -1 0 5870 0 -1 2350
box -6 -8 26 268
use FILL  FILL87750x35250
timestamp 0
transform 1 0 5850 0 1 2350
box -6 -8 26 268
use FILL  FILL87750x50850
timestamp 0
transform 1 0 5850 0 1 3390
box -6 -8 26 268
use FILL  FILL87750x54750
timestamp 0
transform -1 0 5870 0 -1 3910
box -6 -8 26 268
use FILL  FILL87750x70350
timestamp 0
transform -1 0 5870 0 -1 4950
box -6 -8 26 268
use FILL  FILL87750x74250
timestamp 0
transform 1 0 5850 0 1 4950
box -6 -8 26 268
use FILL  FILL87750x82050
timestamp 0
transform 1 0 5850 0 1 5470
box -6 -8 26 268
use FILL  FILL88050x150
timestamp 0
transform -1 0 5890 0 -1 270
box -6 -8 26 268
use FILL  FILL88050x15750
timestamp 0
transform -1 0 5890 0 -1 1310
box -6 -8 26 268
use FILL  FILL88050x19650
timestamp 0
transform 1 0 5870 0 1 1310
box -6 -8 26 268
use FILL  FILL88050x23550
timestamp 0
transform -1 0 5890 0 -1 1830
box -6 -8 26 268
use FILL  FILL88050x31350
timestamp 0
transform -1 0 5890 0 -1 2350
box -6 -8 26 268
use FILL  FILL88050x35250
timestamp 0
transform 1 0 5870 0 1 2350
box -6 -8 26 268
use FILL  FILL88050x50850
timestamp 0
transform 1 0 5870 0 1 3390
box -6 -8 26 268
use FILL  FILL88050x54750
timestamp 0
transform -1 0 5890 0 -1 3910
box -6 -8 26 268
use FILL  FILL88050x70350
timestamp 0
transform -1 0 5890 0 -1 4950
box -6 -8 26 268
use FILL  FILL88050x74250
timestamp 0
transform 1 0 5870 0 1 4950
box -6 -8 26 268
use FILL  FILL88050x78150
timestamp 0
transform -1 0 5890 0 -1 5470
box -6 -8 26 268
use FILL  FILL88050x82050
timestamp 0
transform 1 0 5870 0 1 5470
box -6 -8 26 268
use FILL  FILL88350x150
timestamp 0
transform -1 0 5910 0 -1 270
box -6 -8 26 268
use FILL  FILL88350x15750
timestamp 0
transform -1 0 5910 0 -1 1310
box -6 -8 26 268
use FILL  FILL88350x19650
timestamp 0
transform 1 0 5890 0 1 1310
box -6 -8 26 268
use FILL  FILL88350x23550
timestamp 0
transform -1 0 5910 0 -1 1830
box -6 -8 26 268
use FILL  FILL88350x31350
timestamp 0
transform -1 0 5910 0 -1 2350
box -6 -8 26 268
use FILL  FILL88350x35250
timestamp 0
transform 1 0 5890 0 1 2350
box -6 -8 26 268
use FILL  FILL88350x50850
timestamp 0
transform 1 0 5890 0 1 3390
box -6 -8 26 268
use FILL  FILL88350x54750
timestamp 0
transform -1 0 5910 0 -1 3910
box -6 -8 26 268
use FILL  FILL88350x70350
timestamp 0
transform -1 0 5910 0 -1 4950
box -6 -8 26 268
use FILL  FILL88350x74250
timestamp 0
transform 1 0 5890 0 1 4950
box -6 -8 26 268
use FILL  FILL88350x78150
timestamp 0
transform -1 0 5910 0 -1 5470
box -6 -8 26 268
use FILL  FILL88350x82050
timestamp 0
transform 1 0 5890 0 1 5470
box -6 -8 26 268
use FILL  FILL88650x150
timestamp 0
transform -1 0 5930 0 -1 270
box -6 -8 26 268
use FILL  FILL88650x4050
timestamp 0
transform 1 0 5910 0 1 270
box -6 -8 26 268
use FILL  FILL88650x11850
timestamp 0
transform 1 0 5910 0 1 790
box -6 -8 26 268
use FILL  FILL88650x15750
timestamp 0
transform -1 0 5930 0 -1 1310
box -6 -8 26 268
use FILL  FILL88650x19650
timestamp 0
transform 1 0 5910 0 1 1310
box -6 -8 26 268
use FILL  FILL88650x23550
timestamp 0
transform -1 0 5930 0 -1 1830
box -6 -8 26 268
use FILL  FILL88650x31350
timestamp 0
transform -1 0 5930 0 -1 2350
box -6 -8 26 268
use FILL  FILL88650x35250
timestamp 0
transform 1 0 5910 0 1 2350
box -6 -8 26 268
use FILL  FILL88650x46950
timestamp 0
transform -1 0 5930 0 -1 3390
box -6 -8 26 268
use FILL  FILL88650x50850
timestamp 0
transform 1 0 5910 0 1 3390
box -6 -8 26 268
use FILL  FILL88650x54750
timestamp 0
transform -1 0 5930 0 -1 3910
box -6 -8 26 268
use FILL  FILL88650x70350
timestamp 0
transform -1 0 5930 0 -1 4950
box -6 -8 26 268
use FILL  FILL88650x74250
timestamp 0
transform 1 0 5910 0 1 4950
box -6 -8 26 268
use FILL  FILL88650x78150
timestamp 0
transform -1 0 5930 0 -1 5470
box -6 -8 26 268
use FILL  FILL88650x82050
timestamp 0
transform 1 0 5910 0 1 5470
box -6 -8 26 268
use FILL  FILL88950x150
timestamp 0
transform -1 0 5950 0 -1 270
box -6 -8 26 268
use FILL  FILL88950x4050
timestamp 0
transform 1 0 5930 0 1 270
box -6 -8 26 268
use FILL  FILL88950x11850
timestamp 0
transform 1 0 5930 0 1 790
box -6 -8 26 268
use FILL  FILL88950x15750
timestamp 0
transform -1 0 5950 0 -1 1310
box -6 -8 26 268
use FILL  FILL88950x19650
timestamp 0
transform 1 0 5930 0 1 1310
box -6 -8 26 268
use FILL  FILL88950x23550
timestamp 0
transform -1 0 5950 0 -1 1830
box -6 -8 26 268
use FILL  FILL88950x31350
timestamp 0
transform -1 0 5950 0 -1 2350
box -6 -8 26 268
use FILL  FILL88950x35250
timestamp 0
transform 1 0 5930 0 1 2350
box -6 -8 26 268
use FILL  FILL88950x46950
timestamp 0
transform -1 0 5950 0 -1 3390
box -6 -8 26 268
use FILL  FILL88950x50850
timestamp 0
transform 1 0 5930 0 1 3390
box -6 -8 26 268
use FILL  FILL88950x54750
timestamp 0
transform -1 0 5950 0 -1 3910
box -6 -8 26 268
use FILL  FILL88950x70350
timestamp 0
transform -1 0 5950 0 -1 4950
box -6 -8 26 268
use FILL  FILL88950x74250
timestamp 0
transform 1 0 5930 0 1 4950
box -6 -8 26 268
use FILL  FILL88950x78150
timestamp 0
transform -1 0 5950 0 -1 5470
box -6 -8 26 268
use FILL  FILL88950x82050
timestamp 0
transform 1 0 5930 0 1 5470
box -6 -8 26 268
use FILL  FILL89250x150
timestamp 0
transform -1 0 5970 0 -1 270
box -6 -8 26 268
use FILL  FILL89250x4050
timestamp 0
transform 1 0 5950 0 1 270
box -6 -8 26 268
use FILL  FILL89250x7950
timestamp 0
transform -1 0 5970 0 -1 790
box -6 -8 26 268
use FILL  FILL89250x11850
timestamp 0
transform 1 0 5950 0 1 790
box -6 -8 26 268
use FILL  FILL89250x15750
timestamp 0
transform -1 0 5970 0 -1 1310
box -6 -8 26 268
use FILL  FILL89250x19650
timestamp 0
transform 1 0 5950 0 1 1310
box -6 -8 26 268
use FILL  FILL89250x23550
timestamp 0
transform -1 0 5970 0 -1 1830
box -6 -8 26 268
use FILL  FILL89250x27450
timestamp 0
transform 1 0 5950 0 1 1830
box -6 -8 26 268
use FILL  FILL89250x31350
timestamp 0
transform -1 0 5970 0 -1 2350
box -6 -8 26 268
use FILL  FILL89250x35250
timestamp 0
transform 1 0 5950 0 1 2350
box -6 -8 26 268
use FILL  FILL89250x46950
timestamp 0
transform -1 0 5970 0 -1 3390
box -6 -8 26 268
use FILL  FILL89250x50850
timestamp 0
transform 1 0 5950 0 1 3390
box -6 -8 26 268
use FILL  FILL89250x54750
timestamp 0
transform -1 0 5970 0 -1 3910
box -6 -8 26 268
use FILL  FILL89250x70350
timestamp 0
transform -1 0 5970 0 -1 4950
box -6 -8 26 268
use FILL  FILL89250x74250
timestamp 0
transform 1 0 5950 0 1 4950
box -6 -8 26 268
use FILL  FILL89250x78150
timestamp 0
transform -1 0 5970 0 -1 5470
box -6 -8 26 268
use FILL  FILL89250x82050
timestamp 0
transform 1 0 5950 0 1 5470
box -6 -8 26 268
use FILL  FILL89250x85950
timestamp 0
transform -1 0 5970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__723_
timestamp 0
transform 1 0 1130 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__724_
timestamp 0
transform -1 0 610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__725_
timestamp 0
transform -1 0 1610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__726_
timestamp 0
transform -1 0 1290 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__727_
timestamp 0
transform 1 0 1930 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__728_
timestamp 0
transform -1 0 2010 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__729_
timestamp 0
transform -1 0 730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__730_
timestamp 0
transform -1 0 990 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__731_
timestamp 0
transform 1 0 410 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__732_
timestamp 0
transform -1 0 3090 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__733_
timestamp 0
transform 1 0 1170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__734_
timestamp 0
transform -1 0 1030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__735_
timestamp 0
transform -1 0 470 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__736_
timestamp 0
transform -1 0 550 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__737_
timestamp 0
transform -1 0 1870 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__738_
timestamp 0
transform 1 0 870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__739_
timestamp 0
transform 1 0 470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__740_
timestamp 0
transform -1 0 410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__741_
timestamp 0
transform -1 0 330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__742_
timestamp 0
transform 1 0 690 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__743_
timestamp 0
transform -1 0 290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__744_
timestamp 0
transform -1 0 290 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__745_
timestamp 0
transform -1 0 270 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__746_
timestamp 0
transform 1 0 3470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__747_
timestamp 0
transform -1 0 3190 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__748_
timestamp 0
transform 1 0 3310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__749_
timestamp 0
transform 1 0 3870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__750_
timestamp 0
transform -1 0 3910 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__751_
timestamp 0
transform -1 0 4050 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__752_
timestamp 0
transform 1 0 3990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__753_
timestamp 0
transform -1 0 4210 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__754_
timestamp 0
transform 1 0 4330 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__755_
timestamp 0
transform -1 0 3630 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__756_
timestamp 0
transform -1 0 4330 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__757_
timestamp 0
transform 1 0 4450 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__758_
timestamp 0
transform 1 0 3230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__759_
timestamp 0
transform -1 0 3390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__760_
timestamp 0
transform 1 0 3330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__761_
timestamp 0
transform -1 0 3490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__762_
timestamp 0
transform 1 0 2910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__763_
timestamp 0
transform -1 0 2930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__764_
timestamp 0
transform 1 0 3030 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__765_
timestamp 0
transform -1 0 3330 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__766_
timestamp 0
transform 1 0 2130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__767_
timestamp 0
transform -1 0 2050 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__768_
timestamp 0
transform 1 0 1870 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__769_
timestamp 0
transform -1 0 1550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__770_
timestamp 0
transform 1 0 1770 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__771_
timestamp 0
transform 1 0 1610 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__772_
timestamp 0
transform -1 0 970 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__773_
timestamp 0
transform 1 0 1750 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__774_
timestamp 0
transform -1 0 1230 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__775_
timestamp 0
transform 1 0 670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__776_
timestamp 0
transform 1 0 1370 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__777_
timestamp 0
transform 1 0 790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__778_
timestamp 0
transform -1 0 30 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__779_
timestamp 0
transform 1 0 1710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__780_
timestamp 0
transform -1 0 290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__781_
timestamp 0
transform -1 0 770 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__782_
timestamp 0
transform 1 0 1890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__783_
timestamp 0
transform 1 0 1110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__784_
timestamp 0
transform 1 0 630 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__785_
timestamp 0
transform 1 0 910 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__786_
timestamp 0
transform 1 0 750 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__787_
timestamp 0
transform 1 0 1290 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__788_
timestamp 0
transform 1 0 1730 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__789_
timestamp 0
transform 1 0 1410 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__790_
timestamp 0
transform 1 0 2650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__791_
timestamp 0
transform 1 0 2850 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__792_
timestamp 0
transform 1 0 2770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__793_
timestamp 0
transform 1 0 3110 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__794_
timestamp 0
transform 1 0 3390 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__795_
timestamp 0
transform 1 0 3230 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__796_
timestamp 0
transform -1 0 1210 0 1 790
box -6 -8 26 268
use FILL  FILL_0__797_
timestamp 0
transform 1 0 2390 0 1 790
box -6 -8 26 268
use FILL  FILL_0__798_
timestamp 0
transform 1 0 1550 0 1 790
box -6 -8 26 268
use FILL  FILL_0__799_
timestamp 0
transform 1 0 790 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__800_
timestamp 0
transform 1 0 1090 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__801_
timestamp 0
transform 1 0 930 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__802_
timestamp 0
transform -1 0 3990 0 1 790
box -6 -8 26 268
use FILL  FILL_0__803_
timestamp 0
transform -1 0 3630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__804_
timestamp 0
transform -1 0 3970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__805_
timestamp 0
transform -1 0 4110 0 1 270
box -6 -8 26 268
use FILL  FILL_0__806_
timestamp 0
transform -1 0 3990 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__807_
timestamp 0
transform 1 0 4110 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__808_
timestamp 0
transform -1 0 2290 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__809_
timestamp 0
transform 1 0 2790 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__810_
timestamp 0
transform 1 0 2630 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__811_
timestamp 0
transform 1 0 2150 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__812_
timestamp 0
transform -1 0 1630 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__813_
timestamp 0
transform -1 0 1770 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__814_
timestamp 0
transform -1 0 2070 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__815_
timestamp 0
transform 1 0 2110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__816_
timestamp 0
transform 1 0 2190 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__817_
timestamp 0
transform 1 0 1970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__818_
timestamp 0
transform 1 0 2330 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__819_
timestamp 0
transform -1 0 2050 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__820_
timestamp 0
transform 1 0 1690 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__821_
timestamp 0
transform 1 0 1510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__822_
timestamp 0
transform -1 0 1670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__823_
timestamp 0
transform 1 0 1890 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__824_
timestamp 0
transform -1 0 1870 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__825_
timestamp 0
transform 1 0 2650 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__826_
timestamp 0
transform 1 0 2050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__827_
timestamp 0
transform 1 0 2470 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__828_
timestamp 0
transform -1 0 1890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__829_
timestamp 0
transform -1 0 1110 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__830_
timestamp 0
transform -1 0 2190 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__831_
timestamp 0
transform -1 0 2350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__832_
timestamp 0
transform 1 0 2190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__833_
timestamp 0
transform -1 0 3150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__834_
timestamp 0
transform -1 0 2670 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__835_
timestamp 0
transform -1 0 2490 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__836_
timestamp 0
transform -1 0 2630 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__837_
timestamp 0
transform -1 0 1230 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__838_
timestamp 0
transform 1 0 1710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__839_
timestamp 0
transform -1 0 1290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__840_
timestamp 0
transform -1 0 1570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__841_
timestamp 0
transform -1 0 1410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__842_
timestamp 0
transform 1 0 1070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__843_
timestamp 0
transform 1 0 1190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__844_
timestamp 0
transform -1 0 1370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__845_
timestamp 0
transform 1 0 990 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__846_
timestamp 0
transform 1 0 3390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__847_
timestamp 0
transform 1 0 1370 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__848_
timestamp 0
transform 1 0 2110 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__849_
timestamp 0
transform 1 0 2690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__850_
timestamp 0
transform 1 0 2550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__851_
timestamp 0
transform -1 0 2310 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__852_
timestamp 0
transform 1 0 2390 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__853_
timestamp 0
transform 1 0 2110 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__854_
timestamp 0
transform -1 0 2150 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__855_
timestamp 0
transform -1 0 2010 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__856_
timestamp 0
transform -1 0 2270 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__857_
timestamp 0
transform -1 0 1970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__858_
timestamp 0
transform -1 0 1630 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__859_
timestamp 0
transform -1 0 1550 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__860_
timestamp 0
transform -1 0 1810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__861_
timestamp 0
transform -1 0 3670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__862_
timestamp 0
transform -1 0 2950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__863_
timestamp 0
transform -1 0 2530 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__864_
timestamp 0
transform -1 0 2550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__865_
timestamp 0
transform -1 0 2510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__866_
timestamp 0
transform -1 0 1710 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__867_
timestamp 0
transform 1 0 1630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__868_
timestamp 0
transform -1 0 1470 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__869_
timestamp 0
transform -1 0 1530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__870_
timestamp 0
transform 1 0 1950 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__871_
timestamp 0
transform -1 0 1490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__872_
timestamp 0
transform -1 0 1350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__873_
timestamp 0
transform -1 0 1330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__874_
timestamp 0
transform -1 0 1310 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__875_
timestamp 0
transform -1 0 1090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__876_
timestamp 0
transform 1 0 1110 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__877_
timestamp 0
transform 1 0 170 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__878_
timestamp 0
transform -1 0 970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__879_
timestamp 0
transform -1 0 1810 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__880_
timestamp 0
transform 1 0 1630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__881_
timestamp 0
transform -1 0 2390 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__882_
timestamp 0
transform 1 0 3230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__883_
timestamp 0
transform 1 0 2790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__884_
timestamp 0
transform -1 0 2790 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__885_
timestamp 0
transform -1 0 2290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__886_
timestamp 0
transform 1 0 2670 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__887_
timestamp 0
transform -1 0 2550 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__888_
timestamp 0
transform -1 0 2410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__889_
timestamp 0
transform -1 0 3110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__890_
timestamp 0
transform 1 0 2990 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__891_
timestamp 0
transform 1 0 2630 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__892_
timestamp 0
transform -1 0 2330 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__893_
timestamp 0
transform 1 0 2230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__894_
timestamp 0
transform -1 0 2130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__895_
timestamp 0
transform -1 0 2570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__896_
timestamp 0
transform 1 0 1950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__897_
timestamp 0
transform 1 0 3530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__898_
timestamp 0
transform -1 0 2810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__899_
timestamp 0
transform 1 0 3350 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__900_
timestamp 0
transform 1 0 3390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__901_
timestamp 0
transform 1 0 2950 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__902_
timestamp 0
transform -1 0 2990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__903_
timestamp 0
transform -1 0 2170 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__904_
timestamp 0
transform -1 0 1810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__905_
timestamp 0
transform 1 0 2470 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__906_
timestamp 0
transform -1 0 2130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__907_
timestamp 0
transform -1 0 1970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__908_
timestamp 0
transform -1 0 1690 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__909_
timestamp 0
transform -1 0 1230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__910_
timestamp 0
transform 1 0 1510 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__911_
timestamp 0
transform -1 0 1850 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__912_
timestamp 0
transform -1 0 1850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__913_
timestamp 0
transform -1 0 1690 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__914_
timestamp 0
transform -1 0 1210 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__915_
timestamp 0
transform 1 0 1350 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__916_
timestamp 0
transform 1 0 1030 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__917_
timestamp 0
transform 1 0 710 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__918_
timestamp 0
transform -1 0 3830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__919_
timestamp 0
transform -1 0 2730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__920_
timestamp 0
transform 1 0 2710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__921_
timestamp 0
transform 1 0 1990 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__922_
timestamp 0
transform 1 0 3670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__923_
timestamp 0
transform -1 0 3310 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__924_
timestamp 0
transform 1 0 3130 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__925_
timestamp 0
transform 1 0 3530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__926_
timestamp 0
transform -1 0 3770 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__927_
timestamp 0
transform 1 0 3590 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__928_
timestamp 0
transform -1 0 3490 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__929_
timestamp 0
transform -1 0 3270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__930_
timestamp 0
transform 1 0 3130 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__931_
timestamp 0
transform 1 0 3290 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__932_
timestamp 0
transform -1 0 3350 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__933_
timestamp 0
transform -1 0 2830 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__934_
timestamp 0
transform -1 0 4230 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__935_
timestamp 0
transform 1 0 4910 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__936_
timestamp 0
transform -1 0 4090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__937_
timestamp 0
transform -1 0 4250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__938_
timestamp 0
transform -1 0 4570 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__939_
timestamp 0
transform -1 0 4630 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__940_
timestamp 0
transform 1 0 5050 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__941_
timestamp 0
transform -1 0 4410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__942_
timestamp 0
transform 1 0 4370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__943_
timestamp 0
transform -1 0 3790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__944_
timestamp 0
transform 1 0 4590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__945_
timestamp 0
transform -1 0 4110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__946_
timestamp 0
transform -1 0 4450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__947_
timestamp 0
transform 1 0 4770 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__948_
timestamp 0
transform -1 0 3790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__949_
timestamp 0
transform -1 0 3610 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__950_
timestamp 0
transform -1 0 3190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__951_
timestamp 0
transform -1 0 4290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__952_
timestamp 0
transform 1 0 3930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__953_
timestamp 0
transform -1 0 2870 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__954_
timestamp 0
transform -1 0 2970 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__955_
timestamp 0
transform 1 0 2390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__956_
timestamp 0
transform -1 0 3030 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__957_
timestamp 0
transform -1 0 3450 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__958_
timestamp 0
transform -1 0 3130 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__959_
timestamp 0
transform -1 0 2810 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__960_
timestamp 0
transform -1 0 2850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__961_
timestamp 0
transform 1 0 3270 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__962_
timestamp 0
transform -1 0 2570 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__963_
timestamp 0
transform -1 0 1370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__964_
timestamp 0
transform -1 0 1230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__965_
timestamp 0
transform 1 0 1010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__966_
timestamp 0
transform 1 0 810 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__967_
timestamp 0
transform -1 0 930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__968_
timestamp 0
transform 1 0 150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__969_
timestamp 0
transform -1 0 1510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__970_
timestamp 0
transform 1 0 3010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__971_
timestamp 0
transform 1 0 3170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__972_
timestamp 0
transform 1 0 3610 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__973_
timestamp 0
transform 1 0 3450 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__974_
timestamp 0
transform -1 0 5250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__975_
timestamp 0
transform -1 0 3490 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__976_
timestamp 0
transform 1 0 3610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__977_
timestamp 0
transform 1 0 3910 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__978_
timestamp 0
transform -1 0 4090 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__979_
timestamp 0
transform 1 0 3910 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__980_
timestamp 0
transform -1 0 4150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__981_
timestamp 0
transform 1 0 3970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__982_
timestamp 0
transform 1 0 4050 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__983_
timestamp 0
transform -1 0 4350 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__984_
timestamp 0
transform 1 0 4290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__985_
timestamp 0
transform 1 0 3750 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__986_
timestamp 0
transform 1 0 4450 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__987_
timestamp 0
transform -1 0 5090 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__988_
timestamp 0
transform 1 0 4230 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__989_
timestamp 0
transform -1 0 4390 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__990_
timestamp 0
transform 1 0 4770 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__991_
timestamp 0
transform -1 0 4570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__992_
timestamp 0
transform 1 0 4910 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__993_
timestamp 0
transform -1 0 5090 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__994_
timestamp 0
transform 1 0 4990 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__995_
timestamp 0
transform 1 0 5030 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__996_
timestamp 0
transform 1 0 5250 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__997_
timestamp 0
transform 1 0 4910 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__998_
timestamp 0
transform -1 0 4870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__999_
timestamp 0
transform 1 0 4690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1000_
timestamp 0
transform 1 0 5190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1001_
timestamp 0
transform -1 0 5050 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1002_
timestamp 0
transform -1 0 4530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1003_
timestamp 0
transform -1 0 4770 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1004_
timestamp 0
transform 1 0 4690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1005_
timestamp 0
transform -1 0 4890 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1006_
timestamp 0
transform -1 0 4730 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1007_
timestamp 0
transform -1 0 5190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1008_
timestamp 0
transform 1 0 5210 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1009_
timestamp 0
transform 1 0 5490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1010_
timestamp 0
transform 1 0 4870 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1011_
timestamp 0
transform -1 0 5250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1012_
timestamp 0
transform 1 0 4910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1013_
timestamp 0
transform 1 0 4430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1014_
timestamp 0
transform 1 0 4590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1015_
timestamp 0
transform 1 0 5390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1016_
timestamp 0
transform 1 0 5330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1017_
timestamp 0
transform -1 0 5090 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1018_
timestamp 0
transform -1 0 4930 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1019_
timestamp 0
transform -1 0 4870 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1020_
timestamp 0
transform -1 0 4770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1021_
timestamp 0
transform -1 0 4770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1022_
timestamp 0
transform 1 0 4450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1023_
timestamp 0
transform -1 0 3630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1024_
timestamp 0
transform 1 0 2230 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1025_
timestamp 0
transform -1 0 4310 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1026_
timestamp 0
transform 1 0 3330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1027_
timestamp 0
transform 1 0 3450 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1028_
timestamp 0
transform -1 0 4610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1029_
timestamp 0
transform 1 0 5070 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1030_
timestamp 0
transform -1 0 4150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1031_
timestamp 0
transform -1 0 3990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1032_
timestamp 0
transform 1 0 890 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1033_
timestamp 0
transform 1 0 530 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1034_
timestamp 0
transform 1 0 3810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1035_
timestamp 0
transform 1 0 5350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1036_
timestamp 0
transform 1 0 5470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1037_
timestamp 0
transform 1 0 4930 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1038_
timestamp 0
transform 1 0 5790 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1039_
timestamp 0
transform -1 0 5550 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1040_
timestamp 0
transform 1 0 5370 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1041_
timestamp 0
transform -1 0 4130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1042_
timestamp 0
transform 1 0 4150 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1043_
timestamp 0
transform 1 0 4030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1044_
timestamp 0
transform -1 0 3890 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1045_
timestamp 0
transform 1 0 3710 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1046_
timestamp 0
transform -1 0 4050 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1047_
timestamp 0
transform 1 0 4190 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1048_
timestamp 0
transform 1 0 4190 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1049_
timestamp 0
transform -1 0 3750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1050_
timestamp 0
transform -1 0 3890 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1051_
timestamp 0
transform 1 0 4330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1052_
timestamp 0
transform -1 0 5230 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1053_
timestamp 0
transform 1 0 5150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1054_
timestamp 0
transform -1 0 4950 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1055_
timestamp 0
transform -1 0 5090 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1056_
timestamp 0
transform 1 0 5310 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1057_
timestamp 0
transform 1 0 5130 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1058_
timestamp 0
transform -1 0 5610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1059_
timestamp 0
transform -1 0 5590 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1060_
timestamp 0
transform -1 0 4990 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1061_
timestamp 0
transform 1 0 5450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1062_
timestamp 0
transform 1 0 5690 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1063_
timestamp 0
transform 1 0 5750 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1064_
timestamp 0
transform 1 0 5670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1065_
timestamp 0
transform 1 0 5070 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1066_
timestamp 0
transform -1 0 5390 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1067_
timestamp 0
transform -1 0 5530 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1068_
timestamp 0
transform 1 0 4630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1069_
timestamp 0
transform 1 0 4750 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1070_
timestamp 0
transform 1 0 4810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1071_
timestamp 0
transform 1 0 5510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1072_
timestamp 0
transform 1 0 5530 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1073_
timestamp 0
transform 1 0 5350 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1074_
timestamp 0
transform 1 0 5630 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1075_
timestamp 0
transform -1 0 5370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1076_
timestamp 0
transform -1 0 5670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1077_
timestamp 0
transform 1 0 5670 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1078_
timestamp 0
transform 1 0 5190 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1079_
timestamp 0
transform 1 0 5670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1080_
timestamp 0
transform 1 0 5810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1081_
timestamp 0
transform 1 0 5490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1082_
timestamp 0
transform 1 0 5630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1083_
timestamp 0
transform -1 0 5670 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1084_
timestamp 0
transform 1 0 5670 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1085_
timestamp 0
transform -1 0 5730 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1086_
timestamp 0
transform -1 0 5570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1087_
timestamp 0
transform -1 0 5510 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1088_
timestamp 0
transform 1 0 5010 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1089_
timestamp 0
transform 1 0 5170 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1090_
timestamp 0
transform -1 0 5730 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1091_
timestamp 0
transform 1 0 5790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1092_
timestamp 0
transform 1 0 5330 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1093_
timestamp 0
transform 1 0 4550 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1094_
timestamp 0
transform -1 0 3770 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1095_
timestamp 0
transform 1 0 1570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1096_
timestamp 0
transform -1 0 1550 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1097_
timestamp 0
transform 1 0 3770 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1098_
timestamp 0
transform -1 0 4290 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1099_
timestamp 0
transform -1 0 4430 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1100_
timestamp 0
transform 1 0 4110 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1101_
timestamp 0
transform -1 0 5530 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1102_
timestamp 0
transform 1 0 5350 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1103_
timestamp 0
transform 1 0 4490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1104_
timestamp 0
transform 1 0 5830 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1105_
timestamp 0
transform -1 0 5870 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1106_
timestamp 0
transform -1 0 5710 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1107_
timestamp 0
transform -1 0 3770 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1108_
timestamp 0
transform 1 0 4130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1109_
timestamp 0
transform -1 0 4770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1110_
timestamp 0
transform -1 0 4330 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1111_
timestamp 0
transform 1 0 4410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1112_
timestamp 0
transform 1 0 4510 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1113_
timestamp 0
transform 1 0 5810 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1114_
timestamp 0
transform 1 0 5070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1115_
timestamp 0
transform 1 0 4790 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1116_
timestamp 0
transform -1 0 4510 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1117_
timestamp 0
transform 1 0 4630 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1118_
timestamp 0
transform -1 0 4930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1119_
timestamp 0
transform 1 0 5550 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1120_
timestamp 0
transform 1 0 5410 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1121_
timestamp 0
transform -1 0 5230 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1122_
timestamp 0
transform 1 0 5530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1123_
timestamp 0
transform 1 0 5530 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1124_
timestamp 0
transform 1 0 5030 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1125_
timestamp 0
transform -1 0 5390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1126_
timestamp 0
transform 1 0 5390 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1127_
timestamp 0
transform 1 0 5030 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1128_
timestamp 0
transform 1 0 5690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1129_
timestamp 0
transform 1 0 5550 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1130_
timestamp 0
transform 1 0 5670 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1131_
timestamp 0
transform 1 0 5210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1132_
timestamp 0
transform 1 0 5830 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1133_
timestamp 0
transform 1 0 5670 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1134_
timestamp 0
transform 1 0 5690 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1135_
timestamp 0
transform 1 0 5530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1136_
timestamp 0
transform 1 0 5750 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1137_
timestamp 0
transform -1 0 5650 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1138_
timestamp 0
transform -1 0 5390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1139_
timestamp 0
transform 1 0 5170 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1140_
timestamp 0
transform 1 0 5510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1141_
timestamp 0
transform 1 0 5330 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1142_
timestamp 0
transform 1 0 5470 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1143_
timestamp 0
transform -1 0 5690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1144_
timestamp 0
transform -1 0 5370 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1145_
timestamp 0
transform 1 0 5250 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1146_
timestamp 0
transform 1 0 4570 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1147_
timestamp 0
transform -1 0 3950 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1148_
timestamp 0
transform -1 0 5150 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1149_
timestamp 0
transform -1 0 4990 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1150_
timestamp 0
transform 1 0 4570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1151_
timestamp 0
transform 1 0 4390 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1152_
timestamp 0
transform -1 0 5250 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1153_
timestamp 0
transform -1 0 3110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1154_
timestamp 0
transform -1 0 3490 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1155_
timestamp 0
transform 1 0 3990 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1156_
timestamp 0
transform -1 0 3410 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1157_
timestamp 0
transform 1 0 3530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1158_
timestamp 0
transform 1 0 3230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1159_
timestamp 0
transform 1 0 4370 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1160_
timestamp 0
transform 1 0 4270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1161_
timestamp 0
transform -1 0 4230 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1162_
timestamp 0
transform 1 0 3550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1163_
timestamp 0
transform -1 0 3730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1164_
timestamp 0
transform -1 0 4750 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1165_
timestamp 0
transform 1 0 4890 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1166_
timestamp 0
transform -1 0 4250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1167_
timestamp 0
transform -1 0 4570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1168_
timestamp 0
transform -1 0 4890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1169_
timestamp 0
transform 1 0 4390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1170_
timestamp 0
transform -1 0 4290 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1171_
timestamp 0
transform 1 0 4670 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1172_
timestamp 0
transform 1 0 4510 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1173_
timestamp 0
transform 1 0 4710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1174_
timestamp 0
transform 1 0 4850 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1175_
timestamp 0
transform 1 0 5010 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1176_
timestamp 0
transform -1 0 5070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1177_
timestamp 0
transform 1 0 5190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1178_
timestamp 0
transform 1 0 5790 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1179_
timestamp 0
transform -1 0 5730 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1180_
timestamp 0
transform 1 0 5550 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1181_
timestamp 0
transform -1 0 5410 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1182_
timestamp 0
transform -1 0 4790 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1183_
timestamp 0
transform 1 0 4110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1184_
timestamp 0
transform -1 0 4270 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1185_
timestamp 0
transform -1 0 1330 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1186_
timestamp 0
transform 1 0 5450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1187_
timestamp 0
transform -1 0 5330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1188_
timestamp 0
transform 1 0 5730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1189_
timestamp 0
transform 1 0 5590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1190_
timestamp 0
transform -1 0 5650 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1191_
timestamp 0
transform 1 0 5150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1192_
timestamp 0
transform -1 0 4450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1193_
timestamp 0
transform -1 0 4090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1194_
timestamp 0
transform 1 0 5430 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1195_
timestamp 0
transform 1 0 5210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1196_
timestamp 0
transform -1 0 4030 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1197_
timestamp 0
transform -1 0 3850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1198_
timestamp 0
transform 1 0 3870 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1199_
timestamp 0
transform 1 0 3750 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1200_
timestamp 0
transform 1 0 3850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1201_
timestamp 0
transform -1 0 4590 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1202_
timestamp 0
transform 1 0 4730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1203_
timestamp 0
transform 1 0 5370 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1204_
timestamp 0
transform 1 0 5270 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1205_
timestamp 0
transform 1 0 5250 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1206_
timestamp 0
transform 1 0 5090 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1207_
timestamp 0
transform -1 0 5130 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1208_
timestamp 0
transform -1 0 4970 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1209_
timestamp 0
transform -1 0 4970 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1210_
timestamp 0
transform 1 0 4810 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1211_
timestamp 0
transform 1 0 4750 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1212_
timestamp 0
transform -1 0 4710 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1213_
timestamp 0
transform 1 0 3950 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1214_
timestamp 0
transform -1 0 4910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1215_
timestamp 0
transform 1 0 4090 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1216_
timestamp 0
transform -1 0 5370 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1217_
timestamp 0
transform 1 0 5190 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1218_
timestamp 0
transform -1 0 4610 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1219_
timestamp 0
transform 1 0 1690 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1220_
timestamp 0
transform 1 0 610 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1221_
timestamp 0
transform 1 0 5090 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1222_
timestamp 0
transform 1 0 4090 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1223_
timestamp 0
transform 1 0 3910 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1224_
timestamp 0
transform 1 0 3390 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1225_
timestamp 0
transform 1 0 3690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1226_
timestamp 0
transform -1 0 3710 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1227_
timestamp 0
transform 1 0 3810 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1228_
timestamp 0
transform -1 0 3550 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1229_
timestamp 0
transform -1 0 4230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1230_
timestamp 0
transform 1 0 4890 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1231_
timestamp 0
transform 1 0 4670 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1232_
timestamp 0
transform -1 0 4530 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1233_
timestamp 0
transform -1 0 4670 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1234_
timestamp 0
transform -1 0 4530 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1235_
timestamp 0
transform -1 0 4370 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1236_
timestamp 0
transform 1 0 750 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1237_
timestamp 0
transform -1 0 4350 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1238_
timestamp 0
transform 1 0 5690 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1239_
timestamp 0
transform 1 0 5250 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1240_
timestamp 0
transform -1 0 5430 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1241_
timestamp 0
transform 1 0 4790 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1242_
timestamp 0
transform 1 0 4870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1243_
timestamp 0
transform -1 0 3930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1244_
timestamp 0
transform 1 0 3570 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1245_
timestamp 0
transform -1 0 3770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1246_
timestamp 0
transform 1 0 3970 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1247_
timestamp 0
transform 1 0 4050 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1248_
timestamp 0
transform 1 0 4090 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1249_
timestamp 0
transform 1 0 4610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1250_
timestamp 0
transform 1 0 5030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1251_
timestamp 0
transform -1 0 5490 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1252_
timestamp 0
transform -1 0 5050 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1253_
timestamp 0
transform 1 0 4750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1254_
timestamp 0
transform 1 0 4870 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1255_
timestamp 0
transform 1 0 4690 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1256_
timestamp 0
transform -1 0 4250 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1257_
timestamp 0
transform -1 0 4430 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1258_
timestamp 0
transform 1 0 4250 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1259_
timestamp 0
transform 1 0 4410 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1260_
timestamp 0
transform 1 0 1750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1261_
timestamp 0
transform 1 0 1190 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1262_
timestamp 0
transform -1 0 1510 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1263_
timestamp 0
transform -1 0 1370 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1264_
timestamp 0
transform -1 0 910 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1265_
timestamp 0
transform -1 0 1290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1266_
timestamp 0
transform -1 0 1430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1267_
timestamp 0
transform -1 0 1290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1268_
timestamp 0
transform -1 0 1250 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1269_
timestamp 0
transform -1 0 950 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1270_
timestamp 0
transform -1 0 1070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1271_
timestamp 0
transform 1 0 1070 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1272_
timestamp 0
transform -1 0 930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1273_
timestamp 0
transform 1 0 590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1274_
timestamp 0
transform -1 0 770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1275_
timestamp 0
transform -1 0 1130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1276_
timestamp 0
transform -1 0 770 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1277_
timestamp 0
transform 1 0 550 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1278_
timestamp 0
transform -1 0 430 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1279_
timestamp 0
transform -1 0 570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1280_
timestamp 0
transform 1 0 930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1281_
timestamp 0
transform -1 0 790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1282_
timestamp 0
transform 1 0 710 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1283_
timestamp 0
transform 1 0 850 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1284_
timestamp 0
transform 1 0 570 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1285_
timestamp 0
transform -1 0 330 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1286_
timestamp 0
transform 1 0 250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1287_
timestamp 0
transform -1 0 270 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1288_
timestamp 0
transform 1 0 710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1289_
timestamp 0
transform 1 0 10 0 -1 5470
box -6 -8 26 268
use FILL  FILL_0__1290_
timestamp 0
transform 1 0 130 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0__1291_
timestamp 0
transform 1 0 10 0 1 5470
box -6 -8 26 268
use FILL  FILL_0__1292_
timestamp 0
transform -1 0 30 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1293_
timestamp 0
transform -1 0 570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1294_
timestamp 0
transform -1 0 410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1295_
timestamp 0
transform 1 0 150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1296_
timestamp 0
transform 1 0 10 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1297_
timestamp 0
transform 1 0 130 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1298_
timestamp 0
transform 1 0 430 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1299_
timestamp 0
transform 1 0 390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1300_
timestamp 0
transform -1 0 410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1301_
timestamp 0
transform 1 0 270 0 1 4950
box -6 -8 26 268
use FILL  FILL_0__1302_
timestamp 0
transform -1 0 510 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1303_
timestamp 0
transform 1 0 670 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1304_
timestamp 0
transform -1 0 350 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1305_
timestamp 0
transform -1 0 450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1306_
timestamp 0
transform -1 0 290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0__1307_
timestamp 0
transform 1 0 150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1308_
timestamp 0
transform 1 0 270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1309_
timestamp 0
transform 1 0 470 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1310_
timestamp 0
transform 1 0 250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1311_
timestamp 0
transform -1 0 30 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1312_
timestamp 0
transform -1 0 390 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1313_
timestamp 0
transform -1 0 30 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1314_
timestamp 0
transform -1 0 170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1315_
timestamp 0
transform -1 0 190 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1316_
timestamp 0
transform 1 0 10 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1317_
timestamp 0
transform -1 0 310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1318_
timestamp 0
transform -1 0 1170 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1319_
timestamp 0
transform 1 0 1190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1320_
timestamp 0
transform -1 0 1090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1321_
timestamp 0
transform -1 0 890 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1322_
timestamp 0
transform -1 0 190 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1323_
timestamp 0
transform 1 0 250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1324_
timestamp 0
transform -1 0 270 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1325_
timestamp 0
transform 1 0 1690 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1326_
timestamp 0
transform 1 0 170 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1327_
timestamp 0
transform 1 0 770 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1328_
timestamp 0
transform 1 0 910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1329_
timestamp 0
transform -1 0 30 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1330_
timestamp 0
transform 1 0 570 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1331_
timestamp 0
transform -1 0 30 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1332_
timestamp 0
transform 1 0 570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1333_
timestamp 0
transform 1 0 730 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1334_
timestamp 0
transform -1 0 2590 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1335_
timestamp 0
transform 1 0 2730 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1336_
timestamp 0
transform -1 0 2430 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1337_
timestamp 0
transform -1 0 2170 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1338_
timestamp 0
transform 1 0 2150 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1339_
timestamp 0
transform -1 0 2310 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1340_
timestamp 0
transform -1 0 2010 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1341_
timestamp 0
transform -1 0 1850 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1342_
timestamp 0
transform 1 0 2350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1343_
timestamp 0
transform 1 0 3430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1344_
timestamp 0
transform 1 0 3570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1345_
timestamp 0
transform 1 0 2950 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1346_
timestamp 0
transform 1 0 2790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1347_
timestamp 0
transform -1 0 2530 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1348_
timestamp 0
transform -1 0 2170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1349_
timestamp 0
transform -1 0 1330 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1350_
timestamp 0
transform -1 0 1710 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1351_
timestamp 0
transform -1 0 430 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1352_
timestamp 0
transform -1 0 2030 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1353_
timestamp 0
transform -1 0 2650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1354_
timestamp 0
transform -1 0 1870 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1355_
timestamp 0
transform -1 0 1190 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1356_
timestamp 0
transform -1 0 1050 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1357_
timestamp 0
transform -1 0 770 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1358_
timestamp 0
transform 1 0 630 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1359_
timestamp 0
transform 1 0 550 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1360_
timestamp 0
transform 1 0 890 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1361_
timestamp 0
transform -1 0 730 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1362_
timestamp 0
transform -1 0 510 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1363_
timestamp 0
transform -1 0 230 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1364_
timestamp 0
transform 1 0 150 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1365_
timestamp 0
transform 1 0 130 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1366_
timestamp 0
transform -1 0 30 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1367_
timestamp 0
transform -1 0 30 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1368_
timestamp 0
transform -1 0 30 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1369_
timestamp 0
transform 1 0 170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1370_
timestamp 0
transform -1 0 30 0 -1 1310
box -6 -8 26 268
use FILL  FILL_0__1371_
timestamp 0
transform -1 0 2810 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1372_
timestamp 0
transform 1 0 290 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1373_
timestamp 0
transform -1 0 370 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1374_
timestamp 0
transform -1 0 470 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1375_
timestamp 0
transform -1 0 3950 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1376_
timestamp 0
transform 1 0 4070 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1377_
timestamp 0
transform -1 0 3670 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1378_
timestamp 0
transform 1 0 3770 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1379_
timestamp 0
transform -1 0 2950 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1380_
timestamp 0
transform -1 0 3130 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1381_
timestamp 0
transform 1 0 3230 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1382_
timestamp 0
transform -1 0 3090 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1383_
timestamp 0
transform -1 0 2950 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1384_
timestamp 0
transform 1 0 3490 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1385_
timestamp 0
transform 1 0 4210 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1386_
timestamp 0
transform -1 0 3970 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1387_
timestamp 0
transform -1 0 3830 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1388_
timestamp 0
transform 1 0 3850 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1389_
timestamp 0
transform -1 0 3530 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1390_
timestamp 0
transform 1 0 3670 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1391_
timestamp 0
transform 1 0 3330 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1392_
timestamp 0
transform -1 0 3670 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1393_
timestamp 0
transform -1 0 3550 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1394_
timestamp 0
transform -1 0 3370 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1395_
timestamp 0
transform -1 0 3250 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1396_
timestamp 0
transform -1 0 2570 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1397_
timestamp 0
transform 1 0 2250 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1398_
timestamp 0
transform 1 0 2670 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1399_
timestamp 0
transform 1 0 2210 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1400_
timestamp 0
transform -1 0 1730 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1401_
timestamp 0
transform -1 0 2110 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1402_
timestamp 0
transform -1 0 2410 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1403_
timestamp 0
transform -1 0 1970 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1404_
timestamp 0
transform -1 0 1870 0 1 790
box -6 -8 26 268
use FILL  FILL_0__1405_
timestamp 0
transform -1 0 3410 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1406_
timestamp 0
transform 1 0 1430 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1407_
timestamp 0
transform 1 0 3470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1408_
timestamp 0
transform 1 0 3310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0__1409_
timestamp 0
transform 1 0 3310 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1410_
timestamp 0
transform -1 0 3610 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1411_
timestamp 0
transform 1 0 3430 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1412_
timestamp 0
transform 1 0 2830 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1413_
timestamp 0
transform 1 0 2930 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1414_
timestamp 0
transform 1 0 2950 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1415_
timestamp 0
transform 1 0 1830 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1416_
timestamp 0
transform -1 0 1490 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1417_
timestamp 0
transform 1 0 1430 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1418_
timestamp 0
transform -1 0 850 0 1 1310
box -6 -8 26 268
use FILL  FILL_0__1419_
timestamp 0
transform 1 0 3070 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1420_
timestamp 0
transform 1 0 3210 0 1 2350
box -6 -8 26 268
use FILL  FILL_0__1421_
timestamp 0
transform -1 0 3010 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1422_
timestamp 0
transform 1 0 3130 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1423_
timestamp 0
transform -1 0 2410 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1424_
timestamp 0
transform -1 0 2790 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1425_
timestamp 0
transform 1 0 1130 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1426_
timestamp 0
transform -1 0 1290 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1427_
timestamp 0
transform 1 0 1870 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1428_
timestamp 0
transform -1 0 2150 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1429_
timestamp 0
transform -1 0 2310 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1430_
timestamp 0
transform 1 0 2370 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1431_
timestamp 0
transform -1 0 2710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1432_
timestamp 0
transform 1 0 2050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1433_
timestamp 0
transform -1 0 2230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1434_
timestamp 0
transform -1 0 2210 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1435_
timestamp 0
transform 1 0 2030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1436_
timestamp 0
transform -1 0 2190 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1437_
timestamp 0
transform -1 0 2570 0 1 1830
box -6 -8 26 268
use FILL  FILL_0__1438_
timestamp 0
transform -1 0 2530 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1439_
timestamp 0
transform -1 0 2670 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1440_
timestamp 0
transform -1 0 2470 0 1 2870
box -6 -8 26 268
use FILL  FILL_0__1441_
timestamp 0
transform 1 0 2530 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0__1442_
timestamp 0
transform -1 0 1470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1443_
timestamp 0
transform 1 0 1590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0__1444_
timestamp 0
transform -1 0 2630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1445_
timestamp 0
transform -1 0 2770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1446_
timestamp 0
transform -1 0 3070 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1447_
timestamp 0
transform -1 0 3090 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1448_
timestamp 0
transform -1 0 3210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0__1449_
timestamp 0
transform -1 0 3490 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1450_
timestamp 0
transform -1 0 2390 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1451_
timestamp 0
transform -1 0 2650 0 1 3390
box -6 -8 26 268
use FILL  FILL_0__1527_
timestamp 0
transform 1 0 5490 0 1 270
box -6 -8 26 268
use FILL  FILL_0__1528_
timestamp 0
transform 1 0 3590 0 -1 3390
box -6 -8 26 268
use FILL  FILL_0__1529_
timestamp 0
transform 1 0 4490 0 1 3910
box -6 -8 26 268
use FILL  FILL_0__1530_
timestamp 0
transform 1 0 5350 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0__1531_
timestamp 0
transform 1 0 5830 0 1 4430
box -6 -8 26 268
use FILL  FILL_0__1532_
timestamp 0
transform 1 0 890 0 -1 790
box -6 -8 26 268
use FILL  FILL_0__1533_
timestamp 0
transform -1 0 430 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1534_
timestamp 0
transform -1 0 290 0 -1 270
box -6 -8 26 268
use FILL  FILL_0__1535_
timestamp 0
transform -1 0 30 0 1 790
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert0
timestamp 0
transform -1 0 1030 0 1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert1
timestamp 0
transform 1 0 2950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert2
timestamp 0
transform -1 0 1070 0 1 790
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert3
timestamp 0
transform -1 0 970 0 1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert4
timestamp 0
transform 1 0 1570 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert5
timestamp 0
transform -1 0 2270 0 1 790
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert6
timestamp 0
transform 1 0 2930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert15
timestamp 0
transform -1 0 2670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert16
timestamp 0
transform -1 0 2850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert17
timestamp 0
transform -1 0 3950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert18
timestamp 0
transform 1 0 4250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert19
timestamp 0
transform -1 0 450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert20
timestamp 0
transform 1 0 1070 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert21
timestamp 0
transform -1 0 430 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert22
timestamp 0
transform -1 0 810 0 1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert23
timestamp 0
transform 1 0 2270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert24
timestamp 0
transform 1 0 2710 0 1 1830
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert25
timestamp 0
transform 1 0 3210 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert26
timestamp 0
transform -1 0 3110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert27
timestamp 0
transform -1 0 2830 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert28
timestamp 0
transform -1 0 2850 0 1 2870
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert29
timestamp 0
transform 1 0 1310 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert30
timestamp 0
transform 1 0 4630 0 1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert31
timestamp 0
transform -1 0 2950 0 1 3910
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert32
timestamp 0
transform 1 0 4610 0 1 3390
box -6 -8 26 268
use FILL  FILL_0_BUFX2_insert33
timestamp 0
transform -1 0 2790 0 1 3910
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert7
timestamp 0
transform 1 0 750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert8
timestamp 0
transform -1 0 30 0 -1 1830
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert9
timestamp 0
transform 1 0 2250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert10
timestamp 0
transform -1 0 30 0 1 1830
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert11
timestamp 0
transform 1 0 150 0 1 790
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert12
timestamp 0
transform 1 0 2270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert13
timestamp 0
transform 1 0 1850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_0_CLKBUF1_insert14
timestamp 0
transform 1 0 2530 0 1 790
box -6 -8 26 268
use FILL  FILL_1__723_
timestamp 0
transform 1 0 1150 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__724_
timestamp 0
transform -1 0 630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__725_
timestamp 0
transform -1 0 1630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__726_
timestamp 0
transform -1 0 1310 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__727_
timestamp 0
transform 1 0 1950 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__728_
timestamp 0
transform -1 0 2030 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__729_
timestamp 0
transform -1 0 750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__730_
timestamp 0
transform -1 0 1010 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__731_
timestamp 0
transform 1 0 430 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__732_
timestamp 0
transform -1 0 3110 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__733_
timestamp 0
transform 1 0 1190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__734_
timestamp 0
transform -1 0 1050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__735_
timestamp 0
transform -1 0 490 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__736_
timestamp 0
transform -1 0 570 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__737_
timestamp 0
transform -1 0 1890 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__738_
timestamp 0
transform 1 0 890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__739_
timestamp 0
transform 1 0 490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__740_
timestamp 0
transform -1 0 430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__741_
timestamp 0
transform -1 0 350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__742_
timestamp 0
transform 1 0 710 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__743_
timestamp 0
transform -1 0 310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__744_
timestamp 0
transform -1 0 310 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__745_
timestamp 0
transform -1 0 290 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__746_
timestamp 0
transform 1 0 3490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__747_
timestamp 0
transform -1 0 3210 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__748_
timestamp 0
transform 1 0 3330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__749_
timestamp 0
transform 1 0 3890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__750_
timestamp 0
transform -1 0 3930 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__751_
timestamp 0
transform -1 0 4070 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__752_
timestamp 0
transform 1 0 4010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__753_
timestamp 0
transform -1 0 4230 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__754_
timestamp 0
transform 1 0 4350 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__755_
timestamp 0
transform -1 0 3650 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__756_
timestamp 0
transform -1 0 4350 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__757_
timestamp 0
transform 1 0 4470 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__758_
timestamp 0
transform 1 0 3250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__759_
timestamp 0
transform -1 0 3410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__760_
timestamp 0
transform 1 0 3350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__761_
timestamp 0
transform -1 0 3510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__762_
timestamp 0
transform 1 0 2930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__763_
timestamp 0
transform -1 0 2950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__764_
timestamp 0
transform 1 0 3050 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__765_
timestamp 0
transform -1 0 3350 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__766_
timestamp 0
transform 1 0 2150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__767_
timestamp 0
transform -1 0 2070 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__768_
timestamp 0
transform 1 0 1890 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__769_
timestamp 0
transform -1 0 1570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__770_
timestamp 0
transform 1 0 1790 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__771_
timestamp 0
transform 1 0 1630 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__772_
timestamp 0
transform -1 0 990 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__773_
timestamp 0
transform 1 0 1770 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__774_
timestamp 0
transform -1 0 1250 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__775_
timestamp 0
transform 1 0 690 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__776_
timestamp 0
transform 1 0 1390 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__777_
timestamp 0
transform 1 0 810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__778_
timestamp 0
transform -1 0 50 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__779_
timestamp 0
transform 1 0 1730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__780_
timestamp 0
transform -1 0 310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__781_
timestamp 0
transform -1 0 790 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__782_
timestamp 0
transform 1 0 1910 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__783_
timestamp 0
transform 1 0 1130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__784_
timestamp 0
transform 1 0 650 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__785_
timestamp 0
transform 1 0 930 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__786_
timestamp 0
transform 1 0 770 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__787_
timestamp 0
transform 1 0 1310 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__788_
timestamp 0
transform 1 0 1750 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__789_
timestamp 0
transform 1 0 1430 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__790_
timestamp 0
transform 1 0 2670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__791_
timestamp 0
transform 1 0 2870 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__792_
timestamp 0
transform 1 0 2790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__793_
timestamp 0
transform 1 0 3130 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__794_
timestamp 0
transform 1 0 3410 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__795_
timestamp 0
transform 1 0 3250 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__796_
timestamp 0
transform -1 0 1230 0 1 790
box -6 -8 26 268
use FILL  FILL_1__797_
timestamp 0
transform 1 0 2410 0 1 790
box -6 -8 26 268
use FILL  FILL_1__798_
timestamp 0
transform 1 0 1570 0 1 790
box -6 -8 26 268
use FILL  FILL_1__799_
timestamp 0
transform 1 0 810 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__800_
timestamp 0
transform 1 0 1110 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__801_
timestamp 0
transform 1 0 950 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__802_
timestamp 0
transform -1 0 4010 0 1 790
box -6 -8 26 268
use FILL  FILL_1__803_
timestamp 0
transform -1 0 3650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__804_
timestamp 0
transform -1 0 3990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__805_
timestamp 0
transform -1 0 4130 0 1 270
box -6 -8 26 268
use FILL  FILL_1__806_
timestamp 0
transform -1 0 4010 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__807_
timestamp 0
transform 1 0 4130 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__808_
timestamp 0
transform -1 0 2310 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__809_
timestamp 0
transform 1 0 2810 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__810_
timestamp 0
transform 1 0 2650 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__811_
timestamp 0
transform 1 0 2170 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__812_
timestamp 0
transform -1 0 1650 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__813_
timestamp 0
transform -1 0 1790 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__814_
timestamp 0
transform -1 0 2090 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__815_
timestamp 0
transform 1 0 2130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__816_
timestamp 0
transform 1 0 2210 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__817_
timestamp 0
transform 1 0 1990 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__818_
timestamp 0
transform 1 0 2350 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__819_
timestamp 0
transform -1 0 2070 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__820_
timestamp 0
transform 1 0 1710 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__821_
timestamp 0
transform 1 0 1530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__822_
timestamp 0
transform -1 0 1690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__823_
timestamp 0
transform 1 0 1910 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__824_
timestamp 0
transform -1 0 1890 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__825_
timestamp 0
transform 1 0 2670 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__826_
timestamp 0
transform 1 0 2070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__827_
timestamp 0
transform 1 0 2490 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__828_
timestamp 0
transform -1 0 1910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__829_
timestamp 0
transform -1 0 1130 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__830_
timestamp 0
transform -1 0 2210 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__831_
timestamp 0
transform -1 0 2370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__832_
timestamp 0
transform 1 0 2210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__833_
timestamp 0
transform -1 0 3170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__834_
timestamp 0
transform -1 0 2690 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__835_
timestamp 0
transform -1 0 2510 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__836_
timestamp 0
transform -1 0 2650 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__837_
timestamp 0
transform -1 0 1250 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__838_
timestamp 0
transform 1 0 1730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__839_
timestamp 0
transform -1 0 1310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__840_
timestamp 0
transform -1 0 1590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__841_
timestamp 0
transform -1 0 1430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__842_
timestamp 0
transform 1 0 1090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__843_
timestamp 0
transform 1 0 1210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__844_
timestamp 0
transform -1 0 1390 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__845_
timestamp 0
transform 1 0 1010 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__846_
timestamp 0
transform 1 0 3410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__847_
timestamp 0
transform 1 0 1390 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__848_
timestamp 0
transform 1 0 2130 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__849_
timestamp 0
transform 1 0 2710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__850_
timestamp 0
transform 1 0 2570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__851_
timestamp 0
transform -1 0 2330 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__852_
timestamp 0
transform 1 0 2410 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__853_
timestamp 0
transform 1 0 2130 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__854_
timestamp 0
transform -1 0 2170 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__855_
timestamp 0
transform -1 0 2030 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__856_
timestamp 0
transform -1 0 2290 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__857_
timestamp 0
transform -1 0 1990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__858_
timestamp 0
transform -1 0 1650 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__859_
timestamp 0
transform -1 0 1570 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__860_
timestamp 0
transform -1 0 1830 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__861_
timestamp 0
transform -1 0 3690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__862_
timestamp 0
transform -1 0 2970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__863_
timestamp 0
transform -1 0 2550 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__864_
timestamp 0
transform -1 0 2570 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__865_
timestamp 0
transform -1 0 2530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__866_
timestamp 0
transform -1 0 1730 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__867_
timestamp 0
transform 1 0 1650 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__868_
timestamp 0
transform -1 0 1490 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__869_
timestamp 0
transform -1 0 1550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__870_
timestamp 0
transform 1 0 1970 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__871_
timestamp 0
transform -1 0 1510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__872_
timestamp 0
transform -1 0 1370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__873_
timestamp 0
transform -1 0 1350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__874_
timestamp 0
transform -1 0 1330 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__875_
timestamp 0
transform -1 0 1110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__876_
timestamp 0
transform 1 0 1130 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__877_
timestamp 0
transform 1 0 190 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__878_
timestamp 0
transform -1 0 990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__879_
timestamp 0
transform -1 0 1830 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__880_
timestamp 0
transform 1 0 1650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__881_
timestamp 0
transform -1 0 2410 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__882_
timestamp 0
transform 1 0 3250 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__883_
timestamp 0
transform 1 0 2810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__884_
timestamp 0
transform -1 0 2810 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__885_
timestamp 0
transform -1 0 2310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__886_
timestamp 0
transform 1 0 2690 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__887_
timestamp 0
transform -1 0 2570 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__888_
timestamp 0
transform -1 0 2430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__889_
timestamp 0
transform -1 0 3130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__890_
timestamp 0
transform 1 0 3010 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__891_
timestamp 0
transform 1 0 2650 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__892_
timestamp 0
transform -1 0 2350 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__893_
timestamp 0
transform 1 0 2250 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__894_
timestamp 0
transform -1 0 2150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__895_
timestamp 0
transform -1 0 2590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__896_
timestamp 0
transform 1 0 1970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__897_
timestamp 0
transform 1 0 3550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__898_
timestamp 0
transform -1 0 2830 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__899_
timestamp 0
transform 1 0 3370 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__900_
timestamp 0
transform 1 0 3410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__901_
timestamp 0
transform 1 0 2970 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__902_
timestamp 0
transform -1 0 3010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__903_
timestamp 0
transform -1 0 2190 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__904_
timestamp 0
transform -1 0 1830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__905_
timestamp 0
transform 1 0 2490 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__906_
timestamp 0
transform -1 0 2150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__907_
timestamp 0
transform -1 0 1990 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__908_
timestamp 0
transform -1 0 1710 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__909_
timestamp 0
transform -1 0 1250 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__910_
timestamp 0
transform 1 0 1530 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__911_
timestamp 0
transform -1 0 1870 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__912_
timestamp 0
transform -1 0 1870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__913_
timestamp 0
transform -1 0 1710 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__914_
timestamp 0
transform -1 0 1230 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__915_
timestamp 0
transform 1 0 1370 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__916_
timestamp 0
transform 1 0 1050 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__917_
timestamp 0
transform 1 0 730 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__918_
timestamp 0
transform -1 0 3850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__919_
timestamp 0
transform -1 0 2750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__920_
timestamp 0
transform 1 0 2730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__921_
timestamp 0
transform 1 0 2010 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__922_
timestamp 0
transform 1 0 3690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__923_
timestamp 0
transform -1 0 3330 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__924_
timestamp 0
transform 1 0 3150 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__925_
timestamp 0
transform 1 0 3550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__926_
timestamp 0
transform -1 0 3790 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__927_
timestamp 0
transform 1 0 3610 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__928_
timestamp 0
transform -1 0 3510 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__929_
timestamp 0
transform -1 0 3290 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__930_
timestamp 0
transform 1 0 3150 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__931_
timestamp 0
transform 1 0 3310 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__932_
timestamp 0
transform -1 0 3370 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__933_
timestamp 0
transform -1 0 2850 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__934_
timestamp 0
transform -1 0 4250 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__935_
timestamp 0
transform 1 0 4930 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__936_
timestamp 0
transform -1 0 4110 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__937_
timestamp 0
transform -1 0 4270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__938_
timestamp 0
transform -1 0 4590 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__939_
timestamp 0
transform -1 0 4650 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__940_
timestamp 0
transform 1 0 5070 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__941_
timestamp 0
transform -1 0 4430 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__942_
timestamp 0
transform 1 0 4390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__943_
timestamp 0
transform -1 0 3810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__944_
timestamp 0
transform 1 0 4610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__945_
timestamp 0
transform -1 0 4130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__946_
timestamp 0
transform -1 0 4470 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__947_
timestamp 0
transform 1 0 4790 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__948_
timestamp 0
transform -1 0 3810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__949_
timestamp 0
transform -1 0 3630 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__950_
timestamp 0
transform -1 0 3210 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__951_
timestamp 0
transform -1 0 4310 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__952_
timestamp 0
transform 1 0 3950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__953_
timestamp 0
transform -1 0 2890 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__954_
timestamp 0
transform -1 0 2990 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__955_
timestamp 0
transform 1 0 2410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__956_
timestamp 0
transform -1 0 3050 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__957_
timestamp 0
transform -1 0 3470 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__958_
timestamp 0
transform -1 0 3150 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__959_
timestamp 0
transform -1 0 2830 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__960_
timestamp 0
transform -1 0 2870 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__961_
timestamp 0
transform 1 0 3290 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__962_
timestamp 0
transform -1 0 2590 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__963_
timestamp 0
transform -1 0 1390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__964_
timestamp 0
transform -1 0 1250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__965_
timestamp 0
transform 1 0 1030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__966_
timestamp 0
transform 1 0 830 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__967_
timestamp 0
transform -1 0 950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__968_
timestamp 0
transform 1 0 170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__969_
timestamp 0
transform -1 0 1530 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__970_
timestamp 0
transform 1 0 3030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__971_
timestamp 0
transform 1 0 3190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__972_
timestamp 0
transform 1 0 3630 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__973_
timestamp 0
transform 1 0 3470 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__974_
timestamp 0
transform -1 0 5270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__975_
timestamp 0
transform -1 0 3510 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__976_
timestamp 0
transform 1 0 3630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__977_
timestamp 0
transform 1 0 3930 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__978_
timestamp 0
transform -1 0 4110 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__979_
timestamp 0
transform 1 0 3930 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__980_
timestamp 0
transform -1 0 4170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__981_
timestamp 0
transform 1 0 3990 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__982_
timestamp 0
transform 1 0 4070 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__983_
timestamp 0
transform -1 0 4370 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__984_
timestamp 0
transform 1 0 4310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__985_
timestamp 0
transform 1 0 3770 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__986_
timestamp 0
transform 1 0 4470 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__987_
timestamp 0
transform -1 0 5110 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__988_
timestamp 0
transform 1 0 4250 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__989_
timestamp 0
transform -1 0 4410 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__990_
timestamp 0
transform 1 0 4790 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__991_
timestamp 0
transform -1 0 4590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__992_
timestamp 0
transform 1 0 4930 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__993_
timestamp 0
transform -1 0 5110 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__994_
timestamp 0
transform 1 0 5010 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__995_
timestamp 0
transform 1 0 5050 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__996_
timestamp 0
transform 1 0 5270 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__997_
timestamp 0
transform 1 0 4930 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__998_
timestamp 0
transform -1 0 4890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__999_
timestamp 0
transform 1 0 4710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1000_
timestamp 0
transform 1 0 5210 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1001_
timestamp 0
transform -1 0 5070 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1002_
timestamp 0
transform -1 0 4550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1003_
timestamp 0
transform -1 0 4790 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1004_
timestamp 0
transform 1 0 4710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1005_
timestamp 0
transform -1 0 4910 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1006_
timestamp 0
transform -1 0 4750 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1007_
timestamp 0
transform -1 0 5210 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1008_
timestamp 0
transform 1 0 5230 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1009_
timestamp 0
transform 1 0 5510 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1010_
timestamp 0
transform 1 0 4890 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1011_
timestamp 0
transform -1 0 5270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1012_
timestamp 0
transform 1 0 4930 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1013_
timestamp 0
transform 1 0 4450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1014_
timestamp 0
transform 1 0 4610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1015_
timestamp 0
transform 1 0 5410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1016_
timestamp 0
transform 1 0 5350 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1017_
timestamp 0
transform -1 0 5110 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1018_
timestamp 0
transform -1 0 4950 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1019_
timestamp 0
transform -1 0 4890 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1020_
timestamp 0
transform -1 0 4790 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1021_
timestamp 0
transform -1 0 4790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1022_
timestamp 0
transform 1 0 4470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1023_
timestamp 0
transform -1 0 3650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1024_
timestamp 0
transform 1 0 2250 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1025_
timestamp 0
transform -1 0 4330 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1026_
timestamp 0
transform 1 0 3350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1027_
timestamp 0
transform 1 0 3470 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1028_
timestamp 0
transform -1 0 4630 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1029_
timestamp 0
transform 1 0 5090 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1030_
timestamp 0
transform -1 0 4170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1031_
timestamp 0
transform -1 0 4010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1032_
timestamp 0
transform 1 0 910 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1033_
timestamp 0
transform 1 0 550 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1034_
timestamp 0
transform 1 0 3830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1035_
timestamp 0
transform 1 0 5370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1036_
timestamp 0
transform 1 0 5490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1037_
timestamp 0
transform 1 0 4950 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1038_
timestamp 0
transform 1 0 5810 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1039_
timestamp 0
transform -1 0 5570 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1040_
timestamp 0
transform 1 0 5390 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1041_
timestamp 0
transform -1 0 4150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1042_
timestamp 0
transform 1 0 4170 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1043_
timestamp 0
transform 1 0 4050 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1044_
timestamp 0
transform -1 0 3910 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1045_
timestamp 0
transform 1 0 3730 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1046_
timestamp 0
transform -1 0 4070 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1047_
timestamp 0
transform 1 0 4210 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1048_
timestamp 0
transform 1 0 4210 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1049_
timestamp 0
transform -1 0 3770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1050_
timestamp 0
transform -1 0 3910 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1051_
timestamp 0
transform 1 0 4350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1052_
timestamp 0
transform -1 0 5250 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1053_
timestamp 0
transform 1 0 5170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1054_
timestamp 0
transform -1 0 4970 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1055_
timestamp 0
transform -1 0 5110 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1056_
timestamp 0
transform 1 0 5330 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1057_
timestamp 0
transform 1 0 5150 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1058_
timestamp 0
transform -1 0 5630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1059_
timestamp 0
transform -1 0 5610 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1060_
timestamp 0
transform -1 0 5010 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1061_
timestamp 0
transform 1 0 5470 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1062_
timestamp 0
transform 1 0 5710 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1063_
timestamp 0
transform 1 0 5770 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1064_
timestamp 0
transform 1 0 5690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1065_
timestamp 0
transform 1 0 5090 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1066_
timestamp 0
transform -1 0 5410 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1067_
timestamp 0
transform -1 0 5550 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1068_
timestamp 0
transform 1 0 4650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1069_
timestamp 0
transform 1 0 4770 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1070_
timestamp 0
transform 1 0 4830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1071_
timestamp 0
transform 1 0 5530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1072_
timestamp 0
transform 1 0 5550 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1073_
timestamp 0
transform 1 0 5370 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1074_
timestamp 0
transform 1 0 5650 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1075_
timestamp 0
transform -1 0 5390 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1076_
timestamp 0
transform -1 0 5690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1077_
timestamp 0
transform 1 0 5690 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1078_
timestamp 0
transform 1 0 5210 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1079_
timestamp 0
transform 1 0 5690 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1080_
timestamp 0
transform 1 0 5830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1081_
timestamp 0
transform 1 0 5510 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1082_
timestamp 0
transform 1 0 5650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1083_
timestamp 0
transform -1 0 5690 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1084_
timestamp 0
transform 1 0 5690 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1085_
timestamp 0
transform -1 0 5750 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1086_
timestamp 0
transform -1 0 5590 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1087_
timestamp 0
transform -1 0 5530 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1088_
timestamp 0
transform 1 0 5030 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1089_
timestamp 0
transform 1 0 5190 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1090_
timestamp 0
transform -1 0 5750 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1091_
timestamp 0
transform 1 0 5810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1092_
timestamp 0
transform 1 0 5350 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1093_
timestamp 0
transform 1 0 4570 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1094_
timestamp 0
transform -1 0 3790 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1095_
timestamp 0
transform 1 0 1590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1096_
timestamp 0
transform -1 0 1570 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1097_
timestamp 0
transform 1 0 3790 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1098_
timestamp 0
transform -1 0 4310 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1099_
timestamp 0
transform -1 0 4450 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1100_
timestamp 0
transform 1 0 4130 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1101_
timestamp 0
transform -1 0 5550 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1102_
timestamp 0
transform 1 0 5370 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1103_
timestamp 0
transform 1 0 4510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1104_
timestamp 0
transform 1 0 5850 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1105_
timestamp 0
transform -1 0 5890 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1106_
timestamp 0
transform -1 0 5730 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1107_
timestamp 0
transform -1 0 3790 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1108_
timestamp 0
transform 1 0 4150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1109_
timestamp 0
transform -1 0 4790 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1110_
timestamp 0
transform -1 0 4350 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1111_
timestamp 0
transform 1 0 4430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1112_
timestamp 0
transform 1 0 4530 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1113_
timestamp 0
transform 1 0 5830 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1114_
timestamp 0
transform 1 0 5090 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1115_
timestamp 0
transform 1 0 4810 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1116_
timestamp 0
transform -1 0 4530 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1117_
timestamp 0
transform 1 0 4650 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1118_
timestamp 0
transform -1 0 4950 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1119_
timestamp 0
transform 1 0 5570 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1120_
timestamp 0
transform 1 0 5430 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1121_
timestamp 0
transform -1 0 5250 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1122_
timestamp 0
transform 1 0 5550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1123_
timestamp 0
transform 1 0 5550 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1124_
timestamp 0
transform 1 0 5050 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1125_
timestamp 0
transform -1 0 5410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1126_
timestamp 0
transform 1 0 5410 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1127_
timestamp 0
transform 1 0 5050 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1128_
timestamp 0
transform 1 0 5710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1129_
timestamp 0
transform 1 0 5570 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1130_
timestamp 0
transform 1 0 5690 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1131_
timestamp 0
transform 1 0 5230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1132_
timestamp 0
transform 1 0 5850 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1133_
timestamp 0
transform 1 0 5690 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1134_
timestamp 0
transform 1 0 5710 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1135_
timestamp 0
transform 1 0 5550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1136_
timestamp 0
transform 1 0 5770 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1137_
timestamp 0
transform -1 0 5670 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1138_
timestamp 0
transform -1 0 5410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1139_
timestamp 0
transform 1 0 5190 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1140_
timestamp 0
transform 1 0 5530 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1141_
timestamp 0
transform 1 0 5350 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1142_
timestamp 0
transform 1 0 5490 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1143_
timestamp 0
transform -1 0 5710 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1144_
timestamp 0
transform -1 0 5390 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1145_
timestamp 0
transform 1 0 5270 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1146_
timestamp 0
transform 1 0 4590 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1147_
timestamp 0
transform -1 0 3970 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1148_
timestamp 0
transform -1 0 5170 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1149_
timestamp 0
transform -1 0 5010 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1150_
timestamp 0
transform 1 0 4590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1151_
timestamp 0
transform 1 0 4410 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1152_
timestamp 0
transform -1 0 5270 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1153_
timestamp 0
transform -1 0 3130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1154_
timestamp 0
transform -1 0 3510 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1155_
timestamp 0
transform 1 0 4010 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1156_
timestamp 0
transform -1 0 3430 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1157_
timestamp 0
transform 1 0 3550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1158_
timestamp 0
transform 1 0 3250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1159_
timestamp 0
transform 1 0 4390 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1160_
timestamp 0
transform 1 0 4290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1161_
timestamp 0
transform -1 0 4250 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1162_
timestamp 0
transform 1 0 3570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1163_
timestamp 0
transform -1 0 3750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1164_
timestamp 0
transform -1 0 4770 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1165_
timestamp 0
transform 1 0 4910 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1166_
timestamp 0
transform -1 0 4270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1167_
timestamp 0
transform -1 0 4590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1168_
timestamp 0
transform -1 0 4910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1169_
timestamp 0
transform 1 0 4410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1170_
timestamp 0
transform -1 0 4310 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1171_
timestamp 0
transform 1 0 4690 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1172_
timestamp 0
transform 1 0 4530 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1173_
timestamp 0
transform 1 0 4730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1174_
timestamp 0
transform 1 0 4870 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1175_
timestamp 0
transform 1 0 5030 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1176_
timestamp 0
transform -1 0 5090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1177_
timestamp 0
transform 1 0 5210 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1178_
timestamp 0
transform 1 0 5810 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1179_
timestamp 0
transform -1 0 5750 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1180_
timestamp 0
transform 1 0 5570 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1181_
timestamp 0
transform -1 0 5430 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1182_
timestamp 0
transform -1 0 4810 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1183_
timestamp 0
transform 1 0 4130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1184_
timestamp 0
transform -1 0 4290 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1185_
timestamp 0
transform -1 0 1350 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1186_
timestamp 0
transform 1 0 5470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1187_
timestamp 0
transform -1 0 5350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1188_
timestamp 0
transform 1 0 5750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1189_
timestamp 0
transform 1 0 5610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1190_
timestamp 0
transform -1 0 5670 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1191_
timestamp 0
transform 1 0 5170 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1192_
timestamp 0
transform -1 0 4470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1193_
timestamp 0
transform -1 0 4110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1194_
timestamp 0
transform 1 0 5450 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1195_
timestamp 0
transform 1 0 5230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1196_
timestamp 0
transform -1 0 4050 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1197_
timestamp 0
transform -1 0 3870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1198_
timestamp 0
transform 1 0 3890 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1199_
timestamp 0
transform 1 0 3770 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1200_
timestamp 0
transform 1 0 3870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1201_
timestamp 0
transform -1 0 4610 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1202_
timestamp 0
transform 1 0 4750 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1203_
timestamp 0
transform 1 0 5390 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1204_
timestamp 0
transform 1 0 5290 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1205_
timestamp 0
transform 1 0 5270 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1206_
timestamp 0
transform 1 0 5110 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1207_
timestamp 0
transform -1 0 5150 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1208_
timestamp 0
transform -1 0 4990 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1209_
timestamp 0
transform -1 0 4990 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1210_
timestamp 0
transform 1 0 4830 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1211_
timestamp 0
transform 1 0 4770 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1212_
timestamp 0
transform -1 0 4730 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1213_
timestamp 0
transform 1 0 3970 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1214_
timestamp 0
transform -1 0 4930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1215_
timestamp 0
transform 1 0 4110 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1216_
timestamp 0
transform -1 0 5390 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1217_
timestamp 0
transform 1 0 5210 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1218_
timestamp 0
transform -1 0 4630 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1219_
timestamp 0
transform 1 0 1710 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1220_
timestamp 0
transform 1 0 630 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1221_
timestamp 0
transform 1 0 5110 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1222_
timestamp 0
transform 1 0 4110 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1223_
timestamp 0
transform 1 0 3930 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1224_
timestamp 0
transform 1 0 3410 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1225_
timestamp 0
transform 1 0 3710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1226_
timestamp 0
transform -1 0 3730 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1227_
timestamp 0
transform 1 0 3830 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1228_
timestamp 0
transform -1 0 3570 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1229_
timestamp 0
transform -1 0 4250 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1230_
timestamp 0
transform 1 0 4910 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1231_
timestamp 0
transform 1 0 4690 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1232_
timestamp 0
transform -1 0 4550 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1233_
timestamp 0
transform -1 0 4690 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1234_
timestamp 0
transform -1 0 4550 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1235_
timestamp 0
transform -1 0 4390 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1236_
timestamp 0
transform 1 0 770 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1237_
timestamp 0
transform -1 0 4370 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1238_
timestamp 0
transform 1 0 5710 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1239_
timestamp 0
transform 1 0 5270 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1240_
timestamp 0
transform -1 0 5450 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1241_
timestamp 0
transform 1 0 4810 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1242_
timestamp 0
transform 1 0 4890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1243_
timestamp 0
transform -1 0 3950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1244_
timestamp 0
transform 1 0 3590 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1245_
timestamp 0
transform -1 0 3790 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1246_
timestamp 0
transform 1 0 3990 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1247_
timestamp 0
transform 1 0 4070 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1248_
timestamp 0
transform 1 0 4110 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1249_
timestamp 0
transform 1 0 4630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1250_
timestamp 0
transform 1 0 5050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1251_
timestamp 0
transform -1 0 5510 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1252_
timestamp 0
transform -1 0 5070 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1253_
timestamp 0
transform 1 0 4770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1254_
timestamp 0
transform 1 0 4890 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1255_
timestamp 0
transform 1 0 4710 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1256_
timestamp 0
transform -1 0 4270 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1257_
timestamp 0
transform -1 0 4450 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1258_
timestamp 0
transform 1 0 4270 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1259_
timestamp 0
transform 1 0 4430 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1260_
timestamp 0
transform 1 0 1770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1261_
timestamp 0
transform 1 0 1210 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1262_
timestamp 0
transform -1 0 1530 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1263_
timestamp 0
transform -1 0 1390 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1264_
timestamp 0
transform -1 0 930 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1265_
timestamp 0
transform -1 0 1310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1266_
timestamp 0
transform -1 0 1450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1267_
timestamp 0
transform -1 0 1310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1268_
timestamp 0
transform -1 0 1270 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1269_
timestamp 0
transform -1 0 970 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1270_
timestamp 0
transform -1 0 1090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1271_
timestamp 0
transform 1 0 1090 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1272_
timestamp 0
transform -1 0 950 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1273_
timestamp 0
transform 1 0 610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1274_
timestamp 0
transform -1 0 790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1275_
timestamp 0
transform -1 0 1150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1276_
timestamp 0
transform -1 0 790 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1277_
timestamp 0
transform 1 0 570 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1278_
timestamp 0
transform -1 0 450 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1279_
timestamp 0
transform -1 0 590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1280_
timestamp 0
transform 1 0 950 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1281_
timestamp 0
transform -1 0 810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1282_
timestamp 0
transform 1 0 730 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1283_
timestamp 0
transform 1 0 870 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1284_
timestamp 0
transform 1 0 590 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1285_
timestamp 0
transform -1 0 350 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1286_
timestamp 0
transform 1 0 270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1287_
timestamp 0
transform -1 0 290 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1288_
timestamp 0
transform 1 0 730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1289_
timestamp 0
transform 1 0 30 0 -1 5470
box -6 -8 26 268
use FILL  FILL_1__1290_
timestamp 0
transform 1 0 150 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1__1291_
timestamp 0
transform 1 0 30 0 1 5470
box -6 -8 26 268
use FILL  FILL_1__1292_
timestamp 0
transform -1 0 50 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1293_
timestamp 0
transform -1 0 590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1294_
timestamp 0
transform -1 0 430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1295_
timestamp 0
transform 1 0 170 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1296_
timestamp 0
transform 1 0 30 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1297_
timestamp 0
transform 1 0 150 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1298_
timestamp 0
transform 1 0 450 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1299_
timestamp 0
transform 1 0 410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1300_
timestamp 0
transform -1 0 430 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1301_
timestamp 0
transform 1 0 290 0 1 4950
box -6 -8 26 268
use FILL  FILL_1__1302_
timestamp 0
transform -1 0 530 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1303_
timestamp 0
transform 1 0 690 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1304_
timestamp 0
transform -1 0 370 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1305_
timestamp 0
transform -1 0 470 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1306_
timestamp 0
transform -1 0 310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1__1307_
timestamp 0
transform 1 0 170 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1308_
timestamp 0
transform 1 0 290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1309_
timestamp 0
transform 1 0 490 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1310_
timestamp 0
transform 1 0 270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1311_
timestamp 0
transform -1 0 50 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1312_
timestamp 0
transform -1 0 410 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1313_
timestamp 0
transform -1 0 50 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1314_
timestamp 0
transform -1 0 190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1315_
timestamp 0
transform -1 0 210 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1316_
timestamp 0
transform 1 0 30 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1317_
timestamp 0
transform -1 0 330 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1318_
timestamp 0
transform -1 0 1190 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1319_
timestamp 0
transform 1 0 1210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1320_
timestamp 0
transform -1 0 1110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1321_
timestamp 0
transform -1 0 910 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1322_
timestamp 0
transform -1 0 210 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1323_
timestamp 0
transform 1 0 270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1324_
timestamp 0
transform -1 0 290 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1325_
timestamp 0
transform 1 0 1710 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1326_
timestamp 0
transform 1 0 190 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1327_
timestamp 0
transform 1 0 790 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1328_
timestamp 0
transform 1 0 930 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1329_
timestamp 0
transform -1 0 50 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1330_
timestamp 0
transform 1 0 590 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1331_
timestamp 0
transform -1 0 50 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1332_
timestamp 0
transform 1 0 590 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1333_
timestamp 0
transform 1 0 750 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1334_
timestamp 0
transform -1 0 2610 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1335_
timestamp 0
transform 1 0 2750 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1336_
timestamp 0
transform -1 0 2450 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1337_
timestamp 0
transform -1 0 2190 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1338_
timestamp 0
transform 1 0 2170 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1339_
timestamp 0
transform -1 0 2330 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1340_
timestamp 0
transform -1 0 2030 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1341_
timestamp 0
transform -1 0 1870 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1342_
timestamp 0
transform 1 0 2370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1343_
timestamp 0
transform 1 0 3450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1344_
timestamp 0
transform 1 0 3590 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1345_
timestamp 0
transform 1 0 2970 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1346_
timestamp 0
transform 1 0 2810 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1347_
timestamp 0
transform -1 0 2550 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1348_
timestamp 0
transform -1 0 2190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1349_
timestamp 0
transform -1 0 1350 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1350_
timestamp 0
transform -1 0 1730 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1351_
timestamp 0
transform -1 0 450 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1352_
timestamp 0
transform -1 0 2050 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1353_
timestamp 0
transform -1 0 2670 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1354_
timestamp 0
transform -1 0 1890 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1355_
timestamp 0
transform -1 0 1210 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1356_
timestamp 0
transform -1 0 1070 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1357_
timestamp 0
transform -1 0 790 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1358_
timestamp 0
transform 1 0 650 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1359_
timestamp 0
transform 1 0 570 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1360_
timestamp 0
transform 1 0 910 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1361_
timestamp 0
transform -1 0 750 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1362_
timestamp 0
transform -1 0 530 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1363_
timestamp 0
transform -1 0 250 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1364_
timestamp 0
transform 1 0 170 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1365_
timestamp 0
transform 1 0 150 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1366_
timestamp 0
transform -1 0 50 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1367_
timestamp 0
transform -1 0 50 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1368_
timestamp 0
transform -1 0 50 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1369_
timestamp 0
transform 1 0 190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1370_
timestamp 0
transform -1 0 50 0 -1 1310
box -6 -8 26 268
use FILL  FILL_1__1371_
timestamp 0
transform -1 0 2830 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1372_
timestamp 0
transform 1 0 310 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1373_
timestamp 0
transform -1 0 390 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1374_
timestamp 0
transform -1 0 490 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1375_
timestamp 0
transform -1 0 3970 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1376_
timestamp 0
transform 1 0 4090 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1377_
timestamp 0
transform -1 0 3690 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1378_
timestamp 0
transform 1 0 3790 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1379_
timestamp 0
transform -1 0 2970 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1380_
timestamp 0
transform -1 0 3150 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1381_
timestamp 0
transform 1 0 3250 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1382_
timestamp 0
transform -1 0 3110 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1383_
timestamp 0
transform -1 0 2970 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1384_
timestamp 0
transform 1 0 3510 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1385_
timestamp 0
transform 1 0 4230 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1386_
timestamp 0
transform -1 0 3990 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1387_
timestamp 0
transform -1 0 3850 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1388_
timestamp 0
transform 1 0 3870 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1389_
timestamp 0
transform -1 0 3550 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1390_
timestamp 0
transform 1 0 3690 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1391_
timestamp 0
transform 1 0 3350 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1392_
timestamp 0
transform -1 0 3690 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1393_
timestamp 0
transform -1 0 3570 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1394_
timestamp 0
transform -1 0 3390 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1395_
timestamp 0
transform -1 0 3270 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1396_
timestamp 0
transform -1 0 2590 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1397_
timestamp 0
transform 1 0 2270 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1398_
timestamp 0
transform 1 0 2690 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1399_
timestamp 0
transform 1 0 2230 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1400_
timestamp 0
transform -1 0 1750 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1401_
timestamp 0
transform -1 0 2130 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1402_
timestamp 0
transform -1 0 2430 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1403_
timestamp 0
transform -1 0 1990 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1404_
timestamp 0
transform -1 0 1890 0 1 790
box -6 -8 26 268
use FILL  FILL_1__1405_
timestamp 0
transform -1 0 3430 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1406_
timestamp 0
transform 1 0 1450 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1407_
timestamp 0
transform 1 0 3490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1408_
timestamp 0
transform 1 0 3330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1__1409_
timestamp 0
transform 1 0 3330 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1410_
timestamp 0
transform -1 0 3630 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1411_
timestamp 0
transform 1 0 3450 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1412_
timestamp 0
transform 1 0 2850 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1413_
timestamp 0
transform 1 0 2950 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1414_
timestamp 0
transform 1 0 2970 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1415_
timestamp 0
transform 1 0 1850 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1416_
timestamp 0
transform -1 0 1510 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1417_
timestamp 0
transform 1 0 1450 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1418_
timestamp 0
transform -1 0 870 0 1 1310
box -6 -8 26 268
use FILL  FILL_1__1419_
timestamp 0
transform 1 0 3090 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1420_
timestamp 0
transform 1 0 3230 0 1 2350
box -6 -8 26 268
use FILL  FILL_1__1421_
timestamp 0
transform -1 0 3030 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1422_
timestamp 0
transform 1 0 3150 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1423_
timestamp 0
transform -1 0 2430 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1424_
timestamp 0
transform -1 0 2810 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1425_
timestamp 0
transform 1 0 1150 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1426_
timestamp 0
transform -1 0 1310 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1427_
timestamp 0
transform 1 0 1890 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1428_
timestamp 0
transform -1 0 2170 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1429_
timestamp 0
transform -1 0 2330 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1430_
timestamp 0
transform 1 0 2390 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1431_
timestamp 0
transform -1 0 2730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1432_
timestamp 0
transform 1 0 2070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1433_
timestamp 0
transform -1 0 2250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1434_
timestamp 0
transform -1 0 2230 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1435_
timestamp 0
transform 1 0 2050 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1436_
timestamp 0
transform -1 0 2210 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1437_
timestamp 0
transform -1 0 2590 0 1 1830
box -6 -8 26 268
use FILL  FILL_1__1438_
timestamp 0
transform -1 0 2550 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1439_
timestamp 0
transform -1 0 2690 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1440_
timestamp 0
transform -1 0 2490 0 1 2870
box -6 -8 26 268
use FILL  FILL_1__1441_
timestamp 0
transform 1 0 2550 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1__1442_
timestamp 0
transform -1 0 1490 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1443_
timestamp 0
transform 1 0 1610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1__1444_
timestamp 0
transform -1 0 2650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1445_
timestamp 0
transform -1 0 2790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1446_
timestamp 0
transform -1 0 3090 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1447_
timestamp 0
transform -1 0 3110 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1448_
timestamp 0
transform -1 0 3230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1__1449_
timestamp 0
transform -1 0 3510 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1450_
timestamp 0
transform -1 0 2410 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1451_
timestamp 0
transform -1 0 2670 0 1 3390
box -6 -8 26 268
use FILL  FILL_1__1527_
timestamp 0
transform 1 0 5510 0 1 270
box -6 -8 26 268
use FILL  FILL_1__1528_
timestamp 0
transform 1 0 3610 0 -1 3390
box -6 -8 26 268
use FILL  FILL_1__1529_
timestamp 0
transform 1 0 4510 0 1 3910
box -6 -8 26 268
use FILL  FILL_1__1530_
timestamp 0
transform 1 0 5370 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1__1531_
timestamp 0
transform 1 0 5850 0 1 4430
box -6 -8 26 268
use FILL  FILL_1__1532_
timestamp 0
transform 1 0 910 0 -1 790
box -6 -8 26 268
use FILL  FILL_1__1533_
timestamp 0
transform -1 0 450 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1534_
timestamp 0
transform -1 0 310 0 -1 270
box -6 -8 26 268
use FILL  FILL_1__1535_
timestamp 0
transform -1 0 50 0 1 790
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert0
timestamp 0
transform -1 0 1050 0 1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert1
timestamp 0
transform 1 0 2970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert2
timestamp 0
transform -1 0 1090 0 1 790
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert3
timestamp 0
transform -1 0 990 0 1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert4
timestamp 0
transform 1 0 1590 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert5
timestamp 0
transform -1 0 2290 0 1 790
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert6
timestamp 0
transform 1 0 2950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert15
timestamp 0
transform -1 0 2690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert16
timestamp 0
transform -1 0 2870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert17
timestamp 0
transform -1 0 3970 0 -1 4430
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert18
timestamp 0
transform 1 0 4270 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert19
timestamp 0
transform -1 0 470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert20
timestamp 0
transform 1 0 1090 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert21
timestamp 0
transform -1 0 450 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert22
timestamp 0
transform -1 0 830 0 1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert23
timestamp 0
transform 1 0 2290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert24
timestamp 0
transform 1 0 2730 0 1 1830
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert25
timestamp 0
transform 1 0 3230 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert26
timestamp 0
transform -1 0 3130 0 -1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert27
timestamp 0
transform -1 0 2850 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert28
timestamp 0
transform -1 0 2870 0 1 2870
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert29
timestamp 0
transform 1 0 1330 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert30
timestamp 0
transform 1 0 4650 0 1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert31
timestamp 0
transform -1 0 2970 0 1 3910
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert32
timestamp 0
transform 1 0 4630 0 1 3390
box -6 -8 26 268
use FILL  FILL_1_BUFX2_insert33
timestamp 0
transform -1 0 2810 0 1 3910
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert7
timestamp 0
transform 1 0 770 0 -1 5990
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert8
timestamp 0
transform -1 0 50 0 -1 1830
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert9
timestamp 0
transform 1 0 2270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert10
timestamp 0
transform -1 0 50 0 1 1830
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert11
timestamp 0
transform 1 0 170 0 1 790
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert12
timestamp 0
transform 1 0 2290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert13
timestamp 0
transform 1 0 1870 0 -1 3910
box -6 -8 26 268
use FILL  FILL_1_CLKBUF1_insert14
timestamp 0
transform 1 0 2550 0 1 790
box -6 -8 26 268
use FILL  FILL_2__723_
timestamp 0
transform 1 0 1170 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__724_
timestamp 0
transform -1 0 650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__725_
timestamp 0
transform -1 0 1650 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__726_
timestamp 0
transform -1 0 1330 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__727_
timestamp 0
transform 1 0 1970 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__728_
timestamp 0
transform -1 0 2050 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__729_
timestamp 0
transform -1 0 770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__730_
timestamp 0
transform -1 0 1030 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__731_
timestamp 0
transform 1 0 450 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__732_
timestamp 0
transform -1 0 3130 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__733_
timestamp 0
transform 1 0 1210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__734_
timestamp 0
transform -1 0 1070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__735_
timestamp 0
transform -1 0 510 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__736_
timestamp 0
transform -1 0 590 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__737_
timestamp 0
transform -1 0 1910 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__738_
timestamp 0
transform 1 0 910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__739_
timestamp 0
transform 1 0 510 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__740_
timestamp 0
transform -1 0 450 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__741_
timestamp 0
transform -1 0 370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__742_
timestamp 0
transform 1 0 730 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__743_
timestamp 0
transform -1 0 330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__744_
timestamp 0
transform -1 0 330 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__745_
timestamp 0
transform -1 0 310 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__746_
timestamp 0
transform 1 0 3510 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__747_
timestamp 0
transform -1 0 3230 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__748_
timestamp 0
transform 1 0 3350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__749_
timestamp 0
transform 1 0 3910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__750_
timestamp 0
transform -1 0 3950 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__751_
timestamp 0
transform -1 0 4090 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__752_
timestamp 0
transform 1 0 4030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__753_
timestamp 0
transform -1 0 4250 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__754_
timestamp 0
transform 1 0 4370 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__755_
timestamp 0
transform -1 0 3670 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__756_
timestamp 0
transform -1 0 4370 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__757_
timestamp 0
transform 1 0 4490 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__758_
timestamp 0
transform 1 0 3270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__759_
timestamp 0
transform -1 0 3430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__760_
timestamp 0
transform 1 0 3370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__761_
timestamp 0
transform -1 0 3530 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__762_
timestamp 0
transform 1 0 2950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__763_
timestamp 0
transform -1 0 2970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__764_
timestamp 0
transform 1 0 3070 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__765_
timestamp 0
transform -1 0 3370 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__766_
timestamp 0
transform 1 0 2170 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__767_
timestamp 0
transform -1 0 2090 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__768_
timestamp 0
transform 1 0 1910 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__769_
timestamp 0
transform -1 0 1590 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__770_
timestamp 0
transform 1 0 1810 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__771_
timestamp 0
transform 1 0 1650 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__772_
timestamp 0
transform -1 0 1010 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__773_
timestamp 0
transform 1 0 1790 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__774_
timestamp 0
transform -1 0 1270 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__775_
timestamp 0
transform 1 0 710 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__776_
timestamp 0
transform 1 0 1410 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__777_
timestamp 0
transform 1 0 830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__778_
timestamp 0
transform -1 0 70 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__779_
timestamp 0
transform 1 0 1750 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__780_
timestamp 0
transform -1 0 330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__781_
timestamp 0
transform -1 0 810 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__782_
timestamp 0
transform 1 0 1930 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__783_
timestamp 0
transform 1 0 1150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__784_
timestamp 0
transform 1 0 670 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__785_
timestamp 0
transform 1 0 950 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__786_
timestamp 0
transform 1 0 790 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__787_
timestamp 0
transform 1 0 1330 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__788_
timestamp 0
transform 1 0 1770 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__789_
timestamp 0
transform 1 0 1450 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__790_
timestamp 0
transform 1 0 2690 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__791_
timestamp 0
transform 1 0 2890 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__792_
timestamp 0
transform 1 0 2810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__793_
timestamp 0
transform 1 0 3150 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__794_
timestamp 0
transform 1 0 3430 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__795_
timestamp 0
transform 1 0 3270 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__796_
timestamp 0
transform -1 0 1250 0 1 790
box -6 -8 26 268
use FILL  FILL_2__797_
timestamp 0
transform 1 0 2430 0 1 790
box -6 -8 26 268
use FILL  FILL_2__798_
timestamp 0
transform 1 0 1590 0 1 790
box -6 -8 26 268
use FILL  FILL_2__799_
timestamp 0
transform 1 0 830 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__800_
timestamp 0
transform 1 0 1130 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__801_
timestamp 0
transform 1 0 970 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__802_
timestamp 0
transform -1 0 4030 0 1 790
box -6 -8 26 268
use FILL  FILL_2__803_
timestamp 0
transform -1 0 3670 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__804_
timestamp 0
transform -1 0 4010 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__805_
timestamp 0
transform -1 0 4150 0 1 270
box -6 -8 26 268
use FILL  FILL_2__806_
timestamp 0
transform -1 0 4030 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__807_
timestamp 0
transform 1 0 4150 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__808_
timestamp 0
transform -1 0 2330 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__809_
timestamp 0
transform 1 0 2830 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__810_
timestamp 0
transform 1 0 2670 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__811_
timestamp 0
transform 1 0 2190 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__812_
timestamp 0
transform -1 0 1670 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__813_
timestamp 0
transform -1 0 1810 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__814_
timestamp 0
transform -1 0 2110 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__815_
timestamp 0
transform 1 0 2150 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__816_
timestamp 0
transform 1 0 2230 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__817_
timestamp 0
transform 1 0 2010 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__818_
timestamp 0
transform 1 0 2370 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__819_
timestamp 0
transform -1 0 2090 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__820_
timestamp 0
transform 1 0 1730 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__821_
timestamp 0
transform 1 0 1550 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__822_
timestamp 0
transform -1 0 1710 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__823_
timestamp 0
transform 1 0 1930 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__824_
timestamp 0
transform -1 0 1910 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__825_
timestamp 0
transform 1 0 2690 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__826_
timestamp 0
transform 1 0 2090 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__827_
timestamp 0
transform 1 0 2510 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__828_
timestamp 0
transform -1 0 1930 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__829_
timestamp 0
transform -1 0 1150 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__830_
timestamp 0
transform -1 0 2230 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__831_
timestamp 0
transform -1 0 2390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__832_
timestamp 0
transform 1 0 2230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__833_
timestamp 0
transform -1 0 3190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__834_
timestamp 0
transform -1 0 2710 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__835_
timestamp 0
transform -1 0 2530 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__836_
timestamp 0
transform -1 0 2670 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__837_
timestamp 0
transform -1 0 1270 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__838_
timestamp 0
transform 1 0 1750 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__839_
timestamp 0
transform -1 0 1330 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__840_
timestamp 0
transform -1 0 1610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__841_
timestamp 0
transform -1 0 1450 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__842_
timestamp 0
transform 1 0 1110 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__843_
timestamp 0
transform 1 0 1230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__844_
timestamp 0
transform -1 0 1410 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__845_
timestamp 0
transform 1 0 1030 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__846_
timestamp 0
transform 1 0 3430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__847_
timestamp 0
transform 1 0 1410 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__848_
timestamp 0
transform 1 0 2150 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__849_
timestamp 0
transform 1 0 2730 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__850_
timestamp 0
transform 1 0 2590 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__851_
timestamp 0
transform -1 0 2350 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__852_
timestamp 0
transform 1 0 2430 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__853_
timestamp 0
transform 1 0 2150 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__854_
timestamp 0
transform -1 0 2190 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__855_
timestamp 0
transform -1 0 2050 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__856_
timestamp 0
transform -1 0 2310 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__857_
timestamp 0
transform -1 0 2010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__858_
timestamp 0
transform -1 0 1670 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__859_
timestamp 0
transform -1 0 1590 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__860_
timestamp 0
transform -1 0 1850 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__861_
timestamp 0
transform -1 0 3710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__862_
timestamp 0
transform -1 0 2990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__863_
timestamp 0
transform -1 0 2570 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__864_
timestamp 0
transform -1 0 2590 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__865_
timestamp 0
transform -1 0 2550 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__866_
timestamp 0
transform -1 0 1750 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__867_
timestamp 0
transform 1 0 1670 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__868_
timestamp 0
transform -1 0 1510 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__869_
timestamp 0
transform -1 0 1570 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__870_
timestamp 0
transform 1 0 1990 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__871_
timestamp 0
transform -1 0 1530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__872_
timestamp 0
transform -1 0 1390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__873_
timestamp 0
transform -1 0 1370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__874_
timestamp 0
transform -1 0 1350 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__875_
timestamp 0
transform -1 0 1130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__876_
timestamp 0
transform 1 0 1150 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__877_
timestamp 0
transform 1 0 210 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__878_
timestamp 0
transform -1 0 1010 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__879_
timestamp 0
transform -1 0 1850 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__880_
timestamp 0
transform 1 0 1670 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__881_
timestamp 0
transform -1 0 2430 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__882_
timestamp 0
transform 1 0 3270 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__883_
timestamp 0
transform 1 0 2830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__884_
timestamp 0
transform -1 0 2830 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__885_
timestamp 0
transform -1 0 2330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__886_
timestamp 0
transform 1 0 2710 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__887_
timestamp 0
transform -1 0 2590 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__888_
timestamp 0
transform -1 0 2450 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__889_
timestamp 0
transform -1 0 3150 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__890_
timestamp 0
transform 1 0 3030 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__891_
timestamp 0
transform 1 0 2670 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__892_
timestamp 0
transform -1 0 2370 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__893_
timestamp 0
transform 1 0 2270 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__894_
timestamp 0
transform -1 0 2170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__895_
timestamp 0
transform -1 0 2610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__896_
timestamp 0
transform 1 0 1990 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__897_
timestamp 0
transform 1 0 3570 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__898_
timestamp 0
transform -1 0 2850 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__899_
timestamp 0
transform 1 0 3390 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__900_
timestamp 0
transform 1 0 3430 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__901_
timestamp 0
transform 1 0 2990 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__902_
timestamp 0
transform -1 0 3030 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__903_
timestamp 0
transform -1 0 2210 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__904_
timestamp 0
transform -1 0 1850 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__905_
timestamp 0
transform 1 0 2510 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__906_
timestamp 0
transform -1 0 2170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__907_
timestamp 0
transform -1 0 2010 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__908_
timestamp 0
transform -1 0 1730 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__909_
timestamp 0
transform -1 0 1270 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__910_
timestamp 0
transform 1 0 1550 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__911_
timestamp 0
transform -1 0 1890 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__912_
timestamp 0
transform -1 0 1890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__913_
timestamp 0
transform -1 0 1730 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__914_
timestamp 0
transform -1 0 1250 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__915_
timestamp 0
transform 1 0 1390 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__916_
timestamp 0
transform 1 0 1070 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__917_
timestamp 0
transform 1 0 750 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__918_
timestamp 0
transform -1 0 3870 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__919_
timestamp 0
transform -1 0 2770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__920_
timestamp 0
transform 1 0 2750 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__921_
timestamp 0
transform 1 0 2030 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__922_
timestamp 0
transform 1 0 3710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__923_
timestamp 0
transform -1 0 3350 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__924_
timestamp 0
transform 1 0 3170 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__925_
timestamp 0
transform 1 0 3570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__926_
timestamp 0
transform -1 0 3810 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__927_
timestamp 0
transform 1 0 3630 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__928_
timestamp 0
transform -1 0 3530 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__929_
timestamp 0
transform -1 0 3310 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__930_
timestamp 0
transform 1 0 3170 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__931_
timestamp 0
transform 1 0 3330 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__932_
timestamp 0
transform -1 0 3390 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__933_
timestamp 0
transform -1 0 2870 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__934_
timestamp 0
transform -1 0 4270 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__935_
timestamp 0
transform 1 0 4950 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__936_
timestamp 0
transform -1 0 4130 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__937_
timestamp 0
transform -1 0 4290 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__938_
timestamp 0
transform -1 0 4610 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__939_
timestamp 0
transform -1 0 4670 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__940_
timestamp 0
transform 1 0 5090 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__941_
timestamp 0
transform -1 0 4450 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__942_
timestamp 0
transform 1 0 4410 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__943_
timestamp 0
transform -1 0 3830 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__944_
timestamp 0
transform 1 0 4630 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__945_
timestamp 0
transform -1 0 4150 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__946_
timestamp 0
transform -1 0 4490 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__947_
timestamp 0
transform 1 0 4810 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__948_
timestamp 0
transform -1 0 3830 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__949_
timestamp 0
transform -1 0 3650 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__950_
timestamp 0
transform -1 0 3230 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__951_
timestamp 0
transform -1 0 4330 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__952_
timestamp 0
transform 1 0 3970 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__953_
timestamp 0
transform -1 0 2910 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__954_
timestamp 0
transform -1 0 3010 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__955_
timestamp 0
transform 1 0 2430 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__956_
timestamp 0
transform -1 0 3070 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__957_
timestamp 0
transform -1 0 3490 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__958_
timestamp 0
transform -1 0 3170 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__959_
timestamp 0
transform -1 0 2850 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__960_
timestamp 0
transform -1 0 2890 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__961_
timestamp 0
transform 1 0 3310 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__962_
timestamp 0
transform -1 0 2610 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__963_
timestamp 0
transform -1 0 1410 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__964_
timestamp 0
transform -1 0 1270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__965_
timestamp 0
transform 1 0 1050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__966_
timestamp 0
transform 1 0 850 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__967_
timestamp 0
transform -1 0 970 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__968_
timestamp 0
transform 1 0 190 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__969_
timestamp 0
transform -1 0 1550 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__970_
timestamp 0
transform 1 0 3050 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__971_
timestamp 0
transform 1 0 3210 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__972_
timestamp 0
transform 1 0 3650 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__973_
timestamp 0
transform 1 0 3490 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__974_
timestamp 0
transform -1 0 5290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__975_
timestamp 0
transform -1 0 3530 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__976_
timestamp 0
transform 1 0 3650 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__977_
timestamp 0
transform 1 0 3950 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__978_
timestamp 0
transform -1 0 4130 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__979_
timestamp 0
transform 1 0 3950 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__980_
timestamp 0
transform -1 0 4190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__981_
timestamp 0
transform 1 0 4010 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__982_
timestamp 0
transform 1 0 4090 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__983_
timestamp 0
transform -1 0 4390 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__984_
timestamp 0
transform 1 0 4330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__985_
timestamp 0
transform 1 0 3790 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__986_
timestamp 0
transform 1 0 4490 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__987_
timestamp 0
transform -1 0 5130 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__988_
timestamp 0
transform 1 0 4270 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__989_
timestamp 0
transform -1 0 4430 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__990_
timestamp 0
transform 1 0 4810 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__991_
timestamp 0
transform -1 0 4610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__992_
timestamp 0
transform 1 0 4950 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__993_
timestamp 0
transform -1 0 5130 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__994_
timestamp 0
transform 1 0 5030 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__995_
timestamp 0
transform 1 0 5070 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__996_
timestamp 0
transform 1 0 5290 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__997_
timestamp 0
transform 1 0 4950 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__998_
timestamp 0
transform -1 0 4910 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__999_
timestamp 0
transform 1 0 4730 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1000_
timestamp 0
transform 1 0 5230 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1001_
timestamp 0
transform -1 0 5090 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1002_
timestamp 0
transform -1 0 4570 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1003_
timestamp 0
transform -1 0 4810 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1004_
timestamp 0
transform 1 0 4730 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1005_
timestamp 0
transform -1 0 4930 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1006_
timestamp 0
transform -1 0 4770 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1007_
timestamp 0
transform -1 0 5230 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1008_
timestamp 0
transform 1 0 5250 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1009_
timestamp 0
transform 1 0 5530 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1010_
timestamp 0
transform 1 0 4910 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1011_
timestamp 0
transform -1 0 5290 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1012_
timestamp 0
transform 1 0 4950 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1013_
timestamp 0
transform 1 0 4470 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1014_
timestamp 0
transform 1 0 4630 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1015_
timestamp 0
transform 1 0 5430 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1016_
timestamp 0
transform 1 0 5370 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1017_
timestamp 0
transform -1 0 5130 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1018_
timestamp 0
transform -1 0 4970 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1019_
timestamp 0
transform -1 0 4910 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1020_
timestamp 0
transform -1 0 4810 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1021_
timestamp 0
transform -1 0 4810 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1022_
timestamp 0
transform 1 0 4490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1023_
timestamp 0
transform -1 0 3670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1024_
timestamp 0
transform 1 0 2270 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1025_
timestamp 0
transform -1 0 4350 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1026_
timestamp 0
transform 1 0 3370 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1027_
timestamp 0
transform 1 0 3490 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1028_
timestamp 0
transform -1 0 4650 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1029_
timestamp 0
transform 1 0 5110 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1030_
timestamp 0
transform -1 0 4190 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1031_
timestamp 0
transform -1 0 4030 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1032_
timestamp 0
transform 1 0 930 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1033_
timestamp 0
transform 1 0 570 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1034_
timestamp 0
transform 1 0 3850 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1035_
timestamp 0
transform 1 0 5390 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1036_
timestamp 0
transform 1 0 5510 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1037_
timestamp 0
transform 1 0 4970 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1038_
timestamp 0
transform 1 0 5830 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1039_
timestamp 0
transform -1 0 5590 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1040_
timestamp 0
transform 1 0 5410 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1041_
timestamp 0
transform -1 0 4170 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1042_
timestamp 0
transform 1 0 4190 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1043_
timestamp 0
transform 1 0 4070 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1044_
timestamp 0
transform -1 0 3930 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1045_
timestamp 0
transform 1 0 3750 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1046_
timestamp 0
transform -1 0 4090 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1047_
timestamp 0
transform 1 0 4230 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1048_
timestamp 0
transform 1 0 4230 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1049_
timestamp 0
transform -1 0 3790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1050_
timestamp 0
transform -1 0 3930 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1051_
timestamp 0
transform 1 0 4370 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1052_
timestamp 0
transform -1 0 5270 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1053_
timestamp 0
transform 1 0 5190 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1054_
timestamp 0
transform -1 0 4990 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1055_
timestamp 0
transform -1 0 5130 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1056_
timestamp 0
transform 1 0 5350 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1057_
timestamp 0
transform 1 0 5170 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1058_
timestamp 0
transform -1 0 5650 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1059_
timestamp 0
transform -1 0 5630 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1060_
timestamp 0
transform -1 0 5030 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1061_
timestamp 0
transform 1 0 5490 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1062_
timestamp 0
transform 1 0 5730 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1063_
timestamp 0
transform 1 0 5790 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1064_
timestamp 0
transform 1 0 5710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1065_
timestamp 0
transform 1 0 5110 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1066_
timestamp 0
transform -1 0 5430 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1067_
timestamp 0
transform -1 0 5570 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1068_
timestamp 0
transform 1 0 4670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1069_
timestamp 0
transform 1 0 4790 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1070_
timestamp 0
transform 1 0 4850 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1071_
timestamp 0
transform 1 0 5550 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1072_
timestamp 0
transform 1 0 5570 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1073_
timestamp 0
transform 1 0 5390 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1074_
timestamp 0
transform 1 0 5670 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1075_
timestamp 0
transform -1 0 5410 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1076_
timestamp 0
transform -1 0 5710 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1077_
timestamp 0
transform 1 0 5710 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1078_
timestamp 0
transform 1 0 5230 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1079_
timestamp 0
transform 1 0 5710 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1080_
timestamp 0
transform 1 0 5850 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1081_
timestamp 0
transform 1 0 5530 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1082_
timestamp 0
transform 1 0 5670 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1083_
timestamp 0
transform -1 0 5710 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1084_
timestamp 0
transform 1 0 5710 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1085_
timestamp 0
transform -1 0 5770 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1086_
timestamp 0
transform -1 0 5610 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1087_
timestamp 0
transform -1 0 5550 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1088_
timestamp 0
transform 1 0 5050 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1089_
timestamp 0
transform 1 0 5210 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1090_
timestamp 0
transform -1 0 5770 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1091_
timestamp 0
transform 1 0 5830 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1092_
timestamp 0
transform 1 0 5370 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1093_
timestamp 0
transform 1 0 4590 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1094_
timestamp 0
transform -1 0 3810 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1095_
timestamp 0
transform 1 0 1610 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1096_
timestamp 0
transform -1 0 1590 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1097_
timestamp 0
transform 1 0 3810 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1098_
timestamp 0
transform -1 0 4330 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1099_
timestamp 0
transform -1 0 4470 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1100_
timestamp 0
transform 1 0 4150 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1101_
timestamp 0
transform -1 0 5570 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1102_
timestamp 0
transform 1 0 5390 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1103_
timestamp 0
transform 1 0 4530 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1104_
timestamp 0
transform 1 0 5870 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1105_
timestamp 0
transform -1 0 5910 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1106_
timestamp 0
transform -1 0 5750 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1107_
timestamp 0
transform -1 0 3810 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1108_
timestamp 0
transform 1 0 4170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1109_
timestamp 0
transform -1 0 4810 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1110_
timestamp 0
transform -1 0 4370 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1111_
timestamp 0
transform 1 0 4450 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1112_
timestamp 0
transform 1 0 4550 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1113_
timestamp 0
transform 1 0 5850 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1114_
timestamp 0
transform 1 0 5110 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1115_
timestamp 0
transform 1 0 4830 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1116_
timestamp 0
transform -1 0 4550 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1117_
timestamp 0
transform 1 0 4670 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1118_
timestamp 0
transform -1 0 4970 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1119_
timestamp 0
transform 1 0 5590 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1120_
timestamp 0
transform 1 0 5450 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1121_
timestamp 0
transform -1 0 5270 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1122_
timestamp 0
transform 1 0 5570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1123_
timestamp 0
transform 1 0 5570 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1124_
timestamp 0
transform 1 0 5070 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1125_
timestamp 0
transform -1 0 5430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1126_
timestamp 0
transform 1 0 5430 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1127_
timestamp 0
transform 1 0 5070 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1128_
timestamp 0
transform 1 0 5730 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1129_
timestamp 0
transform 1 0 5590 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1130_
timestamp 0
transform 1 0 5710 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1131_
timestamp 0
transform 1 0 5250 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1132_
timestamp 0
transform 1 0 5870 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1133_
timestamp 0
transform 1 0 5710 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1134_
timestamp 0
transform 1 0 5730 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1135_
timestamp 0
transform 1 0 5570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1136_
timestamp 0
transform 1 0 5790 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1137_
timestamp 0
transform -1 0 5690 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1138_
timestamp 0
transform -1 0 5430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1139_
timestamp 0
transform 1 0 5210 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1140_
timestamp 0
transform 1 0 5550 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1141_
timestamp 0
transform 1 0 5370 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1142_
timestamp 0
transform 1 0 5510 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1143_
timestamp 0
transform -1 0 5730 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1144_
timestamp 0
transform -1 0 5410 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1145_
timestamp 0
transform 1 0 5290 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1146_
timestamp 0
transform 1 0 4610 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1147_
timestamp 0
transform -1 0 3990 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1148_
timestamp 0
transform -1 0 5190 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1149_
timestamp 0
transform -1 0 5030 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1150_
timestamp 0
transform 1 0 4610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1151_
timestamp 0
transform 1 0 4430 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1152_
timestamp 0
transform -1 0 5290 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1153_
timestamp 0
transform -1 0 3150 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1154_
timestamp 0
transform -1 0 3530 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1155_
timestamp 0
transform 1 0 4030 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1156_
timestamp 0
transform -1 0 3450 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1157_
timestamp 0
transform 1 0 3570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1158_
timestamp 0
transform 1 0 3270 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1159_
timestamp 0
transform 1 0 4410 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1160_
timestamp 0
transform 1 0 4310 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1161_
timestamp 0
transform -1 0 4270 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1162_
timestamp 0
transform 1 0 3590 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1163_
timestamp 0
transform -1 0 3770 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1164_
timestamp 0
transform -1 0 4790 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1165_
timestamp 0
transform 1 0 4930 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1166_
timestamp 0
transform -1 0 4290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1167_
timestamp 0
transform -1 0 4610 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1168_
timestamp 0
transform -1 0 4930 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1169_
timestamp 0
transform 1 0 4430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1170_
timestamp 0
transform -1 0 4330 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1171_
timestamp 0
transform 1 0 4710 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1172_
timestamp 0
transform 1 0 4550 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1173_
timestamp 0
transform 1 0 4750 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1174_
timestamp 0
transform 1 0 4890 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1175_
timestamp 0
transform 1 0 5050 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1176_
timestamp 0
transform -1 0 5110 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1177_
timestamp 0
transform 1 0 5230 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1178_
timestamp 0
transform 1 0 5830 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1179_
timestamp 0
transform -1 0 5770 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1180_
timestamp 0
transform 1 0 5590 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1181_
timestamp 0
transform -1 0 5450 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1182_
timestamp 0
transform -1 0 4830 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1183_
timestamp 0
transform 1 0 4150 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1184_
timestamp 0
transform -1 0 4310 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1185_
timestamp 0
transform -1 0 1370 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1186_
timestamp 0
transform 1 0 5490 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1187_
timestamp 0
transform -1 0 5370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1188_
timestamp 0
transform 1 0 5770 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1189_
timestamp 0
transform 1 0 5630 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1190_
timestamp 0
transform -1 0 5690 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1191_
timestamp 0
transform 1 0 5190 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1192_
timestamp 0
transform -1 0 4490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1193_
timestamp 0
transform -1 0 4130 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1194_
timestamp 0
transform 1 0 5470 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1195_
timestamp 0
transform 1 0 5250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1196_
timestamp 0
transform -1 0 4070 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1197_
timestamp 0
transform -1 0 3890 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1198_
timestamp 0
transform 1 0 3910 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1199_
timestamp 0
transform 1 0 3790 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1200_
timestamp 0
transform 1 0 3890 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1201_
timestamp 0
transform -1 0 4630 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1202_
timestamp 0
transform 1 0 4770 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1203_
timestamp 0
transform 1 0 5410 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1204_
timestamp 0
transform 1 0 5310 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1205_
timestamp 0
transform 1 0 5290 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1206_
timestamp 0
transform 1 0 5130 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1207_
timestamp 0
transform -1 0 5170 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1208_
timestamp 0
transform -1 0 5010 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1209_
timestamp 0
transform -1 0 5010 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1210_
timestamp 0
transform 1 0 4850 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1211_
timestamp 0
transform 1 0 4790 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1212_
timestamp 0
transform -1 0 4750 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1213_
timestamp 0
transform 1 0 3990 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1214_
timestamp 0
transform -1 0 4950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1215_
timestamp 0
transform 1 0 4130 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1216_
timestamp 0
transform -1 0 5410 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1217_
timestamp 0
transform 1 0 5230 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1218_
timestamp 0
transform -1 0 4650 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1219_
timestamp 0
transform 1 0 1730 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1220_
timestamp 0
transform 1 0 650 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1221_
timestamp 0
transform 1 0 5130 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1222_
timestamp 0
transform 1 0 4130 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1223_
timestamp 0
transform 1 0 3950 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1224_
timestamp 0
transform 1 0 3430 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1225_
timestamp 0
transform 1 0 3730 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1226_
timestamp 0
transform -1 0 3750 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1227_
timestamp 0
transform 1 0 3850 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1228_
timestamp 0
transform -1 0 3590 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1229_
timestamp 0
transform -1 0 4270 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1230_
timestamp 0
transform 1 0 4930 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1231_
timestamp 0
transform 1 0 4710 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1232_
timestamp 0
transform -1 0 4570 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1233_
timestamp 0
transform -1 0 4710 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1234_
timestamp 0
transform -1 0 4570 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1235_
timestamp 0
transform -1 0 4410 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1236_
timestamp 0
transform 1 0 790 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1237_
timestamp 0
transform -1 0 4390 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1238_
timestamp 0
transform 1 0 5730 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1239_
timestamp 0
transform 1 0 5290 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1240_
timestamp 0
transform -1 0 5470 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1241_
timestamp 0
transform 1 0 4830 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1242_
timestamp 0
transform 1 0 4910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1243_
timestamp 0
transform -1 0 3970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1244_
timestamp 0
transform 1 0 3610 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1245_
timestamp 0
transform -1 0 3810 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1246_
timestamp 0
transform 1 0 4010 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1247_
timestamp 0
transform 1 0 4090 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1248_
timestamp 0
transform 1 0 4130 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1249_
timestamp 0
transform 1 0 4650 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1250_
timestamp 0
transform 1 0 5070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1251_
timestamp 0
transform -1 0 5530 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1252_
timestamp 0
transform -1 0 5090 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1253_
timestamp 0
transform 1 0 4790 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1254_
timestamp 0
transform 1 0 4910 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1255_
timestamp 0
transform 1 0 4730 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1256_
timestamp 0
transform -1 0 4290 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1257_
timestamp 0
transform -1 0 4470 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1258_
timestamp 0
transform 1 0 4290 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1259_
timestamp 0
transform 1 0 4450 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1260_
timestamp 0
transform 1 0 1790 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1261_
timestamp 0
transform 1 0 1230 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1262_
timestamp 0
transform -1 0 1550 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1263_
timestamp 0
transform -1 0 1410 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1264_
timestamp 0
transform -1 0 950 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1265_
timestamp 0
transform -1 0 1330 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1266_
timestamp 0
transform -1 0 1470 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1267_
timestamp 0
transform -1 0 1330 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1268_
timestamp 0
transform -1 0 1290 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1269_
timestamp 0
transform -1 0 990 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1270_
timestamp 0
transform -1 0 1110 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1271_
timestamp 0
transform 1 0 1110 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1272_
timestamp 0
transform -1 0 970 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1273_
timestamp 0
transform 1 0 630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1274_
timestamp 0
transform -1 0 810 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1275_
timestamp 0
transform -1 0 1170 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1276_
timestamp 0
transform -1 0 810 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1277_
timestamp 0
transform 1 0 590 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1278_
timestamp 0
transform -1 0 470 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1279_
timestamp 0
transform -1 0 610 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1280_
timestamp 0
transform 1 0 970 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1281_
timestamp 0
transform -1 0 830 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1282_
timestamp 0
transform 1 0 750 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1283_
timestamp 0
transform 1 0 890 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1284_
timestamp 0
transform 1 0 610 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1285_
timestamp 0
transform -1 0 370 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1286_
timestamp 0
transform 1 0 290 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1287_
timestamp 0
transform -1 0 310 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1288_
timestamp 0
transform 1 0 750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1289_
timestamp 0
transform 1 0 50 0 -1 5470
box -6 -8 26 268
use FILL  FILL_2__1290_
timestamp 0
transform 1 0 170 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2__1291_
timestamp 0
transform 1 0 50 0 1 5470
box -6 -8 26 268
use FILL  FILL_2__1292_
timestamp 0
transform -1 0 70 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1293_
timestamp 0
transform -1 0 610 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1294_
timestamp 0
transform -1 0 450 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1295_
timestamp 0
transform 1 0 190 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1296_
timestamp 0
transform 1 0 50 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1297_
timestamp 0
transform 1 0 170 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1298_
timestamp 0
transform 1 0 470 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1299_
timestamp 0
transform 1 0 430 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1300_
timestamp 0
transform -1 0 450 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1301_
timestamp 0
transform 1 0 310 0 1 4950
box -6 -8 26 268
use FILL  FILL_2__1302_
timestamp 0
transform -1 0 550 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1303_
timestamp 0
transform 1 0 710 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1304_
timestamp 0
transform -1 0 390 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1305_
timestamp 0
transform -1 0 490 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1306_
timestamp 0
transform -1 0 330 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2__1307_
timestamp 0
transform 1 0 190 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1308_
timestamp 0
transform 1 0 310 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1309_
timestamp 0
transform 1 0 510 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1310_
timestamp 0
transform 1 0 290 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1311_
timestamp 0
transform -1 0 70 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1312_
timestamp 0
transform -1 0 430 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1313_
timestamp 0
transform -1 0 70 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1314_
timestamp 0
transform -1 0 210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1315_
timestamp 0
transform -1 0 230 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1316_
timestamp 0
transform 1 0 50 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1317_
timestamp 0
transform -1 0 350 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1318_
timestamp 0
transform -1 0 1210 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1319_
timestamp 0
transform 1 0 1230 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1320_
timestamp 0
transform -1 0 1130 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1321_
timestamp 0
transform -1 0 930 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1322_
timestamp 0
transform -1 0 230 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1323_
timestamp 0
transform 1 0 290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1324_
timestamp 0
transform -1 0 310 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1325_
timestamp 0
transform 1 0 1730 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1326_
timestamp 0
transform 1 0 210 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1327_
timestamp 0
transform 1 0 810 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1328_
timestamp 0
transform 1 0 950 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1329_
timestamp 0
transform -1 0 70 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1330_
timestamp 0
transform 1 0 610 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1331_
timestamp 0
transform -1 0 70 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1332_
timestamp 0
transform 1 0 610 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1333_
timestamp 0
transform 1 0 770 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1334_
timestamp 0
transform -1 0 2630 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1335_
timestamp 0
transform 1 0 2770 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1336_
timestamp 0
transform -1 0 2470 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1337_
timestamp 0
transform -1 0 2210 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1338_
timestamp 0
transform 1 0 2190 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1339_
timestamp 0
transform -1 0 2350 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1340_
timestamp 0
transform -1 0 2050 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1341_
timestamp 0
transform -1 0 1890 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1342_
timestamp 0
transform 1 0 2390 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1343_
timestamp 0
transform 1 0 3470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1344_
timestamp 0
transform 1 0 3610 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1345_
timestamp 0
transform 1 0 2990 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1346_
timestamp 0
transform 1 0 2830 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1347_
timestamp 0
transform -1 0 2570 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1348_
timestamp 0
transform -1 0 2210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1349_
timestamp 0
transform -1 0 1370 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1350_
timestamp 0
transform -1 0 1750 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1351_
timestamp 0
transform -1 0 470 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1352_
timestamp 0
transform -1 0 2070 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1353_
timestamp 0
transform -1 0 2690 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1354_
timestamp 0
transform -1 0 1910 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1355_
timestamp 0
transform -1 0 1230 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1356_
timestamp 0
transform -1 0 1090 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1357_
timestamp 0
transform -1 0 810 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1358_
timestamp 0
transform 1 0 670 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1359_
timestamp 0
transform 1 0 590 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1360_
timestamp 0
transform 1 0 930 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1361_
timestamp 0
transform -1 0 770 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1362_
timestamp 0
transform -1 0 550 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1363_
timestamp 0
transform -1 0 270 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1364_
timestamp 0
transform 1 0 190 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1365_
timestamp 0
transform 1 0 170 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1366_
timestamp 0
transform -1 0 70 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1367_
timestamp 0
transform -1 0 70 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1368_
timestamp 0
transform -1 0 70 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1369_
timestamp 0
transform 1 0 210 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1370_
timestamp 0
transform -1 0 70 0 -1 1310
box -6 -8 26 268
use FILL  FILL_2__1371_
timestamp 0
transform -1 0 2850 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1372_
timestamp 0
transform 1 0 330 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1373_
timestamp 0
transform -1 0 410 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1374_
timestamp 0
transform -1 0 510 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1375_
timestamp 0
transform -1 0 3990 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1376_
timestamp 0
transform 1 0 4110 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1377_
timestamp 0
transform -1 0 3710 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1378_
timestamp 0
transform 1 0 3810 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1379_
timestamp 0
transform -1 0 2990 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1380_
timestamp 0
transform -1 0 3170 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1381_
timestamp 0
transform 1 0 3270 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1382_
timestamp 0
transform -1 0 3130 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1383_
timestamp 0
transform -1 0 2990 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1384_
timestamp 0
transform 1 0 3530 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1385_
timestamp 0
transform 1 0 4250 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1386_
timestamp 0
transform -1 0 4010 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1387_
timestamp 0
transform -1 0 3870 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1388_
timestamp 0
transform 1 0 3890 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1389_
timestamp 0
transform -1 0 3570 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1390_
timestamp 0
transform 1 0 3710 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1391_
timestamp 0
transform 1 0 3370 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1392_
timestamp 0
transform -1 0 3710 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1393_
timestamp 0
transform -1 0 3590 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1394_
timestamp 0
transform -1 0 3410 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1395_
timestamp 0
transform -1 0 3290 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1396_
timestamp 0
transform -1 0 2610 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1397_
timestamp 0
transform 1 0 2290 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1398_
timestamp 0
transform 1 0 2710 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1399_
timestamp 0
transform 1 0 2250 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1400_
timestamp 0
transform -1 0 1770 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1401_
timestamp 0
transform -1 0 2150 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1402_
timestamp 0
transform -1 0 2450 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1403_
timestamp 0
transform -1 0 2010 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1404_
timestamp 0
transform -1 0 1910 0 1 790
box -6 -8 26 268
use FILL  FILL_2__1405_
timestamp 0
transform -1 0 3450 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1406_
timestamp 0
transform 1 0 1470 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1407_
timestamp 0
transform 1 0 3510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1408_
timestamp 0
transform 1 0 3350 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2__1409_
timestamp 0
transform 1 0 3350 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1410_
timestamp 0
transform -1 0 3650 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1411_
timestamp 0
transform 1 0 3470 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1412_
timestamp 0
transform 1 0 2870 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1413_
timestamp 0
transform 1 0 2970 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1414_
timestamp 0
transform 1 0 2990 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1415_
timestamp 0
transform 1 0 1870 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1416_
timestamp 0
transform -1 0 1530 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1417_
timestamp 0
transform 1 0 1470 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1418_
timestamp 0
transform -1 0 890 0 1 1310
box -6 -8 26 268
use FILL  FILL_2__1419_
timestamp 0
transform 1 0 3110 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1420_
timestamp 0
transform 1 0 3250 0 1 2350
box -6 -8 26 268
use FILL  FILL_2__1421_
timestamp 0
transform -1 0 3050 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1422_
timestamp 0
transform 1 0 3170 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1423_
timestamp 0
transform -1 0 2450 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1424_
timestamp 0
transform -1 0 2830 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1425_
timestamp 0
transform 1 0 1170 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1426_
timestamp 0
transform -1 0 1330 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1427_
timestamp 0
transform 1 0 1910 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1428_
timestamp 0
transform -1 0 2190 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1429_
timestamp 0
transform -1 0 2350 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1430_
timestamp 0
transform 1 0 2410 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1431_
timestamp 0
transform -1 0 2750 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1432_
timestamp 0
transform 1 0 2090 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1433_
timestamp 0
transform -1 0 2270 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1434_
timestamp 0
transform -1 0 2250 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1435_
timestamp 0
transform 1 0 2070 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1436_
timestamp 0
transform -1 0 2230 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1437_
timestamp 0
transform -1 0 2610 0 1 1830
box -6 -8 26 268
use FILL  FILL_2__1438_
timestamp 0
transform -1 0 2570 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1439_
timestamp 0
transform -1 0 2710 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1440_
timestamp 0
transform -1 0 2510 0 1 2870
box -6 -8 26 268
use FILL  FILL_2__1441_
timestamp 0
transform 1 0 2570 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2__1442_
timestamp 0
transform -1 0 1510 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1443_
timestamp 0
transform 1 0 1630 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2__1444_
timestamp 0
transform -1 0 2670 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1445_
timestamp 0
transform -1 0 2810 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1446_
timestamp 0
transform -1 0 3110 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1447_
timestamp 0
transform -1 0 3130 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1448_
timestamp 0
transform -1 0 3250 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2__1449_
timestamp 0
transform -1 0 3530 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1450_
timestamp 0
transform -1 0 2430 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1451_
timestamp 0
transform -1 0 2690 0 1 3390
box -6 -8 26 268
use FILL  FILL_2__1527_
timestamp 0
transform 1 0 5530 0 1 270
box -6 -8 26 268
use FILL  FILL_2__1528_
timestamp 0
transform 1 0 3630 0 -1 3390
box -6 -8 26 268
use FILL  FILL_2__1529_
timestamp 0
transform 1 0 4530 0 1 3910
box -6 -8 26 268
use FILL  FILL_2__1530_
timestamp 0
transform 1 0 5390 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2__1531_
timestamp 0
transform 1 0 5870 0 1 4430
box -6 -8 26 268
use FILL  FILL_2__1532_
timestamp 0
transform 1 0 930 0 -1 790
box -6 -8 26 268
use FILL  FILL_2__1533_
timestamp 0
transform -1 0 470 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1534_
timestamp 0
transform -1 0 330 0 -1 270
box -6 -8 26 268
use FILL  FILL_2__1535_
timestamp 0
transform -1 0 70 0 1 790
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert0
timestamp 0
transform -1 0 1070 0 1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert1
timestamp 0
transform 1 0 2990 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert2
timestamp 0
transform -1 0 1110 0 1 790
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert3
timestamp 0
transform -1 0 1010 0 1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert4
timestamp 0
transform 1 0 1610 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert5
timestamp 0
transform -1 0 2310 0 1 790
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert6
timestamp 0
transform 1 0 2970 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert15
timestamp 0
transform -1 0 2710 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert16
timestamp 0
transform -1 0 2890 0 -1 4950
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert17
timestamp 0
transform -1 0 3990 0 -1 4430
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert18
timestamp 0
transform 1 0 4290 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert19
timestamp 0
transform -1 0 490 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert20
timestamp 0
transform 1 0 1110 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert21
timestamp 0
transform -1 0 470 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert22
timestamp 0
transform -1 0 850 0 1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert23
timestamp 0
transform 1 0 2310 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert24
timestamp 0
transform 1 0 2750 0 1 1830
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert25
timestamp 0
transform 1 0 3250 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert26
timestamp 0
transform -1 0 3150 0 -1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert27
timestamp 0
transform -1 0 2870 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert28
timestamp 0
transform -1 0 2890 0 1 2870
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert29
timestamp 0
transform 1 0 1350 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert30
timestamp 0
transform 1 0 4670 0 1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert31
timestamp 0
transform -1 0 2990 0 1 3910
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert32
timestamp 0
transform 1 0 4650 0 1 3390
box -6 -8 26 268
use FILL  FILL_2_BUFX2_insert33
timestamp 0
transform -1 0 2830 0 1 3910
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert7
timestamp 0
transform 1 0 790 0 -1 5990
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert8
timestamp 0
transform -1 0 70 0 -1 1830
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert9
timestamp 0
transform 1 0 2290 0 -1 2350
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert10
timestamp 0
transform -1 0 70 0 1 1830
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert11
timestamp 0
transform 1 0 190 0 1 790
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert12
timestamp 0
transform 1 0 2310 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert13
timestamp 0
transform 1 0 1890 0 -1 3910
box -6 -8 26 268
use FILL  FILL_2_CLKBUF1_insert14
timestamp 0
transform 1 0 2570 0 1 790
box -6 -8 26 268
use FILL  FILL_3__726_
timestamp 0
transform -1 0 1350 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__740_
timestamp 0
transform -1 0 470 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__755_
timestamp 0
transform -1 0 3690 0 1 2870
box -6 -8 26 268
use FILL  FILL_3__770_
timestamp 0
transform 1 0 1830 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__784_
timestamp 0
transform 1 0 690 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__799_
timestamp 0
transform 1 0 850 0 -1 270
box -6 -8 26 268
use FILL  FILL_3__814_
timestamp 0
transform -1 0 2130 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__828_
timestamp 0
transform -1 0 1950 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__843_
timestamp 0
transform 1 0 1250 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__858_
timestamp 0
transform -1 0 1690 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__872_
timestamp 0
transform -1 0 1410 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__887_
timestamp 0
transform -1 0 2610 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__901_
timestamp 0
transform 1 0 3010 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__916_
timestamp 0
transform 1 0 1090 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__931_
timestamp 0
transform 1 0 3350 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__945_
timestamp 0
transform -1 0 4170 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__960_
timestamp 0
transform -1 0 2910 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__975_
timestamp 0
transform -1 0 3550 0 -1 5470
box -6 -8 26 268
use FILL  FILL_3__989_
timestamp 0
transform -1 0 4450 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1009_
timestamp 0
transform 1 0 5550 0 -1 4950
box -6 -8 26 268
use FILL  FILL_3__1024_
timestamp 0
transform 1 0 2290 0 -1 5990
box -6 -8 26 268
use FILL  FILL_3__1039_
timestamp 0
transform -1 0 5610 0 1 4950
box -6 -8 26 268
use FILL  FILL_3__1053_
timestamp 0
transform 1 0 5210 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1068_
timestamp 0
transform 1 0 4690 0 -1 3390
box -6 -8 26 268
use FILL  FILL_3__1083_
timestamp 0
transform -1 0 5730 0 1 5470
box -6 -8 26 268
use FILL  FILL_3__1097_
timestamp 0
transform 1 0 3830 0 1 1310
box -6 -8 26 268
use FILL  FILL_3__1112_
timestamp 0
transform 1 0 4570 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1127_
timestamp 0
transform 1 0 5090 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1141_
timestamp 0
transform 1 0 5390 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1156_
timestamp 0
transform -1 0 3470 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1171_
timestamp 0
transform 1 0 4730 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1185_
timestamp 0
transform -1 0 1390 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1200_
timestamp 0
transform 1 0 3910 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1215_
timestamp 0
transform 1 0 4150 0 1 1830
box -6 -8 26 268
use FILL  FILL_3__1229_
timestamp 0
transform -1 0 4290 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3__1244_
timestamp 0
transform 1 0 3630 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1259_
timestamp 0
transform 1 0 4470 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1273_
timestamp 0
transform 1 0 650 0 -1 2350
box -6 -8 26 268
use FILL  FILL_3__1288_
timestamp 0
transform 1 0 770 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1302_
timestamp 0
transform -1 0 570 0 1 4430
box -6 -8 26 268
use FILL  FILL_3__1317_
timestamp 0
transform -1 0 370 0 -1 3910
box -6 -8 26 268
use FILL  FILL_3__1332_
timestamp 0
transform 1 0 630 0 -1 4430
box -6 -8 26 268
use FILL  FILL_3__1346_
timestamp 0
transform 1 0 2850 0 -1 1310
box -6 -8 26 268
use FILL  FILL_3__1361_
timestamp 0
transform -1 0 790 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1376_
timestamp 0
transform 1 0 4130 0 -1 790
box -6 -8 26 268
use FILL  FILL_3__1390_
timestamp 0
transform 1 0 3730 0 1 790
box -6 -8 26 268
use FILL  FILL_3__1405_
timestamp 0
transform -1 0 3470 0 1 270
box -6 -8 26 268
use FILL  FILL_3__1420_
timestamp 0
transform 1 0 3270 0 1 2350
box -6 -8 26 268
use FILL  FILL_3__1434_
timestamp 0
transform -1 0 2270 0 -1 2870
box -6 -8 26 268
use FILL  FILL_3__1449_
timestamp 0
transform -1 0 3550 0 1 3910
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert4
timestamp 0
transform 1 0 1630 0 1 3390
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert19
timestamp 0
transform -1 0 510 0 -1 1830
box -6 -8 26 268
use FILL  FILL_3_BUFX2_insert33
timestamp 0
transform -1 0 2850 0 1 3910
box -6 -8 26 268
<< labels >>
flabel metal1 s 5983 2 6043 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 4876 6036 4884 6044 3 FreeSans 16 90 0 0 Cin[5]
port 2 nsew
flabel metal2 s 4836 6036 4844 6044 3 FreeSans 16 90 0 0 Cin[4]
port 3 nsew
flabel metal2 s 4736 6036 4744 6044 3 FreeSans 16 90 0 0 Cin[3]
port 4 nsew
flabel metal2 s 4696 6036 4704 6044 3 FreeSans 16 90 0 0 Cin[2]
port 5 nsew
flabel metal2 s 3536 6036 3544 6044 3 FreeSans 16 90 0 0 Cin[1]
port 6 nsew
flabel metal2 s 2936 6036 2944 6044 3 FreeSans 16 90 0 0 Cin[0]
port 7 nsew
flabel metal3 s -24 2216 -16 2224 7 FreeSans 16 0 0 0 Rdy
port 8 nsew
flabel metal3 s 6016 396 6024 404 3 FreeSans 16 0 0 0 Vld
port 9 nsew
flabel metal3 s -24 3856 -16 3864 7 FreeSans 16 0 0 0 Xin[3]
port 10 nsew
flabel metal3 s -24 3816 -16 3824 7 FreeSans 16 0 0 0 Xin[2]
port 11 nsew
flabel metal3 s -24 3776 -16 3784 7 FreeSans 16 0 0 0 Xin[1]
port 12 nsew
flabel metal3 s -24 2996 -16 3004 7 FreeSans 16 0 0 0 Xin[0]
port 13 nsew
flabel metal3 s 6016 4556 6024 4564 3 FreeSans 16 0 0 0 Xout[3]
port 14 nsew
flabel metal3 s 6016 4296 6024 4304 3 FreeSans 16 0 0 0 Xout[2]
port 15 nsew
flabel metal3 s 6016 4036 6024 4044 3 FreeSans 16 0 0 0 Xout[1]
port 16 nsew
flabel metal3 s 6016 3256 6024 3264 3 FreeSans 16 0 0 0 Xout[0]
port 17 nsew
flabel metal2 s 1916 -24 1924 -16 7 FreeSans 16 270 0 0 Yin[3]
port 18 nsew
flabel metal2 s 2916 -24 2924 -16 7 FreeSans 16 270 0 0 Yin[2]
port 19 nsew
flabel metal2 s 3396 -24 3404 -16 7 FreeSans 16 270 0 0 Yin[1]
port 20 nsew
flabel metal2 s 3496 -24 3504 -16 7 FreeSans 16 270 0 0 Yin[0]
port 21 nsew
flabel metal2 s 96 -24 104 -16 7 FreeSans 16 270 0 0 Yout[3]
port 22 nsew
flabel metal2 s 356 -24 364 -16 7 FreeSans 16 270 0 0 Yout[2]
port 23 nsew
flabel metal2 s 496 -24 504 -16 7 FreeSans 16 270 0 0 Yout[1]
port 24 nsew
flabel metal2 s 976 -24 984 -16 7 FreeSans 16 270 0 0 Yout[0]
port 25 nsew
flabel metal2 s 816 6036 824 6044 3 FreeSans 16 90 0 0 clk
port 26 nsew
<< properties >>
string FIXED_BBOX -40 -40 6020 6040
<< end >>
