* NGSPICE file created from cpu.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A Y vdd gnd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR D S R CLK Q vdd gnd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A Y vdd gnd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A Y vdd gnd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 D CLK Q vdd gnd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A Y vdd gnd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S Y vdd gnd
.ends

.subckt cpu gnd vdd AB[15] AB[14] AB[13] AB[12] AB[11] AB[10] AB[9] AB[8] AB[7] AB[6]
+ AB[5] AB[4] AB[3] AB[2] AB[1] AB[0] DI[7] DI[6] DI[5] DI[4] DI[3] DI[2] DI[1] DI[0]
+ DO[7] DO[6] DO[5] DO[4] DO[3] DO[2] DO[1] DO[0] IRQ NMI RDY WE clk reset
XFILL_0__2877_ gnd vdd FILL
XFILL_3__2586_ gnd vdd FILL
XFILL_6__2295_ gnd vdd FILL
X_3155_ _3196_/A _3170_/B vdd gnd INVX1
XFILL_0__1828_ gnd vdd FILL
XFILL_0__1759_ gnd vdd FILL
X_3086_ _3086_/A _3577_/Q _3087_/B vdd gnd XOR2X1
X_2106_ _2294_/A _2441_/B _2106_/C _2107_/B vdd gnd OAI21X1
X_2037_ _2922_/A _2931_/A vdd gnd INVX1
XFILL_4__2000_ gnd vdd FILL
XFILL_3__3207_ gnd vdd FILL
XFILL_0__3429_ gnd vdd FILL
XFILL_1__2222_ gnd vdd FILL
XFILL_3__3138_ gnd vdd FILL
XFILL_7__1990_ gnd vdd FILL
XFILL_3__3069_ gnd vdd FILL
XFILL_1__2153_ gnd vdd FILL
X_2939_ reset _2957_/C _2940_/A vdd gnd NOR2X1
XFILL_1__2084_ gnd vdd FILL
XFILL_4__2902_ gnd vdd FILL
XFILL_7__2611_ gnd vdd FILL
XFILL_4__2833_ gnd vdd FILL
XFILL_7__3591_ gnd vdd FILL
XFILL_9__3458_ gnd vdd FILL
XFILL_7__2542_ gnd vdd FILL
XFILL_4__2764_ gnd vdd FILL
XFILL_8_CLKBUF1_insert33 gnd vdd FILL
XFILL_1__2986_ gnd vdd FILL
XFILL_7__2473_ gnd vdd FILL
XFILL_4__1715_ gnd vdd FILL
XFILL_1__1937_ gnd vdd FILL
XFILL_4__2695_ gnd vdd FILL
XFILL_1__1868_ gnd vdd FILL
XFILL_2__3380_ gnd vdd FILL
XFILL_2__2400_ gnd vdd FILL
XFILL_1__1799_ gnd vdd FILL
XFILL_1__3538_ gnd vdd FILL
XFILL_2__2331_ gnd vdd FILL
XFILL_7__3025_ gnd vdd FILL
XFILL_5__2040_ gnd vdd FILL
XFILL_1__3469_ gnd vdd FILL
XFILL_2__2262_ gnd vdd FILL
XFILL_4__3178_ gnd vdd FILL
XFILL_2__2193_ gnd vdd FILL
XFILL_4__2129_ gnd vdd FILL
XFILL_8__2720_ gnd vdd FILL
XFILL_5__2942_ gnd vdd FILL
XFILL_8__2651_ gnd vdd FILL
XFILL_7__2809_ gnd vdd FILL
XFILL_5__2873_ gnd vdd FILL
XFILL_5__1824_ gnd vdd FILL
XFILL_8__2582_ gnd vdd FILL
XFILL_5__1755_ gnd vdd FILL
XFILL_2__1977_ gnd vdd FILL
XFILL_0__2800_ gnd vdd FILL
XFILL_8__3203_ gnd vdd FILL
XFILL_5__3425_ gnd vdd FILL
XFILL_0__2731_ gnd vdd FILL
XFILL_8__3134_ gnd vdd FILL
XFILL_3__2440_ gnd vdd FILL
XFILL_3__2371_ gnd vdd FILL
XFILL182250x140550 gnd vdd FILL
XFILL_8__3065_ gnd vdd FILL
XFILL_5__2307_ gnd vdd FILL
XFILL_0__2662_ gnd vdd FILL
XFILL_6__2080_ gnd vdd FILL
XFILL_8__2016_ gnd vdd FILL
XFILL_2__2529_ gnd vdd FILL
XFILL_0__2593_ gnd vdd FILL
XFILL_5__2238_ gnd vdd FILL
XFILL_5__2169_ gnd vdd FILL
XFILL_8__2918_ gnd vdd FILL
XFILL_6__2982_ gnd vdd FILL
XFILL_0__3214_ gnd vdd FILL
XFILL_4_BUFX2_insert3 gnd vdd FILL
XFILL_6__1933_ gnd vdd FILL
XFILL_0__3145_ gnd vdd FILL
XFILL_8__2849_ gnd vdd FILL
XFILL_0__3076_ gnd vdd FILL
XFILL_6__1864_ gnd vdd FILL
X_2724_ _2724_/A _2733_/B _2731_/A vdd gnd NOR2X1
XFILL_6__3603_ gnd vdd FILL
XFILL_0__2027_ gnd vdd FILL
X_2655_ _3244_/Q _2685_/B _2656_/C vdd gnd NAND2X1
XFILL_6__1795_ gnd vdd FILL
XFILL_1__2840_ gnd vdd FILL
XFILL_6__3534_ gnd vdd FILL
XFILL_6__3465_ gnd vdd FILL
X_2586_ _3176_/B _2586_/B _3178_/B _2587_/B vdd gnd NAND3X1
XFILL_6__2416_ gnd vdd FILL
XFILL_3__2707_ gnd vdd FILL
XFILL_1__2771_ gnd vdd FILL
XFILL_4__2480_ gnd vdd FILL
XFILL_0__2929_ gnd vdd FILL
XFILL_6__3396_ gnd vdd FILL
XFILL_1__1722_ gnd vdd FILL
XFILL_3__2638_ gnd vdd FILL
XFILL_6__2347_ gnd vdd FILL
X_3207_ _3215_/A _3207_/B _3207_/C _3351_/D vdd gnd OAI21X1
X_3138_ _3345_/Q _3143_/B _3139_/C vdd gnd NAND2X1
XFILL_4__3101_ gnd vdd FILL
XFILL_6__2278_ gnd vdd FILL
XFILL_3__2569_ gnd vdd FILL
XFILL_4__3032_ gnd vdd FILL
X_3069_ _3069_/A _3071_/B vdd gnd INVX1
XFILL_1__2205_ gnd vdd FILL
XFILL_7__1973_ gnd vdd FILL
XFILL_1__3185_ gnd vdd FILL
XFILL_1__2136_ gnd vdd FILL
XFILL_1__2067_ gnd vdd FILL
XFILL_2__2880_ gnd vdd FILL
XFILL_2__1900_ gnd vdd FILL
XFILL_4__2816_ gnd vdd FILL
XFILL_2__1831_ gnd vdd FILL
XFILL_7__2525_ gnd vdd FILL
XFILL_7_BUFX2_insert7 gnd vdd FILL
XFILL_4__2747_ gnd vdd FILL
XFILL_1__2969_ gnd vdd FILL
XFILL_7__2456_ gnd vdd FILL
XFILL_4__2678_ gnd vdd FILL
XFILL_2__1762_ gnd vdd FILL
XFILL_2__3501_ gnd vdd FILL
XFILL_7__2387_ gnd vdd FILL
XFILL_5__3210_ gnd vdd FILL
XFILL_2__1693_ gnd vdd FILL
XFILL_2__3432_ gnd vdd FILL
XFILL_5__3141_ gnd vdd FILL
XFILL_7__3008_ gnd vdd FILL
XFILL_5__3072_ gnd vdd FILL
XFILL_5__2023_ gnd vdd FILL
XFILL_2__2314_ gnd vdd FILL
XFILL_2__2245_ gnd vdd FILL
XFILL_2__2176_ gnd vdd FILL
XFILL_8__2703_ gnd vdd FILL
XFILL_5__2925_ gnd vdd FILL
XFILL_3__1940_ gnd vdd FILL
XFILL_8__2634_ gnd vdd FILL
XFILL_5__2856_ gnd vdd FILL
XFILL_8__2565_ gnd vdd FILL
XFILL_3__1871_ gnd vdd FILL
XFILL_5__2787_ gnd vdd FILL
XFILL_5__1807_ gnd vdd FILL
X_2440_ _3166_/B _3166_/D _2699_/B vdd gnd NAND2X1
XFILL_8__2496_ gnd vdd FILL
XFILL_5__1738_ gnd vdd FILL
X_2371_ _3273_/Q _2863_/A vdd gnd INVX1
XFILL_3__3541_ gnd vdd FILL
XFILL_3__3472_ gnd vdd FILL
XFILL_6__2201_ gnd vdd FILL
XFILL_8__3117_ gnd vdd FILL
XFILL_5__3408_ gnd vdd FILL
XFILL_3__2423_ gnd vdd FILL
XFILL_0__2714_ gnd vdd FILL
XFILL_6__3181_ gnd vdd FILL
XFILL_6__2132_ gnd vdd FILL
XFILL_0__2645_ gnd vdd FILL
XFILL_3__2354_ gnd vdd FILL
XFILL_8__3048_ gnd vdd FILL
XFILL_6__2063_ gnd vdd FILL
XFILL_0__2576_ gnd vdd FILL
XFILL_3__2285_ gnd vdd FILL
XFILL_5_BUFX2_insert61 gnd vdd FILL
XFILL_5_BUFX2_insert50 gnd vdd FILL
XFILL_5_BUFX2_insert94 gnd vdd FILL
XFILL_6__2965_ gnd vdd FILL
XFILL_4__1980_ gnd vdd FILL
XFILL_5_BUFX2_insert83 gnd vdd FILL
XFILL182850x74250 gnd vdd FILL
XFILL_5_BUFX2_insert72 gnd vdd FILL
XFILL_0__3128_ gnd vdd FILL
XFILL_6__2896_ gnd vdd FILL
XFILL_6__1916_ gnd vdd FILL
XFILL_0__3059_ gnd vdd FILL
XFILL_6__1847_ gnd vdd FILL
X_2707_ _3248_/Q _2725_/D _2725_/C _2708_/D vdd gnd NAND3X1
XFILL_6__3517_ gnd vdd FILL
XFILL_7__2310_ gnd vdd FILL
XFILL_6__1778_ gnd vdd FILL
XFILL_4__3581_ gnd vdd FILL
XFILL_4__2601_ gnd vdd FILL
X_2638_ _2638_/A _2638_/B _2638_/C _2638_/D _2639_/C vdd gnd AOI22X1
XFILL_1__2823_ gnd vdd FILL
XFILL_4__2532_ gnd vdd FILL
X_2569_ _2569_/A _2569_/B _3297_/D _2570_/C vdd gnd OAI21X1
XFILL_6__3448_ gnd vdd FILL
XFILL_7__2241_ gnd vdd FILL
XFILL_1__2754_ gnd vdd FILL
XFILL_6__3379_ gnd vdd FILL
XFILL_7__2172_ gnd vdd FILL
XFILL_1__1705_ gnd vdd FILL
XFILL_4__2463_ gnd vdd FILL
XFILL_4__2394_ gnd vdd FILL
XFILL_1__2685_ gnd vdd FILL
XFILL_4__3015_ gnd vdd FILL
XFILL_2__2030_ gnd vdd FILL
XFILL_7__1956_ gnd vdd FILL
XFILL_1__3168_ gnd vdd FILL
XFILL_1__3099_ gnd vdd FILL
XFILL_7__1887_ gnd vdd FILL
XFILL_1__2119_ gnd vdd FILL
XFILL_5__2710_ gnd vdd FILL
XFILL_2__2932_ gnd vdd FILL
XFILL_5__2641_ gnd vdd FILL
XFILL_2__2863_ gnd vdd FILL
XFILL_7__3557_ gnd vdd FILL
XFILL_8__2350_ gnd vdd FILL
XFILL_5__2572_ gnd vdd FILL
XFILL_7__3488_ gnd vdd FILL
XFILL_2__2794_ gnd vdd FILL
XFILL_8__2281_ gnd vdd FILL
XFILL_2__1814_ gnd vdd FILL
XFILL_7__2508_ gnd vdd FILL
XFILL_2__1745_ gnd vdd FILL
XFILL_7__2439_ gnd vdd FILL
XFILL_5__3124_ gnd vdd FILL
XFILL_2__3415_ gnd vdd FILL
XFILL_0__2430_ gnd vdd FILL
XFILL_0__2361_ gnd vdd FILL
XFILL_5__3055_ gnd vdd FILL
XFILL_5__2006_ gnd vdd FILL
XFILL_3__2070_ gnd vdd FILL
X_1940_ _3318_/Q _3029_/B _1941_/B vdd gnd NAND2X1
XFILL_2__2228_ gnd vdd FILL
XFILL_8__1996_ gnd vdd FILL
XFILL_0__2292_ gnd vdd FILL
X_1871_ _1871_/A _1872_/C vdd gnd INVX1
XFILL_2__2159_ gnd vdd FILL
XFILL182850x148350 gnd vdd FILL
XFILL_6__2750_ gnd vdd FILL
XFILL_5__2908_ gnd vdd FILL
XFILL_3__2972_ gnd vdd FILL
X_3541_ _3553_/B _3555_/B _3541_/C _3569_/D vdd gnd OAI21X1
XFILL_6__1701_ gnd vdd FILL
XFILL_6__2681_ gnd vdd FILL
XFILL_8__2617_ gnd vdd FILL
XFILL_5__2839_ gnd vdd FILL
XFILL_8__3597_ gnd vdd FILL
XFILL_3__1923_ gnd vdd FILL
X_3472_ _3472_/A _3472_/B _3473_/C vdd gnd NAND2X1
XFILL184350x124950 gnd vdd FILL
XFILL_3__1854_ gnd vdd FILL
XFILL_8__2548_ gnd vdd FILL
X_2423_ _2423_/A _2515_/A _2428_/C vdd gnd NAND2X1
XFILL_8__2479_ gnd vdd FILL
X_2354_ _3270_/Q _2837_/A vdd gnd INVX1
XFILL_3__1785_ gnd vdd FILL
XFILL_3__3524_ gnd vdd FILL
XFILL_3__3455_ gnd vdd FILL
X_2285_ _2285_/A _2285_/B _2286_/C vdd gnd AND2X2
XFILL_3__3386_ gnd vdd FILL
XFILL_1__2470_ gnd vdd FILL
XFILL_6__3164_ gnd vdd FILL
XFILL_3__2406_ gnd vdd FILL
XFILL_6__3095_ gnd vdd FILL
XFILL_3__2337_ gnd vdd FILL
XFILL_6__2115_ gnd vdd FILL
XFILL_0__2628_ gnd vdd FILL
XBUFX2_insert0 _1773_/Y _3166_/B vdd gnd BUFX2
XFILL_6__2046_ gnd vdd FILL
XFILL_0__2559_ gnd vdd FILL
XFILL_3__2268_ gnd vdd FILL
XFILL_3__2199_ gnd vdd FILL
XFILL_7__2790_ gnd vdd FILL
XFILL_1__3022_ gnd vdd FILL
XFILL_7__1810_ gnd vdd FILL
XFILL_6__2948_ gnd vdd FILL
XFILL_7__1741_ gnd vdd FILL
XFILL_4__1963_ gnd vdd FILL
XFILL_7__3411_ gnd vdd FILL
XFILL_6__2879_ gnd vdd FILL
XFILL_4__1894_ gnd vdd FILL
XFILL_1__2806_ gnd vdd FILL
XFILL_4__3564_ gnd vdd FILL
XFILL_9__3209_ gnd vdd FILL
XFILL_4__3495_ gnd vdd FILL
XFILL_7__2224_ gnd vdd FILL
XFILL_4__2515_ gnd vdd FILL
XFILL_3_CLKBUF1_insert34 gnd vdd FILL
XFILL_4__2446_ gnd vdd FILL
XFILL_1__2737_ gnd vdd FILL
XFILL_1_BUFX2_insert70 gnd vdd FILL
XFILL_1_BUFX2_insert92 gnd vdd FILL
XFILL_7__2155_ gnd vdd FILL
XFILL_1_BUFX2_insert81 gnd vdd FILL
XFILL_1__2668_ gnd vdd FILL
XFILL_7__2086_ gnd vdd FILL
XFILL_4__2377_ gnd vdd FILL
XFILL_2__3200_ gnd vdd FILL
XFILL_2__3131_ gnd vdd FILL
XFILL_1__2599_ gnd vdd FILL
XFILL_2__3062_ gnd vdd FILL
XFILL_8__1850_ gnd vdd FILL
XFILL_2__2013_ gnd vdd FILL
XFILL_7__2988_ gnd vdd FILL
XFILL_8__1781_ gnd vdd FILL
XFILL_7__1939_ gnd vdd FILL
XFILL_8__3520_ gnd vdd FILL
XFILL_8__3451_ gnd vdd FILL
XFILL_2__2915_ gnd vdd FILL
XFILL_8__3382_ gnd vdd FILL
XFILL_8__2402_ gnd vdd FILL
XFILL_0__1930_ gnd vdd FILL
XFILL_8__2333_ gnd vdd FILL
XFILL_5__2624_ gnd vdd FILL
XFILL_2__2846_ gnd vdd FILL
XFILL_0__1861_ gnd vdd FILL
XFILL_5__2555_ gnd vdd FILL
XFILL_8__2264_ gnd vdd FILL
XFILL_0__3600_ gnd vdd FILL
XFILL_2__2777_ gnd vdd FILL
XFILL_8__2195_ gnd vdd FILL
XFILL_0__1792_ gnd vdd FILL
XFILL_5__2486_ gnd vdd FILL
XFILL_2__1728_ gnd vdd FILL
XFILL_0__3531_ gnd vdd FILL
X_2070_ _2958_/A _3173_/B _2242_/A _2347_/B vdd gnd OAI21X1
XFILL_0__3462_ gnd vdd FILL
XFILL_5__3107_ gnd vdd FILL
XFILL_3__3171_ gnd vdd FILL
XFILL_0__2413_ gnd vdd FILL
XFILL_0__3393_ gnd vdd FILL
XFILL_5__3038_ gnd vdd FILL
XFILL_3__2122_ gnd vdd FILL
X_2972_ _3260_/Q _3264_/Q _2973_/B vdd gnd NOR2X1
XFILL_0__2344_ gnd vdd FILL
XFILL_3__2053_ gnd vdd FILL
XFILL_0__2275_ gnd vdd FILL
X_1923_ _3219_/A _2700_/B _2527_/C vdd gnd NOR2X1
XFILL_8__1979_ gnd vdd FILL
XFILL184350x136650 gnd vdd FILL
XFILL_6__2802_ gnd vdd FILL
X_1854_ _1883_/A _1863_/B _1862_/B vdd gnd NOR2X1
XFILL_6__2733_ gnd vdd FILL
XFILL_3__2955_ gnd vdd FILL
X_1785_ _2221_/A _3156_/B _3192_/A _3194_/A vdd gnd OAI21X1
X_3524_ _3524_/A _3537_/C vdd gnd INVX1
XFILL_1__1970_ gnd vdd FILL
XFILL_6__2664_ gnd vdd FILL
XFILL_3__1906_ gnd vdd FILL
X_3455_ _3484_/B _3469_/B _3455_/C _3471_/A _3461_/A vdd gnd AOI22X1
XFILL_3__2886_ gnd vdd FILL
XFILL_6__2595_ gnd vdd FILL
XFILL_3__1837_ gnd vdd FILL
X_2406_ _2795_/A _2409_/C _2717_/C _2406_/D _2407_/C vdd gnd OAI22X1
X_3386_ _3514_/B _3387_/B _3514_/A _3387_/C vdd gnd OAI21X1
XFILL_3__1768_ gnd vdd FILL
XFILL_3__3507_ gnd vdd FILL
X_2337_ _2337_/A _2337_/B _2337_/C _3237_/D vdd gnd NAND3X1
XFILL_4__2300_ gnd vdd FILL
X_2268_ _2894_/A _2268_/B _2269_/B vdd gnd NOR2X1
XFILL_6__3216_ gnd vdd FILL
XFILL_4__2231_ gnd vdd FILL
XFILL_3__1699_ gnd vdd FILL
XFILL_1__2522_ gnd vdd FILL
XFILL_3__3438_ gnd vdd FILL
XFILL_1__2453_ gnd vdd FILL
XFILL_6__3147_ gnd vdd FILL
XFILL_4__2162_ gnd vdd FILL
XFILL_3__3369_ gnd vdd FILL
X_2199_ _2293_/A _2199_/B _2199_/C _2346_/A vdd gnd OAI21X1
XFILL_6__3078_ gnd vdd FILL
XFILL_1__2384_ gnd vdd FILL
XFILL_4__2093_ gnd vdd FILL
XFILL_7__2911_ gnd vdd FILL
XFILL_6__2029_ gnd vdd FILL
XFILL_7__2842_ gnd vdd FILL
XFILL_1__3005_ gnd vdd FILL
XFILL_7__2773_ gnd vdd FILL
XFILL_4__2995_ gnd vdd FILL
XFILL_7__1724_ gnd vdd FILL
XFILL_4__1946_ gnd vdd FILL
XFILL_4__1877_ gnd vdd FILL
XFILL_2__2700_ gnd vdd FILL
XFILL184650x70350 gnd vdd FILL
XFILL_4__3547_ gnd vdd FILL
XFILL_5__2340_ gnd vdd FILL
XFILL_2__2631_ gnd vdd FILL
XFILL_2__2562_ gnd vdd FILL
XFILL_4__3478_ gnd vdd FILL
XFILL_5__2271_ gnd vdd FILL
XFILL_7__2207_ gnd vdd FILL
XFILL_7__3187_ gnd vdd FILL
XFILL_2__2493_ gnd vdd FILL
XFILL_7__2138_ gnd vdd FILL
XFILL_4__2429_ gnd vdd FILL
XFILL_6_BUFX2_insert27 gnd vdd FILL
XFILL_6_BUFX2_insert16 gnd vdd FILL
XFILL_8__2951_ gnd vdd FILL
XFILL_6_BUFX2_insert49 gnd vdd FILL
XFILL_7__2069_ gnd vdd FILL
XFILL_2__3114_ gnd vdd FILL
XFILL_8__2882_ gnd vdd FILL
XFILL_8__1902_ gnd vdd FILL
XFILL_2__3045_ gnd vdd FILL
XFILL_8__1833_ gnd vdd FILL
XFILL_0__2060_ gnd vdd FILL
XFILL_8__1764_ gnd vdd FILL
XFILL_8__3503_ gnd vdd FILL
XFILL_5__1986_ gnd vdd FILL
XFILL_8__1695_ gnd vdd FILL
XFILL_8__3434_ gnd vdd FILL
XFILL_3__2740_ gnd vdd FILL
XFILL_0__2962_ gnd vdd FILL
XFILL_8__3365_ gnd vdd FILL
XFILL_5__2607_ gnd vdd FILL
XFILL_3__2671_ gnd vdd FILL
XFILL_2__2829_ gnd vdd FILL
XFILL_0__2893_ gnd vdd FILL
XFILL_5__3587_ gnd vdd FILL
XFILL_6__2380_ gnd vdd FILL
XFILL_8__2316_ gnd vdd FILL
X_3240_ _3240_/D vdd _3291_/R _3355_/CLK _3240_/Q vdd gnd DFFSR
XFILL_0__1913_ gnd vdd FILL
X_3171_ _3171_/A _3171_/B _3172_/A vdd gnd NOR2X1
XFILL_0__1844_ gnd vdd FILL
XFILL_8__2247_ gnd vdd FILL
XFILL_5__2538_ gnd vdd FILL
X_2122_ _2122_/A _2344_/B _2319_/A vdd gnd NAND2X1
XFILL_5__2469_ gnd vdd FILL
XFILL_0__1775_ gnd vdd FILL
XFILL_0__3514_ gnd vdd FILL
XFILL_6__3001_ gnd vdd FILL
XFILL_8__2178_ gnd vdd FILL
X_2053_ _3166_/C _3195_/B _2374_/C _2075_/A vdd gnd OAI21X1
XFILL_3__3223_ gnd vdd FILL
XFILL_0__3445_ gnd vdd FILL
XFILL_3__3154_ gnd vdd FILL
XFILL184350x148350 gnd vdd FILL
XFILL_0__3376_ gnd vdd FILL
XFILL_3__2105_ gnd vdd FILL
XFILL184050x156150 gnd vdd FILL
XFILL_0__2327_ gnd vdd FILL
XFILL_3__3085_ gnd vdd FILL
XFILL_3__2036_ gnd vdd FILL
X_2955_ reset _2957_/C _3306_/Q _2956_/C vdd gnd OAI21X1
XFILL_0__2258_ gnd vdd FILL
X_2886_ _2886_/A _2897_/C _2931_/B _2886_/D _3282_/D vdd gnd OAI22X1
X_1906_ _3174_/A _1910_/C vdd gnd INVX1
XFILL_0__2189_ gnd vdd FILL
XFILL_4__1800_ gnd vdd FILL
X_1837_ _1987_/A _3152_/C _3088_/S vdd gnd NAND2X1
XFILL_6__2716_ gnd vdd FILL
XFILL_4__2780_ gnd vdd FILL
X_3507_ _3555_/A _3554_/A vdd gnd INVX1
X_1768_ _3313_/Q _3007_/B _1769_/B vdd gnd NAND2X1
XFILL_3__2938_ gnd vdd FILL
XFILL_4__1731_ gnd vdd FILL
XFILL_6__2647_ gnd vdd FILL
XFILL_3__2869_ gnd vdd FILL
XFILL_1__1953_ gnd vdd FILL
X_1699_ _2768_/A DI[3] _1699_/C _2948_/A vdd gnd OAI21X1
XFILL_6__2578_ gnd vdd FILL
XFILL_4__3401_ gnd vdd FILL
X_3438_ _3438_/A _3449_/A vdd gnd INVX1
XFILL_1__1884_ gnd vdd FILL
XFILL_7__3110_ gnd vdd FILL
X_3369_ _3369_/A _3369_/B _3369_/Y vdd gnd NOR2X1
XFILL_7__3041_ gnd vdd FILL
XFILL_1__3554_ gnd vdd FILL
XFILL_1__3485_ gnd vdd FILL
XFILL_4__2214_ gnd vdd FILL
XFILL_1__2505_ gnd vdd FILL
XFILL_4__3194_ gnd vdd FILL
XFILL_4__2145_ gnd vdd FILL
XFILL_1__2436_ gnd vdd FILL
XFILL_1__2367_ gnd vdd FILL
XFILL184050x35250 gnd vdd FILL
XFILL_4__2076_ gnd vdd FILL
XFILL_1__2298_ gnd vdd FILL
XFILL_7__2825_ gnd vdd FILL
XFILL184650x82050 gnd vdd FILL
XFILL_7__2756_ gnd vdd FILL
XFILL_5__1840_ gnd vdd FILL
XFILL_4__2978_ gnd vdd FILL
XFILL_5__1771_ gnd vdd FILL
XFILL_7__1707_ gnd vdd FILL
XFILL_4__1929_ gnd vdd FILL
XFILL_5__3510_ gnd vdd FILL
XFILL_2__1993_ gnd vdd FILL
XFILL_7__2687_ gnd vdd FILL
XFILL_5__3441_ gnd vdd FILL
XFILL_8__3150_ gnd vdd FILL
XFILL_8__3081_ gnd vdd FILL
XFILL_5__3372_ gnd vdd FILL
XFILL_8__2101_ gnd vdd FILL
XFILL_2__2614_ gnd vdd FILL
XFILL_8__2032_ gnd vdd FILL
XFILL_5__2323_ gnd vdd FILL
XFILL_2__3594_ gnd vdd FILL
XFILL_5__2254_ gnd vdd FILL
XFILL_2__2545_ gnd vdd FILL
XFILL_2__2476_ gnd vdd FILL
XFILL_5__2185_ gnd vdd FILL
XFILL_8__2934_ gnd vdd FILL
XFILL_0__3230_ gnd vdd FILL
XFILL_0__3161_ gnd vdd FILL
XFILL_0__2112_ gnd vdd FILL
XFILL_8__2865_ gnd vdd FILL
XFILL_2__3028_ gnd vdd FILL
XFILL_6__1880_ gnd vdd FILL
XFILL_8__2796_ gnd vdd FILL
XFILL_0__3092_ gnd vdd FILL
XFILL_8__1816_ gnd vdd FILL
X_2740_ _2744_/B _2751_/B _2757_/A _2752_/A vdd gnd OAI21X1
XFILL_0__2043_ gnd vdd FILL
XFILL_8__1747_ gnd vdd FILL
X_2671_ _2676_/B _2671_/B _2686_/D _2674_/B vdd gnd OAI21X1
XFILL_6__3550_ gnd vdd FILL
XFILL_5__1969_ gnd vdd FILL
XFILL_6__2501_ gnd vdd FILL
XFILL_6__3481_ gnd vdd FILL
XFILL_8__3417_ gnd vdd FILL
XFILL_3__2723_ gnd vdd FILL
XFILL_2_BUFX2_insert25 gnd vdd FILL
XFILL_2_BUFX2_insert14 gnd vdd FILL
XFILL_2_BUFX2_insert58 gnd vdd FILL
XFILL_0__2945_ gnd vdd FILL
XFILL_2_BUFX2_insert47 gnd vdd FILL
XFILL_6__2432_ gnd vdd FILL
XFILL_2_BUFX2_insert69 gnd vdd FILL
XFILL_6__2363_ gnd vdd FILL
X_3223_ _3582_/A _3227_/B _3224_/C vdd gnd NAND2X1
XFILL_3__2654_ gnd vdd FILL
XFILL_0__2876_ gnd vdd FILL
XFILL_3__2585_ gnd vdd FILL
XFILL_0__1827_ gnd vdd FILL
X_3154_ _3154_/A _3154_/B _3196_/A vdd gnd NOR2X1
XFILL_6__2294_ gnd vdd FILL
X_3085_ _3568_/Q _3085_/B _3086_/A vdd gnd NOR2X1
XFILL_0__1758_ gnd vdd FILL
X_2105_ _2294_/A _2438_/A _2106_/C vdd gnd NAND2X1
X_2036_ _2890_/A _2864_/A _2922_/A vdd gnd NAND2X1
XFILL_0__1689_ gnd vdd FILL
XFILL_3__3206_ gnd vdd FILL
XFILL_0__3428_ gnd vdd FILL
XFILL_1__2221_ gnd vdd FILL
XFILL_3__3137_ gnd vdd FILL
XFILL_3__3068_ gnd vdd FILL
XFILL_1__2152_ gnd vdd FILL
XFILL_1__2083_ gnd vdd FILL
XFILL_4__2901_ gnd vdd FILL
XFILL_3__2019_ gnd vdd FILL
X_2938_ _2938_/A _3157_/C _3022_/A _2957_/C vdd gnd OAI21X1
XFILL_7__3590_ gnd vdd FILL
XFILL_7__2610_ gnd vdd FILL
XFILL_4__2832_ gnd vdd FILL
X_2869_ _3007_/C _2957_/B _2869_/C _3276_/D vdd gnd OAI21X1
XFILL_7__2541_ gnd vdd FILL
XFILL_4__2763_ gnd vdd FILL
XFILL_8_CLKBUF1_insert34 gnd vdd FILL
XFILL_1__2985_ gnd vdd FILL
XFILL_7__2472_ gnd vdd FILL
XFILL_4__1714_ gnd vdd FILL
XFILL_1__1936_ gnd vdd FILL
XFILL_4__2694_ gnd vdd FILL
XFILL_1__1867_ gnd vdd FILL
XFILL_1_BUFX2_insert0 gnd vdd FILL
XFILL_1__1798_ gnd vdd FILL
XFILL_1__3537_ gnd vdd FILL
XFILL_2__2330_ gnd vdd FILL
XFILL_7__3024_ gnd vdd FILL
XFILL_2__2261_ gnd vdd FILL
XFILL_1__3468_ gnd vdd FILL
XFILL_4__3177_ gnd vdd FILL
XFILL_1__3399_ gnd vdd FILL
XFILL_1__2419_ gnd vdd FILL
XFILL_4__2128_ gnd vdd FILL
XFILL_2__2192_ gnd vdd FILL
XFILL_5__2941_ gnd vdd FILL
XFILL_4__2059_ gnd vdd FILL
XFILL_8__2650_ gnd vdd FILL
XFILL_7__2808_ gnd vdd FILL
XFILL_5__2872_ gnd vdd FILL
XFILL_5__1823_ gnd vdd FILL
XFILL_8__2581_ gnd vdd FILL
XFILL_7__2739_ gnd vdd FILL
XFILL_5__1754_ gnd vdd FILL
XFILL_2__1976_ gnd vdd FILL
XFILL_9_BUFX2_insert53 gnd vdd FILL
XFILL_8__3202_ gnd vdd FILL
XFILL_8__3133_ gnd vdd FILL
XFILL_5__3424_ gnd vdd FILL
XFILL_0__2730_ gnd vdd FILL
XFILL_9_BUFX2_insert97 gnd vdd FILL
XFILL_3__2370_ gnd vdd FILL
XFILL_5__2306_ gnd vdd FILL
XFILL_8__3064_ gnd vdd FILL
XFILL_0__2661_ gnd vdd FILL
XFILL_8__2015_ gnd vdd FILL
XFILL_2__2528_ gnd vdd FILL
XFILL_0__2592_ gnd vdd FILL
XFILL_5__2237_ gnd vdd FILL
XFILL_5__2168_ gnd vdd FILL
XFILL_2__2459_ gnd vdd FILL
XFILL_8__2917_ gnd vdd FILL
XFILL_6__2981_ gnd vdd FILL
XFILL_0__3213_ gnd vdd FILL
XFILL_4_BUFX2_insert4 gnd vdd FILL
XFILL_5__2099_ gnd vdd FILL
XFILL_8__2848_ gnd vdd FILL
XFILL_6__1932_ gnd vdd FILL
XFILL_0__3144_ gnd vdd FILL
XFILL_0__3075_ gnd vdd FILL
XFILL_6__1863_ gnd vdd FILL
X_2723_ _2778_/A _2723_/B _2723_/C _3249_/D vdd gnd OAI21X1
XFILL_0__2026_ gnd vdd FILL
XFILL_6__3602_ gnd vdd FILL
XFILL_8__2779_ gnd vdd FILL
XFILL_6__1794_ gnd vdd FILL
X_2654_ _3243_/Q _2685_/B _2656_/A vdd gnd NAND2X1
XFILL_6__3533_ gnd vdd FILL
X_2585_ _3147_/C _2702_/B _3167_/B _2587_/A vdd gnd OAI21X1
XFILL_6__3464_ gnd vdd FILL
XFILL_6__2415_ gnd vdd FILL
XFILL_3__2706_ gnd vdd FILL
XFILL_1__2770_ gnd vdd FILL
XFILL_0__2928_ gnd vdd FILL
XFILL_6__3395_ gnd vdd FILL
XFILL_1__1721_ gnd vdd FILL
XFILL_3__2637_ gnd vdd FILL
XFILL_0__2859_ gnd vdd FILL
XFILL_6__2346_ gnd vdd FILL
X_3206_ _3214_/A _3214_/B _3351_/Q _3207_/C vdd gnd OAI21X1
XFILL_4__3100_ gnd vdd FILL
X_3137_ _3137_/A _3143_/B _3137_/C _3344_/D vdd gnd OAI21X1
XFILL_6__2277_ gnd vdd FILL
XFILL_3__2568_ gnd vdd FILL
XFILL_3__2499_ gnd vdd FILL
XFILL_4__3031_ gnd vdd FILL
X_3068_ _3568_/Q _3085_/B _3084_/B _3069_/A vdd gnd OAI21X1
X_2019_ _2161_/B _2889_/A _2889_/C _2845_/A vdd gnd OAI21X1
XFILL_1__2204_ gnd vdd FILL
XFILL_7__1972_ gnd vdd FILL
XFILL_1__3184_ gnd vdd FILL
XFILL_1__2135_ gnd vdd FILL
XFILL_1__2066_ gnd vdd FILL
XFILL_4__2815_ gnd vdd FILL
XFILL_7_BUFX2_insert8 gnd vdd FILL
XFILL_7__2524_ gnd vdd FILL
XFILL_2__1830_ gnd vdd FILL
XFILL_7__2455_ gnd vdd FILL
XFILL_4__2746_ gnd vdd FILL
XFILL_1__2968_ gnd vdd FILL
XFILL_2__1761_ gnd vdd FILL
XFILL_4__2677_ gnd vdd FILL
XFILL_1__2899_ gnd vdd FILL
XFILL_2__3500_ gnd vdd FILL
XFILL_1__1919_ gnd vdd FILL
XFILL_7__2386_ gnd vdd FILL
XFILL_2__1692_ gnd vdd FILL
XFILL_2__3431_ gnd vdd FILL
XFILL_5__3140_ gnd vdd FILL
XFILL_7__3007_ gnd vdd FILL
XFILL_5__3071_ gnd vdd FILL
XFILL_5__2022_ gnd vdd FILL
XFILL_2__2313_ gnd vdd FILL
XFILL_4__3229_ gnd vdd FILL
XFILL_2__2244_ gnd vdd FILL
XFILL_2__2175_ gnd vdd FILL
XFILL_8__2702_ gnd vdd FILL
XFILL_5__2924_ gnd vdd FILL
XFILL_8__2633_ gnd vdd FILL
XFILL_5__2855_ gnd vdd FILL
XFILL_8__2564_ gnd vdd FILL
XFILL_3__1870_ gnd vdd FILL
XFILL_5__2786_ gnd vdd FILL
XFILL_5__1806_ gnd vdd FILL
XFILL_8__2495_ gnd vdd FILL
XFILL_5__1737_ gnd vdd FILL
XFILL_2__1959_ gnd vdd FILL
X_2370_ _2861_/A _2579_/B _2370_/C _3514_/B vdd gnd OAI21X1
XFILL_3__3540_ gnd vdd FILL
XFILL_3__3471_ gnd vdd FILL
XFILL_5__3407_ gnd vdd FILL
XFILL_6__2200_ gnd vdd FILL
XFILL_8__3116_ gnd vdd FILL
XFILL_3__2422_ gnd vdd FILL
XFILL_0__2713_ gnd vdd FILL
XFILL_6__3180_ gnd vdd FILL
XFILL_8__3047_ gnd vdd FILL
XFILL_6__2131_ gnd vdd FILL
XFILL_0__2644_ gnd vdd FILL
XFILL_3__2353_ gnd vdd FILL
XFILL_6__2062_ gnd vdd FILL
XFILL_0__2575_ gnd vdd FILL
XFILL_3__2284_ gnd vdd FILL
XFILL_9__2811_ gnd vdd FILL
XFILL_5_BUFX2_insert51 gnd vdd FILL
XFILL_5_BUFX2_insert62 gnd vdd FILL
XFILL_6__2964_ gnd vdd FILL
XFILL_5_BUFX2_insert40 gnd vdd FILL
XFILL_5_BUFX2_insert95 gnd vdd FILL
XFILL_5_BUFX2_insert84 gnd vdd FILL
XFILL_5_BUFX2_insert73 gnd vdd FILL
XFILL_6__1915_ gnd vdd FILL
XFILL_0__3127_ gnd vdd FILL
XFILL_6__2895_ gnd vdd FILL
XFILL_0__3058_ gnd vdd FILL
X_2706_ _2706_/A _2706_/B _2706_/C _2711_/D vdd gnd AOI21X1
XFILL_6__1846_ gnd vdd FILL
XFILL_6__1777_ gnd vdd FILL
X_2637_ _3242_/Q _2685_/B _2638_/C vdd gnd NAND2X1
XFILL_0__2009_ gnd vdd FILL
XFILL_6__3516_ gnd vdd FILL
XFILL_3__1999_ gnd vdd FILL
XFILL_4__3580_ gnd vdd FILL
XFILL_4__2600_ gnd vdd FILL
XFILL_1__2822_ gnd vdd FILL
XFILL_4__2531_ gnd vdd FILL
X_2568_ _3577_/Q _2570_/A vdd gnd INVX1
XFILL_6__3447_ gnd vdd FILL
X_2499_ _2499_/A _2519_/C _2499_/C _3211_/B vdd gnd AOI21X1
XFILL_7__2240_ gnd vdd FILL
XFILL_1__2753_ gnd vdd FILL
XFILL_6__3378_ gnd vdd FILL
XFILL_7__2171_ gnd vdd FILL
XFILL_1__1704_ gnd vdd FILL
XFILL_4__2462_ gnd vdd FILL
XFILL_4__2393_ gnd vdd FILL
XFILL_6__2329_ gnd vdd FILL
XFILL_1__2684_ gnd vdd FILL
XFILL_4__3014_ gnd vdd FILL
XFILL_7__1955_ gnd vdd FILL
XFILL_1__3167_ gnd vdd FILL
XFILL_1__3098_ gnd vdd FILL
XFILL_1__2118_ gnd vdd FILL
XFILL_7__1886_ gnd vdd FILL
XFILL_2__2931_ gnd vdd FILL
XFILL_1__2049_ gnd vdd FILL
XFILL_7__3556_ gnd vdd FILL
XFILL_5__2640_ gnd vdd FILL
XFILL_2__2862_ gnd vdd FILL
XFILL_7__2507_ gnd vdd FILL
XFILL_5__2571_ gnd vdd FILL
XFILL_7__3487_ gnd vdd FILL
XFILL_2__2793_ gnd vdd FILL
XFILL_8__2280_ gnd vdd FILL
XFILL_4__2729_ gnd vdd FILL
XFILL_2__1813_ gnd vdd FILL
XFILL_2__1744_ gnd vdd FILL
XFILL_7__2438_ gnd vdd FILL
XFILL_7__2369_ gnd vdd FILL
XFILL_5__3123_ gnd vdd FILL
XFILL_2__3414_ gnd vdd FILL
XFILL_0__2360_ gnd vdd FILL
XFILL_5__3054_ gnd vdd FILL
XFILL_5__2005_ gnd vdd FILL
XFILL_0__2291_ gnd vdd FILL
XFILL_2__2227_ gnd vdd FILL
XFILL_8__1995_ gnd vdd FILL
X_1870_ _3286_/Q _2913_/A vdd gnd INVX1
XFILL_2__2158_ gnd vdd FILL
XFILL_2__2089_ gnd vdd FILL
XFILL_5__2907_ gnd vdd FILL
X_3540_ _3569_/Q _3553_/B _3541_/C vdd gnd NAND2X1
XFILL_6__1700_ gnd vdd FILL
XFILL_3__2971_ gnd vdd FILL
XFILL184650x7950 gnd vdd FILL
XFILL_6__2680_ gnd vdd FILL
XFILL_8__2616_ gnd vdd FILL
XFILL_5__2838_ gnd vdd FILL
XFILL_8__3596_ gnd vdd FILL
XFILL_3__1922_ gnd vdd FILL
X_3471_ _3471_/A _3471_/B _3521_/A _3472_/A vdd gnd AOI21X1
XFILL_3__1853_ gnd vdd FILL
XFILL_8__2547_ gnd vdd FILL
X_2422_ _2422_/A _2422_/B _2422_/C _3601_/A vdd gnd NAND3X1
XFILL_8__2478_ gnd vdd FILL
XFILL_5__2769_ gnd vdd FILL
XFILL_3__3523_ gnd vdd FILL
X_2353_ _2353_/A _2353_/B _3238_/D vdd gnd OR2X2
XFILL_3__1784_ gnd vdd FILL
XFILL_6__3232_ gnd vdd FILL
XFILL_3__3454_ gnd vdd FILL
X_2284_ _2284_/A _2332_/B _2285_/A vdd gnd AND2X2
XFILL_6__3163_ gnd vdd FILL
XFILL_3__3385_ gnd vdd FILL
XFILL_6__2114_ gnd vdd FILL
XFILL_3__2405_ gnd vdd FILL
XFILL_6__3094_ gnd vdd FILL
XFILL_3__2336_ gnd vdd FILL
XFILL_0__2627_ gnd vdd FILL
XBUFX2_insert1 _1773_/Y _2058_/B vdd gnd BUFX2
XFILL_6__2045_ gnd vdd FILL
XFILL_0__2558_ gnd vdd FILL
XFILL_3__2267_ gnd vdd FILL
XFILL_0__2489_ gnd vdd FILL
XFILL_3__2198_ gnd vdd FILL
XFILL_1__3021_ gnd vdd FILL
XFILL_6__2947_ gnd vdd FILL
XFILL_7__1740_ gnd vdd FILL
X_1999_ _2006_/A _3291_/D _1999_/C _2249_/A vdd gnd OAI21X1
XFILL_6__2878_ gnd vdd FILL
XFILL_4__1962_ gnd vdd FILL
XFILL_7__3410_ gnd vdd FILL
XFILL_6__1829_ gnd vdd FILL
XFILL_4__1893_ gnd vdd FILL
XFILL_1__2805_ gnd vdd FILL
XFILL_4__3563_ gnd vdd FILL
XFILL_4__3494_ gnd vdd FILL
XFILL_7__2223_ gnd vdd FILL
XFILL_4__2514_ gnd vdd FILL
XFILL_3_CLKBUF1_insert35 gnd vdd FILL
XFILL_1_BUFX2_insert60 gnd vdd FILL
XFILL_1__2736_ gnd vdd FILL
XFILL_4__2445_ gnd vdd FILL
XFILL_1_BUFX2_insert93 gnd vdd FILL
XFILL_1_BUFX2_insert82 gnd vdd FILL
XFILL_7__2154_ gnd vdd FILL
XFILL_1__2667_ gnd vdd FILL
XFILL_1_BUFX2_insert71 gnd vdd FILL
XFILL_7__2085_ gnd vdd FILL
XFILL_4__2376_ gnd vdd FILL
XFILL_2__3130_ gnd vdd FILL
XFILL_1__2598_ gnd vdd FILL
XFILL_2__3061_ gnd vdd FILL
XFILL_2__2012_ gnd vdd FILL
XFILL_7__2987_ gnd vdd FILL
XFILL_8__1780_ gnd vdd FILL
XFILL_1__3219_ gnd vdd FILL
XFILL_7__1938_ gnd vdd FILL
XFILL_8__3450_ gnd vdd FILL
XFILL_7__1869_ gnd vdd FILL
XFILL_8__2401_ gnd vdd FILL
XFILL_2__2914_ gnd vdd FILL
XFILL_8__3381_ gnd vdd FILL
XFILL_5__2623_ gnd vdd FILL
XFILL_2__2845_ gnd vdd FILL
XFILL_7__3539_ gnd vdd FILL
XFILL_8__2332_ gnd vdd FILL
XFILL_0__1860_ gnd vdd FILL
XFILL_8__2263_ gnd vdd FILL
XFILL_5__2554_ gnd vdd FILL
XFILL_5__2485_ gnd vdd FILL
XFILL_2__2776_ gnd vdd FILL
XFILL_8__2194_ gnd vdd FILL
XFILL_0__1791_ gnd vdd FILL
XFILL_2__1727_ gnd vdd FILL
XFILL_0__3530_ gnd vdd FILL
XFILL_0__3461_ gnd vdd FILL
XFILL_5__3106_ gnd vdd FILL
XFILL_0__2412_ gnd vdd FILL
XFILL_3__3170_ gnd vdd FILL
XFILL_0__3392_ gnd vdd FILL
XFILL_5__3037_ gnd vdd FILL
XFILL_3__2121_ gnd vdd FILL
X_2971_ _2971_/A _2971_/B _2971_/C _3308_/D vdd gnd OAI21X1
XFILL_0__2343_ gnd vdd FILL
XFILL_3__2052_ gnd vdd FILL
XFILL_8__1978_ gnd vdd FILL
XFILL_0__2274_ gnd vdd FILL
X_1922_ _3357_/Q _3219_/A vdd gnd INVX1
XFILL_6__2801_ gnd vdd FILL
X_1853_ _3151_/C _3182_/B _3178_/B _1863_/B vdd gnd OAI21X1
XFILL_6__2732_ gnd vdd FILL
XFILL_3__2954_ gnd vdd FILL
X_1784_ _3190_/B _3156_/B vdd gnd INVX2
X_3523_ _3523_/A _3523_/B _3562_/B vdd gnd XOR2X1
XFILL_8__3579_ gnd vdd FILL
XFILL_3__1905_ gnd vdd FILL
XFILL_6__2663_ gnd vdd FILL
X_3454_ _3468_/A _3521_/B _3469_/B vdd gnd NAND2X1
XFILL_3__2885_ gnd vdd FILL
XFILL_6__2594_ gnd vdd FILL
X_2405_ _2423_/A _2416_/A vdd gnd INVX1
XFILL_3__1836_ gnd vdd FILL
X_3385_ _3442_/B _3514_/A vdd gnd INVX4
XFILL_3__1767_ gnd vdd FILL
XFILL_3__3506_ gnd vdd FILL
X_2336_ _2336_/A _2336_/B _2337_/B vdd gnd NOR2X1
XFILL_0__1989_ gnd vdd FILL
XFILL_6__3215_ gnd vdd FILL
X_2267_ _2843_/C _2911_/A _2269_/A vdd gnd NAND2X1
XFILL_3__3437_ gnd vdd FILL
XFILL_1__2521_ gnd vdd FILL
XFILL_4__2230_ gnd vdd FILL
XFILL_3__1698_ gnd vdd FILL
XFILL_1__2452_ gnd vdd FILL
XFILL_6__3146_ gnd vdd FILL
XFILL_4__2161_ gnd vdd FILL
XFILL_6__3077_ gnd vdd FILL
XFILL_3__3368_ gnd vdd FILL
X_2198_ _2293_/A _3160_/A _3151_/A _2199_/C vdd gnd NAND3X1
XFILL_6__2028_ gnd vdd FILL
XFILL_1__2383_ gnd vdd FILL
XFILL_3__2319_ gnd vdd FILL
XFILL_4__2092_ gnd vdd FILL
XFILL_7__2910_ gnd vdd FILL
XFILL_7__2841_ gnd vdd FILL
XFILL_1__3004_ gnd vdd FILL
XFILL_7__2772_ gnd vdd FILL
XFILL_4__2994_ gnd vdd FILL
XFILL_9__2708_ gnd vdd FILL
XFILL_7__1723_ gnd vdd FILL
XFILL_4__1945_ gnd vdd FILL
XFILL_4__1876_ gnd vdd FILL
XFILL_4__3546_ gnd vdd FILL
XFILL_2__2630_ gnd vdd FILL
XFILL_2__2561_ gnd vdd FILL
XFILL_4__3477_ gnd vdd FILL
XFILL_5__2270_ gnd vdd FILL
XFILL_7__2206_ gnd vdd FILL
XFILL184650x89850 gnd vdd FILL
XFILL_1__2719_ gnd vdd FILL
XFILL_7__3186_ gnd vdd FILL
XFILL_4__2428_ gnd vdd FILL
XFILL_2__2492_ gnd vdd FILL
XFILL_7__2137_ gnd vdd FILL
XFILL_4__2359_ gnd vdd FILL
XFILL_6_BUFX2_insert17 gnd vdd FILL
XFILL_8__2950_ gnd vdd FILL
XFILL_7__2068_ gnd vdd FILL
XFILL_6_BUFX2_insert39 gnd vdd FILL
XFILL_2__3113_ gnd vdd FILL
XFILL_8__2881_ gnd vdd FILL
XFILL_8__1901_ gnd vdd FILL
XFILL_2__3044_ gnd vdd FILL
XFILL_8__1832_ gnd vdd FILL
XFILL_8__1763_ gnd vdd FILL
XFILL_8__3502_ gnd vdd FILL
XFILL_5__1985_ gnd vdd FILL
XFILL_8__1694_ gnd vdd FILL
XFILL_8__3433_ gnd vdd FILL
XFILL181650x140550 gnd vdd FILL
XFILL_0__2961_ gnd vdd FILL
XFILL_8__3364_ gnd vdd FILL
XFILL_8__2315_ gnd vdd FILL
XFILL_5__3586_ gnd vdd FILL
XFILL_0__1912_ gnd vdd FILL
XFILL_5__2606_ gnd vdd FILL
XFILL_3__2670_ gnd vdd FILL
XFILL_2__2828_ gnd vdd FILL
XFILL_0__2892_ gnd vdd FILL
XFILL_5__2537_ gnd vdd FILL
XFILL_0__1843_ gnd vdd FILL
XFILL_8__2246_ gnd vdd FILL
X_3170_ _3170_/A _3170_/B _3214_/A vdd gnd NOR2X1
XFILL_2__2759_ gnd vdd FILL
XFILL_8__2177_ gnd vdd FILL
XFILL_5__2468_ gnd vdd FILL
X_2121_ _2342_/A _2289_/B _2121_/C _2122_/A vdd gnd OAI21X1
XFILL_0__1774_ gnd vdd FILL
XFILL_0__3513_ gnd vdd FILL
XFILL_6__3000_ gnd vdd FILL
XFILL_5__2399_ gnd vdd FILL
X_2052_ _3171_/A _2052_/B _2374_/C vdd gnd NOR2X1
XFILL_3__3222_ gnd vdd FILL
XFILL_0__3444_ gnd vdd FILL
XFILL_3__3153_ gnd vdd FILL
XFILL_3__2104_ gnd vdd FILL
XFILL_0__3375_ gnd vdd FILL
XFILL_3__3084_ gnd vdd FILL
XFILL_0__2326_ gnd vdd FILL
XCLKBUF1_insert30 clk _3363_/CLK vdd gnd CLKBUF1
XFILL_3__2035_ gnd vdd FILL
X_2954_ _3079_/A _2956_/B _2954_/C _3305_/D vdd gnd OAI21X1
X_2885_ _2895_/A _2885_/B _2886_/D vdd gnd OR2X2
XFILL_0__2257_ gnd vdd FILL
X_1905_ _2433_/B _3158_/A vdd gnd INVX1
XFILL_0__2188_ gnd vdd FILL
X_1836_ _3025_/A _1843_/A vdd gnd INVX1
X_1767_ _3276_/Q _3007_/C vdd gnd INVX1
XFILL_6__2715_ gnd vdd FILL
X_3506_ _3508_/A _3506_/B _3529_/C _3555_/A vdd gnd OAI21X1
XFILL_4__1730_ gnd vdd FILL
XFILL_3__2937_ gnd vdd FILL
XFILL_6__2646_ gnd vdd FILL
XFILL_3__2868_ gnd vdd FILL
XFILL_9__2355_ gnd vdd FILL
XFILL_1__1952_ gnd vdd FILL
X_1698_ _3197_/C _3293_/Q _1699_/C vdd gnd OR2X2
XFILL_4__3400_ gnd vdd FILL
X_3437_ _3442_/A _3439_/B vdd gnd INVX1
XFILL_6__2577_ gnd vdd FILL
XFILL_3__1819_ gnd vdd FILL
XFILL_1__1883_ gnd vdd FILL
XFILL_3__2799_ gnd vdd FILL
X_3368_ _3368_/A _3368_/B _3368_/C _3369_/B vdd gnd NAND3X1
XFILL_1__3553_ gnd vdd FILL
XFILL_7__3040_ gnd vdd FILL
X_2319_ _2319_/A _2319_/B _2321_/B vdd gnd OR2X2
X_3299_ _3299_/D _3577_/CLK _3299_/Q vdd gnd DFFPOSX1
XFILL_1__2504_ gnd vdd FILL
XFILL_1__3484_ gnd vdd FILL
XFILL_6__3129_ gnd vdd FILL
XFILL_4__2213_ gnd vdd FILL
XFILL_4__3193_ gnd vdd FILL
XFILL_4__2144_ gnd vdd FILL
XFILL184350x19650 gnd vdd FILL
XFILL_1__2435_ gnd vdd FILL
XFILL_1__2366_ gnd vdd FILL
XFILL_4__2075_ gnd vdd FILL
XFILL_1__2297_ gnd vdd FILL
XFILL_7__2824_ gnd vdd FILL
XFILL181950x74250 gnd vdd FILL
XFILL_7__2755_ gnd vdd FILL
XFILL_4__2977_ gnd vdd FILL
XFILL_5__1770_ gnd vdd FILL
XFILL_7__1706_ gnd vdd FILL
XFILL_7__2686_ gnd vdd FILL
XFILL_4__1928_ gnd vdd FILL
XFILL_2__1992_ gnd vdd FILL
XFILL_4__1859_ gnd vdd FILL
XFILL_5__3440_ gnd vdd FILL
XFILL_8__3080_ gnd vdd FILL
XFILL_5__3371_ gnd vdd FILL
XFILL_2__2613_ gnd vdd FILL
XFILL_8__2100_ gnd vdd FILL
XFILL_4__3529_ gnd vdd FILL
XFILL_5__2322_ gnd vdd FILL
XFILL_8__2031_ gnd vdd FILL
XFILL_2__3593_ gnd vdd FILL
XFILL_5__2253_ gnd vdd FILL
XFILL_2__2544_ gnd vdd FILL
XFILL_2__2475_ gnd vdd FILL
XFILL_7__3169_ gnd vdd FILL
XFILL_5__2184_ gnd vdd FILL
XFILL_8__2933_ gnd vdd FILL
XFILL_0__3160_ gnd vdd FILL
XFILL_8__2864_ gnd vdd FILL
XFILL_0__2111_ gnd vdd FILL
XFILL_0__3091_ gnd vdd FILL
XFILL_2__3027_ gnd vdd FILL
XFILL_8__2795_ gnd vdd FILL
XFILL_8__1815_ gnd vdd FILL
XFILL_0__2042_ gnd vdd FILL
XFILL_8__1746_ gnd vdd FILL
X_2670_ _3577_/Q _2670_/B _2670_/C _2686_/D vdd gnd AOI21X1
XFILL_5__1968_ gnd vdd FILL
XFILL_6__3480_ gnd vdd FILL
XFILL_6__2500_ gnd vdd FILL
XFILL_2_BUFX2_insert26 gnd vdd FILL
XFILL_8__3416_ gnd vdd FILL
XFILL_5__1899_ gnd vdd FILL
XFILL_3__2722_ gnd vdd FILL
XFILL_2_BUFX2_insert15 gnd vdd FILL
XFILL_6__2431_ gnd vdd FILL
XFILL_2_BUFX2_insert59 gnd vdd FILL
XFILL_2_BUFX2_insert48 gnd vdd FILL
XFILL_0__2944_ gnd vdd FILL
XFILL_3__2653_ gnd vdd FILL
XFILL_6__2362_ gnd vdd FILL
XFILL_0__2875_ gnd vdd FILL
X_3222_ _3359_/Q _3224_/A vdd gnd INVX1
XFILL_3__2584_ gnd vdd FILL
X_3153_ _3187_/A _3153_/B _3192_/B _3154_/A vdd gnd NAND3X1
XFILL_8__2229_ gnd vdd FILL
XFILL_6__2293_ gnd vdd FILL
XFILL_0__1826_ gnd vdd FILL
X_2104_ _2104_/A _2438_/A vdd gnd INVX1
X_3084_ _3084_/A _3084_/B _3084_/C _3087_/A vdd gnd OAI21X1
XFILL_0__1757_ gnd vdd FILL
X_2035_ _2957_/A _2948_/A _2035_/C _2864_/A vdd gnd AOI21X1
XFILL_3__3205_ gnd vdd FILL
XFILL_0__1688_ gnd vdd FILL
XFILL_0__3427_ gnd vdd FILL
XFILL_9__2973_ gnd vdd FILL
XFILL_1__2220_ gnd vdd FILL
XFILL_3__3136_ gnd vdd FILL
XFILL_3__3067_ gnd vdd FILL
XFILL_1__2151_ gnd vdd FILL
XFILL_4__2900_ gnd vdd FILL
XFILL_3__2018_ gnd vdd FILL
XFILL_0__2309_ gnd vdd FILL
XFILL_1__2082_ gnd vdd FILL
X_2937_ _3147_/C _3298_/Q _3298_/D vdd gnd AND2X2
X_2868_ _2868_/A _2868_/B _2957_/B _2869_/C vdd gnd OAI21X1
XFILL_4__2831_ gnd vdd FILL
XFILL_7__2540_ gnd vdd FILL
X_2799_ _2813_/C _2803_/D _2799_/C _3262_/D vdd gnd OAI21X1
X_1819_ _2621_/B _3189_/C _3043_/A _1831_/D _3451_/B vdd gnd OAI22X1
XFILL_4__2762_ gnd vdd FILL
XFILL_8_CLKBUF1_insert35 gnd vdd FILL
XFILL_1__2984_ gnd vdd FILL
XFILL_7__2471_ gnd vdd FILL
XFILL_4__1713_ gnd vdd FILL
XFILL_1__1935_ gnd vdd FILL
XFILL_4__2693_ gnd vdd FILL
XFILL_6__2629_ gnd vdd FILL
XFILL_1__1866_ gnd vdd FILL
XFILL_7__3023_ gnd vdd FILL
XFILL_1_BUFX2_insert1 gnd vdd FILL
XFILL_1__1797_ gnd vdd FILL
XFILL_1__3536_ gnd vdd FILL
XFILL_1__3467_ gnd vdd FILL
XFILL_2__2260_ gnd vdd FILL
XFILL_1__2418_ gnd vdd FILL
XFILL_4__3176_ gnd vdd FILL
XFILL_1__3398_ gnd vdd FILL
XFILL_2__2191_ gnd vdd FILL
XFILL_4__2127_ gnd vdd FILL
XFILL_5__2940_ gnd vdd FILL
XFILL_1__2349_ gnd vdd FILL
XFILL_4__2058_ gnd vdd FILL
XFILL_8__2580_ gnd vdd FILL
XFILL_7__2807_ gnd vdd FILL
XFILL_5__2871_ gnd vdd FILL
XFILL_5__1822_ gnd vdd FILL
XFILL_5__1753_ gnd vdd FILL
XFILL_7__2738_ gnd vdd FILL
XFILL_2__1975_ gnd vdd FILL
XFILL_7__2669_ gnd vdd FILL
XFILL_8__3201_ gnd vdd FILL
XFILL_8__3132_ gnd vdd FILL
XFILL_5__3423_ gnd vdd FILL
XFILL_5__2305_ gnd vdd FILL
XFILL_0__2660_ gnd vdd FILL
XFILL_8__3063_ gnd vdd FILL
XFILL_8__2014_ gnd vdd FILL
XFILL_2__2527_ gnd vdd FILL
XFILL_0__2591_ gnd vdd FILL
XFILL_5__2236_ gnd vdd FILL
XFILL_5__2167_ gnd vdd FILL
XFILL_2__2458_ gnd vdd FILL
XFILL_2__2389_ gnd vdd FILL
XFILL_0__3212_ gnd vdd FILL
XFILL_8__2916_ gnd vdd FILL
XFILL_6__2980_ gnd vdd FILL
XFILL_4_BUFX2_insert5 gnd vdd FILL
XFILL_5__2098_ gnd vdd FILL
XFILL_0__3143_ gnd vdd FILL
XFILL_8__2847_ gnd vdd FILL
XFILL183150x140550 gnd vdd FILL
XFILL_6__1931_ gnd vdd FILL
XFILL_6__1862_ gnd vdd FILL
XFILL_0__3074_ gnd vdd FILL
X_2722_ _2722_/A _2732_/A _2723_/B vdd gnd XOR2X1
XFILL_0__2025_ gnd vdd FILL
XFILL_6__3601_ gnd vdd FILL
XFILL_8__2778_ gnd vdd FILL
XFILL_6__3532_ gnd vdd FILL
XFILL_8__1729_ gnd vdd FILL
XFILL_6__1793_ gnd vdd FILL
X_2653_ _2653_/A _2653_/B _2653_/C _2659_/D vdd gnd AOI21X1
X_2584_ _2589_/A _3166_/B _2589_/D _3167_/B vdd gnd OAI21X1
XFILL_6__3463_ gnd vdd FILL
XFILL_3__2705_ gnd vdd FILL
XFILL_0__2927_ gnd vdd FILL
XFILL_6__3394_ gnd vdd FILL
XFILL_6__2414_ gnd vdd FILL
XFILL_1__1720_ gnd vdd FILL
XFILL_6__2345_ gnd vdd FILL
XFILL_3__2636_ gnd vdd FILL
XFILL_0__2858_ gnd vdd FILL
X_3205_ _3215_/A _3205_/B _3205_/C _3350_/D vdd gnd OAI21X1
XFILL_3__2567_ gnd vdd FILL
X_3136_ _3344_/Q _3143_/B _3137_/C vdd gnd NAND2X1
XFILL_0__2789_ gnd vdd FILL
XFILL_6__2276_ gnd vdd FILL
XFILL_0__1809_ gnd vdd FILL
X_3067_ _3339_/Q _3278_/Q _3568_/Q _3084_/B vdd gnd NAND3X1
XFILL_3__2498_ gnd vdd FILL
X_2018_ _2033_/A _2952_/A _2018_/C _2889_/A vdd gnd OAI21X1
XFILL_4__3030_ gnd vdd FILL
XFILL_3__3119_ gnd vdd FILL
XFILL_1__2203_ gnd vdd FILL
XFILL_1__3183_ gnd vdd FILL
XFILL_7__1971_ gnd vdd FILL
XFILL_1__2134_ gnd vdd FILL
XFILL_1__2065_ gnd vdd FILL
XFILL_4__2814_ gnd vdd FILL
XFILL_7_BUFX2_insert9 gnd vdd FILL
XFILL_7__2523_ gnd vdd FILL
XFILL_7__2454_ gnd vdd FILL
XFILL_4__2745_ gnd vdd FILL
XFILL_2__1760_ gnd vdd FILL
XFILL_1__2967_ gnd vdd FILL
XFILL_4__2676_ gnd vdd FILL
XFILL_1__1918_ gnd vdd FILL
XFILL_1__2898_ gnd vdd FILL
XFILL_7__2385_ gnd vdd FILL
XFILL_2__1691_ gnd vdd FILL
XFILL_2__3430_ gnd vdd FILL
XFILL_1__1849_ gnd vdd FILL
XFILL_1__3519_ gnd vdd FILL
XFILL_7__3006_ gnd vdd FILL
XFILL_2__2312_ gnd vdd FILL
XFILL_5__3070_ gnd vdd FILL
XFILL_5__2021_ gnd vdd FILL
XFILL_4__3228_ gnd vdd FILL
XFILL_2__2243_ gnd vdd FILL
XFILL_4__3159_ gnd vdd FILL
XFILL_2__2174_ gnd vdd FILL
XFILL_8__2701_ gnd vdd FILL
XFILL_5__2923_ gnd vdd FILL
XFILL_8__2632_ gnd vdd FILL
XFILL_5__2854_ gnd vdd FILL
XFILL_8__2563_ gnd vdd FILL
XFILL_5__2785_ gnd vdd FILL
XFILL_8__2494_ gnd vdd FILL
XFILL_5__1805_ gnd vdd FILL
XFILL_5__1736_ gnd vdd FILL
XFILL_2__1958_ gnd vdd FILL
XFILL183750x70350 gnd vdd FILL
XFILL_3__3470_ gnd vdd FILL
XFILL_5__3406_ gnd vdd FILL
XFILL_2__1889_ gnd vdd FILL
XFILL_8__3115_ gnd vdd FILL
XFILL_3__2421_ gnd vdd FILL
XFILL_0__2712_ gnd vdd FILL
XFILL_8__3046_ gnd vdd FILL
XFILL_6__2130_ gnd vdd FILL
XFILL_0__2643_ gnd vdd FILL
XFILL_2__3559_ gnd vdd FILL
XFILL_3__2352_ gnd vdd FILL
XFILL_6__2061_ gnd vdd FILL
XFILL_3__2283_ gnd vdd FILL
XFILL_5__2219_ gnd vdd FILL
XFILL_0__2574_ gnd vdd FILL
XFILL_5__3199_ gnd vdd FILL
XFILL_6__2963_ gnd vdd FILL
XFILL_5_BUFX2_insert52 gnd vdd FILL
XFILL_5_BUFX2_insert41 gnd vdd FILL
XFILL_0__3126_ gnd vdd FILL
XFILL_5_BUFX2_insert85 gnd vdd FILL
XFILL_5_BUFX2_insert63 gnd vdd FILL
XFILL_5_BUFX2_insert74 gnd vdd FILL
XFILL_6__1914_ gnd vdd FILL
XFILL_5_BUFX2_insert96 gnd vdd FILL
XFILL_6__2894_ gnd vdd FILL
XFILL_0__3057_ gnd vdd FILL
XFILL_6__1845_ gnd vdd FILL
X_2705_ _2711_/B _2751_/B _2708_/C _2706_/C vdd gnd OAI21X1
X_2636_ _3241_/Q _2685_/B _2638_/A vdd gnd NAND2X1
XFILL_6__1776_ gnd vdd FILL
XFILL_0__2008_ gnd vdd FILL
XFILL_6__3515_ gnd vdd FILL
XFILL_3__1998_ gnd vdd FILL
XFILL_1__2821_ gnd vdd FILL
XFILL_4__2530_ gnd vdd FILL
X_2567_ _3254_/Q _2773_/A vdd gnd INVX1
XFILL_9__3224_ gnd vdd FILL
XFILL_6__3446_ gnd vdd FILL
X_2498_ _2659_/B _2574_/B _2498_/C _2499_/C vdd gnd OAI21X1
XFILL_4__2461_ gnd vdd FILL
XFILL_1__2752_ gnd vdd FILL
XFILL_6__3377_ gnd vdd FILL
XFILL_7__2170_ gnd vdd FILL
XFILL_1__1703_ gnd vdd FILL
XFILL_1__2683_ gnd vdd FILL
XFILL_3__2619_ gnd vdd FILL
XFILL_6__2328_ gnd vdd FILL
XFILL_3__3599_ gnd vdd FILL
XFILL_4__2392_ gnd vdd FILL
XFILL_6__2259_ gnd vdd FILL
X_3119_ _3121_/A _3125_/B _3335_/Q _3120_/C vdd gnd OAI21X1
XFILL_4__3013_ gnd vdd FILL
XFILL_7__1954_ gnd vdd FILL
XFILL_1__3166_ gnd vdd FILL
XFILL_1__3097_ gnd vdd FILL
XFILL_1__2117_ gnd vdd FILL
XFILL_7__1885_ gnd vdd FILL
XFILL_2__2930_ gnd vdd FILL
XFILL_1__2048_ gnd vdd FILL
XFILL_7__3555_ gnd vdd FILL
XFILL_2__2861_ gnd vdd FILL
XFILL_7__2506_ gnd vdd FILL
XFILL_5__2570_ gnd vdd FILL
XFILL_7__3486_ gnd vdd FILL
XFILL_2__2792_ gnd vdd FILL
XFILL_2__1812_ gnd vdd FILL
XFILL_4__2728_ gnd vdd FILL
XFILL_2__1743_ gnd vdd FILL
XFILL_7__2437_ gnd vdd FILL
XFILL_7__2368_ gnd vdd FILL
XFILL_4__2659_ gnd vdd FILL
XFILL_2__3413_ gnd vdd FILL
XFILL_5__3122_ gnd vdd FILL
XFILL_7__2299_ gnd vdd FILL
XFILL_5__3053_ gnd vdd FILL
XFILL_5__2004_ gnd vdd FILL
XFILL_2__2226_ gnd vdd FILL
XFILL_0__2290_ gnd vdd FILL
XFILL_8__1994_ gnd vdd FILL
XFILL183150x35250 gnd vdd FILL
XFILL_2__2157_ gnd vdd FILL
XFILL_3__2970_ gnd vdd FILL
XFILL_2__2088_ gnd vdd FILL
XFILL_5__2906_ gnd vdd FILL
XFILL_3__1921_ gnd vdd FILL
XFILL_8__2615_ gnd vdd FILL
XFILL_5__2837_ gnd vdd FILL
XFILL_8__3595_ gnd vdd FILL
X_3470_ _3470_/A _3470_/B _3472_/B vdd gnd NAND2X1
XFILL_3__1852_ gnd vdd FILL
XFILL_8__2546_ gnd vdd FILL
X_2421_ _3576_/Q _2427_/B _2421_/C _2422_/B vdd gnd AOI21X1
XFILL_3__1783_ gnd vdd FILL
XFILL_5__2768_ gnd vdd FILL
XFILL_8__2477_ gnd vdd FILL
XFILL_3__3522_ gnd vdd FILL
X_2352_ _2352_/A _2352_/B _2352_/C _2353_/A vdd gnd NAND3X1
XFILL_5__1719_ gnd vdd FILL
XFILL_5__2699_ gnd vdd FILL
XFILL183750x148350 gnd vdd FILL
X_2283_ _2328_/A _2283_/B _2286_/B vdd gnd NOR2X1
XFILL_6__3231_ gnd vdd FILL
XFILL_3__3453_ gnd vdd FILL
XFILL_6__3162_ gnd vdd FILL
XFILL_3__3384_ gnd vdd FILL
XFILL_3__2404_ gnd vdd FILL
XFILL_6__2113_ gnd vdd FILL
XFILL_8__3029_ gnd vdd FILL
XFILL_6__3093_ gnd vdd FILL
XFILL_3__2335_ gnd vdd FILL
XBUFX2_insert2 _1773_/Y _1987_/A vdd gnd BUFX2
XFILL_0__2626_ gnd vdd FILL
XFILL_6__2044_ gnd vdd FILL
XFILL_0__2557_ gnd vdd FILL
XFILL_3__2266_ gnd vdd FILL
XFILL_3__2197_ gnd vdd FILL
XFILL_0__2488_ gnd vdd FILL
XFILL_1__3020_ gnd vdd FILL
XFILL_6__2946_ gnd vdd FILL
XFILL_0__3109_ gnd vdd FILL
X_1998_ _2006_/A _1998_/B _2702_/B _1999_/C vdd gnd AOI21X1
XFILL_6__2877_ gnd vdd FILL
XFILL_4__1961_ gnd vdd FILL
XFILL_4__1892_ gnd vdd FILL
XFILL_6__1828_ gnd vdd FILL
XFILL_4__3562_ gnd vdd FILL
XFILL_6__1759_ gnd vdd FILL
X_3599_ _3599_/A DO[4] vdd gnd BUFX2
X_2619_ _2639_/A _2639_/B _2630_/A vdd gnd NAND2X1
XFILL_1__2804_ gnd vdd FILL
XFILL_4__2513_ gnd vdd FILL
XFILL_4__3493_ gnd vdd FILL
XFILL_6__3429_ gnd vdd FILL
XFILL_7__2222_ gnd vdd FILL
XFILL_1__2735_ gnd vdd FILL
XFILL_1_BUFX2_insert61 gnd vdd FILL
XFILL_1_BUFX2_insert50 gnd vdd FILL
XFILL_7__2153_ gnd vdd FILL
XFILL_4__2444_ gnd vdd FILL
XFILL_1_BUFX2_insert94 gnd vdd FILL
XFILL_1_BUFX2_insert83 gnd vdd FILL
XFILL_3_CLKBUF1_insert36 gnd vdd FILL
XFILL_4__2375_ gnd vdd FILL
XFILL_1_BUFX2_insert72 gnd vdd FILL
XFILL_1__2666_ gnd vdd FILL
XFILL_7__2084_ gnd vdd FILL
XFILL_1__2597_ gnd vdd FILL
XFILL_2__3060_ gnd vdd FILL
XFILL_2__2011_ gnd vdd FILL
XFILL_7__2986_ gnd vdd FILL
XFILL_1__3218_ gnd vdd FILL
XFILL_7__1937_ gnd vdd FILL
XFILL_1__3149_ gnd vdd FILL
XFILL_7__1868_ gnd vdd FILL
XFILL_8__2400_ gnd vdd FILL
XFILL_2__2913_ gnd vdd FILL
XFILL_8__3380_ gnd vdd FILL
XFILL_7__1799_ gnd vdd FILL
XFILL_5__2622_ gnd vdd FILL
XFILL_2__2844_ gnd vdd FILL
XFILL_7__3538_ gnd vdd FILL
XFILL_8__2331_ gnd vdd FILL
XFILL_7__3469_ gnd vdd FILL
XFILL_8__2262_ gnd vdd FILL
XFILL_5__2553_ gnd vdd FILL
XFILL_5__2484_ gnd vdd FILL
XFILL_2__2775_ gnd vdd FILL
XFILL_8__2193_ gnd vdd FILL
XFILL_2__1726_ gnd vdd FILL
XFILL_0__1790_ gnd vdd FILL
XFILL_0__3460_ gnd vdd FILL
XFILL_5__3105_ gnd vdd FILL
XFILL_0__3391_ gnd vdd FILL
XFILL_3__2120_ gnd vdd FILL
XFILL_0__2411_ gnd vdd FILL
XFILL_5__3036_ gnd vdd FILL
XFILL_0__2342_ gnd vdd FILL
X_2970_ _3308_/Q _2971_/A _2971_/C vdd gnd NAND2X1
XFILL_3__2051_ gnd vdd FILL
XFILL_8__1977_ gnd vdd FILL
XFILL_0__2273_ gnd vdd FILL
X_1921_ _2468_/A _1927_/B vdd gnd INVX1
XFILL_2__2209_ gnd vdd FILL
XFILL_2__3189_ gnd vdd FILL
XFILL_6__2800_ gnd vdd FILL
X_1852_ _1888_/A _1891_/A _3182_/B vdd gnd NAND2X1
XFILL_6__2731_ gnd vdd FILL
XFILL_3__2953_ gnd vdd FILL
X_1783_ _2442_/A _1783_/B _3190_/B vdd gnd NOR2X1
XFILL_3__2884_ gnd vdd FILL
X_3522_ _3522_/A _3522_/B _3539_/D vdd gnd XOR2X1
XFILL_3__1904_ gnd vdd FILL
XFILL_6__2662_ gnd vdd FILL
X_3453_ _3484_/B _3453_/B _3471_/A vdd gnd NAND2X1
XFILL_8__2529_ gnd vdd FILL
XFILL_6__2593_ gnd vdd FILL
XFILL_3__1835_ gnd vdd FILL
X_2404_ _2404_/A _2404_/B _2404_/C _3598_/A vdd gnd NAND3X1
X_3384_ _3384_/A _3384_/B _3384_/C _3519_/A vdd gnd OAI21X1
XFILL_3__1766_ gnd vdd FILL
XFILL_3__3505_ gnd vdd FILL
XFILL_3__1697_ gnd vdd FILL
X_2335_ _2335_/A _2335_/B _2337_/C vdd gnd AND2X2
XFILL_0__1988_ gnd vdd FILL
XFILL_6__3214_ gnd vdd FILL
X_2266_ _2921_/A _2911_/A vdd gnd INVX1
XFILL_3__3436_ gnd vdd FILL
XFILL_1__2520_ gnd vdd FILL
X_2197_ _2197_/A _2336_/B _2322_/A vdd gnd NOR2X1
XFILL_1__2451_ gnd vdd FILL
XFILL_6__3145_ gnd vdd FILL
XFILL_4__2160_ gnd vdd FILL
XFILL_6__3076_ gnd vdd FILL
XFILL_3__3367_ gnd vdd FILL
XFILL_0__2609_ gnd vdd FILL
XFILL_6__2027_ gnd vdd FILL
XFILL_3__2318_ gnd vdd FILL
XFILL_1__2382_ gnd vdd FILL
XFILL_0__3589_ gnd vdd FILL
XFILL_4__2091_ gnd vdd FILL
XFILL_3__2249_ gnd vdd FILL
XFILL_7__2840_ gnd vdd FILL
XFILL_1__3003_ gnd vdd FILL
XFILL_7__2771_ gnd vdd FILL
XFILL_6__2929_ gnd vdd FILL
XFILL_4__2993_ gnd vdd FILL
XFILL_7__1722_ gnd vdd FILL
XFILL_4__1944_ gnd vdd FILL
XFILL_4__1875_ gnd vdd FILL
XFILL_4__3545_ gnd vdd FILL
XFILL_4__3476_ gnd vdd FILL
XFILL_2__2560_ gnd vdd FILL
XFILL_7__2205_ gnd vdd FILL
XFILL_2__2491_ gnd vdd FILL
XFILL_1__2718_ gnd vdd FILL
XFILL_7__3185_ gnd vdd FILL
XFILL_4__2427_ gnd vdd FILL
XFILL_7__2136_ gnd vdd FILL
XFILL_1__2649_ gnd vdd FILL
XFILL_6_BUFX2_insert18 gnd vdd FILL
XFILL_4__2358_ gnd vdd FILL
XFILL_7__2067_ gnd vdd FILL
XFILL_4__2289_ gnd vdd FILL
XFILL_2__3112_ gnd vdd FILL
XFILL_8__2880_ gnd vdd FILL
XFILL_8__1900_ gnd vdd FILL
XFILL_2__3043_ gnd vdd FILL
XFILL_8__1831_ gnd vdd FILL
XFILL_8__3501_ gnd vdd FILL
XFILL_7__2969_ gnd vdd FILL
XFILL_8__1762_ gnd vdd FILL
XFILL_5__1984_ gnd vdd FILL
XFILL_8__1693_ gnd vdd FILL
XFILL_8__3432_ gnd vdd FILL
XFILL_0__2960_ gnd vdd FILL
XFILL_8__2314_ gnd vdd FILL
XFILL_0__1911_ gnd vdd FILL
XFILL_5__3585_ gnd vdd FILL
XFILL_5__2605_ gnd vdd FILL
XFILL_0__2891_ gnd vdd FILL
XFILL_2__2827_ gnd vdd FILL
XFILL_5__2536_ gnd vdd FILL
XFILL_0__1842_ gnd vdd FILL
XFILL_8__2245_ gnd vdd FILL
XFILL_2__2758_ gnd vdd FILL
XFILL_2__1709_ gnd vdd FILL
XFILL_5__2467_ gnd vdd FILL
XFILL_8__2176_ gnd vdd FILL
X_2120_ _2221_/A _2448_/B _2342_/A _2121_/C vdd gnd OAI21X1
XFILL_0__1773_ gnd vdd FILL
XFILL_0__3512_ gnd vdd FILL
XFILL_5__2398_ gnd vdd FILL
X_2051_ _2108_/A _3156_/B _2449_/C _2052_/B vdd gnd OAI21X1
XFILL_2__2689_ gnd vdd FILL
XFILL_3__3221_ gnd vdd FILL
XFILL_0__3443_ gnd vdd FILL
XFILL_3__3152_ gnd vdd FILL
XFILL_0__3374_ gnd vdd FILL
XFILL_3__3083_ gnd vdd FILL
XFILL_3__2103_ gnd vdd FILL
XFILL_3__2034_ gnd vdd FILL
X_2953_ reset _2957_/C _3305_/Q _2954_/C vdd gnd OAI21X1
XFILL_5__3019_ gnd vdd FILL
XFILL_0__2325_ gnd vdd FILL
XCLKBUF1_insert31 clk _3362_/CLK vdd gnd CLKBUF1
XFILL_0__2256_ gnd vdd FILL
X_1904_ _2221_/A _3189_/A _2433_/B vdd gnd NOR2X1
X_2884_ _2936_/B _2920_/A _2884_/C _3281_/D vdd gnd OAI21X1
XFILL_9__3472_ gnd vdd FILL
XFILL_0__2187_ gnd vdd FILL
X_1835_ _3187_/A _3176_/A _3176_/B _3025_/A vdd gnd NAND3X1
X_1766_ _2108_/A _3173_/B _2072_/B vdd gnd NOR2X1
XFILL_6__2714_ gnd vdd FILL
XFILL_3__2936_ gnd vdd FILL
X_3505_ _3505_/A _3506_/B vdd gnd INVX1
XFILL_1__1951_ gnd vdd FILL
XFILL_6__2645_ gnd vdd FILL
XFILL_3__2867_ gnd vdd FILL
X_1697_ _2985_/A _3292_/D vdd gnd INVX1
X_3436_ _3442_/A _3445_/A _3436_/C _3455_/C _3441_/B vdd gnd AOI22X1
XFILL_6__2576_ gnd vdd FILL
XFILL_1__1882_ gnd vdd FILL
XFILL_3__1818_ gnd vdd FILL
XFILL_3__2798_ gnd vdd FILL
X_3367_ _3571_/Q _3572_/Q _3368_/C vdd gnd NOR2X1
XFILL_1__3552_ gnd vdd FILL
X_2318_ _2318_/A _2318_/B _2318_/C _2321_/C vdd gnd NAND3X1
XFILL_3__1749_ gnd vdd FILL
XFILL_1__2503_ gnd vdd FILL
X_3298_ _3298_/D _3362_/R vdd _3362_/CLK _3298_/Q vdd gnd DFFSR
XFILL_1__3483_ gnd vdd FILL
X_2249_ _2249_/A _2930_/A _2921_/A vdd gnd NOR2X1
XFILL_6__3128_ gnd vdd FILL
XFILL_3__3419_ gnd vdd FILL
XFILL_4__2212_ gnd vdd FILL
XFILL_4__3192_ gnd vdd FILL
XFILL_4__2143_ gnd vdd FILL
XFILL_1__2434_ gnd vdd FILL
XFILL_6__3059_ gnd vdd FILL
XFILL_1__2365_ gnd vdd FILL
XFILL_4__2074_ gnd vdd FILL
XFILL_7__2823_ gnd vdd FILL
XFILL_1__2296_ gnd vdd FILL
XFILL_7__2754_ gnd vdd FILL
XFILL_4__2976_ gnd vdd FILL
XFILL_7__1705_ gnd vdd FILL
XFILL_7__2685_ gnd vdd FILL
XFILL_4__1927_ gnd vdd FILL
XFILL_2__1991_ gnd vdd FILL
XFILL_4__1858_ gnd vdd FILL
XFILL_5__3370_ gnd vdd FILL
XFILL_2__3592_ gnd vdd FILL
XFILL_2__2612_ gnd vdd FILL
XFILL_4__1789_ gnd vdd FILL
XFILL_4__3528_ gnd vdd FILL
XFILL_8__2030_ gnd vdd FILL
XFILL_5__2321_ gnd vdd FILL
XFILL_2__2543_ gnd vdd FILL
XFILL_4__3459_ gnd vdd FILL
XFILL_5__2252_ gnd vdd FILL
XFILL_5__2183_ gnd vdd FILL
XFILL_2__2474_ gnd vdd FILL
XFILL_7__3168_ gnd vdd FILL
XFILL_7__3099_ gnd vdd FILL
XFILL_7__2119_ gnd vdd FILL
XFILL_8__2932_ gnd vdd FILL
XFILL_8__2863_ gnd vdd FILL
XFILL_0__2110_ gnd vdd FILL
XFILL_0__3090_ gnd vdd FILL
XFILL_8__2794_ gnd vdd FILL
XFILL_2__3026_ gnd vdd FILL
XFILL_8__1814_ gnd vdd FILL
XFILL_0__2041_ gnd vdd FILL
XFILL_8__1745_ gnd vdd FILL
XFILL_5__1967_ gnd vdd FILL
XFILL_8__3415_ gnd vdd FILL
XFILL_5__1898_ gnd vdd FILL
XFILL_6__2430_ gnd vdd FILL
XFILL_3__2721_ gnd vdd FILL
XFILL_2_BUFX2_insert27 gnd vdd FILL
XFILL_2_BUFX2_insert16 gnd vdd FILL
XFILL_2_BUFX2_insert49 gnd vdd FILL
XFILL_0__2943_ gnd vdd FILL
XFILL_3__2652_ gnd vdd FILL
XFILL_6__2361_ gnd vdd FILL
XFILL_0__2874_ gnd vdd FILL
X_3221_ _3221_/A _3227_/B _3221_/C _3358_/D vdd gnd OAI21X1
XFILL_5__3499_ gnd vdd FILL
XFILL_0__1825_ gnd vdd FILL
XFILL_8__2228_ gnd vdd FILL
XFILL_3__2583_ gnd vdd FILL
X_3152_ _3166_/C _3165_/A _3152_/C _3153_/B vdd gnd OAI21X1
XFILL_5__2519_ gnd vdd FILL
XFILL_6__2292_ gnd vdd FILL
X_2103_ _3160_/B _3146_/A _2104_/A vdd gnd NAND2X1
X_3083_ _3083_/A _3083_/B _3084_/C vdd gnd NAND2X1
XFILL_0__1756_ gnd vdd FILL
XFILL_8__2159_ gnd vdd FILL
X_2034_ _2957_/A _3302_/Q _2889_/C _2035_/C vdd gnd OAI21X1
XFILL_3__3204_ gnd vdd FILL
XFILL_3__3135_ gnd vdd FILL
XFILL_0__3426_ gnd vdd FILL
XFILL_1__2150_ gnd vdd FILL
XFILL_3__3066_ gnd vdd FILL
XFILL_0__2308_ gnd vdd FILL
XFILL_9__1854_ gnd vdd FILL
X_2936_ _3023_/A _2936_/B _2936_/C _2936_/D _3289_/D vdd gnd AOI22X1
XFILL_3__2017_ gnd vdd FILL
XFILL_1__2081_ gnd vdd FILL
X_2867_ _2867_/A _2887_/B _2868_/A vdd gnd AND2X2
XFILL_0__2239_ gnd vdd FILL
XFILL_4__2830_ gnd vdd FILL
X_1818_ _3291_/D _3043_/A vdd gnd INVX2
X_2798_ _2902_/A _2798_/B _2803_/D vdd gnd OR2X2
XFILL_4__2761_ gnd vdd FILL
XFILL_3__2919_ gnd vdd FILL
XFILL_1__2983_ gnd vdd FILL
XFILL_7__2470_ gnd vdd FILL
XFILL_4__1712_ gnd vdd FILL
X_1749_ _2430_/A _2430_/B _2437_/A _1750_/A vdd gnd OAI21X1
XFILL_8_CLKBUF1_insert36 gnd vdd FILL
XFILL_4__2692_ gnd vdd FILL
XFILL_1__1934_ gnd vdd FILL
XFILL_6__2628_ gnd vdd FILL
XFILL_1__1865_ gnd vdd FILL
X_3419_ _3442_/B _3420_/A _3466_/B _3420_/C vdd gnd OAI21X1
XFILL_6__2559_ gnd vdd FILL
XFILL_7__3022_ gnd vdd FILL
XFILL_1_BUFX2_insert2 gnd vdd FILL
XFILL_1__1796_ gnd vdd FILL
XFILL_1__3535_ gnd vdd FILL
XFILL_1__3466_ gnd vdd FILL
XFILL_1__2417_ gnd vdd FILL
XFILL_4__3175_ gnd vdd FILL
XFILL_1__3397_ gnd vdd FILL
XFILL_2__2190_ gnd vdd FILL
XFILL_4__2126_ gnd vdd FILL
XFILL_1__2348_ gnd vdd FILL
XFILL_4__2057_ gnd vdd FILL
XFILL_1__2279_ gnd vdd FILL
XFILL_5__2870_ gnd vdd FILL
XFILL_7__2806_ gnd vdd FILL
XFILL_5__1821_ gnd vdd FILL
XFILL_7__2737_ gnd vdd FILL
XFILL_4__2959_ gnd vdd FILL
XFILL_5__1752_ gnd vdd FILL
XFILL_2__1974_ gnd vdd FILL
XFILL_7__2668_ gnd vdd FILL
XFILL_7__2599_ gnd vdd FILL
XFILL_8__3200_ gnd vdd FILL
XFILL_8__3131_ gnd vdd FILL
XFILL_5__3422_ gnd vdd FILL
XFILL_8__3062_ gnd vdd FILL
XFILL_5__2304_ gnd vdd FILL
XFILL_8__2013_ gnd vdd FILL
XFILL_0__2590_ gnd vdd FILL
XFILL_2__2526_ gnd vdd FILL
XFILL_5__2235_ gnd vdd FILL
XFILL_2__2457_ gnd vdd FILL
XFILL_5__2166_ gnd vdd FILL
XFILL_2__2388_ gnd vdd FILL
XFILL_0__3211_ gnd vdd FILL
XFILL_5__2097_ gnd vdd FILL
XFILL_8__2915_ gnd vdd FILL
XFILL_4_BUFX2_insert6 gnd vdd FILL
XFILL_0__3142_ gnd vdd FILL
XFILL_8__2846_ gnd vdd FILL
XFILL_6__1930_ gnd vdd FILL
XFILL_2__3009_ gnd vdd FILL
XFILL_0__3073_ gnd vdd FILL
XFILL_6__1861_ gnd vdd FILL
X_2721_ _2732_/C _2721_/B _2722_/A vdd gnd NAND2X1
XFILL_0__2024_ gnd vdd FILL
XFILL_6__3600_ gnd vdd FILL
XFILL_8__2777_ gnd vdd FILL
XFILL_6__3531_ gnd vdd FILL
XFILL_5__2999_ gnd vdd FILL
XFILL_6__1792_ gnd vdd FILL
XFILL_8__1728_ gnd vdd FILL
X_2652_ _2659_/B _2671_/B _2656_/D _2653_/C vdd gnd OAI21X1
X_2583_ _3165_/A _3166_/A _2583_/C _2609_/A vdd gnd AOI21X1
XFILL_6__3462_ gnd vdd FILL
XFILL_3__2704_ gnd vdd FILL
XFILL_0__2926_ gnd vdd FILL
XFILL_6__3393_ gnd vdd FILL
XFILL_6__2413_ gnd vdd FILL
XFILL_6__2344_ gnd vdd FILL
X_3204_ _3214_/A _3214_/B _3350_/Q _3205_/C vdd gnd OAI21X1
XFILL_3__2635_ gnd vdd FILL
XFILL_0__2857_ gnd vdd FILL
XFILL_3__2566_ gnd vdd FILL
X_3135_ _3135_/A _3143_/B _3135_/C _3343_/D vdd gnd OAI21X1
XFILL_0__2788_ gnd vdd FILL
XFILL_6__2275_ gnd vdd FILL
XFILL_0__1808_ gnd vdd FILL
X_3066_ _3090_/A _3137_/A _3066_/C _3319_/D vdd gnd OAI21X1
XFILL_3__2497_ gnd vdd FILL
XFILL_0__1739_ gnd vdd FILL
X_2017_ _2033_/A _3304_/Q _2018_/C vdd gnd NAND2X1
XFILL_1__2202_ gnd vdd FILL
XFILL_3__3118_ gnd vdd FILL
XFILL_0__3409_ gnd vdd FILL
XFILL_1__3182_ gnd vdd FILL
XFILL_7__1970_ gnd vdd FILL
XFILL_3__3049_ gnd vdd FILL
XFILL_1__2133_ gnd vdd FILL
X_2919_ _2919_/A _2919_/B _2919_/C _3287_/D vdd gnd AOI21X1
XFILL_1__2064_ gnd vdd FILL
XFILL_4__2813_ gnd vdd FILL
XFILL_7__2522_ gnd vdd FILL
XFILL_7__2453_ gnd vdd FILL
XFILL_4__2744_ gnd vdd FILL
XFILL_1__2966_ gnd vdd FILL
XFILL_9__3369_ gnd vdd FILL
XFILL_4__2675_ gnd vdd FILL
XFILL_1__1917_ gnd vdd FILL
XFILL_1__2897_ gnd vdd FILL
XFILL_7__2384_ gnd vdd FILL
XFILL_2__1690_ gnd vdd FILL
XFILL_1__1848_ gnd vdd FILL
XFILL_1__1779_ gnd vdd FILL
XFILL_1__3518_ gnd vdd FILL
XFILL_2__2311_ gnd vdd FILL
XFILL_7__3005_ gnd vdd FILL
XFILL_5__2020_ gnd vdd FILL
XFILL_4__3227_ gnd vdd FILL
XFILL_1__3449_ gnd vdd FILL
XFILL_2__2242_ gnd vdd FILL
XFILL_4__3158_ gnd vdd FILL
XFILL_2__2173_ gnd vdd FILL
XFILL_4__2109_ gnd vdd FILL
XFILL_4__3089_ gnd vdd FILL
XFILL_8__2700_ gnd vdd FILL
XFILL_5__2922_ gnd vdd FILL
XFILL_8__2631_ gnd vdd FILL
XFILL_5__2853_ gnd vdd FILL
XFILL_5__1804_ gnd vdd FILL
XFILL_8__2562_ gnd vdd FILL
XFILL_5__2784_ gnd vdd FILL
XFILL_8__2493_ gnd vdd FILL
XFILL_5__1735_ gnd vdd FILL
XFILL_2__1957_ gnd vdd FILL
XFILL_5__3405_ gnd vdd FILL
XFILL_2__1888_ gnd vdd FILL
XFILL_8__3114_ gnd vdd FILL
XFILL_3__2420_ gnd vdd FILL
XFILL_0__2711_ gnd vdd FILL
XFILL_8__3045_ gnd vdd FILL
XFILL_3__2351_ gnd vdd FILL
XFILL_0__2642_ gnd vdd FILL
XFILL_2__3558_ gnd vdd FILL
XFILL_6__2060_ gnd vdd FILL
XFILL_0__2573_ gnd vdd FILL
XFILL_2__3489_ gnd vdd FILL
XFILL_3__2282_ gnd vdd FILL
XFILL_5__2218_ gnd vdd FILL
XFILL_2__2509_ gnd vdd FILL
XFILL_5__3198_ gnd vdd FILL
XFILL_5__2149_ gnd vdd FILL
XFILL_5_BUFX2_insert20 gnd vdd FILL
XFILL_6__2962_ gnd vdd FILL
XFILL_5_BUFX2_insert42 gnd vdd FILL
XFILL_5_BUFX2_insert53 gnd vdd FILL
XFILL_0__3125_ gnd vdd FILL
XFILL_5_BUFX2_insert64 gnd vdd FILL
XFILL_5_BUFX2_insert75 gnd vdd FILL
XFILL_6__1913_ gnd vdd FILL
XFILL_5_BUFX2_insert86 gnd vdd FILL
XFILL_5_BUFX2_insert97 gnd vdd FILL
XFILL_8__2829_ gnd vdd FILL
XFILL_6__2893_ gnd vdd FILL
XFILL_0__3056_ gnd vdd FILL
XFILL_6__1844_ gnd vdd FILL
X_2704_ _2704_/A _2704_/B _2704_/C _2708_/C vdd gnd NOR3X1
XFILL_6__1775_ gnd vdd FILL
X_2635_ _2635_/A _2635_/B _2635_/C _2641_/D vdd gnd AOI21X1
XFILL_0__2007_ gnd vdd FILL
XFILL_1__2820_ gnd vdd FILL
XFILL_6__3514_ gnd vdd FILL
XFILL_3__1997_ gnd vdd FILL
XFILL_6__3445_ gnd vdd FILL
X_2566_ _2768_/B _2574_/B _2566_/C _3585_/A vdd gnd OAI21X1
X_2497_ _2497_/A _2497_/B _2498_/C vdd gnd AND2X2
XFILL_4__2460_ gnd vdd FILL
XFILL_1__2751_ gnd vdd FILL
XFILL_0__2909_ gnd vdd FILL
XFILL_6__3376_ gnd vdd FILL
XFILL_1__1702_ gnd vdd FILL
XFILL_1__2682_ gnd vdd FILL
XFILL_3__2618_ gnd vdd FILL
XFILL_9__2105_ gnd vdd FILL
XFILL_6__2327_ gnd vdd FILL
XFILL_3__3598_ gnd vdd FILL
XFILL_4__2391_ gnd vdd FILL
X_3118_ _3135_/A _3126_/B _3118_/C _3334_/D vdd gnd OAI21X1
XFILL_6__2258_ gnd vdd FILL
XFILL_3__2549_ gnd vdd FILL
XFILL_6__2189_ gnd vdd FILL
XFILL_4__3012_ gnd vdd FILL
X_3049_ _3050_/A _3050_/B _3052_/D vdd gnd NAND2X1
XFILL_7__1953_ gnd vdd FILL
XFILL_1__3165_ gnd vdd FILL
XFILL_1__2116_ gnd vdd FILL
XFILL_1__3096_ gnd vdd FILL
XFILL_7__1884_ gnd vdd FILL
XFILL_1__2047_ gnd vdd FILL
XFILL_7__3554_ gnd vdd FILL
XFILL_2__2860_ gnd vdd FILL
XFILL_7__2505_ gnd vdd FILL
XFILL_7__3485_ gnd vdd FILL
XFILL_2__2791_ gnd vdd FILL
XFILL_4__2727_ gnd vdd FILL
XFILL_2__1811_ gnd vdd FILL
XFILL_1__2949_ gnd vdd FILL
XFILL_2__1742_ gnd vdd FILL
XFILL_7__2436_ gnd vdd FILL
XFILL_7__2367_ gnd vdd FILL
XFILL_4__2658_ gnd vdd FILL
XFILL_2__3412_ gnd vdd FILL
XFILL_4__2589_ gnd vdd FILL
XFILL_5__3121_ gnd vdd FILL
XFILL_7__2298_ gnd vdd FILL
XFILL_5__3052_ gnd vdd FILL
XFILL_5__2003_ gnd vdd FILL
XFILL_2__2225_ gnd vdd FILL
XFILL_8__1993_ gnd vdd FILL
XFILL_2__2156_ gnd vdd FILL
XFILL_5__2905_ gnd vdd FILL
XFILL_2__2087_ gnd vdd FILL
XFILL_3__1920_ gnd vdd FILL
XFILL_8__3594_ gnd vdd FILL
XFILL_8__2614_ gnd vdd FILL
XFILL_5__2836_ gnd vdd FILL
XFILL_8__2545_ gnd vdd FILL
X_2420_ _2668_/B _2426_/B _2420_/C _2421_/C vdd gnd OAI21X1
XFILL_3__1851_ gnd vdd FILL
XFILL_5__2767_ gnd vdd FILL
XFILL_2__2989_ gnd vdd FILL
XFILL_8__2476_ gnd vdd FILL
XFILL_5__1718_ gnd vdd FILL
XFILL_3__1782_ gnd vdd FILL
XFILL_3__3521_ gnd vdd FILL
X_2351_ _2351_/A _2351_/B _2352_/C vdd gnd NOR2X1
XFILL_5__2698_ gnd vdd FILL
X_2282_ _2282_/A _2286_/A vdd gnd INVX1
XFILL_6__3230_ gnd vdd FILL
XFILL_3__3452_ gnd vdd FILL
XFILL_6__3161_ gnd vdd FILL
XFILL_6__2112_ gnd vdd FILL
XFILL_3__3383_ gnd vdd FILL
XFILL_3__2403_ gnd vdd FILL
XFILL_8__3028_ gnd vdd FILL
XFILL_6__3092_ gnd vdd FILL
XFILL_3__2334_ gnd vdd FILL
XFILL_0__2625_ gnd vdd FILL
XFILL_6__2043_ gnd vdd FILL
XBUFX2_insert3 _1773_/Y _3160_/B vdd gnd BUFX2
XFILL_0__2556_ gnd vdd FILL
XFILL_3__2265_ gnd vdd FILL
XFILL_0__2487_ gnd vdd FILL
XFILL_3__2196_ gnd vdd FILL
XFILL_9__2723_ gnd vdd FILL
XFILL_6__2945_ gnd vdd FILL
X_1997_ _3310_/Q _2008_/A _2623_/B _2702_/B vdd gnd OAI21X1
XFILL_0__3108_ gnd vdd FILL
XFILL_6__2876_ gnd vdd FILL
XFILL_4__1960_ gnd vdd FILL
XFILL_0__3039_ gnd vdd FILL
XFILL_6__1827_ gnd vdd FILL
XFILL_4__1891_ gnd vdd FILL
XFILL_4__3561_ gnd vdd FILL
X_3598_ _3598_/A DO[3] vdd gnd BUFX2
X_2618_ _2639_/A _2639_/B _2621_/C vdd gnd NOR2X1
XFILL_6__1758_ gnd vdd FILL
XFILL_1__2803_ gnd vdd FILL
XFILL_6__1689_ gnd vdd FILL
X_2549_ _3360_/Q _2691_/A _2549_/C _2550_/C vdd gnd AOI21X1
XFILL_4__2512_ gnd vdd FILL
XFILL_4__3492_ gnd vdd FILL
XFILL_6__3428_ gnd vdd FILL
XFILL_1__2734_ gnd vdd FILL
XFILL_7__2221_ gnd vdd FILL
XFILL_1_BUFX2_insert51 gnd vdd FILL
XFILL_7__2152_ gnd vdd FILL
XFILL_1_BUFX2_insert40 gnd vdd FILL
XFILL_4__2443_ gnd vdd FILL
XFILL_3_CLKBUF1_insert37 gnd vdd FILL
XFILL_1_BUFX2_insert95 gnd vdd FILL
XFILL_1_BUFX2_insert84 gnd vdd FILL
XFILL_1_BUFX2_insert62 gnd vdd FILL
XFILL_1_BUFX2_insert73 gnd vdd FILL
XFILL_4__2374_ gnd vdd FILL
XFILL_1__2665_ gnd vdd FILL
XFILL_7__2083_ gnd vdd FILL
XFILL_1__2596_ gnd vdd FILL
XFILL_2__2010_ gnd vdd FILL
XFILL_1_CLKBUF1_insert30 gnd vdd FILL
XFILL_7__2985_ gnd vdd FILL
XFILL_1__3217_ gnd vdd FILL
XFILL_7__1936_ gnd vdd FILL
XFILL_1__3148_ gnd vdd FILL
XFILL_7__1867_ gnd vdd FILL
XFILL_1__3079_ gnd vdd FILL
XFILL_2__2912_ gnd vdd FILL
XFILL_5__2621_ gnd vdd FILL
XFILL_7__1798_ gnd vdd FILL
XFILL_2__2843_ gnd vdd FILL
XFILL_7__3537_ gnd vdd FILL
XFILL_8__2330_ gnd vdd FILL
XFILL_7__3468_ gnd vdd FILL
XFILL_8__2261_ gnd vdd FILL
XFILL_5__2552_ gnd vdd FILL
XFILL_7__2419_ gnd vdd FILL
XFILL_5__2483_ gnd vdd FILL
XFILL_2__2774_ gnd vdd FILL
XFILL_7__3399_ gnd vdd FILL
XFILL_8__2192_ gnd vdd FILL
XFILL_2__1725_ gnd vdd FILL
XFILL_5__3104_ gnd vdd FILL
XFILL_0__3390_ gnd vdd FILL
XFILL_0__2410_ gnd vdd FILL
XFILL_5__3035_ gnd vdd FILL
XFILL_0__2341_ gnd vdd FILL
XFILL_3__2050_ gnd vdd FILL
XFILL_8__1976_ gnd vdd FILL
XFILL_0__2272_ gnd vdd FILL
X_1920_ _1920_/A _1920_/B _1920_/C _2468_/A vdd gnd NAND3X1
XFILL_2__2208_ gnd vdd FILL
XFILL_2__3188_ gnd vdd FILL
XFILL_2__2139_ gnd vdd FILL
X_1851_ _3235_/Q _3236_/Q _1888_/A vdd gnd NOR2X1
XFILL_6__2730_ gnd vdd FILL
XFILL_3__2952_ gnd vdd FILL
X_3521_ _3521_/A _3521_/B _3522_/B vdd gnd NAND2X1
X_1782_ _1987_/A _1782_/B _3192_/A vdd gnd NAND2X1
XFILL_6__2661_ gnd vdd FILL
XFILL_5__2819_ gnd vdd FILL
XFILL_3__2883_ gnd vdd FILL
XFILL_9__2370_ gnd vdd FILL
XFILL_3__1903_ gnd vdd FILL
X_3452_ _3485_/A _3493_/B _3493_/A _3497_/A vdd gnd OAI21X1
XFILL_8__2528_ gnd vdd FILL
XFILL_3__1834_ gnd vdd FILL
XFILL_6__2592_ gnd vdd FILL
X_3383_ _3565_/A _3383_/B _3459_/A _3384_/A vdd gnd OAI21X1
X_2403_ _3573_/Q _2427_/B _2403_/C _2404_/B vdd gnd AOI21X1
XFILL_8__2459_ gnd vdd FILL
X_2334_ _2334_/A _2334_/B _2335_/A vdd gnd NOR2X1
XFILL_3__1765_ gnd vdd FILL
XFILL_3__3504_ gnd vdd FILL
XFILL_3__1696_ gnd vdd FILL
XFILL_6__3213_ gnd vdd FILL
XFILL_0__1987_ gnd vdd FILL
X_2265_ _2894_/A _2933_/B _2792_/C _2269_/C vdd gnd OAI21X1
XFILL_3__3435_ gnd vdd FILL
XFILL_8_BUFX2_insert90 gnd vdd FILL
X_2196_ _2896_/B _2196_/B _2196_/C _2197_/A vdd gnd OAI21X1
XFILL_1__2450_ gnd vdd FILL
XFILL_6__3144_ gnd vdd FILL
XFILL_6__3075_ gnd vdd FILL
XFILL_3__3366_ gnd vdd FILL
XFILL_1__2381_ gnd vdd FILL
XFILL_0__2608_ gnd vdd FILL
XFILL_6__2026_ gnd vdd FILL
XFILL_3__2317_ gnd vdd FILL
XFILL_4__2090_ gnd vdd FILL
XFILL_0__3588_ gnd vdd FILL
XFILL_3__2248_ gnd vdd FILL
XFILL_0__2539_ gnd vdd FILL
XFILL_3__2179_ gnd vdd FILL
XFILL_1__3002_ gnd vdd FILL
XFILL_7__2770_ gnd vdd FILL
XFILL_6__2928_ gnd vdd FILL
XFILL_4__2992_ gnd vdd FILL
XFILL_7__1721_ gnd vdd FILL
XFILL_4__1943_ gnd vdd FILL
XFILL_6__2859_ gnd vdd FILL
XFILL_4__1874_ gnd vdd FILL
XFILL_4__3544_ gnd vdd FILL
XFILL_4__3475_ gnd vdd FILL
XFILL_7__2204_ gnd vdd FILL
XFILL_4__2426_ gnd vdd FILL
XFILL_2__2490_ gnd vdd FILL
XFILL_7__3184_ gnd vdd FILL
XFILL_1__2717_ gnd vdd FILL
XFILL_7__2135_ gnd vdd FILL
XFILL_1__2648_ gnd vdd FILL
XFILL_7__2066_ gnd vdd FILL
XFILL_4__2357_ gnd vdd FILL
XFILL_1__2579_ gnd vdd FILL
XFILL_4__2288_ gnd vdd FILL
XFILL_6_BUFX2_insert19 gnd vdd FILL
XFILL_2__3111_ gnd vdd FILL
XFILL_2__3042_ gnd vdd FILL
XFILL_8__1830_ gnd vdd FILL
XFILL_7__2968_ gnd vdd FILL
XFILL_8__1761_ gnd vdd FILL
XFILL_8__3500_ gnd vdd FILL
XFILL_7__1919_ gnd vdd FILL
XFILL_5__1983_ gnd vdd FILL
XFILL_7__2899_ gnd vdd FILL
XFILL_8__1692_ gnd vdd FILL
XFILL_8__3431_ gnd vdd FILL
XFILL_8__2313_ gnd vdd FILL
XFILL_5__3584_ gnd vdd FILL
XFILL_5__2604_ gnd vdd FILL
XFILL_0__1910_ gnd vdd FILL
XFILL_0__2890_ gnd vdd FILL
XFILL_2__2826_ gnd vdd FILL
XFILL_5__2535_ gnd vdd FILL
XFILL_8__2244_ gnd vdd FILL
XFILL_2__2757_ gnd vdd FILL
XFILL_0__1841_ gnd vdd FILL
XFILL_0__1772_ gnd vdd FILL
XFILL_2__1708_ gnd vdd FILL
XFILL_5__2466_ gnd vdd FILL
XFILL_8__2175_ gnd vdd FILL
XFILL_0__3511_ gnd vdd FILL
XFILL_5__2397_ gnd vdd FILL
XFILL_2__2688_ gnd vdd FILL
XFILL_3__3220_ gnd vdd FILL
X_2050_ _3157_/A _3144_/A _2449_/C vdd gnd NAND2X1
XFILL_0__3442_ gnd vdd FILL
XFILL182550x140550 gnd vdd FILL
XFILL_3__3151_ gnd vdd FILL
XFILL_3__3082_ gnd vdd FILL
XFILL_0__3373_ gnd vdd FILL
XFILL_5__3018_ gnd vdd FILL
XFILL_3__2102_ gnd vdd FILL
XFILL_3__2033_ gnd vdd FILL
X_2952_ _2952_/A _2956_/B _2952_/C _3304_/D vdd gnd OAI21X1
XFILL_0__2324_ gnd vdd FILL
XFILL_0__2255_ gnd vdd FILL
XCLKBUF1_insert32 clk _3284_/CLK vdd gnd CLKBUF1
X_1903_ _1903_/A _1903_/B _1986_/A vdd gnd NOR2X1
X_2883_ _2906_/A _2906_/B _3281_/Q _2884_/C vdd gnd OAI21X1
XFILL_8__1959_ gnd vdd FILL
XFILL_0__2186_ gnd vdd FILL
XFILL_6__2713_ gnd vdd FILL
X_1834_ _2602_/A _3157_/B _3176_/B vdd gnd NAND2X1
XFILL_3__2935_ gnd vdd FILL
X_1765_ _3166_/C _3165_/A _1765_/Y vdd gnd NAND2X1
X_3504_ _3514_/A _3514_/B _3508_/B _3505_/A vdd gnd OAI21X1
XFILL_1__1950_ gnd vdd FILL
XFILL_6__2644_ gnd vdd FILL
XFILL_3__2866_ gnd vdd FILL
X_3435_ _3442_/A _3438_/A _3453_/B _3436_/C vdd gnd NAND3X1
XFILL_6__2575_ gnd vdd FILL
X_1696_ _2768_/A DI[2] _1696_/C _2985_/A vdd gnd OAI21X1
XFILL_1__1881_ gnd vdd FILL
XFILL_3__2797_ gnd vdd FILL
XFILL_3__1817_ gnd vdd FILL
X_3366_ _3577_/Q _3576_/Q _3368_/B vdd gnd NOR2X1
XFILL_3__1748_ gnd vdd FILL
XFILL_1__3551_ gnd vdd FILL
X_2317_ _2317_/A _2324_/A vdd gnd INVX1
X_3297_ _3297_/D vdd _3353_/R _3578_/CLK _3297_/Q vdd gnd DFFSR
X_2248_ _2932_/A _2930_/A vdd gnd INVX1
XFILL_1__2502_ gnd vdd FILL
XFILL_1__3482_ gnd vdd FILL
XFILL_6__3127_ gnd vdd FILL
XFILL_3__3418_ gnd vdd FILL
XFILL_4__2211_ gnd vdd FILL
XFILL_4__3191_ gnd vdd FILL
X_2179_ _2179_/A _2889_/C _2915_/A vdd gnd AND2X2
XFILL_4__2142_ gnd vdd FILL
XFILL_1__2433_ gnd vdd FILL
XFILL_6__3058_ gnd vdd FILL
XFILL_1__2364_ gnd vdd FILL
XFILL_1__2295_ gnd vdd FILL
XFILL_4__2073_ gnd vdd FILL
XFILL_6__2009_ gnd vdd FILL
XFILL_7__2822_ gnd vdd FILL
XFILL_7__2753_ gnd vdd FILL
XFILL_4__2975_ gnd vdd FILL
XFILL_7__1704_ gnd vdd FILL
XFILL_7__2684_ gnd vdd FILL
XFILL_4__1926_ gnd vdd FILL
XFILL_2__1990_ gnd vdd FILL
XFILL_4__1857_ gnd vdd FILL
XFILL_4__3527_ gnd vdd FILL
XFILL_2__3591_ gnd vdd FILL
XFILL_5__2320_ gnd vdd FILL
XFILL_2__2611_ gnd vdd FILL
XFILL_4__1788_ gnd vdd FILL
XFILL_2__2542_ gnd vdd FILL
XFILL_4__3458_ gnd vdd FILL
XFILL_5__2251_ gnd vdd FILL
XFILL_7__3167_ gnd vdd FILL
XFILL_4__3389_ gnd vdd FILL
XFILL_5__2182_ gnd vdd FILL
XFILL_7__2118_ gnd vdd FILL
XFILL_2__2473_ gnd vdd FILL
XFILL_4__2409_ gnd vdd FILL
XFILL_7__3098_ gnd vdd FILL
XFILL_8__2931_ gnd vdd FILL
XFILL_7__2049_ gnd vdd FILL
XFILL_8__2862_ gnd vdd FILL
XFILL_8__1813_ gnd vdd FILL
XFILL_0__2040_ gnd vdd FILL
XFILL_8__2793_ gnd vdd FILL
XFILL_2__3025_ gnd vdd FILL
XFILL_8__1744_ gnd vdd FILL
XFILL_5__1966_ gnd vdd FILL
XFILL_8__3414_ gnd vdd FILL
XFILL_5__1897_ gnd vdd FILL
XFILL_2_BUFX2_insert17 gnd vdd FILL
XFILL_3__2720_ gnd vdd FILL
XFILL_0__2942_ gnd vdd FILL
XFILL_2_BUFX2_insert39 gnd vdd FILL
XFILL_3__2651_ gnd vdd FILL
XFILL_6__2360_ gnd vdd FILL
XFILL_2__2809_ gnd vdd FILL
XFILL_0__2873_ gnd vdd FILL
X_3220_ _3581_/A _3227_/B _3221_/C vdd gnd NAND2X1
XFILL_5__3498_ gnd vdd FILL
XFILL_8__2227_ gnd vdd FILL
XFILL_0__1824_ gnd vdd FILL
XFILL_5__2518_ gnd vdd FILL
X_3151_ _3151_/A _3151_/B _3151_/C _3192_/B vdd gnd OAI21X1
XFILL_3__2582_ gnd vdd FILL
XFILL_6__2291_ gnd vdd FILL
XFILL_5__2449_ gnd vdd FILL
X_2102_ _3160_/B _3190_/B _2441_/B vdd gnd NAND2X1
X_3082_ _3090_/A _3141_/A _3082_/C _3321_/D vdd gnd OAI21X1
XFILL_0__1755_ gnd vdd FILL
XFILL_8__2158_ gnd vdd FILL
X_2033_ _2033_/A _2957_/A vdd gnd INVX1
XFILL_8__2089_ gnd vdd FILL
XFILL_3__3203_ gnd vdd FILL
XFILL_3__3134_ gnd vdd FILL
XFILL_0__3425_ gnd vdd FILL
XFILL_3__3065_ gnd vdd FILL
XFILL_0__2307_ gnd vdd FILL
XFILL182250x35250 gnd vdd FILL
X_2935_ _2935_/A _2935_/B _2936_/D vdd gnd NOR2X1
XFILL_1__2080_ gnd vdd FILL
XFILL_3__2016_ gnd vdd FILL
X_2866_ _2866_/A _2919_/B _2866_/C _3275_/D vdd gnd AOI21X1
XFILL_0__2238_ gnd vdd FILL
XFILL_0__2169_ gnd vdd FILL
X_1817_ _3240_/Q _2621_/B vdd gnd INVX2
X_2797_ _2910_/B _2797_/B _2813_/C vdd gnd NAND2X1
XFILL_4__2760_ gnd vdd FILL
XFILL_3__2918_ gnd vdd FILL
XFILL_8_CLKBUF1_insert37 gnd vdd FILL
XFILL_1__2982_ gnd vdd FILL
XFILL_4__1711_ gnd vdd FILL
X_1748_ _3160_/C _2430_/B vdd gnd INVX1
XFILL_4__2691_ gnd vdd FILL
XFILL_6__2627_ gnd vdd FILL
XFILL_3__2849_ gnd vdd FILL
XFILL_1__1933_ gnd vdd FILL
XFILL_9__2267_ gnd vdd FILL
X_3418_ _3418_/A _3418_/B _3418_/C _3508_/A vdd gnd OAI21X1
XFILL_1__1864_ gnd vdd FILL
XFILL_6__2558_ gnd vdd FILL
XFILL_6__2489_ gnd vdd FILL
X_3349_ _3349_/D vdd _3355_/R _3355_/CLK _3349_/Q vdd gnd DFFSR
XFILL_1__3603_ gnd vdd FILL
XFILL_7__3021_ gnd vdd FILL
XFILL_1_BUFX2_insert3 gnd vdd FILL
XFILL_1__1795_ gnd vdd FILL
XFILL_1__3534_ gnd vdd FILL
XFILL_6_CLKBUF1_insert30 gnd vdd FILL
XFILL_1__3465_ gnd vdd FILL
XFILL_1__2416_ gnd vdd FILL
XFILL_4__3174_ gnd vdd FILL
XFILL_1__3396_ gnd vdd FILL
XFILL_4__2125_ gnd vdd FILL
XFILL_1__2347_ gnd vdd FILL
XFILL_4__2056_ gnd vdd FILL
XFILL_1__2278_ gnd vdd FILL
XFILL_7__2805_ gnd vdd FILL
XFILL_5__1820_ gnd vdd FILL
XFILL_7__2736_ gnd vdd FILL
XFILL_4__2958_ gnd vdd FILL
XFILL_5__1751_ gnd vdd FILL
XFILL_2__1973_ gnd vdd FILL
XFILL_7__2667_ gnd vdd FILL
XFILL_4__1909_ gnd vdd FILL
XFILL_4__2889_ gnd vdd FILL
XFILL_5__3421_ gnd vdd FILL
XFILL_7__2598_ gnd vdd FILL
XFILL_8__3130_ gnd vdd FILL
XFILL_8__3061_ gnd vdd FILL
XFILL_8__2012_ gnd vdd FILL
XFILL_5__2303_ gnd vdd FILL
XFILL_7__3219_ gnd vdd FILL
XFILL_2__2525_ gnd vdd FILL
XFILL_5__2234_ gnd vdd FILL
XFILL_2__2456_ gnd vdd FILL
XFILL_5__2165_ gnd vdd FILL
XFILL_2__2387_ gnd vdd FILL
XFILL_0__3210_ gnd vdd FILL
XFILL_5__2096_ gnd vdd FILL
XFILL_8__2914_ gnd vdd FILL
XFILL_0__3141_ gnd vdd FILL
XFILL_8__2845_ gnd vdd FILL
XFILL_4_BUFX2_insert7 gnd vdd FILL
XFILL_6__1860_ gnd vdd FILL
XFILL_2__3008_ gnd vdd FILL
XFILL_0__3072_ gnd vdd FILL
X_2720_ _2720_/A _2720_/B _2720_/C _2732_/A vdd gnd NAND3X1
XFILL_8__2776_ gnd vdd FILL
XFILL_0__2023_ gnd vdd FILL
XFILL_5__2998_ gnd vdd FILL
XFILL_6__1791_ gnd vdd FILL
XFILL_8__1727_ gnd vdd FILL
X_2651_ _3575_/Q _2670_/B _2651_/C _2656_/D vdd gnd AOI21X1
XFILL_6__3530_ gnd vdd FILL
XFILL_5__1949_ gnd vdd FILL
X_2582_ _2700_/B _2582_/B _2582_/C _2583_/C vdd gnd OAI21X1
XFILL_6__3461_ gnd vdd FILL
XFILL_3__2703_ gnd vdd FILL
XFILL_0__2925_ gnd vdd FILL
XFILL184650x124950 gnd vdd FILL
XFILL_6__3392_ gnd vdd FILL
XFILL_6__2412_ gnd vdd FILL
XFILL184050x140550 gnd vdd FILL
XFILL_6__2343_ gnd vdd FILL
X_3203_ _3215_/A _3203_/B _3203_/C _3349_/D vdd gnd OAI21X1
XFILL_3__2634_ gnd vdd FILL
XFILL_0__2856_ gnd vdd FILL
XFILL_3__2565_ gnd vdd FILL
X_3134_ _3343_/Q _3143_/B _3135_/C vdd gnd NAND2X1
XFILL_6__2274_ gnd vdd FILL
XFILL_0__2787_ gnd vdd FILL
XFILL_0__1807_ gnd vdd FILL
X_3065_ _3319_/Q _3090_/A _3066_/C vdd gnd NAND2X1
XFILL_3__2496_ gnd vdd FILL
XFILL_0__1738_ gnd vdd FILL
X_2016_ _2033_/A _2950_/A _2016_/C _2161_/B vdd gnd OAI21X1
XFILL_0__3408_ gnd vdd FILL
XFILL_1__2201_ gnd vdd FILL
XFILL_3__3117_ gnd vdd FILL
XFILL_9__2885_ gnd vdd FILL
XFILL_1__3181_ gnd vdd FILL
XFILL_3__3048_ gnd vdd FILL
XFILL_1__2132_ gnd vdd FILL
X_2918_ _2923_/A _2918_/B _2919_/C vdd gnd NOR2X1
XFILL_1__2063_ gnd vdd FILL
X_2849_ _2900_/A _2926_/C _2850_/A vdd gnd NOR2X1
XFILL_4__2812_ gnd vdd FILL
XFILL_6__1989_ gnd vdd FILL
XFILL_7__2521_ gnd vdd FILL
XFILL_4__2743_ gnd vdd FILL
XFILL_1__2965_ gnd vdd FILL
XFILL_7__2452_ gnd vdd FILL
XFILL_1__1916_ gnd vdd FILL
XFILL_7__2383_ gnd vdd FILL
XFILL_4__2674_ gnd vdd FILL
XFILL_1__2896_ gnd vdd FILL
XFILL_1__1847_ gnd vdd FILL
XFILL_1__1778_ gnd vdd FILL
XFILL_1__3517_ gnd vdd FILL
XFILL_2__2310_ gnd vdd FILL
XFILL_7__3004_ gnd vdd FILL
XFILL_4__3226_ gnd vdd FILL
XFILL_1__3448_ gnd vdd FILL
XFILL_2__2241_ gnd vdd FILL
XFILL_4__3157_ gnd vdd FILL
XFILL_1__3379_ gnd vdd FILL
XFILL_2__2172_ gnd vdd FILL
XFILL_4__2108_ gnd vdd FILL
XFILL_4__3088_ gnd vdd FILL
XFILL_5__2921_ gnd vdd FILL
XFILL_4__2039_ gnd vdd FILL
XFILL_8__2630_ gnd vdd FILL
XFILL_5__2852_ gnd vdd FILL
XFILL_5__1803_ gnd vdd FILL
XFILL_8__2561_ gnd vdd FILL
XFILL_5__2783_ gnd vdd FILL
XFILL_8__2492_ gnd vdd FILL
XFILL_7__2719_ gnd vdd FILL
XFILL_5__1734_ gnd vdd FILL
XFILL_2__1956_ gnd vdd FILL
XFILL_8__3113_ gnd vdd FILL
XFILL_5__3404_ gnd vdd FILL
XFILL_2__1887_ gnd vdd FILL
XFILL_0__2710_ gnd vdd FILL
XFILL_2__3557_ gnd vdd FILL
XFILL_8__3044_ gnd vdd FILL
XFILL_3__2350_ gnd vdd FILL
XFILL_0__2641_ gnd vdd FILL
XFILL_0__2572_ gnd vdd FILL
XFILL_2__2508_ gnd vdd FILL
XFILL_2__3488_ gnd vdd FILL
XFILL_5__2217_ gnd vdd FILL
XFILL_3__2281_ gnd vdd FILL
XFILL_5__3197_ gnd vdd FILL
XFILL_5__2148_ gnd vdd FILL
XFILL_2__2439_ gnd vdd FILL
XFILL_5_BUFX2_insert10 gnd vdd FILL
XFILL_5__2079_ gnd vdd FILL
XFILL_5_BUFX2_insert21 gnd vdd FILL
XFILL_6__2961_ gnd vdd FILL
XFILL_5_BUFX2_insert43 gnd vdd FILL
XFILL_0__3124_ gnd vdd FILL
XFILL_6__2892_ gnd vdd FILL
XFILL_5_BUFX2_insert65 gnd vdd FILL
XFILL_6__1912_ gnd vdd FILL
XFILL_5_BUFX2_insert54 gnd vdd FILL
XFILL_5_BUFX2_insert76 gnd vdd FILL
XFILL_8__2828_ gnd vdd FILL
XFILL_6__1843_ gnd vdd FILL
XFILL_5_BUFX2_insert87 gnd vdd FILL
XFILL184650x136650 gnd vdd FILL
XFILL_0__3055_ gnd vdd FILL
X_2703_ _2771_/A _2703_/B _2703_/C _2704_/B vdd gnd NAND3X1
XFILL_8__2759_ gnd vdd FILL
XFILL184350x144450 gnd vdd FILL
XFILL_0__2006_ gnd vdd FILL
XFILL_6__1774_ gnd vdd FILL
X_2634_ _2641_/B _2671_/B _2638_/D _2635_/C vdd gnd OAI21X1
XFILL_6__3513_ gnd vdd FILL
X_2565_ _2565_/A _3296_/D _2565_/C _2566_/C vdd gnd AOI21X1
XFILL_3__1996_ gnd vdd FILL
XFILL_6__3444_ gnd vdd FILL
X_2496_ _3353_/Q _2538_/B _2496_/C _2497_/B vdd gnd AOI21X1
XFILL_1__2750_ gnd vdd FILL
XFILL_0__2908_ gnd vdd FILL
XFILL_6__3375_ gnd vdd FILL
XFILL_1__1701_ gnd vdd FILL
XFILL_1__2681_ gnd vdd FILL
XFILL_3__2617_ gnd vdd FILL
XFILL_0__2839_ gnd vdd FILL
XFILL_6__2326_ gnd vdd FILL
XFILL_4__2390_ gnd vdd FILL
XFILL_3__3597_ gnd vdd FILL
X_3117_ _3125_/A _3125_/B _3334_/Q _3118_/C vdd gnd OAI21X1
XFILL_6__2257_ gnd vdd FILL
XFILL_3__2548_ gnd vdd FILL
XFILL_3__2479_ gnd vdd FILL
XFILL_6__2188_ gnd vdd FILL
XFILL_4__3011_ gnd vdd FILL
X_3048_ _3048_/A _3050_/A vdd gnd INVX1
XFILL_7__1952_ gnd vdd FILL
XFILL_1__3164_ gnd vdd FILL
XFILL_1__2115_ gnd vdd FILL
XFILL_1__3095_ gnd vdd FILL
XFILL_7__1883_ gnd vdd FILL
XFILL_1__2046_ gnd vdd FILL
XFILL_7__3553_ gnd vdd FILL
XFILL_7__3484_ gnd vdd FILL
XFILL_7__2504_ gnd vdd FILL
XFILL_2__1810_ gnd vdd FILL
XFILL_2__2790_ gnd vdd FILL
XFILL_4__2726_ gnd vdd FILL
XFILL_7__2435_ gnd vdd FILL
XFILL_1__2948_ gnd vdd FILL
XFILL_4__2657_ gnd vdd FILL
XFILL_2__1741_ gnd vdd FILL
XFILL_1__2879_ gnd vdd FILL
XFILL_7__2366_ gnd vdd FILL
XFILL_2__3411_ gnd vdd FILL
XFILL_7__2297_ gnd vdd FILL
XFILL_4__2588_ gnd vdd FILL
XFILL_5__3120_ gnd vdd FILL
XFILL_5__3051_ gnd vdd FILL
XFILL_5__2002_ gnd vdd FILL
XFILL_4__3209_ gnd vdd FILL
XFILL_8__1992_ gnd vdd FILL
XFILL_2__2224_ gnd vdd FILL
XFILL_2__2155_ gnd vdd FILL
XFILL_5__2904_ gnd vdd FILL
XFILL_2__2086_ gnd vdd FILL
XFILL_8__3593_ gnd vdd FILL
XFILL_8__2613_ gnd vdd FILL
XFILL_5__2835_ gnd vdd FILL
XFILL_8__2544_ gnd vdd FILL
XFILL_5__2766_ gnd vdd FILL
XFILL_3__1850_ gnd vdd FILL
XFILL_2__2988_ gnd vdd FILL
XFILL_8__2475_ gnd vdd FILL
XFILL_5__1717_ gnd vdd FILL
XFILL_3__1781_ gnd vdd FILL
XFILL_2__1939_ gnd vdd FILL
XFILL_3__3520_ gnd vdd FILL
X_2350_ _2350_/A _2350_/B _2350_/C _2351_/B vdd gnd NAND3X1
XFILL_5__2697_ gnd vdd FILL
XFILL_3__3451_ gnd vdd FILL
X_2281_ _2315_/C _2281_/B _2281_/C _2326_/A vdd gnd NAND3X1
XFILL_3__2402_ gnd vdd FILL
XFILL_6__3160_ gnd vdd FILL
XFILL_6__3091_ gnd vdd FILL
XFILL_3__3382_ gnd vdd FILL
XFILL_8__3027_ gnd vdd FILL
XFILL_6__2111_ gnd vdd FILL
XFILL_0__2624_ gnd vdd FILL
XFILL_6__2042_ gnd vdd FILL
XFILL_3__2333_ gnd vdd FILL
XFILL_3__2264_ gnd vdd FILL
XFILL_0__2555_ gnd vdd FILL
XBUFX2_insert4 RDY _2767_/A vdd gnd BUFX2
XFILL_0__2486_ gnd vdd FILL
XFILL_3__2195_ gnd vdd FILL
XFILL184350x156150 gnd vdd FILL
XFILL184650x148350 gnd vdd FILL
XFILL_6__2944_ gnd vdd FILL
X_1996_ _3256_/Q _2623_/B vdd gnd INVX1
XFILL_0__3107_ gnd vdd FILL
XFILL_6__2875_ gnd vdd FILL
XFILL_0__3038_ gnd vdd FILL
XFILL_4__1890_ gnd vdd FILL
XFILL_6__1826_ gnd vdd FILL
XFILL_6__1757_ gnd vdd FILL
XFILL_3__1979_ gnd vdd FILL
XFILL_4__3560_ gnd vdd FILL
X_3597_ _3597_/A DO[2] vdd gnd BUFX2
X_2617_ _2621_/B _2671_/B _2617_/C _2639_/A vdd gnd OAI21X1
XFILL_1__2802_ gnd vdd FILL
XFILL_4__2511_ gnd vdd FILL
XFILL_6__1688_ gnd vdd FILL
X_2548_ _3063_/C _2570_/B _2548_/C _2549_/C vdd gnd OAI21X1
XFILL_4__3491_ gnd vdd FILL
XFILL_6__3427_ gnd vdd FILL
XFILL_7__2220_ gnd vdd FILL
XFILL_1__2733_ gnd vdd FILL
XFILL_7__2151_ gnd vdd FILL
X_2479_ _2479_/A _2503_/B _2482_/A vdd gnd NAND2X1
XFILL_1_BUFX2_insert52 gnd vdd FILL
XFILL_4__2442_ gnd vdd FILL
XFILL_1_BUFX2_insert41 gnd vdd FILL
XFILL_3_CLKBUF1_insert38 gnd vdd FILL
XFILL_6__2309_ gnd vdd FILL
XFILL_1_BUFX2_insert85 gnd vdd FILL
XFILL_1_BUFX2_insert63 gnd vdd FILL
XFILL_1_BUFX2_insert74 gnd vdd FILL
XFILL_4__2373_ gnd vdd FILL
XFILL_1__2664_ gnd vdd FILL
XFILL_1_BUFX2_insert96 gnd vdd FILL
XFILL_7__2082_ gnd vdd FILL
XFILL_1__2595_ gnd vdd FILL
XFILL_1__3216_ gnd vdd FILL
XFILL_1_CLKBUF1_insert31 gnd vdd FILL
XFILL_7__2984_ gnd vdd FILL
XFILL_7__1935_ gnd vdd FILL
XFILL_1__3147_ gnd vdd FILL
XFILL_7__1866_ gnd vdd FILL
XFILL_1__3078_ gnd vdd FILL
XFILL_2__2911_ gnd vdd FILL
XFILL_1__2029_ gnd vdd FILL
XFILL_5__2620_ gnd vdd FILL
XFILL_7__1797_ gnd vdd FILL
XFILL_2__2842_ gnd vdd FILL
XFILL_7__3536_ gnd vdd FILL
XFILL_5__2551_ gnd vdd FILL
XFILL_7__3467_ gnd vdd FILL
XFILL_8__2260_ gnd vdd FILL
XFILL_2__2773_ gnd vdd FILL
XFILL_7__3398_ gnd vdd FILL
XFILL_8__2191_ gnd vdd FILL
XFILL_7__2418_ gnd vdd FILL
XFILL_5__2482_ gnd vdd FILL
XFILL_4__2709_ gnd vdd FILL
XFILL_2__1724_ gnd vdd FILL
XFILL_7__2349_ gnd vdd FILL
XFILL_5__3103_ gnd vdd FILL
XFILL_5__3034_ gnd vdd FILL
XFILL_0__2340_ gnd vdd FILL
XFILL_0__2271_ gnd vdd FILL
XFILL_8__1975_ gnd vdd FILL
XFILL_2__2207_ gnd vdd FILL
XFILL_2__3187_ gnd vdd FILL
X_1850_ _3189_/B _3151_/C vdd gnd INVX1
XFILL_2__2138_ gnd vdd FILL
X_1781_ _3144_/B _3160_/C _3189_/C vdd gnd NAND2X1
XFILL_3__2951_ gnd vdd FILL
X_3520_ _3523_/B _3523_/A _3520_/C _3522_/A vdd gnd OAI21X1
XFILL_2__2069_ gnd vdd FILL
XFILL_6__2660_ gnd vdd FILL
XFILL_5__2818_ gnd vdd FILL
XFILL_3__2882_ gnd vdd FILL
XFILL_3__1902_ gnd vdd FILL
X_3451_ _3514_/B _3451_/B _3451_/C _3493_/B vdd gnd AOI21X1
XFILL_8__2527_ gnd vdd FILL
XFILL_6__2591_ gnd vdd FILL
XFILL_3__1833_ gnd vdd FILL
X_3382_ _3521_/A _3459_/A vdd gnd INVX2
X_2402_ _2641_/B _2426_/B _2402_/C _2403_/C vdd gnd OAI21X1
XFILL_8__2458_ gnd vdd FILL
XFILL_5__2749_ gnd vdd FILL
XFILL_3__3503_ gnd vdd FILL
X_2333_ _2333_/A _2333_/B _2334_/B vdd gnd OR2X2
XFILL_3__1764_ gnd vdd FILL
XFILL_0__1986_ gnd vdd FILL
XFILL_3__1695_ gnd vdd FILL
XFILL_8__2389_ gnd vdd FILL
XFILL_6__3212_ gnd vdd FILL
XFILL_6__3143_ gnd vdd FILL
X_2264_ _2264_/A _2264_/B _2273_/C vdd gnd NOR2X1
XFILL_3__3434_ gnd vdd FILL
XFILL_8_BUFX2_insert91 gnd vdd FILL
X_2195_ _2933_/C _2871_/C _2896_/B vdd gnd NAND2X1
XFILL_3__3365_ gnd vdd FILL
XFILL_8_BUFX2_insert80 gnd vdd FILL
XFILL_6__3074_ gnd vdd FILL
XFILL_0__3587_ gnd vdd FILL
XFILL_1__2380_ gnd vdd FILL
XFILL_3__2316_ gnd vdd FILL
XFILL_0__2607_ gnd vdd FILL
XFILL_6__2025_ gnd vdd FILL
XFILL_0__2538_ gnd vdd FILL
XFILL_3__2247_ gnd vdd FILL
XFILL_0__2469_ gnd vdd FILL
XFILL_3__2178_ gnd vdd FILL
XFILL_1__3001_ gnd vdd FILL
XFILL_6__2927_ gnd vdd FILL
XFILL_4__2991_ gnd vdd FILL
XFILL_7__1720_ gnd vdd FILL
X_1979_ _1979_/A _1979_/B _1979_/C _2515_/A vdd gnd NAND3X1
XFILL_4__1942_ gnd vdd FILL
XFILL_4__1873_ gnd vdd FILL
XFILL_6__2858_ gnd vdd FILL
XFILL_6__2789_ gnd vdd FILL
XFILL_6__1809_ gnd vdd FILL
XFILL_4__3543_ gnd vdd FILL
XFILL_4__3474_ gnd vdd FILL
XFILL_7__2203_ gnd vdd FILL
XFILL_4__2425_ gnd vdd FILL
XFILL_1__2716_ gnd vdd FILL
XFILL_7__3183_ gnd vdd FILL
XFILL_7__2134_ gnd vdd FILL
XFILL_1__2647_ gnd vdd FILL
XFILL_7__2065_ gnd vdd FILL
XFILL_4__2356_ gnd vdd FILL
XFILL_1__2578_ gnd vdd FILL
XFILL_2__3110_ gnd vdd FILL
XFILL_4__2287_ gnd vdd FILL
XFILL_2__3041_ gnd vdd FILL
XFILL_8__1760_ gnd vdd FILL
XFILL_7__2967_ gnd vdd FILL
XFILL_7__1918_ gnd vdd FILL
XFILL_5__1982_ gnd vdd FILL
XFILL_7__2898_ gnd vdd FILL
XFILL_8__1691_ gnd vdd FILL
XFILL_8__3430_ gnd vdd FILL
XFILL_7__1849_ gnd vdd FILL
XFILL_2__2825_ gnd vdd FILL
XFILL_7__3519_ gnd vdd FILL
XFILL_8__2312_ gnd vdd FILL
XFILL_5__3583_ gnd vdd FILL
XFILL_5__2603_ gnd vdd FILL
XFILL_8__2243_ gnd vdd FILL
XFILL_5__2534_ gnd vdd FILL
XFILL_0__1840_ gnd vdd FILL
XFILL_5__2465_ gnd vdd FILL
XFILL_2__2756_ gnd vdd FILL
XFILL_0__1771_ gnd vdd FILL
XFILL_2__1707_ gnd vdd FILL
XFILL_8__2174_ gnd vdd FILL
XFILL_2__2687_ gnd vdd FILL
XFILL_0__3510_ gnd vdd FILL
XFILL_5__2396_ gnd vdd FILL
XFILL_0__3441_ gnd vdd FILL
XFILL_3__3150_ gnd vdd FILL
XFILL_3__3081_ gnd vdd FILL
XFILL_5__3017_ gnd vdd FILL
XFILL_0__3372_ gnd vdd FILL
XFILL_3__2101_ gnd vdd FILL
X_2951_ reset _2957_/C _3304_/Q _2952_/C vdd gnd OAI21X1
XFILL_3__2032_ gnd vdd FILL
XFILL_0__2323_ gnd vdd FILL
XFILL_0__2254_ gnd vdd FILL
XCLKBUF1_insert33 clk _3313_/CLK vdd gnd CLKBUF1
X_1902_ _1902_/A _1902_/B _1902_/C _1903_/B vdd gnd NAND3X1
XFILL_8__1958_ gnd vdd FILL
X_2882_ _2885_/B _2882_/B _2882_/C _3280_/D vdd gnd OAI21X1
XFILL_0__2185_ gnd vdd FILL
XFILL_8__1889_ gnd vdd FILL
XFILL_6__2712_ gnd vdd FILL
X_1833_ _2058_/B _2048_/B _3176_/A vdd gnd NAND2X1
XFILL_3__2934_ gnd vdd FILL
X_1764_ _3237_/Q _3165_/A vdd gnd INVX4
XFILL_8__3559_ gnd vdd FILL
X_3503_ _3508_/B _3508_/A _3529_/C vdd gnd NAND2X1
XFILL_6__2643_ gnd vdd FILL
XFILL_3__2865_ gnd vdd FILL
X_3434_ _3434_/A _3521_/A _3441_/C vdd gnd NAND2X1
X_1695_ _3566_/A _3292_/Q _1696_/C vdd gnd OR2X2
XFILL_6__2574_ gnd vdd FILL
XFILL_1__1880_ gnd vdd FILL
XFILL_3__2796_ gnd vdd FILL
XFILL_3__1816_ gnd vdd FILL
X_3365_ _3575_/Q _3574_/Q _3368_/A vdd gnd NOR2X1
XFILL_3__1747_ gnd vdd FILL
XFILL_1__3550_ gnd vdd FILL
XFILL_0__1969_ gnd vdd FILL
X_3296_ _3296_/D vdd _3355_/R _3578_/CLK _3296_/Q vdd gnd DFFSR
X_2316_ _2345_/A _2327_/B _2317_/A vdd gnd NAND2X1
XFILL_1__3481_ gnd vdd FILL
XFILL_3__3417_ gnd vdd FILL
XFILL_4__2210_ gnd vdd FILL
XFILL_1__2501_ gnd vdd FILL
X_2247_ _2894_/A _2247_/B _2306_/A vdd gnd NAND2X1
XFILL_6__3126_ gnd vdd FILL
XFILL_1__2432_ gnd vdd FILL
XFILL_4__3190_ gnd vdd FILL
XFILL_6__3057_ gnd vdd FILL
XFILL_4__2141_ gnd vdd FILL
X_2178_ _2293_/A _3160_/B _3151_/A _2184_/B vdd gnd NAND3X1
XFILL_4__2072_ gnd vdd FILL
XFILL_1__2363_ gnd vdd FILL
XFILL_6__2008_ gnd vdd FILL
XFILL_1__2294_ gnd vdd FILL
XFILL_7__2821_ gnd vdd FILL
XFILL_7__2752_ gnd vdd FILL
XFILL_4__2974_ gnd vdd FILL
XFILL_7__1703_ gnd vdd FILL
XFILL_7__2683_ gnd vdd FILL
XFILL_4__1925_ gnd vdd FILL
XFILL_4__1856_ gnd vdd FILL
XFILL_4__1787_ gnd vdd FILL
XFILL_4__3526_ gnd vdd FILL
XFILL_2__3590_ gnd vdd FILL
XFILL_2__2610_ gnd vdd FILL
XFILL_2__2541_ gnd vdd FILL
XFILL_5__2250_ gnd vdd FILL
XFILL_4__3457_ gnd vdd FILL
XFILL_7__3166_ gnd vdd FILL
XFILL_4__3388_ gnd vdd FILL
XFILL_5__2181_ gnd vdd FILL
XFILL_7__2117_ gnd vdd FILL
XFILL_2__2472_ gnd vdd FILL
XFILL_4__2408_ gnd vdd FILL
XFILL_7__3097_ gnd vdd FILL
XFILL_4__2339_ gnd vdd FILL
XFILL_8__2930_ gnd vdd FILL
XFILL_7__2048_ gnd vdd FILL
XFILL_8__2861_ gnd vdd FILL
XFILL_2__3024_ gnd vdd FILL
XFILL_8__1812_ gnd vdd FILL
XFILL_8__2792_ gnd vdd FILL
XFILL_8__1743_ gnd vdd FILL
XFILL_5__1965_ gnd vdd FILL
XFILL_8__3413_ gnd vdd FILL
XFILL_5__1896_ gnd vdd FILL
XFILL_2_BUFX2_insert18 gnd vdd FILL
XFILL_0__2941_ gnd vdd FILL
XFILL_3__2650_ gnd vdd FILL
XFILL_2__2808_ gnd vdd FILL
XFILL_5__3566_ gnd vdd FILL
XFILL_0__2872_ gnd vdd FILL
XFILL_3__2581_ gnd vdd FILL
XFILL_5__3497_ gnd vdd FILL
XFILL_8__2226_ gnd vdd FILL
XFILL_0__1823_ gnd vdd FILL
XFILL_6__2290_ gnd vdd FILL
XFILL_5__2517_ gnd vdd FILL
X_3150_ _3150_/A _3179_/A _3179_/C _3154_/B vdd gnd NAND3X1
XFILL_2__2739_ gnd vdd FILL
X_3081_ _3321_/Q _3090_/A _3082_/C vdd gnd NAND2X1
X_2101_ _2294_/A _2437_/C _2101_/C _2349_/B vdd gnd OAI21X1
XFILL_0__1754_ gnd vdd FILL
XFILL_5__2448_ gnd vdd FILL
X_2032_ _2889_/C _2161_/B _2932_/B vdd gnd NAND2X1
XFILL_8__2157_ gnd vdd FILL
XFILL_5__2379_ gnd vdd FILL
XFILL_8__2088_ gnd vdd FILL
XFILL_3__3202_ gnd vdd FILL
XFILL_3__3133_ gnd vdd FILL
XFILL_0__3424_ gnd vdd FILL
XFILL_0__2306_ gnd vdd FILL
XFILL_3__3064_ gnd vdd FILL
X_2934_ _2934_/A _2934_/B _2934_/C _2935_/B vdd gnd NAND3X1
XFILL_3__2015_ gnd vdd FILL
X_2865_ _2865_/A _2887_/A _2865_/C _2865_/D _3274_/D vdd gnd OAI22X1
XFILL_0__2237_ gnd vdd FILL
XFILL_0__2168_ gnd vdd FILL
X_1816_ _2612_/B _3189_/C _3016_/A _1831_/D _3484_/B vdd gnd OAI22X1
X_2796_ _2906_/A _2906_/B _3262_/Q _2799_/C vdd gnd OAI21X1
XFILL_3__2917_ gnd vdd FILL
XFILL_9__3384_ gnd vdd FILL
XFILL_1__2981_ gnd vdd FILL
XFILL_4__1710_ gnd vdd FILL
X_1747_ _2594_/B _2442_/A _3160_/C vdd gnd NOR2X1
XFILL_4__2690_ gnd vdd FILL
XFILL_6__2626_ gnd vdd FILL
XFILL_0__2099_ gnd vdd FILL
XFILL_3__2848_ gnd vdd FILL
XFILL_8_CLKBUF1_insert38 gnd vdd FILL
XFILL_1__1932_ gnd vdd FILL
X_3417_ _3421_/B _3417_/B _3459_/A _3418_/A vdd gnd OAI21X1
XFILL_1__1863_ gnd vdd FILL
XFILL_6__2557_ gnd vdd FILL
XFILL_1__3602_ gnd vdd FILL
XFILL_6__2488_ gnd vdd FILL
X_3348_ _3348_/D vdd _3362_/R _3363_/CLK _3348_/Q vdd gnd DFFSR
XFILL_3__2779_ gnd vdd FILL
XFILL_1__3533_ gnd vdd FILL
XFILL_7__3020_ gnd vdd FILL
XFILL_1__1794_ gnd vdd FILL
XFILL_1_BUFX2_insert4 gnd vdd FILL
X_3279_ _3279_/D vdd _3313_/R _3313_/CLK _3279_/Q vdd gnd DFFSR
XFILL_6_CLKBUF1_insert31 gnd vdd FILL
XFILL_1__3464_ gnd vdd FILL
XFILL_4__3173_ gnd vdd FILL
XFILL_6__3109_ gnd vdd FILL
XFILL_1__3395_ gnd vdd FILL
XFILL_1__2415_ gnd vdd FILL
XFILL_4__2124_ gnd vdd FILL
XFILL_1__2346_ gnd vdd FILL
XFILL_4__2055_ gnd vdd FILL
XFILL_1__2277_ gnd vdd FILL
XFILL_7__2804_ gnd vdd FILL
XFILL_7__2735_ gnd vdd FILL
XFILL_4__2957_ gnd vdd FILL
XFILL_5__1750_ gnd vdd FILL
XFILL_2__1972_ gnd vdd FILL
XFILL_7__2666_ gnd vdd FILL
XFILL_4__1908_ gnd vdd FILL
XFILL_5__3420_ gnd vdd FILL
XFILL_4__2888_ gnd vdd FILL
XFILL_9_BUFX2_insert24 gnd vdd FILL
XFILL_7__2597_ gnd vdd FILL
XFILL_4__1839_ gnd vdd FILL
XFILL_9_BUFX2_insert68 gnd vdd FILL
XFILL_8__3060_ gnd vdd FILL
XFILL_8__2011_ gnd vdd FILL
XFILL_4__3509_ gnd vdd FILL
XFILL_5__2302_ gnd vdd FILL
XFILL_7__3218_ gnd vdd FILL
XFILL_2__2524_ gnd vdd FILL
XFILL_5__2233_ gnd vdd FILL
XFILL_2__2455_ gnd vdd FILL
XFILL_7__3149_ gnd vdd FILL
XFILL_5__2164_ gnd vdd FILL
XFILL_8__2913_ gnd vdd FILL
XFILL_2__2386_ gnd vdd FILL
XFILL_5__2095_ gnd vdd FILL
XFILL_0__3140_ gnd vdd FILL
XFILL_8__2844_ gnd vdd FILL
XFILL_4_BUFX2_insert8 gnd vdd FILL
XFILL_2__3007_ gnd vdd FILL
XFILL_0__3071_ gnd vdd FILL
XFILL_8__2775_ gnd vdd FILL
XFILL_0__2022_ gnd vdd FILL
XFILL_5__2997_ gnd vdd FILL
XFILL_8__1726_ gnd vdd FILL
XFILL_6__1790_ gnd vdd FILL
X_2650_ _2650_/A _2748_/B _2669_/C _2651_/C vdd gnd OAI21X1
XFILL_5__1948_ gnd vdd FILL
X_2581_ _3160_/C _3146_/A _2701_/B _2582_/C vdd gnd OAI21X1
XFILL_5__1879_ gnd vdd FILL
XFILL_6__3460_ gnd vdd FILL
XFILL_3__2702_ gnd vdd FILL
XFILL_0__2924_ gnd vdd FILL
XFILL_6__3391_ gnd vdd FILL
XFILL_3__2633_ gnd vdd FILL
XFILL_6__2411_ gnd vdd FILL
XFILL_5__3549_ gnd vdd FILL
XFILL_0__2855_ gnd vdd FILL
XFILL_6__2342_ gnd vdd FILL
X_3202_ _3214_/A _3214_/B _3349_/Q _3203_/C vdd gnd OAI21X1
XFILL_6__2273_ gnd vdd FILL
XFILL_3__2564_ gnd vdd FILL
XFILL_0__1806_ gnd vdd FILL
X_3133_ _3133_/A _3143_/B _3133_/C _3342_/D vdd gnd OAI21X1
XFILL_0__2786_ gnd vdd FILL
XFILL_8__2209_ gnd vdd FILL
XFILL_3__2495_ gnd vdd FILL
XFILL_8__3189_ gnd vdd FILL
X_3064_ _3294_/D _3088_/S _3064_/C _3137_/A vdd gnd OAI21X1
XFILL_0__1737_ gnd vdd FILL
X_2015_ _2025_/A _3303_/Q _2016_/C vdd gnd NAND2X1
XFILL_0__3407_ gnd vdd FILL
XFILL_1__2200_ gnd vdd FILL
XFILL_3__3116_ gnd vdd FILL
XFILL_1__3180_ gnd vdd FILL
XFILL_3__3047_ gnd vdd FILL
XFILL_1__2131_ gnd vdd FILL
X_2917_ _2928_/B _2917_/B _2917_/C _2918_/B vdd gnd OAI21X1
XFILL_1__2062_ gnd vdd FILL
XFILL_9__1766_ gnd vdd FILL
X_2848_ _2932_/B _2881_/A _2926_/C vdd gnd NAND2X1
XFILL_4__2811_ gnd vdd FILL
XFILL_6__1988_ gnd vdd FILL
XFILL_7__2520_ gnd vdd FILL
X_2779_ _3255_/Q _2780_/B vdd gnd INVX1
XFILL_4__2742_ gnd vdd FILL
XFILL_1__2964_ gnd vdd FILL
XFILL_7__2451_ gnd vdd FILL
XFILL_7__2382_ gnd vdd FILL
XFILL_1__1915_ gnd vdd FILL
XFILL_6__3589_ gnd vdd FILL
XFILL_6__2609_ gnd vdd FILL
XFILL_4__2673_ gnd vdd FILL
XFILL_1__2895_ gnd vdd FILL
XFILL_1__1846_ gnd vdd FILL
XFILL_1__1777_ gnd vdd FILL
XFILL_1__3516_ gnd vdd FILL
XFILL_7__3003_ gnd vdd FILL
XFILL_1__3447_ gnd vdd FILL
XFILL_2__2240_ gnd vdd FILL
XFILL_4__3225_ gnd vdd FILL
XFILL_4__3156_ gnd vdd FILL
XFILL_1__3378_ gnd vdd FILL
XFILL_2__2171_ gnd vdd FILL
XFILL_4__3087_ gnd vdd FILL
XFILL_4__2107_ gnd vdd FILL
XFILL_4__2038_ gnd vdd FILL
XFILL184650x85950 gnd vdd FILL
XFILL_1__2329_ gnd vdd FILL
XFILL_5__2920_ gnd vdd FILL
XFILL_5__2851_ gnd vdd FILL
XFILL_8__2560_ gnd vdd FILL
XFILL_5__1802_ gnd vdd FILL
XFILL_8__2491_ gnd vdd FILL
XFILL_7__2718_ gnd vdd FILL
XFILL_5__2782_ gnd vdd FILL
XFILL_2__1955_ gnd vdd FILL
XFILL_5__1733_ gnd vdd FILL
XFILL_7__2649_ gnd vdd FILL
XFILL_8__3112_ gnd vdd FILL
XFILL_5__3403_ gnd vdd FILL
XFILL_2__1886_ gnd vdd FILL
XFILL_8__3043_ gnd vdd FILL
XFILL_2__3556_ gnd vdd FILL
XFILL_0__2640_ gnd vdd FILL
XFILL_2__2507_ gnd vdd FILL
XFILL_0__2571_ gnd vdd FILL
XFILL_2__3487_ gnd vdd FILL
XFILL_5__2216_ gnd vdd FILL
XFILL_3__2280_ gnd vdd FILL
XFILL_5__3196_ gnd vdd FILL
XFILL_5__2147_ gnd vdd FILL
XFILL_2__2438_ gnd vdd FILL
XFILL_2__2369_ gnd vdd FILL
XFILL_5__2078_ gnd vdd FILL
XFILL_6__2960_ gnd vdd FILL
XFILL_5_BUFX2_insert22 gnd vdd FILL
XFILL_5_BUFX2_insert11 gnd vdd FILL
XFILL_5_BUFX2_insert44 gnd vdd FILL
XFILL_0__3123_ gnd vdd FILL
XFILL_6__2891_ gnd vdd FILL
XFILL_8__2827_ gnd vdd FILL
XFILL_5_BUFX2_insert66 gnd vdd FILL
XFILL_6__1911_ gnd vdd FILL
XFILL_5_BUFX2_insert55 gnd vdd FILL
XFILL_5_BUFX2_insert77 gnd vdd FILL
XFILL_0__3054_ gnd vdd FILL
XFILL_6__1842_ gnd vdd FILL
XFILL_5_BUFX2_insert88 gnd vdd FILL
X_2702_ _3357_/Q _2702_/B _2993_/B _2703_/C vdd gnd NAND3X1
XFILL_0__2005_ gnd vdd FILL
XFILL_8__2758_ gnd vdd FILL
XFILL_8__1709_ gnd vdd FILL
XFILL_8__2689_ gnd vdd FILL
XFILL_6__1773_ gnd vdd FILL
X_2633_ _3573_/Q _2670_/B _2633_/C _2638_/D vdd gnd AOI21X1
XFILL_6__3512_ gnd vdd FILL
XFILL_3__1995_ gnd vdd FILL
X_2564_ _3230_/A _2572_/B _2564_/C _2565_/C vdd gnd OAI21X1
XFILL_6__3443_ gnd vdd FILL
XFILL_1__1700_ gnd vdd FILL
X_2495_ _2952_/A _2510_/B _2650_/A _2570_/B _2496_/C vdd gnd OAI22X1
XFILL_0__2907_ gnd vdd FILL
XFILL_6__3374_ gnd vdd FILL
XFILL_1__2680_ gnd vdd FILL
XFILL_3__2616_ gnd vdd FILL
XFILL_0__2838_ gnd vdd FILL
XFILL_6__2325_ gnd vdd FILL
XFILL_3__3596_ gnd vdd FILL
X_3116_ _3133_/A _3126_/B _3116_/C _3333_/D vdd gnd OAI21X1
XFILL_6__2256_ gnd vdd FILL
XFILL_0__2769_ gnd vdd FILL
XFILL_3__2547_ gnd vdd FILL
XFILL_6__2187_ gnd vdd FILL
XFILL_3__2478_ gnd vdd FILL
XFILL_4__3010_ gnd vdd FILL
X_3047_ _3056_/B _3572_/Q _3048_/A vdd gnd XNOR2X1
XFILL_1__3232_ gnd vdd FILL
XFILL_7__1951_ gnd vdd FILL
XFILL_1__3163_ gnd vdd FILL
XFILL_1__2114_ gnd vdd FILL
XFILL_1__3094_ gnd vdd FILL
XFILL_7__1882_ gnd vdd FILL
XFILL_1__2045_ gnd vdd FILL
XFILL184350x15750 gnd vdd FILL
XFILL_7__3552_ gnd vdd FILL
XFILL_7__3483_ gnd vdd FILL
XFILL_7__2503_ gnd vdd FILL
XFILL_4__2725_ gnd vdd FILL
XFILL_7__2434_ gnd vdd FILL
XFILL_1__2947_ gnd vdd FILL
XFILL_2__1740_ gnd vdd FILL
XFILL_4__2656_ gnd vdd FILL
XFILL_1__2878_ gnd vdd FILL
XFILL_7__2365_ gnd vdd FILL
XFILL_2__3410_ gnd vdd FILL
XFILL_7__2296_ gnd vdd FILL
XFILL_1__1829_ gnd vdd FILL
XFILL_4__2587_ gnd vdd FILL
XFILL_5__3050_ gnd vdd FILL
XFILL184650x97650 gnd vdd FILL
XFILL_5__2001_ gnd vdd FILL
XFILL_4__3208_ gnd vdd FILL
XFILL_8__1991_ gnd vdd FILL
XFILL_2__2223_ gnd vdd FILL
XFILL_4__3139_ gnd vdd FILL
XFILL_2__2154_ gnd vdd FILL
XFILL_5__2903_ gnd vdd FILL
XFILL_2__2085_ gnd vdd FILL
XFILL_8__3592_ gnd vdd FILL
XFILL_8__2612_ gnd vdd FILL
XFILL_5__2834_ gnd vdd FILL
XFILL_8__2543_ gnd vdd FILL
XFILL_5__2765_ gnd vdd FILL
XFILL181950x140550 gnd vdd FILL
XFILL_2__2987_ gnd vdd FILL
XFILL_3__1780_ gnd vdd FILL
XFILL_8__2474_ gnd vdd FILL
XFILL_5__1716_ gnd vdd FILL
XFILL_2__1938_ gnd vdd FILL
XFILL_5__2696_ gnd vdd FILL
XFILL_3__3450_ gnd vdd FILL
X_2280_ _2352_/B _2280_/B _2281_/B vdd gnd AND2X2
XFILL_2__1869_ gnd vdd FILL
XFILL_3__2401_ gnd vdd FILL
XFILL_6__3090_ gnd vdd FILL
XFILL_3__3381_ gnd vdd FILL
XFILL_8__3026_ gnd vdd FILL
XFILL_0__2623_ gnd vdd FILL
XFILL_6__2110_ gnd vdd FILL
XFILL_6__2041_ gnd vdd FILL
XFILL_2__3539_ gnd vdd FILL
XFILL_3__2332_ gnd vdd FILL
XFILL_3__2263_ gnd vdd FILL
XBUFX2_insert5 RDY _2294_/A vdd gnd BUFX2
XFILL_0__2554_ gnd vdd FILL
XFILL_0__2485_ gnd vdd FILL
XFILL_5__3179_ gnd vdd FILL
XFILL_3__2194_ gnd vdd FILL
XFILL_6__2943_ gnd vdd FILL
XFILL_0__3106_ gnd vdd FILL
X_1995_ IRQ _2008_/A vdd gnd INVX1
XFILL_6__2874_ gnd vdd FILL
XFILL_0__3037_ gnd vdd FILL
XFILL_6__1825_ gnd vdd FILL
XFILL_6__1756_ gnd vdd FILL
X_2616_ _3571_/Q _2670_/B _2616_/C _2617_/C vdd gnd AOI21X1
XFILL_3__1978_ gnd vdd FILL
X_3596_ _3596_/A DO[1] vdd gnd BUFX2
XFILL_1__2801_ gnd vdd FILL
XFILL_4__2510_ gnd vdd FILL
X_2547_ _2569_/A _2569_/B _3294_/D _2548_/C vdd gnd OAI21X1
XFILL_9__3135_ gnd vdd FILL
XFILL_4__3490_ gnd vdd FILL
XFILL_6__3426_ gnd vdd FILL
X_2478_ _2691_/A _2565_/A _2503_/B vdd gnd NOR2X1
XFILL_1__2732_ gnd vdd FILL
XFILL_1_BUFX2_insert20 gnd vdd FILL
XFILL_7__2150_ gnd vdd FILL
XFILL_1_BUFX2_insert42 gnd vdd FILL
XFILL_4__2441_ gnd vdd FILL
XFILL_1__2663_ gnd vdd FILL
XFILL_3_CLKBUF1_insert28 gnd vdd FILL
XFILL_4__2372_ gnd vdd FILL
XFILL_7__2081_ gnd vdd FILL
XFILL_1_BUFX2_insert64 gnd vdd FILL
XFILL_6__2308_ gnd vdd FILL
XFILL_3__3579_ gnd vdd FILL
XFILL_1_BUFX2_insert75 gnd vdd FILL
XFILL_1_BUFX2_insert53 gnd vdd FILL
XFILL_1_BUFX2_insert86 gnd vdd FILL
XFILL_1_BUFX2_insert97 gnd vdd FILL
XFILL_1__2594_ gnd vdd FILL
XFILL_6__2239_ gnd vdd FILL
XFILL_1_CLKBUF1_insert32 gnd vdd FILL
XFILL_1__3215_ gnd vdd FILL
XFILL184350x27450 gnd vdd FILL
XFILL_7__2983_ gnd vdd FILL
XFILL181350x35250 gnd vdd FILL
XFILL_7__1934_ gnd vdd FILL
XFILL_1__3146_ gnd vdd FILL
XFILL_7__1865_ gnd vdd FILL
XFILL_1__3077_ gnd vdd FILL
XFILL_2__2910_ gnd vdd FILL
XFILL_1__2028_ gnd vdd FILL
XFILL_7__3535_ gnd vdd FILL
XFILL_7__1796_ gnd vdd FILL
XFILL_2__2841_ gnd vdd FILL
XFILL_5__2550_ gnd vdd FILL
XFILL_7__3466_ gnd vdd FILL
XFILL_4__2708_ gnd vdd FILL
XFILL_2__2772_ gnd vdd FILL
XFILL_7__3397_ gnd vdd FILL
XFILL_8__2190_ gnd vdd FILL
XFILL_7__2417_ gnd vdd FILL
XFILL_5__2481_ gnd vdd FILL
XFILL_2__1723_ gnd vdd FILL
XFILL_7__2348_ gnd vdd FILL
XFILL_4__2639_ gnd vdd FILL
XFILL_5__3102_ gnd vdd FILL
XFILL_7__2279_ gnd vdd FILL
XFILL_5__3033_ gnd vdd FILL
XFILL_0__2270_ gnd vdd FILL
XFILL_2__2206_ gnd vdd FILL
XFILL_8__1974_ gnd vdd FILL
XFILL_2__3186_ gnd vdd FILL
XFILL_2__2137_ gnd vdd FILL
X_1780_ _3290_/D _3016_/A vdd gnd INVX1
XFILL_2__2068_ gnd vdd FILL
XFILL_3__2950_ gnd vdd FILL
XFILL_5__2817_ gnd vdd FILL
XFILL_3__2881_ gnd vdd FILL
XFILL_3__1901_ gnd vdd FILL
X_3450_ _3514_/B _3451_/B _3514_/A _3451_/C vdd gnd OAI21X1
XFILL_3__1832_ gnd vdd FILL
XFILL_6__2590_ gnd vdd FILL
XFILL_8__2526_ gnd vdd FILL
X_3381_ _3445_/A _3387_/B _3381_/C _3455_/C _3384_/B vdd gnd AOI22X1
X_2401_ _3309_/Q _2425_/B _2402_/C vdd gnd NAND2X1
XFILL_8__2457_ gnd vdd FILL
XFILL_5__2748_ gnd vdd FILL
XFILL_3__3502_ gnd vdd FILL
XFILL_0__1985_ gnd vdd FILL
X_2332_ _2332_/A _2332_/B _2332_/C _2333_/A vdd gnd NAND3X1
XFILL_3__1763_ gnd vdd FILL
XFILL_5__2679_ gnd vdd FILL
XFILL_8__2388_ gnd vdd FILL
XFILL_3__1694_ gnd vdd FILL
XFILL_6__3211_ gnd vdd FILL
XFILL_6__3142_ gnd vdd FILL
XFILL_3__3433_ gnd vdd FILL
X_2263_ _2896_/B _2307_/A _2263_/C _2264_/B vdd gnd NAND3X1
XFILL_8_BUFX2_insert92 gnd vdd FILL
X_2194_ _2910_/A _2871_/C vdd gnd INVX1
XFILL_3__3364_ gnd vdd FILL
XFILL_8_BUFX2_insert81 gnd vdd FILL
XFILL_8_BUFX2_insert70 gnd vdd FILL
XFILL_8__3009_ gnd vdd FILL
XFILL_3__2315_ gnd vdd FILL
XFILL_6__3073_ gnd vdd FILL
XFILL_0__3586_ gnd vdd FILL
XFILL_0__2606_ gnd vdd FILL
XFILL_6__2024_ gnd vdd FILL
XFILL_0__2537_ gnd vdd FILL
XFILL_3__2246_ gnd vdd FILL
XFILL_1__3000_ gnd vdd FILL
XFILL_3__2177_ gnd vdd FILL
XFILL_0__2468_ gnd vdd FILL
XFILL_0__2399_ gnd vdd FILL
XFILL_6__2926_ gnd vdd FILL
XFILL_4__2990_ gnd vdd FILL
XFILL_9__2635_ gnd vdd FILL
X_1978_ _3322_/Q _3029_/B _1979_/B vdd gnd NAND2X1
XFILL_4__1941_ gnd vdd FILL
XFILL_6__2857_ gnd vdd FILL
XFILL_4__1872_ gnd vdd FILL
XFILL_6__1808_ gnd vdd FILL
XFILL_6__2788_ gnd vdd FILL
XFILL_6__1739_ gnd vdd FILL
X_3579_ _3579_/A AB[0] vdd gnd BUFX2
XFILL_4__3542_ gnd vdd FILL
XFILL_4__3473_ gnd vdd FILL
XFILL_6__3409_ gnd vdd FILL
XFILL_7__2202_ gnd vdd FILL
XFILL_4__2424_ gnd vdd FILL
XFILL_1__2715_ gnd vdd FILL
XFILL_7__3182_ gnd vdd FILL
XFILL_7__2133_ gnd vdd FILL
XFILL_1__2646_ gnd vdd FILL
XFILL_1__2577_ gnd vdd FILL
XFILL_7__2064_ gnd vdd FILL
XFILL_4__2355_ gnd vdd FILL
XFILL184350x39150 gnd vdd FILL
XFILL_4__2286_ gnd vdd FILL
XFILL_2__3040_ gnd vdd FILL
XFILL_7__2966_ gnd vdd FILL
XFILL_1__3129_ gnd vdd FILL
XFILL_7__1917_ gnd vdd FILL
XFILL_5__1981_ gnd vdd FILL
XFILL_7__2897_ gnd vdd FILL
XFILL_8__1690_ gnd vdd FILL
XFILL_7__1848_ gnd vdd FILL
XFILL_5__2602_ gnd vdd FILL
XFILL_7__1779_ gnd vdd FILL
XFILL_2__2824_ gnd vdd FILL
XFILL_7__3518_ gnd vdd FILL
XFILL_8__2311_ gnd vdd FILL
XFILL_5__3582_ gnd vdd FILL
XFILL_7__3449_ gnd vdd FILL
XFILL_8__2242_ gnd vdd FILL
XFILL_5__2533_ gnd vdd FILL
XFILL_5__2464_ gnd vdd FILL
XFILL_2__2755_ gnd vdd FILL
XFILL_0__1770_ gnd vdd FILL
XFILL_8__2173_ gnd vdd FILL
XFILL_2__1706_ gnd vdd FILL
XFILL_2__2686_ gnd vdd FILL
XFILL_5__2395_ gnd vdd FILL
XFILL_0__3440_ gnd vdd FILL
XFILL_0__3371_ gnd vdd FILL
XFILL_3__2100_ gnd vdd FILL
XFILL_3__3080_ gnd vdd FILL
XFILL_5__3016_ gnd vdd FILL
XFILL_0__2322_ gnd vdd FILL
X_2950_ _2950_/A _2956_/B _2950_/C _3303_/D vdd gnd OAI21X1
XFILL_3__2031_ gnd vdd FILL
XCLKBUF1_insert34 clk _3576_/CLK vdd gnd CLKBUF1
XFILL_8__1957_ gnd vdd FILL
X_2881_ _2881_/A _2909_/C _2881_/C _2933_/A _2882_/B vdd gnd AOI22X1
XFILL_0__2253_ gnd vdd FILL
X_1901_ _2938_/A _3157_/C _1902_/B vdd gnd NOR2X1
XFILL_0__2184_ gnd vdd FILL
X_1832_ _2589_/A _1987_/A _2602_/B _3187_/A vdd gnd OAI21X1
XFILL_2__3169_ gnd vdd FILL
XFILL183450x140550 gnd vdd FILL
XFILL_8__1888_ gnd vdd FILL
XFILL_6__2711_ gnd vdd FILL
XFILL_3__2933_ gnd vdd FILL
X_1763_ _1858_/B _1794_/A _3173_/B vdd gnd NAND2X1
X_3502_ _3502_/A _3552_/B _3502_/C _3554_/B vdd gnd OAI21X1
XFILL_8__3558_ gnd vdd FILL
X_1694_ _3022_/A _1694_/Y vdd gnd INVX8
XFILL_6__2642_ gnd vdd FILL
X_3433_ _3525_/B _3483_/B vdd gnd INVX1
XFILL_3__2864_ gnd vdd FILL
XFILL_8__2509_ gnd vdd FILL
XFILL_6__2573_ gnd vdd FILL
XFILL_8__3489_ gnd vdd FILL
XFILL_3__2795_ gnd vdd FILL
XFILL_3__1815_ gnd vdd FILL
X_3364_ _3570_/Q _3573_/Q _3369_/A vdd gnd OR2X2
XFILL_3__1746_ gnd vdd FILL
XFILL_0__1968_ gnd vdd FILL
X_2315_ _2315_/A _2315_/B _2315_/C _2325_/A vdd gnd OAI21X1
X_3295_ _3295_/D vdd _3355_/R _3355_/CLK _3295_/Q vdd gnd DFFSR
XFILL_1__3480_ gnd vdd FILL
XFILL_3__3416_ gnd vdd FILL
XFILL_0__1899_ gnd vdd FILL
XFILL_1__2500_ gnd vdd FILL
X_2246_ _2246_/A _2246_/B _2246_/C _2315_/C vdd gnd AOI21X1
XFILL_6__3125_ gnd vdd FILL
XFILL_1__2431_ gnd vdd FILL
XFILL_6__3056_ gnd vdd FILL
X_2177_ _2177_/A _2246_/A _2184_/A vdd gnd NAND2X1
XFILL_4__2140_ gnd vdd FILL
XFILL_1__2362_ gnd vdd FILL
XFILL_4__2071_ gnd vdd FILL
XFILL_6__2007_ gnd vdd FILL
XFILL_3__2229_ gnd vdd FILL
XFILL_1__2293_ gnd vdd FILL
XFILL_7__2820_ gnd vdd FILL
XFILL_7__2751_ gnd vdd FILL
XFILL_6__2909_ gnd vdd FILL
XFILL_4__2973_ gnd vdd FILL
XFILL_7__1702_ gnd vdd FILL
XFILL_7__2682_ gnd vdd FILL
XFILL_4__1924_ gnd vdd FILL
XFILL_4_BUFX2_insert90 gnd vdd FILL
XFILL_4__1855_ gnd vdd FILL
XFILL_4__1786_ gnd vdd FILL
XFILL_4__3525_ gnd vdd FILL
XFILL_2__2540_ gnd vdd FILL
XFILL_4__3456_ gnd vdd FILL
XFILL_2__2471_ gnd vdd FILL
XFILL_7__3165_ gnd vdd FILL
XFILL_5__2180_ gnd vdd FILL
XFILL_4__3387_ gnd vdd FILL
XFILL_7__2116_ gnd vdd FILL
XFILL_4__2407_ gnd vdd FILL
XFILL_7__3096_ gnd vdd FILL
XFILL_4__2338_ gnd vdd FILL
XFILL_1__2629_ gnd vdd FILL
XFILL_7__2047_ gnd vdd FILL
XFILL_8__2860_ gnd vdd FILL
XFILL_4__2269_ gnd vdd FILL
XFILL_2__3023_ gnd vdd FILL
XFILL_8__1811_ gnd vdd FILL
XFILL_8__2791_ gnd vdd FILL
XFILL_7__2949_ gnd vdd FILL
XFILL_8__1742_ gnd vdd FILL
XFILL_5__1964_ gnd vdd FILL
XFILL_8__3412_ gnd vdd FILL
XFILL_5__1895_ gnd vdd FILL
XFILL_0__2940_ gnd vdd FILL
XFILL_5__3565_ gnd vdd FILL
XFILL_2_BUFX2_insert19 gnd vdd FILL
XFILL_3__2580_ gnd vdd FILL
XFILL_2__2807_ gnd vdd FILL
XFILL_0__2871_ gnd vdd FILL
XFILL_5__2516_ gnd vdd FILL
XFILL_5__3496_ gnd vdd FILL
XFILL_8__2225_ gnd vdd FILL
XFILL_2__2738_ gnd vdd FILL
XFILL_0__1822_ gnd vdd FILL
X_3080_ _3080_/A _3141_/A vdd gnd INVX1
XFILL_8__2156_ gnd vdd FILL
XFILL_5__2447_ gnd vdd FILL
XFILL_0__1753_ gnd vdd FILL
X_2100_ _2294_/A _2288_/B _2101_/C vdd gnd NAND2X1
X_2031_ _2031_/A _2077_/A vdd gnd INVX1
XFILL_5__2378_ gnd vdd FILL
XFILL_2__2669_ gnd vdd FILL
XFILL_8__2087_ gnd vdd FILL
XFILL_3__3201_ gnd vdd FILL
XFILL_3__3132_ gnd vdd FILL
XFILL_0__3423_ gnd vdd FILL
X_2933_ _2933_/A _2933_/B _2933_/C _2934_/B vdd gnd OAI21X1
XFILL_0__2305_ gnd vdd FILL
XFILL_3__3063_ gnd vdd FILL
XFILL_8__2989_ gnd vdd FILL
XFILL_3__2014_ gnd vdd FILL
XFILL_0__2236_ gnd vdd FILL
X_2864_ _2864_/A _2915_/A _2864_/C _2865_/C vdd gnd OAI21X1
X_2795_ _2795_/A _2898_/B _2795_/C _3261_/D vdd gnd OAI21X1
XFILL_0__2167_ gnd vdd FILL
X_1815_ _1815_/A _1815_/B _1815_/C _1831_/D vdd gnd NAND3X1
X_1746_ _3233_/Q _1756_/A _2442_/A vdd gnd NAND2X1
XFILL_0__2098_ gnd vdd FILL
XFILL_3__2916_ gnd vdd FILL
XFILL_8_CLKBUF1_insert28 gnd vdd FILL
XFILL_1__2980_ gnd vdd FILL
XFILL_6__2625_ gnd vdd FILL
XFILL_3__2847_ gnd vdd FILL
XFILL_1__1931_ gnd vdd FILL
XFILL_1__1862_ gnd vdd FILL
X_3416_ _3445_/A _3420_/A _3416_/C _3455_/C _3418_/B vdd gnd AOI22X1
XFILL_6__2556_ gnd vdd FILL
X_3347_ _3347_/D vdd _3347_/R _3573_/CLK _3347_/Q vdd gnd DFFSR
XFILL_1__3601_ gnd vdd FILL
XFILL_6__2487_ gnd vdd FILL
XFILL_1__1793_ gnd vdd FILL
XFILL_3__2778_ gnd vdd FILL
XFILL_1__3532_ gnd vdd FILL
XFILL_3__1729_ gnd vdd FILL
XFILL_6_CLKBUF1_insert32 gnd vdd FILL
X_3278_ _3278_/D vdd _3353_/R _3313_/CLK _3278_/Q vdd gnd DFFSR
XFILL_1_BUFX2_insert5 gnd vdd FILL
XFILL_6__3108_ gnd vdd FILL
XFILL_1__3463_ gnd vdd FILL
XFILL_4__3172_ gnd vdd FILL
X_2229_ _2229_/A _2441_/C vdd gnd INVX1
XFILL_1__3394_ gnd vdd FILL
XFILL_1__2414_ gnd vdd FILL
XFILL_4__2123_ gnd vdd FILL
XFILL_6__3039_ gnd vdd FILL
XFILL_1__2345_ gnd vdd FILL
XFILL_4__2054_ gnd vdd FILL
XFILL_7__2803_ gnd vdd FILL
XFILL_1__2276_ gnd vdd FILL
XFILL_7__2734_ gnd vdd FILL
XFILL_4__2956_ gnd vdd FILL
XFILL_7__2665_ gnd vdd FILL
XFILL_4__2887_ gnd vdd FILL
XFILL_4__1907_ gnd vdd FILL
XFILL_2__1971_ gnd vdd FILL
XFILL_4__1838_ gnd vdd FILL
XFILL_7__2596_ gnd vdd FILL
XFILL_4__1769_ gnd vdd FILL
XFILL_8__2010_ gnd vdd FILL
XFILL_4__3508_ gnd vdd FILL
XFILL_5__2301_ gnd vdd FILL
XFILL_7__3217_ gnd vdd FILL
XFILL_4__3439_ gnd vdd FILL
XFILL_5__2232_ gnd vdd FILL
XFILL_2__2523_ gnd vdd FILL
XFILL_2__2454_ gnd vdd FILL
XFILL_7__3148_ gnd vdd FILL
XFILL_5__2163_ gnd vdd FILL
XFILL_7__3079_ gnd vdd FILL
XFILL_8__2912_ gnd vdd FILL
XFILL_2__2385_ gnd vdd FILL
XFILL_5__2094_ gnd vdd FILL
XFILL_8__2843_ gnd vdd FILL
XFILL_4_BUFX2_insert9 gnd vdd FILL
XFILL_2__3006_ gnd vdd FILL
XFILL_0__3070_ gnd vdd FILL
XFILL_8__2774_ gnd vdd FILL
XFILL_0__2021_ gnd vdd FILL
XFILL_5__2996_ gnd vdd FILL
XFILL_8__1725_ gnd vdd FILL
XFILL_5__1947_ gnd vdd FILL
X_2580_ reset _2580_/Y vdd gnd INVX8
XFILL_5__1878_ gnd vdd FILL
XFILL_3__2701_ gnd vdd FILL
XFILL_6__2410_ gnd vdd FILL
XFILL_0__2923_ gnd vdd FILL
XFILL_6__3390_ gnd vdd FILL
XFILL_3__2632_ gnd vdd FILL
XFILL_5__3548_ gnd vdd FILL
XFILL_0__2854_ gnd vdd FILL
XFILL_6__2341_ gnd vdd FILL
X_3201_ _3215_/A _3201_/B _3201_/C _3348_/D vdd gnd OAI21X1
XFILL_5__3479_ gnd vdd FILL
X_3132_ _3342_/Q _3143_/B _3133_/C vdd gnd NAND2X1
XFILL_6__2272_ gnd vdd FILL
XFILL_8__2208_ gnd vdd FILL
XFILL_0__1805_ gnd vdd FILL
XFILL_3__2563_ gnd vdd FILL
XFILL_0__2785_ gnd vdd FILL
XFILL_3__2494_ gnd vdd FILL
XFILL_8__3188_ gnd vdd FILL
XFILL_8__2139_ gnd vdd FILL
XFILL_0__1736_ gnd vdd FILL
X_3063_ _3165_/A _3063_/B _3063_/C _3064_/C vdd gnd OAI21X1
X_2014_ _2824_/A _2910_/A _2270_/A vdd gnd NOR2X1
XFILL_0__3406_ gnd vdd FILL
XFILL_3__3115_ gnd vdd FILL
XFILL_1__2130_ gnd vdd FILL
XFILL_3__3046_ gnd vdd FILL
X_2916_ _2920_/A _2916_/B _2916_/C _2923_/A vdd gnd OAI21X1
XFILL_1__2061_ gnd vdd FILL
X_2847_ _2910_/B _2887_/B _2900_/A vdd gnd NAND2X1
XFILL_0__2219_ gnd vdd FILL
XFILL_6__1987_ gnd vdd FILL
XFILL_0__3199_ gnd vdd FILL
XFILL_4__2810_ gnd vdd FILL
XFILL_4__2741_ gnd vdd FILL
X_2778_ _2778_/A _2778_/B _2778_/C _3254_/D vdd gnd OAI21X1
XFILL_1__2963_ gnd vdd FILL
XFILL_7__2450_ gnd vdd FILL
X_1729_ _3237_/Q _3166_/C _1729_/Y vdd gnd NAND2X1
XFILL_7__2381_ gnd vdd FILL
XFILL_1__1914_ gnd vdd FILL
XFILL_6__3588_ gnd vdd FILL
XFILL_4__2672_ gnd vdd FILL
XFILL_6__2608_ gnd vdd FILL
XFILL_1__2894_ gnd vdd FILL
XFILL_6__2539_ gnd vdd FILL
XFILL_1__1845_ gnd vdd FILL
XFILL_7__3002_ gnd vdd FILL
XFILL_1__1776_ gnd vdd FILL
XFILL_1__3515_ gnd vdd FILL
XFILL_4__3224_ gnd vdd FILL
XFILL_1__3446_ gnd vdd FILL
XFILL_4__3155_ gnd vdd FILL
XFILL_1__3377_ gnd vdd FILL
XFILL_2__2170_ gnd vdd FILL
XFILL_4__3086_ gnd vdd FILL
XFILL_4__2106_ gnd vdd FILL
XFILL_4__2037_ gnd vdd FILL
XFILL_1__2328_ gnd vdd FILL
XFILL_1__2259_ gnd vdd FILL
XFILL_5__2850_ gnd vdd FILL
XFILL_5__2781_ gnd vdd FILL
XFILL_5__1801_ gnd vdd FILL
XFILL_7__2717_ gnd vdd FILL
XFILL_4__2939_ gnd vdd FILL
XFILL_8__2490_ gnd vdd FILL
XFILL_5__1732_ gnd vdd FILL
XFILL_2__1954_ gnd vdd FILL
XFILL_7__2648_ gnd vdd FILL
XFILL_7__2579_ gnd vdd FILL
XFILL_8__3111_ gnd vdd FILL
XFILL_5__3402_ gnd vdd FILL
XFILL_2__1885_ gnd vdd FILL
XFILL_2__3555_ gnd vdd FILL
XFILL_8__3042_ gnd vdd FILL
XFILL_2__2506_ gnd vdd FILL
XFILL_0__2570_ gnd vdd FILL
XFILL_2__3486_ gnd vdd FILL
XFILL_5__2215_ gnd vdd FILL
XFILL_5__3195_ gnd vdd FILL
XFILL_5__2146_ gnd vdd FILL
XFILL_2__2437_ gnd vdd FILL
XFILL_2__2368_ gnd vdd FILL
XFILL_5_BUFX2_insert23 gnd vdd FILL
XFILL_5__2077_ gnd vdd FILL
XFILL_5_BUFX2_insert12 gnd vdd FILL
XFILL_0__3122_ gnd vdd FILL
XFILL_6__2890_ gnd vdd FILL
XFILL_5_BUFX2_insert56 gnd vdd FILL
XFILL_8__2826_ gnd vdd FILL
XFILL_2__2299_ gnd vdd FILL
XFILL_5_BUFX2_insert45 gnd vdd FILL
XFILL_5_BUFX2_insert67 gnd vdd FILL
XFILL_6__1910_ gnd vdd FILL
XFILL_0__3053_ gnd vdd FILL
XFILL_5_BUFX2_insert78 gnd vdd FILL
X_2701_ _3571_/Q _2701_/B _3166_/D _2703_/B vdd gnd NAND3X1
XFILL_6__1841_ gnd vdd FILL
XFILL_5_BUFX2_insert89 gnd vdd FILL
XFILL_0__2004_ gnd vdd FILL
XFILL_8__2757_ gnd vdd FILL
XFILL_6__3511_ gnd vdd FILL
XFILL_5__2979_ gnd vdd FILL
XFILL_6__1772_ gnd vdd FILL
XFILL_8__1708_ gnd vdd FILL
XFILL_8__2688_ gnd vdd FILL
X_2632_ _2632_/A _2748_/B _2728_/A _2633_/C vdd gnd OAI21X1
XFILL_3__1994_ gnd vdd FILL
X_2563_ _2563_/A _3576_/Q _2760_/B _2564_/C vdd gnd AOI21X1
XFILL_6__3442_ gnd vdd FILL
XFILL_6__3373_ gnd vdd FILL
XFILL_0__2906_ gnd vdd FILL
X_2494_ _2563_/A _2570_/B vdd gnd INVX2
XFILL_6__2324_ gnd vdd FILL
XFILL_3__3595_ gnd vdd FILL
XFILL_3__2615_ gnd vdd FILL
XFILL_0__2837_ gnd vdd FILL
XFILL_3__2546_ gnd vdd FILL
X_3115_ _3115_/A _3125_/B _3333_/Q _3116_/C vdd gnd OAI21X1
XFILL_6__2255_ gnd vdd FILL
XFILL_0__2768_ gnd vdd FILL
XFILL_6__2186_ gnd vdd FILL
X_3046_ _3090_/A _3131_/A _3046_/C _3316_/D vdd gnd OAI21X1
XFILL_0__1719_ gnd vdd FILL
XFILL_3__2477_ gnd vdd FILL
XFILL_0__2699_ gnd vdd FILL
XFILL_1__3231_ gnd vdd FILL
XFILL_7__1950_ gnd vdd FILL
XFILL_1__3162_ gnd vdd FILL
XFILL_1__3093_ gnd vdd FILL
XFILL_7__1881_ gnd vdd FILL
XFILL_1__2113_ gnd vdd FILL
XFILL_3__3029_ gnd vdd FILL
XFILL_1__2044_ gnd vdd FILL
XFILL_9__2797_ gnd vdd FILL
XFILL_7__3551_ gnd vdd FILL
XFILL_7__3482_ gnd vdd FILL
XFILL_7__2502_ gnd vdd FILL
XFILL_4__2724_ gnd vdd FILL
XFILL_7__2433_ gnd vdd FILL
XFILL_1__2946_ gnd vdd FILL
XFILL_4__2655_ gnd vdd FILL
XFILL_1__2877_ gnd vdd FILL
XFILL_7__2364_ gnd vdd FILL
XFILL_7__2295_ gnd vdd FILL
XFILL_4__2586_ gnd vdd FILL
XFILL_1__1828_ gnd vdd FILL
XFILL_1__1759_ gnd vdd FILL
XFILL_5__2000_ gnd vdd FILL
XFILL_4__3207_ gnd vdd FILL
XFILL_4__3138_ gnd vdd FILL
XFILL_1__3429_ gnd vdd FILL
XFILL_8__1990_ gnd vdd FILL
XFILL_2__2222_ gnd vdd FILL
XFILL_2__2153_ gnd vdd FILL
XFILL_4__3069_ gnd vdd FILL
XFILL_5__2902_ gnd vdd FILL
XFILL_2__2084_ gnd vdd FILL
XFILL_8__2611_ gnd vdd FILL
XFILL_5__2833_ gnd vdd FILL
XFILL_8__3591_ gnd vdd FILL
XFILL_8__2542_ gnd vdd FILL
XFILL_8__2473_ gnd vdd FILL
XFILL_5__2764_ gnd vdd FILL
XFILL_2__2986_ gnd vdd FILL
XFILL_5__2695_ gnd vdd FILL
XFILL_5__1715_ gnd vdd FILL
XFILL_2__1937_ gnd vdd FILL
XFILL_2__1868_ gnd vdd FILL
XFILL_3__2400_ gnd vdd FILL
XFILL_3__3380_ gnd vdd FILL
XFILL_2__1799_ gnd vdd FILL
XFILL_8__3025_ gnd vdd FILL
XFILL_0__2622_ gnd vdd FILL
XFILL_6__2040_ gnd vdd FILL
XFILL_2__3538_ gnd vdd FILL
XFILL_3__2331_ gnd vdd FILL
XFILL_2__3469_ gnd vdd FILL
XFILL_3__2262_ gnd vdd FILL
XBUFX2_insert6 RDY _2786_/A vdd gnd BUFX2
XFILL_0__2553_ gnd vdd FILL
XFILL_0__2484_ gnd vdd FILL
XFILL_5__3178_ gnd vdd FILL
XFILL_3__2193_ gnd vdd FILL
XFILL_5__2129_ gnd vdd FILL
XFILL_6__2942_ gnd vdd FILL
XFILL_0__3105_ gnd vdd FILL
X_1994_ _3300_/Q _1998_/B vdd gnd INVX1
XFILL_8__2809_ gnd vdd FILL
XFILL_6__2873_ gnd vdd FILL
XFILL_0__3036_ gnd vdd FILL
XFILL_6__1824_ gnd vdd FILL
XFILL_6__1755_ gnd vdd FILL
X_2615_ _3298_/Q _2728_/A _2615_/C _2616_/C vdd gnd OAI21X1
XFILL_3__1977_ gnd vdd FILL
XFILL_1__2800_ gnd vdd FILL
X_3595_ _3595_/A DO[0] vdd gnd BUFX2
XFILL_6__3425_ gnd vdd FILL
X_2546_ _3574_/Q _3063_/C vdd gnd INVX1
XFILL_1_BUFX2_insert10 gnd vdd FILL
XFILL_1__2731_ gnd vdd FILL
XFILL_4__2440_ gnd vdd FILL
X_2477_ _2569_/B _2569_/A _2565_/A vdd gnd OR2X2
XFILL_1_BUFX2_insert21 gnd vdd FILL
XFILL_1_BUFX2_insert43 gnd vdd FILL
XFILL_6_BUFX2_insert0 gnd vdd FILL
XFILL_1__2662_ gnd vdd FILL
XFILL_4__2371_ gnd vdd FILL
XFILL_7__2080_ gnd vdd FILL
XFILL_9__2016_ gnd vdd FILL
XFILL_6__2307_ gnd vdd FILL
XFILL_3_CLKBUF1_insert29 gnd vdd FILL
XFILL_1_BUFX2_insert65 gnd vdd FILL
XFILL_1_BUFX2_insert54 gnd vdd FILL
XFILL_1_BUFX2_insert76 gnd vdd FILL
XFILL_6__2238_ gnd vdd FILL
XFILL_1_BUFX2_insert87 gnd vdd FILL
XFILL_3__2529_ gnd vdd FILL
XFILL_1__2593_ gnd vdd FILL
X_3029_ _3127_/A _3029_/B _3090_/A vdd gnd NAND2X1
XFILL_6__2169_ gnd vdd FILL
XFILL_7__2982_ gnd vdd FILL
XFILL_1__3214_ gnd vdd FILL
XFILL_1_CLKBUF1_insert33 gnd vdd FILL
XFILL_7__1933_ gnd vdd FILL
XFILL_1__3145_ gnd vdd FILL
XFILL_1__3076_ gnd vdd FILL
XFILL_7__1864_ gnd vdd FILL
XFILL_1__2027_ gnd vdd FILL
XFILL_7__3603_ gnd vdd FILL
XFILL_7__1795_ gnd vdd FILL
XFILL_7__3534_ gnd vdd FILL
XFILL_2__2840_ gnd vdd FILL
XFILL_7__3465_ gnd vdd FILL
XFILL_4__2707_ gnd vdd FILL
XFILL_2__2771_ gnd vdd FILL
XFILL_1__2929_ gnd vdd FILL
XFILL_7__3396_ gnd vdd FILL
XFILL_7__2416_ gnd vdd FILL
XFILL_2__1722_ gnd vdd FILL
XFILL_5__2480_ gnd vdd FILL
XFILL_7__2347_ gnd vdd FILL
XFILL_4__2638_ gnd vdd FILL
XFILL_4__2569_ gnd vdd FILL
XFILL_5__3101_ gnd vdd FILL
XFILL_7__2278_ gnd vdd FILL
XFILL_5__3032_ gnd vdd FILL
XFILL_2__2205_ gnd vdd FILL
XFILL_8__1973_ gnd vdd FILL
XFILL_2__3185_ gnd vdd FILL
XFILL_2__2136_ gnd vdd FILL
XFILL_2__2067_ gnd vdd FILL
XFILL_3__1900_ gnd vdd FILL
XFILL_3__2880_ gnd vdd FILL
XFILL_5__2816_ gnd vdd FILL
XFILL_8__2525_ gnd vdd FILL
XBUFX2_insert90 _3027_/Y _3125_/A vdd gnd BUFX2
XFILL_3__1831_ gnd vdd FILL
X_2400_ _2872_/B _3077_/C _3250_/Q _2404_/A vdd gnd OAI21X1
XFILL_5__2747_ gnd vdd FILL
X_3380_ _3565_/A _3383_/B _3381_/C vdd gnd NAND2X1
XFILL_2__2969_ gnd vdd FILL
XFILL_8__2456_ gnd vdd FILL
XFILL_3__1762_ gnd vdd FILL
XFILL_3__3501_ gnd vdd FILL
XFILL_8__2387_ gnd vdd FILL
X_2331_ _2331_/A _2331_/B _2331_/C _2333_/B vdd gnd NAND3X1
XFILL_0__1984_ gnd vdd FILL
XFILL_5__2678_ gnd vdd FILL
X_2262_ _2270_/A _2794_/A _2307_/A vdd gnd NAND2X1
XFILL_6__3210_ gnd vdd FILL
XFILL_3__1693_ gnd vdd FILL
XFILL_6__3141_ gnd vdd FILL
XFILL_3__3432_ gnd vdd FILL
XFILL_8_BUFX2_insert60 gnd vdd FILL
XFILL_8_BUFX2_insert93 gnd vdd FILL
XFILL_8_BUFX2_insert82 gnd vdd FILL
X_2193_ _2340_/A _3151_/B _2342_/A _2196_/C vdd gnd MUX2X1
XFILL_8_BUFX2_insert71 gnd vdd FILL
XFILL_8__3008_ gnd vdd FILL
XFILL_6__3072_ gnd vdd FILL
XFILL_3__2314_ gnd vdd FILL
XFILL_0__3585_ gnd vdd FILL
XFILL_0__2605_ gnd vdd FILL
XFILL_6__2023_ gnd vdd FILL
XFILL_0__2536_ gnd vdd FILL
XFILL_3__2245_ gnd vdd FILL
XFILL_0__2467_ gnd vdd FILL
XFILL_3__2176_ gnd vdd FILL
XFILL_0__2398_ gnd vdd FILL
XFILL_6__2925_ gnd vdd FILL
XFILL_4__1940_ gnd vdd FILL
X_1977_ _3338_/Q _3110_/A _3127_/B _3347_/Q _1979_/C vdd gnd AOI22X1
XFILL_6__2856_ gnd vdd FILL
XFILL_4__1871_ gnd vdd FILL
XFILL_0__3019_ gnd vdd FILL
XFILL_6__1807_ gnd vdd FILL
XFILL_6__2787_ gnd vdd FILL
XFILL_4__3541_ gnd vdd FILL
X_3578_ _3578_/D vdd _3578_/R _3578_/CLK _3578_/Q vdd gnd DFFSR
XFILL_6__1738_ gnd vdd FILL
X_2529_ _2565_/A _3291_/D _2529_/C _2530_/C vdd gnd AOI21X1
XFILL_4__3472_ gnd vdd FILL
XFILL_6__3408_ gnd vdd FILL
XFILL_7__2201_ gnd vdd FILL
XFILL_1__2714_ gnd vdd FILL
XFILL_7__3181_ gnd vdd FILL
XFILL_4__2423_ gnd vdd FILL
XFILL_7__2132_ gnd vdd FILL
XFILL_4__2354_ gnd vdd FILL
XFILL_1__2645_ gnd vdd FILL
XFILL_1__2576_ gnd vdd FILL
XFILL_7__2063_ gnd vdd FILL
XFILL_4__2285_ gnd vdd FILL
XFILL_7__2965_ gnd vdd FILL
XFILL_1__3128_ gnd vdd FILL
XFILL_7__2896_ gnd vdd FILL
XFILL_7__1916_ gnd vdd FILL
XFILL_5__1980_ gnd vdd FILL
XFILL_7__1847_ gnd vdd FILL
XFILL_1__3059_ gnd vdd FILL
XFILL_7__1778_ gnd vdd FILL
XFILL_5__2601_ gnd vdd FILL
XFILL_7__3517_ gnd vdd FILL
XFILL_2__2823_ gnd vdd FILL
XFILL_8__2310_ gnd vdd FILL
XFILL_5__3581_ gnd vdd FILL
XFILL_7__3448_ gnd vdd FILL
XFILL_8__2241_ gnd vdd FILL
XFILL_5__2532_ gnd vdd FILL
XFILL_5__2463_ gnd vdd FILL
XFILL_2__2754_ gnd vdd FILL
XFILL_7__3379_ gnd vdd FILL
XFILL_8__2172_ gnd vdd FILL
XFILL_2__1705_ gnd vdd FILL
XFILL_2__2685_ gnd vdd FILL
XFILL_5__2394_ gnd vdd FILL
XFILL_0__3370_ gnd vdd FILL
XFILL_5__3015_ gnd vdd FILL
XFILL_0__2321_ gnd vdd FILL
XFILL_3__2030_ gnd vdd FILL
XCLKBUF1_insert35 clk _3573_/CLK vdd gnd CLKBUF1
XFILL_8__1956_ gnd vdd FILL
X_2880_ _2880_/A _2895_/A _2881_/C vdd gnd NOR2X1
XFILL_0__2252_ gnd vdd FILL
XFILL_2__3168_ gnd vdd FILL
X_1900_ _2292_/B _3156_/B _3157_/C vdd gnd NOR2X1
XFILL_0__2183_ gnd vdd FILL
X_1831_ _2676_/B _3189_/C _2993_/A _1831_/D _3387_/B vdd gnd OAI22X1
XFILL_2__2119_ gnd vdd FILL
XFILL_2__3099_ gnd vdd FILL
XFILL_8__1887_ gnd vdd FILL
XFILL_6__2710_ gnd vdd FILL
XFILL_3__2932_ gnd vdd FILL
X_1762_ _3234_/Q _1762_/B _1794_/A vdd gnd NOR2X1
XFILL_6__2641_ gnd vdd FILL
XFILL_3__2863_ gnd vdd FILL
X_3501_ _3528_/C _3502_/C vdd gnd INVX1
XFILL_8__3557_ gnd vdd FILL
X_1693_ _2767_/A _1693_/B _1693_/C _3291_/D vdd gnd OAI21X1
X_3432_ _3432_/A _3432_/B _3500_/C _3525_/B vdd gnd OAI21X1
XFILL_9__2281_ gnd vdd FILL
XFILL_6__2572_ gnd vdd FILL
XFILL_3__1814_ gnd vdd FILL
XFILL_8__2508_ gnd vdd FILL
XFILL_8__3488_ gnd vdd FILL
XFILL183150x167850 gnd vdd FILL
XFILL_3__2794_ gnd vdd FILL
X_3363_ _3363_/D vdd _3363_/R _3363_/CLK _3363_/Q vdd gnd DFFSR
XFILL_3__1745_ gnd vdd FILL
XFILL_8__2439_ gnd vdd FILL
XFILL_0__1967_ gnd vdd FILL
X_3294_ _3294_/D vdd _3355_/R _3578_/CLK _3294_/Q vdd gnd DFFSR
X_2314_ _2314_/A _2314_/B _2314_/C _2315_/B vdd gnd NAND3X1
XFILL_3__3415_ gnd vdd FILL
XFILL_0__1898_ gnd vdd FILL
X_2245_ _2245_/A _2245_/B _2245_/C _2246_/C vdd gnd NAND3X1
XFILL_6__3124_ gnd vdd FILL
X_2176_ _2176_/A _2176_/B _2246_/A vdd gnd NOR2X1
XFILL_1__2430_ gnd vdd FILL
XFILL_6__3055_ gnd vdd FILL
XFILL_1__2361_ gnd vdd FILL
XFILL_6__2006_ gnd vdd FILL
XFILL_4__2070_ gnd vdd FILL
XFILL_0__3499_ gnd vdd FILL
XFILL_3__2228_ gnd vdd FILL
XFILL_0__2519_ gnd vdd FILL
XFILL_1__2292_ gnd vdd FILL
XFILL_3__2159_ gnd vdd FILL
XFILL_7__2750_ gnd vdd FILL
XFILL_6__2908_ gnd vdd FILL
XFILL_4__2972_ gnd vdd FILL
XFILL_7__1701_ gnd vdd FILL
XFILL_4__1923_ gnd vdd FILL
XFILL_7__2681_ gnd vdd FILL
XFILL_6__2839_ gnd vdd FILL
XFILL_4_BUFX2_insert91 gnd vdd FILL
XFILL_4_BUFX2_insert80 gnd vdd FILL
XFILL_4__1854_ gnd vdd FILL
XFILL_4__1785_ gnd vdd FILL
XFILL_4__3524_ gnd vdd FILL
XFILL_4__3455_ gnd vdd FILL
XFILL_2__2470_ gnd vdd FILL
XFILL_7__3164_ gnd vdd FILL
XFILL_4__2406_ gnd vdd FILL
XFILL_7__3095_ gnd vdd FILL
XFILL_4__3386_ gnd vdd FILL
XFILL_7__2115_ gnd vdd FILL
XFILL_1__2628_ gnd vdd FILL
XFILL_4__2337_ gnd vdd FILL
XFILL_7__2046_ gnd vdd FILL
XFILL_4__2268_ gnd vdd FILL
XFILL_1__2559_ gnd vdd FILL
XFILL_8__2790_ gnd vdd FILL
XFILL_2__3022_ gnd vdd FILL
XFILL_8__1810_ gnd vdd FILL
XFILL_4__2199_ gnd vdd FILL
XFILL_8__1741_ gnd vdd FILL
XFILL_7__2948_ gnd vdd FILL
XFILL_5__1963_ gnd vdd FILL
XFILL_7__2879_ gnd vdd FILL
XFILL_8__3411_ gnd vdd FILL
XFILL_5__1894_ gnd vdd FILL
XFILL_5__3564_ gnd vdd FILL
XFILL_0__2870_ gnd vdd FILL
XFILL_2__2806_ gnd vdd FILL
XFILL_5__2515_ gnd vdd FILL
XFILL_5__3495_ gnd vdd FILL
XFILL_0__1821_ gnd vdd FILL
XFILL_8__2224_ gnd vdd FILL
XFILL_2__2737_ gnd vdd FILL
XFILL_8__2155_ gnd vdd FILL
XFILL_5__2446_ gnd vdd FILL
XFILL_0__1752_ gnd vdd FILL
X_2030_ _2331_/B _2338_/B _2338_/A _2031_/A vdd gnd NAND3X1
XFILL_5__2377_ gnd vdd FILL
XFILL_2__2668_ gnd vdd FILL
XFILL_3__3200_ gnd vdd FILL
XFILL_0__3422_ gnd vdd FILL
XFILL_8__2086_ gnd vdd FILL
XFILL_2__2599_ gnd vdd FILL
XFILL_3__3131_ gnd vdd FILL
XFILL_3__3062_ gnd vdd FILL
X_2932_ _2932_/A _2932_/B _2932_/C _2934_/C vdd gnd NAND3X1
XFILL_3__2013_ gnd vdd FILL
XFILL_0__2304_ gnd vdd FILL
XFILL_8__2988_ gnd vdd FILL
XFILL_0__2235_ gnd vdd FILL
XFILL_9__1781_ gnd vdd FILL
XFILL_8__1939_ gnd vdd FILL
X_2863_ _2863_/A _2957_/B _2863_/C _3273_/D vdd gnd OAI21X1
XFILL_0__2166_ gnd vdd FILL
X_2794_ _2794_/A _2794_/B _2795_/C vdd gnd NAND2X1
X_1814_ _1814_/A _3174_/A _1815_/B vdd gnd NOR2X1
XFILL_0__2097_ gnd vdd FILL
X_1745_ _3157_/A _2048_/B _2437_/A vdd gnd NAND2X1
XFILL_3__2915_ gnd vdd FILL
XFILL_1__1930_ gnd vdd FILL
XFILL_6__2624_ gnd vdd FILL
XFILL_3__2846_ gnd vdd FILL
XFILL_8_CLKBUF1_insert29 gnd vdd FILL
XFILL_6__2555_ gnd vdd FILL
X_3415_ _3421_/B _3417_/B _3416_/C vdd gnd NAND2X1
XFILL_1__1861_ gnd vdd FILL
XFILL_3__2777_ gnd vdd FILL
X_3346_ _3346_/D vdd _3346_/R _3346_/CLK _3346_/Q vdd gnd DFFSR
XFILL_0__2999_ gnd vdd FILL
XFILL_1__3600_ gnd vdd FILL
XFILL_1__1792_ gnd vdd FILL
XFILL_6__2486_ gnd vdd FILL
XFILL_3__1728_ gnd vdd FILL
XFILL_1__3531_ gnd vdd FILL
XFILL_6_CLKBUF1_insert33 gnd vdd FILL
X_3277_ _3277_/D vdd _3282_/R _3284_/CLK _3277_/Q vdd gnd DFFSR
XFILL_1_BUFX2_insert6 gnd vdd FILL
XFILL_6__3107_ gnd vdd FILL
XFILL_1__3462_ gnd vdd FILL
X_2228_ _2228_/A _2228_/B _3234_/D vdd gnd OR2X2
XFILL_4__3171_ gnd vdd FILL
XFILL_1__3393_ gnd vdd FILL
XFILL_4__2122_ gnd vdd FILL
X_2159_ _2304_/C _3233_/D vdd gnd INVX1
XFILL_1__2413_ gnd vdd FILL
XFILL_6__3038_ gnd vdd FILL
XFILL_1__2344_ gnd vdd FILL
XFILL_4__2053_ gnd vdd FILL
XFILL_7__2802_ gnd vdd FILL
XFILL_1__2275_ gnd vdd FILL
XFILL_7__2733_ gnd vdd FILL
XFILL_4__2955_ gnd vdd FILL
XFILL_7__2664_ gnd vdd FILL
XFILL_4__2886_ gnd vdd FILL
XFILL_2__1970_ gnd vdd FILL
XFILL_4__1906_ gnd vdd FILL
XFILL_7__2595_ gnd vdd FILL
XFILL_4__1837_ gnd vdd FILL
XFILL_4__1768_ gnd vdd FILL
XFILL_5__2300_ gnd vdd FILL
XFILL_4__3507_ gnd vdd FILL
XFILL_7__3216_ gnd vdd FILL
XFILL_4__1699_ gnd vdd FILL
XFILL_2__2522_ gnd vdd FILL
XFILL_4__3438_ gnd vdd FILL
XFILL_7__3147_ gnd vdd FILL
XFILL_5__2231_ gnd vdd FILL
XFILL_5__2162_ gnd vdd FILL
XFILL_4__3369_ gnd vdd FILL
XFILL_2__2453_ gnd vdd FILL
XFILL_7__3078_ gnd vdd FILL
XFILL_2__2384_ gnd vdd FILL
XFILL_8__2911_ gnd vdd FILL
XFILL_7__2029_ gnd vdd FILL
XFILL_5__2093_ gnd vdd FILL
XFILL_8__2842_ gnd vdd FILL
XFILL_2__3005_ gnd vdd FILL
XFILL_8__2773_ gnd vdd FILL
XFILL_0__2020_ gnd vdd FILL
XFILL_5__2995_ gnd vdd FILL
XFILL_8__1724_ gnd vdd FILL
XFILL_5__1946_ gnd vdd FILL
XFILL_5__1877_ gnd vdd FILL
XFILL_3__2700_ gnd vdd FILL
XFILL_0__2922_ gnd vdd FILL
XFILL_3__2631_ gnd vdd FILL
XFILL_5__3547_ gnd vdd FILL
XFILL_0__2853_ gnd vdd FILL
XFILL_6__2340_ gnd vdd FILL
X_3200_ _3214_/A _3214_/B _3348_/Q _3201_/C vdd gnd OAI21X1
XFILL_5__3478_ gnd vdd FILL
X_3131_ _3131_/A _3143_/B _3131_/C _3341_/D vdd gnd OAI21X1
XFILL_6__2271_ gnd vdd FILL
XFILL_8__2207_ gnd vdd FILL
XFILL_0__1804_ gnd vdd FILL
XFILL_3__2562_ gnd vdd FILL
XFILL_0__2784_ gnd vdd FILL
XFILL_3__2493_ gnd vdd FILL
XFILL_8__3187_ gnd vdd FILL
XFILL_5__2429_ gnd vdd FILL
X_3062_ _3090_/A _3135_/A _3062_/C _3318_/D vdd gnd OAI21X1
XFILL_0__1735_ gnd vdd FILL
XFILL_8__2138_ gnd vdd FILL
X_2013_ _2854_/A _2890_/A _2910_/A vdd gnd NAND2X1
XFILL_8__2069_ gnd vdd FILL
XFILL_3__3114_ gnd vdd FILL
XFILL_0__3405_ gnd vdd FILL
XFILL_3__3045_ gnd vdd FILL
X_2915_ _2915_/A _2932_/B _2915_/C _2916_/B vdd gnd OAI21X1
XFILL_1__2060_ gnd vdd FILL
X_2846_ _2928_/B _2908_/A _2846_/C _2858_/A vdd gnd OAI21X1
XFILL_6__1986_ gnd vdd FILL
XFILL_0__2218_ gnd vdd FILL
XFILL_0__3198_ gnd vdd FILL
XFILL_0__2149_ gnd vdd FILL
X_2777_ _3254_/Q _2778_/A _2778_/C vdd gnd NAND2X1
XFILL_4__2740_ gnd vdd FILL
XFILL_1__2962_ gnd vdd FILL
X_1728_ _3238_/Q _3166_/C vdd gnd INVX2
XFILL_4__2671_ gnd vdd FILL
XFILL_1__2893_ gnd vdd FILL
XFILL_6__3587_ gnd vdd FILL
XFILL_7__2380_ gnd vdd FILL
XFILL_1__1913_ gnd vdd FILL
XFILL_6__2607_ gnd vdd FILL
XFILL_3__2829_ gnd vdd FILL
XFILL_1__1844_ gnd vdd FILL
XFILL_6__2538_ gnd vdd FILL
XFILL_6__2469_ gnd vdd FILL
X_3329_ _3329_/D vdd _3346_/R _3346_/CLK _3329_/Q vdd gnd DFFSR
XFILL_7__3001_ gnd vdd FILL
XFILL_1__1775_ gnd vdd FILL
XFILL_9__2178_ gnd vdd FILL
XFILL_1__3514_ gnd vdd FILL
XFILL_4__3223_ gnd vdd FILL
XFILL_1__3445_ gnd vdd FILL
XFILL_4__3154_ gnd vdd FILL
XFILL_1__3376_ gnd vdd FILL
XFILL_4__3085_ gnd vdd FILL
XFILL_4__2105_ gnd vdd FILL
XFILL_4__2036_ gnd vdd FILL
XFILL_1__2327_ gnd vdd FILL
XFILL_1__2258_ gnd vdd FILL
XFILL_1__2189_ gnd vdd FILL
XFILL_7__2716_ gnd vdd FILL
XFILL_5__2780_ gnd vdd FILL
XFILL_5__1800_ gnd vdd FILL
XFILL_4__2938_ gnd vdd FILL
XFILL_5__1731_ gnd vdd FILL
XFILL_2__1953_ gnd vdd FILL
XFILL_7__2647_ gnd vdd FILL
XFILL_7__2578_ gnd vdd FILL
XFILL_4__2869_ gnd vdd FILL
XFILL_8__3110_ gnd vdd FILL
XFILL_5__3401_ gnd vdd FILL
XFILL_2__1884_ gnd vdd FILL
XFILL_8__3041_ gnd vdd FILL
XFILL_2__3554_ gnd vdd FILL
XFILL_2__3485_ gnd vdd FILL
XFILL_5__2214_ gnd vdd FILL
XFILL_2__2505_ gnd vdd FILL
XFILL_5__3194_ gnd vdd FILL
XFILL_2__2436_ gnd vdd FILL
XFILL_5__2145_ gnd vdd FILL
XFILL_5__2076_ gnd vdd FILL
XFILL_2__2367_ gnd vdd FILL
XFILL_2__2298_ gnd vdd FILL
XFILL_5_BUFX2_insert24 gnd vdd FILL
XFILL_5_BUFX2_insert13 gnd vdd FILL
XFILL_5_BUFX2_insert57 gnd vdd FILL
XFILL_0__3121_ gnd vdd FILL
XFILL_8__2825_ gnd vdd FILL
XFILL_5_BUFX2_insert68 gnd vdd FILL
XFILL_5_BUFX2_insert46 gnd vdd FILL
XFILL_5_BUFX2_insert79 gnd vdd FILL
XFILL_0__3052_ gnd vdd FILL
X_2700_ _3219_/A _2700_/B _2711_/B _2746_/B _2704_/A vdd gnd OAI22X1
XFILL_6__1840_ gnd vdd FILL
XFILL_0__2003_ gnd vdd FILL
XFILL_6__1771_ gnd vdd FILL
XFILL_8__2756_ gnd vdd FILL
XFILL_6__3510_ gnd vdd FILL
XFILL_5__2978_ gnd vdd FILL
XFILL_3__1993_ gnd vdd FILL
XFILL_8__1707_ gnd vdd FILL
XFILL_8__2687_ gnd vdd FILL
X_2631_ _2770_/C _2748_/B vdd gnd INVX2
XFILL_5__1929_ gnd vdd FILL
X_2562_ _3253_/Q _2768_/B vdd gnd INVX1
XFILL_6__3441_ gnd vdd FILL
XFILL_9__3150_ gnd vdd FILL
XFILL_0__2905_ gnd vdd FILL
XFILL_6__3372_ gnd vdd FILL
X_2493_ _3353_/Q _2650_/A vdd gnd INVX1
XFILL_6__2323_ gnd vdd FILL
XFILL_3__3594_ gnd vdd FILL
XFILL_3__2614_ gnd vdd FILL
XFILL_0__2836_ gnd vdd FILL
XFILL_3__2545_ gnd vdd FILL
X_3114_ _3131_/A _3126_/B _3114_/C _3332_/D vdd gnd OAI21X1
XFILL_6__2254_ gnd vdd FILL
XFILL_0__2767_ gnd vdd FILL
XFILL_6__2185_ gnd vdd FILL
X_3045_ _3316_/Q _3090_/A _3046_/C vdd gnd NAND2X1
XFILL_3__2476_ gnd vdd FILL
XFILL_0__1718_ gnd vdd FILL
XFILL_0__2698_ gnd vdd FILL
XFILL_1__3230_ gnd vdd FILL
XFILL_1__3161_ gnd vdd FILL
XFILL_1__2112_ gnd vdd FILL
XFILL_3__3028_ gnd vdd FILL
XFILL_7__1880_ gnd vdd FILL
XFILL_1__3092_ gnd vdd FILL
XFILL_1__2043_ gnd vdd FILL
XFILL_7__3550_ gnd vdd FILL
X_2829_ _2835_/A _2832_/B vdd gnd INVX1
XFILL_6__1969_ gnd vdd FILL
XFILL_7__3481_ gnd vdd FILL
XFILL_7__2501_ gnd vdd FILL
XFILL_1__2945_ gnd vdd FILL
XFILL_4__2723_ gnd vdd FILL
XFILL_7__2432_ gnd vdd FILL
XFILL_7__2363_ gnd vdd FILL
XFILL_4__2654_ gnd vdd FILL
XFILL_1__2876_ gnd vdd FILL
XFILL_4__2585_ gnd vdd FILL
XFILL_1__1827_ gnd vdd FILL
XFILL_7__2294_ gnd vdd FILL
XFILL_1__1758_ gnd vdd FILL
XFILL_1__1689_ gnd vdd FILL
XFILL_4__3206_ gnd vdd FILL
XFILL_4__3137_ gnd vdd FILL
XFILL_1__3428_ gnd vdd FILL
XFILL_2__2221_ gnd vdd FILL
XFILL_2__2152_ gnd vdd FILL
XFILL_4__3068_ gnd vdd FILL
XFILL_2__2083_ gnd vdd FILL
XFILL_5__2901_ gnd vdd FILL
XFILL_4__2019_ gnd vdd FILL
XFILL_8__2610_ gnd vdd FILL
XFILL_5__2832_ gnd vdd FILL
XFILL_8__3590_ gnd vdd FILL
XFILL_8__2541_ gnd vdd FILL
XFILL_8__2472_ gnd vdd FILL
XFILL_5__2763_ gnd vdd FILL
XFILL_2__2985_ gnd vdd FILL
XFILL_5__2694_ gnd vdd FILL
XFILL_5__1714_ gnd vdd FILL
XFILL_2__1936_ gnd vdd FILL
XFILL_2__1867_ gnd vdd FILL
XFILL_2__3537_ gnd vdd FILL
XFILL_3__2330_ gnd vdd FILL
XFILL_8__3024_ gnd vdd FILL
XFILL_0__2621_ gnd vdd FILL
XFILL_2__1798_ gnd vdd FILL
XFILL_0__2552_ gnd vdd FILL
XFILL_2__3468_ gnd vdd FILL
XFILL_3__2261_ gnd vdd FILL
XBUFX2_insert7 RDY _3197_/C vdd gnd BUFX2
XFILL_5__3177_ gnd vdd FILL
XFILL182850x140550 gnd vdd FILL
XFILL_2__3399_ gnd vdd FILL
XFILL_2__2419_ gnd vdd FILL
XFILL_0__2483_ gnd vdd FILL
XFILL_5__2128_ gnd vdd FILL
XFILL_3__2192_ gnd vdd FILL
XFILL_6__2941_ gnd vdd FILL
XFILL_5__2059_ gnd vdd FILL
XFILL_0__3104_ gnd vdd FILL
X_1993_ _2906_/A _2888_/B _1993_/Y vdd gnd NOR2X1
XFILL_8__2808_ gnd vdd FILL
XFILL_6__2872_ gnd vdd FILL
XFILL_0__3035_ gnd vdd FILL
XFILL_6__1823_ gnd vdd FILL
XFILL_8__2739_ gnd vdd FILL
XFILL_6__1754_ gnd vdd FILL
X_2614_ _3349_/Q _2770_/C _2615_/C vdd gnd NAND2X1
XFILL_3__1976_ gnd vdd FILL
X_3594_ _3594_/A AB[9] vdd gnd BUFX2
XFILL_6__3424_ gnd vdd FILL
X_2545_ _3360_/Q _3226_/A vdd gnd INVX1
X_2476_ _2508_/B _2479_/A vdd gnd INVX1
XFILL_1__2730_ gnd vdd FILL
XFILL_1_BUFX2_insert22 gnd vdd FILL
XFILL_1_BUFX2_insert11 gnd vdd FILL
XFILL_6_BUFX2_insert1 gnd vdd FILL
XFILL_1__2661_ gnd vdd FILL
XFILL_0__2819_ gnd vdd FILL
XFILL_4__2370_ gnd vdd FILL
XFILL_6__2306_ gnd vdd FILL
XFILL_1_BUFX2_insert66 gnd vdd FILL
XFILL_1_BUFX2_insert44 gnd vdd FILL
XFILL_1_BUFX2_insert55 gnd vdd FILL
XFILL_1_BUFX2_insert77 gnd vdd FILL
XFILL_6__2237_ gnd vdd FILL
XFILL_1_BUFX2_insert88 gnd vdd FILL
XFILL_3__2528_ gnd vdd FILL
XFILL_1__2592_ gnd vdd FILL
XFILL_3__2459_ gnd vdd FILL
X_3028_ _3111_/A _3127_/A vdd gnd INVX1
XFILL_6__2168_ gnd vdd FILL
XFILL_7__2981_ gnd vdd FILL
XFILL_1__3213_ gnd vdd FILL
XFILL_6__2099_ gnd vdd FILL
XFILL_1_CLKBUF1_insert34 gnd vdd FILL
XFILL_7__1932_ gnd vdd FILL
XFILL_1__3144_ gnd vdd FILL
XFILL_1__3075_ gnd vdd FILL
XFILL_7__1863_ gnd vdd FILL
XFILL_1__2026_ gnd vdd FILL
XFILL_7__3602_ gnd vdd FILL
XFILL_7__1794_ gnd vdd FILL
XFILL_7__3533_ gnd vdd FILL
XFILL_7__3464_ gnd vdd FILL
XFILL_4__2706_ gnd vdd FILL
XFILL_2__2770_ gnd vdd FILL
XFILL_1__2928_ gnd vdd FILL
XFILL_7__3395_ gnd vdd FILL
XFILL_7__2415_ gnd vdd FILL
XFILL_2__1721_ gnd vdd FILL
XFILL_7__2346_ gnd vdd FILL
XFILL_4__2637_ gnd vdd FILL
XFILL_1__2859_ gnd vdd FILL
XFILL_4__2568_ gnd vdd FILL
XFILL_5__3100_ gnd vdd FILL
XFILL_4__2499_ gnd vdd FILL
XFILL_7__2277_ gnd vdd FILL
XFILL_5__3031_ gnd vdd FILL
XFILL_2__2204_ gnd vdd FILL
XFILL_8__1972_ gnd vdd FILL
XFILL_2__3184_ gnd vdd FILL
XFILL_2__2135_ gnd vdd FILL
XFILL_2__2066_ gnd vdd FILL
XFILL_5__2815_ gnd vdd FILL
XFILL_8__2524_ gnd vdd FILL
XBUFX2_insert91 _3027_/Y _3111_/A vdd gnd BUFX2
XBUFX2_insert80 _1694_/Y _2242_/A vdd gnd BUFX2
XFILL_5__2746_ gnd vdd FILL
XFILL_3__1830_ gnd vdd FILL
XFILL_2__2968_ gnd vdd FILL
XFILL_8__2455_ gnd vdd FILL
XFILL_3__1761_ gnd vdd FILL
XFILL_3__3500_ gnd vdd FILL
XFILL_2__1919_ gnd vdd FILL
X_2330_ _2330_/A _2330_/B _2331_/C vdd gnd AND2X2
XFILL_8__2386_ gnd vdd FILL
XFILL_5__2677_ gnd vdd FILL
XFILL_0__1983_ gnd vdd FILL
XFILL_2__2899_ gnd vdd FILL
XFILL_3__3431_ gnd vdd FILL
X_2261_ _2798_/B _2261_/B _2794_/A vdd gnd NOR2X1
XFILL_3__1692_ gnd vdd FILL
XFILL_6__3140_ gnd vdd FILL
XFILL_8_BUFX2_insert50 gnd vdd FILL
XFILL_8_BUFX2_insert61 gnd vdd FILL
XFILL_8_BUFX2_insert94 gnd vdd FILL
XFILL_8_BUFX2_insert83 gnd vdd FILL
XFILL_6__3071_ gnd vdd FILL
X_2192_ _3237_/Q _2448_/B _3151_/B vdd gnd NOR2X1
XFILL_0__2604_ gnd vdd FILL
XFILL_8_BUFX2_insert72 gnd vdd FILL
XFILL_6__2022_ gnd vdd FILL
XFILL_8__3007_ gnd vdd FILL
XFILL_3__2313_ gnd vdd FILL
XFILL_0__3584_ gnd vdd FILL
XFILL_3__2244_ gnd vdd FILL
XFILL_0__2535_ gnd vdd FILL
XFILL_5__3229_ gnd vdd FILL
XFILL_0__2466_ gnd vdd FILL
XFILL_3__2175_ gnd vdd FILL
XFILL_0__2397_ gnd vdd FILL
XFILL_6__2924_ gnd vdd FILL
X_1976_ _3330_/Q _3092_/A _1979_/A vdd gnd NAND2X1
XFILL_6__2855_ gnd vdd FILL
XFILL_4__1870_ gnd vdd FILL
XFILL_0__3018_ gnd vdd FILL
XFILL_6__1806_ gnd vdd FILL
XFILL_6__2786_ gnd vdd FILL
XFILL_4__3540_ gnd vdd FILL
X_3577_ _3577_/D vdd _3578_/R _3577_/CLK _3577_/Q vdd gnd DFFSR
XFILL_6__1737_ gnd vdd FILL
XFILL_3__1959_ gnd vdd FILL
X_2528_ _3219_/A _2572_/B _2528_/C _2529_/C vdd gnd OAI21X1
XFILL_4__3471_ gnd vdd FILL
XFILL_6__3407_ gnd vdd FILL
XFILL_7__2200_ gnd vdd FILL
XFILL_1__2713_ gnd vdd FILL
XFILL_7__3180_ gnd vdd FILL
XFILL_4__2422_ gnd vdd FILL
X_2459_ _3290_/D _2502_/B _2502_/C _3348_/Q _2460_/B vdd gnd AOI22X1
XFILL_7__2131_ gnd vdd FILL
XFILL_9__3047_ gnd vdd FILL
XFILL_4__2353_ gnd vdd FILL
XFILL_1__2644_ gnd vdd FILL
XFILL_1__2575_ gnd vdd FILL
XFILL_7__2062_ gnd vdd FILL
XFILL_4__2284_ gnd vdd FILL
XFILL_7__2964_ gnd vdd FILL
XFILL_1__3127_ gnd vdd FILL
XFILL_7__2895_ gnd vdd FILL
XFILL_7__1915_ gnd vdd FILL
XFILL_1__3058_ gnd vdd FILL
XFILL_7__1846_ gnd vdd FILL
XFILL_1__2009_ gnd vdd FILL
XFILL_7__1777_ gnd vdd FILL
XFILL_5__2600_ gnd vdd FILL
XFILL_7__3516_ gnd vdd FILL
XFILL_4__1999_ gnd vdd FILL
XFILL_2__2822_ gnd vdd FILL
XFILL_5__3580_ gnd vdd FILL
XFILL_7__3447_ gnd vdd FILL
XFILL_8__2240_ gnd vdd FILL
XFILL_5__2531_ gnd vdd FILL
XFILL_5__2462_ gnd vdd FILL
XFILL_2__2753_ gnd vdd FILL
XFILL_7__3378_ gnd vdd FILL
XFILL_8__2171_ gnd vdd FILL
XFILL_5__2393_ gnd vdd FILL
XFILL_2__1704_ gnd vdd FILL
XFILL_2__2684_ gnd vdd FILL
XFILL_7__2329_ gnd vdd FILL
XFILL_5__3014_ gnd vdd FILL
XFILL_0__2320_ gnd vdd FILL
XFILL_0__2251_ gnd vdd FILL
XFILL_8__1955_ gnd vdd FILL
XCLKBUF1_insert36 clk _3355_/CLK vdd gnd CLKBUF1
XFILL_2__3167_ gnd vdd FILL
XFILL_0__2182_ gnd vdd FILL
XFILL_2__2118_ gnd vdd FILL
X_1830_ _3246_/Q _2676_/B vdd gnd INVX2
XFILL_2__3098_ gnd vdd FILL
XFILL_8__1886_ gnd vdd FILL
XFILL_3__2931_ gnd vdd FILL
X_3500_ _3525_/B _3525_/A _3500_/C _3528_/C vdd gnd OAI21X1
XFILL_2__2049_ gnd vdd FILL
X_1761_ _3235_/Q _3236_/Q _1858_/B vdd gnd AND2X2
XFILL_6__2640_ gnd vdd FILL
XFILL_3__2862_ gnd vdd FILL
XFILL_8__3556_ gnd vdd FILL
X_1692_ _2767_/A DI[1] _1693_/C vdd gnd NAND2X1
XFILL_8__3487_ gnd vdd FILL
X_3431_ _3431_/A _3431_/B _3432_/B vdd gnd AND2X2
XFILL_8__2507_ gnd vdd FILL
XFILL_6__2571_ gnd vdd FILL
XFILL_3__1813_ gnd vdd FILL
XFILL_3__2793_ gnd vdd FILL
X_3362_ _3362_/D vdd _3362_/R _3362_/CLK _3362_/Q vdd gnd DFFSR
XFILL_5__2729_ gnd vdd FILL
XFILL_8__2438_ gnd vdd FILL
X_2313_ _2313_/A _2313_/B _2314_/B vdd gnd NOR2X1
XFILL_3__1744_ gnd vdd FILL
XFILL_0__1966_ gnd vdd FILL
XFILL184650x132750 gnd vdd FILL
X_3293_ _3293_/D vdd _3353_/R _3578_/CLK _3293_/Q vdd gnd DFFSR
XFILL_8__2369_ gnd vdd FILL
XFILL184350x140550 gnd vdd FILL
XFILL_3__3414_ gnd vdd FILL
X_2244_ _2244_/A _2244_/B _2245_/C vdd gnd NOR2X1
XFILL_0__1897_ gnd vdd FILL
XFILL_6__3123_ gnd vdd FILL
X_2175_ _2278_/A _2437_/C _2374_/C _2176_/B vdd gnd NAND3X1
XFILL_1__2360_ gnd vdd FILL
XFILL_6__3054_ gnd vdd FILL
XFILL_6__2005_ gnd vdd FILL
XFILL_0__2518_ gnd vdd FILL
XFILL_0__3498_ gnd vdd FILL
XFILL_3__2227_ gnd vdd FILL
XFILL_1__2291_ gnd vdd FILL
XFILL_3__2158_ gnd vdd FILL
XFILL_0__2449_ gnd vdd FILL
XFILL_6__2907_ gnd vdd FILL
XFILL_7__1700_ gnd vdd FILL
XFILL_4__2971_ gnd vdd FILL
XFILL_3__2089_ gnd vdd FILL
X_1959_ _1959_/A _1959_/B _1959_/C _2499_/A vdd gnd NAND3X1
XFILL_4__1922_ gnd vdd FILL
XFILL_7__2680_ gnd vdd FILL
XFILL_6__2838_ gnd vdd FILL
XFILL_4_BUFX2_insert92 gnd vdd FILL
XFILL_4_BUFX2_insert81 gnd vdd FILL
XFILL_4_BUFX2_insert70 gnd vdd FILL
XFILL_4__1853_ gnd vdd FILL
XFILL_6__2769_ gnd vdd FILL
XFILL_4__1784_ gnd vdd FILL
XFILL_4__3523_ gnd vdd FILL
XFILL_7__3232_ gnd vdd FILL
XFILL_4__3454_ gnd vdd FILL
XFILL_4__2405_ gnd vdd FILL
XFILL_7__3163_ gnd vdd FILL
XFILL_7__3094_ gnd vdd FILL
XFILL_4__3385_ gnd vdd FILL
XFILL_7__2114_ gnd vdd FILL
XFILL_1__2627_ gnd vdd FILL
XFILL_7__2045_ gnd vdd FILL
XFILL_4__2336_ gnd vdd FILL
XFILL_4__2267_ gnd vdd FILL
XFILL_1__2558_ gnd vdd FILL
XFILL_1__2489_ gnd vdd FILL
XFILL_2__3021_ gnd vdd FILL
XFILL_4__2198_ gnd vdd FILL
XFILL_7__2947_ gnd vdd FILL
XFILL_8__1740_ gnd vdd FILL
XFILL_5__1962_ gnd vdd FILL
XFILL_7__2878_ gnd vdd FILL
XFILL_8__3410_ gnd vdd FILL
XFILL_7__1829_ gnd vdd FILL
XFILL_5__1893_ gnd vdd FILL
XFILL_5__3563_ gnd vdd FILL
XFILL_2__2805_ gnd vdd FILL
XFILL_0__1820_ gnd vdd FILL
XFILL_5__2514_ gnd vdd FILL
XFILL_5__3494_ gnd vdd FILL
XFILL_2__2736_ gnd vdd FILL
XFILL_8__2223_ gnd vdd FILL
XFILL_8__2154_ gnd vdd FILL
XFILL_0__1751_ gnd vdd FILL
XFILL_5__2445_ gnd vdd FILL
XFILL_5__2376_ gnd vdd FILL
XFILL_2__2667_ gnd vdd FILL
XFILL_8__2085_ gnd vdd FILL
XFILL_0__3421_ gnd vdd FILL
XFILL_2__2598_ gnd vdd FILL
XFILL_3__3130_ gnd vdd FILL
XFILL_3__3061_ gnd vdd FILL
X_2931_ _2931_/A _2931_/B _2931_/C _2934_/A vdd gnd NAND3X1
XFILL_3__2012_ gnd vdd FILL
XFILL_0__2303_ gnd vdd FILL
XFILL_2__3219_ gnd vdd FILL
XFILL_8__2987_ gnd vdd FILL
XFILL_0__2234_ gnd vdd FILL
XFILL_8__1938_ gnd vdd FILL
X_2862_ _2862_/A _2863_/C vdd gnd INVX1
XFILL_8__1869_ gnd vdd FILL
XFILL_0__2165_ gnd vdd FILL
X_2793_ _2821_/A _2794_/B vdd gnd INVX1
X_1813_ _3237_/Q _2446_/B _1841_/B _1814_/A vdd gnd OAI21X1
XFILL_3__2914_ gnd vdd FILL
XFILL_0__2096_ gnd vdd FILL
X_1744_ _2594_/A _2057_/A _2048_/B vdd gnd NOR2X1
XFILL_8__3539_ gnd vdd FILL
XFILL_6__2623_ gnd vdd FILL
XFILL_3__2845_ gnd vdd FILL
XFILL184350x152250 gnd vdd FILL
XFILL184650x144450 gnd vdd FILL
X_3414_ _3453_/B _3420_/A _3417_/B vdd gnd AND2X2
XFILL_6__2554_ gnd vdd FILL
XFILL_1__1860_ gnd vdd FILL
XFILL184050x160050 gnd vdd FILL
XFILL_3__2776_ gnd vdd FILL
X_3345_ _3345_/D vdd _3345_/R _3576_/CLK _3345_/Q vdd gnd DFFSR
XFILL_0__2998_ gnd vdd FILL
XFILL_1__1791_ gnd vdd FILL
XFILL_6__2485_ gnd vdd FILL
XFILL_3__1727_ gnd vdd FILL
X_3276_ _3276_/D vdd _3289_/R _3307_/CLK _3276_/Q vdd gnd DFFSR
XFILL_1__3530_ gnd vdd FILL
XFILL_0__1949_ gnd vdd FILL
XFILL_6_CLKBUF1_insert34 gnd vdd FILL
XFILL_1__3461_ gnd vdd FILL
X_2227_ _2296_/B _2304_/A _2228_/A vdd gnd NAND2X1
XFILL_1_BUFX2_insert7 gnd vdd FILL
XFILL_6__3106_ gnd vdd FILL
XFILL_1__2412_ gnd vdd FILL
XFILL_4__3170_ gnd vdd FILL
XFILL_1__3392_ gnd vdd FILL
X_2158_ _2228_/B _2158_/B _2282_/A _2304_/C vdd gnd NOR3X1
XFILL_4__2121_ gnd vdd FILL
XFILL_6__3037_ gnd vdd FILL
XFILL_1__2343_ gnd vdd FILL
X_2089_ _2212_/A _3189_/A _2298_/A _2090_/C vdd gnd OAI21X1
XFILL_4__2052_ gnd vdd FILL
XFILL_1__2274_ gnd vdd FILL
XFILL_7__2801_ gnd vdd FILL
XFILL_7__2732_ gnd vdd FILL
XFILL_4__2954_ gnd vdd FILL
XFILL_7__2663_ gnd vdd FILL
XFILL_4__2885_ gnd vdd FILL
XFILL_4__1905_ gnd vdd FILL
XFILL_4__1836_ gnd vdd FILL
XFILL_7__2594_ gnd vdd FILL
XFILL_4__1767_ gnd vdd FILL
XFILL_4__3506_ gnd vdd FILL
XFILL_1__1989_ gnd vdd FILL
XFILL_7__3215_ gnd vdd FILL
XFILL_2__2521_ gnd vdd FILL
XFILL_4__1698_ gnd vdd FILL
XFILL_4__3437_ gnd vdd FILL
XFILL_7__3146_ gnd vdd FILL
XFILL_5__2230_ gnd vdd FILL
XFILL_5__2161_ gnd vdd FILL
XFILL_4__3368_ gnd vdd FILL
XFILL_2__2452_ gnd vdd FILL
XFILL_7__3077_ gnd vdd FILL
XFILL_2__2383_ gnd vdd FILL
XFILL_4__2319_ gnd vdd FILL
XFILL_8__2910_ gnd vdd FILL
XFILL_0_BUFX2_insert90 gnd vdd FILL
XFILL_7__2028_ gnd vdd FILL
XFILL_5__2092_ gnd vdd FILL
XFILL_8__2841_ gnd vdd FILL
XFILL_2__3004_ gnd vdd FILL
XFILL_8__2772_ gnd vdd FILL
XFILL_5__2994_ gnd vdd FILL
XFILL_8__1723_ gnd vdd FILL
XFILL_5__1945_ gnd vdd FILL
XFILL_5__1876_ gnd vdd FILL
XFILL_0__2921_ gnd vdd FILL
XFILL_3__2630_ gnd vdd FILL
XFILL_5__3546_ gnd vdd FILL
XFILL_0__2852_ gnd vdd FILL
XFILL_5__3477_ gnd vdd FILL
X_3130_ _3341_/Q _3143_/B _3131_/C vdd gnd NAND2X1
XFILL_6__2270_ gnd vdd FILL
XFILL_0__2783_ gnd vdd FILL
XFILL_8__2206_ gnd vdd FILL
XFILL_0__1803_ gnd vdd FILL
XFILL_3__2561_ gnd vdd FILL
XFILL_5__2428_ gnd vdd FILL
XFILL_3__2492_ gnd vdd FILL
XFILL_2__2719_ gnd vdd FILL
XFILL_8__3186_ gnd vdd FILL
XFILL_0__1734_ gnd vdd FILL
X_3061_ _3318_/Q _3090_/A _3062_/C vdd gnd NAND2X1
XFILL_8__2137_ gnd vdd FILL
XFILL_5__2359_ gnd vdd FILL
X_2012_ _2889_/C _2179_/A _2890_/A vdd gnd NAND2X1
XFILL_8__2068_ gnd vdd FILL
XFILL_3__3113_ gnd vdd FILL
XFILL_0__3404_ gnd vdd FILL
XFILL_3__3044_ gnd vdd FILL
X_2914_ _3287_/Q _2919_/A vdd gnd INVX1
XFILL_9__3502_ gnd vdd FILL
XFILL184650x156150 gnd vdd FILL
X_2845_ _2845_/A _2851_/A _2908_/A vdd gnd NAND2X1
XFILL_0__2217_ gnd vdd FILL
XFILL_6__1985_ gnd vdd FILL
XFILL_0__3197_ gnd vdd FILL
XFILL_0__2148_ gnd vdd FILL
X_2776_ _2776_/A _2776_/B _2778_/B vdd gnd XOR2X1
XFILL_0__2079_ gnd vdd FILL
XFILL_1__2961_ gnd vdd FILL
X_1727_ _1891_/A _2123_/B _3147_/B vdd gnd NAND2X1
XFILL_6__2606_ gnd vdd FILL
XFILL_4__2670_ gnd vdd FILL
XFILL_3__2828_ gnd vdd FILL
XFILL_1__2892_ gnd vdd FILL
XFILL_6__3586_ gnd vdd FILL
XFILL_1__1912_ gnd vdd FILL
XFILL_1__1843_ gnd vdd FILL
XFILL_6__2537_ gnd vdd FILL
X_3328_ _3328_/D vdd _3347_/R _3573_/CLK _3328_/Q vdd gnd DFFSR
XFILL_6__2468_ gnd vdd FILL
XFILL_3__2759_ gnd vdd FILL
XFILL_7__3000_ gnd vdd FILL
XFILL_1__1774_ gnd vdd FILL
XFILL_1__3513_ gnd vdd FILL
X_3259_ _3259_/D vdd _3313_/R _3313_/CLK _3259_/Q vdd gnd DFFSR
XFILL_6__2399_ gnd vdd FILL
XFILL_4__3222_ gnd vdd FILL
XFILL_1__3444_ gnd vdd FILL
XFILL_1__3375_ gnd vdd FILL
XFILL_4__3153_ gnd vdd FILL
XFILL_4__2104_ gnd vdd FILL
XFILL_4__3084_ gnd vdd FILL
XFILL_4__2035_ gnd vdd FILL
XFILL_1__2326_ gnd vdd FILL
XFILL_1__2257_ gnd vdd FILL
XFILL_1__2188_ gnd vdd FILL
XFILL_7__2715_ gnd vdd FILL
XFILL_5__1730_ gnd vdd FILL
XFILL_4__2937_ gnd vdd FILL
XFILL_2__1952_ gnd vdd FILL
XFILL_7__2646_ gnd vdd FILL
XFILL_4__2868_ gnd vdd FILL
XFILL_5__3400_ gnd vdd FILL
XFILL_7__2577_ gnd vdd FILL
XFILL_4__2799_ gnd vdd FILL
XFILL_4__1819_ gnd vdd FILL
XFILL_2__1883_ gnd vdd FILL
XFILL_8__3040_ gnd vdd FILL
XFILL_2__3553_ gnd vdd FILL
XFILL_2__3484_ gnd vdd FILL
XFILL_5__2213_ gnd vdd FILL
XFILL_2__2504_ gnd vdd FILL
XFILL_7__3129_ gnd vdd FILL
XFILL_5__3193_ gnd vdd FILL
XFILL_2__2435_ gnd vdd FILL
XFILL_5__2144_ gnd vdd FILL
XFILL_5__2075_ gnd vdd FILL
XFILL_2__2366_ gnd vdd FILL
XFILL_0__3120_ gnd vdd FILL
XFILL_2__2297_ gnd vdd FILL
XFILL_5_BUFX2_insert25 gnd vdd FILL
XFILL_5_BUFX2_insert14 gnd vdd FILL
XFILL_5_BUFX2_insert58 gnd vdd FILL
XFILL_8__2824_ gnd vdd FILL
XFILL_5_BUFX2_insert47 gnd vdd FILL
XFILL_0__3051_ gnd vdd FILL
XFILL_8__2755_ gnd vdd FILL
XFILL_5_BUFX2_insert69 gnd vdd FILL
XFILL_0__2002_ gnd vdd FILL
XFILL_5__2977_ gnd vdd FILL
XFILL_6__1770_ gnd vdd FILL
XFILL_8__1706_ gnd vdd FILL
X_2630_ _2630_/A _2635_/A vdd gnd INVX1
XFILL_5__1928_ gnd vdd FILL
XFILL_3__1992_ gnd vdd FILL
XFILL_8__2686_ gnd vdd FILL
XFILL182250x163950 gnd vdd FILL
X_2561_ _2751_/A _2574_/B _2561_/C _3584_/A vdd gnd OAI21X1
XFILL_5__1859_ gnd vdd FILL
XFILL_6__3440_ gnd vdd FILL
X_2492_ _2508_/B _2511_/A _3575_/Q _2497_/A vdd gnd OAI21X1
XFILL_0__2904_ gnd vdd FILL
XFILL_6__3371_ gnd vdd FILL
XFILL_5__3529_ gnd vdd FILL
XFILL_6__2322_ gnd vdd FILL
XFILL_3__3593_ gnd vdd FILL
XFILL_3__2613_ gnd vdd FILL
XFILL_0__2835_ gnd vdd FILL
XFILL_9__2031_ gnd vdd FILL
XFILL_3__2544_ gnd vdd FILL
X_3113_ _3121_/A _3125_/B _3332_/Q _3114_/C vdd gnd OAI21X1
XFILL_6__2253_ gnd vdd FILL
XFILL_0__2766_ gnd vdd FILL
XFILL_8__3169_ gnd vdd FILL
X_3044_ _3044_/A _3131_/A vdd gnd INVX1
XFILL_3__2475_ gnd vdd FILL
XFILL_6__2184_ gnd vdd FILL
XFILL_0__1717_ gnd vdd FILL
XFILL_0__2697_ gnd vdd FILL
XFILL_1__3160_ gnd vdd FILL
XFILL_1__3091_ gnd vdd FILL
XFILL_3__3027_ gnd vdd FILL
XFILL_1__2111_ gnd vdd FILL
XFILL_1__2042_ gnd vdd FILL
XFILL_6__1968_ gnd vdd FILL
X_2828_ _2828_/A _2933_/C _2835_/A vdd gnd AND2X2
XFILL_7__2500_ gnd vdd FILL
XFILL_7__3480_ gnd vdd FILL
XFILL_6__1899_ gnd vdd FILL
XFILL_4__2722_ gnd vdd FILL
X_2759_ _2759_/A _2759_/B _3296_/D _2762_/A vdd gnd OAI21X1
XFILL_1__2944_ gnd vdd FILL
XFILL_7__2431_ gnd vdd FILL
XFILL_7__2362_ gnd vdd FILL
XFILL_4__2653_ gnd vdd FILL
XFILL_1__2875_ gnd vdd FILL
XFILL_4__2584_ gnd vdd FILL
XFILL_7__2293_ gnd vdd FILL
XFILL_1__1826_ gnd vdd FILL
XFILL_1__1757_ gnd vdd FILL
XFILL_4__3205_ gnd vdd FILL
XFILL_1__1688_ gnd vdd FILL
XFILL_4__3136_ gnd vdd FILL
XFILL_1__3427_ gnd vdd FILL
XFILL_2__2220_ gnd vdd FILL
XFILL_2__2151_ gnd vdd FILL
XFILL_1__2309_ gnd vdd FILL
XFILL_4__3067_ gnd vdd FILL
XFILL_2__2082_ gnd vdd FILL
XFILL_5__2900_ gnd vdd FILL
XFILL_4__2018_ gnd vdd FILL
XFILL_5__2831_ gnd vdd FILL
XFILL_8__2540_ gnd vdd FILL
XFILL_8__2471_ gnd vdd FILL
XFILL_5__2762_ gnd vdd FILL
XFILL_2__2984_ gnd vdd FILL
XFILL_5__2693_ gnd vdd FILL
XFILL_5__1713_ gnd vdd FILL
XFILL_7__2629_ gnd vdd FILL
XFILL_2__1935_ gnd vdd FILL
XFILL_2__1866_ gnd vdd FILL
XFILL_8__3023_ gnd vdd FILL
XFILL_2__3536_ gnd vdd FILL
XFILL_0__2620_ gnd vdd FILL
XFILL_2__1797_ gnd vdd FILL
XFILL_0__2551_ gnd vdd FILL
XFILL_2__3467_ gnd vdd FILL
XFILL_3__2260_ gnd vdd FILL
XBUFX2_insert8 RDY _2675_/A vdd gnd BUFX2
XFILL_5__3176_ gnd vdd FILL
XFILL_2__3398_ gnd vdd FILL
XFILL_3__2191_ gnd vdd FILL
XFILL_2__2418_ gnd vdd FILL
XFILL_0__2482_ gnd vdd FILL
XFILL_5__2127_ gnd vdd FILL
XFILL_2__2349_ gnd vdd FILL
XFILL_6__2940_ gnd vdd FILL
XFILL_5__2058_ gnd vdd FILL
XFILL_0__3103_ gnd vdd FILL
XFILL_6__2871_ gnd vdd FILL
X_1992_ _2199_/B _2786_/A _2338_/B vdd gnd OR2X2
XFILL_8__2807_ gnd vdd FILL
XFILL_0__3034_ gnd vdd FILL
XFILL_6__1822_ gnd vdd FILL
XFILL_8__2738_ gnd vdd FILL
X_3593_ _3593_/A AB[8] vdd gnd BUFX2
XFILL_6__1753_ gnd vdd FILL
X_2613_ _2685_/B _2671_/B vdd gnd INVX2
XFILL_8__2669_ gnd vdd FILL
XFILL_3__1975_ gnd vdd FILL
X_2544_ _3251_/Q _2744_/B vdd gnd INVX1
XFILL_6__3423_ gnd vdd FILL
X_2475_ _3205_/B _3587_/A vdd gnd INVX1
XFILL_1_BUFX2_insert23 gnd vdd FILL
XFILL_1_BUFX2_insert12 gnd vdd FILL
XFILL_1__2660_ gnd vdd FILL
XFILL_0__2818_ gnd vdd FILL
XFILL_6__2305_ gnd vdd FILL
XFILL_1_BUFX2_insert56 gnd vdd FILL
XFILL_1__2591_ gnd vdd FILL
XFILL_6_BUFX2_insert2 gnd vdd FILL
XFILL_1_BUFX2_insert45 gnd vdd FILL
XFILL_1_BUFX2_insert67 gnd vdd FILL
XFILL_1_BUFX2_insert78 gnd vdd FILL
XFILL_6__2236_ gnd vdd FILL
XFILL_3__2527_ gnd vdd FILL
XFILL_1_BUFX2_insert89 gnd vdd FILL
XFILL_3__2458_ gnd vdd FILL
XFILL_0__2749_ gnd vdd FILL
X_3027_ _3027_/A _3027_/B _3566_/A _3027_/Y vdd gnd OAI21X1
XFILL_6__2167_ gnd vdd FILL
XFILL_7__2980_ gnd vdd FILL
XFILL_3__2389_ gnd vdd FILL
XFILL_1__3212_ gnd vdd FILL
XFILL_6__2098_ gnd vdd FILL
XFILL_1_CLKBUF1_insert35 gnd vdd FILL
XFILL_1__3143_ gnd vdd FILL
XFILL_7__1931_ gnd vdd FILL
XFILL_7__1862_ gnd vdd FILL
XFILL_1__3074_ gnd vdd FILL
XFILL_7__3601_ gnd vdd FILL
XFILL_1__2025_ gnd vdd FILL
XFILL_7__1793_ gnd vdd FILL
XFILL_7__3532_ gnd vdd FILL
XFILL_7__3463_ gnd vdd FILL
XFILL_7__2414_ gnd vdd FILL
XFILL_4__2705_ gnd vdd FILL
XFILL_1__2927_ gnd vdd FILL
XFILL_7__3394_ gnd vdd FILL
XFILL_2__1720_ gnd vdd FILL
XFILL_4__2636_ gnd vdd FILL
XFILL_1__2858_ gnd vdd FILL
XFILL_7__2345_ gnd vdd FILL
XFILL_7__2276_ gnd vdd FILL
XFILL_1__1809_ gnd vdd FILL
XFILL_4__2567_ gnd vdd FILL
XFILL_1__2789_ gnd vdd FILL
XFILL_4__2498_ gnd vdd FILL
XFILL_5__3030_ gnd vdd FILL
XFILL_2__2203_ gnd vdd FILL
XFILL_8__1971_ gnd vdd FILL
XFILL_4__3119_ gnd vdd FILL
XFILL_2__3183_ gnd vdd FILL
XFILL_2__2134_ gnd vdd FILL
XFILL_2__2065_ gnd vdd FILL
XFILL_5__2814_ gnd vdd FILL
XFILL_8__2523_ gnd vdd FILL
XBUFX2_insert92 _3027_/Y _3115_/A vdd gnd BUFX2
XBUFX2_insert81 _1858_/Y _3147_/C vdd gnd BUFX2
XFILL_5__2745_ gnd vdd FILL
XBUFX2_insert70 _1765_/Y _2108_/A vdd gnd BUFX2
XFILL_3__1760_ gnd vdd FILL
XFILL_2__2967_ gnd vdd FILL
XFILL_8__2454_ gnd vdd FILL
XFILL_2__1918_ gnd vdd FILL
XFILL_8__2385_ gnd vdd FILL
XFILL_0__1982_ gnd vdd FILL
XFILL_5__2676_ gnd vdd FILL
XFILL_3__3430_ gnd vdd FILL
X_2260_ _2933_/B _2899_/A _2798_/B vdd gnd NAND2X1
XFILL_2__2898_ gnd vdd FILL
XFILL_3__1691_ gnd vdd FILL
XFILL_8_BUFX2_insert51 gnd vdd FILL
XFILL_8_BUFX2_insert40 gnd vdd FILL
XFILL_2__1849_ gnd vdd FILL
XFILL_8_BUFX2_insert84 gnd vdd FILL
XFILL_8_BUFX2_insert62 gnd vdd FILL
XFILL_8__3006_ gnd vdd FILL
X_2191_ _2191_/A _2196_/B vdd gnd INVX1
XFILL_8_BUFX2_insert73 gnd vdd FILL
XFILL_6__3070_ gnd vdd FILL
XFILL_0__2603_ gnd vdd FILL
XFILL_8_BUFX2_insert95 gnd vdd FILL
XFILL_6__2021_ gnd vdd FILL
XFILL_2__3519_ gnd vdd FILL
XFILL_3__2312_ gnd vdd FILL
XFILL_0__3583_ gnd vdd FILL
XFILL_5__3228_ gnd vdd FILL
XFILL_3__2243_ gnd vdd FILL
XFILL_0__2534_ gnd vdd FILL
XFILL_0__2465_ gnd vdd FILL
XFILL_5__3159_ gnd vdd FILL
XFILL_3__2174_ gnd vdd FILL
XFILL_6__2923_ gnd vdd FILL
XFILL_0__2396_ gnd vdd FILL
XFILL183750x150 gnd vdd FILL
X_1975_ _1986_/A _1975_/B _1975_/C _3404_/B vdd gnd OAI21X1
XFILL_6__2854_ gnd vdd FILL
XFILL_0__3017_ gnd vdd FILL
XFILL_6__2785_ gnd vdd FILL
XFILL_6__1805_ gnd vdd FILL
XFILL_6__1736_ gnd vdd FILL
XFILL_3__1958_ gnd vdd FILL
X_3576_ _3576_/D vdd _3578_/R _3576_/CLK _3576_/Q vdd gnd DFFSR
X_2527_ _2563_/A _3571_/Q _2527_/C _2528_/C vdd gnd AOI21X1
XFILL_4__3470_ gnd vdd FILL
XFILL_6__3406_ gnd vdd FILL
XFILL_3__1889_ gnd vdd FILL
X_2458_ _2508_/B _2511_/A _3570_/Q _2460_/A vdd gnd OAI21X1
XFILL_1__2712_ gnd vdd FILL
XFILL_4__2421_ gnd vdd FILL
XFILL_7__2130_ gnd vdd FILL
XFILL_3__3559_ gnd vdd FILL
XFILL_4__2352_ gnd vdd FILL
X_2389_ _3312_/Q _2425_/B _2390_/C vdd gnd NAND2X1
XFILL_1__2643_ gnd vdd FILL
XFILL_7__2061_ gnd vdd FILL
XFILL_1__2574_ gnd vdd FILL
XFILL_4__2283_ gnd vdd FILL
XFILL_6__2219_ gnd vdd FILL
XFILL_6__3199_ gnd vdd FILL
XFILL_7__2963_ gnd vdd FILL
XFILL_1__3126_ gnd vdd FILL
XFILL_7__2894_ gnd vdd FILL
XFILL_7__1914_ gnd vdd FILL
XFILL_1__3057_ gnd vdd FILL
XFILL_7__1845_ gnd vdd FILL
XFILL_1__2008_ gnd vdd FILL
XFILL_7__3515_ gnd vdd FILL
XFILL_7__1776_ gnd vdd FILL
XFILL_4__1998_ gnd vdd FILL
XFILL_2__2821_ gnd vdd FILL
XFILL_5__2530_ gnd vdd FILL
XFILL_7__3446_ gnd vdd FILL
XFILL_2__2752_ gnd vdd FILL
XFILL_7__3377_ gnd vdd FILL
XFILL_8__2170_ gnd vdd FILL
XFILL_2__1703_ gnd vdd FILL
XFILL_5__2461_ gnd vdd FILL
XFILL_7__2328_ gnd vdd FILL
XFILL_4__3599_ gnd vdd FILL
XFILL_5__2392_ gnd vdd FILL
XFILL_2__2683_ gnd vdd FILL
XFILL_4__2619_ gnd vdd FILL
XFILL_7__2259_ gnd vdd FILL
XFILL_5__3013_ gnd vdd FILL
XFILL_0__2250_ gnd vdd FILL
XCLKBUF1_insert37 clk _3307_/CLK vdd gnd CLKBUF1
XFILL_8__1954_ gnd vdd FILL
XFILL_2__3166_ gnd vdd FILL
XFILL_0__2181_ gnd vdd FILL
XFILL_2__2117_ gnd vdd FILL
XFILL_8__1885_ gnd vdd FILL
XFILL_2__3097_ gnd vdd FILL
X_1760_ _3007_/B _3280_/Q _3274_/Q _1771_/B vdd gnd AOI21X1
XFILL_3__2930_ gnd vdd FILL
XFILL_2__2048_ gnd vdd FILL
XFILL_3__2861_ gnd vdd FILL
XFILL_8__3555_ gnd vdd FILL
X_1691_ _3291_/Q _1693_/B vdd gnd INVX1
XFILL_8__3486_ gnd vdd FILL
X_3430_ _3485_/A _3431_/B vdd gnd INVX1
XFILL_8__2506_ gnd vdd FILL
XFILL_6__2570_ gnd vdd FILL
XFILL_3__1812_ gnd vdd FILL
XFILL_3__2792_ gnd vdd FILL
X_3361_ _3361_/D vdd _3363_/R _3363_/CLK _3361_/Q vdd gnd DFFSR
XFILL_5__2728_ gnd vdd FILL
XFILL_8__2437_ gnd vdd FILL
X_2312_ _2312_/A _2312_/B _2312_/C _2313_/B vdd gnd OAI21X1
XFILL_3__1743_ gnd vdd FILL
XFILL_5__2659_ gnd vdd FILL
XFILL_0__1965_ gnd vdd FILL
X_3292_ _3292_/D vdd _3355_/R _3578_/CLK _3292_/Q vdd gnd DFFSR
XFILL_8__2368_ gnd vdd FILL
XFILL_6__3122_ gnd vdd FILL
XFILL_3__3413_ gnd vdd FILL
X_2243_ _3022_/A _2968_/A _2341_/C _2244_/A vdd gnd OAI21X1
XFILL_8__2299_ gnd vdd FILL
XFILL_0__1896_ gnd vdd FILL
X_2174_ _2276_/A _3189_/A _3176_/B _2177_/A vdd gnd OAI21X1
XFILL_6__3053_ gnd vdd FILL
XFILL_0__3566_ gnd vdd FILL
XFILL184050x167850 gnd vdd FILL
XFILL_6__2004_ gnd vdd FILL
XFILL_0__2517_ gnd vdd FILL
XFILL_0__3497_ gnd vdd FILL
XFILL_3__2226_ gnd vdd FILL
XFILL_1__2290_ gnd vdd FILL
XFILL_3__2157_ gnd vdd FILL
XFILL_0__2448_ gnd vdd FILL
XFILL_0__2379_ gnd vdd FILL
XFILL_6__2906_ gnd vdd FILL
XFILL_4__2970_ gnd vdd FILL
XFILL_3__2088_ gnd vdd FILL
X_1958_ _3320_/Q _3029_/B _1959_/B vdd gnd NAND2X1
XFILL_6__2837_ gnd vdd FILL
XFILL_4_BUFX2_insert60 gnd vdd FILL
XFILL_4__1921_ gnd vdd FILL
XFILL_4_BUFX2_insert93 gnd vdd FILL
XFILL_4_BUFX2_insert82 gnd vdd FILL
X_1889_ _3237_/Q _3183_/B _3281_/Q _2960_/B _1898_/A vdd gnd OAI22X1
XFILL_4__1852_ gnd vdd FILL
XFILL_4_BUFX2_insert71 gnd vdd FILL
XFILL_9__2546_ gnd vdd FILL
XFILL_6__2768_ gnd vdd FILL
XFILL_6__1719_ gnd vdd FILL
XFILL_4__1783_ gnd vdd FILL
XFILL_6__2699_ gnd vdd FILL
X_3559_ _3576_/Q _3560_/A _3560_/C vdd gnd NAND2X1
XFILL_4__3522_ gnd vdd FILL
XFILL_7__3231_ gnd vdd FILL
XFILL184350x11850 gnd vdd FILL
XFILL_4__3453_ gnd vdd FILL
XFILL_4__2404_ gnd vdd FILL
XFILL_7__3162_ gnd vdd FILL
XFILL_7__3093_ gnd vdd FILL
XFILL_4__3384_ gnd vdd FILL
XFILL_7__2113_ gnd vdd FILL
XFILL_1__2626_ gnd vdd FILL
XFILL_7__2044_ gnd vdd FILL
XFILL_4__2335_ gnd vdd FILL
XFILL_4__2266_ gnd vdd FILL
XFILL_1__2557_ gnd vdd FILL
XFILL_1__2488_ gnd vdd FILL
XFILL_4__2197_ gnd vdd FILL
XFILL_2__3020_ gnd vdd FILL
XFILL_7__2946_ gnd vdd FILL
XFILL_1__3109_ gnd vdd FILL
XFILL_5__1961_ gnd vdd FILL
XFILL_7__2877_ gnd vdd FILL
XFILL_5__1892_ gnd vdd FILL
XFILL_7__1828_ gnd vdd FILL
XFILL_7__1759_ gnd vdd FILL
XFILL_2__2804_ gnd vdd FILL
XFILL_5__3562_ gnd vdd FILL
XFILL_5__3493_ gnd vdd FILL
XFILL_7__3429_ gnd vdd FILL
XFILL_8__2222_ gnd vdd FILL
XFILL_5__2513_ gnd vdd FILL
XFILL_2__2735_ gnd vdd FILL
XFILL_5__2444_ gnd vdd FILL
XFILL_8__2153_ gnd vdd FILL
XFILL_0__1750_ gnd vdd FILL
XFILL_2__2666_ gnd vdd FILL
XFILL_8__2084_ gnd vdd FILL
XFILL_5__2375_ gnd vdd FILL
XFILL_0__3420_ gnd vdd FILL
XFILL_2__2597_ gnd vdd FILL
XFILL_3__3060_ gnd vdd FILL
X_2930_ _2930_/A _2933_/A _2931_/C vdd gnd NOR2X1
XFILL_3__2011_ gnd vdd FILL
XFILL_0__2302_ gnd vdd FILL
XFILL_2__3218_ gnd vdd FILL
XFILL_8__2986_ gnd vdd FILL
XFILL_0__2233_ gnd vdd FILL
X_2861_ _2861_/A _2919_/B _2861_/C _2861_/D _3272_/D vdd gnd AOI22X1
XFILL_8__1937_ gnd vdd FILL
XFILL_2__3149_ gnd vdd FILL
XFILL_8__1868_ gnd vdd FILL
XFILL_0__2164_ gnd vdd FILL
X_2792_ _2992_/A _2898_/B _2792_/C _2821_/A _3260_/D vdd gnd OAI22X1
X_1812_ _3152_/C _3149_/C _2379_/A _1841_/B vdd gnd OAI21X1
XFILL_3__2913_ gnd vdd FILL
XFILL_8__1799_ gnd vdd FILL
XFILL_0__2095_ gnd vdd FILL
X_1743_ _3235_/Q _3236_/Q _2057_/A vdd gnd NAND2X1
XFILL_8__3538_ gnd vdd FILL
XFILL_6__2622_ gnd vdd FILL
XFILL_3__2844_ gnd vdd FILL
X_3413_ _3521_/A _3413_/B _3418_/C vdd gnd NAND2X1
XFILL_6__2553_ gnd vdd FILL
XFILL_8__3469_ gnd vdd FILL
XFILL_3__2775_ gnd vdd FILL
X_3344_ _3344_/D vdd _3345_/R _3577_/CLK _3344_/Q vdd gnd DFFSR
XFILL_0__2997_ gnd vdd FILL
XFILL_9__2193_ gnd vdd FILL
XFILL_6__2484_ gnd vdd FILL
XFILL_3__1726_ gnd vdd FILL
XFILL_1__1790_ gnd vdd FILL
X_3275_ _3275_/D vdd _3346_/R _3346_/CLK _3275_/Q vdd gnd DFFSR
XFILL_0__1948_ gnd vdd FILL
XFILL_1__3460_ gnd vdd FILL
X_2226_ _2327_/A _2226_/B _2296_/B vdd gnd AND2X2
XFILL_1_BUFX2_insert8 gnd vdd FILL
XFILL_6_CLKBUF1_insert35 gnd vdd FILL
XFILL_0__1879_ gnd vdd FILL
XFILL_6__3105_ gnd vdd FILL
XFILL_1__2411_ gnd vdd FILL
XFILL_1__3391_ gnd vdd FILL
XFILL_6__3036_ gnd vdd FILL
X_2157_ _2352_/A _2157_/B _2285_/B _2228_/B vdd gnd NAND3X1
XFILL_4__2120_ gnd vdd FILL
XFILL_0__3549_ gnd vdd FILL
X_2088_ _2212_/A _3145_/B _3144_/C vdd gnd NOR2X1
XFILL_4__2051_ gnd vdd FILL
XFILL_1__2342_ gnd vdd FILL
XFILL_1__2273_ gnd vdd FILL
XFILL_3__2209_ gnd vdd FILL
XFILL_7__2800_ gnd vdd FILL
XFILL_3__3189_ gnd vdd FILL
XFILL_7__2731_ gnd vdd FILL
XFILL_4__2953_ gnd vdd FILL
XFILL_4__1904_ gnd vdd FILL
XFILL_7__2662_ gnd vdd FILL
XFILL_4__2884_ gnd vdd FILL
XFILL_7__2593_ gnd vdd FILL
XFILL184350x23550 gnd vdd FILL
XFILL_4__1835_ gnd vdd FILL
XFILL_4__1766_ gnd vdd FILL
XFILL_9_BUFX2_insert39 gnd vdd FILL
XFILL_4__3505_ gnd vdd FILL
XFILL_1__1988_ gnd vdd FILL
XFILL_4__1697_ gnd vdd FILL
XFILL_7__3214_ gnd vdd FILL
XFILL_2__2520_ gnd vdd FILL
XFILL_4__3436_ gnd vdd FILL
XFILL_7__3145_ gnd vdd FILL
XFILL_5__2160_ gnd vdd FILL
XFILL_4__3367_ gnd vdd FILL
XFILL_2__2451_ gnd vdd FILL
XFILL_7__3076_ gnd vdd FILL
XFILL_4__2318_ gnd vdd FILL
XFILL_2__2382_ gnd vdd FILL
XFILL_1__3589_ gnd vdd FILL
XFILL_1__2609_ gnd vdd FILL
XFILL_0_BUFX2_insert91 gnd vdd FILL
XFILL_7__2027_ gnd vdd FILL
XFILL_0_BUFX2_insert80 gnd vdd FILL
XFILL_5__2091_ gnd vdd FILL
XFILL_8__2840_ gnd vdd FILL
XFILL_4__2249_ gnd vdd FILL
XFILL_2__3003_ gnd vdd FILL
XFILL_8__2771_ gnd vdd FILL
XFILL_7__2929_ gnd vdd FILL
XFILL_5__2993_ gnd vdd FILL
XFILL_8__1722_ gnd vdd FILL
XFILL_5__1944_ gnd vdd FILL
XFILL_5__1875_ gnd vdd FILL
XFILL_0__2920_ gnd vdd FILL
XFILL_5__3545_ gnd vdd FILL
XFILL_0__2851_ gnd vdd FILL
XFILL_3__2560_ gnd vdd FILL
XFILL_5__3476_ gnd vdd FILL
XFILL_8__2205_ gnd vdd FILL
XFILL_2__2718_ gnd vdd FILL
XFILL_0__2782_ gnd vdd FILL
XFILL_0__1802_ gnd vdd FILL
XFILL_8__3185_ gnd vdd FILL
X_3060_ _3293_/D _3088_/S _3060_/C _3060_/D _3135_/A vdd gnd OAI22X1
XFILL_5__2427_ gnd vdd FILL
XFILL_3__2491_ gnd vdd FILL
XFILL_8__2136_ gnd vdd FILL
XFILL_0__1733_ gnd vdd FILL
X_2011_ _2022_/A _2985_/A _2011_/C _2179_/A vdd gnd OAI21X1
XFILL_5__2358_ gnd vdd FILL
XFILL_2__2649_ gnd vdd FILL
XFILL_8__2067_ gnd vdd FILL
XFILL_3__3112_ gnd vdd FILL
XFILL_0__3403_ gnd vdd FILL
XFILL_5__2289_ gnd vdd FILL
XFILL_3__3043_ gnd vdd FILL
X_2913_ _2913_/A _2936_/B _2913_/C _2913_/D _3286_/D vdd gnd AOI22X1
XFILL_8__2969_ gnd vdd FILL
X_2844_ _2851_/A _2844_/B _2846_/C vdd gnd NAND2X1
XFILL_0__2216_ gnd vdd FILL
XFILL_6__1984_ gnd vdd FILL
XFILL_9__1693_ gnd vdd FILL
XFILL_0__3196_ gnd vdd FILL
XFILL_0__2147_ gnd vdd FILL
X_2775_ _2775_/A _2775_/B _2775_/C _2776_/A vdd gnd NAND3X1
XFILL_0__2078_ gnd vdd FILL
XFILL_1__2960_ gnd vdd FILL
X_1726_ _3234_/Q _3233_/Q _1891_/A vdd gnd NOR2X1
XFILL_6__2605_ gnd vdd FILL
XFILL_1__2891_ gnd vdd FILL
XFILL_3__2827_ gnd vdd FILL
XFILL_1__1911_ gnd vdd FILL
XFILL_6__3585_ gnd vdd FILL
XFILL_1__1842_ gnd vdd FILL
XFILL_6__2536_ gnd vdd FILL
X_3327_ _3327_/D vdd _3353_/R _3577_/CLK _3327_/Q vdd gnd DFFSR
XFILL_6__2467_ gnd vdd FILL
XFILL_3__2758_ gnd vdd FILL
XFILL_1__3512_ gnd vdd FILL
XFILL_3__1709_ gnd vdd FILL
XFILL_3__2689_ gnd vdd FILL
XFILL_1__1773_ gnd vdd FILL
X_3258_ _3258_/D vdd _3313_/R _3284_/CLK _3258_/Q vdd gnd DFFSR
XFILL_6__2398_ gnd vdd FILL
XFILL_4__3221_ gnd vdd FILL
XFILL_1__3443_ gnd vdd FILL
X_2209_ _2346_/A _2209_/B _2210_/A vdd gnd NOR2X1
XFILL_4__3152_ gnd vdd FILL
X_3189_ _3189_/A _3189_/B _3189_/C _3194_/B vdd gnd OAI21X1
XFILL_1__3374_ gnd vdd FILL
XFILL_4__2103_ gnd vdd FILL
XFILL_6__3019_ gnd vdd FILL
XFILL_4__3083_ gnd vdd FILL
XFILL_1__2325_ gnd vdd FILL
XFILL_4__2034_ gnd vdd FILL
XFILL_1__2256_ gnd vdd FILL
XFILL_1__2187_ gnd vdd FILL
XFILL184350x35250 gnd vdd FILL
XFILL_7__2714_ gnd vdd FILL
XFILL_4__2936_ gnd vdd FILL
XFILL_4__2867_ gnd vdd FILL
XFILL_2__1951_ gnd vdd FILL
XFILL_7__2645_ gnd vdd FILL
XFILL_7__2576_ gnd vdd FILL
XFILL_2__1882_ gnd vdd FILL
XFILL_4__1818_ gnd vdd FILL
XFILL_4__2798_ gnd vdd FILL
XFILL_4__1749_ gnd vdd FILL
XFILL_2__3552_ gnd vdd FILL
XFILL_2__3483_ gnd vdd FILL
XFILL_4__3419_ gnd vdd FILL
XFILL_2__2503_ gnd vdd FILL
XFILL_5__2212_ gnd vdd FILL
XFILL_7__3128_ gnd vdd FILL
XFILL_5__3192_ gnd vdd FILL
XFILL_2__2434_ gnd vdd FILL
XFILL_7__3059_ gnd vdd FILL
XFILL_5__2143_ gnd vdd FILL
XFILL_5__2074_ gnd vdd FILL
XFILL_2__2365_ gnd vdd FILL
XFILL_5_BUFX2_insert26 gnd vdd FILL
XFILL_2__2296_ gnd vdd FILL
XFILL_5_BUFX2_insert15 gnd vdd FILL
XFILL_5_BUFX2_insert59 gnd vdd FILL
XFILL_8__2823_ gnd vdd FILL
XFILL_5_BUFX2_insert48 gnd vdd FILL
XFILL_0__3050_ gnd vdd FILL
XFILL_8__2754_ gnd vdd FILL
XFILL_0__2001_ gnd vdd FILL
XFILL_5__2976_ gnd vdd FILL
XFILL_8__1705_ gnd vdd FILL
XFILL_5__1927_ gnd vdd FILL
XFILL_3__1991_ gnd vdd FILL
XFILL_8__2685_ gnd vdd FILL
X_2560_ _2560_/A _2561_/C vdd gnd INVX1
X_2491_ _3209_/B _3589_/A vdd gnd INVX1
XFILL_5__1858_ gnd vdd FILL
XFILL_0__2903_ gnd vdd FILL
XFILL_6__3370_ gnd vdd FILL
XFILL_3__2612_ gnd vdd FILL
XFILL_5__1789_ gnd vdd FILL
XFILL_0__2834_ gnd vdd FILL
XFILL_5__3528_ gnd vdd FILL
XFILL_6__2321_ gnd vdd FILL
XFILL_3__3592_ gnd vdd FILL
XFILL_5__3459_ gnd vdd FILL
XFILL_6__2252_ gnd vdd FILL
XFILL_3__2543_ gnd vdd FILL
X_3112_ _3129_/A _3126_/B _3112_/C _3331_/D vdd gnd OAI21X1
XFILL_3__2474_ gnd vdd FILL
XFILL_0__2765_ gnd vdd FILL
XFILL_8__3168_ gnd vdd FILL
XFILL_8__3099_ gnd vdd FILL
X_3043_ _3043_/A _3088_/S _3043_/C _3044_/A vdd gnd OAI21X1
XFILL_6__2183_ gnd vdd FILL
XFILL_8__2119_ gnd vdd FILL
XFILL_0__2696_ gnd vdd FILL
XFILL_0__1716_ gnd vdd FILL
XFILL_1__3090_ gnd vdd FILL
XFILL_3__3026_ gnd vdd FILL
XFILL_1__2110_ gnd vdd FILL
XFILL_1__2041_ gnd vdd FILL
XFILL_6__1967_ gnd vdd FILL
X_2827_ _2887_/B _2875_/A _2828_/A vdd gnd NOR2X1
XFILL_0__3179_ gnd vdd FILL
XFILL_6__1898_ gnd vdd FILL
XFILL_4__2721_ gnd vdd FILL
X_2758_ _2768_/B _2773_/B _2766_/A vdd gnd NOR2X1
XFILL_1__2943_ gnd vdd FILL
X_1709_ _3079_/A _3296_/D vdd gnd INVX1
XFILL_7__2430_ gnd vdd FILL
XFILL_7__2361_ gnd vdd FILL
X_2689_ _2706_/B _2689_/B _2696_/B vdd gnd NOR2X1
XFILL_4__2652_ gnd vdd FILL
XFILL_1__2874_ gnd vdd FILL
XFILL_4__2583_ gnd vdd FILL
XFILL_6__2519_ gnd vdd FILL
XFILL_6__3499_ gnd vdd FILL
XFILL_1__1825_ gnd vdd FILL
XFILL_7__2292_ gnd vdd FILL
XFILL_1__1756_ gnd vdd FILL
XFILL_4__3204_ gnd vdd FILL
XFILL_1__3426_ gnd vdd FILL
XFILL_4__3135_ gnd vdd FILL
XFILL_4__3066_ gnd vdd FILL
XFILL_2__2150_ gnd vdd FILL
XFILL_4__2017_ gnd vdd FILL
XFILL_2__2081_ gnd vdd FILL
XFILL_1__2308_ gnd vdd FILL
XFILL_1__2239_ gnd vdd FILL
XFILL_5__2830_ gnd vdd FILL
XFILL_5__2761_ gnd vdd FILL
XFILL_2__2983_ gnd vdd FILL
XFILL_8__2470_ gnd vdd FILL
XFILL_5__1712_ gnd vdd FILL
XFILL_4__2919_ gnd vdd FILL
XFILL_5__2692_ gnd vdd FILL
XFILL_2__1934_ gnd vdd FILL
XFILL_7__2628_ gnd vdd FILL
XFILL_2__1865_ gnd vdd FILL
XFILL_7__2559_ gnd vdd FILL
XFILL_2__1796_ gnd vdd FILL
XFILL_2__3535_ gnd vdd FILL
XFILL_8__3022_ gnd vdd FILL
XFILL_0__2550_ gnd vdd FILL
XFILL_2__3466_ gnd vdd FILL
XBUFX2_insert9 RDY _2278_/A vdd gnd BUFX2
XFILL_5__3175_ gnd vdd FILL
XFILL_2__3397_ gnd vdd FILL
XFILL_3__2190_ gnd vdd FILL
XFILL_2__2417_ gnd vdd FILL
XFILL_5__2126_ gnd vdd FILL
XFILL_0__2481_ gnd vdd FILL
XFILL_2__2348_ gnd vdd FILL
XFILL_5__2057_ gnd vdd FILL
XFILL_6__2870_ gnd vdd FILL
XFILL_0__3102_ gnd vdd FILL
XFILL_8__2806_ gnd vdd FILL
XFILL_2__2279_ gnd vdd FILL
X_1991_ _2242_/A _1991_/B _1991_/C _2066_/A _2331_/B vdd gnd AOI22X1
XFILL_0__3033_ gnd vdd FILL
XFILL_6__1821_ gnd vdd FILL
XFILL_8__2737_ gnd vdd FILL
XFILL183750x140550 gnd vdd FILL
XFILL_5__2959_ gnd vdd FILL
X_3592_ _3592_/A AB[7] vdd gnd BUFX2
XFILL_6__1752_ gnd vdd FILL
X_2612_ _3197_/C _2612_/B _2612_/C _2612_/D _3239_/D vdd gnd OAI22X1
XFILL_8__2668_ gnd vdd FILL
XFILL_3__1974_ gnd vdd FILL
X_2543_ _2734_/B _2574_/B _2543_/C _3582_/A vdd gnd OAI21X1
XFILL_6__3422_ gnd vdd FILL
XFILL_8__2599_ gnd vdd FILL
X_2474_ _2474_/A _2519_/C _2474_/C _3205_/B vdd gnd AOI21X1
XFILL_9__3062_ gnd vdd FILL
XFILL_6__2304_ gnd vdd FILL
XFILL_1_BUFX2_insert24 gnd vdd FILL
XFILL_1_BUFX2_insert13 gnd vdd FILL
XFILL_1_BUFX2_insert57 gnd vdd FILL
XFILL_0__2817_ gnd vdd FILL
XFILL_1_BUFX2_insert68 gnd vdd FILL
XFILL_1_BUFX2_insert46 gnd vdd FILL
XFILL_6_BUFX2_insert3 gnd vdd FILL
XFILL_1__2590_ gnd vdd FILL
XFILL_3__2526_ gnd vdd FILL
XFILL_1_BUFX2_insert79 gnd vdd FILL
XFILL_6__2235_ gnd vdd FILL
XFILL_0__2748_ gnd vdd FILL
XFILL_6__2166_ gnd vdd FILL
XFILL_3__2457_ gnd vdd FILL
X_3026_ _3026_/A _3027_/B vdd gnd INVX1
XFILL_3__2388_ gnd vdd FILL
XFILL_0__2679_ gnd vdd FILL
XFILL_1__3211_ gnd vdd FILL
XFILL_6__2097_ gnd vdd FILL
XFILL_1__3142_ gnd vdd FILL
XFILL_7__1930_ gnd vdd FILL
XFILL_1_CLKBUF1_insert36 gnd vdd FILL
XFILL_3__3009_ gnd vdd FILL
XFILL_1__3073_ gnd vdd FILL
XFILL_7__3600_ gnd vdd FILL
XFILL_7__1861_ gnd vdd FILL
XFILL_1__2024_ gnd vdd FILL
XFILL_6__2999_ gnd vdd FILL
XFILL_7__1792_ gnd vdd FILL
XFILL_7__3531_ gnd vdd FILL
XFILL_7__3462_ gnd vdd FILL
XFILL_4__2704_ gnd vdd FILL
XFILL_7__2413_ gnd vdd FILL
XFILL_1__2926_ gnd vdd FILL
XFILL_7__3393_ gnd vdd FILL
XFILL_4__2635_ gnd vdd FILL
XFILL_1__2857_ gnd vdd FILL
XFILL_7__2344_ gnd vdd FILL
XFILL_7__2275_ gnd vdd FILL
XFILL_1__1808_ gnd vdd FILL
XFILL_4__2566_ gnd vdd FILL
XFILL_1__2788_ gnd vdd FILL
XFILL_4__2497_ gnd vdd FILL
XFILL_1__1739_ gnd vdd FILL
XFILL_4__3118_ gnd vdd FILL
XFILL_1__3409_ gnd vdd FILL
XFILL_2__2202_ gnd vdd FILL
XFILL_2__3182_ gnd vdd FILL
XFILL_8__1970_ gnd vdd FILL
XFILL_2__2133_ gnd vdd FILL
XFILL_4__3049_ gnd vdd FILL
XFILL_2__2064_ gnd vdd FILL
XFILL_5__2813_ gnd vdd FILL
XBUFX2_insert60 _1993_/Y _2298_/D vdd gnd BUFX2
XFILL_8__2522_ gnd vdd FILL
XBUFX2_insert93 _3027_/Y _3121_/A vdd gnd BUFX2
XBUFX2_insert82 _1858_/Y _3006_/B vdd gnd BUFX2
XFILL_5__2744_ gnd vdd FILL
XBUFX2_insert71 _1765_/Y _2221_/A vdd gnd BUFX2
XFILL_2__2966_ gnd vdd FILL
XFILL_8__2453_ gnd vdd FILL
XFILL_5__2675_ gnd vdd FILL
XFILL_2__1917_ gnd vdd FILL
XFILL_2__2897_ gnd vdd FILL
XFILL_8__2384_ gnd vdd FILL
XFILL_3__1690_ gnd vdd FILL
XFILL_0__1981_ gnd vdd FILL
XFILL_2__1848_ gnd vdd FILL
X_2190_ _2786_/A _3192_/A _2821_/A _2190_/D _2336_/B vdd gnd OAI22X1
XFILL_8_BUFX2_insert41 gnd vdd FILL
XFILL_8_BUFX2_insert85 gnd vdd FILL
XFILL_8_BUFX2_insert63 gnd vdd FILL
XFILL_8_BUFX2_insert74 gnd vdd FILL
XFILL_8__3005_ gnd vdd FILL
XFILL_0__2602_ gnd vdd FILL
XFILL_8_BUFX2_insert52 gnd vdd FILL
XFILL_2__1779_ gnd vdd FILL
XFILL_8_BUFX2_insert96 gnd vdd FILL
XFILL_6__2020_ gnd vdd FILL
XFILL_2__3518_ gnd vdd FILL
XFILL_3__2311_ gnd vdd FILL
XFILL_0__3582_ gnd vdd FILL
XFILL_5__3227_ gnd vdd FILL
XFILL_2__3449_ gnd vdd FILL
XFILL_3__2242_ gnd vdd FILL
XFILL_0__2533_ gnd vdd FILL
XFILL_0__2464_ gnd vdd FILL
XFILL_5__3158_ gnd vdd FILL
XFILL_5__3089_ gnd vdd FILL
XFILL_3__2173_ gnd vdd FILL
XFILL_5__2109_ gnd vdd FILL
XFILL_6__2922_ gnd vdd FILL
XFILL_0__2395_ gnd vdd FILL
X_1974_ _1985_/A _3576_/Q _1974_/C _1975_/C vdd gnd AOI21X1
XFILL_6__2853_ gnd vdd FILL
XFILL_6__2784_ gnd vdd FILL
XFILL_0__3016_ gnd vdd FILL
XFILL_6__1804_ gnd vdd FILL
XFILL_6__1735_ gnd vdd FILL
XFILL_3__1957_ gnd vdd FILL
X_3575_ _3575_/D vdd _3578_/R _3576_/CLK _3575_/Q vdd gnd DFFSR
X_2526_ _2538_/B _2572_/B vdd gnd INVX2
XFILL_6__3405_ gnd vdd FILL
XFILL_4__2420_ gnd vdd FILL
X_2457_ _2457_/A _2457_/B _2574_/B vdd gnd NAND2X1
XFILL_3__1888_ gnd vdd FILL
XFILL_1__2711_ gnd vdd FILL
XFILL_1__2642_ gnd vdd FILL
XFILL_3__3558_ gnd vdd FILL
XFILL_4__2351_ gnd vdd FILL
X_2388_ _2872_/B _3077_/C _3248_/Q _2392_/A vdd gnd OAI21X1
XFILL_7__2060_ gnd vdd FILL
XFILL_3__3489_ gnd vdd FILL
XFILL_4__2282_ gnd vdd FILL
XFILL_3__2509_ gnd vdd FILL
XFILL_1__2573_ gnd vdd FILL
XFILL_6__2218_ gnd vdd FILL
XFILL_6__3198_ gnd vdd FILL
X_3009_ _3009_/A _3013_/C _3010_/B vdd gnd NAND2X1
XFILL_6__2149_ gnd vdd FILL
XFILL_7__2962_ gnd vdd FILL
XFILL_1__3125_ gnd vdd FILL
XFILL_7__2893_ gnd vdd FILL
XFILL_7__1913_ gnd vdd FILL
XFILL_1__3056_ gnd vdd FILL
XFILL_7__1844_ gnd vdd FILL
XFILL_1__2007_ gnd vdd FILL
XFILL_7__3514_ gnd vdd FILL
XFILL_7__1775_ gnd vdd FILL
XFILL_4__1997_ gnd vdd FILL
XFILL_2__2820_ gnd vdd FILL
XFILL_7__3445_ gnd vdd FILL
XFILL_2__2751_ gnd vdd FILL
XFILL_1__2909_ gnd vdd FILL
XFILL_7__3376_ gnd vdd FILL
XFILL_2__1702_ gnd vdd FILL
XFILL_5__2460_ gnd vdd FILL
XFILL_7__2327_ gnd vdd FILL
XFILL_4__3598_ gnd vdd FILL
XFILL_5__2391_ gnd vdd FILL
XFILL_2__2682_ gnd vdd FILL
XFILL_4__2618_ gnd vdd FILL
XFILL_4__2549_ gnd vdd FILL
XFILL_7__2258_ gnd vdd FILL
XFILL_7__2189_ gnd vdd FILL
XFILL_5__3012_ gnd vdd FILL
XCLKBUF1_insert38 clk _3577_/CLK vdd gnd CLKBUF1
XFILL_8__1953_ gnd vdd FILL
XFILL_2__3165_ gnd vdd FILL
XFILL_0__2180_ gnd vdd FILL
XFILL_2__3096_ gnd vdd FILL
XFILL_2__2116_ gnd vdd FILL
XFILL_8__1884_ gnd vdd FILL
XFILL_2__2047_ gnd vdd FILL
XFILL_3__2860_ gnd vdd FILL
XFILL_8__3554_ gnd vdd FILL
X_1690_ _2675_/A _1690_/B _1690_/C _3290_/D vdd gnd OAI21X1
XFILL_8__3485_ gnd vdd FILL
XFILL_3__2791_ gnd vdd FILL
XFILL_8__2505_ gnd vdd FILL
XFILL_3__1811_ gnd vdd FILL
XFILL_3__1742_ gnd vdd FILL
X_3360_ _3360_/D vdd _3363_/R _3363_/CLK _3360_/Q vdd gnd DFFSR
XFILL_5__2727_ gnd vdd FILL
XFILL_8__2436_ gnd vdd FILL
XFILL_2__2949_ gnd vdd FILL
X_2311_ _2311_/A _2312_/B vdd gnd INVX1
XFILL_0__1964_ gnd vdd FILL
XFILL_5__2658_ gnd vdd FILL
XFILL_8__2367_ gnd vdd FILL
X_3291_ _3291_/D vdd _3291_/R _3355_/CLK _3291_/Q vdd gnd DFFSR
XFILL_5__2589_ gnd vdd FILL
XFILL_6__3121_ gnd vdd FILL
XFILL_3__3412_ gnd vdd FILL
XFILL_8__2298_ gnd vdd FILL
X_2242_ _2242_/A _2242_/B _2242_/C _2341_/C vdd gnd OAI21X1
XFILL_0__1895_ gnd vdd FILL
X_2173_ _2339_/C _2335_/B _2323_/A vdd gnd NAND2X1
XFILL_6__3052_ gnd vdd FILL
XFILL_0__3565_ gnd vdd FILL
XFILL_6__2003_ gnd vdd FILL
XFILL_0__2516_ gnd vdd FILL
XFILL_0__3496_ gnd vdd FILL
XFILL_3__2225_ gnd vdd FILL
XFILL_3__2156_ gnd vdd FILL
XFILL_0__2447_ gnd vdd FILL
XFILL_0__2378_ gnd vdd FILL
XFILL_6__2905_ gnd vdd FILL
XFILL_3__2087_ gnd vdd FILL
XFILL_6__2836_ gnd vdd FILL
X_1957_ _3336_/Q _3110_/A _3127_/B _3345_/Q _1959_/C vdd gnd AOI22X1
XFILL_4_BUFX2_insert50 gnd vdd FILL
XFILL_4__1920_ gnd vdd FILL
XFILL_4_BUFX2_insert61 gnd vdd FILL
XFILL_4_BUFX2_insert94 gnd vdd FILL
XFILL_4_BUFX2_insert83 gnd vdd FILL
X_1888_ _1888_/A _1888_/B _3183_/B vdd gnd NAND2X1
XFILL_4__1851_ gnd vdd FILL
XFILL_4_BUFX2_insert72 gnd vdd FILL
XFILL_6__2767_ gnd vdd FILL
XFILL_3__2989_ gnd vdd FILL
X_3558_ _3560_/A _3558_/B _3558_/C _3575_/D vdd gnd OAI21X1
XFILL_6__1718_ gnd vdd FILL
XFILL_6__2698_ gnd vdd FILL
XFILL_4__1782_ gnd vdd FILL
XFILL_4__3521_ gnd vdd FILL
X_2509_ _3355_/Q _2669_/A vdd gnd INVX1
XFILL_7__3230_ gnd vdd FILL
X_3489_ _3493_/B _3491_/B vdd gnd INVX1
XFILL_4__3452_ gnd vdd FILL
XFILL_7__3161_ gnd vdd FILL
XFILL_4__3383_ gnd vdd FILL
XFILL_4__2403_ gnd vdd FILL
XFILL_7__2112_ gnd vdd FILL
XFILL_7__3092_ gnd vdd FILL
XFILL_4__2334_ gnd vdd FILL
XFILL_1__2625_ gnd vdd FILL
XFILL_7__2043_ gnd vdd FILL
XFILL_1__2556_ gnd vdd FILL
XFILL_4__2265_ gnd vdd FILL
XFILL_4__2196_ gnd vdd FILL
XFILL_1__2487_ gnd vdd FILL
XFILL_7__2945_ gnd vdd FILL
XFILL_1__3108_ gnd vdd FILL
XFILL_5__1960_ gnd vdd FILL
XFILL_7__2876_ gnd vdd FILL
XFILL_5__1891_ gnd vdd FILL
XFILL_1__3039_ gnd vdd FILL
XFILL_7__1827_ gnd vdd FILL
XFILL_7__1758_ gnd vdd FILL
XFILL_2__2803_ gnd vdd FILL
XFILL_5__3561_ gnd vdd FILL
XFILL_5__3492_ gnd vdd FILL
XFILL_7__3428_ gnd vdd FILL
XFILL_7__1689_ gnd vdd FILL
XFILL_8__2221_ gnd vdd FILL
XFILL_5__2512_ gnd vdd FILL
XFILL_2__2734_ gnd vdd FILL
XFILL_5__2443_ gnd vdd FILL
XFILL_8__2152_ gnd vdd FILL
XFILL_2__2665_ gnd vdd FILL
XFILL_8__2083_ gnd vdd FILL
XFILL_5__2374_ gnd vdd FILL
XFILL_2__2596_ gnd vdd FILL
XFILL_0__2301_ gnd vdd FILL
XFILL_3__2010_ gnd vdd FILL
XFILL_8__2985_ gnd vdd FILL
XFILL_2__3217_ gnd vdd FILL
X_2860_ _2860_/A _2866_/C _2861_/D vdd gnd AND2X2
XFILL_8__1936_ gnd vdd FILL
XFILL_2__3148_ gnd vdd FILL
XFILL_0__2232_ gnd vdd FILL
XFILL_0__2163_ gnd vdd FILL
X_1811_ _2435_/A _2289_/B _3174_/A vdd gnd OR2X2
XFILL_8__1867_ gnd vdd FILL
X_2791_ _3260_/Q _2992_/A vdd gnd INVX1
XFILL_2__3079_ gnd vdd FILL
XFILL_3__2912_ gnd vdd FILL
X_1742_ _2430_/A _2446_/B _2167_/A _1750_/B vdd gnd OAI21X1
XFILL_8__1798_ gnd vdd FILL
XFILL_0__2094_ gnd vdd FILL
XFILL_8__3537_ gnd vdd FILL
XFILL_6__2621_ gnd vdd FILL
XFILL_3__2843_ gnd vdd FILL
X_3412_ _3509_/C _3511_/A _3535_/A vdd gnd NAND2X1
XFILL_6__2552_ gnd vdd FILL
XFILL_8__3468_ gnd vdd FILL
XFILL_6__2483_ gnd vdd FILL
XFILL_3__2774_ gnd vdd FILL
X_3343_ _3343_/D vdd _3347_/R _3573_/CLK _3343_/Q vdd gnd DFFSR
XFILL_8__3399_ gnd vdd FILL
XFILL_0__2996_ gnd vdd FILL
XFILL_8__2419_ gnd vdd FILL
XFILL_3__1725_ gnd vdd FILL
XFILL_0__1947_ gnd vdd FILL
X_3274_ _3274_/D vdd _3282_/R _3284_/CLK _3274_/Q vdd gnd DFFSR
XFILL_0__1878_ gnd vdd FILL
XFILL_1_BUFX2_insert9 gnd vdd FILL
X_2225_ _2247_/B _2797_/B _2225_/C _2226_/B vdd gnd AOI21X1
XFILL_6__3104_ gnd vdd FILL
XFILL_6_CLKBUF1_insert36 gnd vdd FILL
XFILL_1__2410_ gnd vdd FILL
XFILL_1__3390_ gnd vdd FILL
XFILL_6__3035_ gnd vdd FILL
X_2156_ _2156_/A _2319_/B _2157_/B vdd gnd NOR2X1
XFILL_0__3548_ gnd vdd FILL
X_2087_ _2298_/A _3163_/A _2087_/C _2284_/A vdd gnd AOI21X1
XFILL_1__2341_ gnd vdd FILL
XFILL_4__2050_ gnd vdd FILL
XFILL_0__3479_ gnd vdd FILL
XFILL_1__2272_ gnd vdd FILL
XFILL_3__2208_ gnd vdd FILL
XFILL_3__3188_ gnd vdd FILL
XFILL_3__2139_ gnd vdd FILL
XFILL_7__2730_ gnd vdd FILL
XFILL_4__2952_ gnd vdd FILL
X_2989_ _3276_/Q _3023_/B _2990_/C vdd gnd NOR2X1
XFILL_4__1903_ gnd vdd FILL
XFILL_7__2661_ gnd vdd FILL
XFILL_6__2819_ gnd vdd FILL
XFILL_4__2883_ gnd vdd FILL
XFILL_7__2592_ gnd vdd FILL
XFILL_4__1834_ gnd vdd FILL
XFILL_4__1765_ gnd vdd FILL
XFILL_4__3504_ gnd vdd FILL
XFILL_1__1987_ gnd vdd FILL
XFILL_4__1696_ gnd vdd FILL
XFILL_7__3213_ gnd vdd FILL
XFILL_4__3435_ gnd vdd FILL
XFILL_2__2450_ gnd vdd FILL
XFILL_7__3144_ gnd vdd FILL
XFILL_4__3366_ gnd vdd FILL
XFILL_7__3075_ gnd vdd FILL
XFILL_4__2317_ gnd vdd FILL
XFILL_2__2381_ gnd vdd FILL
XFILL_5__2090_ gnd vdd FILL
XFILL_1__3588_ gnd vdd FILL
XFILL_1__2608_ gnd vdd FILL
XFILL_4__2248_ gnd vdd FILL
XFILL_7__2026_ gnd vdd FILL
XFILL_0_BUFX2_insert92 gnd vdd FILL
XFILL_0_BUFX2_insert81 gnd vdd FILL
XFILL_1__2539_ gnd vdd FILL
XFILL_0_BUFX2_insert70 gnd vdd FILL
XFILL_4__2179_ gnd vdd FILL
XFILL_2__3002_ gnd vdd FILL
XFILL_8__2770_ gnd vdd FILL
XFILL_7__2928_ gnd vdd FILL
XFILL_5__2992_ gnd vdd FILL
XFILL_8__1721_ gnd vdd FILL
XFILL_7__2859_ gnd vdd FILL
XFILL_5__1943_ gnd vdd FILL
XFILL_5__1874_ gnd vdd FILL
XFILL_5__3544_ gnd vdd FILL
XFILL_0__2850_ gnd vdd FILL
XFILL_5__3475_ gnd vdd FILL
XFILL_8__2204_ gnd vdd FILL
XFILL_0__2781_ gnd vdd FILL
XFILL_0__1801_ gnd vdd FILL
XFILL_8__3184_ gnd vdd FILL
XFILL_2__2717_ gnd vdd FILL
XFILL_5__2426_ gnd vdd FILL
XFILL_3__2490_ gnd vdd FILL
XFILL_8__2135_ gnd vdd FILL
XFILL_0__1732_ gnd vdd FILL
X_2010_ _2022_/A _3301_/Q _2011_/C vdd gnd NAND2X1
XFILL_2__2648_ gnd vdd FILL
XFILL_5__2357_ gnd vdd FILL
XFILL_2__2579_ gnd vdd FILL
XFILL_0__3402_ gnd vdd FILL
XFILL_8__2066_ gnd vdd FILL
XFILL_3__3111_ gnd vdd FILL
XFILL_5__2288_ gnd vdd FILL
XFILL_3__3042_ gnd vdd FILL
X_2912_ _2935_/A _2912_/B _2913_/D vdd gnd NOR2X1
XFILL_0__2215_ gnd vdd FILL
XFILL_8__2968_ gnd vdd FILL
X_2843_ _2933_/A _2895_/A _2843_/C _2844_/B vdd gnd OAI21X1
XFILL_8__2899_ gnd vdd FILL
XFILL_8__1919_ gnd vdd FILL
XFILL_0__3195_ gnd vdd FILL
XFILL_6__1983_ gnd vdd FILL
XFILL_0__2146_ gnd vdd FILL
X_2774_ _2774_/A _2775_/B vdd gnd INVX1
XFILL_0__2077_ gnd vdd FILL
X_1725_ _1725_/A _2279_/A vdd gnd INVX1
XFILL_6__2604_ gnd vdd FILL
XFILL_1__1910_ gnd vdd FILL
XFILL_1__2890_ gnd vdd FILL
XFILL_3__2826_ gnd vdd FILL
XFILL_6__3584_ gnd vdd FILL
XFILL_6__2535_ gnd vdd FILL
XFILL_1__1841_ gnd vdd FILL
X_3326_ _3326_/D vdd _3345_/R _3576_/CLK _3326_/Q vdd gnd DFFSR
XFILL_1__1772_ gnd vdd FILL
XFILL_6__2466_ gnd vdd FILL
XFILL_3__2757_ gnd vdd FILL
XFILL_1__3511_ gnd vdd FILL
XFILL_0__2979_ gnd vdd FILL
XFILL_3__1708_ gnd vdd FILL
XFILL_3__2688_ gnd vdd FILL
X_3257_ _3257_/D vdd _3282_/R _3284_/CLK _3257_/Q vdd gnd DFFSR
XFILL_6__2397_ gnd vdd FILL
XFILL_4__3220_ gnd vdd FILL
XFILL_1__3442_ gnd vdd FILL
X_2208_ _2786_/A _2700_/B _2208_/C _2235_/C _2209_/B vdd gnd OAI22X1
XFILL_4__3151_ gnd vdd FILL
X_3188_ _3188_/A _3191_/A vdd gnd INVX1
XFILL_1__3373_ gnd vdd FILL
X_2139_ _2212_/A _2448_/B _2342_/A _2140_/C vdd gnd OAI21X1
XFILL_4__2102_ gnd vdd FILL
XFILL_4__3082_ gnd vdd FILL
XFILL_6__3018_ gnd vdd FILL
XFILL_1__2324_ gnd vdd FILL
XFILL_4__2033_ gnd vdd FILL
XFILL184650x19650 gnd vdd FILL
XFILL_1__2255_ gnd vdd FILL
XFILL_1__2186_ gnd vdd FILL
XFILL_7__2713_ gnd vdd FILL
XFILL_4__2935_ gnd vdd FILL
XFILL_7__2644_ gnd vdd FILL
XFILL_4__2866_ gnd vdd FILL
XFILL_2__1950_ gnd vdd FILL
XFILL_2__1881_ gnd vdd FILL
XFILL_7__2575_ gnd vdd FILL
XFILL_4__1817_ gnd vdd FILL
XFILL_4__2797_ gnd vdd FILL
XFILL_4__1748_ gnd vdd FILL
XFILL_2__3551_ gnd vdd FILL
XFILL_2__3482_ gnd vdd FILL
XFILL_4__3418_ gnd vdd FILL
XFILL_5__2211_ gnd vdd FILL
XFILL_2__2502_ gnd vdd FILL
XFILL_5__3191_ gnd vdd FILL
XFILL_7__3127_ gnd vdd FILL
XFILL_5__2142_ gnd vdd FILL
XFILL_2__2433_ gnd vdd FILL
XFILL_7__3058_ gnd vdd FILL
XFILL_2__2364_ gnd vdd FILL
XFILL_5__2073_ gnd vdd FILL
XFILL_7__2009_ gnd vdd FILL
XFILL_2__2295_ gnd vdd FILL
XFILL_5_BUFX2_insert16 gnd vdd FILL
XFILL_5_BUFX2_insert49 gnd vdd FILL
XFILL_8__2822_ gnd vdd FILL
XFILL_5_BUFX2_insert27 gnd vdd FILL
XFILL_8__2753_ gnd vdd FILL
XFILL_0__2000_ gnd vdd FILL
XFILL_5__2975_ gnd vdd FILL
XFILL_8__1704_ gnd vdd FILL
XFILL_5__1926_ gnd vdd FILL
XFILL_3__1990_ gnd vdd FILL
XFILL_8__2684_ gnd vdd FILL
XFILL_5__1857_ gnd vdd FILL
X_2490_ _2490_/A _2519_/C _2490_/C _3209_/B vdd gnd AOI21X1
XFILL_0__2902_ gnd vdd FILL
XFILL_3__2611_ gnd vdd FILL
XFILL_5__1788_ gnd vdd FILL
XFILL_5__3527_ gnd vdd FILL
XFILL_0__2833_ gnd vdd FILL
XFILL_3__3591_ gnd vdd FILL
XFILL_6__2320_ gnd vdd FILL
X_3111_ _3111_/A _3125_/B _3331_/Q _3112_/C vdd gnd OAI21X1
XFILL_5__3458_ gnd vdd FILL
XFILL_6__2251_ gnd vdd FILL
XFILL_3__2542_ gnd vdd FILL
XFILL_3__2473_ gnd vdd FILL
XFILL_0__2764_ gnd vdd FILL
XFILL_8__3167_ gnd vdd FILL
XFILL_5__2409_ gnd vdd FILL
XFILL_8__3098_ gnd vdd FILL
XFILL_5__3389_ gnd vdd FILL
XFILL_6__2182_ gnd vdd FILL
X_3042_ _3571_/Q _3042_/B _3042_/C _3043_/C vdd gnd OAI21X1
XFILL_8__2118_ gnd vdd FILL
XFILL_0__2695_ gnd vdd FILL
XFILL_0__1715_ gnd vdd FILL
XFILL183150x163950 gnd vdd FILL
XFILL_8__2049_ gnd vdd FILL
XFILL_3__3025_ gnd vdd FILL
XFILL_1__2040_ gnd vdd FILL
XFILL_6__1966_ gnd vdd FILL
X_2826_ _2960_/A _2885_/B _2826_/C _3269_/D vdd gnd AOI21X1
XFILL_0__3178_ gnd vdd FILL
XFILL_0__2129_ gnd vdd FILL
XFILL_6__1897_ gnd vdd FILL
XFILL_4__2720_ gnd vdd FILL
X_2757_ _2757_/A _2757_/B _2757_/C _2757_/D _2775_/A vdd gnd AOI22X1
XFILL_1__2942_ gnd vdd FILL
X_1708_ _2768_/A DI[6] _1708_/C _3079_/A vdd gnd OAI21X1
X_2688_ _2741_/C _2741_/B _2689_/B vdd gnd OR2X2
XFILL_7__2360_ gnd vdd FILL
XFILL_4__2651_ gnd vdd FILL
XFILL_3__2809_ gnd vdd FILL
XFILL_1__2873_ gnd vdd FILL
XFILL_6__2518_ gnd vdd FILL
XFILL_4__2582_ gnd vdd FILL
XFILL_6__3498_ gnd vdd FILL
XFILL_1__1824_ gnd vdd FILL
XFILL_7__2291_ gnd vdd FILL
XFILL_1__1755_ gnd vdd FILL
X_3309_ _3309_/D vdd _3353_/R _3313_/CLK _3309_/Q vdd gnd DFFSR
XFILL_6__2449_ gnd vdd FILL
XFILL_4__3203_ gnd vdd FILL
XFILL_1__3425_ gnd vdd FILL
XFILL_4__3134_ gnd vdd FILL
XFILL_4__3065_ gnd vdd FILL
XFILL_2__2080_ gnd vdd FILL
XFILL_4__2016_ gnd vdd FILL
XFILL_1__2307_ gnd vdd FILL
XFILL_1__2238_ gnd vdd FILL
XFILL_1__2169_ gnd vdd FILL
XFILL_5__2760_ gnd vdd FILL
XFILL_4__2918_ gnd vdd FILL
XFILL_2__2982_ gnd vdd FILL
XFILL_5__1711_ gnd vdd FILL
XFILL_3_BUFX2_insert0 gnd vdd FILL
XFILL_5__2691_ gnd vdd FILL
XFILL_2__1933_ gnd vdd FILL
XFILL_7__2627_ gnd vdd FILL
XFILL_4__2849_ gnd vdd FILL
XFILL_7__2558_ gnd vdd FILL
XFILL_2__1864_ gnd vdd FILL
XFILL_7__2489_ gnd vdd FILL
XFILL_2__3603_ gnd vdd FILL
XFILL_2__1795_ gnd vdd FILL
XFILL_2__3534_ gnd vdd FILL
XFILL_8__3021_ gnd vdd FILL
XFILL_2__3465_ gnd vdd FILL
XFILL_5__3174_ gnd vdd FILL
XFILL_0__2480_ gnd vdd FILL
XFILL_2__3396_ gnd vdd FILL
XFILL_2__2416_ gnd vdd FILL
XFILL_5__2125_ gnd vdd FILL
XFILL_2__2347_ gnd vdd FILL
X_1990_ _2063_/B _3022_/A _1991_/C vdd gnd AND2X2
XFILL_5__2056_ gnd vdd FILL
XFILL_2__2278_ gnd vdd FILL
XFILL_8__2805_ gnd vdd FILL
XFILL_0__3101_ gnd vdd FILL
XFILL_0__3032_ gnd vdd FILL
XFILL_6__1820_ gnd vdd FILL
XFILL_8__2736_ gnd vdd FILL
X_3591_ _3591_/A AB[6] vdd gnd BUFX2
XFILL_5__2958_ gnd vdd FILL
XFILL_6__1751_ gnd vdd FILL
X_2611_ _3197_/C _2611_/B _2612_/D vdd gnd NAND2X1
XFILL_8__2667_ gnd vdd FILL
XFILL_5__2889_ gnd vdd FILL
XFILL_3__1973_ gnd vdd FILL
X_2542_ _2542_/A _2543_/C vdd gnd INVX1
XFILL_5__1909_ gnd vdd FILL
XFILL_6__3421_ gnd vdd FILL
XFILL_8__2598_ gnd vdd FILL
X_2473_ _2627_/A _2574_/B _2473_/C _2474_/C vdd gnd OAI21X1
XFILL183150x175650 gnd vdd FILL
XFILL183450x167850 gnd vdd FILL
XFILL_6__2303_ gnd vdd FILL
XFILL_1_BUFX2_insert25 gnd vdd FILL
XFILL_1_BUFX2_insert14 gnd vdd FILL
XFILL_1_BUFX2_insert58 gnd vdd FILL
XFILL_0__2816_ gnd vdd FILL
XFILL_3__2525_ gnd vdd FILL
XFILL_8__3219_ gnd vdd FILL
XFILL_1_BUFX2_insert47 gnd vdd FILL
XFILL_6_BUFX2_insert4 gnd vdd FILL
XFILL_6__2234_ gnd vdd FILL
XFILL_0__2747_ gnd vdd FILL
XFILL_1_BUFX2_insert69 gnd vdd FILL
XFILL_6__2165_ gnd vdd FILL
X_3025_ _3025_/A _3025_/B _3026_/A vdd gnd NOR2X1
XFILL_3__2456_ gnd vdd FILL
XFILL_3__2387_ gnd vdd FILL
XFILL_1__3210_ gnd vdd FILL
XFILL_0__2678_ gnd vdd FILL
XFILL_9__2914_ gnd vdd FILL
XFILL_6__2096_ gnd vdd FILL
XFILL_1_CLKBUF1_insert37 gnd vdd FILL
XFILL_1__3141_ gnd vdd FILL
XFILL_7__1860_ gnd vdd FILL
XFILL_1__3072_ gnd vdd FILL
XFILL_1__2023_ gnd vdd FILL
XFILL_3__3008_ gnd vdd FILL
XFILL_6__2998_ gnd vdd FILL
XFILL_7__1791_ gnd vdd FILL
XFILL_7__3530_ gnd vdd FILL
XFILL_6__1949_ gnd vdd FILL
X_2809_ _2973_/A _2887_/A _2809_/C _2815_/B _3265_/D vdd gnd OAI22X1
XFILL_7__3461_ gnd vdd FILL
XFILL_7__2412_ gnd vdd FILL
XFILL_4__2703_ gnd vdd FILL
XFILL_1__2925_ gnd vdd FILL
XFILL_7__3392_ gnd vdd FILL
XFILL_4__2634_ gnd vdd FILL
XFILL_1__2856_ gnd vdd FILL
XFILL_7__2343_ gnd vdd FILL
XFILL_7__2274_ gnd vdd FILL
XFILL_1__1807_ gnd vdd FILL
XFILL_4__2565_ gnd vdd FILL
XFILL_1__2787_ gnd vdd FILL
XFILL_4__2496_ gnd vdd FILL
XFILL_1__1738_ gnd vdd FILL
XFILL_4__3117_ gnd vdd FILL
XFILL_1__3408_ gnd vdd FILL
XFILL_2__2201_ gnd vdd FILL
XFILL_2__3181_ gnd vdd FILL
XFILL_2__2132_ gnd vdd FILL
XFILL_4__3048_ gnd vdd FILL
XFILL_2__2063_ gnd vdd FILL
XFILL_5__2812_ gnd vdd FILL
XFILL_7__1989_ gnd vdd FILL
XBUFX2_insert50 _3307_/Q _2022_/A vdd gnd BUFX2
XFILL_8__2521_ gnd vdd FILL
XBUFX2_insert61 _1993_/Y _2957_/B vdd gnd BUFX2
XBUFX2_insert83 _1858_/Y _2968_/A vdd gnd BUFX2
XFILL_8__2452_ gnd vdd FILL
XFILL_5__2743_ gnd vdd FILL
XBUFX2_insert72 _1765_/Y _2781_/A vdd gnd BUFX2
XBUFX2_insert94 _2083_/Y _2305_/A vdd gnd BUFX2
XFILL_2__2965_ gnd vdd FILL
XFILL_5__2674_ gnd vdd FILL
XFILL_2__2896_ gnd vdd FILL
XFILL_2__1916_ gnd vdd FILL
XFILL_0__1980_ gnd vdd FILL
XFILL_8__2383_ gnd vdd FILL
XFILL_2__1847_ gnd vdd FILL
XFILL_8_BUFX2_insert20 gnd vdd FILL
XFILL_8_BUFX2_insert42 gnd vdd FILL
XFILL_8_BUFX2_insert64 gnd vdd FILL
XFILL_8__3004_ gnd vdd FILL
XFILL_2__1778_ gnd vdd FILL
XFILL_0__3581_ gnd vdd FILL
XFILL_8_BUFX2_insert75 gnd vdd FILL
XFILL_8_BUFX2_insert53 gnd vdd FILL
XFILL_0__2601_ gnd vdd FILL
XFILL_8_BUFX2_insert97 gnd vdd FILL
XFILL_2__3517_ gnd vdd FILL
XFILL_3__2310_ gnd vdd FILL
XFILL_0__2532_ gnd vdd FILL
XFILL_5__3226_ gnd vdd FILL
XFILL_8_BUFX2_insert86 gnd vdd FILL
XFILL_2__3448_ gnd vdd FILL
XFILL_3__2241_ gnd vdd FILL
XFILL_3__2172_ gnd vdd FILL
XFILL_0__2463_ gnd vdd FILL
XFILL_5__3157_ gnd vdd FILL
XFILL_2__3379_ gnd vdd FILL
XFILL_5__3088_ gnd vdd FILL
XFILL_0__2394_ gnd vdd FILL
XFILL_5__2108_ gnd vdd FILL
XFILL_6__2921_ gnd vdd FILL
XFILL_5__2039_ gnd vdd FILL
X_1973_ _3079_/A _1984_/B _1973_/C _1974_/C vdd gnd OAI21X1
XFILL_6__2852_ gnd vdd FILL
XFILL_9__2561_ gnd vdd FILL
XFILL_0__3015_ gnd vdd FILL
XFILL_6__2783_ gnd vdd FILL
XFILL_6__1803_ gnd vdd FILL
XFILL_8__2719_ gnd vdd FILL
XFILL_6__1734_ gnd vdd FILL
XFILL_3__1956_ gnd vdd FILL
X_3574_ _3574_/D vdd _3578_/R _3577_/CLK _3574_/Q vdd gnd DFFSR
XFILL_6__3404_ gnd vdd FILL
X_2525_ _3248_/Q _2711_/B vdd gnd INVX1
XFILL_3__1887_ gnd vdd FILL
X_2456_ _2502_/C _2456_/B _2457_/B vdd gnd NOR2X1
XFILL_1__2710_ gnd vdd FILL
XFILL_1__2641_ gnd vdd FILL
XFILL_3__3557_ gnd vdd FILL
X_2387_ _2423_/A _2468_/A _2392_/C vdd gnd NAND2X1
XFILL_4__2350_ gnd vdd FILL
XFILL_3__3488_ gnd vdd FILL
XFILL_6__2217_ gnd vdd FILL
XFILL_4__2281_ gnd vdd FILL
XFILL_1__2572_ gnd vdd FILL
XFILL_3__2508_ gnd vdd FILL
XFILL_6__3197_ gnd vdd FILL
XFILL_3__2439_ gnd vdd FILL
X_3008_ _3260_/Q _3262_/Q _3013_/C vdd gnd NOR2X1
XFILL_6__2148_ gnd vdd FILL
XFILL_6__2079_ gnd vdd FILL
XFILL_7__2961_ gnd vdd FILL
XFILL_7__1912_ gnd vdd FILL
XFILL_1__3124_ gnd vdd FILL
XFILL_7__2892_ gnd vdd FILL
XFILL_1__3055_ gnd vdd FILL
XFILL_7__1843_ gnd vdd FILL
XFILL_1__2006_ gnd vdd FILL
XFILL_7__1774_ gnd vdd FILL
XFILL_7__3513_ gnd vdd FILL
XFILL_4__1996_ gnd vdd FILL
XFILL_7__3444_ gnd vdd FILL
XFILL_2__2750_ gnd vdd FILL
XFILL_1__2908_ gnd vdd FILL
XFILL_7__3375_ gnd vdd FILL
XFILL_2__1701_ gnd vdd FILL
XFILL_7__2326_ gnd vdd FILL
XFILL_5__2390_ gnd vdd FILL
XFILL_4__3597_ gnd vdd FILL
XFILL_2__2681_ gnd vdd FILL
XFILL_4__2617_ gnd vdd FILL
XFILL_1__2839_ gnd vdd FILL
XFILL_4__2548_ gnd vdd FILL
XFILL_7__2257_ gnd vdd FILL
XFILL_7__2188_ gnd vdd FILL
XFILL_5__3011_ gnd vdd FILL
XFILL_4__2479_ gnd vdd FILL
XCLKBUF1_insert28 clk _3346_/CLK vdd gnd CLKBUF1
XFILL_8__1952_ gnd vdd FILL
XFILL_2__3164_ gnd vdd FILL
XFILL_2__3095_ gnd vdd FILL
XFILL_2__2115_ gnd vdd FILL
XFILL_8__1883_ gnd vdd FILL
XFILL_2__2046_ gnd vdd FILL
XFILL183450x35250 gnd vdd FILL
XFILL_8__3553_ gnd vdd FILL
XFILL_8__2504_ gnd vdd FILL
XFILL_8__3484_ gnd vdd FILL
XFILL_3__2790_ gnd vdd FILL
XFILL_5__2726_ gnd vdd FILL
XFILL_3__1810_ gnd vdd FILL
XFILL_2__2948_ gnd vdd FILL
XFILL_3__1741_ gnd vdd FILL
XFILL_8__2435_ gnd vdd FILL
X_2310_ _2310_/A _2310_/B _2313_/A vdd gnd NAND2X1
XFILL_0__1963_ gnd vdd FILL
X_3290_ _3290_/D vdd _3355_/R _3355_/CLK _3290_/Q vdd gnd DFFSR
XFILL_8__2366_ gnd vdd FILL
XFILL_5__2657_ gnd vdd FILL
XFILL_2__2879_ gnd vdd FILL
X_2241_ _2329_/A _2244_/B vdd gnd INVX1
XFILL_5__2588_ gnd vdd FILL
XFILL_6__3120_ gnd vdd FILL
XFILL_3__3411_ gnd vdd FILL
XFILL_8__2297_ gnd vdd FILL
XFILL_0__1894_ gnd vdd FILL
X_2172_ _2814_/A _2172_/B _2172_/C _2298_/D _2339_/C vdd gnd AOI22X1
XFILL_6__3051_ gnd vdd FILL
XFILL_0__3564_ gnd vdd FILL
XFILL_6__2002_ gnd vdd FILL
XFILL_5__3209_ gnd vdd FILL
XFILL_0__2515_ gnd vdd FILL
XFILL_0__3495_ gnd vdd FILL
XFILL_3__2224_ gnd vdd FILL
XFILL_3__2155_ gnd vdd FILL
XFILL_0__2446_ gnd vdd FILL
XFILL_3__2086_ gnd vdd FILL
XFILL_0__2377_ gnd vdd FILL
XFILL_6__2904_ gnd vdd FILL
X_1956_ _3328_/Q _3092_/A _1959_/A vdd gnd NAND2X1
XFILL_6__2835_ gnd vdd FILL
XFILL_4_BUFX2_insert51 gnd vdd FILL
XFILL_4_BUFX2_insert40 gnd vdd FILL
XFILL_4_BUFX2_insert84 gnd vdd FILL
XFILL_4_BUFX2_insert62 gnd vdd FILL
XFILL_4_BUFX2_insert73 gnd vdd FILL
X_1887_ _2072_/B _2960_/B vdd gnd INVX1
XFILL_4__1850_ gnd vdd FILL
XFILL_4_BUFX2_insert95 gnd vdd FILL
XFILL_6__2766_ gnd vdd FILL
X_3557_ _3575_/Q _3560_/A _3558_/C vdd gnd NAND2X1
XFILL_4__3520_ gnd vdd FILL
XFILL_3__2988_ gnd vdd FILL
XFILL_6__1717_ gnd vdd FILL
XFILL_6__2697_ gnd vdd FILL
XFILL_4__1781_ gnd vdd FILL
XFILL_3__1939_ gnd vdd FILL
X_2508_ _3577_/Q _2508_/B _2512_/A vdd gnd NAND2X1
X_3488_ _3545_/A _3488_/B _3544_/C _3492_/B vdd gnd OAI21X1
XFILL_4__3451_ gnd vdd FILL
XFILL_7__3160_ gnd vdd FILL
XFILL_4__3382_ gnd vdd FILL
XFILL_4__2402_ gnd vdd FILL
XFILL_7__2111_ gnd vdd FILL
X_2439_ _2439_/A _2523_/A _2508_/B vdd gnd NAND2X1
XFILL_7__3091_ gnd vdd FILL
XFILL_4__2333_ gnd vdd FILL
XFILL_1__2624_ gnd vdd FILL
XFILL_7__2042_ gnd vdd FILL
XFILL_1__2555_ gnd vdd FILL
XFILL_4__2264_ gnd vdd FILL
XFILL_4__2195_ gnd vdd FILL
XFILL_1__2486_ gnd vdd FILL
XFILL_7__2944_ gnd vdd FILL
XFILL_1__3107_ gnd vdd FILL
XFILL_7__2875_ gnd vdd FILL
XFILL_5__1890_ gnd vdd FILL
XFILL_7__1826_ gnd vdd FILL
XFILL_1__3038_ gnd vdd FILL
XFILL_7__1757_ gnd vdd FILL
XFILL_4__1979_ gnd vdd FILL
XFILL_5__3560_ gnd vdd FILL
XFILL_2__2802_ gnd vdd FILL
XFILL_7__1688_ gnd vdd FILL
XFILL_5__3491_ gnd vdd FILL
XFILL_7__3427_ gnd vdd FILL
XFILL_8__2220_ gnd vdd FILL
XFILL_5__2511_ gnd vdd FILL
XFILL_2__2733_ gnd vdd FILL
XFILL_5__2442_ gnd vdd FILL
XFILL_8__2151_ gnd vdd FILL
XFILL_2__2664_ gnd vdd FILL
XFILL_7__2309_ gnd vdd FILL
XFILL_8__2082_ gnd vdd FILL
XFILL_5__2373_ gnd vdd FILL
XFILL_2__2595_ gnd vdd FILL
XFILL_0__2300_ gnd vdd FILL
XFILL_8__2984_ gnd vdd FILL
XFILL_2__3216_ gnd vdd FILL
XFILL_8__1935_ gnd vdd FILL
XFILL_2__3147_ gnd vdd FILL
XFILL_0__2231_ gnd vdd FILL
XFILL_0__2162_ gnd vdd FILL
X_1810_ _2453_/A _2781_/B _1810_/C _2435_/A vdd gnd OAI21X1
XFILL_8__1866_ gnd vdd FILL
X_2790_ _2814_/A _2933_/B _2790_/C _3259_/D vdd gnd OAI21X1
XFILL_2__3078_ gnd vdd FILL
XFILL_3__2911_ gnd vdd FILL
XFILL_2__2029_ gnd vdd FILL
XFILL_6__2620_ gnd vdd FILL
XFILL_8__1797_ gnd vdd FILL
X_1741_ _2379_/A _3152_/C _2167_/A vdd gnd NAND2X1
XFILL_0__2093_ gnd vdd FILL
XFILL_3__2842_ gnd vdd FILL
XFILL_8__3536_ gnd vdd FILL
XFILL_8__3467_ gnd vdd FILL
X_3411_ _3411_/A _3428_/B _3411_/C _3509_/C vdd gnd OAI21X1
XFILL_6__2551_ gnd vdd FILL
X_3342_ _3342_/D vdd _3345_/R _3576_/CLK _3342_/Q vdd gnd DFFSR
XFILL_8__2418_ gnd vdd FILL
XFILL_6__2482_ gnd vdd FILL
XFILL_5__2709_ gnd vdd FILL
XFILL_3__2773_ gnd vdd FILL
XFILL_8__3398_ gnd vdd FILL
XFILL_0__2995_ gnd vdd FILL
XFILL_3__1724_ gnd vdd FILL
X_3273_ _3273_/D vdd _3346_/R _3346_/CLK _3273_/Q vdd gnd DFFSR
XFILL_0__1946_ gnd vdd FILL
XFILL_8__2349_ gnd vdd FILL
XFILL_0__1877_ gnd vdd FILL
X_2224_ _2224_/A _2320_/B _2345_/B _2225_/C vdd gnd NAND3X1
XFILL_6_CLKBUF1_insert37 gnd vdd FILL
XFILL_6__3103_ gnd vdd FILL
X_2155_ _2330_/A _2155_/B _2319_/B vdd gnd NAND2X1
XFILL_6__3034_ gnd vdd FILL
XFILL_0__3547_ gnd vdd FILL
X_2086_ _2305_/A _2312_/C _2087_/C vdd gnd NOR2X1
XFILL_1__2340_ gnd vdd FILL
XFILL_0__3478_ gnd vdd FILL
XFILL_1__2271_ gnd vdd FILL
XFILL_3__2207_ gnd vdd FILL
XFILL_4_CLKBUF1_insert30 gnd vdd FILL
XFILL_3__3187_ gnd vdd FILL
XFILL_0__2429_ gnd vdd FILL
XFILL_3__2138_ gnd vdd FILL
XFILL_4__2951_ gnd vdd FILL
X_2988_ _2988_/A _2988_/B _2988_/C _3310_/D vdd gnd OAI21X1
XFILL_3__2069_ gnd vdd FILL
X_1939_ _3334_/Q _3110_/A _3127_/B _3343_/Q _1941_/C vdd gnd AOI22X1
XFILL_4__1902_ gnd vdd FILL
XFILL_7__2660_ gnd vdd FILL
XFILL_6__2818_ gnd vdd FILL
XFILL_4__2882_ gnd vdd FILL
XFILL_7__2591_ gnd vdd FILL
XFILL_6__2749_ gnd vdd FILL
XFILL_4__1833_ gnd vdd FILL
XFILL_9__2458_ gnd vdd FILL
XFILL_4__1764_ gnd vdd FILL
XFILL_4__3503_ gnd vdd FILL
XFILL_1__1986_ gnd vdd FILL
XFILL_7__3212_ gnd vdd FILL
XFILL_4__3434_ gnd vdd FILL
XFILL_4__1695_ gnd vdd FILL
XFILL_7__3143_ gnd vdd FILL
XFILL_7__3074_ gnd vdd FILL
XFILL_4__3365_ gnd vdd FILL
XFILL_1__2607_ gnd vdd FILL
XFILL_7__2025_ gnd vdd FILL
XFILL_0_BUFX2_insert60 gnd vdd FILL
XFILL_1__3587_ gnd vdd FILL
XFILL_2__2380_ gnd vdd FILL
XFILL_4__2316_ gnd vdd FILL
XFILL_0_BUFX2_insert93 gnd vdd FILL
XFILL_0_BUFX2_insert82 gnd vdd FILL
XFILL_4__2247_ gnd vdd FILL
XFILL_1__2538_ gnd vdd FILL
XFILL_0_BUFX2_insert71 gnd vdd FILL
XFILL_1__2469_ gnd vdd FILL
XFILL_2__3001_ gnd vdd FILL
XFILL_4__2178_ gnd vdd FILL
XFILL_5__2991_ gnd vdd FILL
XFILL_8__1720_ gnd vdd FILL
XFILL_7__2927_ gnd vdd FILL
XFILL_5__1942_ gnd vdd FILL
XFILL_7__2858_ gnd vdd FILL
XFILL_5__1873_ gnd vdd FILL
XFILL_7__2789_ gnd vdd FILL
XFILL_7__1809_ gnd vdd FILL
XFILL_5__3543_ gnd vdd FILL
XFILL_5__3474_ gnd vdd FILL
XFILL_8__2203_ gnd vdd FILL
XFILL_2__2716_ gnd vdd FILL
XFILL_0__2780_ gnd vdd FILL
XFILL_0__1800_ gnd vdd FILL
XFILL_8__3183_ gnd vdd FILL
XFILL_5__2425_ gnd vdd FILL
XFILL_8__2134_ gnd vdd FILL
XFILL_0__1731_ gnd vdd FILL
XFILL_5__2356_ gnd vdd FILL
XFILL_2__2647_ gnd vdd FILL
XFILL_2__2578_ gnd vdd FILL
XFILL_0__3401_ gnd vdd FILL
XFILL_8__2065_ gnd vdd FILL
XFILL_3__3110_ gnd vdd FILL
XFILL_5__2287_ gnd vdd FILL
XFILL_3__3041_ gnd vdd FILL
X_2911_ _2911_/A _2911_/B _2922_/B _2912_/B vdd gnd OAI21X1
XFILL_0__2214_ gnd vdd FILL
XFILL_8__2967_ gnd vdd FILL
XFILL_8__1918_ gnd vdd FILL
X_2842_ _2915_/A _2921_/A _2895_/A vdd gnd NAND2X1
XFILL_8__2898_ gnd vdd FILL
XFILL_6__1982_ gnd vdd FILL
XFILL_0__3194_ gnd vdd FILL
XFILL_0__2145_ gnd vdd FILL
X_2773_ _2773_/A _2773_/B _2773_/C _2776_/B vdd gnd OAI21X1
XFILL_8__1849_ gnd vdd FILL
XFILL_0__2076_ gnd vdd FILL
X_1724_ _3157_/A _1846_/B _1725_/A vdd gnd NAND2X1
XFILL_6__3583_ gnd vdd FILL
XFILL_6__2603_ gnd vdd FILL
XFILL_3__2825_ gnd vdd FILL
XFILL_8__3519_ gnd vdd FILL
XFILL_6__2534_ gnd vdd FILL
XFILL_3__2756_ gnd vdd FILL
XFILL_1__1840_ gnd vdd FILL
X_3325_ _3325_/D vdd _3345_/R _3577_/CLK _3325_/Q vdd gnd DFFSR
XFILL_0__2978_ gnd vdd FILL
XFILL_1__1771_ gnd vdd FILL
XFILL_3__1707_ gnd vdd FILL
XFILL_6__2465_ gnd vdd FILL
XFILL_0__1929_ gnd vdd FILL
XFILL_1__3510_ gnd vdd FILL
XFILL_6__2396_ gnd vdd FILL
X_3256_ _3256_/D vdd _3363_/R _3363_/CLK _3256_/Q vdd gnd DFFSR
XFILL_3__2687_ gnd vdd FILL
X_2207_ _2786_/A _3163_/A _2208_/C vdd gnd NAND2X1
XFILL_1__3441_ gnd vdd FILL
X_3187_ _3187_/A _3193_/A vdd gnd INVX1
XFILL_4__3150_ gnd vdd FILL
XFILL_1__3372_ gnd vdd FILL
XFILL_4__2101_ gnd vdd FILL
X_2138_ _3176_/A _2433_/A vdd gnd INVX1
XFILL_4__3081_ gnd vdd FILL
XFILL_6__3017_ gnd vdd FILL
XFILL_1__2323_ gnd vdd FILL
X_2069_ _2966_/B _2958_/A _3022_/A _2347_/A vdd gnd OAI21X1
XFILL_4__2032_ gnd vdd FILL
XFILL_9__1958_ gnd vdd FILL
XFILL_1__2254_ gnd vdd FILL
XFILL_1__2185_ gnd vdd FILL
XFILL_7__2712_ gnd vdd FILL
XFILL_4__2934_ gnd vdd FILL
XFILL_7__2643_ gnd vdd FILL
XFILL_4__2865_ gnd vdd FILL
XFILL_2__1880_ gnd vdd FILL
XFILL_4__1816_ gnd vdd FILL
XFILL_7__2574_ gnd vdd FILL
XFILL_4__2796_ gnd vdd FILL
XFILL_2__3550_ gnd vdd FILL
XFILL_4__1747_ gnd vdd FILL
XFILL_1__1969_ gnd vdd FILL
XFILL_2__2501_ gnd vdd FILL
XFILL_2__3481_ gnd vdd FILL
XFILL_7__3126_ gnd vdd FILL
XFILL_4__3417_ gnd vdd FILL
XFILL_5__2210_ gnd vdd FILL
XFILL_5__3190_ gnd vdd FILL
XFILL_5__2141_ gnd vdd FILL
XFILL_2__2432_ gnd vdd FILL
XFILL_7__3057_ gnd vdd FILL
XFILL_2__2363_ gnd vdd FILL
XFILL_5__2072_ gnd vdd FILL
XFILL_7__2008_ gnd vdd FILL
XFILL_5_BUFX2_insert17 gnd vdd FILL
XFILL_2__2294_ gnd vdd FILL
XFILL_8__2821_ gnd vdd FILL
XFILL_5_BUFX2_insert39 gnd vdd FILL
XFILL_8__2752_ gnd vdd FILL
XFILL_5__2974_ gnd vdd FILL
XFILL_8__1703_ gnd vdd FILL
XFILL_8__2683_ gnd vdd FILL
XFILL_5__1925_ gnd vdd FILL
XFILL_5__1856_ gnd vdd FILL
XFILL_0__2901_ gnd vdd FILL
XFILL_3__2610_ gnd vdd FILL
XFILL_5__1787_ gnd vdd FILL
XFILL_5__3526_ gnd vdd FILL
XFILL_0__2832_ gnd vdd FILL
XFILL_3__3590_ gnd vdd FILL
XFILL_6__2250_ gnd vdd FILL
X_3110_ _3110_/A _3125_/B vdd gnd INVX2
XFILL_5__3457_ gnd vdd FILL
XFILL_3__2541_ gnd vdd FILL
XFILL_3__2472_ gnd vdd FILL
XFILL_0__2763_ gnd vdd FILL
XFILL_8__3166_ gnd vdd FILL
XFILL_5__2408_ gnd vdd FILL
XFILL_5__3388_ gnd vdd FILL
XFILL_6__2181_ gnd vdd FILL
XFILL_8__3097_ gnd vdd FILL
XFILL_8__2117_ gnd vdd FILL
X_3041_ _3077_/C _3041_/B _3042_/C vdd gnd NOR2X1
XFILL_0__2694_ gnd vdd FILL
XFILL_0__1714_ gnd vdd FILL
XFILL_5__2339_ gnd vdd FILL
XFILL_8__2048_ gnd vdd FILL
XFILL_3__3024_ gnd vdd FILL
XFILL_6__1965_ gnd vdd FILL
X_2825_ _2885_/B _2835_/B _2826_/C vdd gnd NOR2X1
XFILL_0__3177_ gnd vdd FILL
XFILL_0__2128_ gnd vdd FILL
XFILL_9__3413_ gnd vdd FILL
XFILL_6__1896_ gnd vdd FILL
X_2756_ _3252_/Q _2756_/B _2757_/D vdd gnd NAND2X1
XFILL_1__2941_ gnd vdd FILL
X_1707_ _3566_/A _3296_/Q _1708_/C vdd gnd OR2X2
X_2687_ _2687_/A _2687_/B _2741_/B vdd gnd NAND2X1
XFILL_0__2059_ gnd vdd FILL
XFILL_4__2650_ gnd vdd FILL
XFILL_3__2808_ gnd vdd FILL
XFILL_6__3566_ gnd vdd FILL
XFILL_1__2872_ gnd vdd FILL
XFILL_6__3497_ gnd vdd FILL
XFILL_1__1823_ gnd vdd FILL
XFILL_7__2290_ gnd vdd FILL
XFILL_6__2517_ gnd vdd FILL
XFILL_4__2581_ gnd vdd FILL
XFILL_3__2739_ gnd vdd FILL
XFILL_6__2448_ gnd vdd FILL
X_3308_ _3308_/D vdd _3353_/R _3578_/CLK _3308_/Q vdd gnd DFFSR
XFILL_1__1754_ gnd vdd FILL
X_3239_ _3239_/D vdd _3362_/R _3363_/CLK _3239_/Q vdd gnd DFFSR
XFILL_6__2379_ gnd vdd FILL
XFILL_4__3202_ gnd vdd FILL
XFILL_1__3424_ gnd vdd FILL
XFILL_4__3133_ gnd vdd FILL
XFILL_4__3064_ gnd vdd FILL
XFILL_1__2306_ gnd vdd FILL
XFILL_4__2015_ gnd vdd FILL
XFILL_1__2237_ gnd vdd FILL
XFILL_1__2168_ gnd vdd FILL
XFILL_4__2917_ gnd vdd FILL
XFILL_2__2981_ gnd vdd FILL
XFILL_5__1710_ gnd vdd FILL
XFILL_3_BUFX2_insert1 gnd vdd FILL
XFILL_1__2099_ gnd vdd FILL
XFILL_2__1932_ gnd vdd FILL
XFILL_5__2690_ gnd vdd FILL
XFILL_7__2626_ gnd vdd FILL
XFILL_4__2848_ gnd vdd FILL
XFILL_7__2557_ gnd vdd FILL
XFILL_2__1863_ gnd vdd FILL
XFILL_2__3602_ gnd vdd FILL
XFILL_4__2779_ gnd vdd FILL
XFILL_7__2488_ gnd vdd FILL
XFILL_8__3020_ gnd vdd FILL
XFILL_2__1794_ gnd vdd FILL
XFILL_2__3533_ gnd vdd FILL
XFILL_2__3464_ gnd vdd FILL
XFILL181350x109350 gnd vdd FILL
XFILL_7__3109_ gnd vdd FILL
XFILL_2__2415_ gnd vdd FILL
XFILL_5__3173_ gnd vdd FILL
XFILL_2__3395_ gnd vdd FILL
XFILL_5__2124_ gnd vdd FILL
XFILL_2__2346_ gnd vdd FILL
XFILL_5__2055_ gnd vdd FILL
XFILL_2__2277_ gnd vdd FILL
XFILL_0__3100_ gnd vdd FILL
XFILL_8__2804_ gnd vdd FILL
XFILL_0__3031_ gnd vdd FILL
XFILL_5__2957_ gnd vdd FILL
XFILL_6__1750_ gnd vdd FILL
XFILL_8__2735_ gnd vdd FILL
XFILL_3__1972_ gnd vdd FILL
X_3590_ _3590_/A AB[5] vdd gnd BUFX2
X_2610_ _2639_/B _2611_/B vdd gnd INVX1
XFILL_8__2666_ gnd vdd FILL
XFILL_5__1908_ gnd vdd FILL
XFILL_5__2888_ gnd vdd FILL
XFILL_8__2597_ gnd vdd FILL
X_2541_ _2948_/A _2541_/B _2541_/C _2542_/A vdd gnd OAI21X1
XFILL_6__3420_ gnd vdd FILL
XFILL_5__1839_ gnd vdd FILL
X_2472_ _2472_/A _2472_/B _2473_/C vdd gnd AND2X2
XFILL_5__3509_ gnd vdd FILL
XFILL_6__2302_ gnd vdd FILL
XFILL_1_BUFX2_insert15 gnd vdd FILL
XFILL_1_BUFX2_insert26 gnd vdd FILL
XFILL_1_BUFX2_insert59 gnd vdd FILL
XFILL_1_BUFX2_insert48 gnd vdd FILL
XFILL_0__2815_ gnd vdd FILL
XFILL_6_BUFX2_insert5 gnd vdd FILL
XFILL_3__2524_ gnd vdd FILL
XFILL_8__3218_ gnd vdd FILL
XFILL184650x140550 gnd vdd FILL
XFILL_6__2233_ gnd vdd FILL
XFILL_0__2746_ gnd vdd FILL
XFILL_8__3149_ gnd vdd FILL
XFILL_6__2164_ gnd vdd FILL
X_3024_ _3024_/A _3145_/B _3088_/S _3025_/B vdd gnd OAI21X1
XFILL_3__2455_ gnd vdd FILL
XFILL_3__2386_ gnd vdd FILL
XFILL_0__2677_ gnd vdd FILL
XFILL_6__2095_ gnd vdd FILL
XFILL_1__3140_ gnd vdd FILL
XFILL_1_CLKBUF1_insert38 gnd vdd FILL
XFILL_3__3007_ gnd vdd FILL
XFILL_1__3071_ gnd vdd FILL
XFILL_1__2022_ gnd vdd FILL
XFILL_0__3229_ gnd vdd FILL
XFILL_6__2997_ gnd vdd FILL
XFILL_7__1790_ gnd vdd FILL
XFILL_6__1948_ gnd vdd FILL
X_2808_ _3265_/Q _2973_/A vdd gnd INVX1
XFILL_6__1879_ gnd vdd FILL
XFILL_7__3460_ gnd vdd FILL
XFILL_4__2702_ gnd vdd FILL
X_2739_ _3294_/D _2772_/B _2739_/C _2757_/A vdd gnd AOI21X1
XFILL_1__2924_ gnd vdd FILL
XFILL_7__3391_ gnd vdd FILL
XFILL_7__2411_ gnd vdd FILL
XFILL_7__2342_ gnd vdd FILL
XFILL_4__2633_ gnd vdd FILL
XFILL_6__3549_ gnd vdd FILL
XFILL_1__2855_ gnd vdd FILL
XFILL_4__2564_ gnd vdd FILL
XFILL_7__2273_ gnd vdd FILL
XFILL_1__2786_ gnd vdd FILL
XFILL_1__1806_ gnd vdd FILL
XFILL_4__2495_ gnd vdd FILL
XFILL_1__1737_ gnd vdd FILL
XFILL_4__3116_ gnd vdd FILL
XFILL_1__3407_ gnd vdd FILL
XFILL_2__2200_ gnd vdd FILL
XFILL_2__3180_ gnd vdd FILL
XFILL_9_BUFX2_insert9 gnd vdd FILL
XFILL_2__2131_ gnd vdd FILL
XFILL_4__3047_ gnd vdd FILL
XFILL_2__2062_ gnd vdd FILL
XFILL_5__2811_ gnd vdd FILL
XFILL_7__1988_ gnd vdd FILL
XBUFX2_insert51 _3307_/Q _2033_/A vdd gnd BUFX2
XBUFX2_insert40 _1734_/Y _2430_/A vdd gnd BUFX2
XFILL_8__2520_ gnd vdd FILL
XBUFX2_insert84 _1858_/Y _2888_/B vdd gnd BUFX2
XBUFX2_insert62 _1993_/Y _2897_/C vdd gnd BUFX2
XBUFX2_insert73 _1694_/Y _2814_/A vdd gnd BUFX2
XFILL_8__2451_ gnd vdd FILL
XFILL_5__2742_ gnd vdd FILL
XBUFX2_insert95 _2083_/Y _2885_/B vdd gnd BUFX2
XFILL_2__2964_ gnd vdd FILL
XFILL_7__2609_ gnd vdd FILL
XFILL_5__2673_ gnd vdd FILL
XFILL_2__2895_ gnd vdd FILL
XFILL_8__2382_ gnd vdd FILL
XFILL_2__1915_ gnd vdd FILL
XFILL_7__3589_ gnd vdd FILL
XFILL_2__1846_ gnd vdd FILL
XFILL_8_BUFX2_insert21 gnd vdd FILL
XFILL_8_BUFX2_insert10 gnd vdd FILL
XFILL_2__3516_ gnd vdd FILL
XFILL_8__3003_ gnd vdd FILL
XFILL_8_BUFX2_insert43 gnd vdd FILL
XFILL_2__1777_ gnd vdd FILL
XFILL_0__3580_ gnd vdd FILL
XFILL_8_BUFX2_insert65 gnd vdd FILL
XFILL_0__2600_ gnd vdd FILL
XFILL_8_BUFX2_insert54 gnd vdd FILL
XFILL_8_BUFX2_insert76 gnd vdd FILL
XFILL_8_BUFX2_insert87 gnd vdd FILL
XFILL_0__2531_ gnd vdd FILL
XFILL_5__3225_ gnd vdd FILL
XFILL_2__3447_ gnd vdd FILL
XFILL_3__2240_ gnd vdd FILL
XFILL_5__3156_ gnd vdd FILL
XFILL_2__3378_ gnd vdd FILL
XFILL_3__2171_ gnd vdd FILL
XFILL_0__2462_ gnd vdd FILL
XFILL_5__2107_ gnd vdd FILL
XFILL_5__3087_ gnd vdd FILL
XFILL_0__2393_ gnd vdd FILL
XFILL_2__2329_ gnd vdd FILL
XFILL_6__2920_ gnd vdd FILL
XFILL_5__2038_ gnd vdd FILL
XFILL_6__2851_ gnd vdd FILL
X_1972_ _2760_/B _1973_/C vdd gnd INVX1
XFILL_6__1802_ gnd vdd FILL
XFILL_0__3014_ gnd vdd FILL
XFILL_8__2718_ gnd vdd FILL
XFILL_6__2782_ gnd vdd FILL
XFILL_6__1733_ gnd vdd FILL
X_3573_ _3573_/D vdd _3578_/R _3573_/CLK _3573_/Q vdd gnd DFFSR
XFILL_3__1955_ gnd vdd FILL
XFILL_8__2649_ gnd vdd FILL
XFILL_6__3403_ gnd vdd FILL
XFILL_3__1886_ gnd vdd FILL
X_2524_ _3216_/A _3216_/B _3593_/A vdd gnd OR2X2
XFILL184650x152250 gnd vdd FILL
X_2455_ _2510_/B _2455_/B _2456_/B vdd gnd NAND2X1
XFILL184350x160050 gnd vdd FILL
X_2386_ _2386_/A _2386_/B _2386_/C _3595_/A vdd gnd NAND3X1
XFILL_1__2640_ gnd vdd FILL
XFILL_3__3556_ gnd vdd FILL
XFILL_3__3487_ gnd vdd FILL
XFILL_6__2216_ gnd vdd FILL
XFILL_4__2280_ gnd vdd FILL
XFILL_3__2507_ gnd vdd FILL
XFILL_1__2571_ gnd vdd FILL
XFILL_6__3196_ gnd vdd FILL
XFILL_0__2729_ gnd vdd FILL
XFILL_3__2438_ gnd vdd FILL
X_3007_ _3007_/A _3007_/B _3007_/C _3015_/A vdd gnd NAND3X1
XFILL_6__2147_ gnd vdd FILL
XFILL_6__2078_ gnd vdd FILL
XFILL_7__2960_ gnd vdd FILL
XFILL_3__2369_ gnd vdd FILL
XFILL_1__3123_ gnd vdd FILL
XFILL_7__1911_ gnd vdd FILL
XFILL_7__2891_ gnd vdd FILL
XFILL_1__3054_ gnd vdd FILL
XFILL_7__1842_ gnd vdd FILL
XFILL_1__2005_ gnd vdd FILL
XFILL_7__1773_ gnd vdd FILL
XFILL_7__3512_ gnd vdd FILL
XFILL_4__1995_ gnd vdd FILL
XFILL_7__3443_ gnd vdd FILL
XFILL_1__2907_ gnd vdd FILL
XFILL_7__3374_ gnd vdd FILL
XFILL_2__1700_ gnd vdd FILL
XFILL_2__2680_ gnd vdd FILL
XFILL_4__2616_ gnd vdd FILL
XFILL_1__2838_ gnd vdd FILL
XFILL_7__2325_ gnd vdd FILL
XFILL_4__3596_ gnd vdd FILL
XFILL_7__2256_ gnd vdd FILL
XFILL_4__2547_ gnd vdd FILL
XFILL_4__2478_ gnd vdd FILL
XFILL_1__2769_ gnd vdd FILL
XFILL_5__3010_ gnd vdd FILL
XFILL_7__2187_ gnd vdd FILL
XFILL_2__3232_ gnd vdd FILL
XCLKBUF1_insert29 clk _3578_/CLK vdd gnd CLKBUF1
XFILL_8__1951_ gnd vdd FILL
XFILL_2__3163_ gnd vdd FILL
XFILL_2__3094_ gnd vdd FILL
XFILL_2__2114_ gnd vdd FILL
XFILL_8__1882_ gnd vdd FILL
XFILL_2__2045_ gnd vdd FILL
XFILL_8__3552_ gnd vdd FILL
XFILL_8__2503_ gnd vdd FILL
XFILL_8__3483_ gnd vdd FILL
XFILL_5__2725_ gnd vdd FILL
XFILL_2__2947_ gnd vdd FILL
XFILL_3__1740_ gnd vdd FILL
XFILL_8__2434_ gnd vdd FILL
XFILL_0__1962_ gnd vdd FILL
XFILL_8__2365_ gnd vdd FILL
XFILL_5__2656_ gnd vdd FILL
XFILL_3__3410_ gnd vdd FILL
XFILL_2__2878_ gnd vdd FILL
X_2240_ _2278_/A _2240_/B _2240_/C _2329_/A vdd gnd OAI21X1
XFILL_5__2587_ gnd vdd FILL
XFILL_8__2296_ gnd vdd FILL
XFILL_2__1829_ gnd vdd FILL
XFILL_0__1893_ gnd vdd FILL
X_2171_ _2297_/A _2312_/A _2172_/C vdd gnd NOR2X1
XFILL_6__3050_ gnd vdd FILL
XFILL_6__2001_ gnd vdd FILL
XFILL_0__3563_ gnd vdd FILL
XFILL_5__3208_ gnd vdd FILL
XFILL_0__3494_ gnd vdd FILL
XFILL_3__2223_ gnd vdd FILL
XFILL_0__2514_ gnd vdd FILL
XFILL_5__3139_ gnd vdd FILL
XFILL_0__2445_ gnd vdd FILL
XFILL_3__2154_ gnd vdd FILL
XFILL_3__2085_ gnd vdd FILL
XFILL_0__2376_ gnd vdd FILL
XFILL_6__2903_ gnd vdd FILL
X_1955_ _1986_/A _2412_/B _1955_/C _3421_/B vdd gnd OAI21X1
XFILL_6__2834_ gnd vdd FILL
XFILL_4_BUFX2_insert41 gnd vdd FILL
XFILL_4_BUFX2_insert63 gnd vdd FILL
XFILL_4_BUFX2_insert74 gnd vdd FILL
X_1886_ _2240_/B _3148_/B _1902_/A vdd gnd NOR2X1
XFILL_4_BUFX2_insert52 gnd vdd FILL
XFILL_4_BUFX2_insert96 gnd vdd FILL
XFILL_4_BUFX2_insert85 gnd vdd FILL
XFILL_3__2987_ gnd vdd FILL
XFILL_4__1780_ gnd vdd FILL
XFILL_6__2765_ gnd vdd FILL
XFILL_3__1938_ gnd vdd FILL
X_3556_ _3556_/A _3556_/B _3556_/C _3574_/D vdd gnd OAI21X1
XFILL_6__2696_ gnd vdd FILL
XFILL_6__1716_ gnd vdd FILL
X_2507_ _3213_/B _3591_/A vdd gnd INVX1
X_3487_ _3544_/B _3544_/A _3488_/B vdd gnd NOR2X1
XFILL_4__3450_ gnd vdd FILL
XFILL_3__1869_ gnd vdd FILL
XFILL_4__3381_ gnd vdd FILL
XFILL_4__2401_ gnd vdd FILL
X_2438_ _2438_/A _2438_/B _2439_/A vdd gnd NOR2X1
XFILL_7__2110_ gnd vdd FILL
XFILL_7__3090_ gnd vdd FILL
XFILL_3__3539_ gnd vdd FILL
XFILL_4__2332_ gnd vdd FILL
X_2369_ _3314_/Q _2691_/A _2373_/B _2370_/C vdd gnd AOI21X1
XFILL_1__2623_ gnd vdd FILL
XFILL_7__2041_ gnd vdd FILL
XFILL_1__2554_ gnd vdd FILL
XFILL_4__2263_ gnd vdd FILL
XFILL_6__3179_ gnd vdd FILL
XFILL_4__2194_ gnd vdd FILL
XFILL_1__2485_ gnd vdd FILL
XFILL_7__2943_ gnd vdd FILL
XFILL_1__3106_ gnd vdd FILL
XFILL_7__2874_ gnd vdd FILL
XFILL_1__3037_ gnd vdd FILL
XFILL_7__1825_ gnd vdd FILL
XFILL_7__1756_ gnd vdd FILL
XFILL_4__1978_ gnd vdd FILL
XFILL_2__2801_ gnd vdd FILL
XFILL_5__2510_ gnd vdd FILL
XFILL_5__3490_ gnd vdd FILL
XFILL_7__3426_ gnd vdd FILL
XFILL_2__2732_ gnd vdd FILL
XFILL_8__2150_ gnd vdd FILL
XFILL_5__2441_ gnd vdd FILL
XFILL_5__2372_ gnd vdd FILL
XFILL_4__3579_ gnd vdd FILL
XFILL_2__2663_ gnd vdd FILL
XFILL_8__2081_ gnd vdd FILL
XFILL_7__2308_ gnd vdd FILL
XFILL_2__2594_ gnd vdd FILL
XFILL_7__2239_ gnd vdd FILL
XFILL_8__2983_ gnd vdd FILL
XFILL_2__3215_ gnd vdd FILL
XFILL_8__1934_ gnd vdd FILL
XFILL_2__3146_ gnd vdd FILL
XFILL_0__2230_ gnd vdd FILL
XFILL_0__2161_ gnd vdd FILL
XFILL_8__1865_ gnd vdd FILL
XFILL_2__3077_ gnd vdd FILL
XFILL_3__2910_ gnd vdd FILL
XFILL_2__2028_ gnd vdd FILL
X_1740_ _1933_/C _2442_/B _3152_/C vdd gnd NOR2X1
XFILL_0__2092_ gnd vdd FILL
XFILL_8__1796_ gnd vdd FILL
XFILL_3__2841_ gnd vdd FILL
XFILL_8__3535_ gnd vdd FILL
XFILL_8__3466_ gnd vdd FILL
X_3410_ _3442_/B _3411_/A _3466_/B _3411_/C vdd gnd OAI21X1
XFILL_6__2550_ gnd vdd FILL
XFILL182550x163950 gnd vdd FILL
X_3341_ _3341_/D vdd _3345_/R _3576_/CLK _3341_/Q vdd gnd DFFSR
XFILL_8__2417_ gnd vdd FILL
XFILL_6__2481_ gnd vdd FILL
XFILL_5__2708_ gnd vdd FILL
XFILL_3__2772_ gnd vdd FILL
XFILL_8__3397_ gnd vdd FILL
XFILL_0__2994_ gnd vdd FILL
XFILL_3__1723_ gnd vdd FILL
XFILL_5__2639_ gnd vdd FILL
X_3272_ _3272_/D vdd _3346_/R _3307_/CLK _3272_/Q vdd gnd DFFSR
XFILL_8__2348_ gnd vdd FILL
XFILL_0__1945_ gnd vdd FILL
XFILL_0__1876_ gnd vdd FILL
XFILL_6__3102_ gnd vdd FILL
XFILL_8__2279_ gnd vdd FILL
X_2223_ _3144_/B _3149_/C _2223_/C _2224_/A vdd gnd NAND3X1
XFILL_6_CLKBUF1_insert38 gnd vdd FILL
X_2154_ _2347_/C _2154_/B _2155_/B vdd gnd NOR2X1
XFILL_0__3546_ gnd vdd FILL
XFILL_6__3033_ gnd vdd FILL
X_2085_ _2894_/A _2270_/A _2312_/C vdd gnd NAND2X1
XFILL_0__3477_ gnd vdd FILL
XFILL_1__2270_ gnd vdd FILL
XFILL_3__2206_ gnd vdd FILL
XFILL_3__3186_ gnd vdd FILL
XFILL_0__2428_ gnd vdd FILL
XFILL_3__2137_ gnd vdd FILL
XFILL_0__2359_ gnd vdd FILL
XFILL_4_CLKBUF1_insert31 gnd vdd FILL
XFILL_4__2950_ gnd vdd FILL
X_2987_ _3310_/Q _2988_/A _2988_/C vdd gnd NAND2X1
XFILL_3__2068_ gnd vdd FILL
X_1938_ _3326_/Q _3092_/A _1941_/A vdd gnd NAND2X1
XFILL_4__2881_ gnd vdd FILL
XFILL_4__1901_ gnd vdd FILL
XFILL_6__2817_ gnd vdd FILL
X_1869_ _3340_/Q _3127_/B _1881_/A vdd gnd NAND2X1
XFILL_4__1832_ gnd vdd FILL
XFILL_7__2590_ gnd vdd FILL
XFILL_6__2748_ gnd vdd FILL
XFILL_4__1763_ gnd vdd FILL
XFILL_4__3502_ gnd vdd FILL
X_3539_ _3539_/A _3553_/B _3539_/C _3539_/D _3568_/D vdd gnd AOI22X1
XFILL_1__1985_ gnd vdd FILL
XFILL_4__1694_ gnd vdd FILL
XFILL_7__3211_ gnd vdd FILL
XFILL_6__2679_ gnd vdd FILL
XFILL_4__3433_ gnd vdd FILL
XFILL_7__3142_ gnd vdd FILL
XFILL_7__3073_ gnd vdd FILL
XFILL_4__3364_ gnd vdd FILL
XFILL_1__2606_ gnd vdd FILL
XFILL_0_BUFX2_insert50 gnd vdd FILL
XFILL_7__2024_ gnd vdd FILL
XFILL_4__2315_ gnd vdd FILL
XFILL_1__3586_ gnd vdd FILL
XFILL_0_BUFX2_insert61 gnd vdd FILL
XFILL_0_BUFX2_insert83 gnd vdd FILL
XFILL_4__2246_ gnd vdd FILL
XFILL_1__2537_ gnd vdd FILL
XFILL_0_BUFX2_insert72 gnd vdd FILL
XFILL_0_BUFX2_insert94 gnd vdd FILL
XFILL_1__2468_ gnd vdd FILL
XFILL_2__3000_ gnd vdd FILL
XFILL_4__2177_ gnd vdd FILL
XFILL_7__2926_ gnd vdd FILL
XFILL_5__2990_ gnd vdd FILL
XFILL_1__2399_ gnd vdd FILL
XFILL_5__1941_ gnd vdd FILL
XFILL_7__2857_ gnd vdd FILL
XFILL_5__1872_ gnd vdd FILL
XFILL_7__2788_ gnd vdd FILL
XFILL_7__1808_ gnd vdd FILL
XFILL_7__1739_ gnd vdd FILL
XFILL_5__3542_ gnd vdd FILL
XFILL_5__3473_ gnd vdd FILL
XFILL_7__3409_ gnd vdd FILL
XFILL_8__2202_ gnd vdd FILL
XFILL_5__2424_ gnd vdd FILL
XFILL_2__2715_ gnd vdd FILL
XFILL_8__3182_ gnd vdd FILL
XFILL_8__2133_ gnd vdd FILL
XFILL_0__1730_ gnd vdd FILL
XFILL_2__2646_ gnd vdd FILL
XFILL_8__2064_ gnd vdd FILL
XFILL_5__2355_ gnd vdd FILL
XFILL_0__3400_ gnd vdd FILL
XFILL_2__2577_ gnd vdd FILL
XFILL_5__2286_ gnd vdd FILL
XFILL_3__3040_ gnd vdd FILL
X_2910_ _2910_/A _2910_/B _2931_/B _2911_/B vdd gnd NAND3X1
XFILL_0__2213_ gnd vdd FILL
XFILL_8__2966_ gnd vdd FILL
X_2841_ _2841_/A _2919_/B _2862_/A _2841_/D _3271_/D vdd gnd AOI22X1
XFILL_2__3129_ gnd vdd FILL
XFILL_8__1917_ gnd vdd FILL
XFILL_8__2897_ gnd vdd FILL
XFILL_6__1981_ gnd vdd FILL
XFILL_0__3193_ gnd vdd FILL
XFILL_0__2144_ gnd vdd FILL
XFILL_8__1848_ gnd vdd FILL
X_2772_ _3297_/D _2772_/B _2772_/C _2773_/C vdd gnd AOI21X1
XFILL_0__2075_ gnd vdd FILL
X_1723_ _2594_/A _1783_/B _1846_/B vdd gnd NOR2X1
XFILL_8__3518_ gnd vdd FILL
XFILL_9__2311_ gnd vdd FILL
XFILL_6__2602_ gnd vdd FILL
XFILL_6__3582_ gnd vdd FILL
XFILL_8__1779_ gnd vdd FILL
XFILL_3__2824_ gnd vdd FILL
XFILL_6__2533_ gnd vdd FILL
XFILL_8__3449_ gnd vdd FILL
XFILL_3__2755_ gnd vdd FILL
X_3324_ _3324_/D vdd _3345_/R _3577_/CLK _3324_/Q vdd gnd DFFSR
XFILL_0__2977_ gnd vdd FILL
XFILL_1__1770_ gnd vdd FILL
XFILL_3__1706_ gnd vdd FILL
XFILL_6__2464_ gnd vdd FILL
XFILL_0__1928_ gnd vdd FILL
XFILL_6__2395_ gnd vdd FILL
X_3255_ NMI vdd _3363_/R _3363_/CLK _3255_/Q vdd gnd DFFSR
XFILL_3__2686_ gnd vdd FILL
XFILL_1__3440_ gnd vdd FILL
X_2206_ _2206_/A _3257_/Q _2235_/C vdd gnd XOR2X1
XFILL_0__1859_ gnd vdd FILL
X_3186_ _3186_/A _3186_/B _3186_/C _3196_/D vdd gnd OAI21X1
XFILL_4__3080_ gnd vdd FILL
XFILL_1__3371_ gnd vdd FILL
X_2137_ _2342_/A _2279_/A _2137_/C _2144_/B vdd gnd OAI21X1
XFILL_4__2100_ gnd vdd FILL
XFILL_0__3529_ gnd vdd FILL
XFILL_6__3016_ gnd vdd FILL
XFILL_1__2322_ gnd vdd FILL
XFILL_4__2031_ gnd vdd FILL
X_2068_ _2242_/A _2240_/B _2068_/C _2329_/B vdd gnd OAI21X1
XFILL_1__2253_ gnd vdd FILL
XFILL_3__3169_ gnd vdd FILL
XFILL_1__2184_ gnd vdd FILL
XFILL_7__2711_ gnd vdd FILL
XFILL_4__2933_ gnd vdd FILL
XFILL_7__2642_ gnd vdd FILL
XFILL_4__2864_ gnd vdd FILL
XFILL_4__2795_ gnd vdd FILL
XFILL_7__2573_ gnd vdd FILL
XFILL_4__1815_ gnd vdd FILL
XFILL_4__1746_ gnd vdd FILL
XFILL_1__1968_ gnd vdd FILL
XFILL_2__2500_ gnd vdd FILL
XFILL_2__3480_ gnd vdd FILL
XFILL_7__3125_ gnd vdd FILL
XFILL_4__3416_ gnd vdd FILL
XFILL_1__1899_ gnd vdd FILL
XFILL_5__2140_ gnd vdd FILL
XFILL_2__2431_ gnd vdd FILL
XFILL_2__2362_ gnd vdd FILL
XFILL_7__3056_ gnd vdd FILL
XFILL_5__2071_ gnd vdd FILL
XFILL_7__2007_ gnd vdd FILL
XFILL_8__2820_ gnd vdd FILL
XFILL_4__2229_ gnd vdd FILL
XFILL_2__2293_ gnd vdd FILL
XFILL_5_BUFX2_insert18 gnd vdd FILL
XFILL_8__2751_ gnd vdd FILL
XFILL_7__2909_ gnd vdd FILL
XFILL_5__2973_ gnd vdd FILL
XFILL_8__1702_ gnd vdd FILL
XFILL_8__2682_ gnd vdd FILL
XFILL_5__1924_ gnd vdd FILL
XFILL_5__1855_ gnd vdd FILL
XFILL_0__2900_ gnd vdd FILL
XFILL_5__1786_ gnd vdd FILL
XFILL_5__3525_ gnd vdd FILL
XFILL_0__2831_ gnd vdd FILL
XFILL_3__2540_ gnd vdd FILL
XFILL_5__3456_ gnd vdd FILL
XFILL_0__2762_ gnd vdd FILL
XFILL_6__2180_ gnd vdd FILL
XFILL_3__2471_ gnd vdd FILL
XFILL_0__1713_ gnd vdd FILL
XFILL_8__3165_ gnd vdd FILL
XFILL_5__2407_ gnd vdd FILL
XFILL_8__3096_ gnd vdd FILL
XFILL_5__3387_ gnd vdd FILL
X_3040_ _3050_/B _3041_/B vdd gnd INVX1
XFILL_8__2116_ gnd vdd FILL
XFILL_0__2693_ gnd vdd FILL
XFILL_2__2629_ gnd vdd FILL
XFILL_5__2338_ gnd vdd FILL
XFILL_8__2047_ gnd vdd FILL
XFILL_5__2269_ gnd vdd FILL
XFILL_3__3023_ gnd vdd FILL
XFILL181950x7950 gnd vdd FILL
XFILL_8__2949_ gnd vdd FILL
X_2824_ _2824_/A _2824_/B _2835_/B vdd gnd NOR2X1
XFILL_6__1964_ gnd vdd FILL
XFILL_0__3176_ gnd vdd FILL
XFILL182550x35250 gnd vdd FILL
XFILL184050x163950 gnd vdd FILL
XFILL_0__2127_ gnd vdd FILL
X_2755_ _3251_/Q _2756_/B _2757_/B vdd gnd NAND2X1
XFILL_6__1895_ gnd vdd FILL
XFILL_1__2940_ gnd vdd FILL
X_1706_ _2952_/A _3295_/D vdd gnd INVX1
XFILL_0__2058_ gnd vdd FILL
X_2686_ _2686_/A _2686_/B _2686_/C _2686_/D _2687_/B vdd gnd AOI22X1
XFILL_3__2807_ gnd vdd FILL
XFILL_1__2871_ gnd vdd FILL
XFILL_6__3565_ gnd vdd FILL
XFILL_6__3496_ gnd vdd FILL
XFILL_4__2580_ gnd vdd FILL
XFILL_6__2516_ gnd vdd FILL
XFILL_1__1822_ gnd vdd FILL
X_3307_ _3307_/D vdd _3346_/R _3307_/CLK _3307_/Q vdd gnd DFFSR
XFILL_6__2447_ gnd vdd FILL
XFILL_3__2738_ gnd vdd FILL
XFILL_1__1753_ gnd vdd FILL
XFILL_3__2669_ gnd vdd FILL
X_3238_ _3238_/D vdd _3313_/R _3284_/CLK _3238_/Q vdd gnd DFFSR
XFILL_6__2378_ gnd vdd FILL
XFILL_4__3201_ gnd vdd FILL
XFILL_4__3132_ gnd vdd FILL
XFILL_1__3423_ gnd vdd FILL
X_3169_ _3169_/A _3169_/B _3169_/C _3170_/A vdd gnd NAND3X1
XFILL_1__2305_ gnd vdd FILL
XFILL_4__3063_ gnd vdd FILL
XFILL_4__2014_ gnd vdd FILL
XFILL_1__2236_ gnd vdd FILL
XFILL_1__2167_ gnd vdd FILL
XFILL_4__2916_ gnd vdd FILL
XFILL_2__2980_ gnd vdd FILL
XFILL_1__2098_ gnd vdd FILL
XFILL_3_BUFX2_insert2 gnd vdd FILL
XFILL_2__1931_ gnd vdd FILL
XFILL_7__2625_ gnd vdd FILL
XFILL_2__1862_ gnd vdd FILL
XFILL_4__2847_ gnd vdd FILL
XFILL_7__2556_ gnd vdd FILL
XFILL_2__3601_ gnd vdd FILL
XFILL_4__2778_ gnd vdd FILL
XFILL_7__2487_ gnd vdd FILL
XFILL_4__1729_ gnd vdd FILL
XFILL_2__1793_ gnd vdd FILL
XFILL_2__3532_ gnd vdd FILL
XFILL_2__3463_ gnd vdd FILL
XFILL_7__3108_ gnd vdd FILL
XFILL_2__2414_ gnd vdd FILL
XFILL_5__3172_ gnd vdd FILL
XFILL_7__3039_ gnd vdd FILL
XFILL_2__3394_ gnd vdd FILL
XFILL_5__2123_ gnd vdd FILL
XFILL_5__2054_ gnd vdd FILL
XFILL_2__2345_ gnd vdd FILL
XFILL_2__2276_ gnd vdd FILL
XFILL_8__2803_ gnd vdd FILL
XFILL_0__3030_ gnd vdd FILL
XFILL_8__2734_ gnd vdd FILL
XFILL_5__2956_ gnd vdd FILL
XFILL_5__1907_ gnd vdd FILL
XFILL_3__1971_ gnd vdd FILL
XFILL_8__2665_ gnd vdd FILL
XFILL_5__2887_ gnd vdd FILL
X_2540_ _2540_/A _2540_/B _2541_/C vdd gnd AND2X2
XFILL_8__2596_ gnd vdd FILL
XFILL_5__1838_ gnd vdd FILL
X_2471_ _3292_/D _2502_/B _2502_/C _3350_/Q _2472_/B vdd gnd AOI22X1
XFILL_5__1769_ gnd vdd FILL
XFILL_5__3508_ gnd vdd FILL
XFILL_6__2301_ gnd vdd FILL
XFILL_1_BUFX2_insert16 gnd vdd FILL
XFILL_1_BUFX2_insert49 gnd vdd FILL
XFILL_0__2814_ gnd vdd FILL
XFILL_6_BUFX2_insert6 gnd vdd FILL
XFILL183450x150 gnd vdd FILL
XFILL_8__3217_ gnd vdd FILL
XFILL_1_BUFX2_insert27 gnd vdd FILL
XFILL_3__2523_ gnd vdd FILL
XFILL_5__3439_ gnd vdd FILL
XFILL_3__2454_ gnd vdd FILL
XFILL_0__2745_ gnd vdd FILL
XFILL_8__3148_ gnd vdd FILL
XFILL_6__2232_ gnd vdd FILL
XFILL_6__2163_ gnd vdd FILL
X_3023_ _3023_/A _3023_/B _3027_/A vdd gnd NOR2X1
XFILL_0__2676_ gnd vdd FILL
XFILL_8__3079_ gnd vdd FILL
XFILL_3__2385_ gnd vdd FILL
XFILL_6__2094_ gnd vdd FILL
XFILL_1_CLKBUF1_insert28 gnd vdd FILL
XFILL184350x167850 gnd vdd FILL
XFILL184050x175650 gnd vdd FILL
XFILL_3__3006_ gnd vdd FILL
XFILL_1__3070_ gnd vdd FILL
XFILL_1__2021_ gnd vdd FILL
XFILL_0__3228_ gnd vdd FILL
XFILL_6__2996_ gnd vdd FILL
XFILL_6__1947_ gnd vdd FILL
X_2807_ _2813_/C _2809_/C _2807_/C _3264_/D vdd gnd OAI21X1
XFILL_0__3159_ gnd vdd FILL
XFILL_6__1878_ gnd vdd FILL
XFILL_4__2701_ gnd vdd FILL
X_2738_ _2738_/A _2738_/B _2739_/C vdd gnd OR2X2
XFILL_1__2923_ gnd vdd FILL
XFILL_7__3390_ gnd vdd FILL
XFILL_7__2410_ gnd vdd FILL
XFILL_6__3548_ gnd vdd FILL
XFILL_7__2341_ gnd vdd FILL
XFILL_4__2632_ gnd vdd FILL
X_2669_ _2669_/A _2748_/B _2669_/C _2670_/C vdd gnd OAI21X1
XFILL_1__2854_ gnd vdd FILL
XFILL_4__2563_ gnd vdd FILL
XFILL_6__3479_ gnd vdd FILL
XFILL_7__2272_ gnd vdd FILL
XFILL_1__2785_ gnd vdd FILL
XFILL_9__2208_ gnd vdd FILL
XFILL_1__1805_ gnd vdd FILL
XFILL_4__2494_ gnd vdd FILL
XFILL_1__1736_ gnd vdd FILL
XFILL_4__3115_ gnd vdd FILL
XFILL_1__3406_ gnd vdd FILL
XFILL_4__3046_ gnd vdd FILL
XFILL_2__2130_ gnd vdd FILL
XFILL184050x54750 gnd vdd FILL
XFILL_2__2061_ gnd vdd FILL
XFILL_1__2219_ gnd vdd FILL
XFILL_5__2810_ gnd vdd FILL
XFILL_7__1987_ gnd vdd FILL
XFILL_1__3199_ gnd vdd FILL
XBUFX2_insert41 _1734_/Y _2292_/B vdd gnd BUFX2
XBUFX2_insert63 _1993_/Y _2898_/B vdd gnd BUFX2
XBUFX2_insert74 _1694_/Y _2298_/A vdd gnd BUFX2
XFILL_8__2450_ gnd vdd FILL
XFILL_5__2741_ gnd vdd FILL
XBUFX2_insert52 _1733_/Y _2379_/A vdd gnd BUFX2
XBUFX2_insert96 _2083_/Y _2919_/B vdd gnd BUFX2
XBUFX2_insert85 _1858_/Y _2906_/B vdd gnd BUFX2
XFILL_2__2963_ gnd vdd FILL
XFILL_5__2672_ gnd vdd FILL
XFILL_7__2608_ gnd vdd FILL
XFILL_2__2894_ gnd vdd FILL
XFILL_8__2381_ gnd vdd FILL
XFILL_2__1914_ gnd vdd FILL
XFILL_7__3588_ gnd vdd FILL
XFILL_2__1845_ gnd vdd FILL
XFILL_7__2539_ gnd vdd FILL
XFILL_8_BUFX2_insert22 gnd vdd FILL
XFILL_8_BUFX2_insert11 gnd vdd FILL
XFILL_2__1776_ gnd vdd FILL
XFILL_2__3515_ gnd vdd FILL
XFILL_8__3002_ gnd vdd FILL
XFILL_8_BUFX2_insert66 gnd vdd FILL
XFILL_8_BUFX2_insert44 gnd vdd FILL
XFILL_8_BUFX2_insert55 gnd vdd FILL
XFILL_8_BUFX2_insert88 gnd vdd FILL
XFILL_0__2530_ gnd vdd FILL
XFILL_5__3224_ gnd vdd FILL
XFILL_8_BUFX2_insert77 gnd vdd FILL
XFILL_2__3446_ gnd vdd FILL
XFILL_5__3155_ gnd vdd FILL
XFILL_2__3377_ gnd vdd FILL
XFILL_3__2170_ gnd vdd FILL
XFILL_0__2461_ gnd vdd FILL
XFILL_5__2106_ gnd vdd FILL
XFILL_5__3086_ gnd vdd FILL
XFILL_2__2328_ gnd vdd FILL
XFILL_0__2392_ gnd vdd FILL
XFILL_5__2037_ gnd vdd FILL
XFILL_6__2850_ gnd vdd FILL
XFILL_2__2259_ gnd vdd FILL
X_1971_ _3230_/A _2700_/B _2760_/B vdd gnd NOR2X1
XFILL_0__3013_ gnd vdd FILL
XFILL_6__1801_ gnd vdd FILL
XFILL_6__2781_ gnd vdd FILL
XFILL_8__2717_ gnd vdd FILL
X_3572_ _3572_/D vdd _3578_/R _3573_/CLK _3572_/Q vdd gnd DFFSR
XFILL_5__2939_ gnd vdd FILL
XFILL_6__1732_ gnd vdd FILL
XFILL_8__2648_ gnd vdd FILL
XFILL_3__1954_ gnd vdd FILL
X_2523_ _2523_/A _2523_/B _2523_/C _3216_/B vdd gnd NAND3X1
XFILL_8__2579_ gnd vdd FILL
XFILL_6__3402_ gnd vdd FILL
XFILL_3__1885_ gnd vdd FILL
X_2454_ _2502_/B _2510_/B vdd gnd INVX1
X_2385_ _3570_/Q _2427_/B _2385_/C _2386_/B vdd gnd AOI21X1
XFILL_3__3555_ gnd vdd FILL
XFILL_1__2570_ gnd vdd FILL
XFILL_3__3486_ gnd vdd FILL
XFILL_6__2215_ gnd vdd FILL
XFILL_3__2506_ gnd vdd FILL
XFILL184350x179550 gnd vdd FILL
XFILL_6__3195_ gnd vdd FILL
XFILL_0__2728_ gnd vdd FILL
XFILL_3__2437_ gnd vdd FILL
X_3006_ _3282_/Q _3006_/B _3010_/C vdd gnd NOR2X1
XFILL_6__2146_ gnd vdd FILL
XFILL_3__2368_ gnd vdd FILL
XFILL_0__2659_ gnd vdd FILL
XFILL_6__2077_ gnd vdd FILL
XFILL_1__3122_ gnd vdd FILL
XFILL_3__2299_ gnd vdd FILL
XFILL_7__1910_ gnd vdd FILL
XFILL_7__2890_ gnd vdd FILL
XFILL_9__2826_ gnd vdd FILL
XFILL_1__3053_ gnd vdd FILL
XFILL_7__1841_ gnd vdd FILL
XFILL_1__2004_ gnd vdd FILL
XFILL_6__2979_ gnd vdd FILL
XFILL_7__1772_ gnd vdd FILL
XFILL_7__3511_ gnd vdd FILL
XFILL_4__1994_ gnd vdd FILL
XFILL_7__3442_ gnd vdd FILL
XFILL_7__3373_ gnd vdd FILL
XFILL_1__2906_ gnd vdd FILL
XFILL_4__2615_ gnd vdd FILL
XFILL_1__2837_ gnd vdd FILL
XFILL_7__2324_ gnd vdd FILL
XFILL_4__3595_ gnd vdd FILL
XFILL_7__2255_ gnd vdd FILL
XFILL_4__2546_ gnd vdd FILL
XFILL_1__2768_ gnd vdd FILL
XFILL_4__2477_ gnd vdd FILL
XFILL_7__2186_ gnd vdd FILL
XFILL181050x74250 gnd vdd FILL
XFILL_1__1719_ gnd vdd FILL
XFILL_1__2699_ gnd vdd FILL
XFILL_2__3231_ gnd vdd FILL
XFILL_8__1950_ gnd vdd FILL
XFILL_2__3162_ gnd vdd FILL
XFILL_2__2113_ gnd vdd FILL
XFILL_4__3029_ gnd vdd FILL
XFILL_2__3093_ gnd vdd FILL
XFILL_8__1881_ gnd vdd FILL
XFILL_2__2044_ gnd vdd FILL
XFILL_8__3551_ gnd vdd FILL
XFILL_8__2502_ gnd vdd FILL
XFILL_8__3482_ gnd vdd FILL
XFILL_5__2724_ gnd vdd FILL
XFILL_2__2946_ gnd vdd FILL
XFILL_8__2433_ gnd vdd FILL
XFILL_8__2364_ gnd vdd FILL
XFILL_0__1961_ gnd vdd FILL
XFILL_5__2655_ gnd vdd FILL
XFILL_2__2877_ gnd vdd FILL
XFILL_0__1892_ gnd vdd FILL
XFILL_5__2586_ gnd vdd FILL
XFILL_8__2295_ gnd vdd FILL
XFILL_2__1828_ gnd vdd FILL
X_2170_ _2823_/B _2875_/A _2297_/A vdd gnd NAND2X1
XFILL_2__1759_ gnd vdd FILL
XFILL_6__2000_ gnd vdd FILL
XFILL_0__3562_ gnd vdd FILL
XFILL_5__3207_ gnd vdd FILL
XFILL_0__3493_ gnd vdd FILL
XFILL_2__3429_ gnd vdd FILL
XFILL_3__2222_ gnd vdd FILL
XFILL_0__2513_ gnd vdd FILL
XFILL_5__3138_ gnd vdd FILL
XFILL_0__2444_ gnd vdd FILL
XFILL_5__3069_ gnd vdd FILL
XFILL_3__2153_ gnd vdd FILL
XFILL_6__2902_ gnd vdd FILL
XFILL_3__2084_ gnd vdd FILL
XFILL_0__2375_ gnd vdd FILL
X_1954_ _1985_/A _3574_/Q _1954_/C _1955_/C vdd gnd AOI21X1
XFILL_4_BUFX2_insert20 gnd vdd FILL
XFILL_6__2833_ gnd vdd FILL
XFILL_4_BUFX2_insert42 gnd vdd FILL
XFILL_4_BUFX2_insert64 gnd vdd FILL
X_1885_ _1885_/A _2240_/B vdd gnd INVX1
XFILL_6__2764_ gnd vdd FILL
XFILL_4_BUFX2_insert75 gnd vdd FILL
XFILL_4_BUFX2_insert53 gnd vdd FILL
XFILL_4_BUFX2_insert97 gnd vdd FILL
XFILL_3__2986_ gnd vdd FILL
XFILL_9__2473_ gnd vdd FILL
XFILL_6__1715_ gnd vdd FILL
XFILL_4_BUFX2_insert86 gnd vdd FILL
X_3555_ _3555_/A _3555_/B _3566_/A _3556_/B vdd gnd OAI21X1
XFILL_3__1937_ gnd vdd FILL
XFILL_6__2695_ gnd vdd FILL
X_3486_ _3543_/C _3545_/A vdd gnd INVX1
X_2506_ _2506_/A _2519_/C _2506_/C _3213_/B vdd gnd AOI21X1
XFILL_3__1868_ gnd vdd FILL
X_2437_ _2437_/A _3158_/B _2437_/C _2438_/B vdd gnd NAND3X1
XFILL_4__3380_ gnd vdd FILL
XFILL_4__2400_ gnd vdd FILL
XFILL_3__1799_ gnd vdd FILL
XFILL_3__3538_ gnd vdd FILL
XFILL_4__2331_ gnd vdd FILL
X_2368_ _3063_/B _2429_/A _2426_/B _2373_/B vdd gnd NAND3X1
XFILL_1__2622_ gnd vdd FILL
XFILL_7__2040_ gnd vdd FILL
XFILL_4__2262_ gnd vdd FILL
X_2299_ _2299_/A _3145_/B _2341_/A _2300_/C vdd gnd OAI21X1
XFILL_1__2553_ gnd vdd FILL
XFILL_3__3469_ gnd vdd FILL
XFILL_1__2484_ gnd vdd FILL
XFILL_6__3178_ gnd vdd FILL
XFILL_4__2193_ gnd vdd FILL
XFILL_6__2129_ gnd vdd FILL
XFILL_7__2942_ gnd vdd FILL
XFILL_1__3105_ gnd vdd FILL
XFILL_7__2873_ gnd vdd FILL
XFILL_1__3036_ gnd vdd FILL
XFILL_7__1824_ gnd vdd FILL
XFILL184350x43050 gnd vdd FILL
XFILL_7__1755_ gnd vdd FILL
XFILL_4__1977_ gnd vdd FILL
XFILL_2__2800_ gnd vdd FILL
XFILL_7__3425_ gnd vdd FILL
XFILL_2__2731_ gnd vdd FILL
XFILL_5__2440_ gnd vdd FILL
XFILL_5__2371_ gnd vdd FILL
XFILL_7__2307_ gnd vdd FILL
XFILL_2__2662_ gnd vdd FILL
XFILL_8__2080_ gnd vdd FILL
XFILL_4__2529_ gnd vdd FILL
XFILL_2__2593_ gnd vdd FILL
XFILL_7__2238_ gnd vdd FILL
XFILL_7__2169_ gnd vdd FILL
XFILL_8__2982_ gnd vdd FILL
XFILL_2__3214_ gnd vdd FILL
XFILL_8__1933_ gnd vdd FILL
XFILL_2__3145_ gnd vdd FILL
XFILL_0__2160_ gnd vdd FILL
XFILL_2__3076_ gnd vdd FILL
XFILL_8__1864_ gnd vdd FILL
XFILL_2__2027_ gnd vdd FILL
XFILL_8__3603_ gnd vdd FILL
XFILL_0__2091_ gnd vdd FILL
XFILL_8__1795_ gnd vdd FILL
XFILL_3__2840_ gnd vdd FILL
XFILL_8__3534_ gnd vdd FILL
XFILL_8__3465_ gnd vdd FILL
X_3340_ _3340_/D vdd _3346_/R _3346_/CLK _3340_/Q vdd gnd DFFSR
XFILL_8__2416_ gnd vdd FILL
XFILL_5__2707_ gnd vdd FILL
XFILL_3__2771_ gnd vdd FILL
XFILL_6__2480_ gnd vdd FILL
XFILL_2__2929_ gnd vdd FILL
XFILL_8__3396_ gnd vdd FILL
XFILL_0__2993_ gnd vdd FILL
XFILL_3__1722_ gnd vdd FILL
XFILL_5__2638_ gnd vdd FILL
X_3271_ _3271_/D vdd _3289_/R _3307_/CLK _3271_/Q vdd gnd DFFSR
XFILL_8__2347_ gnd vdd FILL
XFILL_0__1944_ gnd vdd FILL
XFILL_0__1875_ gnd vdd FILL
XFILL_6__3101_ gnd vdd FILL
XFILL_8__2278_ gnd vdd FILL
X_2222_ _2294_/A _3177_/B _2223_/C _2320_/B vdd gnd OAI21X1
XFILL_5__2569_ gnd vdd FILL
XFILL_6_CLKBUF1_insert28 gnd vdd FILL
X_2153_ _2341_/A _2167_/A _2153_/C _2347_/C vdd gnd OAI21X1
XFILL_0__3545_ gnd vdd FILL
XFILL_6__3032_ gnd vdd FILL
X_2084_ _2932_/B _2894_/A vdd gnd INVX2
XFILL_0__3476_ gnd vdd FILL
XFILL_3__2205_ gnd vdd FILL
XFILL_3__3185_ gnd vdd FILL
XFILL_0__2427_ gnd vdd FILL
XFILL_3__2136_ gnd vdd FILL
XFILL_4_CLKBUF1_insert32 gnd vdd FILL
XFILL_0__2358_ gnd vdd FILL
X_2986_ _2986_/A _2986_/B _2986_/C _2988_/B vdd gnd AOI21X1
XFILL_3__2067_ gnd vdd FILL
XFILL_4__2880_ gnd vdd FILL
XFILL_6__2816_ gnd vdd FILL
X_1937_ _1986_/A _1937_/B _1937_/C _3438_/A vdd gnd OAI21X1
XFILL_4__1900_ gnd vdd FILL
XFILL_0__2289_ gnd vdd FILL
X_1868_ _1879_/C _1878_/B _3127_/B vdd gnd NOR2X1
XFILL_4__1831_ gnd vdd FILL
XFILL_6__2747_ gnd vdd FILL
X_3538_ _3562_/B _3538_/B _3553_/B _3539_/C vdd gnd AOI21X1
XFILL_3__2969_ gnd vdd FILL
X_1799_ _2299_/A _3147_/B _3148_/B vdd gnd NOR2X1
XFILL_6__2678_ gnd vdd FILL
XFILL_4__1762_ gnd vdd FILL
XFILL_4__3501_ gnd vdd FILL
XFILL_1__1984_ gnd vdd FILL
XFILL_7__3210_ gnd vdd FILL
XFILL_4__1693_ gnd vdd FILL
X_3469_ _3484_/B _3469_/B _3470_/A vdd gnd NAND2X1
XFILL_4__3432_ gnd vdd FILL
XFILL_7__3141_ gnd vdd FILL
XFILL_7__3072_ gnd vdd FILL
XFILL_1__2605_ gnd vdd FILL
XFILL_0_BUFX2_insert51 gnd vdd FILL
XFILL_7__2023_ gnd vdd FILL
XFILL_0_BUFX2_insert40 gnd vdd FILL
XFILL_4__2314_ gnd vdd FILL
XFILL_1__3585_ gnd vdd FILL
XFILL_0_BUFX2_insert84 gnd vdd FILL
XFILL_0_BUFX2_insert62 gnd vdd FILL
XFILL_0_BUFX2_insert73 gnd vdd FILL
XFILL_4__2245_ gnd vdd FILL
XFILL_1__2536_ gnd vdd FILL
XFILL_0_BUFX2_insert95 gnd vdd FILL
XFILL_1__2467_ gnd vdd FILL
XFILL_1__2398_ gnd vdd FILL
XFILL_4__2176_ gnd vdd FILL
XFILL_7__2925_ gnd vdd FILL
XFILL_5__1940_ gnd vdd FILL
XFILL_7__2856_ gnd vdd FILL
XFILL_5__1871_ gnd vdd FILL
XFILL_1__3019_ gnd vdd FILL
XFILL_7__2787_ gnd vdd FILL
XFILL_7__1807_ gnd vdd FILL
XFILL_7__1738_ gnd vdd FILL
XFILL_5__3541_ gnd vdd FILL
XFILL_5__3472_ gnd vdd FILL
XFILL_7__3408_ gnd vdd FILL
XFILL_8__2201_ gnd vdd FILL
XFILL_5__2423_ gnd vdd FILL
XFILL_2__2714_ gnd vdd FILL
XFILL_8__3181_ gnd vdd FILL
XFILL_8__2132_ gnd vdd FILL
XFILL_2__2645_ gnd vdd FILL
XFILL_5__2354_ gnd vdd FILL
XFILL_8__2063_ gnd vdd FILL
XFILL_2__2576_ gnd vdd FILL
XFILL_5__2285_ gnd vdd FILL
XFILL_8__2965_ gnd vdd FILL
X_2840_ _2921_/A _2867_/A _2933_/B _2841_/D vdd gnd OAI21X1
XFILL_8__1916_ gnd vdd FILL
XFILL_6__1980_ gnd vdd FILL
XFILL_0__2212_ gnd vdd FILL
XFILL_0__3192_ gnd vdd FILL
XFILL_2__3128_ gnd vdd FILL
XFILL_8__2896_ gnd vdd FILL
XFILL_0__2143_ gnd vdd FILL
XFILL_2__3059_ gnd vdd FILL
XFILL_8__1847_ gnd vdd FILL
X_2771_ _2771_/A _2771_/B _2771_/C _2772_/C vdd gnd NAND3X1
XFILL_0__2074_ gnd vdd FILL
XFILL_8__1778_ gnd vdd FILL
X_1722_ _3234_/Q _3233_/Q _2594_/A vdd gnd NAND2X1
XFILL_8__3517_ gnd vdd FILL
XFILL_6__3581_ gnd vdd FILL
XFILL_6__2601_ gnd vdd FILL
XFILL_3__2823_ gnd vdd FILL
XFILL_6__2532_ gnd vdd FILL
XFILL_8__3448_ gnd vdd FILL
XFILL_3__2754_ gnd vdd FILL
X_3323_ _3323_/D vdd _3346_/R _3346_/CLK _3323_/Q vdd gnd DFFSR
XFILL_0__2976_ gnd vdd FILL
XFILL_8__3379_ gnd vdd FILL
XFILL_3__1705_ gnd vdd FILL
XFILL_6__2463_ gnd vdd FILL
XFILL_0__1927_ gnd vdd FILL
XFILL_6__2394_ gnd vdd FILL
X_3254_ _3254_/D vdd _3291_/R _3362_/CLK _3254_/Q vdd gnd DFFSR
XFILL_3__2685_ gnd vdd FILL
X_2205_ _3258_/Q _2205_/B _2205_/C _2206_/A vdd gnd OAI21X1
XFILL_0__1858_ gnd vdd FILL
X_3185_ _3185_/A _3185_/B _3185_/C _3186_/B vdd gnd NAND3X1
XFILL_6__3015_ gnd vdd FILL
XFILL_1__3370_ gnd vdd FILL
X_2136_ _2221_/A _3183_/B _2342_/A _2137_/C vdd gnd OAI21X1
XFILL_0__1789_ gnd vdd FILL
XFILL_7_BUFX2_insert90 gnd vdd FILL
XFILL_0__3528_ gnd vdd FILL
XFILL_4__2030_ gnd vdd FILL
XFILL_1__2321_ gnd vdd FILL
X_2067_ _2276_/A _3173_/B _2242_/A _2068_/C vdd gnd OAI21X1
XFILL_0__3459_ gnd vdd FILL
XFILL_1__2252_ gnd vdd FILL
XFILL_3__3168_ gnd vdd FILL
XFILL_3__3099_ gnd vdd FILL
XFILL_1__2183_ gnd vdd FILL
XFILL_3__2119_ gnd vdd FILL
XFILL_7__2710_ gnd vdd FILL
XFILL_4__2932_ gnd vdd FILL
X_2969_ _2969_/A _3372_/Y _2969_/C _2971_/B vdd gnd AOI21X1
XFILL_7__2641_ gnd vdd FILL
XFILL_4__2863_ gnd vdd FILL
XFILL_7__2572_ gnd vdd FILL
XFILL_4__2794_ gnd vdd FILL
XFILL_4__1814_ gnd vdd FILL
XFILL_4__1745_ gnd vdd FILL
XFILL_1__1967_ gnd vdd FILL
XFILL_7__3124_ gnd vdd FILL
XFILL_4__3415_ gnd vdd FILL
XFILL_1__1898_ gnd vdd FILL
XFILL_2__2430_ gnd vdd FILL
XFILL_2__2361_ gnd vdd FILL
XFILL_7__3055_ gnd vdd FILL
XFILL_7__2006_ gnd vdd FILL
XFILL_5__2070_ gnd vdd FILL
XFILL_1__2519_ gnd vdd FILL
XFILL_2__2292_ gnd vdd FILL
XFILL_1__3499_ gnd vdd FILL
XFILL_4__2228_ gnd vdd FILL
XFILL_4__2159_ gnd vdd FILL
XFILL_5_BUFX2_insert19 gnd vdd FILL
XFILL_8__2750_ gnd vdd FILL
XFILL_7__2908_ gnd vdd FILL
XFILL_5__2972_ gnd vdd FILL
XFILL_8__1701_ gnd vdd FILL
XFILL_8__2681_ gnd vdd FILL
XFILL_7__2839_ gnd vdd FILL
XFILL_5__1923_ gnd vdd FILL
XFILL_5__1854_ gnd vdd FILL
XFILL_5__3524_ gnd vdd FILL
XFILL_5__1785_ gnd vdd FILL
XFILL_0__2830_ gnd vdd FILL
XFILL_5__3455_ gnd vdd FILL
XFILL_0__2761_ gnd vdd FILL
XFILL_8__3164_ gnd vdd FILL
XFILL_5__3386_ gnd vdd FILL
XFILL_8__2115_ gnd vdd FILL
XFILL_3__2470_ gnd vdd FILL
XFILL_0__1712_ gnd vdd FILL
XFILL_5__2406_ gnd vdd FILL
XFILL_8__3095_ gnd vdd FILL
XFILL_5__2337_ gnd vdd FILL
XFILL_0__2692_ gnd vdd FILL
XFILL_2__2628_ gnd vdd FILL
XFILL_8__2046_ gnd vdd FILL
XFILL_2__2559_ gnd vdd FILL
XFILL_5__2268_ gnd vdd FILL
XFILL_9__1810_ gnd vdd FILL
XFILL_5__2199_ gnd vdd FILL
XFILL_3__3022_ gnd vdd FILL
XFILL_8__2948_ gnd vdd FILL
X_2823_ _2915_/A _2823_/B _2823_/C _2824_/B vdd gnd NAND3X1
XFILL_8__2879_ gnd vdd FILL
XFILL_6__1963_ gnd vdd FILL
XFILL_0__3175_ gnd vdd FILL
XFILL183750x160050 gnd vdd FILL
XFILL_0__2126_ gnd vdd FILL
X_2754_ _2778_/A _2754_/B _2754_/C _3252_/D vdd gnd OAI21X1
XFILL_6__1894_ gnd vdd FILL
X_1705_ _2768_/A DI[5] _1705_/C _2952_/A vdd gnd OAI21X1
XFILL_0__2057_ gnd vdd FILL
X_2685_ _3246_/Q _2685_/B _2686_/C vdd gnd NAND2X1
XFILL_1__2870_ gnd vdd FILL
XFILL_3__2806_ gnd vdd FILL
XFILL_6__3564_ gnd vdd FILL
XFILL_6__3495_ gnd vdd FILL
XFILL_1__1821_ gnd vdd FILL
XFILL_6__2515_ gnd vdd FILL
X_3306_ _3306_/D _3346_/CLK _3306_/Q vdd gnd DFFPOSX1
XFILL_6__2446_ gnd vdd FILL
XFILL_3__2737_ gnd vdd FILL
XFILL_0__2959_ gnd vdd FILL
XFILL_1__1752_ gnd vdd FILL
XFILL_3__2668_ gnd vdd FILL
X_3237_ _3237_/D vdd _3313_/R _3284_/CLK _3237_/Q vdd gnd DFFSR
XFILL_6__2377_ gnd vdd FILL
XFILL_4__3200_ gnd vdd FILL
XFILL_4__3131_ gnd vdd FILL
XFILL_1__3422_ gnd vdd FILL
XFILL_3__2599_ gnd vdd FILL
X_3168_ _3168_/A _3174_/A _3169_/B vdd gnd NOR2X1
X_2119_ _2298_/A _3171_/A _2191_/A _2288_/C _2344_/B vdd gnd AOI22X1
XFILL_4__3062_ gnd vdd FILL
X_3099_ _3121_/A _3107_/B _3326_/Q _3100_/C vdd gnd OAI21X1
XFILL_1__2304_ gnd vdd FILL
XFILL_4__2013_ gnd vdd FILL
XFILL_9__2988_ gnd vdd FILL
XFILL_1__2235_ gnd vdd FILL
XFILL_1__2166_ gnd vdd FILL
XFILL_4__2915_ gnd vdd FILL
XFILL_1__2097_ gnd vdd FILL
XFILL_3_BUFX2_insert3 gnd vdd FILL
XFILL_7__2624_ gnd vdd FILL
XFILL_4__2846_ gnd vdd FILL
XFILL_2__1930_ gnd vdd FILL
XFILL_2__1861_ gnd vdd FILL
XFILL_7__2555_ gnd vdd FILL
XFILL_2__3600_ gnd vdd FILL
XFILL_7__2486_ gnd vdd FILL
XFILL_4__2777_ gnd vdd FILL
XFILL_1__2999_ gnd vdd FILL
XFILL_2__1792_ gnd vdd FILL
XFILL_4__1728_ gnd vdd FILL
XFILL_2__3531_ gnd vdd FILL
XFILL182550x7950 gnd vdd FILL
XFILL_2__3462_ gnd vdd FILL
XFILL_7__3107_ gnd vdd FILL
XFILL_5__3171_ gnd vdd FILL
XFILL_2__2413_ gnd vdd FILL
XFILL_2__3393_ gnd vdd FILL
XFILL_7__3038_ gnd vdd FILL
XFILL_5__2122_ gnd vdd FILL
XFILL_2__2344_ gnd vdd FILL
XFILL_5__2053_ gnd vdd FILL
XFILL_2__2275_ gnd vdd FILL
XFILL_8__2802_ gnd vdd FILL
XFILL182250x109350 gnd vdd FILL
XFILL_8__2733_ gnd vdd FILL
XFILL_5__2955_ gnd vdd FILL
XFILL_3__1970_ gnd vdd FILL
XFILL_8__2664_ gnd vdd FILL
XFILL_5__1906_ gnd vdd FILL
XFILL_5__2886_ gnd vdd FILL
XFILL_8__2595_ gnd vdd FILL
X_2470_ _2508_/B _2511_/A _3572_/Q _2472_/A vdd gnd OAI21X1
XFILL_5__1837_ gnd vdd FILL
XFILL_5__1768_ gnd vdd FILL
XFILL_5__3507_ gnd vdd FILL
XFILL_0__2813_ gnd vdd FILL
XFILL_6__2300_ gnd vdd FILL
XFILL_8__3216_ gnd vdd FILL
XFILL_5__3438_ gnd vdd FILL
XFILL_1_BUFX2_insert17 gnd vdd FILL
XFILL_1_BUFX2_insert39 gnd vdd FILL
XFILL_6__2231_ gnd vdd FILL
XFILL_6_BUFX2_insert7 gnd vdd FILL
XFILL_5__1699_ gnd vdd FILL
XFILL_3__2522_ gnd vdd FILL
XFILL_3__2453_ gnd vdd FILL
XFILL_8__3147_ gnd vdd FILL
XFILL_0__2744_ gnd vdd FILL
XFILL_6__2162_ gnd vdd FILL
XFILL_8__3078_ gnd vdd FILL
XFILL_5__3369_ gnd vdd FILL
X_3022_ _3022_/A _3022_/B _3022_/C _3314_/D vdd gnd OAI21X1
XFILL_0__2675_ gnd vdd FILL
XFILL_8__2029_ gnd vdd FILL
XFILL_3__2384_ gnd vdd FILL
XFILL_6__2093_ gnd vdd FILL
XFILL_1_CLKBUF1_insert29 gnd vdd FILL
XFILL_3__3005_ gnd vdd FILL
XFILL_1__2020_ gnd vdd FILL
XFILL_6__2995_ gnd vdd FILL
XFILL_0__3227_ gnd vdd FILL
XFILL_6__1946_ gnd vdd FILL
X_2806_ _2851_/A _2881_/A _2809_/C vdd gnd NAND2X1
XFILL_0__3158_ gnd vdd FILL
XFILL_0__3089_ gnd vdd FILL
XFILL_6__1877_ gnd vdd FILL
XFILL_4__2700_ gnd vdd FILL
X_2737_ _3226_/A _2748_/B _2737_/C _2738_/A vdd gnd OAI21X1
XFILL_0__2109_ gnd vdd FILL
XFILL_1__2922_ gnd vdd FILL
X_2668_ _2675_/A _2668_/B _2668_/C _2668_/D _3245_/D vdd gnd OAI22X1
XFILL_6__3547_ gnd vdd FILL
XFILL_7__2340_ gnd vdd FILL
XFILL_4__2631_ gnd vdd FILL
XFILL_1__2853_ gnd vdd FILL
X_2599_ _2599_/A _2599_/B _2751_/B _2601_/A vdd gnd NAND3X1
XFILL_4__2562_ gnd vdd FILL
XFILL_6__3478_ gnd vdd FILL
XFILL_1__2784_ gnd vdd FILL
XFILL_7__2271_ gnd vdd FILL
XFILL_1__1804_ gnd vdd FILL
XFILL_4__2493_ gnd vdd FILL
XFILL_1__1735_ gnd vdd FILL
XFILL_6__2429_ gnd vdd FILL
XFILL_1__3405_ gnd vdd FILL
XFILL_4__3114_ gnd vdd FILL
XFILL_4__3045_ gnd vdd FILL
XFILL_2__2060_ gnd vdd FILL
XFILL_1__2218_ gnd vdd FILL
XFILL_7__1986_ gnd vdd FILL
XFILL_1__3198_ gnd vdd FILL
XBUFX2_insert20 _2580_/Y _3289_/R vdd gnd BUFX2
XFILL_1__2149_ gnd vdd FILL
XBUFX2_insert42 _1734_/Y _3024_/A vdd gnd BUFX2
XFILL_5__2740_ gnd vdd FILL
XBUFX2_insert64 _1993_/Y _2887_/A vdd gnd BUFX2
XFILL_2__2962_ gnd vdd FILL
XBUFX2_insert75 _1694_/Y _2778_/A vdd gnd BUFX2
XBUFX2_insert53 _1733_/Y _3160_/A vdd gnd BUFX2
XBUFX2_insert97 _2083_/Y _2936_/B vdd gnd BUFX2
XFILL_7__3587_ gnd vdd FILL
XFILL_8__2380_ gnd vdd FILL
XFILL_2__1913_ gnd vdd FILL
XFILL_7__2607_ gnd vdd FILL
XFILL_5__2671_ gnd vdd FILL
XBUFX2_insert86 _1729_/Y _3147_/A vdd gnd BUFX2
XFILL_4__2829_ gnd vdd FILL
XFILL_2__2893_ gnd vdd FILL
XFILL_7__2538_ gnd vdd FILL
XFILL_2__1844_ gnd vdd FILL
XFILL_8_BUFX2_insert23 gnd vdd FILL
XFILL_8_BUFX2_insert12 gnd vdd FILL
XFILL_7__2469_ gnd vdd FILL
XFILL_2__1775_ gnd vdd FILL
XFILL_2__3514_ gnd vdd FILL
XFILL_8_BUFX2_insert56 gnd vdd FILL
XFILL_8__3001_ gnd vdd FILL
XFILL_8_BUFX2_insert45 gnd vdd FILL
XFILL_8_BUFX2_insert67 gnd vdd FILL
XFILL_8_BUFX2_insert78 gnd vdd FILL
XFILL_5__3223_ gnd vdd FILL
XFILL_8_BUFX2_insert89 gnd vdd FILL
XFILL_2__3445_ gnd vdd FILL
XFILL_5__3154_ gnd vdd FILL
XFILL_2__3376_ gnd vdd FILL
XFILL_0__2460_ gnd vdd FILL
XFILL_5__2105_ gnd vdd FILL
XFILL_2__2327_ gnd vdd FILL
XFILL_5__3085_ gnd vdd FILL
XFILL_0__2391_ gnd vdd FILL
XFILL_5__2036_ gnd vdd FILL
X_1970_ _3362_/Q _3230_/A vdd gnd INVX1
XFILL_2__2258_ gnd vdd FILL
XFILL_2__2189_ gnd vdd FILL
XFILL_0__3012_ gnd vdd FILL
XFILL_6__1800_ gnd vdd FILL
XFILL_8__2716_ gnd vdd FILL
XFILL_6__2780_ gnd vdd FILL
X_3571_ _3571_/D vdd _3578_/R _3573_/CLK _3571_/Q vdd gnd DFFSR
XFILL_5__2938_ gnd vdd FILL
XFILL_6__1731_ gnd vdd FILL
XFILL_8__2647_ gnd vdd FILL
XFILL_5__2869_ gnd vdd FILL
XFILL_3__1953_ gnd vdd FILL
X_2522_ _2565_/A _3290_/D _2522_/C _2523_/C vdd gnd AOI21X1
XFILL_8__2578_ gnd vdd FILL
XFILL_6__3401_ gnd vdd FILL
XFILL_3__1884_ gnd vdd FILL
X_2453_ _2453_/A _3183_/B _3156_/C _2502_/B vdd gnd OAI21X1
XFILL_3__3554_ gnd vdd FILL
X_2384_ _2612_/B _2426_/B _2384_/C _2385_/C vdd gnd OAI21X1
XFILL_3__2505_ gnd vdd FILL
XFILL_3__3485_ gnd vdd FILL
XFILL_6__2214_ gnd vdd FILL
XFILL_6__3194_ gnd vdd FILL
XFILL_0__2727_ gnd vdd FILL
X_3005_ _3005_/A _3005_/B _3005_/C _3312_/D vdd gnd OAI21X1
XFILL_6__2145_ gnd vdd FILL
XFILL_3__2436_ gnd vdd FILL
XFILL_3__2367_ gnd vdd FILL
XFILL_0__2658_ gnd vdd FILL
XFILL_6__2076_ gnd vdd FILL
XFILL_0__2589_ gnd vdd FILL
XFILL_1__3121_ gnd vdd FILL
XFILL_3__2298_ gnd vdd FILL
XFILL_7__1840_ gnd vdd FILL
XFILL_1__3052_ gnd vdd FILL
XFILL_1__2003_ gnd vdd FILL
XFILL_6__2978_ gnd vdd FILL
XFILL_7__1771_ gnd vdd FILL
XFILL_9__1707_ gnd vdd FILL
XFILL_6__1929_ gnd vdd FILL
XFILL_7__3510_ gnd vdd FILL
XFILL_4__1993_ gnd vdd FILL
XFILL_7__3441_ gnd vdd FILL
XFILL184650x15750 gnd vdd FILL
XFILL_1__2905_ gnd vdd FILL
XFILL_7__3372_ gnd vdd FILL
XFILL_4__2614_ gnd vdd FILL
XFILL_1__2836_ gnd vdd FILL
XFILL_7__2323_ gnd vdd FILL
XFILL_4__3594_ gnd vdd FILL
XFILL_7__2254_ gnd vdd FILL
XFILL_4__2545_ gnd vdd FILL
XFILL_4__2476_ gnd vdd FILL
XFILL_1__2767_ gnd vdd FILL
XFILL_7__2185_ gnd vdd FILL
XFILL_1__1718_ gnd vdd FILL
XFILL_1__2698_ gnd vdd FILL
XFILL_2__3230_ gnd vdd FILL
XFILL_2__3161_ gnd vdd FILL
XFILL_2__2112_ gnd vdd FILL
XFILL_4__3028_ gnd vdd FILL
XFILL_8__1880_ gnd vdd FILL
XFILL_2__3092_ gnd vdd FILL
XFILL_2__2043_ gnd vdd FILL
XFILL_8__3550_ gnd vdd FILL
XFILL_7__1969_ gnd vdd FILL
XFILL_8__3481_ gnd vdd FILL
XFILL_8__2501_ gnd vdd FILL
XFILL_5__2723_ gnd vdd FILL
XFILL_8__2432_ gnd vdd FILL
XFILL_2__2945_ gnd vdd FILL
XFILL_5__2654_ gnd vdd FILL
XFILL_2__2876_ gnd vdd FILL
XFILL_0__1960_ gnd vdd FILL
XFILL_8__2363_ gnd vdd FILL
XFILL_2__1827_ gnd vdd FILL
XFILL_0__1891_ gnd vdd FILL
XFILL_5__2585_ gnd vdd FILL
XFILL_8__2294_ gnd vdd FILL
XFILL_2__1758_ gnd vdd FILL
XFILL_0__3561_ gnd vdd FILL
XFILL_2__1689_ gnd vdd FILL
XFILL184350x4050 gnd vdd FILL
XFILL_5__3206_ gnd vdd FILL
XFILL_0__3492_ gnd vdd FILL
XFILL_2__3428_ gnd vdd FILL
XFILL_3__2221_ gnd vdd FILL
XFILL_0__2512_ gnd vdd FILL
XFILL_5__3137_ gnd vdd FILL
XFILL_0__2443_ gnd vdd FILL
XFILL_5__3068_ gnd vdd FILL
XFILL_3__2152_ gnd vdd FILL
XFILL_3__2083_ gnd vdd FILL
XFILL_6__2901_ gnd vdd FILL
XFILL_5__2019_ gnd vdd FILL
XFILL_0__2374_ gnd vdd FILL
X_1953_ _2950_/A _1984_/B _2735_/C _1954_/C vdd gnd OAI21X1
XFILL_6__2832_ gnd vdd FILL
XFILL_4_BUFX2_insert21 gnd vdd FILL
XFILL_4_BUFX2_insert10 gnd vdd FILL
X_1884_ _2430_/A _2430_/B _1884_/C _1903_/A vdd gnd OAI21X1
XFILL_4_BUFX2_insert43 gnd vdd FILL
XFILL_4_BUFX2_insert65 gnd vdd FILL
XFILL_6__2763_ gnd vdd FILL
XFILL_4_BUFX2_insert54 gnd vdd FILL
XFILL_3__2985_ gnd vdd FILL
XFILL_4_BUFX2_insert87 gnd vdd FILL
XFILL_6__1714_ gnd vdd FILL
XFILL_4_BUFX2_insert76 gnd vdd FILL
X_3554_ _3554_/A _3554_/B _3556_/A vdd gnd NOR2X1
XFILL_3__1936_ gnd vdd FILL
XFILL_6__2694_ gnd vdd FILL
X_3485_ _3485_/A _3544_/B _3544_/A _3544_/C vdd gnd OAI21X1
X_2505_ _2668_/B _2574_/B _2505_/C _2506_/C vdd gnd OAI21X1
XFILL_3__1867_ gnd vdd FILL
X_2436_ _2436_/A _2436_/B _2523_/A vdd gnd NOR2X1
XFILL_1__2621_ gnd vdd FILL
XFILL_3__1798_ gnd vdd FILL
XFILL_3__3537_ gnd vdd FILL
XFILL_4__2330_ gnd vdd FILL
X_2367_ _2872_/B _2367_/B _2429_/A vdd gnd NOR2X1
XFILL_3__3468_ gnd vdd FILL
XFILL_4__2261_ gnd vdd FILL
X_2298_ _2298_/A _3144_/C _2308_/B _2298_/D _2327_/B vdd gnd AOI22X1
XFILL_1__2552_ gnd vdd FILL
XFILL_3__2419_ gnd vdd FILL
XFILL_1__2483_ gnd vdd FILL
XFILL_6__3177_ gnd vdd FILL
XFILL_3__3399_ gnd vdd FILL
XFILL_6__2128_ gnd vdd FILL
XFILL_4__2192_ gnd vdd FILL
XFILL_6__2059_ gnd vdd FILL
XFILL_7__2941_ gnd vdd FILL
XFILL_1__3104_ gnd vdd FILL
XFILL_7__2872_ gnd vdd FILL
XFILL_1__3035_ gnd vdd FILL
XFILL_7__1823_ gnd vdd FILL
XFILL184650x27450 gnd vdd FILL
XFILL181650x35250 gnd vdd FILL
XFILL_7__1754_ gnd vdd FILL
XFILL_4__1976_ gnd vdd FILL
XFILL_7__3424_ gnd vdd FILL
XFILL_2__2730_ gnd vdd FILL
XFILL_5__2370_ gnd vdd FILL
XFILL_7__2306_ gnd vdd FILL
XFILL_2__2661_ gnd vdd FILL
XFILL_1__2819_ gnd vdd FILL
XFILL_4__2528_ gnd vdd FILL
XFILL_2__2592_ gnd vdd FILL
XFILL_7__2237_ gnd vdd FILL
XFILL_7__2168_ gnd vdd FILL
XFILL_4__2459_ gnd vdd FILL
XFILL_2__3213_ gnd vdd FILL
XFILL_8__2981_ gnd vdd FILL
XFILL_7__2099_ gnd vdd FILL
XFILL_8__1932_ gnd vdd FILL
XFILL_2__3144_ gnd vdd FILL
XFILL_2__3075_ gnd vdd FILL
XFILL_8__1863_ gnd vdd FILL
XFILL_2__2026_ gnd vdd FILL
XFILL_8__3602_ gnd vdd FILL
XFILL_0__2090_ gnd vdd FILL
XFILL_8__1794_ gnd vdd FILL
XFILL_8__3533_ gnd vdd FILL
XFILL_8__3464_ gnd vdd FILL
XFILL_3__2770_ gnd vdd FILL
XFILL_2__2928_ gnd vdd FILL
XFILL_8__3395_ gnd vdd FILL
XFILL_0__2992_ gnd vdd FILL
XFILL_8__2415_ gnd vdd FILL
XFILL_3__1721_ gnd vdd FILL
XFILL_5__2706_ gnd vdd FILL
X_3270_ _3270_/D vdd _3289_/R _3307_/CLK _3270_/Q vdd gnd DFFSR
XFILL_8__2346_ gnd vdd FILL
XFILL_5__2637_ gnd vdd FILL
XFILL_0__1943_ gnd vdd FILL
XFILL_2__2859_ gnd vdd FILL
XFILL_5__2568_ gnd vdd FILL
X_2221_ _2221_/A _3189_/A _2294_/A _2223_/C vdd gnd OAI21X1
XFILL_0__1874_ gnd vdd FILL
XFILL_6__3100_ gnd vdd FILL
XFILL_8__2277_ gnd vdd FILL
XFILL_6_CLKBUF1_insert29 gnd vdd FILL
X_2152_ _2242_/A _2242_/B _2153_/C vdd gnd NAND2X1
XFILL_5__2499_ gnd vdd FILL
XFILL_0__3544_ gnd vdd FILL
X_2083_ _2957_/B _2083_/Y vdd gnd INVX8
XFILL_6__3031_ gnd vdd FILL
XFILL183450x163950 gnd vdd FILL
XFILL_0__3475_ gnd vdd FILL
XFILL_3__2204_ gnd vdd FILL
XFILL_9__1972_ gnd vdd FILL
XFILL_3__3184_ gnd vdd FILL
XFILL_0__2426_ gnd vdd FILL
XFILL_3__2135_ gnd vdd FILL
XFILL_4_CLKBUF1_insert33 gnd vdd FILL
XFILL_0__2357_ gnd vdd FILL
XFILL_3__2066_ gnd vdd FILL
X_2985_ _2985_/A _2986_/B _3176_/B _2986_/C vdd gnd OAI21X1
XFILL_6__2815_ gnd vdd FILL
X_1936_ _1985_/A _3572_/Q _1936_/C _1937_/C vdd gnd AOI21X1
XFILL_0__2288_ gnd vdd FILL
X_1867_ _1867_/A _3285_/Q _1875_/A _1878_/B vdd gnd MUX2X1
XFILL_4__1830_ gnd vdd FILL
XFILL_6__2746_ gnd vdd FILL
X_1798_ _3063_/B _1806_/A vdd gnd INVX1
XFILL_4__3500_ gnd vdd FILL
X_3537_ _3560_/B _3558_/B _3537_/C _3538_/B vdd gnd AOI21X1
XFILL_3__2968_ gnd vdd FILL
XFILL_4__1761_ gnd vdd FILL
XFILL_6__2677_ gnd vdd FILL
XFILL_3__2899_ gnd vdd FILL
XFILL_3__1919_ gnd vdd FILL
XFILL_4__1692_ gnd vdd FILL
XFILL_1__1983_ gnd vdd FILL
XFILL_7__3140_ gnd vdd FILL
X_3468_ _3468_/A _3468_/B _3468_/S _3470_/B vdd gnd MUX2X1
XFILL_4__3431_ gnd vdd FILL
X_3399_ _3399_/A _3399_/B _3399_/C _3518_/A vdd gnd OAI21X1
X_2419_ _3308_/Q _2425_/B _2420_/C vdd gnd NAND2X1
XFILL_4__2313_ gnd vdd FILL
XFILL_7__3071_ gnd vdd FILL
XFILL_1__3584_ gnd vdd FILL
XFILL_1__2604_ gnd vdd FILL
XFILL_7__2022_ gnd vdd FILL
XFILL_1__2535_ gnd vdd FILL
XFILL_6__3229_ gnd vdd FILL
XFILL_0_BUFX2_insert41 gnd vdd FILL
XFILL_0_BUFX2_insert63 gnd vdd FILL
XFILL_0_BUFX2_insert74 gnd vdd FILL
XFILL_4__2244_ gnd vdd FILL
XFILL_0_BUFX2_insert52 gnd vdd FILL
XFILL_0_BUFX2_insert96 gnd vdd FILL
XFILL_0_BUFX2_insert85 gnd vdd FILL
XFILL_1__2466_ gnd vdd FILL
XFILL_4__2175_ gnd vdd FILL
XFILL184650x39150 gnd vdd FILL
XFILL_1__2397_ gnd vdd FILL
XFILL_7__2924_ gnd vdd FILL
XFILL_5__1870_ gnd vdd FILL
XFILL_7__2855_ gnd vdd FILL
XFILL_7__2786_ gnd vdd FILL
XFILL_1__3018_ gnd vdd FILL
XFILL_7__1806_ gnd vdd FILL
XFILL_7__1737_ gnd vdd FILL
XFILL_4__1959_ gnd vdd FILL
XFILL_5__3540_ gnd vdd FILL
XFILL_5__3471_ gnd vdd FILL
XFILL_7__3407_ gnd vdd FILL
XFILL_8__2200_ gnd vdd FILL
XFILL_5__2422_ gnd vdd FILL
XFILL_2__2713_ gnd vdd FILL
XFILL_8__3180_ gnd vdd FILL
XFILL_8__2131_ gnd vdd FILL
XFILL_2__2644_ gnd vdd FILL
XFILL_5__2353_ gnd vdd FILL
XFILL_8__2062_ gnd vdd FILL
XFILL_2__2575_ gnd vdd FILL
XFILL_5__2284_ gnd vdd FILL
XFILL_8__2964_ gnd vdd FILL
XFILL_2__3127_ gnd vdd FILL
XFILL_0__2211_ gnd vdd FILL
XFILL_8__1915_ gnd vdd FILL
XFILL_0__3191_ gnd vdd FILL
XFILL_8__2895_ gnd vdd FILL
XFILL_0__2142_ gnd vdd FILL
XFILL_2__3058_ gnd vdd FILL
XFILL_8__1846_ gnd vdd FILL
X_2770_ _3577_/Q _2770_/B _2770_/C _3363_/Q _2771_/B vdd gnd AOI22X1
XFILL_0__2073_ gnd vdd FILL
XFILL_8__1777_ gnd vdd FILL
X_1721_ _1739_/B _1793_/B _1783_/B vdd gnd NAND2X1
XFILL_2__2009_ gnd vdd FILL
XFILL_8__3516_ gnd vdd FILL
XFILL_5__1999_ gnd vdd FILL
XFILL_3__2822_ gnd vdd FILL
XFILL_6__3580_ gnd vdd FILL
XFILL_6__2600_ gnd vdd FILL
XFILL_6__2531_ gnd vdd FILL
XFILL_8__3447_ gnd vdd FILL
XFILL_6__2462_ gnd vdd FILL
XFILL_3__2753_ gnd vdd FILL
X_3322_ _3322_/D vdd _3347_/R _3573_/CLK _3322_/Q vdd gnd DFFSR
XFILL_8__3378_ gnd vdd FILL
XFILL_0__2975_ gnd vdd FILL
XFILL_3__1704_ gnd vdd FILL
XFILL_3__2684_ gnd vdd FILL
XFILL183750x167850 gnd vdd FILL
XFILL_0__1926_ gnd vdd FILL
XFILL_6__2393_ gnd vdd FILL
XFILL_8__2329_ gnd vdd FILL
X_3253_ _3253_/D vdd _3291_/R _3362_/CLK _3253_/Q vdd gnd DFFSR
XFILL_0__1857_ gnd vdd FILL
XFILL183450x175650 gnd vdd FILL
X_2204_ _3313_/Q _3311_/Q _3259_/Q _2205_/B vdd gnd MUX2X1
X_3184_ _3184_/A _3184_/B _3185_/C vdd gnd NOR2X1
X_2135_ _2135_/A _2135_/B _2319_/A _2285_/B vdd gnd NOR3X1
XFILL_6__3014_ gnd vdd FILL
XFILL_0__1788_ gnd vdd FILL
XFILL_0__3527_ gnd vdd FILL
XFILL_7_BUFX2_insert91 gnd vdd FILL
X_2066_ _2066_/A _2066_/B _2066_/C _2074_/A vdd gnd OAI21X1
XFILL_7_BUFX2_insert80 gnd vdd FILL
XFILL_1__2320_ gnd vdd FILL
XFILL_0__3458_ gnd vdd FILL
XFILL_1__2251_ gnd vdd FILL
XFILL_3__3167_ gnd vdd FILL
XFILL_0__2409_ gnd vdd FILL
XFILL_3__3098_ gnd vdd FILL
XFILL_0__3389_ gnd vdd FILL
XFILL_1__2182_ gnd vdd FILL
XFILL_3__2118_ gnd vdd FILL
XFILL_4__2931_ gnd vdd FILL
X_2968_ _2968_/A _2968_/B _2968_/C _2969_/C vdd gnd OAI21X1
XFILL_3__2049_ gnd vdd FILL
X_1919_ _3316_/Q _3029_/B _1920_/B vdd gnd NAND2X1
XFILL_7__2640_ gnd vdd FILL
XFILL_4__2862_ gnd vdd FILL
X_2899_ _2899_/A _2915_/A _2900_/B vdd gnd NAND2X1
XFILL_7__2571_ gnd vdd FILL
XFILL_9__3487_ gnd vdd FILL
XFILL_4__2793_ gnd vdd FILL
XFILL_6__2729_ gnd vdd FILL
XFILL_4__1813_ gnd vdd FILL
XFILL_4__1744_ gnd vdd FILL
XFILL_1__1966_ gnd vdd FILL
XFILL_4__3414_ gnd vdd FILL
XFILL_7__3123_ gnd vdd FILL
XFILL_1__1897_ gnd vdd FILL
XFILL_7__3054_ gnd vdd FILL
XFILL_2__2360_ gnd vdd FILL
XFILL_7__2005_ gnd vdd FILL
XFILL_1__3498_ gnd vdd FILL
XFILL_4__2227_ gnd vdd FILL
XFILL_1__2518_ gnd vdd FILL
XFILL_2__2291_ gnd vdd FILL
XFILL_1__2449_ gnd vdd FILL
XFILL_4__2158_ gnd vdd FILL
XFILL_5__2971_ gnd vdd FILL
XFILL_4__2089_ gnd vdd FILL
XFILL_7__2907_ gnd vdd FILL
XFILL_8__1700_ gnd vdd FILL
XFILL_8__2680_ gnd vdd FILL
XFILL_7__2838_ gnd vdd FILL
XFILL_5__1922_ gnd vdd FILL
XFILL_5__1853_ gnd vdd FILL
XFILL_7__2769_ gnd vdd FILL
XFILL_5__1784_ gnd vdd FILL
XFILL_5__3523_ gnd vdd FILL
XFILL_8__3232_ gnd vdd FILL
XFILL_5__3454_ gnd vdd FILL
XFILL_8__3163_ gnd vdd FILL
XFILL_0__2760_ gnd vdd FILL
XFILL_5__3385_ gnd vdd FILL
XFILL_8__2114_ gnd vdd FILL
XFILL_5__2405_ gnd vdd FILL
XFILL_0__1711_ gnd vdd FILL
XFILL_8__3094_ gnd vdd FILL
XFILL_5__2336_ gnd vdd FILL
XFILL_0__2691_ gnd vdd FILL
XFILL_2__2627_ gnd vdd FILL
XFILL_8__2045_ gnd vdd FILL
XFILL_2__2558_ gnd vdd FILL
XFILL_5__2267_ gnd vdd FILL
XFILL_2__2489_ gnd vdd FILL
XFILL_3__3021_ gnd vdd FILL
XFILL_0_BUFX2_insert0 gnd vdd FILL
XFILL_5__2198_ gnd vdd FILL
XFILL_8__2947_ gnd vdd FILL
XFILL_8__2878_ gnd vdd FILL
X_2822_ _3269_/Q _2960_/A vdd gnd INVX1
XFILL_6__1962_ gnd vdd FILL
XFILL_0__3174_ gnd vdd FILL
XFILL_8__1829_ gnd vdd FILL
XFILL_0__2125_ gnd vdd FILL
X_2753_ _2753_/A _2753_/B _2754_/B vdd gnd XOR2X1
XFILL_6__1893_ gnd vdd FILL
XFILL_0__2056_ gnd vdd FILL
X_1704_ _2675_/A _3295_/Q _1705_/C vdd gnd OR2X2
X_2684_ _3245_/Q _2685_/B _2686_/A vdd gnd NAND2X1
XFILL_3__2805_ gnd vdd FILL
XFILL_6__3563_ gnd vdd FILL
XFILL_6__3494_ gnd vdd FILL
XFILL_1__1820_ gnd vdd FILL
XFILL_3__2736_ gnd vdd FILL
XFILL_9__2223_ gnd vdd FILL
XFILL_6__2514_ gnd vdd FILL
X_3305_ _3305_/D _3313_/CLK _3305_/Q vdd gnd DFFPOSX1
XFILL_0__2958_ gnd vdd FILL
XFILL_1__1751_ gnd vdd FILL
XFILL_6__2445_ gnd vdd FILL
XFILL_6__2376_ gnd vdd FILL
XFILL_3__2667_ gnd vdd FILL
XFILL_0__1909_ gnd vdd FILL
XFILL_0__2889_ gnd vdd FILL
X_3236_ _3236_/D _3313_/R vdd _3363_/CLK _3236_/Q vdd gnd DFFSR
XFILL_3__2598_ gnd vdd FILL
XFILL_4__3130_ gnd vdd FILL
XFILL_1__3421_ gnd vdd FILL
X_3167_ _3167_/A _3167_/B _3172_/B _3168_/A vdd gnd NAND3X1
X_3098_ _3133_/A _3108_/B _3098_/C _3325_/D vdd gnd OAI21X1
X_2118_ _2305_/A _2894_/A _2191_/A vdd gnd NOR2X1
XFILL_4__3061_ gnd vdd FILL
XFILL_1__2303_ gnd vdd FILL
X_2049_ _3156_/C _3171_/A vdd gnd INVX1
XFILL_4__2012_ gnd vdd FILL
XFILL_3__3219_ gnd vdd FILL
XFILL_1__2234_ gnd vdd FILL
XFILL_1__2165_ gnd vdd FILL
XFILL_9__1869_ gnd vdd FILL
XFILL_4__2914_ gnd vdd FILL
XFILL_1__2096_ gnd vdd FILL
XFILL_3_BUFX2_insert4 gnd vdd FILL
XFILL_7__2623_ gnd vdd FILL
XFILL_4__2845_ gnd vdd FILL
XFILL_2__1860_ gnd vdd FILL
XFILL_7__2554_ gnd vdd FILL
XFILL_7__2485_ gnd vdd FILL
XFILL_4__2776_ gnd vdd FILL
XFILL_2__3530_ gnd vdd FILL
XFILL_1__2998_ gnd vdd FILL
XFILL_2__1791_ gnd vdd FILL
XFILL_4__1727_ gnd vdd FILL
XFILL_1__1949_ gnd vdd FILL
XFILL_2__3461_ gnd vdd FILL
XFILL_5__3170_ gnd vdd FILL
XFILL_7__3106_ gnd vdd FILL
XFILL_2__3392_ gnd vdd FILL
XFILL_2__2412_ gnd vdd FILL
XFILL_5__2121_ gnd vdd FILL
XFILL_7__3037_ gnd vdd FILL
XFILL_2__2343_ gnd vdd FILL
XFILL_5__2052_ gnd vdd FILL
XFILL_2__2274_ gnd vdd FILL
XFILL_8__2801_ gnd vdd FILL
XFILL_8__2732_ gnd vdd FILL
XFILL_5__2954_ gnd vdd FILL
XFILL_5__1905_ gnd vdd FILL
XFILL_8__2663_ gnd vdd FILL
XFILL_5__2885_ gnd vdd FILL
XFILL_8__2594_ gnd vdd FILL
XFILL_5__1836_ gnd vdd FILL
XFILL_5__1767_ gnd vdd FILL
XFILL_0__2812_ gnd vdd FILL
XFILL_5__3506_ gnd vdd FILL
XFILL_2__1989_ gnd vdd FILL
XFILL_8__3215_ gnd vdd FILL
XFILL_5__1698_ gnd vdd FILL
XFILL_1_BUFX2_insert18 gnd vdd FILL
XFILL_5__3437_ gnd vdd FILL
XFILL_6_BUFX2_insert8 gnd vdd FILL
XFILL_3__2521_ gnd vdd FILL
XFILL_6__2230_ gnd vdd FILL
XFILL_3__2452_ gnd vdd FILL
XFILL_8__3146_ gnd vdd FILL
XFILL_0__2743_ gnd vdd FILL
XFILL_6__2161_ gnd vdd FILL
XFILL_8__3077_ gnd vdd FILL
XFILL_5__3368_ gnd vdd FILL
X_3021_ _3197_/C DI[7] _3022_/C vdd gnd NAND2X1
XFILL_0__2674_ gnd vdd FILL
XFILL_8__2028_ gnd vdd FILL
XFILL_3__2383_ gnd vdd FILL
XFILL_5__2319_ gnd vdd FILL
XFILL_6__2092_ gnd vdd FILL
XFILL_9__2841_ gnd vdd FILL
XFILL_3__3004_ gnd vdd FILL
XFILL_6__2994_ gnd vdd FILL
XFILL_0__3226_ gnd vdd FILL
X_2805_ _2933_/B _2899_/A _2851_/A vdd gnd NOR2X1
XFILL_6__1945_ gnd vdd FILL
XFILL_0__3157_ gnd vdd FILL
XFILL183150x7950 gnd vdd FILL
XFILL_0__2108_ gnd vdd FILL
XFILL_6__1876_ gnd vdd FILL
XFILL_0__3088_ gnd vdd FILL
X_2736_ _3574_/Q _2770_/B _3177_/B _2737_/C vdd gnd AOI21X1
XFILL_1__2921_ gnd vdd FILL
XFILL_0__2039_ gnd vdd FILL
XFILL_4__2630_ gnd vdd FILL
X_2667_ _2675_/A _2673_/B _2668_/D vdd gnd NAND2X1
XFILL_6__3546_ gnd vdd FILL
XFILL_1__2852_ gnd vdd FILL
XFILL_7__2270_ gnd vdd FILL
XFILL_1__1803_ gnd vdd FILL
XFILL_4__2561_ gnd vdd FILL
X_2598_ _2598_/A _2598_/B _2993_/B _2599_/B vdd gnd OAI21X1
XFILL_6__3477_ gnd vdd FILL
XFILL_1__2783_ gnd vdd FILL
XFILL_4__2492_ gnd vdd FILL
XFILL_3__2719_ gnd vdd FILL
XFILL_6__2428_ gnd vdd FILL
XFILL_1__1734_ gnd vdd FILL
XFILL_6__2359_ gnd vdd FILL
X_3219_ _3219_/A _3228_/B _3219_/C _3357_/D vdd gnd OAI21X1
XFILL_1__3404_ gnd vdd FILL
XFILL_4__3113_ gnd vdd FILL
XFILL_4__3044_ gnd vdd FILL
XFILL_1__2217_ gnd vdd FILL
XFILL_7__1985_ gnd vdd FILL
XFILL_1__3197_ gnd vdd FILL
XBUFX2_insert21 _2580_/Y _3282_/R vdd gnd BUFX2
XBUFX2_insert10 RDY _3566_/A vdd gnd BUFX2
XFILL_1__2148_ gnd vdd FILL
XFILL_1__2079_ gnd vdd FILL
XFILL_2__2961_ gnd vdd FILL
XBUFX2_insert43 _1734_/Y _2299_/A vdd gnd BUFX2
XBUFX2_insert65 _3198_/Y _3228_/B vdd gnd BUFX2
XBUFX2_insert54 _1733_/Y _2432_/A vdd gnd BUFX2
XBUFX2_insert87 _1729_/Y _2276_/A vdd gnd BUFX2
XFILL_7__3586_ gnd vdd FILL
XFILL_2__1912_ gnd vdd FILL
XFILL_7__2606_ gnd vdd FILL
XFILL_5__2670_ gnd vdd FILL
XBUFX2_insert76 _1694_/Y _2768_/A vdd gnd BUFX2
XFILL_4__2828_ gnd vdd FILL
XFILL_2__2892_ gnd vdd FILL
XFILL_7__2537_ gnd vdd FILL
XFILL_2__1843_ gnd vdd FILL
XFILL_4__2759_ gnd vdd FILL
XFILL_8_BUFX2_insert24 gnd vdd FILL
XFILL_7__2468_ gnd vdd FILL
XFILL_2__1774_ gnd vdd FILL
XFILL_8_BUFX2_insert13 gnd vdd FILL
XFILL_8_BUFX2_insert57 gnd vdd FILL
XFILL_2__3513_ gnd vdd FILL
XFILL_8__3000_ gnd vdd FILL
XFILL_7__2399_ gnd vdd FILL
XFILL_8_BUFX2_insert46 gnd vdd FILL
XFILL_5__3222_ gnd vdd FILL
XFILL_2__3444_ gnd vdd FILL
XFILL_8_BUFX2_insert79 gnd vdd FILL
XFILL_8_BUFX2_insert68 gnd vdd FILL
XFILL_5__3153_ gnd vdd FILL
XFILL_5__2104_ gnd vdd FILL
XFILL_2__3375_ gnd vdd FILL
XFILL_5__3084_ gnd vdd FILL
XFILL_5__2035_ gnd vdd FILL
XFILL_2__2326_ gnd vdd FILL
XFILL_0__2390_ gnd vdd FILL
XFILL_2__2257_ gnd vdd FILL
XFILL_2__2188_ gnd vdd FILL
XFILL_0__3011_ gnd vdd FILL
XFILL_8__2715_ gnd vdd FILL
X_3570_ _3570_/D vdd _3578_/R _3573_/CLK _3570_/Q vdd gnd DFFSR
XFILL_6__1730_ gnd vdd FILL
XFILL_3__1952_ gnd vdd FILL
XFILL_5__2937_ gnd vdd FILL
XFILL_8__2646_ gnd vdd FILL
XFILL_5__2868_ gnd vdd FILL
X_2521_ _3030_/C _2570_/B _2521_/C _2522_/C vdd gnd OAI21X1
XFILL_6__3400_ gnd vdd FILL
XFILL_8__2577_ gnd vdd FILL
XFILL_5__1819_ gnd vdd FILL
XFILL_3__1883_ gnd vdd FILL
XFILL_5__2799_ gnd vdd FILL
X_2452_ _2519_/C _2455_/B vdd gnd INVX1
XFILL_3__3553_ gnd vdd FILL
X_2383_ _3313_/Q _2425_/B _2384_/C vdd gnd NAND2X1
XFILL_3__2504_ gnd vdd FILL
XFILL_3__3484_ gnd vdd FILL
XFILL_8__3129_ gnd vdd FILL
XFILL_6__2213_ gnd vdd FILL
XFILL_0__2726_ gnd vdd FILL
XFILL_6__3193_ gnd vdd FILL
X_3004_ _3312_/Q _3005_/A _3005_/C vdd gnd NAND2X1
XFILL_6__2144_ gnd vdd FILL
XFILL_3__2435_ gnd vdd FILL
XFILL_3__2366_ gnd vdd FILL
XFILL_0__2657_ gnd vdd FILL
XFILL_6__2075_ gnd vdd FILL
XFILL_0__2588_ gnd vdd FILL
XFILL_1__3120_ gnd vdd FILL
XFILL_3__2297_ gnd vdd FILL
XFILL_1__3051_ gnd vdd FILL
XFILL_1__2002_ gnd vdd FILL
XFILL_0__3209_ gnd vdd FILL
XFILL_6__2977_ gnd vdd FILL
XFILL_7__1770_ gnd vdd FILL
XFILL_6__1928_ gnd vdd FILL
XFILL_4__1992_ gnd vdd FILL
XFILL_6__1859_ gnd vdd FILL
XFILL_7__3440_ gnd vdd FILL
X_2719_ _3249_/Q _2725_/D _2725_/C _2720_/B vdd gnd NAND3X1
XFILL_1__2904_ gnd vdd FILL
XFILL_7__3371_ gnd vdd FILL
XFILL_4__3593_ gnd vdd FILL
XFILL_4__2613_ gnd vdd FILL
XFILL_1__2835_ gnd vdd FILL
XFILL_6__3529_ gnd vdd FILL
XFILL_7__2322_ gnd vdd FILL
XFILL_4__2544_ gnd vdd FILL
XFILL_7__2253_ gnd vdd FILL
XFILL_1__2766_ gnd vdd FILL
XFILL_4__2475_ gnd vdd FILL
XFILL_7__2184_ gnd vdd FILL
XFILL_1__1717_ gnd vdd FILL
XFILL_1__2697_ gnd vdd FILL
XFILL_2__3160_ gnd vdd FILL
XFILL_2__2111_ gnd vdd FILL
XFILL_2__3091_ gnd vdd FILL
XFILL_4__3027_ gnd vdd FILL
XFILL_2__2042_ gnd vdd FILL
XFILL_7__1968_ gnd vdd FILL
XFILL_8__3480_ gnd vdd FILL
XFILL_8__2500_ gnd vdd FILL
XFILL_7__1899_ gnd vdd FILL
XFILL_5__2722_ gnd vdd FILL
XFILL_8__2431_ gnd vdd FILL
XFILL_2__2944_ gnd vdd FILL
XFILL_5__2653_ gnd vdd FILL
XFILL_8__2362_ gnd vdd FILL
XFILL_2__2875_ gnd vdd FILL
XFILL_5__2584_ gnd vdd FILL
XFILL_0__1890_ gnd vdd FILL
XFILL_8__2293_ gnd vdd FILL
XFILL_2__1826_ gnd vdd FILL
XFILL_0__3560_ gnd vdd FILL
XFILL_2__1757_ gnd vdd FILL
XFILL_5__3205_ gnd vdd FILL
XFILL_0__2511_ gnd vdd FILL
XFILL_2__1688_ gnd vdd FILL
XFILL_0__3491_ gnd vdd FILL
XFILL_2__3427_ gnd vdd FILL
XFILL_3__2220_ gnd vdd FILL
XFILL_5__3136_ gnd vdd FILL
XFILL_3__2151_ gnd vdd FILL
XFILL_0__2442_ gnd vdd FILL
XFILL_2__2309_ gnd vdd FILL
XFILL_5__3067_ gnd vdd FILL
XFILL_0__2373_ gnd vdd FILL
XFILL_6__2900_ gnd vdd FILL
XFILL_5__2018_ gnd vdd FILL
XFILL_3__2082_ gnd vdd FILL
X_1952_ _3360_/Q _2691_/A _2735_/C vdd gnd NAND2X1
XFILL_6__2831_ gnd vdd FILL
XFILL_4_BUFX2_insert22 gnd vdd FILL
X_1883_ _1883_/A _1884_/C vdd gnd INVX1
XFILL_4_BUFX2_insert11 gnd vdd FILL
XFILL_4_BUFX2_insert66 gnd vdd FILL
XFILL_4_BUFX2_insert44 gnd vdd FILL
XFILL_4_BUFX2_insert55 gnd vdd FILL
XFILL_6__2762_ gnd vdd FILL
XFILL_3__2984_ gnd vdd FILL
XFILL_4_BUFX2_insert88 gnd vdd FILL
XFILL_6__1713_ gnd vdd FILL
XFILL_4_BUFX2_insert77 gnd vdd FILL
X_3553_ _3574_/Q _3553_/B _3556_/C vdd gnd NAND2X1
XFILL_3__1935_ gnd vdd FILL
XFILL_6__2693_ gnd vdd FILL
XFILL_8__2629_ gnd vdd FILL
X_3484_ _3514_/B _3484_/B _3484_/C _3544_/B vdd gnd AOI21X1
X_2504_ _3576_/Q _2508_/B _2504_/C _2505_/C vdd gnd AOI21X1
XFILL_3__1866_ gnd vdd FILL
X_2435_ _2435_/A _2435_/B _2436_/B vdd gnd OR2X2
XFILL_1__2620_ gnd vdd FILL
XFILL_3__1797_ gnd vdd FILL
XFILL_3__3536_ gnd vdd FILL
X_2366_ _2407_/A _2426_/B vdd gnd INVX2
XFILL_3__3467_ gnd vdd FILL
XFILL_4__2260_ gnd vdd FILL
X_2297_ _2297_/A _2297_/B _2308_/B vdd gnd NOR2X1
XFILL_1__2551_ gnd vdd FILL
XFILL_3__2418_ gnd vdd FILL
XFILL_1__2482_ gnd vdd FILL
XFILL_0__2709_ gnd vdd FILL
XFILL_6__3176_ gnd vdd FILL
XFILL_3__3398_ gnd vdd FILL
XFILL_4__2191_ gnd vdd FILL
XFILL_6__2127_ gnd vdd FILL
XFILL_7__2940_ gnd vdd FILL
XFILL_3__2349_ gnd vdd FILL
XFILL_6__2058_ gnd vdd FILL
XFILL_1__3103_ gnd vdd FILL
XFILL_7__2871_ gnd vdd FILL
XFILL_1__3034_ gnd vdd FILL
XFILL_9__2738_ gnd vdd FILL
XFILL_7__1822_ gnd vdd FILL
XFILL_7__1753_ gnd vdd FILL
XFILL_4__1975_ gnd vdd FILL
XFILL_7__3423_ gnd vdd FILL
XFILL_2__2660_ gnd vdd FILL
XFILL_7__2305_ gnd vdd FILL
XFILL_1__2818_ gnd vdd FILL
XFILL_4__2527_ gnd vdd FILL
XFILL_2__2591_ gnd vdd FILL
XFILL_7__2236_ gnd vdd FILL
XFILL_1__2749_ gnd vdd FILL
XFILL_7__2167_ gnd vdd FILL
XFILL_4__2458_ gnd vdd FILL
XFILL_4__2389_ gnd vdd FILL
XFILL_2__3212_ gnd vdd FILL
XFILL_7__2098_ gnd vdd FILL
XFILL_8__2980_ gnd vdd FILL
XFILL_2__3143_ gnd vdd FILL
XFILL_8__1931_ gnd vdd FILL
XFILL_8__1862_ gnd vdd FILL
XFILL_2__3074_ gnd vdd FILL
XFILL_2__2025_ gnd vdd FILL
XFILL_8__3601_ gnd vdd FILL
XFILL_8__3532_ gnd vdd FILL
XFILL_8__1793_ gnd vdd FILL
XFILL_8__3463_ gnd vdd FILL
XFILL_5__2705_ gnd vdd FILL
XFILL_2__2927_ gnd vdd FILL
XFILL_8__3394_ gnd vdd FILL
XFILL_0__2991_ gnd vdd FILL
XFILL_8__2414_ gnd vdd FILL
XFILL_3__1720_ gnd vdd FILL
XFILL_0__1942_ gnd vdd FILL
XFILL_8__2345_ gnd vdd FILL
XFILL_5__2636_ gnd vdd FILL
XFILL_2__2858_ gnd vdd FILL
X_2220_ _2278_/A _2367_/B _2220_/C _2345_/B vdd gnd OAI21X1
XFILL_5__2567_ gnd vdd FILL
XFILL_0__1873_ gnd vdd FILL
XFILL_2__2789_ gnd vdd FILL
XFILL_8__2276_ gnd vdd FILL
XFILL_2__1809_ gnd vdd FILL
X_2151_ _2958_/A _2781_/B _2242_/B vdd gnd NOR2X1
XFILL_5__2498_ gnd vdd FILL
XFILL_0__3543_ gnd vdd FILL
X_2082_ _2298_/A _3157_/C _2305_/B _2298_/D _2339_/B vdd gnd AOI22X1
XFILL_6__3030_ gnd vdd FILL
XFILL_0__3474_ gnd vdd FILL
XFILL_3__2203_ gnd vdd FILL
XFILL_5__3119_ gnd vdd FILL
XFILL_0__2425_ gnd vdd FILL
XFILL_3__3183_ gnd vdd FILL
XFILL_3__2134_ gnd vdd FILL
XFILL_4_CLKBUF1_insert34 gnd vdd FILL
XFILL_3__2065_ gnd vdd FILL
XFILL_0__2356_ gnd vdd FILL
X_2984_ _3056_/A _3148_/B _2984_/C _2986_/A vdd gnd OAI21X1
XFILL_0__2287_ gnd vdd FILL
X_1935_ _2985_/A _1984_/B _2715_/C _1936_/C vdd gnd OAI21X1
XFILL_6__2814_ gnd vdd FILL
X_1866_ _1874_/B _1873_/B _1873_/A _1867_/A vdd gnd NAND3X1
XFILL_6__2745_ gnd vdd FILL
X_1797_ _3166_/C _3152_/C _3063_/B vdd gnd NAND2X1
X_3536_ _3536_/A _3536_/B _3560_/B vdd gnd NAND2X1
XFILL_4__1760_ gnd vdd FILL
XFILL_3__2967_ gnd vdd FILL
XFILL_1__1982_ gnd vdd FILL
XFILL_6__2676_ gnd vdd FILL
XFILL_3__1918_ gnd vdd FILL
XFILL_3__2898_ gnd vdd FILL
XFILL_4__1691_ gnd vdd FILL
XFILL_4__3430_ gnd vdd FILL
X_3467_ _3521_/A _3467_/B _3543_/C vdd gnd NOR2X1
XFILL_3__1849_ gnd vdd FILL
X_3398_ _3404_/B _3398_/B _3459_/A _3399_/A vdd gnd OAI21X1
X_2418_ _2872_/B _3077_/C _3253_/Q _2422_/A vdd gnd OAI21X1
XFILL_3__3519_ gnd vdd FILL
XFILL_4__2312_ gnd vdd FILL
XFILL_7__3070_ gnd vdd FILL
X_2349_ _2349_/A _2349_/B _2350_/B vdd gnd NOR2X1
XFILL_1__3583_ gnd vdd FILL
XFILL_1__2603_ gnd vdd FILL
XFILL_0_BUFX2_insert20 gnd vdd FILL
XFILL_7__2021_ gnd vdd FILL
XFILL_0_BUFX2_insert42 gnd vdd FILL
XFILL_1__2534_ gnd vdd FILL
XFILL_6__3228_ gnd vdd FILL
XFILL_0_BUFX2_insert64 gnd vdd FILL
XFILL_4__2243_ gnd vdd FILL
XFILL_0_BUFX2_insert75 gnd vdd FILL
XFILL_0_BUFX2_insert53 gnd vdd FILL
XFILL_6__3159_ gnd vdd FILL
XFILL_0_BUFX2_insert97 gnd vdd FILL
XFILL_4__2174_ gnd vdd FILL
XFILL_1__2465_ gnd vdd FILL
XFILL_0_BUFX2_insert86 gnd vdd FILL
XFILL_1__2396_ gnd vdd FILL
XFILL_7__2923_ gnd vdd FILL
XFILL_7__2854_ gnd vdd FILL
XFILL_1__3017_ gnd vdd FILL
XFILL_7__1805_ gnd vdd FILL
XFILL_7__2785_ gnd vdd FILL
XFILL_7__1736_ gnd vdd FILL
XFILL_4__1958_ gnd vdd FILL
XFILL_5__3470_ gnd vdd FILL
XFILL_7__3406_ gnd vdd FILL
XFILL_4__1889_ gnd vdd FILL
XFILL_5__2421_ gnd vdd FILL
XFILL_2__2712_ gnd vdd FILL
XFILL_8__2130_ gnd vdd FILL
XFILL_2__2643_ gnd vdd FILL
XFILL_4__3559_ gnd vdd FILL
XFILL_5__2352_ gnd vdd FILL
XFILL_8__2061_ gnd vdd FILL
XFILL_2__2574_ gnd vdd FILL
XFILL_5__2283_ gnd vdd FILL
XFILL_7__2219_ gnd vdd FILL
XFILL181350x117150 gnd vdd FILL
XFILL181650x109350 gnd vdd FILL
XFILL_7__3199_ gnd vdd FILL
XFILL_8__2963_ gnd vdd FILL
XFILL_2__3126_ gnd vdd FILL
XFILL_0__2210_ gnd vdd FILL
XFILL_8__1914_ gnd vdd FILL
XFILL_0__3190_ gnd vdd FILL
XFILL_8__2894_ gnd vdd FILL
XFILL_0__2141_ gnd vdd FILL
XFILL_2__3057_ gnd vdd FILL
XFILL_8__1845_ gnd vdd FILL
XFILL_0__2072_ gnd vdd FILL
X_1720_ _3235_/Q _1739_/B vdd gnd INVX1
XFILL_8__1776_ gnd vdd FILL
XFILL_2__2008_ gnd vdd FILL
XFILL_8__3515_ gnd vdd FILL
XFILL_5__1998_ gnd vdd FILL
XFILL_3__2821_ gnd vdd FILL
XFILL_8__3446_ gnd vdd FILL
XFILL_6__2530_ gnd vdd FILL
X_3321_ _3321_/D vdd _3346_/R _3346_/CLK _3321_/Q vdd gnd DFFSR
XFILL_6__2461_ gnd vdd FILL
XFILL_3__2752_ gnd vdd FILL
XFILL_8__3377_ gnd vdd FILL
XFILL_0__2974_ gnd vdd FILL
XFILL_3__1703_ gnd vdd FILL
XFILL_3__2683_ gnd vdd FILL
XFILL_5__2619_ gnd vdd FILL
XFILL_8__2328_ gnd vdd FILL
XFILL_5__3599_ gnd vdd FILL
XFILL_6__2392_ gnd vdd FILL
XFILL_0__1925_ gnd vdd FILL
X_3252_ _3252_/D vdd _3291_/R _3355_/CLK _3252_/Q vdd gnd DFFSR
XFILL_8__2259_ gnd vdd FILL
X_2203_ _2203_/A _2203_/B _3258_/Q _2205_/C vdd gnd OAI21X1
XFILL_0__1856_ gnd vdd FILL
X_3183_ _3237_/Q _3183_/B _3183_/C _3184_/A vdd gnd OAI21X1
X_2134_ _2700_/B _2134_/B _3022_/A _2717_/B _2135_/B vdd gnd OAI22X1
XFILL_6__3013_ gnd vdd FILL
XFILL_0__1787_ gnd vdd FILL
XFILL_0__3526_ gnd vdd FILL
XFILL_7_BUFX2_insert92 gnd vdd FILL
X_2065_ _2786_/A _2275_/B _2279_/A _2066_/C vdd gnd NAND3X1
XFILL_7_BUFX2_insert81 gnd vdd FILL
XFILL_7_BUFX2_insert70 gnd vdd FILL
XFILL_1__2250_ gnd vdd FILL
XFILL_0__3457_ gnd vdd FILL
XFILL_3__3166_ gnd vdd FILL
XFILL_0__3388_ gnd vdd FILL
XFILL_1__2181_ gnd vdd FILL
XFILL_0__2408_ gnd vdd FILL
XFILL_3__3097_ gnd vdd FILL
XFILL_3__2117_ gnd vdd FILL
XFILL_0__2339_ gnd vdd FILL
XFILL_4__2930_ gnd vdd FILL
X_2967_ _3260_/Q _3576_/Q _2968_/B vdd gnd NAND2X1
XFILL_3__2048_ gnd vdd FILL
X_1918_ _3332_/Q _3110_/A _3127_/B _3341_/Q _1920_/C vdd gnd AOI22X1
X_2898_ _2898_/A _2898_/B _2898_/C _3284_/D vdd gnd OAI21X1
XFILL_4__2861_ gnd vdd FILL
X_1849_ _3166_/C _3165_/A _3189_/B vdd gnd NOR2X1
XFILL_7__2570_ gnd vdd FILL
XFILL_4__2792_ gnd vdd FILL
XFILL_4__1812_ gnd vdd FILL
XFILL_6__2728_ gnd vdd FILL
XFILL_4__1743_ gnd vdd FILL
XFILL_1__1965_ gnd vdd FILL
X_3519_ _3519_/A _3519_/B _3520_/C _3523_/B vdd gnd OAI21X1
XFILL_6__2659_ gnd vdd FILL
XFILL_4__3413_ gnd vdd FILL
XFILL_1__1896_ gnd vdd FILL
XFILL_7__3122_ gnd vdd FILL
XFILL_7__3053_ gnd vdd FILL
XFILL_7__2004_ gnd vdd FILL
XFILL_1__3566_ gnd vdd FILL
XFILL_1__3497_ gnd vdd FILL
XFILL_4__2226_ gnd vdd FILL
XFILL_2__2290_ gnd vdd FILL
XFILL_1__2517_ gnd vdd FILL
XFILL_1__2448_ gnd vdd FILL
XFILL_4__2157_ gnd vdd FILL
XFILL_7__2906_ gnd vdd FILL
XFILL_5__2970_ gnd vdd FILL
XFILL_4__2088_ gnd vdd FILL
XFILL_1__2379_ gnd vdd FILL
XFILL_5__1921_ gnd vdd FILL
XFILL_7__2837_ gnd vdd FILL
XFILL_5__1852_ gnd vdd FILL
XFILL_7__2768_ gnd vdd FILL
XFILL_7__1719_ gnd vdd FILL
XFILL_5__1783_ gnd vdd FILL
XFILL_5__3522_ gnd vdd FILL
XFILL_7__2699_ gnd vdd FILL
XFILL_8__3231_ gnd vdd FILL
XFILL_5__3453_ gnd vdd FILL
XFILL_8__3162_ gnd vdd FILL
XFILL_5__3384_ gnd vdd FILL
XFILL_5__2404_ gnd vdd FILL
XFILL_8__2113_ gnd vdd FILL
XFILL_0__1710_ gnd vdd FILL
XFILL_0__2690_ gnd vdd FILL
XFILL_8__3093_ gnd vdd FILL
XFILL_5__2335_ gnd vdd FILL
XFILL_2__2626_ gnd vdd FILL
XFILL_8__2044_ gnd vdd FILL
XFILL_2__2557_ gnd vdd FILL
XFILL_5__2266_ gnd vdd FILL
XFILL_2__2488_ gnd vdd FILL
XFILL_5__2197_ gnd vdd FILL
XFILL_3__3020_ gnd vdd FILL
XFILL_0_BUFX2_insert1 gnd vdd FILL
XFILL_8__2946_ gnd vdd FILL
XFILL_2__3109_ gnd vdd FILL
X_2821_ _2821_/A _2926_/B _2821_/C _3268_/D vdd gnd OAI21X1
XFILL_8__2877_ gnd vdd FILL
XFILL_6__1961_ gnd vdd FILL
XFILL_0__3173_ gnd vdd FILL
XFILL_0__2124_ gnd vdd FILL
XFILL_6__1892_ gnd vdd FILL
X_2752_ _2752_/A _2775_/C _2753_/A vdd gnd NAND2X1
XFILL_8__1828_ gnd vdd FILL
X_1703_ _2950_/A _3294_/D vdd gnd INVX1
XFILL_0__2055_ gnd vdd FILL
XFILL_6__3562_ gnd vdd FILL
XFILL_8__1759_ gnd vdd FILL
X_2683_ _2697_/B _2751_/B _2708_/A _2706_/B vdd gnd OAI21X1
XFILL_3__2804_ gnd vdd FILL
XFILL_6__2513_ gnd vdd FILL
XFILL_6__3493_ gnd vdd FILL
XFILL_8__3429_ gnd vdd FILL
XFILL_3__2735_ gnd vdd FILL
X_3304_ _3304_/D _3346_/CLK _3304_/Q vdd gnd DFFPOSX1
XFILL_0__2957_ gnd vdd FILL
XFILL_1__1750_ gnd vdd FILL
XFILL_6__2444_ gnd vdd FILL
XFILL184650x160050 gnd vdd FILL
XFILL_6__2375_ gnd vdd FILL
X_3235_ _3235_/D vdd _3363_/R _3363_/CLK _3235_/Q vdd gnd DFFSR
XFILL_3__2666_ gnd vdd FILL
XFILL_0__1908_ gnd vdd FILL
XFILL_0__2888_ gnd vdd FILL
XFILL_3__2597_ gnd vdd FILL
XFILL_1__3420_ gnd vdd FILL
XFILL_0__1839_ gnd vdd FILL
X_3166_ _3166_/A _3166_/B _3166_/C _3166_/D _3172_/B vdd gnd AOI22X1
X_3097_ _3115_/A _3107_/B _3325_/Q _3098_/C vdd gnd OAI21X1
X_2117_ _2890_/A _2864_/A _2288_/C vdd gnd NOR2X1
XFILL_4__3060_ gnd vdd FILL
XFILL_0__3509_ gnd vdd FILL
XFILL_1__2302_ gnd vdd FILL
X_2048_ _2379_/A _2048_/B _3156_/C vdd gnd NAND2X1
XFILL_4__2011_ gnd vdd FILL
XFILL_3__3218_ gnd vdd FILL
XFILL_1__2233_ gnd vdd FILL
XFILL_3__3149_ gnd vdd FILL
XFILL_1__2164_ gnd vdd FILL
XFILL_1__2095_ gnd vdd FILL
XFILL_4__2913_ gnd vdd FILL
XFILL_3_BUFX2_insert5 gnd vdd FILL
XFILL_7__2622_ gnd vdd FILL
XFILL_4__2844_ gnd vdd FILL
XFILL_7__2553_ gnd vdd FILL
XFILL_3_BUFX2_insert90 gnd vdd FILL
XFILL_7__2484_ gnd vdd FILL
XFILL_4__2775_ gnd vdd FILL
XFILL_2__1790_ gnd vdd FILL
XFILL_1__2997_ gnd vdd FILL
XFILL_4__1726_ gnd vdd FILL
XFILL_1__1948_ gnd vdd FILL
XFILL_1__1879_ gnd vdd FILL
XFILL_7__3105_ gnd vdd FILL
XFILL_2__3460_ gnd vdd FILL
XFILL_2__3391_ gnd vdd FILL
XFILL_5__2120_ gnd vdd FILL
XFILL_2__2411_ gnd vdd FILL
XFILL_1__3549_ gnd vdd FILL
XFILL_7__3036_ gnd vdd FILL
XFILL_2__2342_ gnd vdd FILL
XFILL_5__2051_ gnd vdd FILL
XFILL_2__2273_ gnd vdd FILL
XFILL_8__2800_ gnd vdd FILL
XFILL_4__2209_ gnd vdd FILL
XFILL_4__3189_ gnd vdd FILL
XFILL_8__2731_ gnd vdd FILL
XFILL_5__2953_ gnd vdd FILL
XFILL_8__2662_ gnd vdd FILL
XFILL_5__2884_ gnd vdd FILL
XFILL_5__1904_ gnd vdd FILL
XFILL_8__2593_ gnd vdd FILL
XFILL_5__1835_ gnd vdd FILL
XFILL_5__1766_ gnd vdd FILL
XFILL_0__2811_ gnd vdd FILL
XFILL_5__3505_ gnd vdd FILL
XFILL_5__1697_ gnd vdd FILL
XFILL_2__1988_ gnd vdd FILL
XFILL_8__3214_ gnd vdd FILL
XFILL_5__3436_ gnd vdd FILL
XFILL183150x109350 gnd vdd FILL
XFILL_3__2520_ gnd vdd FILL
XFILL_1_BUFX2_insert19 gnd vdd FILL
XFILL_3__2451_ gnd vdd FILL
XFILL_6_BUFX2_insert9 gnd vdd FILL
XFILL_8__3145_ gnd vdd FILL
XFILL_0__2742_ gnd vdd FILL
XFILL_6__2160_ gnd vdd FILL
XFILL_8__3076_ gnd vdd FILL
XFILL_5__3367_ gnd vdd FILL
XFILL_3__2382_ gnd vdd FILL
X_3020_ _3314_/Q _3022_/B vdd gnd INVX1
XFILL_2__2609_ gnd vdd FILL
XFILL_0__2673_ gnd vdd FILL
XFILL_8__2027_ gnd vdd FILL
XFILL_5__2318_ gnd vdd FILL
XFILL_2__3589_ gnd vdd FILL
XFILL_6__2091_ gnd vdd FILL
XFILL_5__2249_ gnd vdd FILL
XFILL_3__3003_ gnd vdd FILL
XFILL_8__2929_ gnd vdd FILL
XFILL_6__2993_ gnd vdd FILL
XFILL_9__1722_ gnd vdd FILL
XFILL_0__3225_ gnd vdd FILL
X_2804_ _2906_/A _3006_/B _3264_/Q _2807_/C vdd gnd OAI21X1
XFILL_0__3156_ gnd vdd FILL
XFILL_6__1944_ gnd vdd FILL
XFILL_0__2107_ gnd vdd FILL
XFILL_6__1875_ gnd vdd FILL
XFILL_0__3087_ gnd vdd FILL
X_2735_ _2744_/B _2746_/B _2735_/C _2738_/B vdd gnd OAI21X1
XFILL_1__2920_ gnd vdd FILL
XFILL_0__2038_ gnd vdd FILL
X_2666_ _2674_/A _2674_/C _2673_/B vdd gnd NAND2X1
XFILL_6__3545_ gnd vdd FILL
XFILL_1__2851_ gnd vdd FILL
XFILL_6__3476_ gnd vdd FILL
XFILL_4__2560_ gnd vdd FILL
XFILL_1__1802_ gnd vdd FILL
X_2597_ _2612_/B _2702_/B _2598_/A vdd gnd NOR2X1
XFILL_6__2427_ gnd vdd FILL
XFILL_4__2491_ gnd vdd FILL
XFILL_3__2718_ gnd vdd FILL
XFILL_1__2782_ gnd vdd FILL
XFILL_1__1733_ gnd vdd FILL
XFILL_3__2649_ gnd vdd FILL
XFILL_6__2358_ gnd vdd FILL
X_3218_ _3594_/A _3228_/B _3219_/C vdd gnd NAND2X1
XFILL_1__3403_ gnd vdd FILL
X_3149_ _3166_/C _3165_/A _3149_/C _3150_/A vdd gnd OAI21X1
XFILL_6__2289_ gnd vdd FILL
XFILL_4__3112_ gnd vdd FILL
XFILL_4__3043_ gnd vdd FILL
XFILL_1__2216_ gnd vdd FILL
XFILL_7__1984_ gnd vdd FILL
XFILL_1__3196_ gnd vdd FILL
XFILL_1__2147_ gnd vdd FILL
XBUFX2_insert22 _2580_/Y _3355_/R vdd gnd BUFX2
XBUFX2_insert11 RDY _3022_/A vdd gnd BUFX2
XFILL_1__2078_ gnd vdd FILL
XFILL_2__2960_ gnd vdd FILL
XBUFX2_insert66 _3198_/Y _3232_/B vdd gnd BUFX2
XBUFX2_insert44 _1716_/Y _2701_/B vdd gnd BUFX2
XBUFX2_insert55 _1733_/Y _2589_/A vdd gnd BUFX2
XBUFX2_insert88 _1729_/Y _2212_/A vdd gnd BUFX2
XFILL_2__1911_ gnd vdd FILL
XFILL_7__3585_ gnd vdd FILL
XFILL_7__2605_ gnd vdd FILL
XBUFX2_insert77 _1694_/Y _2293_/A vdd gnd BUFX2
XFILL_2__2891_ gnd vdd FILL
XFILL_4__2827_ gnd vdd FILL
XFILL_7__2536_ gnd vdd FILL
XFILL_2__1842_ gnd vdd FILL
XFILL_4__2758_ gnd vdd FILL
XFILL_4__1709_ gnd vdd FILL
XFILL_7__2467_ gnd vdd FILL
XFILL_2__1773_ gnd vdd FILL
XFILL_8_BUFX2_insert14 gnd vdd FILL
XFILL_8_BUFX2_insert58 gnd vdd FILL
XFILL_2__3512_ gnd vdd FILL
XFILL_7__2398_ gnd vdd FILL
XFILL_4__2689_ gnd vdd FILL
XFILL_5__3221_ gnd vdd FILL
XFILL_8_BUFX2_insert25 gnd vdd FILL
XFILL_8_BUFX2_insert47 gnd vdd FILL
XFILL_2__3443_ gnd vdd FILL
XFILL_8_BUFX2_insert69 gnd vdd FILL
XFILL_5__3152_ gnd vdd FILL
XFILL_2__3374_ gnd vdd FILL
XFILL_7__3019_ gnd vdd FILL
XFILL_5__3083_ gnd vdd FILL
XFILL_5__2103_ gnd vdd FILL
XFILL_5__2034_ gnd vdd FILL
XFILL_2__2325_ gnd vdd FILL
XFILL_2__2256_ gnd vdd FILL
XFILL_0__3010_ gnd vdd FILL
XFILL_2__2187_ gnd vdd FILL
XFILL_8__2714_ gnd vdd FILL
XFILL_5__2936_ gnd vdd FILL
XFILL_3__1951_ gnd vdd FILL
XFILL_8__2645_ gnd vdd FILL
XFILL_5__2867_ gnd vdd FILL
XFILL_8__2576_ gnd vdd FILL
X_2520_ _3570_/Q _3030_/C vdd gnd INVX1
XFILL_5__2798_ gnd vdd FILL
XFILL_3__1882_ gnd vdd FILL
XFILL_5__1818_ gnd vdd FILL
X_2451_ _2510_/D _2502_/C vdd gnd INVX2
XFILL_5__1749_ gnd vdd FILL
XFILL182850x163950 gnd vdd FILL
XFILL_3__3552_ gnd vdd FILL
X_2382_ _2795_/A _2409_/C _2717_/C _2425_/B vdd gnd OAI21X1
XFILL_3__2503_ gnd vdd FILL
XFILL_3__3483_ gnd vdd FILL
XFILL_8__3128_ gnd vdd FILL
XFILL_5__3419_ gnd vdd FILL
XFILL_6__2212_ gnd vdd FILL
XFILL_0__2725_ gnd vdd FILL
XFILL_6__3192_ gnd vdd FILL
X_3003_ _3003_/A _3369_/Y _3003_/S _3005_/B vdd gnd MUX2X1
XFILL_6__2143_ gnd vdd FILL
XFILL_3__2434_ gnd vdd FILL
XFILL_8__3059_ gnd vdd FILL
XFILL_3__2365_ gnd vdd FILL
XFILL_0__2656_ gnd vdd FILL
XFILL_6__2074_ gnd vdd FILL
XFILL_0__2587_ gnd vdd FILL
XFILL_3__2296_ gnd vdd FILL
XFILL_1__3050_ gnd vdd FILL
XFILL_1__2001_ gnd vdd FILL
XFILL_0__3208_ gnd vdd FILL
XFILL_6__2976_ gnd vdd FILL
XFILL_0__3139_ gnd vdd FILL
XFILL_6__1927_ gnd vdd FILL
XFILL_4__1991_ gnd vdd FILL
XFILL_6__1858_ gnd vdd FILL
X_2718_ _2718_/A _2718_/B _2718_/C _2720_/C vdd gnd NOR3X1
XFILL_1__2903_ gnd vdd FILL
XFILL_7__3370_ gnd vdd FILL
XFILL_6__3528_ gnd vdd FILL
XFILL_7__2321_ gnd vdd FILL
XFILL_4__3592_ gnd vdd FILL
XFILL_4__2612_ gnd vdd FILL
XFILL_6__1789_ gnd vdd FILL
X_2649_ _2741_/C _2653_/A vdd gnd INVX1
XFILL_1__2834_ gnd vdd FILL
XFILL_4__2543_ gnd vdd FILL
XFILL_6__3459_ gnd vdd FILL
XFILL_7__2252_ gnd vdd FILL
XFILL_1__2765_ gnd vdd FILL
XFILL_7__2183_ gnd vdd FILL
XFILL_9__2119_ gnd vdd FILL
XFILL_4__2474_ gnd vdd FILL
XFILL_1__1716_ gnd vdd FILL
XFILL_1__2696_ gnd vdd FILL
XFILL_2__3090_ gnd vdd FILL
XFILL_2__2110_ gnd vdd FILL
XFILL_2__2041_ gnd vdd FILL
XFILL_4__3026_ gnd vdd FILL
XFILL_7__1967_ gnd vdd FILL
XFILL_1__3179_ gnd vdd FILL
XFILL_7__1898_ gnd vdd FILL
XFILL_8__2430_ gnd vdd FILL
XFILL_5__2721_ gnd vdd FILL
XFILL_2__2943_ gnd vdd FILL
XFILL_5__2652_ gnd vdd FILL
XFILL_8__2361_ gnd vdd FILL
XFILL_2__2874_ gnd vdd FILL
XFILL_7__3499_ gnd vdd FILL
XFILL_2__1825_ gnd vdd FILL
XFILL_5__2583_ gnd vdd FILL
XFILL_7__2519_ gnd vdd FILL
XFILL_8__2292_ gnd vdd FILL
XFILL_2__1756_ gnd vdd FILL
XFILL_5__3204_ gnd vdd FILL
XFILL_0__2510_ gnd vdd FILL
XFILL_5__3135_ gnd vdd FILL
XFILL_0__3490_ gnd vdd FILL
XFILL_2__3426_ gnd vdd FILL
XFILL_3__2150_ gnd vdd FILL
XFILL_0__2441_ gnd vdd FILL
XFILL_0__2372_ gnd vdd FILL
XFILL_5__3066_ gnd vdd FILL
XFILL_2__2308_ gnd vdd FILL
XFILL_5__2017_ gnd vdd FILL
XFILL_3__2081_ gnd vdd FILL
XFILL_6__2830_ gnd vdd FILL
X_1951_ _2490_/A _2412_/B vdd gnd INVX1
XFILL_2__2239_ gnd vdd FILL
XFILL_4_BUFX2_insert23 gnd vdd FILL
X_1882_ _2462_/A _1916_/B vdd gnd INVX1
XFILL_4_BUFX2_insert12 gnd vdd FILL
XFILL_4_BUFX2_insert56 gnd vdd FILL
XFILL_4_BUFX2_insert45 gnd vdd FILL
XFILL_6__2761_ gnd vdd FILL
XFILL_5__2919_ gnd vdd FILL
X_3552_ _3552_/A _3552_/B _3552_/C _3573_/D vdd gnd OAI21X1
XFILL_3__2983_ gnd vdd FILL
XFILL_4_BUFX2_insert78 gnd vdd FILL
XFILL_6__1712_ gnd vdd FILL
XFILL_6__2692_ gnd vdd FILL
XFILL_8__2628_ gnd vdd FILL
XFILL_4_BUFX2_insert67 gnd vdd FILL
XFILL_4_BUFX2_insert89 gnd vdd FILL
X_2503_ _3084_/A _2503_/B _2503_/C _2504_/C vdd gnd OAI21X1
XFILL_3__1934_ gnd vdd FILL
XFILL_3__1865_ gnd vdd FILL
X_3483_ _3525_/A _3483_/B _3552_/B vdd gnd XOR2X1
XFILL_8__2559_ gnd vdd FILL
X_2434_ _2434_/A _3183_/C _2434_/C _2436_/A vdd gnd NAND3X1
X_2365_ _2966_/A _3189_/A _2365_/C _2407_/A vdd gnd OAI21X1
XFILL_3__1796_ gnd vdd FILL
XFILL_3__3535_ gnd vdd FILL
XFILL_3__3466_ gnd vdd FILL
X_2296_ _2296_/A _2296_/B _2303_/A vdd gnd NAND2X1
XFILL_1__2550_ gnd vdd FILL
XFILL_3__2417_ gnd vdd FILL
XFILL_1__2481_ gnd vdd FILL
XFILL_0__2708_ gnd vdd FILL
XFILL_6__3175_ gnd vdd FILL
XFILL_3__3397_ gnd vdd FILL
XFILL_4__2190_ gnd vdd FILL
XFILL_6__2126_ gnd vdd FILL
XFILL_0__2639_ gnd vdd FILL
XFILL_3__2348_ gnd vdd FILL
XFILL_6__2057_ gnd vdd FILL
XFILL_1__3102_ gnd vdd FILL
XFILL_3__2279_ gnd vdd FILL
XFILL_7__2870_ gnd vdd FILL
XFILL_1__3033_ gnd vdd FILL
XFILL_7__1821_ gnd vdd FILL
XFILL_6__2959_ gnd vdd FILL
XFILL_7__1752_ gnd vdd FILL
XFILL_8_BUFX2_insert0 gnd vdd FILL
XFILL_4__1974_ gnd vdd FILL
XFILL_7__3422_ gnd vdd FILL
XFILL_1__2817_ gnd vdd FILL
XFILL_7__2304_ gnd vdd FILL
XFILL_7__2235_ gnd vdd FILL
XFILL_2__2590_ gnd vdd FILL
XFILL_4__2526_ gnd vdd FILL
XFILL_4__2457_ gnd vdd FILL
XFILL_1__2748_ gnd vdd FILL
XFILL_7__2166_ gnd vdd FILL
XFILL_1__2679_ gnd vdd FILL
XFILL_4__2388_ gnd vdd FILL
XFILL_2__3211_ gnd vdd FILL
XFILL_7__2097_ gnd vdd FILL
XFILL_8__1930_ gnd vdd FILL
XFILL_2__3142_ gnd vdd FILL
XFILL_4__3009_ gnd vdd FILL
XFILL_2__3073_ gnd vdd FILL
XFILL_8__1861_ gnd vdd FILL
XFILL_2__2024_ gnd vdd FILL
XFILL_7__2999_ gnd vdd FILL
XFILL_8__3600_ gnd vdd FILL
XFILL_8__1792_ gnd vdd FILL
XFILL_8__3531_ gnd vdd FILL
XFILL_8__3462_ gnd vdd FILL
XFILL_5__2704_ gnd vdd FILL
XFILL_2__2926_ gnd vdd FILL
XFILL_0__2990_ gnd vdd FILL
XFILL_8__3393_ gnd vdd FILL
XFILL_8__2413_ gnd vdd FILL
XFILL_0__1941_ gnd vdd FILL
XFILL_8__2344_ gnd vdd FILL
XFILL_5__2635_ gnd vdd FILL
XFILL_2__2857_ gnd vdd FILL
XFILL_5__2566_ gnd vdd FILL
XFILL_0__1872_ gnd vdd FILL
XFILL_2__2788_ gnd vdd FILL
XFILL_8__2275_ gnd vdd FILL
XFILL_2__1808_ gnd vdd FILL
X_2150_ _2278_/A _3176_/B _2150_/C _2154_/B vdd gnd OAI21X1
XFILL_5__2497_ gnd vdd FILL
XFILL_2__1739_ gnd vdd FILL
XFILL_0__3542_ gnd vdd FILL
X_2081_ _2081_/A _2902_/A _2305_/B vdd gnd NOR2X1
XFILL_0__3473_ gnd vdd FILL
XFILL_2__3409_ gnd vdd FILL
XFILL_3__2202_ gnd vdd FILL
XFILL_5__3118_ gnd vdd FILL
XFILL_0__2424_ gnd vdd FILL
XFILL_3__3182_ gnd vdd FILL
XFILL_5__3049_ gnd vdd FILL
XFILL_3__2133_ gnd vdd FILL
XFILL_4_CLKBUF1_insert35 gnd vdd FILL
XFILL_3__2064_ gnd vdd FILL
X_2983_ _3017_/A _2986_/B vdd gnd INVX1
XFILL_0__2355_ gnd vdd FILL
XFILL_0__2286_ gnd vdd FILL
X_1934_ _3358_/Q _2691_/A _2715_/C vdd gnd NAND2X1
XFILL_6__2813_ gnd vdd FILL
X_1865_ _3287_/Q _2993_/B _1873_/B vdd gnd NAND2X1
XFILL_6__2744_ gnd vdd FILL
XFILL184050x171750 gnd vdd FILL
XFILL184350x163950 gnd vdd FILL
XFILL_3__2966_ gnd vdd FILL
X_1796_ _1796_/A _1796_/B _1815_/C vdd gnd NOR2X1
X_3535_ _3535_/A _3535_/B _3535_/C _3536_/A vdd gnd NAND3X1
XFILL_3__1917_ gnd vdd FILL
XFILL_9__2384_ gnd vdd FILL
XFILL_1__1981_ gnd vdd FILL
XFILL_6__2675_ gnd vdd FILL
X_3466_ _3514_/A _3466_/B _3466_/C _3467_/B vdd gnd OAI21X1
XFILL_3__2897_ gnd vdd FILL
XFILL_4__1690_ gnd vdd FILL
X_2417_ _2423_/A _2506_/A _2422_/C vdd gnd NAND2X1
XFILL_3__1848_ gnd vdd FILL
X_3397_ _3445_/A _3403_/A _3397_/C _3455_/C _3399_/B vdd gnd AOI22X1
XFILL_3__1779_ gnd vdd FILL
XFILL_3__3518_ gnd vdd FILL
XFILL_4__2311_ gnd vdd FILL
X_2348_ _2348_/A _2348_/B _2350_/C vdd gnd AND2X2
XFILL_1__2602_ gnd vdd FILL
XFILL_1__3582_ gnd vdd FILL
XFILL_7__2020_ gnd vdd FILL
XFILL_0_BUFX2_insert21 gnd vdd FILL
X_2279_ _2279_/A _2279_/B _2279_/C _2280_/B vdd gnd AOI21X1
XFILL_0_BUFX2_insert10 gnd vdd FILL
XFILL_1__2533_ gnd vdd FILL
XFILL_6__3227_ gnd vdd FILL
XFILL_3__3449_ gnd vdd FILL
XFILL_4__2242_ gnd vdd FILL
XFILL_0_BUFX2_insert43 gnd vdd FILL
XFILL_0_BUFX2_insert65 gnd vdd FILL
XFILL_0_BUFX2_insert54 gnd vdd FILL
XFILL_6__3158_ gnd vdd FILL
XFILL_4__2173_ gnd vdd FILL
XFILL_1__2464_ gnd vdd FILL
XFILL_0_BUFX2_insert87 gnd vdd FILL
XFILL_0_BUFX2_insert76 gnd vdd FILL
XFILL_6__2109_ gnd vdd FILL
XFILL_6__3089_ gnd vdd FILL
XFILL_1__2395_ gnd vdd FILL
XFILL_7__2922_ gnd vdd FILL
XFILL_7__2853_ gnd vdd FILL
XFILL_1__3016_ gnd vdd FILL
XFILL_7__1804_ gnd vdd FILL
XFILL_7__2784_ gnd vdd FILL
XFILL_7__1735_ gnd vdd FILL
XFILL_4__1957_ gnd vdd FILL
XFILL_7__3405_ gnd vdd FILL
XFILL_4__1888_ gnd vdd FILL
XFILL_2__2711_ gnd vdd FILL
XFILL_5__2420_ gnd vdd FILL
XFILL_4__3558_ gnd vdd FILL
XFILL_5__2351_ gnd vdd FILL
XFILL_2__2642_ gnd vdd FILL
XFILL_4__2509_ gnd vdd FILL
XFILL_8__2060_ gnd vdd FILL
XFILL_2__2573_ gnd vdd FILL
XFILL_4__3489_ gnd vdd FILL
XFILL_5__2282_ gnd vdd FILL
XFILL_7__2218_ gnd vdd FILL
XFILL_7__3198_ gnd vdd FILL
XFILL_7__2149_ gnd vdd FILL
XFILL_8__2962_ gnd vdd FILL
XFILL_2__3125_ gnd vdd FILL
XFILL_8__2893_ gnd vdd FILL
XFILL_8__1913_ gnd vdd FILL
XFILL_0__2140_ gnd vdd FILL
XFILL_8__1844_ gnd vdd FILL
XFILL_2__3056_ gnd vdd FILL
XFILL_0__2071_ gnd vdd FILL
XFILL_8__1775_ gnd vdd FILL
XFILL_2__2007_ gnd vdd FILL
XFILL_3__2820_ gnd vdd FILL
XFILL_8__3514_ gnd vdd FILL
XFILL_5__1997_ gnd vdd FILL
XFILL_8__3445_ gnd vdd FILL
X_3320_ _3320_/D vdd _3347_/R _3573_/CLK _3320_/Q vdd gnd DFFSR
XFILL_6__2460_ gnd vdd FILL
XFILL_3__2751_ gnd vdd FILL
XFILL_2__2909_ gnd vdd FILL
XFILL_8__3376_ gnd vdd FILL
XFILL_0__2973_ gnd vdd FILL
XFILL_3__1702_ gnd vdd FILL
XFILL_3__2682_ gnd vdd FILL
XFILL_5__2618_ gnd vdd FILL
XFILL_8__2327_ gnd vdd FILL
XFILL_5__3598_ gnd vdd FILL
XFILL_6__2391_ gnd vdd FILL
X_3251_ _3251_/D vdd _3362_/R _3362_/CLK _3251_/Q vdd gnd DFFSR
XFILL_0__1924_ gnd vdd FILL
XFILL_8__2258_ gnd vdd FILL
X_2202_ _3259_/Q _2202_/B _2203_/B vdd gnd NOR2X1
XFILL_0__1855_ gnd vdd FILL
XFILL_5__2549_ gnd vdd FILL
X_3182_ _3238_/Q _3182_/B _3182_/C _3184_/B vdd gnd OAI21X1
X_2133_ _3022_/A _2582_/B _2134_/B vdd gnd NAND2X1
XFILL_0__3525_ gnd vdd FILL
XFILL_8__2189_ gnd vdd FILL
XFILL_6__3012_ gnd vdd FILL
XFILL_0__1786_ gnd vdd FILL
XFILL_7_BUFX2_insert82 gnd vdd FILL
XFILL_7_BUFX2_insert60 gnd vdd FILL
X_2064_ _3282_/Q _2066_/A _2275_/B vdd gnd NOR2X1
XFILL_7_BUFX2_insert71 gnd vdd FILL
XFILL_0__3456_ gnd vdd FILL
XFILL_7_BUFX2_insert93 gnd vdd FILL
XFILL_3__3165_ gnd vdd FILL
XFILL_1__2180_ gnd vdd FILL
XFILL_0__3387_ gnd vdd FILL
XFILL_3__2116_ gnd vdd FILL
XFILL_0__2407_ gnd vdd FILL
XFILL184350x175650 gnd vdd FILL
XFILL184650x167850 gnd vdd FILL
XFILL_3__3096_ gnd vdd FILL
XFILL_0__2338_ gnd vdd FILL
XFILL_9__1884_ gnd vdd FILL
X_2966_ _2966_/A _2966_/B _3296_/D _2968_/C vdd gnd OAI21X1
XFILL_3__2047_ gnd vdd FILL
XFILL_4__2860_ gnd vdd FILL
XFILL_0__2269_ gnd vdd FILL
X_1917_ _3324_/Q _3092_/A _1920_/A vdd gnd NAND2X1
X_2897_ _2897_/A _2897_/B _2897_/C _2898_/C vdd gnd OAI21X1
X_1848_ _3144_/B _3149_/C _3178_/B vdd gnd NAND2X1
XFILL_4__1811_ gnd vdd FILL
XFILL_4__2791_ gnd vdd FILL
XFILL_6__2727_ gnd vdd FILL
XFILL_3__2949_ gnd vdd FILL
XFILL_4__1742_ gnd vdd FILL
X_1779_ _3239_/Q _2612_/B vdd gnd INVX2
XFILL_6__2658_ gnd vdd FILL
X_3518_ _3518_/A _3518_/B _3534_/B _3534_/A _3523_/A vdd gnd AOI22X1
XFILL_1__1964_ gnd vdd FILL
XFILL_4__3412_ gnd vdd FILL
X_3449_ _3449_/A _3459_/A _3449_/C _3449_/D _3493_/A vdd gnd OAI22X1
XFILL_6__2589_ gnd vdd FILL
XFILL_1__1895_ gnd vdd FILL
XFILL_7__3121_ gnd vdd FILL
XFILL_7__3052_ gnd vdd FILL
XFILL_7__2003_ gnd vdd FILL
XFILL_1__3565_ gnd vdd FILL
XFILL_1__3496_ gnd vdd FILL
XFILL_1__2516_ gnd vdd FILL
XFILL_4__2225_ gnd vdd FILL
XFILL_1__2447_ gnd vdd FILL
XFILL_4__2156_ gnd vdd FILL
XFILL_7__2905_ gnd vdd FILL
XFILL_4__2087_ gnd vdd FILL
XFILL_1__2378_ gnd vdd FILL
XFILL_5__1920_ gnd vdd FILL
XFILL_7__2836_ gnd vdd FILL
XFILL_5__1851_ gnd vdd FILL
XFILL_7__2767_ gnd vdd FILL
XFILL_4__2989_ gnd vdd FILL
XFILL_7__1718_ gnd vdd FILL
XFILL_5__1782_ gnd vdd FILL
XFILL_5__3521_ gnd vdd FILL
XFILL_7__2698_ gnd vdd FILL
XFILL_8__3230_ gnd vdd FILL
XFILL_5__3452_ gnd vdd FILL
XFILL_5__2403_ gnd vdd FILL
XFILL_8__3161_ gnd vdd FILL
XFILL_8__2112_ gnd vdd FILL
XFILL_8__3092_ gnd vdd FILL
XFILL_5__3383_ gnd vdd FILL
XFILL_2__2625_ gnd vdd FILL
XFILL_8__2043_ gnd vdd FILL
XFILL_5__2334_ gnd vdd FILL
XFILL_5__2265_ gnd vdd FILL
XFILL_2__2556_ gnd vdd FILL
XFILL_2__2487_ gnd vdd FILL
XFILL_5__2196_ gnd vdd FILL
XFILL_0_BUFX2_insert2 gnd vdd FILL
XFILL_8__2945_ gnd vdd FILL
XFILL_6__1960_ gnd vdd FILL
X_2820_ _2927_/B _2926_/B vdd gnd INVX1
XFILL_2__3108_ gnd vdd FILL
XFILL_8__2876_ gnd vdd FILL
XFILL_0__3172_ gnd vdd FILL
XFILL_2__3039_ gnd vdd FILL
XFILL_8__1827_ gnd vdd FILL
XFILL_6__1891_ gnd vdd FILL
XFILL_0__2123_ gnd vdd FILL
X_2751_ _2751_/A _2751_/B _2757_/C _2753_/B vdd gnd OAI21X1
XFILL_0__2054_ gnd vdd FILL
X_1702_ _2768_/A DI[4] _1702_/C _2950_/A vdd gnd OAI21X1
X_2682_ _2682_/A _2682_/B _2682_/C _2708_/A vdd gnd NOR3X1
XFILL_6__3561_ gnd vdd FILL
XFILL_8__1758_ gnd vdd FILL
XFILL_3__2803_ gnd vdd FILL
XFILL_8__1689_ gnd vdd FILL
XFILL_6__2512_ gnd vdd FILL
XFILL_6__3492_ gnd vdd FILL
XFILL_8__3428_ gnd vdd FILL
XFILL_3__2734_ gnd vdd FILL
XFILL_0__2956_ gnd vdd FILL
X_3303_ _3303_/D _3346_/CLK _3303_/Q vdd gnd DFFPOSX1
XFILL184650x150 gnd vdd FILL
XFILL_6__2443_ gnd vdd FILL
XFILL_6__2374_ gnd vdd FILL
X_3234_ _3234_/D vdd _3363_/R _3363_/CLK _3234_/Q vdd gnd DFFSR
XFILL_0__1907_ gnd vdd FILL
XFILL_3__2665_ gnd vdd FILL
XFILL_0__2887_ gnd vdd FILL
XFILL_3__2596_ gnd vdd FILL
XFILL_0__1838_ gnd vdd FILL
X_3165_ _3165_/A _3166_/A _3167_/A vdd gnd NAND2X1
XFILL184650x179550 gnd vdd FILL
X_3096_ _3131_/A _3108_/B _3096_/C _3324_/D vdd gnd OAI21X1
XFILL_0__1769_ gnd vdd FILL
X_2116_ _2786_/A _2340_/A _2116_/C _2352_/A vdd gnd OAI21X1
XFILL_4__2010_ gnd vdd FILL
XFILL_0__3508_ gnd vdd FILL
XFILL_1__2301_ gnd vdd FILL
X_2047_ _2375_/A _3195_/B vdd gnd INVX1
XFILL_3__3217_ gnd vdd FILL
XFILL_0__3439_ gnd vdd FILL
XFILL_1__2232_ gnd vdd FILL
XFILL_3__3148_ gnd vdd FILL
XFILL_1__2163_ gnd vdd FILL
XFILL_3__3079_ gnd vdd FILL
XFILL_4__2912_ gnd vdd FILL
X_2949_ reset _2957_/C _3303_/Q _2950_/C vdd gnd OAI21X1
XFILL_1__2094_ gnd vdd FILL
XFILL_7__2621_ gnd vdd FILL
XFILL_4__2843_ gnd vdd FILL
XFILL_3_BUFX2_insert6 gnd vdd FILL
XFILL_7__2552_ gnd vdd FILL
XFILL_4__2774_ gnd vdd FILL
XFILL_3_BUFX2_insert91 gnd vdd FILL
XFILL_1__2996_ gnd vdd FILL
XFILL_3_BUFX2_insert80 gnd vdd FILL
XFILL_7__2483_ gnd vdd FILL
XFILL_4__1725_ gnd vdd FILL
XFILL_1__1947_ gnd vdd FILL
XFILL_9__3399_ gnd vdd FILL
XFILL_1__1878_ gnd vdd FILL
XFILL_7__3104_ gnd vdd FILL
XFILL_2__3390_ gnd vdd FILL
XFILL_2__2410_ gnd vdd FILL
XFILL_1__3548_ gnd vdd FILL
XFILL_7__3035_ gnd vdd FILL
XFILL_2__2341_ gnd vdd FILL
XFILL184050x74250 gnd vdd FILL
XFILL_5__2050_ gnd vdd FILL
XFILL_1__3479_ gnd vdd FILL
XFILL_2__2272_ gnd vdd FILL
XFILL_4__2208_ gnd vdd FILL
XFILL_4__3188_ gnd vdd FILL
XFILL_4__2139_ gnd vdd FILL
XFILL_8__2730_ gnd vdd FILL
XFILL_5__2952_ gnd vdd FILL
XFILL_8__2661_ gnd vdd FILL
XFILL_7__2819_ gnd vdd FILL
XFILL_5__2883_ gnd vdd FILL
XFILL_5__1903_ gnd vdd FILL
XFILL_5__1834_ gnd vdd FILL
XFILL_8__2592_ gnd vdd FILL
XFILL_5__1765_ gnd vdd FILL
XFILL_5__3504_ gnd vdd FILL
XFILL_0__2810_ gnd vdd FILL
XFILL_5__1696_ gnd vdd FILL
XFILL_8__3213_ gnd vdd FILL
XFILL_2__1987_ gnd vdd FILL
XFILL_5__3435_ gnd vdd FILL
XFILL_0__2741_ gnd vdd FILL
XFILL_8__3144_ gnd vdd FILL
XFILL_5__3366_ gnd vdd FILL
XFILL_3__2450_ gnd vdd FILL
XFILL_8__3075_ gnd vdd FILL
XFILL_5__2317_ gnd vdd FILL
XFILL_3__2381_ gnd vdd FILL
XFILL_2__3588_ gnd vdd FILL
XFILL_0__2672_ gnd vdd FILL
XFILL_2__2608_ gnd vdd FILL
XFILL_8__2026_ gnd vdd FILL
XFILL_6__2090_ gnd vdd FILL
XFILL_2__2539_ gnd vdd FILL
XFILL_5__2248_ gnd vdd FILL
XFILL_5__2179_ gnd vdd FILL
XFILL_3__3002_ gnd vdd FILL
XFILL_8__2928_ gnd vdd FILL
XFILL_6__2992_ gnd vdd FILL
XFILL_0__3224_ gnd vdd FILL
X_2803_ _3009_/A _2887_/A _2815_/B _2803_/D _3263_/D vdd gnd OAI22X1
XFILL_0__3155_ gnd vdd FILL
XFILL_6__1943_ gnd vdd FILL
XFILL_6__1874_ gnd vdd FILL
XFILL_8__2859_ gnd vdd FILL
XFILL_0__2106_ gnd vdd FILL
XFILL_0__3086_ gnd vdd FILL
X_2734_ _2767_/A _2734_/B _2734_/C _2734_/D _3250_/D vdd gnd OAI22X1
XFILL_0__2037_ gnd vdd FILL
X_2665_ _2674_/A _2674_/C _2668_/C vdd gnd NOR2X1
XFILL_1__2850_ gnd vdd FILL
XFILL_6__3544_ gnd vdd FILL
X_2596_ _2702_/B _3348_/Q _2598_/B vdd gnd AND2X2
XFILL_6__3475_ gnd vdd FILL
XFILL_1__1801_ gnd vdd FILL
XFILL_6__2426_ gnd vdd FILL
XFILL_4__2490_ gnd vdd FILL
XFILL_1__2781_ gnd vdd FILL
XFILL_3__2717_ gnd vdd FILL
XFILL_0__2939_ gnd vdd FILL
XFILL_1__1732_ gnd vdd FILL
XFILL_3__2648_ gnd vdd FILL
X_3217_ _3217_/A _3228_/B _3217_/C _3356_/D vdd gnd OAI21X1
XFILL_6__2357_ gnd vdd FILL
XFILL_4__3111_ gnd vdd FILL
XFILL_3__2579_ gnd vdd FILL
XFILL_1__3402_ gnd vdd FILL
XFILL_6__2288_ gnd vdd FILL
X_3148_ _3180_/A _3148_/B _3179_/A vdd gnd NOR2X1
XFILL_4__3042_ gnd vdd FILL
X_3079_ _3079_/A _3088_/S _3079_/C _3080_/A vdd gnd OAI21X1
XFILL_1__2215_ gnd vdd FILL
XFILL_1__3195_ gnd vdd FILL
XFILL_7__1983_ gnd vdd FILL
XFILL_1__2146_ gnd vdd FILL
XBUFX2_insert23 _2580_/Y _3345_/R vdd gnd BUFX2
XBUFX2_insert12 RDY _2342_/A vdd gnd BUFX2
XBUFX2_insert56 _3374_/Y _3553_/B vdd gnd BUFX2
XFILL_1__2077_ gnd vdd FILL
XBUFX2_insert45 _1716_/Y _3144_/B vdd gnd BUFX2
XFILL_2__2890_ gnd vdd FILL
XBUFX2_insert78 _1694_/Y _2341_/A vdd gnd BUFX2
XFILL_7__3584_ gnd vdd FILL
XFILL_7__2604_ gnd vdd FILL
XBUFX2_insert67 _3198_/Y _3230_/B vdd gnd BUFX2
XBUFX2_insert89 _1729_/Y _2453_/A vdd gnd BUFX2
XFILL_2__1910_ gnd vdd FILL
XFILL_4__2826_ gnd vdd FILL
XFILL_7__2535_ gnd vdd FILL
XFILL_2__1841_ gnd vdd FILL
XFILL_7__2466_ gnd vdd FILL
XFILL_4__2757_ gnd vdd FILL
XFILL_1__2979_ gnd vdd FILL
XFILL_2__1772_ gnd vdd FILL
XFILL_4__1708_ gnd vdd FILL
XFILL_4__2688_ gnd vdd FILL
XFILL_8_BUFX2_insert15 gnd vdd FILL
XFILL_8_BUFX2_insert26 gnd vdd FILL
XFILL_2__3511_ gnd vdd FILL
XFILL_8_BUFX2_insert48 gnd vdd FILL
XFILL_7__2397_ gnd vdd FILL
XFILL_5__3220_ gnd vdd FILL
XFILL_8_BUFX2_insert59 gnd vdd FILL
XFILL_2__3442_ gnd vdd FILL
XFILL_5__3151_ gnd vdd FILL
XFILL_5__3082_ gnd vdd FILL
XFILL_2__3373_ gnd vdd FILL
XFILL_7__3018_ gnd vdd FILL
XFILL_5__2102_ gnd vdd FILL
XFILL_5__2033_ gnd vdd FILL
XFILL_2__2324_ gnd vdd FILL
XFILL_2__2255_ gnd vdd FILL
XFILL_2__2186_ gnd vdd FILL
XFILL_8__2713_ gnd vdd FILL
XFILL_5__2935_ gnd vdd FILL
XFILL_3__1950_ gnd vdd FILL
XFILL_8__2644_ gnd vdd FILL
XFILL_5__2866_ gnd vdd FILL
XFILL_8__2575_ gnd vdd FILL
XFILL_3__1881_ gnd vdd FILL
XFILL_5__2797_ gnd vdd FILL
X_2450_ _2563_/A _2538_/B _2510_/D vdd gnd NOR2X1
XFILL_5__1817_ gnd vdd FILL
XFILL_5__1748_ gnd vdd FILL
XFILL_3__3551_ gnd vdd FILL
X_2381_ _3261_/Q _2795_/A vdd gnd INVX1
XFILL_3__3482_ gnd vdd FILL
XFILL_6__2211_ gnd vdd FILL
XFILL_3__2502_ gnd vdd FILL
XFILL_8__3127_ gnd vdd FILL
XFILL_5__3418_ gnd vdd FILL
XFILL_0__2724_ gnd vdd FILL
XFILL_6__3191_ gnd vdd FILL
XFILL_3__2433_ gnd vdd FILL
XFILL_8__3058_ gnd vdd FILL
X_3002_ _3017_/A _3002_/B _3002_/C _3003_/A vdd gnd OAI21X1
XFILL_6__2142_ gnd vdd FILL
XFILL_0__2655_ gnd vdd FILL
XFILL_6__2073_ gnd vdd FILL
XFILL_3__2364_ gnd vdd FILL
XFILL_3__2295_ gnd vdd FILL
XFILL_0__2586_ gnd vdd FILL
XFILL_8__2009_ gnd vdd FILL
XFILL_1__2000_ gnd vdd FILL
XFILL_0__3207_ gnd vdd FILL
XFILL_6__2975_ gnd vdd FILL
XFILL_4__1990_ gnd vdd FILL
XFILL_0__3138_ gnd vdd FILL
XFILL_6__1926_ gnd vdd FILL
XFILL_6__1857_ gnd vdd FILL
XFILL_0__3069_ gnd vdd FILL
X_2717_ _3056_/A _2717_/B _2717_/C _2718_/B vdd gnd OAI21X1
XFILL_1__2902_ gnd vdd FILL
XFILL_6__1788_ gnd vdd FILL
XFILL_6__3527_ gnd vdd FILL
XFILL_4__3591_ gnd vdd FILL
XFILL_7__2320_ gnd vdd FILL
X_2648_ _2768_/A _2648_/B _2648_/C _3243_/D vdd gnd OAI21X1
XFILL_4__2611_ gnd vdd FILL
XFILL_1__2833_ gnd vdd FILL
X_2579_ _2866_/A _2579_/B _3521_/A vdd gnd NOR2X1
XFILL_4__2542_ gnd vdd FILL
XFILL_6__3458_ gnd vdd FILL
XFILL_7__2251_ gnd vdd FILL
XFILL_1__2764_ gnd vdd FILL
XFILL_6__3389_ gnd vdd FILL
XFILL_7__2182_ gnd vdd FILL
XFILL_4__2473_ gnd vdd FILL
XFILL_1__1715_ gnd vdd FILL
XFILL_6__2409_ gnd vdd FILL
XFILL_1__2695_ gnd vdd FILL
XFILL_4__3025_ gnd vdd FILL
XFILL_2__2040_ gnd vdd FILL
XFILL_7__1966_ gnd vdd FILL
XFILL_1__3178_ gnd vdd FILL
XFILL_7__1897_ gnd vdd FILL
XFILL_1__2129_ gnd vdd FILL
XFILL_2__2942_ gnd vdd FILL
XFILL_5__2720_ gnd vdd FILL
XFILL_8__2360_ gnd vdd FILL
XFILL_5__2651_ gnd vdd FILL
XFILL_4__2809_ gnd vdd FILL
XFILL_2__2873_ gnd vdd FILL
XFILL_5__2582_ gnd vdd FILL
XFILL_7__3498_ gnd vdd FILL
XFILL_2__1824_ gnd vdd FILL
XFILL_7__2518_ gnd vdd FILL
XFILL_8__2291_ gnd vdd FILL
XFILL_2__1755_ gnd vdd FILL
XFILL_7__2449_ gnd vdd FILL
XFILL_5__3203_ gnd vdd FILL
XFILL_5__3134_ gnd vdd FILL
XFILL_2__3425_ gnd vdd FILL
XFILL_0__2440_ gnd vdd FILL
XFILL_0__2371_ gnd vdd FILL
XFILL_5__3065_ gnd vdd FILL
XFILL_2__2307_ gnd vdd FILL
XFILL_3__2080_ gnd vdd FILL
XFILL_5__2016_ gnd vdd FILL
X_1950_ _1950_/A _1950_/B _1950_/C _2490_/A vdd gnd NAND3X1
XFILL_2__2238_ gnd vdd FILL
X_1881_ _1881_/A _1881_/B _1881_/C _2462_/A vdd gnd NAND3X1
XFILL_2__2169_ gnd vdd FILL
XFILL_4_BUFX2_insert24 gnd vdd FILL
XFILL_4_BUFX2_insert13 gnd vdd FILL
XFILL_4_BUFX2_insert57 gnd vdd FILL
XFILL_4_BUFX2_insert46 gnd vdd FILL
XFILL_6__2760_ gnd vdd FILL
XFILL_5__2918_ gnd vdd FILL
X_3551_ _3573_/Q _3552_/A _3552_/C vdd gnd NAND2X1
XFILL_4_BUFX2_insert79 gnd vdd FILL
XFILL_3__2982_ gnd vdd FILL
XFILL_6__1711_ gnd vdd FILL
XFILL_6__2691_ gnd vdd FILL
XFILL_4_BUFX2_insert68 gnd vdd FILL
XFILL_8__2627_ gnd vdd FILL
XFILL_5__2849_ gnd vdd FILL
X_2502_ _3296_/D _2502_/B _2502_/C _3354_/Q _2503_/C vdd gnd AOI22X1
XFILL_3__1933_ gnd vdd FILL
X_3482_ _3482_/A _3482_/B _3526_/A _3497_/B _3525_/A vdd gnd AOI22X1
XFILL_3__1864_ gnd vdd FILL
XFILL_8__2558_ gnd vdd FILL
XFILL_8__2489_ gnd vdd FILL
XFILL_3__3603_ gnd vdd FILL
X_2433_ _2433_/A _2433_/B _2434_/C vdd gnd NOR2X1
XFILL_3__3534_ gnd vdd FILL
X_2364_ _2364_/A _2365_/C vdd gnd INVX1
XFILL_3__1795_ gnd vdd FILL
XFILL_3__3465_ gnd vdd FILL
X_2295_ _2295_/A _2336_/A _2296_/A vdd gnd NOR2X1
XFILL_0__2707_ gnd vdd FILL
XFILL_6__3174_ gnd vdd FILL
XFILL_3__3396_ gnd vdd FILL
XFILL_3__2416_ gnd vdd FILL
XFILL_6__2125_ gnd vdd FILL
XFILL_1__2480_ gnd vdd FILL
XFILL_3__2347_ gnd vdd FILL
XFILL_0__2638_ gnd vdd FILL
XFILL_6__2056_ gnd vdd FILL
XFILL_0__2569_ gnd vdd FILL
XFILL_1__3101_ gnd vdd FILL
XFILL_3__2278_ gnd vdd FILL
XFILL_1__3032_ gnd vdd FILL
XFILL_7__1820_ gnd vdd FILL
XFILL_6__2958_ gnd vdd FILL
XFILL_7__1751_ gnd vdd FILL
XFILL_8_BUFX2_insert1 gnd vdd FILL
XFILL_4__1973_ gnd vdd FILL
XFILL_6__1909_ gnd vdd FILL
XFILL_6__2889_ gnd vdd FILL
XFILL_7__3421_ gnd vdd FILL
XFILL_1__2816_ gnd vdd FILL
XFILL_7__2303_ gnd vdd FILL
XFILL_4__2525_ gnd vdd FILL
XFILL_7__2234_ gnd vdd FILL
XFILL_4__2456_ gnd vdd FILL
XFILL_1__2747_ gnd vdd FILL
XFILL_7__2165_ gnd vdd FILL
XFILL_1__2678_ gnd vdd FILL
XFILL_4__2387_ gnd vdd FILL
XFILL_2__3210_ gnd vdd FILL
XFILL_7__2096_ gnd vdd FILL
XFILL_2__3141_ gnd vdd FILL
XFILL_8__1860_ gnd vdd FILL
XFILL_4__3008_ gnd vdd FILL
XFILL_2__3072_ gnd vdd FILL
XFILL_2__2023_ gnd vdd FILL
XFILL_7__2998_ gnd vdd FILL
XFILL_8__1791_ gnd vdd FILL
XFILL_8__3530_ gnd vdd FILL
XFILL_7__1949_ gnd vdd FILL
XFILL_8__3461_ gnd vdd FILL
XFILL_5__2703_ gnd vdd FILL
XFILL_2__2925_ gnd vdd FILL
XFILL_8__3392_ gnd vdd FILL
XFILL_8__2412_ gnd vdd FILL
XFILL_0__1940_ gnd vdd FILL
XFILL_2__2856_ gnd vdd FILL
XFILL182250x105450 gnd vdd FILL
XFILL_8__2343_ gnd vdd FILL
XFILL_5__2634_ gnd vdd FILL
XFILL_0__1871_ gnd vdd FILL
XFILL_8__2274_ gnd vdd FILL
XFILL_2__1807_ gnd vdd FILL
XFILL_5__2565_ gnd vdd FILL
XFILL_2__2787_ gnd vdd FILL
XFILL_5__2496_ gnd vdd FILL
XFILL_2__1738_ gnd vdd FILL
X_2080_ _2933_/B _2845_/A _2081_/A vdd gnd NAND2X1
XFILL_0__3541_ gnd vdd FILL
XFILL_0__3472_ gnd vdd FILL
XFILL_2__3408_ gnd vdd FILL
XFILL_3__2201_ gnd vdd FILL
XFILL_5__3117_ gnd vdd FILL
XFILL_0__2423_ gnd vdd FILL
XFILL_3__3181_ gnd vdd FILL
XFILL_5__3048_ gnd vdd FILL
XFILL_3__2132_ gnd vdd FILL
XFILL_0__2354_ gnd vdd FILL
X_2982_ _3267_/Q _2984_/C _3148_/B _2982_/D _2988_/A vdd gnd OAI22X1
XFILL_3__2063_ gnd vdd FILL
XFILL_4_CLKBUF1_insert36 gnd vdd FILL
XFILL_0__2285_ gnd vdd FILL
X_1933_ _2594_/B _2781_/A _1933_/C _2691_/A vdd gnd NOR3X1
XFILL_6__2812_ gnd vdd FILL
XFILL_8__1989_ gnd vdd FILL
X_1864_ _2968_/A _2993_/B vdd gnd INVX2
X_3603_ _3603_/A WE vdd gnd BUFX2
XFILL_6__2743_ gnd vdd FILL
XFILL_3__2965_ gnd vdd FILL
X_1795_ _2108_/A _3189_/A _1984_/B _1796_/B vdd gnd OAI21X1
X_3534_ _3534_/A _3534_/B _3536_/B vdd gnd NAND2X1
XFILL_3__1916_ gnd vdd FILL
XFILL_1__1980_ gnd vdd FILL
XFILL_6__2674_ gnd vdd FILL
X_3465_ _3514_/A _3514_/B _3473_/B _3474_/B vdd gnd OAI21X1
XFILL_3__2896_ gnd vdd FILL
X_2416_ _2416_/A _2416_/B _2416_/C _3600_/A vdd gnd OAI21X1
XFILL_3__1847_ gnd vdd FILL
X_3396_ _3404_/B _3398_/B _3397_/C vdd gnd NAND2X1
XFILL_3__1778_ gnd vdd FILL
XFILL_1__2601_ gnd vdd FILL
XFILL_3__3517_ gnd vdd FILL
XFILL_4__2310_ gnd vdd FILL
X_2347_ _2347_/A _2347_/B _2347_/C _2348_/A vdd gnd AOI21X1
XFILL_1__3581_ gnd vdd FILL
XFILL_0_BUFX2_insert22 gnd vdd FILL
XFILL_4__2241_ gnd vdd FILL
X_2278_ _2278_/A _2449_/C _2329_/C _2279_/C vdd gnd OAI21X1
XFILL_0_BUFX2_insert11 gnd vdd FILL
XFILL_1__2532_ gnd vdd FILL
XFILL_6__3226_ gnd vdd FILL
XFILL_3__3448_ gnd vdd FILL
XFILL_1__2463_ gnd vdd FILL
XFILL_0_BUFX2_insert66 gnd vdd FILL
XFILL_0_BUFX2_insert44 gnd vdd FILL
XFILL_0_BUFX2_insert55 gnd vdd FILL
XFILL_6__3157_ gnd vdd FILL
XFILL_3__3379_ gnd vdd FILL
XFILL_6__3088_ gnd vdd FILL
XFILL_4__2172_ gnd vdd FILL
XFILL_0_BUFX2_insert88 gnd vdd FILL
XFILL183750x7950 gnd vdd FILL
XFILL_6__2108_ gnd vdd FILL
XFILL_0_BUFX2_insert77 gnd vdd FILL
XFILL_6__2039_ gnd vdd FILL
XFILL_1__2394_ gnd vdd FILL
XFILL_7__2921_ gnd vdd FILL
XFILL_7__2852_ gnd vdd FILL
XFILL_1__3015_ gnd vdd FILL
XFILL_7__1803_ gnd vdd FILL
XFILL_7__2783_ gnd vdd FILL
XFILL_7__1734_ gnd vdd FILL
XFILL_4__1956_ gnd vdd FILL
XFILL_7__3404_ gnd vdd FILL
XFILL_4__1887_ gnd vdd FILL
XFILL_2__2710_ gnd vdd FILL
XFILL_4__3557_ gnd vdd FILL
XFILL_5__2350_ gnd vdd FILL
XFILL_2__2641_ gnd vdd FILL
XFILL_2__2572_ gnd vdd FILL
XFILL_4__2508_ gnd vdd FILL
XFILL_4__3488_ gnd vdd FILL
XFILL_7__2217_ gnd vdd FILL
XFILL_5__2281_ gnd vdd FILL
XFILL_7__3197_ gnd vdd FILL
XFILL_7__2148_ gnd vdd FILL
XFILL_4__2439_ gnd vdd FILL
XFILL_7__2079_ gnd vdd FILL
XFILL_8__2961_ gnd vdd FILL
XFILL_2__3124_ gnd vdd FILL
XFILL_8__2892_ gnd vdd FILL
XFILL_8__1912_ gnd vdd FILL
XFILL_2__3055_ gnd vdd FILL
XFILL_8__1843_ gnd vdd FILL
XFILL_2__2006_ gnd vdd FILL
XFILL_0__2070_ gnd vdd FILL
XFILL182550x109350 gnd vdd FILL
XFILL_8__1774_ gnd vdd FILL
XFILL_8__3513_ gnd vdd FILL
XFILL182250x117150 gnd vdd FILL
XFILL_5__1996_ gnd vdd FILL
XFILL_8__3444_ gnd vdd FILL
XFILL_3__2750_ gnd vdd FILL
XFILL_0__2972_ gnd vdd FILL
XFILL_3__1701_ gnd vdd FILL
XFILL_2__2908_ gnd vdd FILL
XFILL_8__3375_ gnd vdd FILL
XFILL_6__2390_ gnd vdd FILL
XFILL_0__1923_ gnd vdd FILL
XFILL_3__2681_ gnd vdd FILL
XFILL_5__2617_ gnd vdd FILL
XFILL_2__2839_ gnd vdd FILL
XFILL_8__2326_ gnd vdd FILL
XFILL_5__3597_ gnd vdd FILL
X_3250_ _3250_/D vdd _3291_/R _3362_/CLK _3250_/Q vdd gnd DFFSR
XFILL_8__2257_ gnd vdd FILL
XFILL_0__1854_ gnd vdd FILL
X_2201_ _3308_/Q _2202_/B vdd gnd INVX1
X_3181_ _3181_/A _3181_/B _3186_/A vdd gnd NAND2X1
XFILL_5__2548_ gnd vdd FILL
X_2132_ _3568_/Q _3314_/Q _2582_/B vdd gnd XOR2X1
XFILL_5__2479_ gnd vdd FILL
XFILL_0__1785_ gnd vdd FILL
XFILL_0__3524_ gnd vdd FILL
XFILL_8__2188_ gnd vdd FILL
XFILL_6__3011_ gnd vdd FILL
XFILL_7_BUFX2_insert61 gnd vdd FILL
XFILL_7_BUFX2_insert50 gnd vdd FILL
XFILL_7_BUFX2_insert83 gnd vdd FILL
X_2063_ _3022_/A _2063_/B _2066_/B vdd gnd NAND2X1
XFILL_7_BUFX2_insert72 gnd vdd FILL
XFILL_0__3455_ gnd vdd FILL
XFILL_7_BUFX2_insert94 gnd vdd FILL
XFILL_3__3164_ gnd vdd FILL
XFILL_0__3386_ gnd vdd FILL
XFILL_3__2115_ gnd vdd FILL
XFILL_0__2406_ gnd vdd FILL
XFILL_3__3095_ gnd vdd FILL
XFILL_0__2337_ gnd vdd FILL
X_2965_ _3279_/Q _2965_/B _2991_/B _2971_/A vdd gnd OAI21X1
XFILL_3__2046_ gnd vdd FILL
XFILL_0__2268_ gnd vdd FILL
X_2896_ _2932_/B _2896_/B _2896_/C _2897_/A vdd gnd OAI21X1
X_1916_ _1986_/A _1916_/B _1916_/C _3521_/B vdd gnd OAI21X1
X_1847_ _2108_/A _2448_/B _3158_/B _1883_/A vdd gnd OAI21X1
XFILL_4__1810_ gnd vdd FILL
XFILL_0__2199_ gnd vdd FILL
XFILL_4__2790_ gnd vdd FILL
XFILL_6__2726_ gnd vdd FILL
X_3517_ _3535_/B _3534_/A vdd gnd INVX1
XFILL_3__2948_ gnd vdd FILL
X_1778_ _1778_/A _1778_/B _3466_/C vdd gnd OR2X2
XFILL_6__2657_ gnd vdd FILL
XFILL_4__1741_ gnd vdd FILL
XFILL_3__2879_ gnd vdd FILL
XFILL_1__1963_ gnd vdd FILL
XFILL_4__3411_ gnd vdd FILL
X_3448_ _3460_/B _3448_/B _3459_/A _3449_/D vdd gnd OAI21X1
XFILL_6__2588_ gnd vdd FILL
XFILL_1__1894_ gnd vdd FILL
XFILL_7__3120_ gnd vdd FILL
X_3379_ _3453_/B _3387_/B _3383_/B vdd gnd AND2X2
XFILL_7__3051_ gnd vdd FILL
XFILL_1__3564_ gnd vdd FILL
XFILL184650x11850 gnd vdd FILL
XFILL_7__2002_ gnd vdd FILL
XFILL_6__3209_ gnd vdd FILL
XFILL_1__2515_ gnd vdd FILL
XFILL_1__3495_ gnd vdd FILL
XFILL_4__2224_ gnd vdd FILL
XFILL_4__2155_ gnd vdd FILL
XFILL_1__2446_ gnd vdd FILL
XFILL_1__2377_ gnd vdd FILL
XFILL_7__2904_ gnd vdd FILL
XFILL_4__2086_ gnd vdd FILL
XFILL_7__2835_ gnd vdd FILL
XFILL_7__2766_ gnd vdd FILL
XFILL_5__1850_ gnd vdd FILL
XFILL_4__2988_ gnd vdd FILL
XFILL_7__1717_ gnd vdd FILL
XFILL_5__1781_ gnd vdd FILL
XFILL_4__1939_ gnd vdd FILL
XFILL_5__3520_ gnd vdd FILL
XFILL_7__2697_ gnd vdd FILL
XFILL_5__3451_ gnd vdd FILL
XFILL_5__2402_ gnd vdd FILL
XFILL_8__3160_ gnd vdd FILL
XFILL_8__3091_ gnd vdd FILL
XFILL_5__3382_ gnd vdd FILL
XFILL_8__2111_ gnd vdd FILL
XFILL_2__2624_ gnd vdd FILL
XFILL_8__2042_ gnd vdd FILL
XFILL_5__2333_ gnd vdd FILL
XFILL_5__2264_ gnd vdd FILL
XFILL_2__2555_ gnd vdd FILL
XFILL_2__2486_ gnd vdd FILL
XFILL_5__2195_ gnd vdd FILL
XFILL_0_BUFX2_insert3 gnd vdd FILL
XFILL_8__2944_ gnd vdd FILL
XFILL_2__3107_ gnd vdd FILL
XFILL_0__3171_ gnd vdd FILL
XFILL_8__2875_ gnd vdd FILL
XFILL_0__2122_ gnd vdd FILL
XFILL_2__3038_ gnd vdd FILL
X_2750_ _3295_/D _2772_/B _2750_/C _2757_/C vdd gnd AOI21X1
XFILL_6__1890_ gnd vdd FILL
XFILL_8__1826_ gnd vdd FILL
X_1701_ _2675_/A _3294_/Q _1702_/C vdd gnd OR2X2
XFILL_0__2053_ gnd vdd FILL
XFILL_8__1757_ gnd vdd FILL
X_2681_ _2771_/A _2681_/B _2681_/C _2682_/B vdd gnd NAND3X1
XFILL_5__1979_ gnd vdd FILL
XFILL_6__3560_ gnd vdd FILL
XFILL_3__2802_ gnd vdd FILL
XFILL_6__2511_ gnd vdd FILL
XFILL_8__1688_ gnd vdd FILL
XFILL_6__3491_ gnd vdd FILL
XFILL_8__3427_ gnd vdd FILL
XFILL_3__2733_ gnd vdd FILL
X_3302_ _3302_/D _3346_/CLK _3302_/Q vdd gnd DFFPOSX1
XFILL_0__2955_ gnd vdd FILL
XFILL_6__2442_ gnd vdd FILL
XFILL_8__2309_ gnd vdd FILL
XFILL_0__2886_ gnd vdd FILL
XFILL_6__2373_ gnd vdd FILL
X_3233_ _3233_/D vdd _3363_/R _3363_/CLK _3233_/Q vdd gnd DFFSR
XFILL_3__2664_ gnd vdd FILL
XFILL_0__1906_ gnd vdd FILL
XFILL_3__2595_ gnd vdd FILL
XFILL_0__1837_ gnd vdd FILL
X_3164_ _3164_/A _3173_/C _3169_/A vdd gnd AND2X2
X_3095_ _3115_/A _3107_/B _3324_/Q _3096_/C vdd gnd OAI21X1
XFILL_0__1768_ gnd vdd FILL
X_2115_ _2886_/A _2115_/B _2786_/A _2116_/C vdd gnd OAI21X1
XFILL_0__3507_ gnd vdd FILL
XFILL_1__2300_ gnd vdd FILL
X_2046_ _3165_/A _3156_/B _2375_/A vdd gnd NOR2X1
XFILL_3__3216_ gnd vdd FILL
XFILL_0__1699_ gnd vdd FILL
XFILL_0__3438_ gnd vdd FILL
XFILL_1__2231_ gnd vdd FILL
XFILL_3__3147_ gnd vdd FILL
XFILL_1__2162_ gnd vdd FILL
XFILL_3__3078_ gnd vdd FILL
XFILL_0__3369_ gnd vdd FILL
XFILL_4__2911_ gnd vdd FILL
X_2948_ _2948_/A _2956_/B _2948_/C _3302_/D vdd gnd OAI21X1
XFILL_3__2029_ gnd vdd FILL
XFILL_1__2093_ gnd vdd FILL
XFILL_7__2620_ gnd vdd FILL
XFILL_4__2842_ gnd vdd FILL
X_2879_ _2906_/A _2888_/B _3280_/Q _2882_/C vdd gnd OAI21X1
XFILL_7__2551_ gnd vdd FILL
XFILL_3_BUFX2_insert7 gnd vdd FILL
XFILL_6__2709_ gnd vdd FILL
XFILL_4__2773_ gnd vdd FILL
XFILL_3_BUFX2_insert92 gnd vdd FILL
XFILL_1__2995_ gnd vdd FILL
XFILL_7__2482_ gnd vdd FILL
XFILL_3_BUFX2_insert81 gnd vdd FILL
XFILL184650x23550 gnd vdd FILL
XFILL_4__1724_ gnd vdd FILL
XFILL_3_BUFX2_insert70 gnd vdd FILL
XFILL_1__1946_ gnd vdd FILL
XFILL_7__3103_ gnd vdd FILL
XFILL_1__1877_ gnd vdd FILL
XFILL_1__3547_ gnd vdd FILL
XFILL_7__3034_ gnd vdd FILL
XFILL_2__2340_ gnd vdd FILL
XFILL184350x58650 gnd vdd FILL
XFILL_1__3478_ gnd vdd FILL
XFILL_2__2271_ gnd vdd FILL
XFILL_4__2207_ gnd vdd FILL
XFILL_4__3187_ gnd vdd FILL
XFILL_1__2429_ gnd vdd FILL
XFILL_4__2138_ gnd vdd FILL
XFILL_4__2069_ gnd vdd FILL
XFILL_5__2951_ gnd vdd FILL
XFILL_8__2660_ gnd vdd FILL
XFILL_7__2818_ gnd vdd FILL
XFILL_5__2882_ gnd vdd FILL
XFILL_5__1902_ gnd vdd FILL
XFILL_8__2591_ gnd vdd FILL
XFILL_5__1833_ gnd vdd FILL
XFILL_7__2749_ gnd vdd FILL
XFILL_5__3503_ gnd vdd FILL
XFILL_5__1764_ gnd vdd FILL
XFILL_2__1986_ gnd vdd FILL
XFILL_5__1695_ gnd vdd FILL
XFILL_8__3212_ gnd vdd FILL
XFILL_8__3143_ gnd vdd FILL
XFILL_5__3434_ gnd vdd FILL
XFILL_0__2740_ gnd vdd FILL
XFILL_5__3365_ gnd vdd FILL
XFILL_8__3074_ gnd vdd FILL
XFILL_2__3587_ gnd vdd FILL
XFILL_3__2380_ gnd vdd FILL
XFILL_5__2316_ gnd vdd FILL
XFILL_2__2607_ gnd vdd FILL
XFILL_0__2671_ gnd vdd FILL
XFILL_8__2025_ gnd vdd FILL
XFILL_2__2538_ gnd vdd FILL
XFILL_5__2247_ gnd vdd FILL
XFILL_3__3001_ gnd vdd FILL
XFILL_2__2469_ gnd vdd FILL
XFILL_5__2178_ gnd vdd FILL
XFILL184050x109350 gnd vdd FILL
XFILL_0__3223_ gnd vdd FILL
XFILL_8__2927_ gnd vdd FILL
XFILL_6__2991_ gnd vdd FILL
XFILL_8__2858_ gnd vdd FILL
X_2802_ _2894_/A _2864_/C _2815_/B vdd gnd NAND2X1
XFILL_6__1942_ gnd vdd FILL
XFILL_0__3154_ gnd vdd FILL
XFILL_6__1873_ gnd vdd FILL
XFILL_0__3085_ gnd vdd FILL
X_2733_ _2741_/A _2733_/B _2767_/A _2734_/C vdd gnd OAI21X1
XFILL_8__1809_ gnd vdd FILL
XFILL_0__2105_ gnd vdd FILL
XFILL_0__2036_ gnd vdd FILL
XFILL_8__2789_ gnd vdd FILL
X_2664_ _2668_/B _2671_/B _2686_/B _2674_/A vdd gnd OAI21X1
XFILL_6__3543_ gnd vdd FILL
X_2595_ _3239_/Q _2770_/B _2670_/B _3570_/Q _2599_/A vdd gnd AOI22X1
XFILL_6__3474_ gnd vdd FILL
XFILL_1__2780_ gnd vdd FILL
XFILL_1__1800_ gnd vdd FILL
XFILL_6__2425_ gnd vdd FILL
XFILL_3__2716_ gnd vdd FILL
XFILL_1__1731_ gnd vdd FILL
XFILL_0__2938_ gnd vdd FILL
XFILL_9__2134_ gnd vdd FILL
XFILL_3__2647_ gnd vdd FILL
XFILL_0__2869_ gnd vdd FILL
XFILL_6__2356_ gnd vdd FILL
X_3216_ _3216_/A _3216_/B _3228_/B _3217_/C vdd gnd OAI21X1
XFILL_3__2578_ gnd vdd FILL
XFILL_4__3110_ gnd vdd FILL
XFILL_1__3401_ gnd vdd FILL
XFILL_6__2287_ gnd vdd FILL
X_3147_ _3147_/A _3147_/B _3147_/C _3180_/A vdd gnd OAI21X1
XFILL_4__3041_ gnd vdd FILL
X_3078_ _3083_/B _3083_/A _3078_/C _3079_/C vdd gnd OAI21X1
X_2029_ _2897_/C _2270_/A _2311_/A _2338_/A vdd gnd NAND3X1
XFILL_1__2214_ gnd vdd FILL
XFILL_7__1982_ gnd vdd FILL
XFILL_1__3194_ gnd vdd FILL
XFILL_1__2145_ gnd vdd FILL
XBUFX2_insert24 _2580_/Y _3353_/R vdd gnd BUFX2
XBUFX2_insert13 _1907_/Y _2717_/C vdd gnd BUFX2
XBUFX2_insert57 _3374_/Y _3550_/A vdd gnd BUFX2
XFILL_1__2076_ gnd vdd FILL
XBUFX2_insert46 _1716_/Y _2602_/A vdd gnd BUFX2
XFILL_7__2603_ gnd vdd FILL
XFILL184650x35250 gnd vdd FILL
XFILL_4__2825_ gnd vdd FILL
XBUFX2_insert79 _1694_/Y _2906_/A vdd gnd BUFX2
XFILL_7__3583_ gnd vdd FILL
XBUFX2_insert68 _3198_/Y _3227_/B vdd gnd BUFX2
XFILL_7__2534_ gnd vdd FILL
XFILL_2__1840_ gnd vdd FILL
XFILL_7__2465_ gnd vdd FILL
XFILL_4__2756_ gnd vdd FILL
XFILL_1__2978_ gnd vdd FILL
XFILL_2__1771_ gnd vdd FILL
XFILL_4__1707_ gnd vdd FILL
XFILL_4__2687_ gnd vdd FILL
XFILL_1__1929_ gnd vdd FILL
XFILL_2__3510_ gnd vdd FILL
XFILL_8_BUFX2_insert49 gnd vdd FILL
XFILL_7__2396_ gnd vdd FILL
XFILL_8_BUFX2_insert27 gnd vdd FILL
XFILL_8_BUFX2_insert16 gnd vdd FILL
XFILL_2__3441_ gnd vdd FILL
XFILL_2__3372_ gnd vdd FILL
XFILL_5__3150_ gnd vdd FILL
XFILL_5__3081_ gnd vdd FILL
XFILL_7__3017_ gnd vdd FILL
XFILL_2__2323_ gnd vdd FILL
XFILL_5__2101_ gnd vdd FILL
XFILL_5__2032_ gnd vdd FILL
XFILL_2__2254_ gnd vdd FILL
XFILL_2__2185_ gnd vdd FILL
XFILL_8__2712_ gnd vdd FILL
XFILL_5__2934_ gnd vdd FILL
XFILL_8__2643_ gnd vdd FILL
XFILL_5__2865_ gnd vdd FILL
XFILL_8__2574_ gnd vdd FILL
XFILL_3__1880_ gnd vdd FILL
XFILL_5__2796_ gnd vdd FILL
XFILL_5__1816_ gnd vdd FILL
XFILL_5__1747_ gnd vdd FILL
XFILL_3__3550_ gnd vdd FILL
XFILL_2__1969_ gnd vdd FILL
X_2380_ _3261_/Q _2409_/C _3003_/S _2427_/B vdd gnd OAI21X1
XFILL_3__3481_ gnd vdd FILL
XFILL_5__3417_ gnd vdd FILL
XFILL_6__2210_ gnd vdd FILL
XFILL_3__2501_ gnd vdd FILL
XFILL_8__3126_ gnd vdd FILL
XFILL_0__2723_ gnd vdd FILL
XFILL_3__2432_ gnd vdd FILL
XFILL_6__3190_ gnd vdd FILL
XFILL_8__3057_ gnd vdd FILL
X_3001_ _3291_/D _3017_/A _3002_/C vdd gnd NAND2X1
XFILL_6__2141_ gnd vdd FILL
XFILL_0__2654_ gnd vdd FILL
XFILL_6__2072_ gnd vdd FILL
XFILL_3__2363_ gnd vdd FILL
XFILL_8__2008_ gnd vdd FILL
XFILL_0__2585_ gnd vdd FILL
XFILL_3__2294_ gnd vdd FILL
XFILL183750x163950 gnd vdd FILL
XFILL183450x171750 gnd vdd FILL
XFILL_9__2752_ gnd vdd FILL
XFILL_6__2974_ gnd vdd FILL
XFILL_0__3206_ gnd vdd FILL
XFILL_0__3137_ gnd vdd FILL
XFILL_6__1925_ gnd vdd FILL
XFILL_0__3068_ gnd vdd FILL
XFILL_6__1856_ gnd vdd FILL
X_2716_ _3572_/Q _3056_/A vdd gnd INVX1
XFILL_1__2901_ gnd vdd FILL
XFILL_0__2019_ gnd vdd FILL
XFILL_6__1787_ gnd vdd FILL
X_2647_ _2741_/C _2653_/B _2648_/B vdd gnd XOR2X1
XFILL_6__3526_ gnd vdd FILL
XFILL_4__3590_ gnd vdd FILL
XFILL_4__2610_ gnd vdd FILL
X_2578_ _3275_/Q _2866_/A vdd gnd INVX1
XFILL_1__2832_ gnd vdd FILL
XFILL_4__2541_ gnd vdd FILL
XFILL_7__2250_ gnd vdd FILL
XFILL_6__3457_ gnd vdd FILL
XFILL_1__2763_ gnd vdd FILL
XFILL_6__3388_ gnd vdd FILL
XFILL_7__2181_ gnd vdd FILL
XFILL_4__2472_ gnd vdd FILL
XFILL_1__2694_ gnd vdd FILL
XFILL_1__1714_ gnd vdd FILL
XFILL_6__2408_ gnd vdd FILL
XFILL_6__2339_ gnd vdd FILL
XFILL_4__3024_ gnd vdd FILL
XFILL_7__1965_ gnd vdd FILL
XFILL_1__3177_ gnd vdd FILL
XFILL_7__1896_ gnd vdd FILL
XFILL_1__2128_ gnd vdd FILL
XFILL_2__2941_ gnd vdd FILL
XFILL_1__2059_ gnd vdd FILL
XFILL_7__3566_ gnd vdd FILL
XFILL_5__2650_ gnd vdd FILL
XFILL_4__2808_ gnd vdd FILL
XFILL_2__2872_ gnd vdd FILL
XFILL_7__2517_ gnd vdd FILL
XFILL_5__2581_ gnd vdd FILL
XFILL_7__3497_ gnd vdd FILL
XFILL_2__1823_ gnd vdd FILL
XFILL_8__2290_ gnd vdd FILL
XFILL_4__2739_ gnd vdd FILL
XFILL_2__1754_ gnd vdd FILL
XFILL_7__2448_ gnd vdd FILL
XFILL_7__2379_ gnd vdd FILL
XFILL_5__3202_ gnd vdd FILL
XFILL_5__3133_ gnd vdd FILL
XFILL_2__3424_ gnd vdd FILL
XFILL_0__2370_ gnd vdd FILL
XFILL_2__2306_ gnd vdd FILL
XFILL_5__3064_ gnd vdd FILL
XFILL_5__2015_ gnd vdd FILL
XFILL_2__2237_ gnd vdd FILL
XFILL_2__2168_ gnd vdd FILL
X_1880_ _3331_/Q _3110_/A _3092_/A _3323_/Q _1881_/C vdd gnd AOI22X1
XFILL_4_BUFX2_insert14 gnd vdd FILL
XFILL_4_BUFX2_insert25 gnd vdd FILL
XFILL_4_BUFX2_insert47 gnd vdd FILL
XFILL_2__2099_ gnd vdd FILL
X_3550_ _3550_/A _3550_/B _3550_/C _3572_/D vdd gnd OAI21X1
XFILL_5__2917_ gnd vdd FILL
XFILL_4_BUFX2_insert58 gnd vdd FILL
XFILL_3__2981_ gnd vdd FILL
XFILL_6__1710_ gnd vdd FILL
XFILL_6__2690_ gnd vdd FILL
XFILL_8__2626_ gnd vdd FILL
XFILL_4_BUFX2_insert69 gnd vdd FILL
XFILL_5__2848_ gnd vdd FILL
XFILL_3__1932_ gnd vdd FILL
X_2501_ _3576_/Q _3084_/A vdd gnd INVX1
X_3481_ _3526_/B _3497_/B vdd gnd INVX1
XFILL_3__1863_ gnd vdd FILL
XFILL_8__2557_ gnd vdd FILL
XFILL_3__3602_ gnd vdd FILL
XFILL_8__2488_ gnd vdd FILL
XFILL_5__2779_ gnd vdd FILL
X_2432_ _2432_/A _2602_/B _2434_/A vdd gnd NAND2X1
XFILL_3__3533_ gnd vdd FILL
X_2363_ _2453_/A _2781_/B _2364_/A vdd gnd NOR2X1
XFILL_3__1794_ gnd vdd FILL
XFILL_8__3109_ gnd vdd FILL
XFILL_3__3464_ gnd vdd FILL
XFILL_0__2706_ gnd vdd FILL
XFILL_6__3173_ gnd vdd FILL
X_2294_ _2294_/A _2294_/B _2342_/C _2295_/A vdd gnd OAI21X1
XFILL183750x175650 gnd vdd FILL
XFILL_3__3395_ gnd vdd FILL
XFILL_3__2415_ gnd vdd FILL
XFILL_6__2124_ gnd vdd FILL
XFILL_3__2346_ gnd vdd FILL
XFILL_0__2637_ gnd vdd FILL
XFILL_6__2055_ gnd vdd FILL
XFILL_0__2568_ gnd vdd FILL
XFILL_1__3100_ gnd vdd FILL
XFILL_3__2277_ gnd vdd FILL
XFILL_1__3031_ gnd vdd FILL
XFILL_0__2499_ gnd vdd FILL
XFILL_6__2957_ gnd vdd FILL
XFILL_7__1750_ gnd vdd FILL
XFILL_8_BUFX2_insert2 gnd vdd FILL
XFILL_6__2888_ gnd vdd FILL
XFILL_4__1972_ gnd vdd FILL
XFILL_6__1908_ gnd vdd FILL
XFILL_7__3420_ gnd vdd FILL
XFILL_6__1839_ gnd vdd FILL
XFILL_6__3509_ gnd vdd FILL
XFILL_1__2815_ gnd vdd FILL
XFILL_7__2302_ gnd vdd FILL
XFILL_4__2524_ gnd vdd FILL
XFILL_7__2233_ gnd vdd FILL
XFILL_4__2455_ gnd vdd FILL
XFILL_1__2746_ gnd vdd FILL
XFILL_7__2164_ gnd vdd FILL
XFILL_1__2677_ gnd vdd FILL
XFILL_4__2386_ gnd vdd FILL
XFILL_7__2095_ gnd vdd FILL
XFILL_2__3140_ gnd vdd FILL
XFILL_4__3007_ gnd vdd FILL
XFILL_2__3071_ gnd vdd FILL
XFILL_2__2022_ gnd vdd FILL
XFILL_7__2997_ gnd vdd FILL
XFILL_1__3229_ gnd vdd FILL
XFILL_8__1790_ gnd vdd FILL
XFILL_7__1948_ gnd vdd FILL
XFILL_8__3460_ gnd vdd FILL
XFILL_7__1879_ gnd vdd FILL
XFILL_5__2702_ gnd vdd FILL
XFILL_8__2411_ gnd vdd FILL
XFILL_2__2924_ gnd vdd FILL
XFILL_8__3391_ gnd vdd FILL
XFILL_5__2633_ gnd vdd FILL
XFILL_7__3549_ gnd vdd FILL
XFILL_2__2855_ gnd vdd FILL
XFILL_8__2342_ gnd vdd FILL
XFILL_0__1870_ gnd vdd FILL
XFILL_8__2273_ gnd vdd FILL
XFILL_5__2564_ gnd vdd FILL
XFILL_2__1806_ gnd vdd FILL
XFILL_2__2786_ gnd vdd FILL
XFILL_5__2495_ gnd vdd FILL
XFILL_2__1737_ gnd vdd FILL
XFILL_0__3540_ gnd vdd FILL
XFILL_0__3471_ gnd vdd FILL
XFILL_2__3407_ gnd vdd FILL
XFILL_3__2200_ gnd vdd FILL
XFILL_3__3180_ gnd vdd FILL
XFILL_5__3116_ gnd vdd FILL
XFILL_0__2422_ gnd vdd FILL
XFILL183150x74250 gnd vdd FILL
XFILL_5__3047_ gnd vdd FILL
XFILL_0__2353_ gnd vdd FILL
XFILL_3__2131_ gnd vdd FILL
XFILL_4_CLKBUF1_insert37 gnd vdd FILL
XFILL_3__2062_ gnd vdd FILL
X_2981_ _2981_/A _3176_/B _2995_/A _2982_/D vdd gnd AOI21X1
X_1932_ _2474_/A _1937_/B vdd gnd INVX1
XFILL_0__2284_ gnd vdd FILL
XFILL_8__1988_ gnd vdd FILL
XFILL_6__2811_ gnd vdd FILL
X_1863_ _1883_/A _1863_/B _3284_/Q _1874_/B vdd gnd OAI21X1
X_3602_ _3602_/A DO[7] vdd gnd BUFX2
XFILL_6__2742_ gnd vdd FILL
XFILL_3__2964_ gnd vdd FILL
X_1794_ _1794_/A _1891_/B _3189_/A vdd gnd NAND2X1
X_3533_ _3533_/A _3535_/C _3558_/B vdd gnd NAND2X1
XFILL_3__1915_ gnd vdd FILL
XFILL_2_CLKBUF1_insert30 gnd vdd FILL
XFILL_8__3589_ gnd vdd FILL
XFILL_8__2609_ gnd vdd FILL
XFILL_6__2673_ gnd vdd FILL
X_3464_ _3466_/B _3468_/B _3464_/C _3473_/B vdd gnd OAI21X1
XFILL_3__2895_ gnd vdd FILL
X_2415_ _2425_/B _2415_/B _2416_/C vdd gnd NOR2X1
XFILL_3__1846_ gnd vdd FILL
X_3395_ _3453_/B _3403_/A _3398_/B vdd gnd AND2X2
XFILL_9__3003_ gnd vdd FILL
XFILL_3__1777_ gnd vdd FILL
XFILL_1__2600_ gnd vdd FILL
XFILL_3__3516_ gnd vdd FILL
XFILL_0__1999_ gnd vdd FILL
X_2346_ _2346_/A _2346_/B _2350_/A vdd gnd NOR2X1
XFILL_1__3580_ gnd vdd FILL
XFILL_6__3225_ gnd vdd FILL
XFILL_0_BUFX2_insert23 gnd vdd FILL
XFILL_3__3447_ gnd vdd FILL
XFILL_4__2240_ gnd vdd FILL
XFILL_0_BUFX2_insert12 gnd vdd FILL
X_2277_ _2341_/A _3171_/B _2277_/C _2329_/C vdd gnd OAI21X1
XFILL_1__2531_ gnd vdd FILL
XFILL_0_BUFX2_insert56 gnd vdd FILL
XFILL_1__2462_ gnd vdd FILL
XFILL_0_BUFX2_insert45 gnd vdd FILL
XFILL_6__3156_ gnd vdd FILL
XFILL_3__3378_ gnd vdd FILL
XFILL_4__2171_ gnd vdd FILL
XFILL_6__3087_ gnd vdd FILL
XFILL_0_BUFX2_insert78 gnd vdd FILL
XFILL_6__2107_ gnd vdd FILL
XFILL_0_BUFX2_insert67 gnd vdd FILL
XFILL_0_BUFX2_insert89 gnd vdd FILL
XFILL_7__2920_ gnd vdd FILL
XFILL_6__2038_ gnd vdd FILL
XFILL_1__2393_ gnd vdd FILL
XFILL_3__2329_ gnd vdd FILL
XFILL_7__2851_ gnd vdd FILL
XFILL_1__3014_ gnd vdd FILL
XFILL_7__2782_ gnd vdd FILL
XFILL_7__1802_ gnd vdd FILL
XFILL_7__1733_ gnd vdd FILL
XFILL_4__1955_ gnd vdd FILL
XFILL_9__2649_ gnd vdd FILL
XFILL_7__3403_ gnd vdd FILL
XFILL_4__1886_ gnd vdd FILL
XFILL_4__3556_ gnd vdd FILL
XFILL_2__2640_ gnd vdd FILL
XFILL_4__2507_ gnd vdd FILL
XFILL_2__2571_ gnd vdd FILL
XFILL_4__3487_ gnd vdd FILL
XFILL_7__2216_ gnd vdd FILL
XFILL_5__2280_ gnd vdd FILL
XFILL_7__3196_ gnd vdd FILL
XFILL_1__2729_ gnd vdd FILL
XFILL_7__2147_ gnd vdd FILL
XFILL_4__2438_ gnd vdd FILL
XFILL_4__2369_ gnd vdd FILL
XFILL_7__2078_ gnd vdd FILL
XFILL_8__2960_ gnd vdd FILL
XFILL_2__3123_ gnd vdd FILL
XFILL_8__2891_ gnd vdd FILL
XFILL_8__1911_ gnd vdd FILL
XFILL_2__3054_ gnd vdd FILL
XFILL_8__1842_ gnd vdd FILL
XFILL_2__2005_ gnd vdd FILL
XFILL_8__3512_ gnd vdd FILL
XFILL_8__1773_ gnd vdd FILL
XFILL_5__1995_ gnd vdd FILL
XFILL_8__3443_ gnd vdd FILL
XFILL_2__2907_ gnd vdd FILL
XFILL_8__3374_ gnd vdd FILL
XFILL_3__1700_ gnd vdd FILL
XFILL_0__2971_ gnd vdd FILL
XFILL_8__2325_ gnd vdd FILL
XFILL_5__3596_ gnd vdd FILL
XFILL184350x7950 gnd vdd FILL
XFILL_0__1922_ gnd vdd FILL
XFILL_3__2680_ gnd vdd FILL
XFILL_5__2616_ gnd vdd FILL
XFILL_2__2838_ gnd vdd FILL
X_2200_ _3259_/Q _3312_/Q _2203_/A vdd gnd AND2X2
XFILL_5__2547_ gnd vdd FILL
XFILL_8__2256_ gnd vdd FILL
X_3180_ _3180_/A _3181_/B vdd gnd INVX1
XFILL_0__1853_ gnd vdd FILL
XFILL_2__2769_ gnd vdd FILL
XFILL_8__2187_ gnd vdd FILL
XFILL_5__2478_ gnd vdd FILL
X_2131_ _2602_/A _3166_/D _2717_/B vdd gnd NAND2X1
XFILL_0__1784_ gnd vdd FILL
XFILL_0__3523_ gnd vdd FILL
XFILL_6__3010_ gnd vdd FILL
X_2062_ _3282_/Q _2814_/A _2075_/B vdd gnd NOR2X1
XFILL_7_BUFX2_insert40 gnd vdd FILL
XFILL_7_BUFX2_insert51 gnd vdd FILL
XFILL_7_BUFX2_insert62 gnd vdd FILL
XFILL_7_BUFX2_insert73 gnd vdd FILL
XFILL_3__3232_ gnd vdd FILL
XFILL_0__3454_ gnd vdd FILL
XFILL_7_BUFX2_insert95 gnd vdd FILL
XFILL_7_BUFX2_insert84 gnd vdd FILL
XFILL_3__3163_ gnd vdd FILL
XFILL_0__3385_ gnd vdd FILL
XFILL_3__2114_ gnd vdd FILL
XFILL_0__2405_ gnd vdd FILL
XFILL_3__3094_ gnd vdd FILL
X_2964_ _2969_/A _2965_/B vdd gnd INVX1
XFILL_0__2336_ gnd vdd FILL
XFILL_0__2267_ gnd vdd FILL
XFILL_3__2045_ gnd vdd FILL
X_1915_ _1985_/A _3570_/Q _1915_/C _1916_/C vdd gnd AOI21X1
X_2895_ _2895_/A _2901_/A _2897_/B vdd gnd NOR2X1
X_1846_ _2058_/B _1846_/B _3158_/B vdd gnd NAND2X1
XFILL_0__2198_ gnd vdd FILL
X_1777_ _1810_/C _1777_/B _1777_/C _1778_/B vdd gnd NAND3X1
XFILL_6__2725_ gnd vdd FILL
X_3516_ _3518_/A _3516_/B _3516_/C _3535_/B vdd gnd OAI21X1
XFILL_3__2947_ gnd vdd FILL
XFILL_4__1740_ gnd vdd FILL
XFILL_6__2656_ gnd vdd FILL
XFILL_3__2878_ gnd vdd FILL
XFILL_1__1962_ gnd vdd FILL
XFILL_4__3410_ gnd vdd FILL
X_3447_ _3468_/S _3447_/B _3448_/B vdd gnd NOR2X1
XFILL_9__2296_ gnd vdd FILL
XFILL_3__1829_ gnd vdd FILL
XFILL_6__2587_ gnd vdd FILL
XFILL_1__1893_ gnd vdd FILL
X_3378_ _3468_/S _3453_/B vdd gnd INVX2
XFILL_1__3563_ gnd vdd FILL
XFILL_7__3050_ gnd vdd FILL
X_2329_ _2329_/A _2329_/B _2329_/C _2334_/A vdd gnd NAND3X1
XFILL_7__2001_ gnd vdd FILL
XFILL_6__3208_ gnd vdd FILL
XFILL_1__2514_ gnd vdd FILL
XFILL_1__3494_ gnd vdd FILL
XFILL_6__3139_ gnd vdd FILL
XFILL_4__2223_ gnd vdd FILL
XFILL_4__2154_ gnd vdd FILL
XFILL_1__2445_ gnd vdd FILL
XFILL_1__2376_ gnd vdd FILL
XFILL_7__2903_ gnd vdd FILL
XFILL_4__2085_ gnd vdd FILL
XFILL_7__2834_ gnd vdd FILL
XFILL_7__2765_ gnd vdd FILL
XFILL_4__2987_ gnd vdd FILL
XFILL_5__1780_ gnd vdd FILL
XFILL_7__2696_ gnd vdd FILL
XFILL_7__1716_ gnd vdd FILL
XFILL_4__1938_ gnd vdd FILL
XFILL_5__3450_ gnd vdd FILL
XFILL_4__1869_ gnd vdd FILL
XFILL_5__2401_ gnd vdd FILL
XFILL_8__3090_ gnd vdd FILL
XFILL_5__3381_ gnd vdd FILL
XFILL_2__2623_ gnd vdd FILL
XFILL_8__2110_ gnd vdd FILL
XFILL_8__2041_ gnd vdd FILL
XFILL_4__3539_ gnd vdd FILL
XFILL_5__2332_ gnd vdd FILL
XFILL_5__2263_ gnd vdd FILL
XFILL_2__2554_ gnd vdd FILL
XFILL_2__2485_ gnd vdd FILL
XFILL_7__3179_ gnd vdd FILL
XFILL_5__2194_ gnd vdd FILL
XFILL_8__2943_ gnd vdd FILL
XFILL_0_BUFX2_insert4 gnd vdd FILL
XFILL_2__3106_ gnd vdd FILL
XFILL_0__3170_ gnd vdd FILL
XFILL_8__2874_ gnd vdd FILL
XFILL_0__2121_ gnd vdd FILL
XFILL_2__3037_ gnd vdd FILL
XFILL_8__1825_ gnd vdd FILL
X_1700_ _2948_/A _3293_/D vdd gnd INVX1
XFILL_0__2052_ gnd vdd FILL
XFILL_8__1756_ gnd vdd FILL
X_2680_ _3356_/Q _2702_/B _2993_/B _2681_/C vdd gnd NAND3X1
XFILL_5__1978_ gnd vdd FILL
XFILL_3__2801_ gnd vdd FILL
XFILL_6__3490_ gnd vdd FILL
XFILL_8__3426_ gnd vdd FILL
XFILL_6__2510_ gnd vdd FILL
X_3301_ _3301_/D _3346_/CLK _3301_/Q vdd gnd DFFPOSX1
XFILL_3__2732_ gnd vdd FILL
XFILL_6__2441_ gnd vdd FILL
XFILL_0__2954_ gnd vdd FILL
XFILL_3__2663_ gnd vdd FILL
XFILL_6__2372_ gnd vdd FILL
XFILL_0__2885_ gnd vdd FILL
XFILL_8__2308_ gnd vdd FILL
XFILL_5__3579_ gnd vdd FILL
X_3232_ _3232_/A _3232_/B _3232_/C _3363_/D vdd gnd OAI21X1
XFILL_0__1905_ gnd vdd FILL
XFILL_0__1836_ gnd vdd FILL
XFILL_8__2239_ gnd vdd FILL
XFILL_3__2594_ gnd vdd FILL
X_3163_ _3163_/A _3194_/A _3164_/A vdd gnd NOR2X1
X_2114_ _3282_/Q _2886_/A vdd gnd INVX1
X_3094_ _3129_/A _3108_/B _3094_/C _3323_/D vdd gnd OAI21X1
XFILL_0__1767_ gnd vdd FILL
X_2045_ _2897_/C _2932_/B _2252_/B _2318_/B vdd gnd NAND3X1
XFILL_0__3506_ gnd vdd FILL
XFILL_3__3215_ gnd vdd FILL
XFILL_0__1698_ gnd vdd FILL
XFILL_0__3437_ gnd vdd FILL
XFILL_1__2230_ gnd vdd FILL
XFILL_1__2161_ gnd vdd FILL
XFILL_3__3146_ gnd vdd FILL
XFILL_3__3077_ gnd vdd FILL
XFILL_0__3368_ gnd vdd FILL
XFILL_4__2910_ gnd vdd FILL
X_2947_ reset _2957_/C _3302_/Q _2948_/C vdd gnd OAI21X1
XFILL_3__2028_ gnd vdd FILL
XFILL_0__2319_ gnd vdd FILL
XFILL_1__2092_ gnd vdd FILL
XFILL_9__1796_ gnd vdd FILL
XFILL_4__2841_ gnd vdd FILL
X_2878_ _3007_/A _2878_/B _2878_/C _3279_/D vdd gnd OAI21X1
XFILL_3_BUFX2_insert8 gnd vdd FILL
XFILL_7__2550_ gnd vdd FILL
X_1829_ _2668_/B _3189_/C _3079_/A _1831_/D _3403_/A vdd gnd OAI22X1
XFILL_6__2708_ gnd vdd FILL
XFILL_4__2772_ gnd vdd FILL
XFILL_3_BUFX2_insert82 gnd vdd FILL
XFILL_3_BUFX2_insert60 gnd vdd FILL
XFILL_1__2994_ gnd vdd FILL
XFILL_7__2481_ gnd vdd FILL
XFILL_4__1723_ gnd vdd FILL
XFILL_3_BUFX2_insert71 gnd vdd FILL
XFILL_3_BUFX2_insert93 gnd vdd FILL
XFILL_1__1945_ gnd vdd FILL
XFILL_6__2639_ gnd vdd FILL
XFILL_1__1876_ gnd vdd FILL
XFILL_7__3102_ gnd vdd FILL
XFILL_7__3033_ gnd vdd FILL
XFILL_1__3546_ gnd vdd FILL
XFILL_1__3477_ gnd vdd FILL
XFILL_2__2270_ gnd vdd FILL
XFILL_4__2206_ gnd vdd FILL
XFILL_1__2428_ gnd vdd FILL
XFILL_4__3186_ gnd vdd FILL
XFILL_4__2137_ gnd vdd FILL
XFILL_1__2359_ gnd vdd FILL
XFILL_5__2950_ gnd vdd FILL
XFILL_4__2068_ gnd vdd FILL
XFILL_5__1901_ gnd vdd FILL
XFILL_7__2817_ gnd vdd FILL
XFILL_5__2881_ gnd vdd FILL
XFILL_8__2590_ gnd vdd FILL
XFILL_5__1832_ gnd vdd FILL
XFILL_7__2748_ gnd vdd FILL
XFILL_5__1763_ gnd vdd FILL
XFILL_5__3502_ gnd vdd FILL
XFILL_2__1985_ gnd vdd FILL
XFILL_7__2679_ gnd vdd FILL
XFILL_5__1694_ gnd vdd FILL
XFILL_8__3211_ gnd vdd FILL
XFILL_8__3142_ gnd vdd FILL
XFILL_5__3433_ gnd vdd FILL
XFILL_5__3364_ gnd vdd FILL
XFILL_5__2315_ gnd vdd FILL
XFILL_8__3073_ gnd vdd FILL
XFILL_2__3586_ gnd vdd FILL
XFILL_2__2606_ gnd vdd FILL
XFILL_0__2670_ gnd vdd FILL
XFILL_8__2024_ gnd vdd FILL
XFILL_2__2537_ gnd vdd FILL
XFILL_5__2246_ gnd vdd FILL
XFILL_3__3000_ gnd vdd FILL
XFILL_5__2177_ gnd vdd FILL
XFILL_2__2468_ gnd vdd FILL
XFILL_2__2399_ gnd vdd FILL
XFILL_0__3222_ gnd vdd FILL
XFILL_8__2926_ gnd vdd FILL
XFILL_6__2990_ gnd vdd FILL
XFILL_6__1941_ gnd vdd FILL
XFILL_8__2857_ gnd vdd FILL
X_2801_ _2888_/B _2801_/B _2864_/C vdd gnd NOR2X1
XFILL_7_CLKBUF1_insert30 gnd vdd FILL
XFILL_0__3153_ gnd vdd FILL
XFILL_0__2104_ gnd vdd FILL
XFILL_6__1872_ gnd vdd FILL
XFILL_0__3084_ gnd vdd FILL
X_2732_ _2732_/A _2732_/B _2732_/C _2741_/A vdd gnd NAND3X1
XFILL_8__1808_ gnd vdd FILL
XFILL_0__2035_ gnd vdd FILL
XFILL_8__2788_ gnd vdd FILL
XFILL_6__3542_ gnd vdd FILL
XFILL_8__1739_ gnd vdd FILL
X_2663_ _3576_/Q _2670_/B _2663_/C _2686_/B vdd gnd AOI21X1
X_2594_ _2594_/A _2594_/B _2781_/A _2770_/B vdd gnd NOR3X1
XFILL_6__3473_ gnd vdd FILL
XFILL_8__3409_ gnd vdd FILL
XFILL_3__2715_ gnd vdd FILL
XFILL_6__2424_ gnd vdd FILL
XFILL_1__1730_ gnd vdd FILL
XFILL_0__2937_ gnd vdd FILL
XFILL_6__2355_ gnd vdd FILL
X_3215_ _3215_/A _3215_/B _3215_/C _3355_/D vdd gnd OAI21X1
XFILL_3__2646_ gnd vdd FILL
XFILL_0__2868_ gnd vdd FILL
XFILL_3__2577_ gnd vdd FILL
XFILL_1__3400_ gnd vdd FILL
XFILL_0__2799_ gnd vdd FILL
XFILL_0__1819_ gnd vdd FILL
XFILL_6__2286_ gnd vdd FILL
X_3146_ _3146_/A _3146_/B _3179_/C vdd gnd NOR2X1
X_3077_ _3083_/B _3083_/A _3077_/C _3078_/C vdd gnd AOI21X1
X_2028_ _2261_/B _2811_/A _2311_/A vdd gnd NOR2X1
XFILL_4__3040_ gnd vdd FILL
XFILL_3__3129_ gnd vdd FILL
XFILL_1__2213_ gnd vdd FILL
XFILL_7__1981_ gnd vdd FILL
XFILL_1__3193_ gnd vdd FILL
XFILL_1__2144_ gnd vdd FILL
XBUFX2_insert14 _1907_/Y _2771_/A vdd gnd BUFX2
XFILL_1__2075_ gnd vdd FILL
XFILL_7__2602_ gnd vdd FILL
XBUFX2_insert25 _2580_/Y _3363_/R vdd gnd BUFX2
XBUFX2_insert47 _1716_/Y _3157_/A vdd gnd BUFX2
XBUFX2_insert58 _3374_/Y _3560_/A vdd gnd BUFX2
XFILL_4__2824_ gnd vdd FILL
XFILL_7__3582_ gnd vdd FILL
XBUFX2_insert69 _1765_/Y _2966_/A vdd gnd BUFX2
XFILL_7__2533_ gnd vdd FILL
XFILL_7__2464_ gnd vdd FILL
XFILL_4__2755_ gnd vdd FILL
XFILL_1__2977_ gnd vdd FILL
XFILL_2__1770_ gnd vdd FILL
XFILL_4__1706_ gnd vdd FILL
XFILL_4__2686_ gnd vdd FILL
XFILL_1__1928_ gnd vdd FILL
XFILL_7__2395_ gnd vdd FILL
XFILL_8_BUFX2_insert17 gnd vdd FILL
XFILL_8_BUFX2_insert39 gnd vdd FILL
XFILL_1__1859_ gnd vdd FILL
XFILL_2__3440_ gnd vdd FILL
XFILL_2__3371_ gnd vdd FILL
XFILL_5__2100_ gnd vdd FILL
XFILL_5__3080_ gnd vdd FILL
XFILL_1__3529_ gnd vdd FILL
XFILL_7__3016_ gnd vdd FILL
XFILL_2__2322_ gnd vdd FILL
XFILL_5__2031_ gnd vdd FILL
XFILL_2__2253_ gnd vdd FILL
XFILL_4__3169_ gnd vdd FILL
XFILL_2__2184_ gnd vdd FILL
XFILL_8__2711_ gnd vdd FILL
XFILL_5__2933_ gnd vdd FILL
XFILL_8__2642_ gnd vdd FILL
XFILL_5__2864_ gnd vdd FILL
XFILL_8__2573_ gnd vdd FILL
XFILL_5__1815_ gnd vdd FILL
XFILL_5__2795_ gnd vdd FILL
XFILL_5__1746_ gnd vdd FILL
XFILL_2__1968_ gnd vdd FILL
XFILL_3__3480_ gnd vdd FILL
XFILL_5__3416_ gnd vdd FILL
XFILL_2__1899_ gnd vdd FILL
XFILL_3__2500_ gnd vdd FILL
XFILL_8__3125_ gnd vdd FILL
XFILL_0__2722_ gnd vdd FILL
XFILL_3__2431_ gnd vdd FILL
XFILL_8__3056_ gnd vdd FILL
X_3000_ _3571_/Q _3369_/Y _3260_/Q _3002_/B vdd gnd MUX2X1
XFILL_6__2140_ gnd vdd FILL
XFILL_0__2653_ gnd vdd FILL
XFILL_3__2362_ gnd vdd FILL
XFILL_6__2071_ gnd vdd FILL
XFILL_8__2007_ gnd vdd FILL
XFILL_0__2584_ gnd vdd FILL
XFILL_5__2229_ gnd vdd FILL
XFILL_3__2293_ gnd vdd FILL
XFILL_8__2909_ gnd vdd FILL
XFILL_6__2973_ gnd vdd FILL
XFILL_0__3205_ gnd vdd FILL
XFILL_0__3136_ gnd vdd FILL
XFILL_6__1924_ gnd vdd FILL
XFILL_0__3067_ gnd vdd FILL
XFILL_6__1855_ gnd vdd FILL
X_2715_ _2715_/A _2746_/B _2715_/C _2718_/C vdd gnd OAI21X1
XFILL_1__2900_ gnd vdd FILL
XFILL_0__2018_ gnd vdd FILL
X_2646_ _2646_/A _2671_/B _2656_/B _2653_/B vdd gnd OAI21X1
XFILL_6__1786_ gnd vdd FILL
XFILL_6__3525_ gnd vdd FILL
XFILL_1__2831_ gnd vdd FILL
XFILL_6__3456_ gnd vdd FILL
X_2577_ _3035_/B _2960_/B _3524_/A vdd gnd NOR2X1
XFILL_4__2540_ gnd vdd FILL
XFILL_4__2471_ gnd vdd FILL
XFILL_9__3165_ gnd vdd FILL
XFILL_1__2762_ gnd vdd FILL
XFILL_6__2407_ gnd vdd FILL
XFILL_7__2180_ gnd vdd FILL
XFILL_6__3387_ gnd vdd FILL
XFILL_1__2693_ gnd vdd FILL
XFILL_1__1713_ gnd vdd FILL
XFILL_3__2629_ gnd vdd FILL
XFILL_6__2338_ gnd vdd FILL
XFILL_6__2269_ gnd vdd FILL
X_3129_ _3129_/A _3143_/B _3129_/C _3340_/D vdd gnd OAI21X1
XFILL_4__3023_ gnd vdd FILL
XFILL_7__1964_ gnd vdd FILL
XFILL_1__3176_ gnd vdd FILL
XFILL_1__2127_ gnd vdd FILL
XFILL_7__1895_ gnd vdd FILL
XFILL_2__2940_ gnd vdd FILL
XFILL_1__2058_ gnd vdd FILL
XFILL_7__3565_ gnd vdd FILL
XFILL_5__2580_ gnd vdd FILL
XFILL_4__2807_ gnd vdd FILL
XFILL_2__2871_ gnd vdd FILL
XFILL_7__2516_ gnd vdd FILL
XFILL_7__3496_ gnd vdd FILL
XFILL_4__2738_ gnd vdd FILL
XFILL_2__1822_ gnd vdd FILL
XFILL_7__2447_ gnd vdd FILL
XFILL_2__1753_ gnd vdd FILL
XFILL_7__2378_ gnd vdd FILL
XFILL_4__2669_ gnd vdd FILL
XFILL_5__3201_ gnd vdd FILL
XFILL_2__3423_ gnd vdd FILL
XFILL_5__3132_ gnd vdd FILL
XFILL_5__3063_ gnd vdd FILL
XFILL_5__2014_ gnd vdd FILL
XFILL_2__2305_ gnd vdd FILL
XFILL181650x117150 gnd vdd FILL
XFILL181950x109350 gnd vdd FILL
XFILL_2__2236_ gnd vdd FILL
XFILL_2__2167_ gnd vdd FILL
XFILL_4_BUFX2_insert15 gnd vdd FILL
XFILL_4_BUFX2_insert26 gnd vdd FILL
XFILL_4_BUFX2_insert48 gnd vdd FILL
XFILL_3__2980_ gnd vdd FILL
XFILL_2__2098_ gnd vdd FILL
XFILL_5__2916_ gnd vdd FILL
XFILL_4_BUFX2_insert59 gnd vdd FILL
XFILL_3__1931_ gnd vdd FILL
XFILL_8__2625_ gnd vdd FILL
X_3480_ _3482_/A _3480_/B _3480_/C _3526_/B vdd gnd OAI21X1
XFILL_5__2847_ gnd vdd FILL
X_2500_ _3211_/B _3590_/A vdd gnd INVX1
XFILL_3__1862_ gnd vdd FILL
XFILL_5__2778_ gnd vdd FILL
XFILL_8__2556_ gnd vdd FILL
X_2431_ _2431_/A _2431_/B _2519_/C vdd gnd OR2X2
XFILL_3__3601_ gnd vdd FILL
XFILL_8__2487_ gnd vdd FILL
XFILL_5__1729_ gnd vdd FILL
XFILL_3__1793_ gnd vdd FILL
X_2362_ _3272_/Q _2861_/A vdd gnd INVX1
XFILL_3__3532_ gnd vdd FILL
X_2293_ _2293_/A _2433_/A _2293_/C _2342_/C vdd gnd OAI21X1
XFILL_8__3108_ gnd vdd FILL
XFILL_3__3463_ gnd vdd FILL
XFILL_0__2705_ gnd vdd FILL
XFILL_6__3172_ gnd vdd FILL
XFILL_3__3394_ gnd vdd FILL
XFILL_3__2414_ gnd vdd FILL
XFILL_6__2123_ gnd vdd FILL
XFILL_8__3039_ gnd vdd FILL
XFILL_3__2345_ gnd vdd FILL
XFILL_0__2636_ gnd vdd FILL
XFILL_6__2054_ gnd vdd FILL
XFILL_0__2567_ gnd vdd FILL
XFILL_3__2276_ gnd vdd FILL
XFILL_0__2498_ gnd vdd FILL
XFILL_1__3030_ gnd vdd FILL
XFILL_6__2956_ gnd vdd FILL
XFILL_8_BUFX2_insert3 gnd vdd FILL
XFILL_0__3119_ gnd vdd FILL
XFILL_6__2887_ gnd vdd FILL
XFILL_6__1907_ gnd vdd FILL
XFILL_4__1971_ gnd vdd FILL
XFILL_6__1838_ gnd vdd FILL
XFILL_7__2301_ gnd vdd FILL
XFILL_6__1769_ gnd vdd FILL
X_2629_ _2778_/A _2629_/B _2629_/C _3241_/D vdd gnd OAI21X1
XFILL_6__3508_ gnd vdd FILL
XFILL_1__2814_ gnd vdd FILL
XFILL_4__2523_ gnd vdd FILL
XFILL_6__3439_ gnd vdd FILL
XFILL_1__2745_ gnd vdd FILL
XFILL_7__2232_ gnd vdd FILL
XFILL_7__2163_ gnd vdd FILL
XFILL_4__2454_ gnd vdd FILL
XFILL_4__2385_ gnd vdd FILL
XFILL_1__2676_ gnd vdd FILL
XFILL_7__2094_ gnd vdd FILL
XFILL_4__3006_ gnd vdd FILL
XFILL_2__3070_ gnd vdd FILL
XFILL_2__2021_ gnd vdd FILL
XFILL_7__2996_ gnd vdd FILL
XFILL_1__3228_ gnd vdd FILL
XFILL_7__1947_ gnd vdd FILL
XFILL_1__3159_ gnd vdd FILL
XFILL_7__1878_ gnd vdd FILL
XFILL_5__2701_ gnd vdd FILL
XFILL_8__2410_ gnd vdd FILL
XFILL_2__2923_ gnd vdd FILL
XFILL_8__3390_ gnd vdd FILL
XFILL_5__2632_ gnd vdd FILL
XFILL_7__3548_ gnd vdd FILL
XFILL_2__2854_ gnd vdd FILL
XFILL_8__2341_ gnd vdd FILL
XFILL_7__3479_ gnd vdd FILL
XFILL_8__2272_ gnd vdd FILL
XFILL_2__1805_ gnd vdd FILL
XFILL_5__2563_ gnd vdd FILL
XFILL_2__2785_ gnd vdd FILL
XFILL_5__2494_ gnd vdd FILL
XFILL_2__1736_ gnd vdd FILL
XFILL_0__3470_ gnd vdd FILL
XFILL_5__3115_ gnd vdd FILL
XFILL_2__3406_ gnd vdd FILL
XFILL_0__2421_ gnd vdd FILL
XFILL_3__2130_ gnd vdd FILL
XFILL_5__3046_ gnd vdd FILL
XFILL183150x105450 gnd vdd FILL
XFILL_0__2352_ gnd vdd FILL
X_2980_ _2980_/A _3148_/B _2984_/C vdd gnd NAND2X1
XFILL_3__2061_ gnd vdd FILL
XFILL_4_CLKBUF1_insert38 gnd vdd FILL
X_1931_ _1931_/A _1931_/B _1931_/C _2474_/A vdd gnd NAND3X1
XFILL_0__2283_ gnd vdd FILL
XFILL_2__2219_ gnd vdd FILL
XFILL_8__1987_ gnd vdd FILL
XFILL_2__3199_ gnd vdd FILL
X_1862_ _2906_/B _1862_/B _1873_/A _1875_/A vdd gnd NAND3X1
XFILL_6__2810_ gnd vdd FILL
X_3601_ _3601_/A DO[6] vdd gnd BUFX2
XFILL_6__2741_ gnd vdd FILL
XFILL_3__2963_ gnd vdd FILL
X_1793_ _3235_/Q _1793_/B _1891_/B vdd gnd NOR2X1
XFILL_6__2672_ gnd vdd FILL
XFILL_3__2894_ gnd vdd FILL
X_3532_ _3532_/A _3532_/B _3533_/A vdd gnd NAND2X1
XFILL_3__1914_ gnd vdd FILL
XFILL_8__3588_ gnd vdd FILL
XFILL_2_CLKBUF1_insert31 gnd vdd FILL
XFILL_8__2608_ gnd vdd FILL
X_3463_ _3484_/C _3464_/C vdd gnd INVX1
XFILL_3__1845_ gnd vdd FILL
XFILL_8__2539_ gnd vdd FILL
X_2414_ _2659_/B _2426_/B _2414_/C _2415_/B vdd gnd OAI21X1
X_3394_ _3521_/A _3565_/A _3399_/C vdd gnd NAND2X1
XFILL_3__1776_ gnd vdd FILL
XFILL_3__3515_ gnd vdd FILL
XFILL_0__1998_ gnd vdd FILL
X_2345_ _2345_/A _2345_/B _2346_/B vdd gnd NAND2X1
XFILL_6__3224_ gnd vdd FILL
XFILL_3__3446_ gnd vdd FILL
XFILL_0_BUFX2_insert24 gnd vdd FILL
X_2276_ _2276_/A _3147_/B _2341_/A _2277_/C vdd gnd OAI21X1
XFILL_1__2530_ gnd vdd FILL
XFILL_0_BUFX2_insert13 gnd vdd FILL
XFILL_0_BUFX2_insert57 gnd vdd FILL
XFILL_1__2461_ gnd vdd FILL
XFILL_0_BUFX2_insert46 gnd vdd FILL
XFILL_6__3155_ gnd vdd FILL
XFILL_3__3377_ gnd vdd FILL
XFILL_4__2170_ gnd vdd FILL
XFILL_0_BUFX2_insert79 gnd vdd FILL
XFILL_6__3086_ gnd vdd FILL
XFILL_0_BUFX2_insert68 gnd vdd FILL
XFILL_0__2619_ gnd vdd FILL
XFILL_6__2106_ gnd vdd FILL
XFILL_6__2037_ gnd vdd FILL
XFILL_3__2328_ gnd vdd FILL
XFILL_0__3599_ gnd vdd FILL
XFILL_1__2392_ gnd vdd FILL
XFILL_3__2259_ gnd vdd FILL
XFILL_7__2850_ gnd vdd FILL
XFILL_1__3013_ gnd vdd FILL
XFILL_7__2781_ gnd vdd FILL
XFILL_7__1801_ gnd vdd FILL
XFILL_6__2939_ gnd vdd FILL
XFILL_7__1732_ gnd vdd FILL
XFILL_4__1954_ gnd vdd FILL
XFILL_7__3402_ gnd vdd FILL
XFILL_4__1885_ gnd vdd FILL
XFILL_4__3555_ gnd vdd FILL
XFILL_4__3486_ gnd vdd FILL
XFILL_7__2215_ gnd vdd FILL
XFILL_4__2506_ gnd vdd FILL
XFILL_2__2570_ gnd vdd FILL
XFILL_7__3195_ gnd vdd FILL
XFILL_1__2728_ gnd vdd FILL
XFILL_4__2437_ gnd vdd FILL
XFILL_7__2146_ gnd vdd FILL
XFILL_1__2659_ gnd vdd FILL
XFILL_7__2077_ gnd vdd FILL
XFILL_4__2368_ gnd vdd FILL
XFILL_4__2299_ gnd vdd FILL
XFILL_2__3122_ gnd vdd FILL
XFILL_8__2890_ gnd vdd FILL
XFILL_8__1910_ gnd vdd FILL
XFILL_2__3053_ gnd vdd FILL
XFILL_8__1841_ gnd vdd FILL
XFILL_2__2004_ gnd vdd FILL
XFILL_8__3511_ gnd vdd FILL
XFILL_5__1994_ gnd vdd FILL
XFILL_7__2979_ gnd vdd FILL
XFILL_8__1772_ gnd vdd FILL
XFILL183750x35250 gnd vdd FILL
XFILL_8__3442_ gnd vdd FILL
XFILL_8__3373_ gnd vdd FILL
XFILL_2__2906_ gnd vdd FILL
XFILL_0__2970_ gnd vdd FILL
XFILL_0__1921_ gnd vdd FILL
XFILL_8__2324_ gnd vdd FILL
XFILL_5__3595_ gnd vdd FILL
XFILL_5__2615_ gnd vdd FILL
XFILL_2__2837_ gnd vdd FILL
XFILL_5__2546_ gnd vdd FILL
XFILL_8__2255_ gnd vdd FILL
XFILL_0__1852_ gnd vdd FILL
XFILL_2__2768_ gnd vdd FILL
XFILL_8__2186_ gnd vdd FILL
XFILL183150x117150 gnd vdd FILL
XFILL183450x109350 gnd vdd FILL
X_2130_ _2331_/A _2348_/B _2135_/A vdd gnd NAND2X1
XFILL_2__1719_ gnd vdd FILL
XFILL_0__1783_ gnd vdd FILL
XFILL_5__2477_ gnd vdd FILL
XFILL_0__3522_ gnd vdd FILL
X_2061_ _2786_/A _2176_/A _2115_/B _2318_/A vdd gnd NAND3X1
XFILL_3__3231_ gnd vdd FILL
XFILL_2__2699_ gnd vdd FILL
XFILL_0__3453_ gnd vdd FILL
XFILL_7_BUFX2_insert63 gnd vdd FILL
XFILL_7_BUFX2_insert74 gnd vdd FILL
XFILL_7_BUFX2_insert52 gnd vdd FILL
XFILL_7_BUFX2_insert41 gnd vdd FILL
XFILL_7_BUFX2_insert96 gnd vdd FILL
XFILL_7_BUFX2_insert85 gnd vdd FILL
XFILL_0__2404_ gnd vdd FILL
XFILL_3__3162_ gnd vdd FILL
XFILL_5__3029_ gnd vdd FILL
XFILL_3__3093_ gnd vdd FILL
XFILL_0__3384_ gnd vdd FILL
XFILL_3__2113_ gnd vdd FILL
XFILL_3__2044_ gnd vdd FILL
X_2963_ _3268_/Q _3023_/B _2969_/A vdd gnd NOR2X1
XFILL_0__2335_ gnd vdd FILL
XFILL_0__2266_ gnd vdd FILL
X_1914_ _3016_/A _1984_/B _2521_/C _1915_/C vdd gnd OAI21X1
X_2894_ _2894_/A _2931_/B _2901_/A vdd gnd NAND2X1
XFILL_0__2197_ gnd vdd FILL
XFILL_9__2502_ gnd vdd FILL
X_1845_ _1858_/B _1888_/B _2448_/B vdd gnd NAND2X1
XFILL_6__2724_ gnd vdd FILL
X_1776_ _1782_/B _3149_/C _1987_/A _1777_/B vdd gnd OAI21X1
X_3515_ _3515_/A _3516_/B vdd gnd INVX1
XFILL_3__2946_ gnd vdd FILL
XFILL_1__1961_ gnd vdd FILL
XFILL_6__2655_ gnd vdd FILL
XFILL_3__2877_ gnd vdd FILL
XFILL_6__2586_ gnd vdd FILL
X_3446_ _3451_/B _3447_/B vdd gnd INVX1
XFILL_1__1892_ gnd vdd FILL
XFILL_3__1828_ gnd vdd FILL
X_3377_ _3468_/S _3445_/A _3455_/C vdd gnd NAND2X1
XFILL_3__1759_ gnd vdd FILL
XFILL_1__3562_ gnd vdd FILL
X_2328_ _2328_/A _2328_/B _2337_/A vdd gnd NOR2X1
XFILL_7__2000_ gnd vdd FILL
XFILL_6__3207_ gnd vdd FILL
XFILL_1__2513_ gnd vdd FILL
XFILL_1__3493_ gnd vdd FILL
XFILL_6__3138_ gnd vdd FILL
XFILL_3__3429_ gnd vdd FILL
X_2259_ _2297_/B _2297_/A _2263_/C vdd gnd OR2X2
XFILL_4__2222_ gnd vdd FILL
XFILL_4__2153_ gnd vdd FILL
XFILL_1__2444_ gnd vdd FILL
XFILL_6__3069_ gnd vdd FILL
XFILL_1__2375_ gnd vdd FILL
XFILL_7__2902_ gnd vdd FILL
XFILL_4__2084_ gnd vdd FILL
XFILL_7__2833_ gnd vdd FILL
XFILL_7__2764_ gnd vdd FILL
XFILL_4__2986_ gnd vdd FILL
XFILL_7__2695_ gnd vdd FILL
XFILL_7__1715_ gnd vdd FILL
XFILL_4__1937_ gnd vdd FILL
XFILL_4__1868_ gnd vdd FILL
XFILL_5__3380_ gnd vdd FILL
XFILL_5__2400_ gnd vdd FILL
XFILL_5__2331_ gnd vdd FILL
XFILL_4__1799_ gnd vdd FILL
XFILL_2__2622_ gnd vdd FILL
XFILL_8__2040_ gnd vdd FILL
XFILL_4__3538_ gnd vdd FILL
XFILL_2__2553_ gnd vdd FILL
XFILL_4__3469_ gnd vdd FILL
XFILL_5__2262_ gnd vdd FILL
XFILL_7__3178_ gnd vdd FILL
XFILL_5__2193_ gnd vdd FILL
XFILL_2__2484_ gnd vdd FILL
XFILL_7__2129_ gnd vdd FILL
XFILL_8__2942_ gnd vdd FILL
XFILL_0_BUFX2_insert5 gnd vdd FILL
XFILL_2__3105_ gnd vdd FILL
XFILL_8__2873_ gnd vdd FILL
XFILL_0__2120_ gnd vdd FILL
XFILL_2__3036_ gnd vdd FILL
XFILL_8__1824_ gnd vdd FILL
XFILL_8__1755_ gnd vdd FILL
XFILL_0__2051_ gnd vdd FILL
XFILL_5__1977_ gnd vdd FILL
XFILL_3__2800_ gnd vdd FILL
XFILL_8__3425_ gnd vdd FILL
X_3300_ _3300_/D _3313_/CLK _3300_/Q vdd gnd DFFPOSX1
XFILL_3__2731_ gnd vdd FILL
XFILL_6__2440_ gnd vdd FILL
XFILL_0__2953_ gnd vdd FILL
XFILL_3__2662_ gnd vdd FILL
XFILL_0__2884_ gnd vdd FILL
XFILL_6__2371_ gnd vdd FILL
XFILL_8__2307_ gnd vdd FILL
X_3231_ _3586_/A _3232_/B _3232_/C vdd gnd NAND2X1
XFILL_0__1904_ gnd vdd FILL
XFILL_8__2238_ gnd vdd FILL
XFILL_5__2529_ gnd vdd FILL
XFILL_3__2593_ gnd vdd FILL
XFILL_0__1835_ gnd vdd FILL
X_3162_ _3162_/A _3173_/C vdd gnd INVX1
X_2113_ _2339_/B _2284_/A _2113_/C _2158_/B vdd gnd NAND3X1
X_3093_ _3111_/A _3107_/B _3323_/Q _3094_/C vdd gnd OAI21X1
XFILL_8__2169_ gnd vdd FILL
XFILL_0__3505_ gnd vdd FILL
XFILL_0__1766_ gnd vdd FILL
X_2044_ _2044_/A _2044_/B _2896_/C _2252_/B vdd gnd OAI21X1
XFILL_0__1697_ gnd vdd FILL
XFILL_3__3214_ gnd vdd FILL
XFILL_0__3436_ gnd vdd FILL
XFILL_3__3145_ gnd vdd FILL
XFILL_1__2160_ gnd vdd FILL
XFILL_0__3367_ gnd vdd FILL
XFILL_3__3076_ gnd vdd FILL
XFILL_0__2318_ gnd vdd FILL
XFILL_3__2027_ gnd vdd FILL
X_2946_ _2985_/A _2956_/B _2946_/C _3301_/D vdd gnd OAI21X1
XFILL_1__2091_ gnd vdd FILL
XFILL_0__2249_ gnd vdd FILL
X_2877_ _3279_/Q _3007_/A vdd gnd INVX1
XFILL_4__2840_ gnd vdd FILL
XFILL_3_BUFX2_insert9 gnd vdd FILL
X_1828_ _3245_/Q _2668_/B vdd gnd INVX2
XFILL_6__2707_ gnd vdd FILL
XFILL_4__2771_ gnd vdd FILL
XFILL_7__2480_ gnd vdd FILL
XFILL_3__2929_ gnd vdd FILL
XFILL_3_BUFX2_insert61 gnd vdd FILL
XFILL_3_BUFX2_insert50 gnd vdd FILL
X_1759_ _3277_/Q _3007_/B vdd gnd INVX1
XFILL_1__2993_ gnd vdd FILL
XFILL_3_BUFX2_insert83 gnd vdd FILL
XFILL_4__1722_ gnd vdd FILL
XFILL_3_BUFX2_insert72 gnd vdd FILL
XFILL_3_BUFX2_insert94 gnd vdd FILL
XFILL_6__2638_ gnd vdd FILL
XFILL_1__1944_ gnd vdd FILL
XFILL_1__1875_ gnd vdd FILL
X_3429_ _3431_/A _3432_/A _3500_/C vdd gnd NAND2X1
XFILL_6__2569_ gnd vdd FILL
XFILL_7__3101_ gnd vdd FILL
XFILL_7__3032_ gnd vdd FILL
XFILL_1__3545_ gnd vdd FILL
XFILL_1__3476_ gnd vdd FILL
XFILL_4__2205_ gnd vdd FILL
XFILL_1__2427_ gnd vdd FILL
XFILL_4__3185_ gnd vdd FILL
XFILL_4__2136_ gnd vdd FILL
XFILL_1__2358_ gnd vdd FILL
XFILL_4__2067_ gnd vdd FILL
XFILL_5__1900_ gnd vdd FILL
XFILL_1__2289_ gnd vdd FILL
XFILL_5__2880_ gnd vdd FILL
XFILL_7__2816_ gnd vdd FILL
XFILL_5__1831_ gnd vdd FILL
XFILL_7__2747_ gnd vdd FILL
XFILL_4__2969_ gnd vdd FILL
XFILL_5__1762_ gnd vdd FILL
XFILL_5__3501_ gnd vdd FILL
XFILL_2__1984_ gnd vdd FILL
XFILL_7__2678_ gnd vdd FILL
XFILL_8__3210_ gnd vdd FILL
XFILL_5__1693_ gnd vdd FILL
XFILL_8__3141_ gnd vdd FILL
XFILL_5__3432_ gnd vdd FILL
XFILL_8__3072_ gnd vdd FILL
XFILL_2__2605_ gnd vdd FILL
XFILL_5__2314_ gnd vdd FILL
XFILL_2__3585_ gnd vdd FILL
XFILL_8__2023_ gnd vdd FILL
XFILL_5__2245_ gnd vdd FILL
XFILL_2__2536_ gnd vdd FILL
XFILL_2__2467_ gnd vdd FILL
XFILL_5__2176_ gnd vdd FILL
XFILL_2__2398_ gnd vdd FILL
XFILL_0__3221_ gnd vdd FILL
XFILL_8__2925_ gnd vdd FILL
XFILL_6__1940_ gnd vdd FILL
XFILL_8__2856_ gnd vdd FILL
X_2800_ _3263_/Q _3009_/A vdd gnd INVX1
XFILL_0__3152_ gnd vdd FILL
XFILL_7_CLKBUF1_insert31 gnd vdd FILL
XFILL_6__1871_ gnd vdd FILL
XFILL_2__3019_ gnd vdd FILL
XFILL_0__3083_ gnd vdd FILL
XFILL_8__1807_ gnd vdd FILL
X_2731_ _2731_/A _2732_/A _2732_/B _2734_/D vdd gnd AOI21X1
XFILL_0__2103_ gnd vdd FILL
XFILL_0__2034_ gnd vdd FILL
XFILL_8__2787_ gnd vdd FILL
XFILL_6__3541_ gnd vdd FILL
XFILL_8__1738_ gnd vdd FILL
X_2662_ _2662_/A _2748_/B _2669_/C _2663_/C vdd gnd OAI21X1
X_2593_ _2756_/B _2751_/B vdd gnd INVX2
XFILL_6__3472_ gnd vdd FILL
XFILL_8__3408_ gnd vdd FILL
XFILL_3__2714_ gnd vdd FILL
XFILL_0__2936_ gnd vdd FILL
XFILL_6__2423_ gnd vdd FILL
XFILL_6__2354_ gnd vdd FILL
X_3214_ _3214_/A _3214_/B _3355_/Q _3215_/C vdd gnd OAI21X1
XFILL_3__2645_ gnd vdd FILL
XFILL_0__2867_ gnd vdd FILL
XFILL_3__2576_ gnd vdd FILL
XFILL_0__2798_ gnd vdd FILL
XFILL_6__2285_ gnd vdd FILL
XFILL_0__1818_ gnd vdd FILL
X_3145_ _3237_/Q _3145_/B _3181_/A _3146_/B vdd gnd OAI21X1
X_3076_ _3084_/B _3576_/Q _3083_/A vdd gnd XNOR2X1
XFILL_0__1749_ gnd vdd FILL
X_2027_ _2933_/B _2857_/A _2811_/A vdd gnd NAND2X1
XFILL_0__3419_ gnd vdd FILL
XFILL182250x74250 gnd vdd FILL
XFILL_1__2212_ gnd vdd FILL
XFILL_3__3128_ gnd vdd FILL
XFILL_7__1980_ gnd vdd FILL
XFILL_1__3192_ gnd vdd FILL
XFILL_3__3059_ gnd vdd FILL
XFILL_1__2143_ gnd vdd FILL
X_2929_ _2929_/A _2929_/B _2936_/C vdd gnd NOR2X1
XFILL_1__2074_ gnd vdd FILL
XBUFX2_insert15 _1907_/Y _2728_/A vdd gnd BUFX2
XBUFX2_insert26 _2580_/Y _3347_/R vdd gnd BUFX2
XBUFX2_insert48 _3307_/Q _2025_/A vdd gnd BUFX2
XFILL_7__2601_ gnd vdd FILL
XBUFX2_insert59 _3374_/Y _3552_/A vdd gnd BUFX2
XFILL_4__2823_ gnd vdd FILL
XFILL_7__3581_ gnd vdd FILL
XFILL_7__2532_ gnd vdd FILL
XFILL_1__2976_ gnd vdd FILL
XFILL_7__2463_ gnd vdd FILL
XFILL_4__2754_ gnd vdd FILL
XFILL_4__1705_ gnd vdd FILL
XFILL_4__2685_ gnd vdd FILL
XFILL_8_BUFX2_insert18 gnd vdd FILL
XFILL_1__1927_ gnd vdd FILL
XFILL_7__2394_ gnd vdd FILL
XFILL_1__1858_ gnd vdd FILL
XFILL_2__3370_ gnd vdd FILL
XFILL_1__1789_ gnd vdd FILL
XFILL_1__3528_ gnd vdd FILL
XFILL_7__3015_ gnd vdd FILL
XFILL_2__2321_ gnd vdd FILL
XFILL_5__2030_ gnd vdd FILL
XFILL_1__3459_ gnd vdd FILL
XFILL_2__2252_ gnd vdd FILL
XFILL_4__3168_ gnd vdd FILL
XFILL_2__2183_ gnd vdd FILL
XFILL_4__2119_ gnd vdd FILL
XFILL_4__3099_ gnd vdd FILL
XFILL_8__2710_ gnd vdd FILL
XFILL_5__2932_ gnd vdd FILL
XFILL_8__2641_ gnd vdd FILL
XFILL_5__2863_ gnd vdd FILL
XFILL_8__2572_ gnd vdd FILL
XFILL_5__1814_ gnd vdd FILL
XFILL_5__2794_ gnd vdd FILL
XFILL_5__1745_ gnd vdd FILL
XFILL_2__1967_ gnd vdd FILL
XFILL_5__3415_ gnd vdd FILL
XFILL_2__1898_ gnd vdd FILL
XFILL_0__2721_ gnd vdd FILL
XFILL_8__3124_ gnd vdd FILL
XFILL_3__2430_ gnd vdd FILL
XFILL_3__2361_ gnd vdd FILL
XFILL_8__3055_ gnd vdd FILL
XFILL_0__2652_ gnd vdd FILL
XFILL_8__2006_ gnd vdd FILL
XFILL_6__2070_ gnd vdd FILL
XFILL_0__2583_ gnd vdd FILL
XFILL_2__3499_ gnd vdd FILL
XFILL_5__2228_ gnd vdd FILL
XFILL_2__2519_ gnd vdd FILL
XFILL_3__2292_ gnd vdd FILL
XFILL_5__2159_ gnd vdd FILL
XFILL_8__2908_ gnd vdd FILL
XFILL_6__2972_ gnd vdd FILL
XFILL_0__3204_ gnd vdd FILL
XFILL_0__3135_ gnd vdd FILL
XFILL_6__1923_ gnd vdd FILL
XFILL_8__2839_ gnd vdd FILL
XFILL_0__3066_ gnd vdd FILL
XFILL_6__1854_ gnd vdd FILL
X_2714_ _3221_/A _3147_/C _2889_/C _2718_/A vdd gnd NOR3X1
XFILL_0__2017_ gnd vdd FILL
XFILL_6__1785_ gnd vdd FILL
X_2645_ _3574_/Q _2670_/B _2645_/C _2656_/B vdd gnd AOI21X1
XFILL184350x171750 gnd vdd FILL
XFILL184650x163950 gnd vdd FILL
XFILL_1__2830_ gnd vdd FILL
XFILL_6__3524_ gnd vdd FILL
XFILL_6__3455_ gnd vdd FILL
X_2576_ _3278_/Q _3035_/B vdd gnd INVX1
XFILL_4__2470_ gnd vdd FILL
XFILL_1__2761_ gnd vdd FILL
XFILL_6__2406_ gnd vdd FILL
XFILL_0__2919_ gnd vdd FILL
XFILL_6__3386_ gnd vdd FILL
XFILL_1__1712_ gnd vdd FILL
XFILL_1__2692_ gnd vdd FILL
XFILL_3__2628_ gnd vdd FILL
XFILL_6__2337_ gnd vdd FILL
XFILL_9__2046_ gnd vdd FILL
X_3128_ _3340_/Q _3143_/B _3129_/C vdd gnd NAND2X1
XFILL_6__2268_ gnd vdd FILL
XFILL_3__2559_ gnd vdd FILL
X_3059_ _3059_/A _3059_/B _3088_/S _3060_/C vdd gnd OAI21X1
XFILL_4__3022_ gnd vdd FILL
XFILL_6__2199_ gnd vdd FILL
XFILL_7__1963_ gnd vdd FILL
XFILL_1__3175_ gnd vdd FILL
XFILL_1__2126_ gnd vdd FILL
XFILL_7__1894_ gnd vdd FILL
XFILL_1__2057_ gnd vdd FILL
XFILL_2__2870_ gnd vdd FILL
XFILL_7__3564_ gnd vdd FILL
XFILL_4__2806_ gnd vdd FILL
XFILL_7__2515_ gnd vdd FILL
XFILL_7__3495_ gnd vdd FILL
XFILL_2__1821_ gnd vdd FILL
XFILL_4__2737_ gnd vdd FILL
XFILL_1__2959_ gnd vdd FILL
XFILL_7__2446_ gnd vdd FILL
XFILL_2__1752_ gnd vdd FILL
XFILL_7__2377_ gnd vdd FILL
XFILL_4__2668_ gnd vdd FILL
XFILL_5__3200_ gnd vdd FILL
XFILL_2__3422_ gnd vdd FILL
XFILL_4__2599_ gnd vdd FILL
XFILL_5__3131_ gnd vdd FILL
XFILL_5__3062_ gnd vdd FILL
XFILL_5_BUFX2_insert0 gnd vdd FILL
XFILL_5__2013_ gnd vdd FILL
XFILL_2__2304_ gnd vdd FILL
XFILL_2__2235_ gnd vdd FILL
XFILL_2__2166_ gnd vdd FILL
XFILL_5__2915_ gnd vdd FILL
XFILL_2__2097_ gnd vdd FILL
XFILL_4_BUFX2_insert27 gnd vdd FILL
XFILL_4_BUFX2_insert16 gnd vdd FILL
XFILL_3__1930_ gnd vdd FILL
XFILL_4_BUFX2_insert49 gnd vdd FILL
XFILL_8__2624_ gnd vdd FILL
XFILL_5__2846_ gnd vdd FILL
XFILL_8__2555_ gnd vdd FILL
XFILL_3__1861_ gnd vdd FILL
X_2430_ _2430_/A _2430_/B _3188_/A _2431_/B vdd gnd OAI21X1
XFILL_5__2777_ gnd vdd FILL
XFILL_2__2999_ gnd vdd FILL
XFILL_3__3600_ gnd vdd FILL
XFILL_3__1792_ gnd vdd FILL
XFILL_8__2486_ gnd vdd FILL
XFILL_5__1728_ gnd vdd FILL
X_2361_ _2841_/A _2579_/B _2361_/C _3468_/A vdd gnd OAI21X1
XFILL_3__3531_ gnd vdd FILL
X_2292_ _3182_/B _2292_/B _2293_/A _2293_/C vdd gnd OAI21X1
XFILL_8__3107_ gnd vdd FILL
XFILL_3__3462_ gnd vdd FILL
XFILL_6__3171_ gnd vdd FILL
XFILL_0__2704_ gnd vdd FILL
XFILL_3__3393_ gnd vdd FILL
XFILL_6__2122_ gnd vdd FILL
XFILL_0__2635_ gnd vdd FILL
XFILL_3__2413_ gnd vdd FILL
XFILL_8__3038_ gnd vdd FILL
XFILL_3__2344_ gnd vdd FILL
XFILL_6__2053_ gnd vdd FILL
XFILL_3__2275_ gnd vdd FILL
XFILL_0__2566_ gnd vdd FILL
XFILL_0__2497_ gnd vdd FILL
XFILL184650x175650 gnd vdd FILL
XFILL_6__2955_ gnd vdd FILL
XFILL_9__2664_ gnd vdd FILL
XFILL_0__3118_ gnd vdd FILL
XFILL_6__2886_ gnd vdd FILL
XFILL_6__1906_ gnd vdd FILL
XFILL_8_BUFX2_insert4 gnd vdd FILL
XFILL_4__1970_ gnd vdd FILL
XFILL_0__3049_ gnd vdd FILL
XFILL_6__1837_ gnd vdd FILL
XFILL_6__3507_ gnd vdd FILL
XFILL_6__1768_ gnd vdd FILL
XFILL_7__2300_ gnd vdd FILL
X_2628_ _2630_/A _2635_/B _2629_/B vdd gnd XOR2X1
XFILL_1__2813_ gnd vdd FILL
X_2559_ _3228_/A _2572_/B _2559_/C _2560_/A vdd gnd OAI21X1
XFILL_6__1699_ gnd vdd FILL
XFILL_4__2522_ gnd vdd FILL
XFILL_6__3438_ gnd vdd FILL
XFILL_7__2231_ gnd vdd FILL
XFILL_1__2744_ gnd vdd FILL
XFILL_7__2162_ gnd vdd FILL
XFILL_6__3369_ gnd vdd FILL
XFILL_4__2453_ gnd vdd FILL
XFILL_4__2384_ gnd vdd FILL
XFILL_1__2675_ gnd vdd FILL
XFILL_7__2093_ gnd vdd FILL
XFILL_2__2020_ gnd vdd FILL
XFILL_4__3005_ gnd vdd FILL
XFILL_1__3227_ gnd vdd FILL
XFILL_7__2995_ gnd vdd FILL
XFILL_7__1946_ gnd vdd FILL
XFILL_1__3158_ gnd vdd FILL
XFILL_1__3089_ gnd vdd FILL
XFILL_7__1877_ gnd vdd FILL
XFILL184050x70350 gnd vdd FILL
XFILL_1__2109_ gnd vdd FILL
XFILL_5__2700_ gnd vdd FILL
XFILL_2__2922_ gnd vdd FILL
XFILL_5__2631_ gnd vdd FILL
XFILL_7__3547_ gnd vdd FILL
XFILL_2__2853_ gnd vdd FILL
XFILL_8__2340_ gnd vdd FILL
XFILL_7__3478_ gnd vdd FILL
XFILL_8__2271_ gnd vdd FILL
XFILL_2__1804_ gnd vdd FILL
XFILL_5__2562_ gnd vdd FILL
XFILL_2__2784_ gnd vdd FILL
XFILL_5__2493_ gnd vdd FILL
XFILL_7__2429_ gnd vdd FILL
XFILL_2__1735_ gnd vdd FILL
XFILL_5__3114_ gnd vdd FILL
XFILL_2__3405_ gnd vdd FILL
XFILL_0__2420_ gnd vdd FILL
XFILL_5__3045_ gnd vdd FILL
XFILL_0__2351_ gnd vdd FILL
XFILL_4_CLKBUF1_insert28 gnd vdd FILL
XFILL_3__2060_ gnd vdd FILL
X_1930_ _3317_/Q _3029_/B _1931_/B vdd gnd NAND2X1
XFILL_8__1986_ gnd vdd FILL
XFILL_0__2282_ gnd vdd FILL
XFILL_2__2218_ gnd vdd FILL
XFILL_2__3198_ gnd vdd FILL
X_1861_ _3025_/A _1861_/B _1861_/C _1873_/A vdd gnd NOR3X1
XFILL_2__2149_ gnd vdd FILL
X_3600_ _3600_/A DO[5] vdd gnd BUFX2
XFILL_6__2740_ gnd vdd FILL
X_3531_ _3531_/A _3531_/B _3535_/C vdd gnd NAND2X1
XFILL_3__2962_ gnd vdd FILL
X_1792_ _3163_/A _2340_/A _1984_/B vdd gnd NOR2X1
XFILL_8__2607_ gnd vdd FILL
XFILL_6__2671_ gnd vdd FILL
XFILL_5__2829_ gnd vdd FILL
XFILL_2_CLKBUF1_insert32 gnd vdd FILL
XFILL_3__2893_ gnd vdd FILL
XFILL_8__3587_ gnd vdd FILL
XFILL_3__1913_ gnd vdd FILL
X_3462_ _3514_/B _3484_/B _3514_/A _3484_/C vdd gnd OAI21X1
XFILL_3__1844_ gnd vdd FILL
XFILL_8__2538_ gnd vdd FILL
X_3393_ _3519_/B _3485_/A _3519_/A _3520_/C vdd gnd OAI21X1
XFILL_8__2469_ gnd vdd FILL
X_2413_ _2413_/A _3575_/Q _3252_/Q _2413_/D _2414_/C vdd gnd AOI22X1
X_2344_ _2344_/A _2344_/B _2344_/C _2351_/A vdd gnd NAND3X1
XFILL_3__1775_ gnd vdd FILL
XFILL_3__3514_ gnd vdd FILL
XFILL_6__3223_ gnd vdd FILL
XFILL_0__1997_ gnd vdd FILL
XFILL_3__3445_ gnd vdd FILL
X_2275_ _2814_/A _2275_/B _2279_/B vdd gnd NOR2X1
XFILL_0_BUFX2_insert14 gnd vdd FILL
XFILL_1__2460_ gnd vdd FILL
XFILL_0_BUFX2_insert25 gnd vdd FILL
XFILL_0_BUFX2_insert47 gnd vdd FILL
XFILL_6__3154_ gnd vdd FILL
XFILL_3__3376_ gnd vdd FILL
XFILL_0_BUFX2_insert58 gnd vdd FILL
XFILL_6__3085_ gnd vdd FILL
XFILL_0__3598_ gnd vdd FILL
XFILL_1__2391_ gnd vdd FILL
XFILL_0__2618_ gnd vdd FILL
XFILL_0_BUFX2_insert69 gnd vdd FILL
XFILL_6__2105_ gnd vdd FILL
XFILL_6__2036_ gnd vdd FILL
XFILL_3__2327_ gnd vdd FILL
XFILL_0__2549_ gnd vdd FILL
XFILL_3__2258_ gnd vdd FILL
XFILL_3__2189_ gnd vdd FILL
XFILL_1__3012_ gnd vdd FILL
XFILL_7__2780_ gnd vdd FILL
XFILL_7__1800_ gnd vdd FILL
XFILL_6__2938_ gnd vdd FILL
XFILL_7__1731_ gnd vdd FILL
XFILL_4__1953_ gnd vdd FILL
XFILL_7__3401_ gnd vdd FILL
XFILL_6__2869_ gnd vdd FILL
XFILL_4__1884_ gnd vdd FILL
XFILL_4__3554_ gnd vdd FILL
XFILL_4__3485_ gnd vdd FILL
XFILL_7__2214_ gnd vdd FILL
XFILL_4__2505_ gnd vdd FILL
XFILL_7__3194_ gnd vdd FILL
XFILL_1__2727_ gnd vdd FILL
XFILL_4__2436_ gnd vdd FILL
XFILL_7__2145_ gnd vdd FILL
XFILL_1__2658_ gnd vdd FILL
XFILL_7__2076_ gnd vdd FILL
XFILL_4__2367_ gnd vdd FILL
XFILL_2__3121_ gnd vdd FILL
XFILL_4__2298_ gnd vdd FILL
XFILL_1__2589_ gnd vdd FILL
XFILL_2__3052_ gnd vdd FILL
XFILL_8__1840_ gnd vdd FILL
XFILL_2__2003_ gnd vdd FILL
XFILL_7__2978_ gnd vdd FILL
XFILL_8__1771_ gnd vdd FILL
XFILL_7__1929_ gnd vdd FILL
XFILL_8__3510_ gnd vdd FILL
XFILL_5__1993_ gnd vdd FILL
XFILL_8__3441_ gnd vdd FILL
XFILL_2__2905_ gnd vdd FILL
XFILL_8__3372_ gnd vdd FILL
XFILL_0__1920_ gnd vdd FILL
XFILL_8__2323_ gnd vdd FILL
XFILL_5__3594_ gnd vdd FILL
XFILL_5__2614_ gnd vdd FILL
XFILL_2__2836_ gnd vdd FILL
XFILL_0__1851_ gnd vdd FILL
XFILL_5__2545_ gnd vdd FILL
XFILL_8__2254_ gnd vdd FILL
XFILL_2__2767_ gnd vdd FILL
XFILL_8__2185_ gnd vdd FILL
XFILL_5__2476_ gnd vdd FILL
XFILL_2__1718_ gnd vdd FILL
XFILL_0__1782_ gnd vdd FILL
XFILL_7_BUFX2_insert20 gnd vdd FILL
XFILL_0__3521_ gnd vdd FILL
X_2060_ _2060_/A _2060_/B _3003_/S _2176_/A vdd gnd NAND3X1
XFILL_2__2698_ gnd vdd FILL
XFILL_3__3230_ gnd vdd FILL
XFILL_0__3452_ gnd vdd FILL
XFILL_7_BUFX2_insert64 gnd vdd FILL
XFILL_7_BUFX2_insert42 gnd vdd FILL
XFILL_7_BUFX2_insert53 gnd vdd FILL
XFILL_7_BUFX2_insert97 gnd vdd FILL
XFILL_0__2403_ gnd vdd FILL
XFILL_7_BUFX2_insert75 gnd vdd FILL
XFILL_3__3161_ gnd vdd FILL
XFILL_7_BUFX2_insert86 gnd vdd FILL
XFILL_3__2112_ gnd vdd FILL
XFILL_5__3028_ gnd vdd FILL
XFILL_3__3092_ gnd vdd FILL
XFILL_0__3383_ gnd vdd FILL
XFILL_3__2043_ gnd vdd FILL
X_2962_ _2995_/A _3023_/B vdd gnd INVX1
XFILL_0__2334_ gnd vdd FILL
XFILL_0__2265_ gnd vdd FILL
XFILL184350x150 gnd vdd FILL
X_1913_ _1913_/A _2521_/C vdd gnd INVX1
X_2893_ _3284_/Q _2898_/A vdd gnd INVX1
XFILL_8__1969_ gnd vdd FILL
XFILL_0__2196_ gnd vdd FILL
XFILL_6__2723_ gnd vdd FILL
X_1844_ _1891_/A _1858_/B _2966_/B vdd gnd NAND2X1
XFILL_3__2945_ gnd vdd FILL
X_1775_ _2057_/A _1933_/C _1782_/B vdd gnd NOR2X1
X_3514_ _3514_/A _3514_/B _3518_/B _3515_/A vdd gnd OAI21X1
XFILL_1__1960_ gnd vdd FILL
XFILL_6__2654_ gnd vdd FILL
X_3445_ _3445_/A _3451_/B _3445_/C _3455_/C _3449_/C vdd gnd AOI22X1
XFILL_3__2876_ gnd vdd FILL
XFILL_6__2585_ gnd vdd FILL
XFILL_3__1827_ gnd vdd FILL
XFILL_1__1891_ gnd vdd FILL
X_3376_ _3468_/A _3445_/A vdd gnd INVX2
XFILL_3__1758_ gnd vdd FILL
XFILL_1__3561_ gnd vdd FILL
X_2327_ _2327_/A _2327_/B _2328_/B vdd gnd NAND2X1
XFILL_1__3492_ gnd vdd FILL
X_2258_ _2853_/A _2297_/B vdd gnd INVX1
XFILL_3__1689_ gnd vdd FILL
XFILL_6__3206_ gnd vdd FILL
XFILL_1__2512_ gnd vdd FILL
XFILL_6__3137_ gnd vdd FILL
XFILL_3__3428_ gnd vdd FILL
XFILL_1__2443_ gnd vdd FILL
XFILL_4__2221_ gnd vdd FILL
X_2189_ _2897_/C _2881_/A _2821_/A vdd gnd NAND2X1
XFILL_4__2152_ gnd vdd FILL
XFILL_4__2083_ gnd vdd FILL
XFILL_6__3068_ gnd vdd FILL
XFILL_1__2374_ gnd vdd FILL
XFILL_7__2901_ gnd vdd FILL
XFILL_6__2019_ gnd vdd FILL
XFILL_7__2832_ gnd vdd FILL
XFILL_7__2763_ gnd vdd FILL
XFILL_4__2985_ gnd vdd FILL
XFILL_7__2694_ gnd vdd FILL
XFILL_7__1714_ gnd vdd FILL
XFILL_4__1936_ gnd vdd FILL
XFILL_4__1867_ gnd vdd FILL
XFILL_4__3537_ gnd vdd FILL
XFILL_5__2330_ gnd vdd FILL
XFILL_2__2621_ gnd vdd FILL
XFILL_4__1798_ gnd vdd FILL
XFILL_2__2552_ gnd vdd FILL
XFILL_4__3468_ gnd vdd FILL
XFILL_5__2261_ gnd vdd FILL
XFILL_7__3177_ gnd vdd FILL
XFILL_4__3399_ gnd vdd FILL
XFILL_4__2419_ gnd vdd FILL
XFILL_2__2483_ gnd vdd FILL
XFILL_7__2128_ gnd vdd FILL
XFILL_5__2192_ gnd vdd FILL
XFILL_8__2941_ gnd vdd FILL
XFILL_0_BUFX2_insert6 gnd vdd FILL
XFILL_7__2059_ gnd vdd FILL
XFILL_2__3104_ gnd vdd FILL
XFILL_8__2872_ gnd vdd FILL
XFILL_8__1823_ gnd vdd FILL
XFILL_2__3035_ gnd vdd FILL
XFILL_0__2050_ gnd vdd FILL
XFILL_8__1754_ gnd vdd FILL
XFILL_5__1976_ gnd vdd FILL
XFILL_8__3424_ gnd vdd FILL
XFILL_3__2730_ gnd vdd FILL
XFILL_0__2952_ gnd vdd FILL
XFILL_3__2661_ gnd vdd FILL
XFILL_2__2819_ gnd vdd FILL
XFILL_0__2883_ gnd vdd FILL
XFILL_6__2370_ gnd vdd FILL
XFILL_8__2306_ gnd vdd FILL
XFILL_0__1903_ gnd vdd FILL
X_3230_ _3230_/A _3230_/B _3230_/C _3362_/D vdd gnd OAI21X1
XFILL_8__2237_ gnd vdd FILL
XFILL_5__2528_ gnd vdd FILL
XFILL_0__1834_ gnd vdd FILL
XFILL_3__2592_ gnd vdd FILL
X_3161_ _3237_/Q _3161_/B _3161_/C _3162_/A vdd gnd OAI21X1
X_2112_ _2112_/A _2320_/C _2113_/C vdd gnd AND2X2
XFILL_5__2459_ gnd vdd FILL
XFILL_0__1765_ gnd vdd FILL
XFILL_8__2168_ gnd vdd FILL
X_3092_ _3092_/A _3107_/B vdd gnd INVX2
XFILL_0__3504_ gnd vdd FILL
X_2043_ _2854_/A _2887_/B _2044_/B vdd gnd NAND2X1
XFILL_0__1696_ gnd vdd FILL
XFILL_3__3213_ gnd vdd FILL
XFILL_8__2099_ gnd vdd FILL
XFILL_0__3435_ gnd vdd FILL
XFILL_3__3144_ gnd vdd FILL
XFILL_0__3366_ gnd vdd FILL
XFILL_3__3075_ gnd vdd FILL
XFILL_0__2317_ gnd vdd FILL
XFILL_9__3602_ gnd vdd FILL
XFILL_3__2026_ gnd vdd FILL
X_2945_ reset _2957_/C _3301_/Q _2946_/C vdd gnd OAI21X1
XFILL_1__2090_ gnd vdd FILL
XFILL_0__2248_ gnd vdd FILL
X_2876_ _3035_/B _2878_/B _2876_/C _2878_/C _3278_/D vdd gnd OAI22X1
XFILL_0__2179_ gnd vdd FILL
X_1827_ _2659_/B _3189_/C _2952_/A _1831_/D _3411_/A vdd gnd OAI22X1
XFILL_3_BUFX2_insert40 gnd vdd FILL
XFILL_6__2706_ gnd vdd FILL
XFILL_4__2770_ gnd vdd FILL
XFILL_3__2928_ gnd vdd FILL
XFILL_3_BUFX2_insert51 gnd vdd FILL
XFILL_3_BUFX2_insert62 gnd vdd FILL
XFILL_1__2992_ gnd vdd FILL
XFILL_3_BUFX2_insert73 gnd vdd FILL
XFILL_4__1721_ gnd vdd FILL
X_1758_ _1846_/B _3144_/A _2432_/A _2448_/C vdd gnd OAI21X1
XFILL_6__2637_ gnd vdd FILL
XFILL_3_BUFX2_insert95 gnd vdd FILL
XFILL_3__2859_ gnd vdd FILL
XFILL_3_BUFX2_insert84 gnd vdd FILL
X_1689_ DI[0] _2675_/A _1690_/C vdd gnd NAND2X1
XFILL_1__1943_ gnd vdd FILL
XFILL_1__1874_ gnd vdd FILL
X_3428_ _3428_/A _3428_/B _3428_/C _3431_/A vdd gnd OAI21X1
XFILL_6__2568_ gnd vdd FILL
XFILL_7__3100_ gnd vdd FILL
XFILL_6__2499_ gnd vdd FILL
X_3359_ _3359_/D vdd _3362_/R _3362_/CLK _3359_/Q vdd gnd DFFSR
XFILL_7__3031_ gnd vdd FILL
XFILL_1__3544_ gnd vdd FILL
XFILL_1__3475_ gnd vdd FILL
XFILL_4__2204_ gnd vdd FILL
XFILL_1__2426_ gnd vdd FILL
XFILL_4__3184_ gnd vdd FILL
XFILL_4__2135_ gnd vdd FILL
XFILL_4__2066_ gnd vdd FILL
XFILL_1__2357_ gnd vdd FILL
XFILL_1__2288_ gnd vdd FILL
XFILL_7__2815_ gnd vdd FILL
XFILL_7__2746_ gnd vdd FILL
XFILL_5__1830_ gnd vdd FILL
XFILL_4__2968_ gnd vdd FILL
XFILL_5__1761_ gnd vdd FILL
XFILL_5__3500_ gnd vdd FILL
XFILL_4__1919_ gnd vdd FILL
XFILL_7__2677_ gnd vdd FILL
XFILL_2__1983_ gnd vdd FILL
XFILL_4__2899_ gnd vdd FILL
XFILL_5__3431_ gnd vdd FILL
XFILL_5__1692_ gnd vdd FILL
XFILL_8__3140_ gnd vdd FILL
XFILL_8__3071_ gnd vdd FILL
XFILL_2__2604_ gnd vdd FILL
XFILL_8__2022_ gnd vdd FILL
XFILL_5__2313_ gnd vdd FILL
XFILL_2__3584_ gnd vdd FILL
XFILL_7__3229_ gnd vdd FILL
XFILL_5__2244_ gnd vdd FILL
XFILL_2__2535_ gnd vdd FILL
XFILL182250x101550 gnd vdd FILL
XFILL_2__2466_ gnd vdd FILL
XFILL_5__2175_ gnd vdd FILL
XFILL_8__2924_ gnd vdd FILL
XFILL_2__2397_ gnd vdd FILL
XFILL_0__3220_ gnd vdd FILL
XFILL_0__3151_ gnd vdd FILL
XFILL_8__2855_ gnd vdd FILL
XFILL_7_CLKBUF1_insert32 gnd vdd FILL
XFILL_0__2102_ gnd vdd FILL
XFILL_0__3082_ gnd vdd FILL
XFILL_6__1870_ gnd vdd FILL
XFILL_8__2786_ gnd vdd FILL
XFILL_2__3018_ gnd vdd FILL
X_2730_ _2734_/B _2773_/B _2730_/C _2732_/B vdd gnd OAI21X1
XFILL_8__1806_ gnd vdd FILL
XFILL_0__2033_ gnd vdd FILL
XFILL_8__1737_ gnd vdd FILL
X_2661_ _3354_/Q _2662_/A vdd gnd INVX1
XFILL_5__1959_ gnd vdd FILL
XFILL_6__3540_ gnd vdd FILL
X_2592_ _2692_/A _2670_/B _2756_/B vdd gnd NOR2X1
XFILL_6__3471_ gnd vdd FILL
XFILL_8__3407_ gnd vdd FILL
XFILL_3__2713_ gnd vdd FILL
XFILL_0__2935_ gnd vdd FILL
XFILL_6__2422_ gnd vdd FILL
XFILL_6__2353_ gnd vdd FILL
X_3213_ _3215_/A _3213_/B _3213_/C _3354_/D vdd gnd OAI21X1
XFILL_3__2644_ gnd vdd FILL
XFILL_0__2866_ gnd vdd FILL
XFILL_3__2575_ gnd vdd FILL
XFILL_0__2797_ gnd vdd FILL
XFILL_6__2284_ gnd vdd FILL
XFILL_0__1817_ gnd vdd FILL
X_3144_ _3144_/A _3144_/B _3144_/C _3181_/A vdd gnd AOI21X1
X_3075_ _3090_/A _3139_/A _3075_/C _3320_/D vdd gnd OAI21X1
XFILL_0__1748_ gnd vdd FILL
X_2026_ _2889_/B _2889_/C _2857_/A vdd gnd AND2X2
XFILL_0__3418_ gnd vdd FILL
XFILL_1__2211_ gnd vdd FILL
XFILL_3__3127_ gnd vdd FILL
XFILL_1__3191_ gnd vdd FILL
XFILL_3__3058_ gnd vdd FILL
XFILL_1__2142_ gnd vdd FILL
X_2928_ _2928_/A _2928_/B _2928_/C _2929_/A vdd gnd OAI21X1
XFILL_1__2073_ gnd vdd FILL
XFILL_3__2009_ gnd vdd FILL
XFILL_7__3580_ gnd vdd FILL
XBUFX2_insert27 _2580_/Y _3291_/R vdd gnd BUFX2
XFILL_7__2600_ gnd vdd FILL
XBUFX2_insert16 _1907_/Y _2669_/C vdd gnd BUFX2
XFILL_9__3516_ gnd vdd FILL
X_2859_ _2859_/A _2921_/A _2885_/B _2866_/C vdd gnd AOI21X1
XBUFX2_insert49 _3307_/Q _2006_/A vdd gnd BUFX2
XFILL_6__1999_ gnd vdd FILL
XFILL_4__2822_ gnd vdd FILL
XFILL_7__2531_ gnd vdd FILL
XFILL_4__2753_ gnd vdd FILL
XFILL_1__2975_ gnd vdd FILL
XFILL_4__1704_ gnd vdd FILL
XFILL_7__2462_ gnd vdd FILL
XFILL_1__1926_ gnd vdd FILL
XFILL_7__2393_ gnd vdd FILL
XFILL_4__2684_ gnd vdd FILL
XFILL_8_BUFX2_insert19 gnd vdd FILL
XFILL_1__1857_ gnd vdd FILL
XFILL_1__1788_ gnd vdd FILL
XFILL_1__3527_ gnd vdd FILL
XFILL_7__3014_ gnd vdd FILL
XFILL_2__2320_ gnd vdd FILL
XFILL_1__3458_ gnd vdd FILL
XFILL_2__2251_ gnd vdd FILL
XFILL_4__3167_ gnd vdd FILL
XFILL_1__3389_ gnd vdd FILL
XFILL_2__2182_ gnd vdd FILL
XFILL_4__2118_ gnd vdd FILL
XFILL_1__2409_ gnd vdd FILL
XFILL_4__3098_ gnd vdd FILL
XFILL_5__2931_ gnd vdd FILL
XFILL_4__2049_ gnd vdd FILL
XFILL_8__2640_ gnd vdd FILL
XFILL_5__2862_ gnd vdd FILL
XFILL_8__2571_ gnd vdd FILL
XFILL_5__1813_ gnd vdd FILL
XFILL_5__2793_ gnd vdd FILL
XFILL_7__2729_ gnd vdd FILL
XFILL_5__1744_ gnd vdd FILL
XFILL_2__1966_ gnd vdd FILL
XFILL_8__3123_ gnd vdd FILL
XFILL182550x105450 gnd vdd FILL
XFILL_5__3414_ gnd vdd FILL
XFILL_2__1897_ gnd vdd FILL
XFILL_0__2720_ gnd vdd FILL
XFILL_3__2360_ gnd vdd FILL
XFILL_8__3054_ gnd vdd FILL
XFILL_0__2651_ gnd vdd FILL
XFILL_8__2005_ gnd vdd FILL
XFILL_2__2518_ gnd vdd FILL
XFILL_0__2582_ gnd vdd FILL
XFILL_2__3498_ gnd vdd FILL
XFILL_5__2227_ gnd vdd FILL
XFILL_3__2291_ gnd vdd FILL
XFILL_5__2158_ gnd vdd FILL
XFILL_2__2449_ gnd vdd FILL
XFILL_8__2907_ gnd vdd FILL
XFILL_6__2971_ gnd vdd FILL
XFILL_5__2089_ gnd vdd FILL
XFILL_0__3203_ gnd vdd FILL
XFILL_0__3134_ gnd vdd FILL
XFILL_6__1922_ gnd vdd FILL
XFILL_8__2838_ gnd vdd FILL
XFILL_0__3065_ gnd vdd FILL
XFILL_6__1853_ gnd vdd FILL
XFILL_0__2016_ gnd vdd FILL
X_2713_ _2759_/A _2759_/B _3292_/D _2720_/A vdd gnd OAI21X1
XFILL_8__2769_ gnd vdd FILL
XFILL182850x35250 gnd vdd FILL
XFILL_6__1784_ gnd vdd FILL
X_2644_ _2644_/A _2748_/B _2669_/C _2645_/C vdd gnd OAI21X1
XFILL_6__3523_ gnd vdd FILL
X_2575_ _3279_/Q _3309_/Q _3339_/D vdd gnd AND2X2
XFILL_6__3454_ gnd vdd FILL
XFILL_6__2405_ gnd vdd FILL
XFILL_1__2760_ gnd vdd FILL
XFILL_0__2918_ gnd vdd FILL
XFILL_6__3385_ gnd vdd FILL
XFILL_1__1711_ gnd vdd FILL
XFILL_1__2691_ gnd vdd FILL
XFILL_3__2627_ gnd vdd FILL
XFILL_0__2849_ gnd vdd FILL
XFILL_6__2336_ gnd vdd FILL
X_3127_ _3127_/A _3127_/B _3143_/B vdd gnd NAND2X1
XFILL_6__2267_ gnd vdd FILL
XFILL_3__2558_ gnd vdd FILL
XFILL_3__2489_ gnd vdd FILL
X_3058_ _3059_/B _3059_/A _3060_/D vdd gnd AND2X2
XFILL_4__3021_ gnd vdd FILL
XFILL_6__2198_ gnd vdd FILL
X_2009_ _2009_/A _3256_/Q _2406_/D _2889_/C vdd gnd OAI21X1
XFILL_7__1962_ gnd vdd FILL
XFILL_1__3174_ gnd vdd FILL
XFILL_1__2125_ gnd vdd FILL
XFILL_7__1893_ gnd vdd FILL
XFILL_1__2056_ gnd vdd FILL
XFILL_4__2805_ gnd vdd FILL
XFILL_7__3563_ gnd vdd FILL
XFILL_7__3494_ gnd vdd FILL
XFILL_2__1820_ gnd vdd FILL
XFILL_7__2514_ gnd vdd FILL
XFILL_4__2736_ gnd vdd FILL
XFILL_7__2445_ gnd vdd FILL
XFILL_1__2958_ gnd vdd FILL
XFILL_2__1751_ gnd vdd FILL
XFILL_4__2667_ gnd vdd FILL
XFILL_1__2889_ gnd vdd FILL
XFILL_7__2376_ gnd vdd FILL
XFILL_1__1909_ gnd vdd FILL
XFILL_2__3421_ gnd vdd FILL
XFILL_4__2598_ gnd vdd FILL
XFILL_5__3130_ gnd vdd FILL
XFILL_5__3061_ gnd vdd FILL
XFILL_5__2012_ gnd vdd FILL
XFILL_2__2303_ gnd vdd FILL
XFILL_4__3219_ gnd vdd FILL
XFILL_5_BUFX2_insert1 gnd vdd FILL
XFILL_2__2234_ gnd vdd FILL
XFILL_2__2165_ gnd vdd FILL
XFILL_5__2914_ gnd vdd FILL
XFILL_4_BUFX2_insert17 gnd vdd FILL
XFILL_4_BUFX2_insert39 gnd vdd FILL
XFILL_2__2096_ gnd vdd FILL
XFILL_8__2623_ gnd vdd FILL
XFILL_5__2845_ gnd vdd FILL
XFILL182850x109350 gnd vdd FILL
XFILL_8__2554_ gnd vdd FILL
XFILL_3__1860_ gnd vdd FILL
XFILL182550x117150 gnd vdd FILL
XFILL_5__2776_ gnd vdd FILL
XFILL_2__2998_ gnd vdd FILL
XFILL_3__1791_ gnd vdd FILL
XFILL_8__2485_ gnd vdd FILL
XFILL_5__1727_ gnd vdd FILL
X_2360_ _3271_/Q _2841_/A vdd gnd INVX1
XFILL_3__3530_ gnd vdd FILL
XFILL_2__1949_ gnd vdd FILL
XFILL_3__3461_ gnd vdd FILL
X_2291_ _3144_/B _3146_/A _2294_/B vdd gnd NAND2X1
XFILL_8__3106_ gnd vdd FILL
XFILL_3__2412_ gnd vdd FILL
XFILL_0__2703_ gnd vdd FILL
XFILL_6__3170_ gnd vdd FILL
XFILL_3__3392_ gnd vdd FILL
XFILL_8__3037_ gnd vdd FILL
XFILL_6__2121_ gnd vdd FILL
XFILL_0__2634_ gnd vdd FILL
XFILL_3__2343_ gnd vdd FILL
XFILL_6__2052_ gnd vdd FILL
XFILL_3__2274_ gnd vdd FILL
XFILL_0__2565_ gnd vdd FILL
XFILL_0__2496_ gnd vdd FILL
XFILL_6__2954_ gnd vdd FILL
XFILL_6__1905_ gnd vdd FILL
XFILL_0__3117_ gnd vdd FILL
XFILL_6__2885_ gnd vdd FILL
XFILL_8_BUFX2_insert5 gnd vdd FILL
XFILL_0__3048_ gnd vdd FILL
XFILL_6__1836_ gnd vdd FILL
XFILL_6__1767_ gnd vdd FILL
XFILL_6__3506_ gnd vdd FILL
XFILL_3__1989_ gnd vdd FILL
X_2627_ _2627_/A _2671_/B _2638_/B _2635_/B vdd gnd OAI21X1
XFILL_1__2812_ gnd vdd FILL
XFILL_4__2521_ gnd vdd FILL
X_2558_ _3361_/Q _2691_/A _2558_/C _2559_/C vdd gnd AOI21X1
XFILL_6__1698_ gnd vdd FILL
XFILL_6__3437_ gnd vdd FILL
X_2489_ _2646_/A _2574_/B _2489_/C _2490_/C vdd gnd OAI21X1
XFILL_1__2743_ gnd vdd FILL
XFILL_7__2230_ gnd vdd FILL
XFILL_7__2161_ gnd vdd FILL
XFILL_6__3368_ gnd vdd FILL
XFILL_4__2452_ gnd vdd FILL
XFILL_4__2383_ gnd vdd FILL
XFILL_6__2319_ gnd vdd FILL
XFILL_1__2674_ gnd vdd FILL
XFILL_7__2092_ gnd vdd FILL
XFILL_4__3004_ gnd vdd FILL
XFILL_1__3226_ gnd vdd FILL
XFILL_7__2994_ gnd vdd FILL
XFILL_7__1945_ gnd vdd FILL
XFILL184350x54750 gnd vdd FILL
XFILL_1__3157_ gnd vdd FILL
XFILL_7__1876_ gnd vdd FILL
XFILL_1__3088_ gnd vdd FILL
XFILL_1__2108_ gnd vdd FILL
XFILL_2__2921_ gnd vdd FILL
XFILL_1__2039_ gnd vdd FILL
XFILL_7__3546_ gnd vdd FILL
XFILL_5__2630_ gnd vdd FILL
XFILL_2__2852_ gnd vdd FILL
XFILL_5__2561_ gnd vdd FILL
XFILL_7__3477_ gnd vdd FILL
XFILL_8__2270_ gnd vdd FILL
XFILL_2__2783_ gnd vdd FILL
XFILL_2__1803_ gnd vdd FILL
XFILL_4__2719_ gnd vdd FILL
XFILL_7__2428_ gnd vdd FILL
XFILL_5__2492_ gnd vdd FILL
XFILL_2__1734_ gnd vdd FILL
XFILL_7__2359_ gnd vdd FILL
XFILL_5__3113_ gnd vdd FILL
XFILL_2__3404_ gnd vdd FILL
XFILL_5__3044_ gnd vdd FILL
XFILL_0__2350_ gnd vdd FILL
XFILL_0__2281_ gnd vdd FILL
XFILL_2__2217_ gnd vdd FILL
XFILL_8__1985_ gnd vdd FILL
XFILL_4_CLKBUF1_insert29 gnd vdd FILL
XFILL_2__3197_ gnd vdd FILL
X_1860_ _1860_/A _3286_/Q _1871_/A _1879_/C vdd gnd AOI21X1
XFILL_2__2148_ gnd vdd FILL
X_1791_ _3189_/C _3163_/A vdd gnd INVX1
XFILL_2__2079_ gnd vdd FILL
X_3530_ _3532_/A _3531_/A vdd gnd INVX1
XFILL_3__2961_ gnd vdd FILL
XFILL_8__2606_ gnd vdd FILL
XFILL_6__2670_ gnd vdd FILL
XFILL_5__2828_ gnd vdd FILL
XFILL_3__2892_ gnd vdd FILL
XFILL_2_CLKBUF1_insert33 gnd vdd FILL
XFILL184050x105450 gnd vdd FILL
XFILL_8__3586_ gnd vdd FILL
XFILL_3__1912_ gnd vdd FILL
X_3461_ _3461_/A _3461_/B _3473_/A _3544_/A vdd gnd OAI21X1
XFILL_3__1843_ gnd vdd FILL
XFILL_8__2537_ gnd vdd FILL
X_3392_ _3568_/Q _3539_/A vdd gnd INVX1
X_2412_ _2416_/A _2412_/B _2412_/C _3599_/A vdd gnd OAI21X1
XFILL_8__2468_ gnd vdd FILL
XFILL_5__2759_ gnd vdd FILL
XFILL_3__3513_ gnd vdd FILL
X_2343_ _2343_/A _2343_/B _2344_/C vdd gnd NOR2X1
XFILL_3__1774_ gnd vdd FILL
XFILL_8__2399_ gnd vdd FILL
XFILL_6__3222_ gnd vdd FILL
XFILL_0__1996_ gnd vdd FILL
XFILL_3__3444_ gnd vdd FILL
X_2274_ _2814_/A _3148_/B _2274_/C _2298_/D _2352_/B vdd gnd AOI22X1
XFILL_6__3153_ gnd vdd FILL
XFILL_0_BUFX2_insert15 gnd vdd FILL
XFILL_6__2104_ gnd vdd FILL
XFILL_0_BUFX2_insert26 gnd vdd FILL
XFILL_0_BUFX2_insert48 gnd vdd FILL
XFILL_3__3375_ gnd vdd FILL
XFILL_0_BUFX2_insert59 gnd vdd FILL
XFILL_6__3084_ gnd vdd FILL
XFILL_3__2326_ gnd vdd FILL
XFILL_1__2390_ gnd vdd FILL
XFILL_0__3597_ gnd vdd FILL
XFILL_0__2617_ gnd vdd FILL
XFILL_6__2035_ gnd vdd FILL
XFILL_0__2548_ gnd vdd FILL
XFILL_3__2257_ gnd vdd FILL
XFILL_3__2188_ gnd vdd FILL
XFILL_0__2479_ gnd vdd FILL
XFILL_1__3011_ gnd vdd FILL
XFILL_7__1730_ gnd vdd FILL
XFILL_6__2937_ gnd vdd FILL
XFILL_6__2868_ gnd vdd FILL
X_1989_ _3568_/Q _3283_/Q _2066_/A vdd gnd OR2X2
XFILL_4__1952_ gnd vdd FILL
XFILL_7__3400_ gnd vdd FILL
XFILL_4__1883_ gnd vdd FILL
XFILL_6__2799_ gnd vdd FILL
XFILL_6__1819_ gnd vdd FILL
XFILL_4__3553_ gnd vdd FILL
XFILL_4__3484_ gnd vdd FILL
XFILL_7__2213_ gnd vdd FILL
XFILL_4__2504_ gnd vdd FILL
XFILL184650x31350 gnd vdd FILL
XFILL_1__2726_ gnd vdd FILL
XFILL_7__3193_ gnd vdd FILL
XFILL_4__2435_ gnd vdd FILL
XFILL_7__2144_ gnd vdd FILL
XFILL_1__2657_ gnd vdd FILL
XFILL_7__2075_ gnd vdd FILL
XFILL_4__2366_ gnd vdd FILL
XFILL_2__3120_ gnd vdd FILL
XFILL_4__2297_ gnd vdd FILL
XFILL_1__2588_ gnd vdd FILL
XFILL181350x74250 gnd vdd FILL
XFILL_2__3051_ gnd vdd FILL
XFILL_2__2002_ gnd vdd FILL
XFILL_7__2977_ gnd vdd FILL
XFILL_8__1770_ gnd vdd FILL
XFILL_1__3209_ gnd vdd FILL
XFILL_7__1928_ gnd vdd FILL
XFILL_5__1992_ gnd vdd FILL
XFILL_8__3440_ gnd vdd FILL
XFILL_7__1859_ gnd vdd FILL
XFILL_2__2904_ gnd vdd FILL
XFILL_8__3371_ gnd vdd FILL
XFILL_5__2613_ gnd vdd FILL
XFILL_2__2835_ gnd vdd FILL
XFILL_7__3529_ gnd vdd FILL
XFILL_8__2322_ gnd vdd FILL
XFILL_5__3593_ gnd vdd FILL
XFILL_8__2253_ gnd vdd FILL
XFILL_5__2544_ gnd vdd FILL
XFILL_0__1850_ gnd vdd FILL
XFILL_5__2475_ gnd vdd FILL
XFILL_2__2766_ gnd vdd FILL
XFILL_8__2184_ gnd vdd FILL
XFILL_2__1717_ gnd vdd FILL
XFILL_2__2697_ gnd vdd FILL
XFILL_0__1781_ gnd vdd FILL
XFILL_0__3520_ gnd vdd FILL
XFILL_7_BUFX2_insert21 gnd vdd FILL
XFILL_7_BUFX2_insert10 gnd vdd FILL
XFILL_0__3451_ gnd vdd FILL
XFILL_7_BUFX2_insert43 gnd vdd FILL
XFILL_7_BUFX2_insert65 gnd vdd FILL
XFILL_7_BUFX2_insert54 gnd vdd FILL
XFILL_0__2402_ gnd vdd FILL
XFILL_7_BUFX2_insert87 gnd vdd FILL
XFILL_3__3160_ gnd vdd FILL
XFILL_7_BUFX2_insert76 gnd vdd FILL
XFILL_3__3091_ gnd vdd FILL
XFILL_0__3382_ gnd vdd FILL
XFILL_5__3027_ gnd vdd FILL
XFILL_3__2111_ gnd vdd FILL
XFILL_3__2042_ gnd vdd FILL
X_2961_ _3260_/Q _3006_/B _2995_/A vdd gnd NOR2X1
XFILL_0__2333_ gnd vdd FILL
XFILL_0__2264_ gnd vdd FILL
XFILL184350x109350 gnd vdd FILL
X_1912_ _3217_/A _2700_/B _1913_/A vdd gnd NOR2X1
XFILL_8__1968_ gnd vdd FILL
X_2892_ _2892_/A _2892_/B _2892_/C _3283_/D vdd gnd OAI21X1
XFILL184050x117150 gnd vdd FILL
XFILL_0__2195_ gnd vdd FILL
XFILL_8__1899_ gnd vdd FILL
X_1843_ _1843_/A _1843_/B _1843_/C _1856_/A vdd gnd NAND3X1
XFILL_6__2722_ gnd vdd FILL
XFILL_3__2944_ gnd vdd FILL
X_1774_ _1933_/C _1783_/B _3149_/C vdd gnd NOR2X1
X_3513_ _3518_/B _3518_/A _3516_/C vdd gnd NAND2X1
XFILL_6__2653_ gnd vdd FILL
X_3444_ _3451_/B _3460_/B _3453_/B _3445_/C vdd gnd NAND3X1
XFILL_3__2875_ gnd vdd FILL
XFILL_6__2584_ gnd vdd FILL
XFILL_1__1890_ gnd vdd FILL
XFILL_3__1826_ gnd vdd FILL
X_3375_ _3521_/A _3466_/C _3384_/C vdd gnd NAND2X1
XFILL_3__1757_ gnd vdd FILL
XFILL_0__1979_ gnd vdd FILL
XFILL_1__3560_ gnd vdd FILL
X_2326_ _2326_/A _2326_/B _2326_/C _3236_/D vdd gnd OAI21X1
XFILL_6__3205_ gnd vdd FILL
XFILL_1__3491_ gnd vdd FILL
XFILL_3__3427_ gnd vdd FILL
X_2257_ _2312_/C _2257_/B _2310_/B _2264_/A vdd gnd NAND3X1
XFILL_4__2220_ gnd vdd FILL
XFILL_1__2511_ gnd vdd FILL
XFILL_3__1688_ gnd vdd FILL
XFILL_6__3136_ gnd vdd FILL
XFILL_1__2442_ gnd vdd FILL
X_2188_ _2824_/A _2922_/A _2881_/A vdd gnd NOR2X1
XFILL_6__3067_ gnd vdd FILL
XFILL_4__2151_ gnd vdd FILL
XFILL_6__2018_ gnd vdd FILL
XFILL_3__2309_ gnd vdd FILL
XFILL_4__2082_ gnd vdd FILL
XFILL_1__2373_ gnd vdd FILL
XFILL_7__2900_ gnd vdd FILL
XFILL_7__2831_ gnd vdd FILL
XFILL_7__2762_ gnd vdd FILL
XFILL_4__2984_ gnd vdd FILL
XFILL_4__1935_ gnd vdd FILL
XFILL_7__2693_ gnd vdd FILL
XFILL_7__1713_ gnd vdd FILL
XFILL184650x43050 gnd vdd FILL
XFILL_4__1866_ gnd vdd FILL
XFILL_4__1797_ gnd vdd FILL
XFILL_4__3536_ gnd vdd FILL
XFILL_2__2620_ gnd vdd FILL
XFILL_2__2551_ gnd vdd FILL
XFILL_4__3467_ gnd vdd FILL
XFILL_5__2260_ gnd vdd FILL
XFILL184350x78150 gnd vdd FILL
XFILL_1__2709_ gnd vdd FILL
XFILL_7__3176_ gnd vdd FILL
XFILL_4__3398_ gnd vdd FILL
XFILL_5__2191_ gnd vdd FILL
XFILL_4__2418_ gnd vdd FILL
XFILL_2__2482_ gnd vdd FILL
XFILL_7__2127_ gnd vdd FILL
XFILL_4__2349_ gnd vdd FILL
XFILL_8__2940_ gnd vdd FILL
XFILL_7__2058_ gnd vdd FILL
XFILL_0_BUFX2_insert7 gnd vdd FILL
XFILL_2__3103_ gnd vdd FILL
XFILL_8__2871_ gnd vdd FILL
XFILL_2__3034_ gnd vdd FILL
XFILL_8__1822_ gnd vdd FILL
XFILL_8__1753_ gnd vdd FILL
XFILL_5__1975_ gnd vdd FILL
XFILL_8__3423_ gnd vdd FILL
XFILL_0__2951_ gnd vdd FILL
XFILL_0__1902_ gnd vdd FILL
XFILL_3__2660_ gnd vdd FILL
XFILL_2__2818_ gnd vdd FILL
XFILL_8__2305_ gnd vdd FILL
XFILL_0__2882_ gnd vdd FILL
XFILL_5__2527_ gnd vdd FILL
XFILL_3__2591_ gnd vdd FILL
XFILL_8__2236_ gnd vdd FILL
XFILL_2__2749_ gnd vdd FILL
XFILL_0__1833_ gnd vdd FILL
X_3160_ _3160_/A _3160_/B _3160_/C _3161_/C vdd gnd OAI21X1
X_3091_ _3127_/A _3092_/A _3108_/B vdd gnd NAND2X1
XFILL_8__2167_ gnd vdd FILL
XFILL_5__2458_ gnd vdd FILL
X_2111_ _2332_/C _2111_/B _2112_/A vdd gnd AND2X2
XFILL_0__1764_ gnd vdd FILL
X_2042_ _2933_/B _2887_/B vdd gnd INVX1
XFILL_0__3503_ gnd vdd FILL
XFILL_5__2389_ gnd vdd FILL
XFILL_0__1695_ gnd vdd FILL
XFILL_3__3212_ gnd vdd FILL
XFILL_8__2098_ gnd vdd FILL
XFILL_3__3143_ gnd vdd FILL
XFILL_0__3434_ gnd vdd FILL
XFILL_0__3365_ gnd vdd FILL
XFILL_3__3074_ gnd vdd FILL
XFILL_0__2316_ gnd vdd FILL
XFILL183750x171750 gnd vdd FILL
XFILL_3__2025_ gnd vdd FILL
X_2944_ _3043_/A _2956_/B _2944_/C _3300_/D vdd gnd OAI21X1
X_2875_ _2875_/A _2878_/B _2933_/C _2878_/C vdd gnd NAND3X1
XFILL_0__2247_ gnd vdd FILL
XFILL_0__2178_ gnd vdd FILL
X_1826_ _3244_/Q _2659_/B vdd gnd INVX2
XFILL_9__2414_ gnd vdd FILL
XFILL_6__2705_ gnd vdd FILL
XFILL_3__2927_ gnd vdd FILL
XFILL_3_BUFX2_insert63 gnd vdd FILL
XFILL_3_BUFX2_insert74 gnd vdd FILL
XFILL_1__2991_ gnd vdd FILL
X_1757_ _2594_/B _1803_/B _3144_/A vdd gnd NOR2X1
XFILL_4__1720_ gnd vdd FILL
XFILL_3_BUFX2_insert52 gnd vdd FILL
XFILL_6__2636_ gnd vdd FILL
XFILL_3_BUFX2_insert41 gnd vdd FILL
XFILL_3_BUFX2_insert96 gnd vdd FILL
XFILL_3__2858_ gnd vdd FILL
XFILL_3_BUFX2_insert85 gnd vdd FILL
XFILL_1__1942_ gnd vdd FILL
X_1688_ _3290_/Q _1690_/B vdd gnd INVX1
XFILL_1__1873_ gnd vdd FILL
X_3427_ _3442_/B _3428_/A _3466_/B _3428_/C vdd gnd OAI21X1
XFILL_3__1809_ gnd vdd FILL
XFILL_6__2567_ gnd vdd FILL
XFILL_3__2789_ gnd vdd FILL
XFILL_6__2498_ gnd vdd FILL
X_3358_ _3358_/D vdd _3363_/R _3362_/CLK _3358_/Q vdd gnd DFFSR
XFILL_1__3543_ gnd vdd FILL
X_2309_ _2915_/A _2933_/C _2854_/A _2310_/A vdd gnd OAI21X1
XFILL_7__3030_ gnd vdd FILL
X_3289_ _3289_/D vdd _3289_/R _3307_/CLK _3289_/Q vdd gnd DFFSR
XFILL_1__3474_ gnd vdd FILL
XFILL_6__3119_ gnd vdd FILL
XFILL_4__2203_ gnd vdd FILL
XFILL_4__3183_ gnd vdd FILL
XFILL_1__2425_ gnd vdd FILL
XFILL_4__2134_ gnd vdd FILL
XFILL_1__2356_ gnd vdd FILL
XFILL_4__2065_ gnd vdd FILL
XFILL_1__2287_ gnd vdd FILL
XFILL_7__2814_ gnd vdd FILL
XFILL_7__2745_ gnd vdd FILL
XFILL_5__1760_ gnd vdd FILL
XFILL_4__2967_ gnd vdd FILL
XFILL_4__1918_ gnd vdd FILL
XFILL_4__2898_ gnd vdd FILL
XFILL_5__1691_ gnd vdd FILL
XFILL_2__1982_ gnd vdd FILL
XFILL_7__2676_ gnd vdd FILL
XFILL_5__3430_ gnd vdd FILL
XFILL_4__1849_ gnd vdd FILL
XFILL_8__3070_ gnd vdd FILL
XFILL_2__2603_ gnd vdd FILL
XFILL_8__2021_ gnd vdd FILL
XFILL_4__3519_ gnd vdd FILL
XFILL_5__2312_ gnd vdd FILL
XFILL_2__3583_ gnd vdd FILL
XFILL_7__3228_ gnd vdd FILL
XFILL_5__2243_ gnd vdd FILL
XFILL_2__2534_ gnd vdd FILL
XFILL_2__2465_ gnd vdd FILL
XFILL_7__3159_ gnd vdd FILL
XFILL_5__2174_ gnd vdd FILL
XFILL_8__2923_ gnd vdd FILL
XFILL_2__2396_ gnd vdd FILL
XFILL_0__3150_ gnd vdd FILL
XFILL_8__2854_ gnd vdd FILL
XFILL_7_CLKBUF1_insert33 gnd vdd FILL
XFILL_0__2101_ gnd vdd FILL
XFILL_0__3081_ gnd vdd FILL
XFILL_2__3017_ gnd vdd FILL
XFILL_8__2785_ gnd vdd FILL
XFILL_8__1805_ gnd vdd FILL
XFILL_0__2032_ gnd vdd FILL
XFILL_8__1736_ gnd vdd FILL
X_2660_ _2660_/A _2741_/C _2674_/C vdd gnd NOR2X1
XFILL_5__1958_ gnd vdd FILL
XFILL_6__3470_ gnd vdd FILL
X_2591_ _3147_/C _2717_/B _2771_/A _2692_/A vdd gnd NAND3X1
XFILL_8__3406_ gnd vdd FILL
XFILL_5__1889_ gnd vdd FILL
XFILL_6__2421_ gnd vdd FILL
XFILL_3__2712_ gnd vdd FILL
XFILL_0__2934_ gnd vdd FILL
XFILL_3__2643_ gnd vdd FILL
XFILL_5__3559_ gnd vdd FILL
XFILL_0__2865_ gnd vdd FILL
XFILL_6__2352_ gnd vdd FILL
XFILL_9__2061_ gnd vdd FILL
X_3212_ _3214_/A _3214_/B _3354_/Q _3213_/C vdd gnd OAI21X1
XFILL_0__1816_ gnd vdd FILL
XFILL_6__2283_ gnd vdd FILL
XFILL_3__2574_ gnd vdd FILL
X_3143_ _3143_/A _3143_/B _3143_/C _3347_/D vdd gnd OAI21X1
XFILL_0__2796_ gnd vdd FILL
XFILL_8__2219_ gnd vdd FILL
XFILL_8__3199_ gnd vdd FILL
X_3074_ _3320_/Q _3090_/A _3075_/C vdd gnd NAND2X1
XFILL_0__1747_ gnd vdd FILL
X_2025_ _2025_/A _3079_/A _2025_/C _2889_/B vdd gnd OAI21X1
XFILL_0__3417_ gnd vdd FILL
XFILL_1__2210_ gnd vdd FILL
XFILL_3__3126_ gnd vdd FILL
XFILL_1__3190_ gnd vdd FILL
XFILL_3__3057_ gnd vdd FILL
XFILL_1__2141_ gnd vdd FILL
X_2927_ _2927_/A _2927_/B _2928_/C vdd gnd NAND2X1
XFILL_1__2072_ gnd vdd FILL
XFILL_3__2008_ gnd vdd FILL
XBUFX2_insert17 _2580_/Y _3313_/R vdd gnd BUFX2
XBUFX2_insert39 _1734_/Y _2958_/A vdd gnd BUFX2
X_2858_ _2858_/A _2858_/B _2861_/C vdd gnd NOR2X1
XFILL_6__1998_ gnd vdd FILL
XFILL_4__2821_ gnd vdd FILL
XFILL_7__2530_ gnd vdd FILL
X_2789_ _3259_/Q _2814_/A _2790_/C vdd gnd NAND2X1
X_1809_ _2123_/A _1891_/B _2781_/B vdd gnd NAND2X1
XFILL_4__2752_ gnd vdd FILL
XFILL_1__2974_ gnd vdd FILL
XFILL_4__1703_ gnd vdd FILL
XFILL_7__2461_ gnd vdd FILL
XFILL_6__3599_ gnd vdd FILL
XFILL_7__2392_ gnd vdd FILL
XFILL_1__1925_ gnd vdd FILL
XFILL_4__2683_ gnd vdd FILL
XFILL_6__2619_ gnd vdd FILL
XFILL_1__1856_ gnd vdd FILL
XFILL_7__3013_ gnd vdd FILL
XFILL_1__1787_ gnd vdd FILL
XFILL_1__3526_ gnd vdd FILL
XFILL_2__2250_ gnd vdd FILL
XFILL_1__3457_ gnd vdd FILL
XFILL_4__3166_ gnd vdd FILL
XFILL_1__2408_ gnd vdd FILL
XFILL_1__3388_ gnd vdd FILL
XFILL_2__2181_ gnd vdd FILL
XFILL_4__3097_ gnd vdd FILL
XFILL_4__2117_ gnd vdd FILL
XFILL_1__2339_ gnd vdd FILL
XFILL_4__2048_ gnd vdd FILL
XFILL_5__2930_ gnd vdd FILL
XFILL_5__2861_ gnd vdd FILL
XFILL_5__2792_ gnd vdd FILL
XFILL_8__2570_ gnd vdd FILL
XFILL_5__1812_ gnd vdd FILL
XFILL_5__1743_ gnd vdd FILL
XFILL_7__2728_ gnd vdd FILL
XFILL_2__1965_ gnd vdd FILL
XFILL_7__2659_ gnd vdd FILL
XFILL_8__3122_ gnd vdd FILL
XFILL_5__3413_ gnd vdd FILL
XFILL_2__1896_ gnd vdd FILL
XFILL_8__3053_ gnd vdd FILL
XFILL_2__3566_ gnd vdd FILL
XFILL_0__2650_ gnd vdd FILL
XFILL_8__2004_ gnd vdd FILL
XFILL_2__2517_ gnd vdd FILL
XFILL_0__2581_ gnd vdd FILL
XFILL_2__3497_ gnd vdd FILL
XFILL_5__2226_ gnd vdd FILL
XFILL_3__2290_ gnd vdd FILL
XFILL_5__2157_ gnd vdd FILL
XFILL_2__2448_ gnd vdd FILL
XFILL_2__2379_ gnd vdd FILL
XFILL_0__3202_ gnd vdd FILL
XFILL_8__2906_ gnd vdd FILL
XFILL_6__2970_ gnd vdd FILL
XFILL_5__2088_ gnd vdd FILL
XFILL_8__2837_ gnd vdd FILL
XFILL_0__3133_ gnd vdd FILL
XFILL_6__1921_ gnd vdd FILL
XFILL_0__3064_ gnd vdd FILL
X_2712_ _3249_/Q _2778_/A _2723_/C vdd gnd NAND2X1
XFILL_6__1852_ gnd vdd FILL
XFILL_0__2015_ gnd vdd FILL
XFILL_8__2768_ gnd vdd FILL
XFILL_8__1719_ gnd vdd FILL
XFILL_6__1783_ gnd vdd FILL
XFILL_8__2699_ gnd vdd FILL
X_2643_ _3352_/Q _2644_/A vdd gnd INVX1
XFILL_6__3522_ gnd vdd FILL
X_2574_ _2773_/A _2574_/B _2574_/C _3586_/A vdd gnd OAI21X1
XFILL_6__3453_ gnd vdd FILL
XFILL_0__2917_ gnd vdd FILL
XFILL_6__3384_ gnd vdd FILL
XFILL_6__2404_ gnd vdd FILL
XFILL_1__1710_ gnd vdd FILL
XFILL_6__2335_ gnd vdd FILL
XFILL_1__2690_ gnd vdd FILL
XFILL_3__2626_ gnd vdd FILL
XFILL_0__2848_ gnd vdd FILL
XFILL_3__2557_ gnd vdd FILL
XFILL_6__2266_ gnd vdd FILL
X_3126_ _3143_/A _3126_/B _3126_/C _3338_/D vdd gnd OAI21X1
XFILL_0__2779_ gnd vdd FILL
XFILL_6__2197_ gnd vdd FILL
XFILL_3__2488_ gnd vdd FILL
X_3057_ _3057_/A _3573_/Q _3059_/A vdd gnd XNOR2X1
XFILL_4__3020_ gnd vdd FILL
X_2008_ _2008_/A _2623_/B _2406_/D vdd gnd NAND2X1
XFILL_3__3109_ gnd vdd FILL
XFILL_7__1961_ gnd vdd FILL
XFILL_1__3173_ gnd vdd FILL
XFILL_1__2124_ gnd vdd FILL
XFILL_7__1892_ gnd vdd FILL
XFILL_1__2055_ gnd vdd FILL
XFILL_4__2804_ gnd vdd FILL
XFILL_7__3562_ gnd vdd FILL
XFILL_7__3493_ gnd vdd FILL
XFILL_7__2513_ gnd vdd FILL
XFILL_4__2735_ gnd vdd FILL
XFILL_7__2444_ gnd vdd FILL
XFILL_1__2957_ gnd vdd FILL
XFILL_2__1750_ gnd vdd FILL
XFILL_4__2666_ gnd vdd FILL
XFILL_1__2888_ gnd vdd FILL
XFILL_7__2375_ gnd vdd FILL
XFILL_1__1908_ gnd vdd FILL
XFILL_2__3420_ gnd vdd FILL
XFILL_1__1839_ gnd vdd FILL
XFILL_4__2597_ gnd vdd FILL
XFILL_5__3060_ gnd vdd FILL
XFILL_2__2302_ gnd vdd FILL
XFILL_5__2011_ gnd vdd FILL
XFILL_1__3509_ gnd vdd FILL
XFILL_4__3218_ gnd vdd FILL
XFILL_5_BUFX2_insert2 gnd vdd FILL
XFILL_2__2233_ gnd vdd FILL
XFILL_4__3149_ gnd vdd FILL
XFILL_2__2164_ gnd vdd FILL
XFILL_5__2913_ gnd vdd FILL
XFILL_4_BUFX2_insert18 gnd vdd FILL
XFILL_2__2095_ gnd vdd FILL
XFILL_8__2622_ gnd vdd FILL
XFILL_5__2844_ gnd vdd FILL
XFILL_8__2553_ gnd vdd FILL
XFILL_5__2775_ gnd vdd FILL
XFILL_2__2997_ gnd vdd FILL
XFILL_8__2484_ gnd vdd FILL
XFILL_5__1726_ gnd vdd FILL
XFILL_3__1790_ gnd vdd FILL
XFILL_2__1948_ gnd vdd FILL
XFILL_2__1879_ gnd vdd FILL
XFILL_3__3460_ gnd vdd FILL
X_2290_ _2290_/A _2344_/A _2336_/A vdd gnd NAND2X1
XFILL_8__3105_ gnd vdd FILL
XFILL_0__2702_ gnd vdd FILL
XFILL_3__2411_ gnd vdd FILL
XFILL_3__3391_ gnd vdd FILL
XFILL_8__3036_ gnd vdd FILL
XFILL_6__2120_ gnd vdd FILL
XFILL_0__2633_ gnd vdd FILL
XFILL_2__3549_ gnd vdd FILL
XFILL_6__2051_ gnd vdd FILL
XFILL_3__2342_ gnd vdd FILL
XFILL_3__2273_ gnd vdd FILL
XFILL_5__2209_ gnd vdd FILL
XFILL_0__2564_ gnd vdd FILL
XFILL_0__2495_ gnd vdd FILL
XFILL_5__3189_ gnd vdd FILL
XFILL_6__2953_ gnd vdd FILL
XFILL_0__3116_ gnd vdd FILL
XFILL_6__1904_ gnd vdd FILL
XFILL_6__2884_ gnd vdd FILL
XFILL_8_BUFX2_insert6 gnd vdd FILL
XFILL_0__3047_ gnd vdd FILL
XFILL_6__1835_ gnd vdd FILL
XFILL_6__1766_ gnd vdd FILL
X_2626_ _3572_/Q _2670_/B _2626_/C _2638_/B vdd gnd AOI21X1
XFILL_1__2811_ gnd vdd FILL
XFILL_6__3505_ gnd vdd FILL
XFILL_3__1988_ gnd vdd FILL
XFILL_6__1697_ gnd vdd FILL
XFILL_4__2520_ gnd vdd FILL
X_2557_ _3071_/A _2570_/B _2557_/C _2558_/C vdd gnd OAI21X1
XFILL_6__3436_ gnd vdd FILL
X_2488_ _2488_/A _2488_/B _2489_/C vdd gnd AND2X2
XFILL_4__2451_ gnd vdd FILL
XFILL_1__2742_ gnd vdd FILL
XFILL_7__2160_ gnd vdd FILL
XFILL_6__3367_ gnd vdd FILL
XFILL_1__2673_ gnd vdd FILL
XFILL_9__3076_ gnd vdd FILL
XFILL_6__2318_ gnd vdd FILL
XFILL_4__2382_ gnd vdd FILL
XFILL_3__3589_ gnd vdd FILL
XFILL_3__2609_ gnd vdd FILL
XFILL_7__2091_ gnd vdd FILL
X_3109_ _3127_/A _3110_/A _3126_/B vdd gnd NAND2X1
XFILL_6__2249_ gnd vdd FILL
XFILL_4__3003_ gnd vdd FILL
XFILL_1__3225_ gnd vdd FILL
XFILL_9__2929_ gnd vdd FILL
XFILL_7__2993_ gnd vdd FILL
XFILL_1__3156_ gnd vdd FILL
XFILL_7__1944_ gnd vdd FILL
XFILL_7__1875_ gnd vdd FILL
XFILL_1__3087_ gnd vdd FILL
XFILL_1__2107_ gnd vdd FILL
XFILL_2__2920_ gnd vdd FILL
XFILL_1__2038_ gnd vdd FILL
XFILL_7__3545_ gnd vdd FILL
XFILL_2__2851_ gnd vdd FILL
XFILL_5__2560_ gnd vdd FILL
XFILL_7__3476_ gnd vdd FILL
XFILL_4__2718_ gnd vdd FILL
XFILL_2__2782_ gnd vdd FILL
XFILL_2__1802_ gnd vdd FILL
XFILL_7__2427_ gnd vdd FILL
XFILL_5__2491_ gnd vdd FILL
XFILL_2__1733_ gnd vdd FILL
XFILL_7__2358_ gnd vdd FILL
XFILL_4__2649_ gnd vdd FILL
XFILL_5__3112_ gnd vdd FILL
XFILL_2__3403_ gnd vdd FILL
XFILL_7__2289_ gnd vdd FILL
XFILL_5__3043_ gnd vdd FILL
XFILL_2__2216_ gnd vdd FILL
XFILL_0__2280_ gnd vdd FILL
XFILL_8__1984_ gnd vdd FILL
XFILL_2__3196_ gnd vdd FILL
XFILL_2__2147_ gnd vdd FILL
XFILL_2__2078_ gnd vdd FILL
X_1790_ _2292_/B _3161_/B _2340_/A vdd gnd NOR2X1
XFILL_3__2960_ gnd vdd FILL
XFILL_8__2605_ gnd vdd FILL
XFILL_2_CLKBUF1_insert34 gnd vdd FILL
XFILL_3__2891_ gnd vdd FILL
XFILL_5__2827_ gnd vdd FILL
XFILL_3__1911_ gnd vdd FILL
XFILL_8__3585_ gnd vdd FILL
X_3460_ _3521_/A _3460_/B _3473_/A vdd gnd NAND2X1
XFILL_3__1842_ gnd vdd FILL
XFILL_8__2536_ gnd vdd FILL
X_3391_ _3552_/A _3391_/B _3391_/C _3567_/D vdd gnd OAI21X1
XFILL_8__2467_ gnd vdd FILL
XFILL_3__1773_ gnd vdd FILL
XFILL_5__2758_ gnd vdd FILL
X_2411_ _2411_/A _2411_/B _2412_/C vdd gnd AND2X2
XFILL_3__3512_ gnd vdd FILL
XFILL_5__1709_ gnd vdd FILL
X_2342_ _2342_/A _3003_/S _2342_/C _2343_/A vdd gnd OAI21X1
XFILL_0__1995_ gnd vdd FILL
XFILL_5__2689_ gnd vdd FILL
XFILL_8__2398_ gnd vdd FILL
XFILL_6__3221_ gnd vdd FILL
XFILL_3__3443_ gnd vdd FILL
X_2273_ _2273_/A _2273_/B _2273_/C _2281_/C vdd gnd NAND3X1
XFILL_6__3152_ gnd vdd FILL
XFILL_3__3374_ gnd vdd FILL
XFILL_0_BUFX2_insert27 gnd vdd FILL
XFILL_6__2103_ gnd vdd FILL
XFILL_0_BUFX2_insert16 gnd vdd FILL
XFILL_0_BUFX2_insert49 gnd vdd FILL
XFILL_8__3019_ gnd vdd FILL
XFILL_6__3083_ gnd vdd FILL
XFILL_3__2325_ gnd vdd FILL
XFILL_0__3596_ gnd vdd FILL
XFILL_0__2616_ gnd vdd FILL
XFILL_6__2034_ gnd vdd FILL
XFILL_0__2547_ gnd vdd FILL
XFILL_3__2256_ gnd vdd FILL
XFILL_1__3010_ gnd vdd FILL
XFILL_3__2187_ gnd vdd FILL
XFILL_0__2478_ gnd vdd FILL
XFILL_6__2936_ gnd vdd FILL
XFILL_6__2867_ gnd vdd FILL
XFILL_4__1951_ gnd vdd FILL
X_1988_ _2449_/B _1991_/B vdd gnd INVX1
XFILL_9__2576_ gnd vdd FILL
XFILL_4__1882_ gnd vdd FILL
XFILL_6__1818_ gnd vdd FILL
XFILL_6__2798_ gnd vdd FILL
X_3589_ _3589_/A AB[4] vdd gnd BUFX2
XFILL_6__1749_ gnd vdd FILL
X_2609_ _2609_/A _2609_/B _2609_/C _2609_/D _2639_/B vdd gnd AOI22X1
XFILL_4__3552_ gnd vdd FILL
XFILL_4__3483_ gnd vdd FILL
XFILL_6__3419_ gnd vdd FILL
XFILL_4__2503_ gnd vdd FILL
XFILL_7__2212_ gnd vdd FILL
XFILL_1__2725_ gnd vdd FILL
XFILL_7__3192_ gnd vdd FILL
XFILL_4__2434_ gnd vdd FILL
XFILL_7__2143_ gnd vdd FILL
XFILL_4__2365_ gnd vdd FILL
XFILL_1__2656_ gnd vdd FILL
XFILL_7__2074_ gnd vdd FILL
XFILL_1__2587_ gnd vdd FILL
XFILL_4__2296_ gnd vdd FILL
XFILL_2__3050_ gnd vdd FILL
XFILL_2__2001_ gnd vdd FILL
XFILL_7__2976_ gnd vdd FILL
XFILL_1__3208_ gnd vdd FILL
XFILL_1__3139_ gnd vdd FILL
XFILL_7__1927_ gnd vdd FILL
XFILL_5__1991_ gnd vdd FILL
XFILL_7__1858_ gnd vdd FILL
XFILL_2__2903_ gnd vdd FILL
XFILL_8__3370_ gnd vdd FILL
XFILL_5__2612_ gnd vdd FILL
XFILL_7__1789_ gnd vdd FILL
XFILL_2__2834_ gnd vdd FILL
XFILL_7__3528_ gnd vdd FILL
XFILL_8__2321_ gnd vdd FILL
XFILL_5__3592_ gnd vdd FILL
XFILL_7__3459_ gnd vdd FILL
XFILL_8__2252_ gnd vdd FILL
XFILL_5__2543_ gnd vdd FILL
XFILL_5__2474_ gnd vdd FILL
XFILL_2__2765_ gnd vdd FILL
XFILL_8__2183_ gnd vdd FILL
XFILL_0__1780_ gnd vdd FILL
XFILL_2__2696_ gnd vdd FILL
XFILL_2__1716_ gnd vdd FILL
XFILL_7_BUFX2_insert22 gnd vdd FILL
XFILL_7_BUFX2_insert11 gnd vdd FILL
XFILL_0__3450_ gnd vdd FILL
XFILL_7_BUFX2_insert44 gnd vdd FILL
XFILL_7_BUFX2_insert55 gnd vdd FILL
XFILL_0__3381_ gnd vdd FILL
XFILL_0__2401_ gnd vdd FILL
XFILL_7_BUFX2_insert88 gnd vdd FILL
XFILL_7_BUFX2_insert66 gnd vdd FILL
XFILL_7_BUFX2_insert77 gnd vdd FILL
XFILL_3__2110_ gnd vdd FILL
XFILL_3__3090_ gnd vdd FILL
XFILL_5__3026_ gnd vdd FILL
XFILL_0__2332_ gnd vdd FILL
XFILL_3__2041_ gnd vdd FILL
X_2960_ _2960_/A _2960_/B _2981_/A _2991_/B vdd gnd OAI21X1
XFILL_8__1967_ gnd vdd FILL
X_2891_ _2933_/C _2927_/A _2891_/C _2892_/B vdd gnd OAI21X1
XFILL_0__2263_ gnd vdd FILL
X_1911_ _3356_/Q _3217_/A vdd gnd INVX1
XFILL_2__3179_ gnd vdd FILL
XFILL_0__2194_ gnd vdd FILL
X_1842_ _1861_/C _1843_/C vdd gnd INVX1
XFILL_8__1898_ gnd vdd FILL
XFILL_6__2721_ gnd vdd FILL
XFILL_3__2943_ gnd vdd FILL
X_1773_ _3238_/Q _3165_/A _1773_/Y vdd gnd NOR2X1
X_3512_ _3532_/A _3532_/B _3535_/A _3534_/B vdd gnd OAI21X1
XFILL_6__2652_ gnd vdd FILL
X_3443_ _3443_/A _3466_/B _3482_/B vdd gnd XOR2X1
XFILL_3__2874_ gnd vdd FILL
XFILL_6__2583_ gnd vdd FILL
XFILL_8__2519_ gnd vdd FILL
XFILL_8__3499_ gnd vdd FILL
XFILL_3__1825_ gnd vdd FILL
X_3374_ _3566_/A _3374_/Y vdd gnd INVX4
XFILL_3__1756_ gnd vdd FILL
XFILL_0__1978_ gnd vdd FILL
X_2325_ _2325_/A _2325_/B _2326_/C vdd gnd NOR2X1
XFILL_6__3204_ gnd vdd FILL
XFILL_1__3490_ gnd vdd FILL
X_2256_ _2305_/A _2288_/C _2257_/B vdd gnd NOR2X1
XFILL_3__3426_ gnd vdd FILL
XFILL_1__2510_ gnd vdd FILL
XFILL_6__3135_ gnd vdd FILL
XFILL_1__2441_ gnd vdd FILL
XFILL_6__3066_ gnd vdd FILL
X_2187_ _2255_/C _2190_/D vdd gnd INVX1
XFILL_4__2150_ gnd vdd FILL
XFILL_1__2372_ gnd vdd FILL
XFILL_6__2017_ gnd vdd FILL
XFILL_4__2081_ gnd vdd FILL
XFILL_3__2308_ gnd vdd FILL
XFILL_0__3579_ gnd vdd FILL
XFILL_3__2239_ gnd vdd FILL
XFILL_7__2830_ gnd vdd FILL
XFILL_7__2761_ gnd vdd FILL
XFILL_6__2919_ gnd vdd FILL
XFILL_4__2983_ gnd vdd FILL
XFILL_7__1712_ gnd vdd FILL
XFILL_7__2692_ gnd vdd FILL
XFILL_4__1934_ gnd vdd FILL
XFILL181950x35250 gnd vdd FILL
XFILL_4__1865_ gnd vdd FILL
XFILL_4__1796_ gnd vdd FILL
XFILL_4__3535_ gnd vdd FILL
XFILL_2__2550_ gnd vdd FILL
XFILL_4__3466_ gnd vdd FILL
XFILL_2__2481_ gnd vdd FILL
XFILL_1__2708_ gnd vdd FILL
XFILL_7__3175_ gnd vdd FILL
XFILL_4__3397_ gnd vdd FILL
XFILL_5__2190_ gnd vdd FILL
XFILL_4__2417_ gnd vdd FILL
XFILL_7__2126_ gnd vdd FILL
XFILL_4__2348_ gnd vdd FILL
XFILL_1__2639_ gnd vdd FILL
XFILL_4__2279_ gnd vdd FILL
XFILL_0_BUFX2_insert8 gnd vdd FILL
XFILL_7__2057_ gnd vdd FILL
XFILL_8__2870_ gnd vdd FILL
XFILL_2__3102_ gnd vdd FILL
XFILL_2__3033_ gnd vdd FILL
XFILL_8__1821_ gnd vdd FILL
XFILL181950x105450 gnd vdd FILL
XFILL_7__2959_ gnd vdd FILL
XFILL_8__1752_ gnd vdd FILL
XFILL_5__1974_ gnd vdd FILL
XFILL_8__3422_ gnd vdd FILL
XFILL_0__2950_ gnd vdd FILL
XFILL_8__2304_ gnd vdd FILL
XFILL_0__1901_ gnd vdd FILL
XFILL_2__2817_ gnd vdd FILL
XFILL_0__2881_ gnd vdd FILL
XFILL_3__2590_ gnd vdd FILL
XFILL_5__2526_ gnd vdd FILL
XFILL_8__2235_ gnd vdd FILL
XFILL_0__1832_ gnd vdd FILL
XFILL_2__2748_ gnd vdd FILL
X_3090_ _3090_/A _3143_/A _3090_/C _3322_/D vdd gnd OAI21X1
XFILL_8__2166_ gnd vdd FILL
XFILL_5__2457_ gnd vdd FILL
XFILL_0__1763_ gnd vdd FILL
X_2110_ _2294_/A _2357_/A _2110_/C _2111_/B vdd gnd OAI21X1
XFILL_0__3502_ gnd vdd FILL
X_2041_ _2932_/A _2890_/A _2044_/A vdd gnd NAND2X1
XFILL_5__2388_ gnd vdd FILL
XFILL_2__2679_ gnd vdd FILL
XFILL_0__3433_ gnd vdd FILL
XFILL_0__1694_ gnd vdd FILL
XFILL_3__3211_ gnd vdd FILL
XFILL_8__2097_ gnd vdd FILL
XFILL_3__3142_ gnd vdd FILL
XFILL_3__3073_ gnd vdd FILL
XFILL_0__3364_ gnd vdd FILL
XFILL_3__2024_ gnd vdd FILL
XFILL_5__3009_ gnd vdd FILL
X_2943_ reset _2957_/C _3300_/Q _2944_/C vdd gnd OAI21X1
XFILL_0__2315_ gnd vdd FILL
XFILL_8__2999_ gnd vdd FILL
XFILL_0__2246_ gnd vdd FILL
XFILL_9__3531_ gnd vdd FILL
X_2874_ _3309_/Q _2933_/B _2876_/C vdd gnd NAND2X1
X_1825_ _2646_/A _3189_/C _2950_/A _1831_/D _3420_/A vdd gnd OAI22X1
XFILL_0__2177_ gnd vdd FILL
XFILL_3_BUFX2_insert20 gnd vdd FILL
XFILL_1__2990_ gnd vdd FILL
X_1756_ _1756_/A _1762_/B _1803_/B vdd gnd NAND2X1
XFILL_6__2704_ gnd vdd FILL
XFILL_3__2926_ gnd vdd FILL
XFILL_3_BUFX2_insert64 gnd vdd FILL
XFILL_3_BUFX2_insert42 gnd vdd FILL
XFILL_3_BUFX2_insert53 gnd vdd FILL
XFILL_6__2635_ gnd vdd FILL
XFILL_3_BUFX2_insert97 gnd vdd FILL
XFILL_1__1941_ gnd vdd FILL
XFILL_3__2857_ gnd vdd FILL
XFILL_3_BUFX2_insert75 gnd vdd FILL
XFILL_3_BUFX2_insert86 gnd vdd FILL
XFILL_1__1872_ gnd vdd FILL
X_3426_ _3426_/A _3426_/B _3426_/C _3432_/A vdd gnd OAI21X1
XFILL_3__1808_ gnd vdd FILL
XFILL_6__2566_ gnd vdd FILL
XFILL_3__2788_ gnd vdd FILL
XFILL_6__2497_ gnd vdd FILL
X_3357_ _3357_/D vdd _3363_/R _3363_/CLK _3357_/Q vdd gnd DFFSR
XFILL_1__3542_ gnd vdd FILL
X_2308_ _2308_/A _2308_/B _2314_/C vdd gnd NOR2X1
XFILL_3__1739_ gnd vdd FILL
X_3288_ _3288_/D vdd _3289_/R _3307_/CLK _3288_/Q vdd gnd DFFSR
XFILL_6__3118_ gnd vdd FILL
XFILL_1__3473_ gnd vdd FILL
XFILL_3__3409_ gnd vdd FILL
XFILL_4__2202_ gnd vdd FILL
X_2239_ _2276_/A _2781_/B _2278_/A _2240_/C vdd gnd OAI21X1
XFILL_4__3182_ gnd vdd FILL
XFILL_1__2424_ gnd vdd FILL
XFILL_4__2133_ gnd vdd FILL
XFILL_6__3049_ gnd vdd FILL
XFILL_1__2355_ gnd vdd FILL
XFILL_4__2064_ gnd vdd FILL
XFILL_7__2813_ gnd vdd FILL
XFILL_1__2286_ gnd vdd FILL
XFILL_7__2744_ gnd vdd FILL
XFILL_4__2966_ gnd vdd FILL
XFILL_7__2675_ gnd vdd FILL
XFILL_4__1917_ gnd vdd FILL
XFILL_4__2897_ gnd vdd FILL
XFILL_5__1690_ gnd vdd FILL
XFILL_2__1981_ gnd vdd FILL
XFILL_4__1848_ gnd vdd FILL
XFILL_2__2602_ gnd vdd FILL
XFILL_4__1779_ gnd vdd FILL
XFILL_8__2020_ gnd vdd FILL
XFILL_4__3518_ gnd vdd FILL
XFILL_5__2311_ gnd vdd FILL
XFILL_2__3582_ gnd vdd FILL
XFILL_7__3227_ gnd vdd FILL
XFILL_4__3449_ gnd vdd FILL
XFILL_5__2242_ gnd vdd FILL
XFILL_2__2533_ gnd vdd FILL
XFILL_5__2173_ gnd vdd FILL
XFILL_2__2464_ gnd vdd FILL
XFILL_7__3158_ gnd vdd FILL
XFILL_7__3089_ gnd vdd FILL
XFILL_2__2395_ gnd vdd FILL
XFILL_7__2109_ gnd vdd FILL
XFILL_8__2922_ gnd vdd FILL
XFILL181950x117150 gnd vdd FILL
XFILL_7_CLKBUF1_insert34 gnd vdd FILL
XFILL_8__2853_ gnd vdd FILL
XFILL_0__2100_ gnd vdd FILL
XFILL_8__2784_ gnd vdd FILL
XFILL_0__3080_ gnd vdd FILL
XFILL_2__3016_ gnd vdd FILL
XFILL_8__1804_ gnd vdd FILL
XFILL183150x101550 gnd vdd FILL
XFILL_0__2031_ gnd vdd FILL
XFILL_8__1735_ gnd vdd FILL
XFILL_5__1957_ gnd vdd FILL
XFILL_8__3405_ gnd vdd FILL
X_2590_ _2700_/B _2699_/B _2726_/C _2670_/B vdd gnd NAND3X1
XFILL_6__2420_ gnd vdd FILL
XFILL_5__1888_ gnd vdd FILL
XFILL_3__2711_ gnd vdd FILL
XFILL_0__2933_ gnd vdd FILL
XFILL_3__2642_ gnd vdd FILL
XFILL_5__3558_ gnd vdd FILL
XFILL_0__2864_ gnd vdd FILL
XFILL_6__2351_ gnd vdd FILL
X_3211_ _3215_/A _3211_/B _3211_/C _3353_/D vdd gnd OAI21X1
X_3142_ _3347_/Q _3143_/B _3143_/C vdd gnd NAND2X1
XFILL_5__3489_ gnd vdd FILL
XFILL_6__2282_ gnd vdd FILL
XFILL_8__2218_ gnd vdd FILL
XFILL_5__2509_ gnd vdd FILL
XFILL_3__2573_ gnd vdd FILL
XFILL_0__1815_ gnd vdd FILL
XFILL_0__2795_ gnd vdd FILL
XFILL_8__3198_ gnd vdd FILL
X_3073_ _3295_/D _3077_/C _3073_/C _3073_/D _3139_/A vdd gnd AOI22X1
XFILL_8__2149_ gnd vdd FILL
XFILL_0__1746_ gnd vdd FILL
X_2024_ _2025_/A _3305_/Q _2025_/C vdd gnd NAND2X1
XFILL_0__3416_ gnd vdd FILL
XFILL_9__1913_ gnd vdd FILL
XFILL_3__3125_ gnd vdd FILL
XFILL_1__2140_ gnd vdd FILL
XFILL_3__3056_ gnd vdd FILL
X_2926_ _2928_/B _2926_/B _2926_/C _2929_/B vdd gnd OAI21X1
XFILL_1__2071_ gnd vdd FILL
XFILL_3__2007_ gnd vdd FILL
XBUFX2_insert18 _2580_/Y _3346_/R vdd gnd BUFX2
X_2857_ _2857_/A _2916_/C _2857_/C _2858_/B vdd gnd OAI21X1
XFILL_6__1997_ gnd vdd FILL
XFILL_0__2229_ gnd vdd FILL
XFILL_4__2820_ gnd vdd FILL
X_1808_ _2594_/A _2123_/A vdd gnd INVX1
X_2788_ _2814_/A _2899_/A _2788_/C _3258_/D vdd gnd OAI21X1
XFILL_4__2751_ gnd vdd FILL
XFILL_3__2909_ gnd vdd FILL
XFILL_1__2973_ gnd vdd FILL
XFILL_4__1702_ gnd vdd FILL
XFILL_7__2460_ gnd vdd FILL
X_1739_ _3236_/Q _1739_/B _2442_/B vdd gnd NAND2X1
XFILL_6__3598_ gnd vdd FILL
XFILL_7__2391_ gnd vdd FILL
XFILL_4__2682_ gnd vdd FILL
XFILL_6__2618_ gnd vdd FILL
XFILL_1__1924_ gnd vdd FILL
X_3409_ _3409_/A _3409_/B _3409_/C _3511_/A vdd gnd OAI21X1
XFILL_6__2549_ gnd vdd FILL
XFILL_1__1855_ gnd vdd FILL
XFILL_7__3012_ gnd vdd FILL
XFILL_1__1786_ gnd vdd FILL
XFILL_1__3525_ gnd vdd FILL
XFILL_1__3456_ gnd vdd FILL
XFILL_4__3165_ gnd vdd FILL
XFILL_1__2407_ gnd vdd FILL
XFILL_2__2180_ gnd vdd FILL
XFILL_4__3096_ gnd vdd FILL
XFILL_1__3387_ gnd vdd FILL
XFILL_4__2116_ gnd vdd FILL
XFILL_1__2338_ gnd vdd FILL
XFILL_4__2047_ gnd vdd FILL
XFILL_1__2269_ gnd vdd FILL
XFILL_5__2860_ gnd vdd FILL
XFILL_5__2791_ gnd vdd FILL
XFILL_7__2727_ gnd vdd FILL
XFILL_5__1811_ gnd vdd FILL
XFILL_4__2949_ gnd vdd FILL
XFILL_5__1742_ gnd vdd FILL
XFILL_2__1964_ gnd vdd FILL
XFILL_7__2658_ gnd vdd FILL
XFILL_7__2589_ gnd vdd FILL
XFILL_8__3121_ gnd vdd FILL
XFILL_5__3412_ gnd vdd FILL
XFILL_2__1895_ gnd vdd FILL
XFILL_8__3052_ gnd vdd FILL
XFILL_2__3565_ gnd vdd FILL
XFILL_0__2580_ gnd vdd FILL
XFILL_8__2003_ gnd vdd FILL
XFILL_2__2516_ gnd vdd FILL
XFILL_2__3496_ gnd vdd FILL
XFILL_5__2225_ gnd vdd FILL
XFILL_5__2156_ gnd vdd FILL
XFILL_2__2447_ gnd vdd FILL
XFILL183450x105450 gnd vdd FILL
XFILL_2__2378_ gnd vdd FILL
XFILL_0__3201_ gnd vdd FILL
XFILL_8__2905_ gnd vdd FILL
XFILL_5__2087_ gnd vdd FILL
XFILL_8__2836_ gnd vdd FILL
XFILL_0__3132_ gnd vdd FILL
XFILL_6__1920_ gnd vdd FILL
XFILL_6__1851_ gnd vdd FILL
X_2711_ _2767_/A _2711_/B _2711_/C _2711_/D _3248_/D vdd gnd OAI22X1
XFILL_0__3063_ gnd vdd FILL
XFILL_0__2014_ gnd vdd FILL
XFILL_8__2767_ gnd vdd FILL
XFILL_5__2989_ gnd vdd FILL
XFILL_6__3521_ gnd vdd FILL
X_2642_ _3243_/Q _2768_/A _2648_/C vdd gnd NAND2X1
XFILL_8__1718_ gnd vdd FILL
XFILL_8__2698_ gnd vdd FILL
XFILL_6__1782_ gnd vdd FILL
X_2573_ _2573_/A _2574_/C vdd gnd INVX1
XFILL_6__3452_ gnd vdd FILL
XFILL_0__2916_ gnd vdd FILL
XFILL_6__3383_ gnd vdd FILL
XFILL_6__2403_ gnd vdd FILL
XFILL_6__2334_ gnd vdd FILL
XFILL_3__2625_ gnd vdd FILL
XFILL_0__2847_ gnd vdd FILL
XFILL_3__2556_ gnd vdd FILL
X_3125_ _3125_/A _3125_/B _3338_/Q _3126_/C vdd gnd OAI21X1
XFILL_6__2265_ gnd vdd FILL
XFILL_0__2778_ gnd vdd FILL
X_3056_ _3056_/A _3056_/B _3056_/C _3059_/B vdd gnd OAI21X1
XFILL_6__2196_ gnd vdd FILL
XFILL_3__2487_ gnd vdd FILL
XFILL_0__1729_ gnd vdd FILL
X_2007_ _3310_/Q _2009_/A vdd gnd INVX1
XFILL_6_BUFX2_insert90 gnd vdd FILL
XFILL_3__3108_ gnd vdd FILL
XFILL_7__1960_ gnd vdd FILL
XFILL_1__3172_ gnd vdd FILL
XFILL_7__1891_ gnd vdd FILL
XFILL_1__2123_ gnd vdd FILL
XFILL_3__3039_ gnd vdd FILL
XFILL_1__2054_ gnd vdd FILL
X_2909_ _2915_/C _2933_/A _2909_/C _2922_/B vdd gnd NAND3X1
XFILL_4__2803_ gnd vdd FILL
XFILL_7__3561_ gnd vdd FILL
XFILL_7__3492_ gnd vdd FILL
XFILL_9__3428_ gnd vdd FILL
XFILL_7__2512_ gnd vdd FILL
XFILL_4__2734_ gnd vdd FILL
XFILL_7__2443_ gnd vdd FILL
XFILL_1__2956_ gnd vdd FILL
XFILL_4__2665_ gnd vdd FILL
XFILL_1__2887_ gnd vdd FILL
XFILL_7__2374_ gnd vdd FILL
XFILL_1__1907_ gnd vdd FILL
XFILL_1__1838_ gnd vdd FILL
XFILL_4__2596_ gnd vdd FILL
XFILL_1__3508_ gnd vdd FILL
XFILL_2__2301_ gnd vdd FILL
XFILL_1__1769_ gnd vdd FILL
XFILL_5__2010_ gnd vdd FILL
XFILL_4__3217_ gnd vdd FILL
XFILL_5_BUFX2_insert3 gnd vdd FILL
XFILL_1__3439_ gnd vdd FILL
XFILL_4__3148_ gnd vdd FILL
XFILL_2__2232_ gnd vdd FILL
XFILL_2__2163_ gnd vdd FILL
XFILL_4__3079_ gnd vdd FILL
XFILL_5__2912_ gnd vdd FILL
XFILL_8__2621_ gnd vdd FILL
XFILL_2__2094_ gnd vdd FILL
XFILL_4_BUFX2_insert19 gnd vdd FILL
XFILL_5__2843_ gnd vdd FILL
XFILL_8__2552_ gnd vdd FILL
XFILL_8__2483_ gnd vdd FILL
XFILL_5__2774_ gnd vdd FILL
XFILL_2__2996_ gnd vdd FILL
XFILL_5__1725_ gnd vdd FILL
XFILL_2__1947_ gnd vdd FILL
XFILL_2__1878_ gnd vdd FILL
XFILL_8__3104_ gnd vdd FILL
XFILL_0__2701_ gnd vdd FILL
XFILL_3__2410_ gnd vdd FILL
XFILL_3__3390_ gnd vdd FILL
XFILL_8__3035_ gnd vdd FILL
XFILL183750x109350 gnd vdd FILL
XFILL_0__2632_ gnd vdd FILL
XFILL_2__3548_ gnd vdd FILL
XFILL183450x117150 gnd vdd FILL
XFILL_3__2341_ gnd vdd FILL
XFILL_6__2050_ gnd vdd FILL
XFILL_2__3479_ gnd vdd FILL
XFILL_3__2272_ gnd vdd FILL
XFILL_5__2208_ gnd vdd FILL
XFILL_0__2563_ gnd vdd FILL
XFILL_0__2494_ gnd vdd FILL
XFILL_5__3188_ gnd vdd FILL
XFILL_5__2139_ gnd vdd FILL
XFILL_6__2952_ gnd vdd FILL
XFILL_0__3115_ gnd vdd FILL
XFILL_6__1903_ gnd vdd FILL
XFILL_8__2819_ gnd vdd FILL
XFILL_6__2883_ gnd vdd FILL
XFILL_8_BUFX2_insert7 gnd vdd FILL
XFILL_0__3046_ gnd vdd FILL
XFILL_6__1834_ gnd vdd FILL
XFILL_6__1765_ gnd vdd FILL
X_2625_ _2728_/A _2625_/B _2625_/C _2626_/C vdd gnd OAI21X1
XFILL_6__3504_ gnd vdd FILL
XFILL_1__2810_ gnd vdd FILL
XFILL_3__1987_ gnd vdd FILL
XFILL_6__3435_ gnd vdd FILL
XFILL_6__1696_ gnd vdd FILL
X_2556_ _2569_/A _2569_/B _3295_/D _2557_/C vdd gnd OAI21X1
X_2487_ _3294_/D _2502_/B _2502_/C _3352_/Q _2488_/B vdd gnd AOI22X1
XFILL_4__2450_ gnd vdd FILL
XFILL_1__2741_ gnd vdd FILL
XFILL_6__3366_ gnd vdd FILL
XFILL_1__2672_ gnd vdd FILL
XFILL_3__2608_ gnd vdd FILL
XFILL_6__2317_ gnd vdd FILL
XFILL_4__2381_ gnd vdd FILL
XFILL_7__2090_ gnd vdd FILL
XFILL_3__3588_ gnd vdd FILL
X_3108_ _3143_/A _3108_/B _3108_/C _3330_/D vdd gnd OAI21X1
XFILL_6__2248_ gnd vdd FILL
XFILL_3__2539_ gnd vdd FILL
XFILL_6__2179_ gnd vdd FILL
X_3039_ _3039_/A _3057_/A _3571_/Q _3050_/B vdd gnd OAI21X1
XFILL_4__3002_ gnd vdd FILL
XFILL_7__2992_ gnd vdd FILL
XFILL_1__3224_ gnd vdd FILL
XFILL_7__1943_ gnd vdd FILL
XFILL_1__3155_ gnd vdd FILL
XFILL_7__1874_ gnd vdd FILL
XFILL_1__3086_ gnd vdd FILL
XFILL_1__2106_ gnd vdd FILL
XFILL_1__2037_ gnd vdd FILL
XFILL_7__3544_ gnd vdd FILL
XFILL_2__2850_ gnd vdd FILL
XFILL_7__3475_ gnd vdd FILL
XFILL_2__2781_ gnd vdd FILL
XFILL_2__1801_ gnd vdd FILL
XFILL_4__2717_ gnd vdd FILL
XFILL_1__2939_ gnd vdd FILL
XFILL_7__2426_ gnd vdd FILL
XFILL_5__2490_ gnd vdd FILL
XFILL_2__1732_ gnd vdd FILL
XFILL_4__2648_ gnd vdd FILL
XFILL_7__2357_ gnd vdd FILL
XFILL_4__2579_ gnd vdd FILL
XFILL_2__3402_ gnd vdd FILL
XFILL_5__3111_ gnd vdd FILL
XFILL_7__2288_ gnd vdd FILL
XFILL_5__3042_ gnd vdd FILL
XFILL_2__2215_ gnd vdd FILL
XFILL_2__3195_ gnd vdd FILL
XFILL_8__1983_ gnd vdd FILL
XFILL_2__2146_ gnd vdd FILL
XFILL_2__2077_ gnd vdd FILL
XFILL_8__3584_ gnd vdd FILL
XFILL_8__2604_ gnd vdd FILL
XFILL_3__1910_ gnd vdd FILL
XFILL_3__2890_ gnd vdd FILL
XFILL_5__2826_ gnd vdd FILL
XFILL_8__2535_ gnd vdd FILL
XFILL_2_CLKBUF1_insert35 gnd vdd FILL
XFILL_5__2757_ gnd vdd FILL
XFILL_3__1841_ gnd vdd FILL
X_2410_ _2413_/A _3574_/Q _3251_/Q _2413_/D _2411_/B vdd gnd AOI22X1
X_3390_ _3567_/Q _3552_/A _3391_/C vdd gnd NAND2X1
XFILL_2__2979_ gnd vdd FILL
XFILL_3__1772_ gnd vdd FILL
XFILL_5__1708_ gnd vdd FILL
XFILL_8__2466_ gnd vdd FILL
XFILL_3__3511_ gnd vdd FILL
XFILL_0__1994_ gnd vdd FILL
XFILL_8__2397_ gnd vdd FILL
X_2341_ _2341_/A _2341_/B _2341_/C _2343_/B vdd gnd OAI21X1
XFILL_5__2688_ gnd vdd FILL
X_2272_ _2272_/A _2273_/B vdd gnd INVX1
XFILL_6__3220_ gnd vdd FILL
XFILL_3__3442_ gnd vdd FILL
XFILL_6__3151_ gnd vdd FILL
XFILL_3__3373_ gnd vdd FILL
XFILL_0_BUFX2_insert17 gnd vdd FILL
XFILL_0_BUFX2_insert39 gnd vdd FILL
XFILL_6__2102_ gnd vdd FILL
XFILL_6__3082_ gnd vdd FILL
XFILL_8__3018_ gnd vdd FILL
XFILL_3__2324_ gnd vdd FILL
XFILL_0__3595_ gnd vdd FILL
XFILL_0__2615_ gnd vdd FILL
XFILL_6__2033_ gnd vdd FILL
XFILL_0__2546_ gnd vdd FILL
XFILL_3__2255_ gnd vdd FILL
XFILL_3__2186_ gnd vdd FILL
XFILL_0__2477_ gnd vdd FILL
XFILL_6__2935_ gnd vdd FILL
X_1987_ _1987_/A _3160_/C _2449_/B vdd gnd NAND2X1
XFILL_6__2866_ gnd vdd FILL
XFILL_4__1950_ gnd vdd FILL
XFILL_0__3029_ gnd vdd FILL
XFILL_4__1881_ gnd vdd FILL
XFILL_6__1817_ gnd vdd FILL
XFILL_6__2797_ gnd vdd FILL
XFILL_4__3551_ gnd vdd FILL
X_3588_ _3588_/A AB[3] vdd gnd BUFX2
XFILL_6__1748_ gnd vdd FILL
X_2608_ _3348_/Q _2770_/C _2670_/B _3570_/Q _2609_/D vdd gnd AOI22X1
XFILL_4__2502_ gnd vdd FILL
X_2539_ _3359_/Q _2691_/A _2563_/A _3573_/Q _2540_/A vdd gnd AOI22X1
XFILL_4__3482_ gnd vdd FILL
XFILL_6__3418_ gnd vdd FILL
XFILL_7__2211_ gnd vdd FILL
XFILL_1__2724_ gnd vdd FILL
XFILL_7__3191_ gnd vdd FILL
XFILL_7__2142_ gnd vdd FILL
XFILL_4__2433_ gnd vdd FILL
XFILL_4__2364_ gnd vdd FILL
XFILL_1__2655_ gnd vdd FILL
XFILL_7__2073_ gnd vdd FILL
XFILL_1__2586_ gnd vdd FILL
XFILL_4__2295_ gnd vdd FILL
XFILL_2__2000_ gnd vdd FILL
XFILL_7__2975_ gnd vdd FILL
XFILL_1__3207_ gnd vdd FILL
XFILL_1__3138_ gnd vdd FILL
XFILL_7__1926_ gnd vdd FILL
XFILL_5__1990_ gnd vdd FILL
XFILL_7__1857_ gnd vdd FILL
XFILL_1__3069_ gnd vdd FILL
XFILL_2__2902_ gnd vdd FILL
XFILL_5__2611_ gnd vdd FILL
XFILL_7__1788_ gnd vdd FILL
XFILL_7__3527_ gnd vdd FILL
XFILL_2__2833_ gnd vdd FILL
XFILL_5__3591_ gnd vdd FILL
XFILL_8__2320_ gnd vdd FILL
XFILL_7__3458_ gnd vdd FILL
XFILL_8__2251_ gnd vdd FILL
XFILL_5__2542_ gnd vdd FILL
XFILL_5__2473_ gnd vdd FILL
XFILL_2__2764_ gnd vdd FILL
XFILL_7__2409_ gnd vdd FILL
XFILL_7__3389_ gnd vdd FILL
XFILL_8__2182_ gnd vdd FILL
XFILL_2__2695_ gnd vdd FILL
XFILL_2__1715_ gnd vdd FILL
XFILL_7_BUFX2_insert12 gnd vdd FILL
XFILL_7_BUFX2_insert23 gnd vdd FILL
XFILL_7_BUFX2_insert56 gnd vdd FILL
XFILL_7_BUFX2_insert45 gnd vdd FILL
XFILL_0__3380_ gnd vdd FILL
XFILL_7_BUFX2_insert78 gnd vdd FILL
XFILL_0__2400_ gnd vdd FILL
XFILL_7_BUFX2_insert67 gnd vdd FILL
XFILL_7_BUFX2_insert89 gnd vdd FILL
XFILL_0__2331_ gnd vdd FILL
XFILL_5__3025_ gnd vdd FILL
XFILL_3__2040_ gnd vdd FILL
XFILL_8__1966_ gnd vdd FILL
X_2890_ _2890_/A _2930_/A _2927_/A vdd gnd NOR2X1
XFILL_0__2262_ gnd vdd FILL
XFILL_2__3178_ gnd vdd FILL
X_1910_ _3158_/A _1910_/B _1910_/C _1985_/A vdd gnd NAND3X1
XFILL_0__2193_ gnd vdd FILL
XFILL_2__2129_ gnd vdd FILL
X_1841_ _1841_/A _1841_/B _1861_/C vdd gnd NAND2X1
XFILL_8__1897_ gnd vdd FILL
XFILL_6__2720_ gnd vdd FILL
XFILL_3__2942_ gnd vdd FILL
X_1772_ _3313_/Q _2865_/A _1772_/C _1777_/C vdd gnd OAI21X1
XFILL_6__2651_ gnd vdd FILL
X_3511_ _3511_/A _3511_/B _3535_/A _3532_/A vdd gnd OAI21X1
XFILL_5__2809_ gnd vdd FILL
XFILL_3__2873_ gnd vdd FILL
XFILL_8__3498_ gnd vdd FILL
X_3442_ _3442_/A _3442_/B _3443_/A vdd gnd NOR2X1
XFILL_3__1824_ gnd vdd FILL
XFILL_8__2518_ gnd vdd FILL
XFILL_6__2582_ gnd vdd FILL
X_3373_ reset _3578_/R vdd gnd INVX4
XFILL_8__2449_ gnd vdd FILL
XFILL_3__1755_ gnd vdd FILL
X_2324_ _2324_/A _2324_/B _2324_/C _2325_/B vdd gnd NAND3X1
XFILL_0__1977_ gnd vdd FILL
XFILL_6__3203_ gnd vdd FILL
X_2255_ _2270_/A _2881_/A _2255_/C _2310_/B vdd gnd OAI21X1
XFILL_3__3425_ gnd vdd FILL
XFILL_6__3134_ gnd vdd FILL
X_2186_ _2910_/B _2928_/A _2255_/C vdd gnd NOR2X1
XFILL_1__2440_ gnd vdd FILL
XFILL_6__3065_ gnd vdd FILL
XFILL_1__2371_ gnd vdd FILL
XFILL_4__2080_ gnd vdd FILL
XFILL_6__2016_ gnd vdd FILL
XFILL_3__2307_ gnd vdd FILL
XFILL_3__2238_ gnd vdd FILL
XFILL_0__2529_ gnd vdd FILL
XFILL_3__2169_ gnd vdd FILL
XFILL_7__2760_ gnd vdd FILL
XFILL_6__2918_ gnd vdd FILL
XFILL_4__2982_ gnd vdd FILL
XFILL_7__1711_ gnd vdd FILL
XFILL_7__2691_ gnd vdd FILL
XFILL_4__1933_ gnd vdd FILL
XFILL_6__2849_ gnd vdd FILL
XFILL_4__1864_ gnd vdd FILL
XFILL_4__3603_ gnd vdd FILL
XFILL_4__1795_ gnd vdd FILL
XFILL_4__3534_ gnd vdd FILL
XFILL_4__3465_ gnd vdd FILL
XFILL_4__2416_ gnd vdd FILL
XFILL_1__2707_ gnd vdd FILL
XFILL_7__3174_ gnd vdd FILL
XFILL_2__2480_ gnd vdd FILL
XFILL_4__3396_ gnd vdd FILL
XFILL_7__2125_ gnd vdd FILL
XFILL_1__2638_ gnd vdd FILL
XFILL_4__2347_ gnd vdd FILL
XFILL_7__2056_ gnd vdd FILL
XFILL_4__2278_ gnd vdd FILL
XFILL_0_BUFX2_insert9 gnd vdd FILL
XFILL_1__2569_ gnd vdd FILL
XFILL_2__3101_ gnd vdd FILL
XFILL_2__3032_ gnd vdd FILL
XFILL_8__1820_ gnd vdd FILL
XFILL_8__1751_ gnd vdd FILL
XFILL_5__1973_ gnd vdd FILL
XFILL_7__2958_ gnd vdd FILL
XFILL_7__2889_ gnd vdd FILL
XFILL_7__1909_ gnd vdd FILL
XFILL_8__3421_ gnd vdd FILL
XFILL_8__2303_ gnd vdd FILL
XFILL_0__1900_ gnd vdd FILL
XFILL_0__2880_ gnd vdd FILL
XFILL_2__2816_ gnd vdd FILL
XFILL_5__2525_ gnd vdd FILL
XFILL_0__1831_ gnd vdd FILL
XFILL_8__2234_ gnd vdd FILL
XFILL_2__2747_ gnd vdd FILL
XFILL_8__2165_ gnd vdd FILL
XFILL_5__2456_ gnd vdd FILL
XFILL_0__1762_ gnd vdd FILL
X_2040_ _2933_/C _2931_/A _2896_/C vdd gnd NAND2X1
XFILL_0__3501_ gnd vdd FILL
XFILL_5__2387_ gnd vdd FILL
XFILL_3__3210_ gnd vdd FILL
XFILL_2__2678_ gnd vdd FILL
XFILL_0__3432_ gnd vdd FILL
XFILL_8__2096_ gnd vdd FILL
XFILL_0__1693_ gnd vdd FILL
XFILL_3__3141_ gnd vdd FILL
XFILL_5__3008_ gnd vdd FILL
XFILL_3__3072_ gnd vdd FILL
XFILL_3__2023_ gnd vdd FILL
X_2942_ _3016_/A _2956_/B _2942_/C _3299_/D vdd gnd OAI21X1
XFILL_0__2314_ gnd vdd FILL
XFILL_8__2998_ gnd vdd FILL
XFILL_0__2245_ gnd vdd FILL
XFILL_8__1949_ gnd vdd FILL
X_2873_ _2873_/A _2878_/B vdd gnd INVX1
XFILL_0__2176_ gnd vdd FILL
X_1824_ _3243_/Q _2646_/A vdd gnd INVX1
XFILL_6__2703_ gnd vdd FILL
XFILL_3__2925_ gnd vdd FILL
X_1755_ _3274_/Q _2865_/A vdd gnd INVX1
XFILL_3_BUFX2_insert21 gnd vdd FILL
XFILL_3_BUFX2_insert10 gnd vdd FILL
XFILL_1__1940_ gnd vdd FILL
XFILL_3_BUFX2_insert43 gnd vdd FILL
XFILL_3_BUFX2_insert65 gnd vdd FILL
XFILL_3_BUFX2_insert54 gnd vdd FILL
XFILL_6__2634_ gnd vdd FILL
XFILL_3__2856_ gnd vdd FILL
XFILL_3_BUFX2_insert87 gnd vdd FILL
XFILL_6__2565_ gnd vdd FILL
XFILL_3_BUFX2_insert76 gnd vdd FILL
XFILL_1__1871_ gnd vdd FILL
XFILL184650x171750 gnd vdd FILL
X_3425_ _3434_/A _3425_/B _3459_/A _3426_/A vdd gnd OAI21X1
XFILL_3__2787_ gnd vdd FILL
XFILL_3__1807_ gnd vdd FILL
XFILL_6__2496_ gnd vdd FILL
X_3356_ _3356_/D vdd _3363_/R _3363_/CLK _3356_/Q vdd gnd DFFSR
XFILL_3__1738_ gnd vdd FILL
X_3287_ _3287_/D vdd _3346_/R _3307_/CLK _3287_/Q vdd gnd DFFSR
X_2307_ _2307_/A _2307_/B _2308_/A vdd gnd NAND2X1
XFILL_1__3541_ gnd vdd FILL
X_2238_ _2242_/C _2238_/B _2245_/B vdd gnd NAND2X1
XFILL_6__3117_ gnd vdd FILL
XFILL_1__3472_ gnd vdd FILL
XFILL_3__3408_ gnd vdd FILL
XFILL_4__2201_ gnd vdd FILL
XFILL_4__3181_ gnd vdd FILL
X_2169_ _2910_/B _2899_/A _2875_/A vdd gnd NOR2X1
XFILL_1__2423_ gnd vdd FILL
XFILL_4__2132_ gnd vdd FILL
XFILL_1__2354_ gnd vdd FILL
XFILL_6__3048_ gnd vdd FILL
XFILL_4__2063_ gnd vdd FILL
XFILL_7__2812_ gnd vdd FILL
XFILL_1__2285_ gnd vdd FILL
XFILL_7__2743_ gnd vdd FILL
XFILL_4__2965_ gnd vdd FILL
XFILL_7__2674_ gnd vdd FILL
XFILL_4__2896_ gnd vdd FILL
XFILL_4__1916_ gnd vdd FILL
XFILL_2__1980_ gnd vdd FILL
XFILL_4__1847_ gnd vdd FILL
XFILL_4__3517_ gnd vdd FILL
XFILL_5__2310_ gnd vdd FILL
XFILL_4__1778_ gnd vdd FILL
XFILL_2__3581_ gnd vdd FILL
XFILL_2__2601_ gnd vdd FILL
XFILL_2__2532_ gnd vdd FILL
XFILL_7__3226_ gnd vdd FILL
XFILL_4__3448_ gnd vdd FILL
XFILL_5__2241_ gnd vdd FILL
XFILL_7__3157_ gnd vdd FILL
XFILL_4__3379_ gnd vdd FILL
XFILL_5__2172_ gnd vdd FILL
XFILL_2__2463_ gnd vdd FILL
XFILL_7__2108_ gnd vdd FILL
XFILL_7__3088_ gnd vdd FILL
XFILL_2__2394_ gnd vdd FILL
XFILL_8__2921_ gnd vdd FILL
XFILL_7__2039_ gnd vdd FILL
XFILL_7_CLKBUF1_insert35 gnd vdd FILL
XFILL_8__2852_ gnd vdd FILL
XFILL_2__3015_ gnd vdd FILL
XFILL_8__2783_ gnd vdd FILL
XFILL_8__1803_ gnd vdd FILL
XFILL_0__2030_ gnd vdd FILL
XFILL_8__1734_ gnd vdd FILL
XFILL_5__1956_ gnd vdd FILL
XFILL_8__3404_ gnd vdd FILL
XFILL_5__1887_ gnd vdd FILL
XFILL_3__2710_ gnd vdd FILL
XFILL_0__2932_ gnd vdd FILL
XFILL_3__2641_ gnd vdd FILL
XFILL_0__2863_ gnd vdd FILL
XFILL_5__3557_ gnd vdd FILL
XFILL_6__2350_ gnd vdd FILL
X_3210_ _3214_/A _3214_/B _3353_/Q _3211_/C vdd gnd OAI21X1
X_3141_ _3141_/A _3143_/B _3141_/C _3346_/D vdd gnd OAI21X1
XFILL_5__3488_ gnd vdd FILL
XFILL_8__2217_ gnd vdd FILL
XFILL_6__2281_ gnd vdd FILL
XFILL_3__2572_ gnd vdd FILL
XFILL_0__1814_ gnd vdd FILL
XFILL_5__2508_ gnd vdd FILL
XFILL_0__2794_ gnd vdd FILL
XFILL_8__3197_ gnd vdd FILL
XFILL_5__2439_ gnd vdd FILL
X_3072_ _3077_/C _3083_/B _3073_/C vdd gnd NOR2X1
XFILL_8__2148_ gnd vdd FILL
XFILL_0__1745_ gnd vdd FILL
XFILL_8__2079_ gnd vdd FILL
X_2023_ _2889_/C _2161_/A _2933_/B vdd gnd NAND2X1
XFILL_3__3124_ gnd vdd FILL
XFILL_0__3415_ gnd vdd FILL
XFILL_3__3055_ gnd vdd FILL
X_2925_ _3289_/Q _3023_/A vdd gnd INVX1
XFILL_3__2006_ gnd vdd FILL
XFILL_1__2070_ gnd vdd FILL
X_2856_ _2868_/B _2857_/C vdd gnd INVX1
XFILL_0__2228_ gnd vdd FILL
XFILL_6__1996_ gnd vdd FILL
XBUFX2_insert19 _2580_/Y _3362_/R vdd gnd BUFX2
X_1807_ _2437_/A _2289_/B vdd gnd INVX1
XFILL_0__2159_ gnd vdd FILL
X_2787_ _3258_/Q _2814_/A _2788_/C vdd gnd NAND2X1
XFILL_4__2750_ gnd vdd FILL
XFILL_3__2908_ gnd vdd FILL
XFILL_1__2972_ gnd vdd FILL
XFILL_4__1701_ gnd vdd FILL
XFILL_4__2681_ gnd vdd FILL
X_1738_ _3151_/A _2446_/B vdd gnd INVX2
XFILL_3__2839_ gnd vdd FILL
XFILL_9__2326_ gnd vdd FILL
XFILL_7__2390_ gnd vdd FILL
XFILL_6__3597_ gnd vdd FILL
XFILL_1__1923_ gnd vdd FILL
XFILL_6__2617_ gnd vdd FILL
X_3408_ _3413_/B _3408_/B _3459_/A _3409_/A vdd gnd OAI21X1
XFILL_1__1854_ gnd vdd FILL
XFILL_6__2548_ gnd vdd FILL
XFILL_6__2479_ gnd vdd FILL
X_3339_ _3339_/D vdd _3353_/R _3577_/CLK _3339_/Q vdd gnd DFFSR
XFILL_7__3011_ gnd vdd FILL
XFILL_1__1785_ gnd vdd FILL
XFILL_1__3524_ gnd vdd FILL
XFILL_1__3455_ gnd vdd FILL
XFILL_4__3164_ gnd vdd FILL
XFILL_1__2406_ gnd vdd FILL
XFILL_4__3095_ gnd vdd FILL
XFILL_1__3386_ gnd vdd FILL
XFILL_4__2115_ gnd vdd FILL
XFILL_1__2337_ gnd vdd FILL
XFILL_4__2046_ gnd vdd FILL
XFILL_1__2268_ gnd vdd FILL
XFILL_5__2790_ gnd vdd FILL
XFILL_7__2726_ gnd vdd FILL
XFILL_5__1810_ gnd vdd FILL
XFILL_1__2199_ gnd vdd FILL
XFILL_4__2948_ gnd vdd FILL
XFILL_5__1741_ gnd vdd FILL
XFILL_2__1963_ gnd vdd FILL
XFILL_7__2657_ gnd vdd FILL
XFILL_5__3411_ gnd vdd FILL
XFILL_4__2879_ gnd vdd FILL
XFILL_7__2588_ gnd vdd FILL
XFILL_8__3120_ gnd vdd FILL
XFILL_2__1894_ gnd vdd FILL
XFILL_8__3051_ gnd vdd FILL
XFILL_8__2002_ gnd vdd FILL
XFILL_2__3564_ gnd vdd FILL
XFILL_2__3495_ gnd vdd FILL
XFILL_7__3209_ gnd vdd FILL
XFILL_5__2224_ gnd vdd FILL
XFILL_2__2515_ gnd vdd FILL
XFILL_2__2446_ gnd vdd FILL
XFILL_5__2155_ gnd vdd FILL
XFILL_5__2086_ gnd vdd FILL
XFILL_2__2377_ gnd vdd FILL
XFILL_0__3200_ gnd vdd FILL
XFILL_8__2904_ gnd vdd FILL
XFILL_0__3131_ gnd vdd FILL
XFILL_8__2835_ gnd vdd FILL
XFILL_0__3062_ gnd vdd FILL
X_2710_ _2724_/A _2733_/B _2767_/A _2711_/C vdd gnd OAI21X1
XFILL_6__1850_ gnd vdd FILL
XFILL_0__2013_ gnd vdd FILL
XFILL_5__2988_ gnd vdd FILL
XFILL_8__2766_ gnd vdd FILL
XFILL_6__1781_ gnd vdd FILL
XFILL_6__3520_ gnd vdd FILL
XFILL_8__1717_ gnd vdd FILL
XFILL_8__2697_ gnd vdd FILL
X_2641_ _2675_/A _2641_/B _2641_/C _2641_/D _3242_/D vdd gnd OAI22X1
XFILL_5__1939_ gnd vdd FILL
X_2572_ _3232_/A _2572_/B _2572_/C _2573_/A vdd gnd OAI21X1
XFILL_6__3451_ gnd vdd FILL
XFILL_0__2915_ gnd vdd FILL
XFILL_6__3382_ gnd vdd FILL
XFILL_6__2402_ gnd vdd FILL
XFILL_2_BUFX2_insert0 gnd vdd FILL
XFILL_9__3091_ gnd vdd FILL
XFILL_6__2333_ gnd vdd FILL
XFILL_3__2624_ gnd vdd FILL
XFILL_0__2846_ gnd vdd FILL
XFILL_3__2555_ gnd vdd FILL
X_3124_ _3141_/A _3126_/B _3124_/C _3337_/D vdd gnd OAI21X1
XFILL_6__2264_ gnd vdd FILL
XFILL_0__2777_ gnd vdd FILL
XFILL_6__2195_ gnd vdd FILL
X_3055_ _3055_/A _3056_/C vdd gnd INVX1
XFILL_3__2486_ gnd vdd FILL
XFILL_0__1728_ gnd vdd FILL
X_2006_ _2006_/A _3293_/D _2006_/C _2854_/A vdd gnd OAI21X1
XFILL_9__2944_ gnd vdd FILL
XFILL_3__3107_ gnd vdd FILL
XFILL_6_BUFX2_insert80 gnd vdd FILL
XFILL_1__3171_ gnd vdd FILL
XFILL_6_BUFX2_insert91 gnd vdd FILL
XFILL_3__3038_ gnd vdd FILL
XFILL_1__2122_ gnd vdd FILL
XFILL_7__1890_ gnd vdd FILL
X_2908_ _2908_/A _2928_/B _2957_/B _2935_/A vdd gnd OAI21X1
XFILL_1__2053_ gnd vdd FILL
XFILL_7__3560_ gnd vdd FILL
XFILL_6__1979_ gnd vdd FILL
X_2839_ _2839_/A _2843_/C _2867_/A vdd gnd NOR2X1
XFILL_4__2802_ gnd vdd FILL
XFILL_7__3491_ gnd vdd FILL
XFILL_7__2511_ gnd vdd FILL
XFILL_4__2733_ gnd vdd FILL
XFILL_1__2955_ gnd vdd FILL
XFILL_7__2442_ gnd vdd FILL
XFILL_7__2373_ gnd vdd FILL
XFILL_4__2664_ gnd vdd FILL
XFILL_1__1906_ gnd vdd FILL
XFILL_1__2886_ gnd vdd FILL
XFILL_4__2595_ gnd vdd FILL
XFILL_1__1837_ gnd vdd FILL
XFILL_1__1768_ gnd vdd FILL
XFILL_1__3507_ gnd vdd FILL
XFILL_2__2300_ gnd vdd FILL
XFILL_4__3216_ gnd vdd FILL
XFILL_5_BUFX2_insert4 gnd vdd FILL
XFILL_1__1699_ gnd vdd FILL
XFILL_1__3438_ gnd vdd FILL
XFILL_4__3147_ gnd vdd FILL
XFILL_2__2231_ gnd vdd FILL
XFILL_2__2162_ gnd vdd FILL
XFILL_1__3369_ gnd vdd FILL
XFILL_4__3078_ gnd vdd FILL
XFILL_5__2911_ gnd vdd FILL
XFILL_4__2029_ gnd vdd FILL
XFILL_8__2620_ gnd vdd FILL
XFILL_2__2093_ gnd vdd FILL
XFILL_5__2842_ gnd vdd FILL
XFILL_8__2551_ gnd vdd FILL
XFILL_8__2482_ gnd vdd FILL
XFILL_7__2709_ gnd vdd FILL
XFILL_5__2773_ gnd vdd FILL
XFILL_2__2995_ gnd vdd FILL
XFILL_5__1724_ gnd vdd FILL
XFILL_2__1946_ gnd vdd FILL
XFILL_2__1877_ gnd vdd FILL
XFILL_0__2700_ gnd vdd FILL
XFILL_8__3103_ gnd vdd FILL
XFILL_2__3547_ gnd vdd FILL
XFILL_8__3034_ gnd vdd FILL
XFILL_3__2340_ gnd vdd FILL
XFILL_0__2631_ gnd vdd FILL
XFILL_0__2562_ gnd vdd FILL
XFILL_2__3478_ gnd vdd FILL
XFILL_3__2271_ gnd vdd FILL
XFILL_5__2207_ gnd vdd FILL
XFILL_5__3187_ gnd vdd FILL
XFILL_0__2493_ gnd vdd FILL
XFILL_5__2138_ gnd vdd FILL
XFILL_2__2429_ gnd vdd FILL
XFILL_6__2951_ gnd vdd FILL
XFILL_5__2069_ gnd vdd FILL
XFILL_0__3114_ gnd vdd FILL
XFILL_6__2882_ gnd vdd FILL
XFILL_6__1902_ gnd vdd FILL
XFILL_8__2818_ gnd vdd FILL
XFILL_8_BUFX2_insert8 gnd vdd FILL
XFILL_9__2591_ gnd vdd FILL
XFILL_0__3045_ gnd vdd FILL
XFILL_8__2749_ gnd vdd FILL
XFILL_6__1833_ gnd vdd FILL
XFILL_6__1764_ gnd vdd FILL
X_2624_ _3350_/Q _2770_/C _2625_/C vdd gnd NAND2X1
XFILL_6__3503_ gnd vdd FILL
XFILL_3__1986_ gnd vdd FILL
XFILL_6__1695_ gnd vdd FILL
XFILL_6__3434_ gnd vdd FILL
X_2555_ _3575_/Q _3071_/A vdd gnd INVX1
X_2486_ _2508_/B _2511_/A _3574_/Q _2488_/A vdd gnd OAI21X1
XFILL_1__2740_ gnd vdd FILL
XFILL_6__3365_ gnd vdd FILL
XFILL_3__2607_ gnd vdd FILL
XFILL_1__2671_ gnd vdd FILL
XFILL_0__2829_ gnd vdd FILL
XFILL_3__3587_ gnd vdd FILL
XFILL_4__2380_ gnd vdd FILL
XFILL_6__2316_ gnd vdd FILL
X_3107_ _3125_/A _3107_/B _3330_/Q _3108_/C vdd gnd OAI21X1
XFILL_6__2247_ gnd vdd FILL
XFILL_3__2538_ gnd vdd FILL
XFILL_3__2469_ gnd vdd FILL
X_3038_ _3569_/Q _3085_/B _3057_/A vdd gnd NOR2X1
XFILL_4__3001_ gnd vdd FILL
XFILL_6__2178_ gnd vdd FILL
XFILL_7__2991_ gnd vdd FILL
XFILL_1__3223_ gnd vdd FILL
XFILL_7__1942_ gnd vdd FILL
XFILL_1__3154_ gnd vdd FILL
XFILL_1__2105_ gnd vdd FILL
XFILL_7__1873_ gnd vdd FILL
XFILL_1__3085_ gnd vdd FILL
XFILL_1__2036_ gnd vdd FILL
XFILL_7__3543_ gnd vdd FILL
XFILL_2__1800_ gnd vdd FILL
XFILL_7__3474_ gnd vdd FILL
XFILL_4__2716_ gnd vdd FILL
XFILL_2__2780_ gnd vdd FILL
XFILL_7__2425_ gnd vdd FILL
XFILL_1__2938_ gnd vdd FILL
XFILL_2__1731_ gnd vdd FILL
XFILL_4__2647_ gnd vdd FILL
XFILL_1__2869_ gnd vdd FILL
XFILL_7__2356_ gnd vdd FILL
XFILL_4__2578_ gnd vdd FILL
XFILL_2__3401_ gnd vdd FILL
XFILL_7__2287_ gnd vdd FILL
XFILL_5__3110_ gnd vdd FILL
XFILL_5__3041_ gnd vdd FILL
XFILL_2__2214_ gnd vdd FILL
XFILL_8__1982_ gnd vdd FILL
XFILL_2__3194_ gnd vdd FILL
XFILL_2__2145_ gnd vdd FILL
XFILL_2__2076_ gnd vdd FILL
XFILL_8__3583_ gnd vdd FILL
XFILL_8__2603_ gnd vdd FILL
XFILL_5__2825_ gnd vdd FILL
XFILL_8__2534_ gnd vdd FILL
XFILL_2_CLKBUF1_insert36 gnd vdd FILL
XFILL_5__2756_ gnd vdd FILL
XFILL_3__1840_ gnd vdd FILL
XFILL_2__2978_ gnd vdd FILL
XFILL_3__1771_ gnd vdd FILL
XFILL_5__1707_ gnd vdd FILL
XFILL_8__2465_ gnd vdd FILL
XFILL_2__1929_ gnd vdd FILL
XFILL_3__3510_ gnd vdd FILL
XFILL_0__1993_ gnd vdd FILL
XFILL_8__2396_ gnd vdd FILL
X_2340_ _2340_/A _2341_/B vdd gnd INVX1
XFILL_5__2687_ gnd vdd FILL
X_2271_ _2307_/B _2314_/A _2271_/C _2272_/A vdd gnd NAND3X1
XFILL_3__3441_ gnd vdd FILL
XFILL_6__3150_ gnd vdd FILL
XFILL_6__3081_ gnd vdd FILL
XFILL_0_BUFX2_insert18 gnd vdd FILL
XFILL_3__3372_ gnd vdd FILL
XFILL_6__2101_ gnd vdd FILL
XFILL184050x150 gnd vdd FILL
XFILL_0__2614_ gnd vdd FILL
XFILL_6__2032_ gnd vdd FILL
XFILL_8__3017_ gnd vdd FILL
XFILL_3__2323_ gnd vdd FILL
XFILL_0__3594_ gnd vdd FILL
XFILL_3__2254_ gnd vdd FILL
XFILL_0__2545_ gnd vdd FILL
XFILL_0__2476_ gnd vdd FILL
XFILL_3__2185_ gnd vdd FILL
XFILL_6__2934_ gnd vdd FILL
X_1986_ _1986_/A _1986_/B _1986_/C _3565_/A vdd gnd OAI21X1
XFILL_6__2865_ gnd vdd FILL
XFILL_0__3028_ gnd vdd FILL
XFILL_4__1880_ gnd vdd FILL
XFILL_6__1816_ gnd vdd FILL
XFILL_6__2796_ gnd vdd FILL
XFILL_4__3550_ gnd vdd FILL
XFILL_3__1969_ gnd vdd FILL
X_3587_ _3587_/A AB[2] vdd gnd BUFX2
XFILL_6__1747_ gnd vdd FILL
X_2607_ _3147_/C _2889_/C _2770_/C vdd gnd NOR2X1
XFILL_4__2501_ gnd vdd FILL
X_2538_ _3359_/Q _2538_/B _2540_/B vdd gnd NAND2X1
XFILL_4__3481_ gnd vdd FILL
XFILL_6__3417_ gnd vdd FILL
XFILL_7__2210_ gnd vdd FILL
XFILL_1__2723_ gnd vdd FILL
XFILL_7__3190_ gnd vdd FILL
XFILL_7__2141_ gnd vdd FILL
X_2469_ _3203_/B _3580_/A vdd gnd INVX1
XFILL_4__2432_ gnd vdd FILL
XFILL_4__2363_ gnd vdd FILL
XFILL_1__2654_ gnd vdd FILL
XFILL_7__2072_ gnd vdd FILL
XFILL_1__2585_ gnd vdd FILL
XFILL_4__2294_ gnd vdd FILL
XFILL_1__3206_ gnd vdd FILL
XFILL_7__2974_ gnd vdd FILL
XFILL_1__3137_ gnd vdd FILL
XFILL_7__1925_ gnd vdd FILL
XFILL_1__3068_ gnd vdd FILL
XFILL_7__1856_ gnd vdd FILL
XFILL_1__2019_ gnd vdd FILL
XFILL_2__2901_ gnd vdd FILL
XFILL_5__3590_ gnd vdd FILL
XFILL_5__2610_ gnd vdd FILL
XFILL_7__1787_ gnd vdd FILL
XFILL_7__3526_ gnd vdd FILL
XFILL_2__2832_ gnd vdd FILL
XFILL_5__2541_ gnd vdd FILL
XFILL_8__2250_ gnd vdd FILL
XFILL_7__3457_ gnd vdd FILL
XFILL_2__2763_ gnd vdd FILL
XFILL_8__2181_ gnd vdd FILL
XFILL_5__2472_ gnd vdd FILL
XFILL_2__1714_ gnd vdd FILL
XFILL_7__2408_ gnd vdd FILL
XFILL_7__3388_ gnd vdd FILL
XFILL_2__2694_ gnd vdd FILL
XFILL_7__2339_ gnd vdd FILL
XFILL_7_BUFX2_insert13 gnd vdd FILL
XFILL_7_BUFX2_insert24 gnd vdd FILL
XFILL_7_BUFX2_insert46 gnd vdd FILL
XFILL_7_BUFX2_insert57 gnd vdd FILL
XFILL_7_BUFX2_insert79 gnd vdd FILL
XFILL_7_BUFX2_insert68 gnd vdd FILL
XFILL182550x101550 gnd vdd FILL
XFILL_0__2330_ gnd vdd FILL
XFILL_5__3024_ gnd vdd FILL
XFILL_8__1965_ gnd vdd FILL
XFILL_0__2261_ gnd vdd FILL
XFILL_2__3177_ gnd vdd FILL
XFILL_2__2128_ gnd vdd FILL
XFILL_0__2192_ gnd vdd FILL
X_1840_ _3165_/A _2091_/B _1841_/A vdd gnd NAND2X1
XFILL_8__1896_ gnd vdd FILL
X_3510_ _3510_/A _3511_/B vdd gnd INVX1
XFILL_3__2941_ gnd vdd FILL
X_1771_ _2448_/C _1771_/B _1771_/C _1772_/C vdd gnd OAI21X1
XFILL_2__2059_ gnd vdd FILL
XFILL_6__2650_ gnd vdd FILL
XFILL_5__2808_ gnd vdd FILL
XFILL_8__3566_ gnd vdd FILL
XFILL_3__2872_ gnd vdd FILL
XFILL_8__3497_ gnd vdd FILL
X_3441_ _3441_/A _3441_/B _3441_/C _3482_/A vdd gnd OAI21X1
XFILL_3__1823_ gnd vdd FILL
XFILL_8__2517_ gnd vdd FILL
XFILL_6__2581_ gnd vdd FILL
X_3372_ _3372_/A _3372_/B _3372_/Y vdd gnd XNOR2X1
XFILL_5__2739_ gnd vdd FILL
XFILL_8__2448_ gnd vdd FILL
X_2323_ _2323_/A _2323_/B _2324_/C vdd gnd NOR2X1
XFILL_3__1754_ gnd vdd FILL
XFILL_0__1976_ gnd vdd FILL
XFILL_8__2379_ gnd vdd FILL
XFILL_6__3202_ gnd vdd FILL
XFILL_6__3133_ gnd vdd FILL
X_2254_ _2254_/A _2273_/A vdd gnd INVX1
XFILL_3__3424_ gnd vdd FILL
X_2185_ _2823_/B _2928_/A vdd gnd INVX1
XFILL_1__2370_ gnd vdd FILL
XFILL_3__2306_ gnd vdd FILL
XFILL_6__3064_ gnd vdd FILL
XFILL_6__2015_ gnd vdd FILL
XFILL_0__2528_ gnd vdd FILL
XFILL_3__2237_ gnd vdd FILL
XFILL_3__2168_ gnd vdd FILL
XFILL_0__2459_ gnd vdd FILL
XFILL_6__2917_ gnd vdd FILL
XFILL_4__2981_ gnd vdd FILL
XFILL_7__1710_ gnd vdd FILL
XFILL_3__2099_ gnd vdd FILL
X_1969_ _2506_/A _1975_/B vdd gnd INVX1
XFILL_4__1932_ gnd vdd FILL
XFILL_7__2690_ gnd vdd FILL
XFILL_6__2848_ gnd vdd FILL
XFILL_4__1863_ gnd vdd FILL
XFILL_4__3602_ gnd vdd FILL
XFILL_6__2779_ gnd vdd FILL
XFILL_4__1794_ gnd vdd FILL
XFILL_4__3533_ gnd vdd FILL
XFILL_4__3464_ gnd vdd FILL
XFILL_4__2415_ gnd vdd FILL
XFILL_1__2706_ gnd vdd FILL
XFILL_7__3173_ gnd vdd FILL
XFILL_4__3395_ gnd vdd FILL
XFILL_7__2124_ gnd vdd FILL
XFILL_1__2637_ gnd vdd FILL
XFILL_4__2346_ gnd vdd FILL
XFILL_7__2055_ gnd vdd FILL
XFILL_2__3100_ gnd vdd FILL
XFILL_4__2277_ gnd vdd FILL
XFILL_1__2568_ gnd vdd FILL
XFILL_1__2499_ gnd vdd FILL
XFILL_2__3031_ gnd vdd FILL
XFILL_7__2957_ gnd vdd FILL
XFILL_8__1750_ gnd vdd FILL
XFILL_5__1972_ gnd vdd FILL
XFILL_7__1908_ gnd vdd FILL
XFILL_7__2888_ gnd vdd FILL
XFILL_8__3420_ gnd vdd FILL
XFILL_7__1839_ gnd vdd FILL
XFILL_7__3509_ gnd vdd FILL
XFILL_8__2302_ gnd vdd FILL
XFILL_2__2815_ gnd vdd FILL
XFILL_5__2524_ gnd vdd FILL
XFILL_0__1830_ gnd vdd FILL
XFILL_8__2233_ gnd vdd FILL
XFILL_2__2746_ gnd vdd FILL
XFILL_8__2164_ gnd vdd FILL
XFILL182850x105450 gnd vdd FILL
XFILL_5__2455_ gnd vdd FILL
XFILL_0__1761_ gnd vdd FILL
XFILL_2__2677_ gnd vdd FILL
XFILL_0__3500_ gnd vdd FILL
XFILL_5__2386_ gnd vdd FILL
XFILL_8__2095_ gnd vdd FILL
XFILL_0__1692_ gnd vdd FILL
XFILL_0__3431_ gnd vdd FILL
XFILL_3__3140_ gnd vdd FILL
XFILL_5__3007_ gnd vdd FILL
XFILL_3__3071_ gnd vdd FILL
XFILL_3__2022_ gnd vdd FILL
X_2941_ reset _2957_/C _3299_/Q _2942_/C vdd gnd OAI21X1
XFILL_0__2313_ gnd vdd FILL
XFILL_2__3229_ gnd vdd FILL
XFILL_8__2997_ gnd vdd FILL
XFILL_0__2244_ gnd vdd FILL
XFILL_8__1948_ gnd vdd FILL
X_2872_ _2993_/B _2872_/B _3022_/A _2873_/A vdd gnd OAI21X1
XFILL_8__1879_ gnd vdd FILL
X_1823_ _2641_/B _3189_/C _2948_/A _1831_/D _3428_/A vdd gnd OAI22X1
XFILL_0__2175_ gnd vdd FILL
XFILL_6__2702_ gnd vdd FILL
XFILL_3__2924_ gnd vdd FILL
XFILL_3_BUFX2_insert22 gnd vdd FILL
XFILL_3_BUFX2_insert11 gnd vdd FILL
X_1754_ _3166_/D _3157_/B _2589_/A _1810_/C vdd gnd OAI21X1
XFILL_8__3549_ gnd vdd FILL
XFILL_3_BUFX2_insert44 gnd vdd FILL
XFILL_3_BUFX2_insert55 gnd vdd FILL
XFILL_6__2633_ gnd vdd FILL
XFILL_3__2855_ gnd vdd FILL
X_3424_ _3445_/A _3428_/A _3424_/C _3455_/C _3426_/B vdd gnd AOI22X1
XFILL_3_BUFX2_insert88 gnd vdd FILL
XFILL_3_BUFX2_insert66 gnd vdd FILL
XFILL_6__2564_ gnd vdd FILL
XFILL_3_BUFX2_insert77 gnd vdd FILL
XFILL_1__1870_ gnd vdd FILL
XFILL_3__2786_ gnd vdd FILL
XFILL_3__1806_ gnd vdd FILL
XFILL_6__2495_ gnd vdd FILL
X_3355_ _3355_/D vdd _3355_/R _3355_/CLK _3355_/Q vdd gnd DFFSR
XFILL_3__1737_ gnd vdd FILL
X_3286_ _3286_/D vdd _3289_/R _3307_/CLK _3286_/Q vdd gnd DFFSR
XFILL_0__1959_ gnd vdd FILL
X_2306_ _2306_/A _2917_/C _2306_/C _2315_/A vdd gnd NAND3X1
XFILL_1__3540_ gnd vdd FILL
XFILL_1__3471_ gnd vdd FILL
XFILL_4__2200_ gnd vdd FILL
X_2237_ _2582_/B _2700_/B _2238_/B vdd gnd NOR2X1
XFILL_6__3116_ gnd vdd FILL
XFILL_3__3407_ gnd vdd FILL
XFILL_1__2422_ gnd vdd FILL
XFILL_4__3180_ gnd vdd FILL
X_2168_ _2889_/C _2889_/B _2899_/A vdd gnd NAND2X1
XFILL_4__2131_ gnd vdd FILL
XFILL_6__3047_ gnd vdd FILL
XFILL_1__2353_ gnd vdd FILL
XFILL_4__2062_ gnd vdd FILL
X_2099_ _3189_/B _3190_/B _2437_/C vdd gnd NAND2X1
XFILL_1__2284_ gnd vdd FILL
XFILL_7__2811_ gnd vdd FILL
XFILL_7__2742_ gnd vdd FILL
XFILL_4__2964_ gnd vdd FILL
XFILL_7__2673_ gnd vdd FILL
XFILL_4__2895_ gnd vdd FILL
XFILL_4__1915_ gnd vdd FILL
XFILL_4__1846_ gnd vdd FILL
XFILL_4__3516_ gnd vdd FILL
XFILL_1__1999_ gnd vdd FILL
XFILL_4__1777_ gnd vdd FILL
XFILL_2__3580_ gnd vdd FILL
XFILL_2__2600_ gnd vdd FILL
XFILL_2__2531_ gnd vdd FILL
XFILL_7__3225_ gnd vdd FILL
XFILL_4__3447_ gnd vdd FILL
XFILL_5__2240_ gnd vdd FILL
XFILL_7__3156_ gnd vdd FILL
XFILL_4__3378_ gnd vdd FILL
XFILL_5__2171_ gnd vdd FILL
XFILL_2__2462_ gnd vdd FILL
XFILL_7__2107_ gnd vdd FILL
XFILL_7__3087_ gnd vdd FILL
XFILL_2__2393_ gnd vdd FILL
XFILL_4__2329_ gnd vdd FILL
XFILL_8__2920_ gnd vdd FILL
XFILL_7__2038_ gnd vdd FILL
XFILL_8__2851_ gnd vdd FILL
XFILL_2__3014_ gnd vdd FILL
XFILL_8__1802_ gnd vdd FILL
XFILL_7_CLKBUF1_insert36 gnd vdd FILL
XFILL_8__2782_ gnd vdd FILL
XFILL_8__1733_ gnd vdd FILL
XFILL_5__1955_ gnd vdd FILL
XFILL_8__3403_ gnd vdd FILL
XFILL_5__1886_ gnd vdd FILL
XFILL_0__2931_ gnd vdd FILL
XFILL182850x117150 gnd vdd FILL
XFILL_3__2640_ gnd vdd FILL
XFILL_0__2862_ gnd vdd FILL
XFILL_5__3556_ gnd vdd FILL
XFILL_3__2571_ gnd vdd FILL
X_3140_ _3346_/Q _3143_/B _3141_/C vdd gnd NAND2X1
XFILL_5__3487_ gnd vdd FILL
XFILL_8__2216_ gnd vdd FILL
XFILL_0__2793_ gnd vdd FILL
XFILL_6__2280_ gnd vdd FILL
XFILL_5__2507_ gnd vdd FILL
XFILL_0__1813_ gnd vdd FILL
XFILL184050x101550 gnd vdd FILL
XFILL_0__1744_ gnd vdd FILL
XFILL_8__3196_ gnd vdd FILL
XFILL_2__2729_ gnd vdd FILL
XFILL_5__2438_ gnd vdd FILL
X_3071_ _3071_/A _3071_/B _3083_/B vdd gnd NOR2X1
XFILL_8__2147_ gnd vdd FILL
XFILL_8__2078_ gnd vdd FILL
X_2022_ _2022_/A _2993_/A _2022_/C _2161_/A vdd gnd OAI21X1
XFILL_5__2369_ gnd vdd FILL
XFILL_3__3123_ gnd vdd FILL
XFILL_0__3414_ gnd vdd FILL
XFILL_3__3054_ gnd vdd FILL
X_2924_ _2924_/A _2936_/B _2924_/C _3288_/D vdd gnd AOI21X1
XFILL_3__2005_ gnd vdd FILL
X_2855_ _2880_/A _2855_/B _2855_/C _2868_/B vdd gnd OAI21X1
XFILL_0__2227_ gnd vdd FILL
XFILL_6__1995_ gnd vdd FILL
XFILL_9__3443_ gnd vdd FILL
XFILL_0__2158_ gnd vdd FILL
X_1806_ _1806_/A _1806_/B _1815_/A vdd gnd NOR2X1
X_2786_ _2786_/A _2786_/B _2801_/B _3257_/D vdd gnd OAI21X1
XFILL_3__2907_ gnd vdd FILL
XFILL_4__1700_ gnd vdd FILL
XFILL_1__2971_ gnd vdd FILL
XFILL_0__2089_ gnd vdd FILL
X_1737_ _2594_/B _1933_/C _3151_/A vdd gnd NOR2X1
XFILL_4__2680_ gnd vdd FILL
XFILL_6__2616_ gnd vdd FILL
XFILL_3__2838_ gnd vdd FILL
XFILL_6__3596_ gnd vdd FILL
XFILL_1__1922_ gnd vdd FILL
X_3407_ _3445_/A _3411_/A _3407_/C _3455_/C _3409_/B vdd gnd AOI22X1
XFILL_1__1853_ gnd vdd FILL
XFILL_6__2547_ gnd vdd FILL
X_3338_ _3338_/D vdd _3347_/R _3573_/CLK _3338_/Q vdd gnd DFFSR
XFILL_6__2478_ gnd vdd FILL
XFILL_3__2769_ gnd vdd FILL
XFILL_7__3010_ gnd vdd FILL
XFILL_1__1784_ gnd vdd FILL
XFILL_1__3523_ gnd vdd FILL
X_3269_ _3269_/D vdd _3282_/R _3313_/CLK _3269_/Q vdd gnd DFFSR
XFILL_4__3232_ gnd vdd FILL
XFILL_1__3454_ gnd vdd FILL
XFILL_4__3163_ gnd vdd FILL
XFILL_1__3385_ gnd vdd FILL
XFILL_4__2114_ gnd vdd FILL
XFILL_1__2405_ gnd vdd FILL
XFILL_4__3094_ gnd vdd FILL
XFILL_1__2336_ gnd vdd FILL
XFILL_4__2045_ gnd vdd FILL
XFILL_1__2267_ gnd vdd FILL
XFILL_1__2198_ gnd vdd FILL
XFILL184350x62550 gnd vdd FILL
XFILL_7__2725_ gnd vdd FILL
XFILL_4__2947_ gnd vdd FILL
XFILL_5__1740_ gnd vdd FILL
XFILL_2__1962_ gnd vdd FILL
XFILL_7__2656_ gnd vdd FILL
XFILL_5__3410_ gnd vdd FILL
XFILL_4__2878_ gnd vdd FILL
XFILL_7__2587_ gnd vdd FILL
XFILL_2__1893_ gnd vdd FILL
XFILL_4__1829_ gnd vdd FILL
XFILL_8__3050_ gnd vdd FILL
XFILL_8__2001_ gnd vdd FILL
XFILL_2__3563_ gnd vdd FILL
XFILL_7__3208_ gnd vdd FILL
XFILL_2__3494_ gnd vdd FILL
XFILL_5__2223_ gnd vdd FILL
XFILL_2__2514_ gnd vdd FILL
XFILL_7__3139_ gnd vdd FILL
XFILL_2__2445_ gnd vdd FILL
XFILL_5__2154_ gnd vdd FILL
XFILL_8__2903_ gnd vdd FILL
XFILL_5__2085_ gnd vdd FILL
XFILL_2__2376_ gnd vdd FILL
XFILL_0__3130_ gnd vdd FILL
XFILL_8__2834_ gnd vdd FILL
XFILL_0__3061_ gnd vdd FILL
XFILL_8__2765_ gnd vdd FILL
XFILL_0__2012_ gnd vdd FILL
XFILL_5__2987_ gnd vdd FILL
XFILL_6__1780_ gnd vdd FILL
XFILL_8__1716_ gnd vdd FILL
X_2640_ _2675_/A _2741_/C _2641_/C vdd gnd NAND2X1
XFILL_5__1938_ gnd vdd FILL
XFILL_8__2696_ gnd vdd FILL
X_2571_ _2571_/A _2571_/B _2572_/C vdd gnd NOR2X1
XFILL_6__3450_ gnd vdd FILL
XFILL_5__1869_ gnd vdd FILL
XFILL184350x105450 gnd vdd FILL
XFILL_0__2914_ gnd vdd FILL
XFILL_6__3381_ gnd vdd FILL
XFILL_6__2401_ gnd vdd FILL
XFILL_2_BUFX2_insert1 gnd vdd FILL
XFILL_5__3539_ gnd vdd FILL
XFILL_6__2332_ gnd vdd FILL
XFILL_3__2623_ gnd vdd FILL
XFILL_0__2845_ gnd vdd FILL
XFILL_3__2554_ gnd vdd FILL
X_3123_ _3125_/A _3125_/B _3337_/Q _3124_/C vdd gnd OAI21X1
XFILL_6__2263_ gnd vdd FILL
XFILL_3__2485_ gnd vdd FILL
XFILL_0__2776_ gnd vdd FILL
XFILL_8__3179_ gnd vdd FILL
X_3054_ _3090_/A _3133_/A _3054_/C _3317_/D vdd gnd OAI21X1
XFILL_6__2194_ gnd vdd FILL
XFILL_0__1727_ gnd vdd FILL
X_2005_ _2006_/A _2005_/B _2702_/B _2006_/C vdd gnd AOI21X1
XFILL_3__3106_ gnd vdd FILL
XFILL_6_BUFX2_insert81 gnd vdd FILL
XFILL_1__3170_ gnd vdd FILL
XFILL_6_BUFX2_insert70 gnd vdd FILL
XFILL_6_BUFX2_insert92 gnd vdd FILL
XFILL_3__3037_ gnd vdd FILL
XFILL_9__1825_ gnd vdd FILL
XFILL_1__2121_ gnd vdd FILL
X_2907_ _2936_/B _2907_/B _2907_/C _3285_/D vdd gnd OAI21X1
XFILL_1__2052_ gnd vdd FILL
XFILL_6__1978_ gnd vdd FILL
X_2838_ _2910_/B _2857_/A _2839_/A vdd gnd NAND2X1
XFILL_4__2801_ gnd vdd FILL
XFILL_7__2510_ gnd vdd FILL
XFILL_7__3490_ gnd vdd FILL
XFILL_4__2732_ gnd vdd FILL
X_2769_ _2769_/A _2769_/B _3253_/D vdd gnd AND2X2
XFILL_1__2954_ gnd vdd FILL
XFILL_7__2441_ gnd vdd FILL
XFILL_7__2372_ gnd vdd FILL
XFILL_6__3579_ gnd vdd FILL
XFILL_1__1905_ gnd vdd FILL
XFILL_4__2663_ gnd vdd FILL
XFILL_1__2885_ gnd vdd FILL
XFILL_4__2594_ gnd vdd FILL
XFILL_1__1836_ gnd vdd FILL
XFILL_1__1767_ gnd vdd FILL
XFILL_1__3506_ gnd vdd FILL
XFILL_4__3215_ gnd vdd FILL
XFILL_5_BUFX2_insert5 gnd vdd FILL
XFILL_2__2230_ gnd vdd FILL
XFILL_1__1698_ gnd vdd FILL
XFILL_1__3437_ gnd vdd FILL
XFILL_4__3146_ gnd vdd FILL
XFILL_2__2161_ gnd vdd FILL
XFILL_4__3077_ gnd vdd FILL
XFILL_1__3368_ gnd vdd FILL
XFILL_1__2319_ gnd vdd FILL
XFILL184350x74250 gnd vdd FILL
XFILL_2__2092_ gnd vdd FILL
XFILL_5__2910_ gnd vdd FILL
XFILL_4__2028_ gnd vdd FILL
XFILL_5__2841_ gnd vdd FILL
XFILL_8__2550_ gnd vdd FILL
XFILL_8__2481_ gnd vdd FILL
XFILL_7__2708_ gnd vdd FILL
XFILL_5__2772_ gnd vdd FILL
XFILL_2__2994_ gnd vdd FILL
XFILL_5__1723_ gnd vdd FILL
XFILL_7__2639_ gnd vdd FILL
XFILL_2__1945_ gnd vdd FILL
XFILL_2__1876_ gnd vdd FILL
XFILL_8__3102_ gnd vdd FILL
XFILL_2__3546_ gnd vdd FILL
XFILL_8__3033_ gnd vdd FILL
XFILL_0__2630_ gnd vdd FILL
XFILL_0__2561_ gnd vdd FILL
XFILL_2__3477_ gnd vdd FILL
XFILL_3__2270_ gnd vdd FILL
XFILL_5__2206_ gnd vdd FILL
XFILL_5__3186_ gnd vdd FILL
XFILL_2__2428_ gnd vdd FILL
XFILL_0__2492_ gnd vdd FILL
XFILL_5__2137_ gnd vdd FILL
XFILL_2__2359_ gnd vdd FILL
XFILL_6__2950_ gnd vdd FILL
XFILL_5__2068_ gnd vdd FILL
XFILL_0__3113_ gnd vdd FILL
XFILL_8__2817_ gnd vdd FILL
XFILL_6__2881_ gnd vdd FILL
XFILL_6__1901_ gnd vdd FILL
XFILL_0__3044_ gnd vdd FILL
XFILL184350x117150 gnd vdd FILL
XFILL184650x109350 gnd vdd FILL
XFILL_8_BUFX2_insert9 gnd vdd FILL
XFILL_6__1832_ gnd vdd FILL
XFILL_8__2748_ gnd vdd FILL
XFILL_6__1763_ gnd vdd FILL
XFILL_8__2679_ gnd vdd FILL
X_2623_ _3298_/Q _2623_/B _2625_/B vdd gnd NOR2X1
XFILL_6__3502_ gnd vdd FILL
XFILL_3__1985_ gnd vdd FILL
XFILL_6__1694_ gnd vdd FILL
X_2554_ _3361_/Q _3228_/A vdd gnd INVX1
XFILL_6__3433_ gnd vdd FILL
X_2485_ _3207_/B _3588_/A vdd gnd INVX1
XFILL_6__3364_ gnd vdd FILL
XFILL_3__2606_ gnd vdd FILL
XFILL_1__2670_ gnd vdd FILL
XFILL_0__2828_ gnd vdd FILL
XFILL_6__2315_ gnd vdd FILL
XFILL_3__3586_ gnd vdd FILL
X_3106_ _3141_/A _3108_/B _3106_/C _3329_/D vdd gnd OAI21X1
XFILL_6__2246_ gnd vdd FILL
XFILL_3__2537_ gnd vdd FILL
XFILL_3__2468_ gnd vdd FILL
XFILL_0__2759_ gnd vdd FILL
X_3037_ _3056_/B _3039_/A vdd gnd INVX1
XFILL_4__3000_ gnd vdd FILL
XFILL_3__2399_ gnd vdd FILL
XFILL_6__2177_ gnd vdd FILL
XFILL_7__2990_ gnd vdd FILL
XFILL_1__3222_ gnd vdd FILL
XFILL_7__1941_ gnd vdd FILL
XFILL_1__3153_ gnd vdd FILL
XFILL_1__2104_ gnd vdd FILL
XFILL_7__1872_ gnd vdd FILL
XFILL_1__3084_ gnd vdd FILL
XFILL_1__2035_ gnd vdd FILL
XFILL_7__3542_ gnd vdd FILL
XFILL_7__3473_ gnd vdd FILL
XFILL_7__2424_ gnd vdd FILL
XFILL_4__2715_ gnd vdd FILL
XFILL_2__1730_ gnd vdd FILL
XFILL_1__2937_ gnd vdd FILL
XFILL_4__2646_ gnd vdd FILL
XFILL_2_BUFX2_insert90 gnd vdd FILL
XFILL_1__2868_ gnd vdd FILL
XFILL_7__2355_ gnd vdd FILL
XFILL_2__3400_ gnd vdd FILL
XFILL_4__2577_ gnd vdd FILL
XFILL_1__1819_ gnd vdd FILL
XFILL_7__2286_ gnd vdd FILL
XFILL_1__2799_ gnd vdd FILL
XFILL_5__3040_ gnd vdd FILL
XFILL_2__2213_ gnd vdd FILL
XFILL_8__1981_ gnd vdd FILL
XFILL_2__3193_ gnd vdd FILL
XFILL_4__3129_ gnd vdd FILL
XFILL_2__2144_ gnd vdd FILL
XFILL_2__2075_ gnd vdd FILL
XFILL_8__2602_ gnd vdd FILL
XFILL_8__3582_ gnd vdd FILL
XFILL_5__2824_ gnd vdd FILL
XFILL_8__2533_ gnd vdd FILL
XFILL_2_CLKBUF1_insert37 gnd vdd FILL
XFILL_5__2755_ gnd vdd FILL
XFILL_2__2977_ gnd vdd FILL
XFILL_3__1770_ gnd vdd FILL
XFILL_5__1706_ gnd vdd FILL
XFILL_8__2464_ gnd vdd FILL
XFILL_2__1928_ gnd vdd FILL
XFILL_8__2395_ gnd vdd FILL
XFILL_0__1992_ gnd vdd FILL
XFILL_5__2686_ gnd vdd FILL
X_2270_ _2270_/A _2311_/A _2305_/B _2271_/C vdd gnd AOI21X1
XFILL_3__3440_ gnd vdd FILL
XFILL_2__1859_ gnd vdd FILL
XFILL_0_CLKBUF1_insert30 gnd vdd FILL
XFILL_6__3080_ gnd vdd FILL
XFILL_8__3016_ gnd vdd FILL
XFILL_3__3371_ gnd vdd FILL
XFILL_0__2613_ gnd vdd FILL
XFILL_0_BUFX2_insert19 gnd vdd FILL
XFILL_6__2100_ gnd vdd FILL
XFILL_2__3529_ gnd vdd FILL
XFILL_3__2322_ gnd vdd FILL
XFILL_6__2031_ gnd vdd FILL
XFILL_0__3593_ gnd vdd FILL
XFILL_3__2253_ gnd vdd FILL
XFILL_0__2544_ gnd vdd FILL
XFILL_0__2475_ gnd vdd FILL
XFILL_5__3169_ gnd vdd FILL
XFILL_3__2184_ gnd vdd FILL
XFILL_6__2933_ gnd vdd FILL
X_1985_ _1985_/A _3577_/Q _1985_/C _1986_/C vdd gnd AOI21X1
XFILL_6__2864_ gnd vdd FILL
XFILL_0__3027_ gnd vdd FILL
XFILL_6__2795_ gnd vdd FILL
XFILL_6__1815_ gnd vdd FILL
XFILL_6__1746_ gnd vdd FILL
X_2606_ _3239_/Q _2685_/B _2609_/C vdd gnd NAND2X1
XFILL_3__1968_ gnd vdd FILL
X_3586_ _3586_/A AB[15] vdd gnd BUFX2
XFILL_4__2500_ gnd vdd FILL
X_2537_ _3250_/Q _2734_/B vdd gnd INVX1
XFILL_4__3480_ gnd vdd FILL
XFILL_6__3416_ gnd vdd FILL
XFILL_3__1899_ gnd vdd FILL
X_2468_ _2468_/A _2519_/C _2468_/C _3203_/B vdd gnd AOI21X1
XFILL_1__2722_ gnd vdd FILL
XFILL_7__2140_ gnd vdd FILL
XFILL_4__2431_ gnd vdd FILL
XFILL_4__2362_ gnd vdd FILL
X_2399_ _2423_/A _2484_/A _2404_/C vdd gnd NAND2X1
XFILL_1__2653_ gnd vdd FILL
XFILL_7__2071_ gnd vdd FILL
XFILL_1__2584_ gnd vdd FILL
XFILL_6__2229_ gnd vdd FILL
XFILL_4__2293_ gnd vdd FILL
XFILL_1__3205_ gnd vdd FILL
XFILL_7__2973_ gnd vdd FILL
XFILL_1__3136_ gnd vdd FILL
XFILL_7__1924_ gnd vdd FILL
XFILL_1__3067_ gnd vdd FILL
XFILL_7__1855_ gnd vdd FILL
XFILL_2__2900_ gnd vdd FILL
XFILL_1__2018_ gnd vdd FILL
XFILL_7__3525_ gnd vdd FILL
XFILL_7__1786_ gnd vdd FILL
XFILL_2__2831_ gnd vdd FILL
XFILL_5__2540_ gnd vdd FILL
XFILL_7__3456_ gnd vdd FILL
XFILL_2__2762_ gnd vdd FILL
XFILL_8__2180_ gnd vdd FILL
XFILL_7__3387_ gnd vdd FILL
XFILL_5__2471_ gnd vdd FILL
XFILL_2__1713_ gnd vdd FILL
XFILL_7__2407_ gnd vdd FILL
XFILL_7__2338_ gnd vdd FILL
XFILL_2__2693_ gnd vdd FILL
XFILL_4__2629_ gnd vdd FILL
XFILL_7__2269_ gnd vdd FILL
XFILL_7_BUFX2_insert25 gnd vdd FILL
XFILL_7_BUFX2_insert47 gnd vdd FILL
XFILL_7_BUFX2_insert14 gnd vdd FILL
XFILL_7_BUFX2_insert58 gnd vdd FILL
XFILL_7_BUFX2_insert69 gnd vdd FILL
XFILL_5__3023_ gnd vdd FILL
XFILL_0__2260_ gnd vdd FILL
XFILL_8__1964_ gnd vdd FILL
XFILL_2__3176_ gnd vdd FILL
XFILL_0__2191_ gnd vdd FILL
XFILL_2__2127_ gnd vdd FILL
XFILL_8__1895_ gnd vdd FILL
X_1770_ _3274_/Q _1770_/B _2072_/B _1771_/C vdd gnd OAI21X1
XFILL_2__2058_ gnd vdd FILL
XFILL_3__2940_ gnd vdd FILL
XFILL_5__2807_ gnd vdd FILL
XFILL_3__2871_ gnd vdd FILL
XFILL_8__3565_ gnd vdd FILL
XFILL_8__3496_ gnd vdd FILL
XFILL_6__2580_ gnd vdd FILL
X_3440_ _3459_/A _3440_/B _3441_/A vdd gnd NAND2X1
XFILL_8__2516_ gnd vdd FILL
XFILL_3__1822_ gnd vdd FILL
X_3371_ _3577_/Q _3567_/Q _3372_/B vdd gnd XNOR2X1
XFILL_8__2447_ gnd vdd FILL
XFILL_5__2738_ gnd vdd FILL
X_2322_ _2322_/A _2323_/B vdd gnd INVX1
XFILL_3__1753_ gnd vdd FILL
XFILL_5__2669_ gnd vdd FILL
XFILL_0__1975_ gnd vdd FILL
XFILL_8__2378_ gnd vdd FILL
XFILL_6__3201_ gnd vdd FILL
XFILL_6__3132_ gnd vdd FILL
X_2253_ _2306_/A _2306_/C _2254_/A vdd gnd NAND2X1
XFILL_3__3423_ gnd vdd FILL
X_2184_ _2184_/A _2184_/B _2184_/C _2328_/A vdd gnd NAND3X1
XFILL_3__2305_ gnd vdd FILL
XFILL_6__3063_ gnd vdd FILL
XFILL_6__2014_ gnd vdd FILL
XFILL_0__2527_ gnd vdd FILL
XFILL_3__2236_ gnd vdd FILL
XFILL_3__2167_ gnd vdd FILL
XFILL_0__2458_ gnd vdd FILL
XFILL_0__2389_ gnd vdd FILL
XFILL_6__2916_ gnd vdd FILL
XFILL_4__2980_ gnd vdd FILL
XFILL_3__2098_ gnd vdd FILL
X_1968_ _1968_/A _1968_/B _1968_/C _2506_/A vdd gnd NAND3X1
XFILL_6__2847_ gnd vdd FILL
XFILL_4__1931_ gnd vdd FILL
XFILL_4__1862_ gnd vdd FILL
X_1899_ _3192_/A _2938_/A vdd gnd INVX1
XFILL_4__3601_ gnd vdd FILL
XFILL_9__2487_ gnd vdd FILL
XFILL_6__2778_ gnd vdd FILL
X_3569_ _3569_/D vdd _3578_/R _3577_/CLK _3569_/Q vdd gnd DFFSR
XFILL_6__1729_ gnd vdd FILL
XFILL_4__1793_ gnd vdd FILL
XFILL_4__3532_ gnd vdd FILL
XFILL_4__3463_ gnd vdd FILL
XFILL_4__2414_ gnd vdd FILL
XFILL_1__2705_ gnd vdd FILL
XFILL_7__3172_ gnd vdd FILL
XFILL_4__3394_ gnd vdd FILL
XFILL_7__2123_ gnd vdd FILL
XFILL_1__2636_ gnd vdd FILL
XFILL_7__2054_ gnd vdd FILL
XFILL_4__2345_ gnd vdd FILL
XFILL_4__2276_ gnd vdd FILL
XFILL_1__2567_ gnd vdd FILL
XFILL_1__2498_ gnd vdd FILL
XFILL_2__3030_ gnd vdd FILL
XFILL_7__2956_ gnd vdd FILL
XFILL_1__3119_ gnd vdd FILL
XFILL_7__1907_ gnd vdd FILL
XFILL_5__1971_ gnd vdd FILL
XFILL_7__2887_ gnd vdd FILL
XFILL_7__1838_ gnd vdd FILL
XFILL_7__1769_ gnd vdd FILL
XFILL_7__3508_ gnd vdd FILL
XFILL_8__2301_ gnd vdd FILL
XFILL_2__2814_ gnd vdd FILL
XFILL_7__3439_ gnd vdd FILL
XFILL_8__2232_ gnd vdd FILL
XFILL_5__2523_ gnd vdd FILL
XFILL_5__2454_ gnd vdd FILL
XFILL_2__2745_ gnd vdd FILL
XFILL_8__2163_ gnd vdd FILL
XFILL_0__1760_ gnd vdd FILL
XFILL_2__2676_ gnd vdd FILL
XFILL_5__2385_ gnd vdd FILL
XFILL_0__1691_ gnd vdd FILL
XFILL_8__2094_ gnd vdd FILL
XFILL_0__3430_ gnd vdd FILL
XFILL_5__3006_ gnd vdd FILL
XFILL_3__3070_ gnd vdd FILL
X_2940_ _2940_/A _2956_/B vdd gnd INVX2
XFILL_3__2021_ gnd vdd FILL
XFILL_0__2312_ gnd vdd FILL
XFILL_8__2996_ gnd vdd FILL
XFILL_2__3228_ gnd vdd FILL
XFILL_8__1947_ gnd vdd FILL
X_2871_ _3007_/B _2898_/B _2871_/C _2871_/D _3277_/D vdd gnd OAI22X1
XFILL_0__2243_ gnd vdd FILL
XFILL_0__2174_ gnd vdd FILL
X_1822_ _3242_/Q _2641_/B vdd gnd INVX2
XFILL_2__3159_ gnd vdd FILL
XFILL_8__1878_ gnd vdd FILL
XFILL_6__2701_ gnd vdd FILL
XFILL_3__2923_ gnd vdd FILL
XFILL_3_BUFX2_insert12 gnd vdd FILL
X_1753_ _2594_/A _2442_/B _3157_/B vdd gnd NOR2X1
XFILL_8__3548_ gnd vdd FILL
XFILL_3_BUFX2_insert23 gnd vdd FILL
XFILL_3_BUFX2_insert56 gnd vdd FILL
XFILL_3_BUFX2_insert45 gnd vdd FILL
XFILL_6__2632_ gnd vdd FILL
XFILL_3__2854_ gnd vdd FILL
X_3423_ _3434_/A _3425_/B _3424_/C vdd gnd NAND2X1
XFILL_3_BUFX2_insert78 gnd vdd FILL
XFILL_3_BUFX2_insert67 gnd vdd FILL
XFILL_6__2563_ gnd vdd FILL
XFILL_3_BUFX2_insert89 gnd vdd FILL
XFILL_8__3479_ gnd vdd FILL
XFILL_3__2785_ gnd vdd FILL
XFILL_3__1805_ gnd vdd FILL
X_3354_ _3354_/D vdd _3355_/R _3578_/CLK _3354_/Q vdd gnd DFFSR
XFILL_6__2494_ gnd vdd FILL
XFILL_3__1736_ gnd vdd FILL
X_3285_ _3285_/D vdd _3289_/R _3307_/CLK _3285_/Q vdd gnd DFFSR
XFILL_0__1958_ gnd vdd FILL
X_2305_ _2305_/A _2305_/B _2917_/C vdd gnd NOR2X1
XFILL_1__3470_ gnd vdd FILL
XFILL_3__3406_ gnd vdd FILL
X_2236_ _2966_/B _2958_/A _2242_/A _2242_/C vdd gnd OAI21X1
XFILL_6__3115_ gnd vdd FILL
XFILL_0__1889_ gnd vdd FILL
XFILL_1__2421_ gnd vdd FILL
XFILL_6__3046_ gnd vdd FILL
X_2167_ _2167_/A _2172_/B vdd gnd INVX1
XFILL_4__2130_ gnd vdd FILL
XFILL_0__3559_ gnd vdd FILL
XFILL_1__2352_ gnd vdd FILL
XFILL_4__2061_ gnd vdd FILL
X_2098_ _2098_/A _2332_/A _2320_/C vdd gnd AND2X2
XFILL_1__2283_ gnd vdd FILL
XFILL_3__2219_ gnd vdd FILL
XFILL_7__2810_ gnd vdd FILL
XFILL_9__1987_ gnd vdd FILL
XFILL_3__3199_ gnd vdd FILL
XFILL_7__2741_ gnd vdd FILL
XFILL_4__2963_ gnd vdd FILL
XFILL_4__1914_ gnd vdd FILL
XFILL_7__2672_ gnd vdd FILL
XFILL_4__2894_ gnd vdd FILL
XFILL_4__1845_ gnd vdd FILL
XFILL_4__1776_ gnd vdd FILL
XFILL_4__3515_ gnd vdd FILL
XFILL_1__1998_ gnd vdd FILL
XFILL_2__2530_ gnd vdd FILL
XFILL_7__3224_ gnd vdd FILL
XFILL_4__3446_ gnd vdd FILL
XFILL_7__3155_ gnd vdd FILL
XFILL_4__3377_ gnd vdd FILL
XFILL_5__2170_ gnd vdd FILL
XFILL_2__2461_ gnd vdd FILL
XFILL_7__2106_ gnd vdd FILL
XFILL_7__3086_ gnd vdd FILL
XFILL_4__2328_ gnd vdd FILL
XFILL_1__3599_ gnd vdd FILL
XFILL_2__2392_ gnd vdd FILL
XFILL_1__2619_ gnd vdd FILL
XFILL_7__2037_ gnd vdd FILL
XFILL_8__2850_ gnd vdd FILL
XFILL_4__2259_ gnd vdd FILL
XFILL_2__3013_ gnd vdd FILL
XFILL_8__1801_ gnd vdd FILL
XFILL_7_CLKBUF1_insert37 gnd vdd FILL
XFILL_8__2781_ gnd vdd FILL
XFILL_7__2939_ gnd vdd FILL
XFILL_8__1732_ gnd vdd FILL
XFILL_5__1954_ gnd vdd FILL
XFILL_8__3402_ gnd vdd FILL
XFILL_5__1885_ gnd vdd FILL
XFILL_0__2930_ gnd vdd FILL
XFILL_5_CLKBUF1_insert30 gnd vdd FILL
XFILL_5__3555_ gnd vdd FILL
XFILL_0__2861_ gnd vdd FILL
XFILL_5__2506_ gnd vdd FILL
XFILL_3__2570_ gnd vdd FILL
XFILL_5__3486_ gnd vdd FILL
XFILL_8__2215_ gnd vdd FILL
XFILL_0__2792_ gnd vdd FILL
XFILL_8__3195_ gnd vdd FILL
XFILL_0__1812_ gnd vdd FILL
XFILL_2__2728_ gnd vdd FILL
X_3070_ _3071_/A _3071_/B _3073_/D vdd gnd NAND2X1
XFILL_8__2146_ gnd vdd FILL
XFILL_0__1743_ gnd vdd FILL
XFILL_5__2437_ gnd vdd FILL
X_2021_ _2022_/A _3306_/Q _2022_/C vdd gnd NAND2X1
XFILL_5__2368_ gnd vdd FILL
XFILL_2__2659_ gnd vdd FILL
XFILL_8__2077_ gnd vdd FILL
XFILL_3__3122_ gnd vdd FILL
XFILL_0__3413_ gnd vdd FILL
XFILL_5__2299_ gnd vdd FILL
XFILL_3__3053_ gnd vdd FILL
X_2923_ _2923_/A _2923_/B _2924_/C vdd gnd NOR2X1
XFILL_3__2004_ gnd vdd FILL
XFILL_8__2979_ gnd vdd FILL
X_2854_ _2854_/A _2932_/B _2915_/C _2855_/B vdd gnd NAND3X1
XFILL_6__1994_ gnd vdd FILL
XFILL_0__2226_ gnd vdd FILL
X_2785_ _2786_/A _2933_/A _2801_/B vdd gnd NAND2X1
XFILL_0__2157_ gnd vdd FILL
X_1805_ _3182_/C _1885_/A _1805_/C _1806_/B vdd gnd NAND3X1
XFILL_0__2088_ gnd vdd FILL
X_1736_ _3234_/Q _1762_/B _1933_/C vdd gnd NAND2X1
XFILL_3__2906_ gnd vdd FILL
XFILL_1__2970_ gnd vdd FILL
XFILL_6__2615_ gnd vdd FILL
XFILL_3__2837_ gnd vdd FILL
XFILL_1__1921_ gnd vdd FILL
XFILL_6__3595_ gnd vdd FILL
X_3406_ _3413_/B _3408_/B _3407_/C vdd gnd NAND2X1
XFILL_1__1852_ gnd vdd FILL
XFILL_6__2546_ gnd vdd FILL
X_3337_ _3337_/D vdd _3346_/R _3573_/CLK _3337_/Q vdd gnd DFFSR
XFILL_3__2768_ gnd vdd FILL
XFILL_6__2477_ gnd vdd FILL
XFILL_1__3522_ gnd vdd FILL
XFILL_3__1719_ gnd vdd FILL
XFILL_1__1783_ gnd vdd FILL
XFILL_3__2699_ gnd vdd FILL
X_3268_ _3268_/D vdd _3282_/R _3284_/CLK _3268_/Q vdd gnd DFFSR
XFILL_4__3231_ gnd vdd FILL
XFILL_1__3453_ gnd vdd FILL
X_2219_ _2299_/A _3156_/B _2278_/A _2220_/C vdd gnd OAI21X1
XFILL_4__3162_ gnd vdd FILL
X_3199_ _3230_/B _3215_/A vdd gnd INVX2
XFILL_1__3384_ gnd vdd FILL
XFILL_1__2404_ gnd vdd FILL
XFILL_4__2113_ gnd vdd FILL
XFILL_6__3029_ gnd vdd FILL
XFILL_4__3093_ gnd vdd FILL
XFILL_1__2335_ gnd vdd FILL
XFILL_4__2044_ gnd vdd FILL
XFILL_1__2266_ gnd vdd FILL
XFILL_1__2197_ gnd vdd FILL
XFILL_7__2724_ gnd vdd FILL
XFILL_4__2946_ gnd vdd FILL
XFILL_7__2655_ gnd vdd FILL
XFILL_4__2877_ gnd vdd FILL
XFILL_2__1961_ gnd vdd FILL
XFILL_2__1892_ gnd vdd FILL
XFILL_7__2586_ gnd vdd FILL
XFILL_4__1828_ gnd vdd FILL
XFILL_4__1759_ gnd vdd FILL
XFILL_8__2000_ gnd vdd FILL
XFILL_2__3562_ gnd vdd FILL
XFILL_7__3207_ gnd vdd FILL
XFILL_2__3493_ gnd vdd FILL
XFILL_4__3429_ gnd vdd FILL
XFILL_5__2222_ gnd vdd FILL
XFILL_2__2513_ gnd vdd FILL
XFILL_7__3138_ gnd vdd FILL
XFILL_2__2444_ gnd vdd FILL
XFILL_7__3069_ gnd vdd FILL
XFILL_5__2153_ gnd vdd FILL
XFILL_8__2902_ gnd vdd FILL
XFILL_5__2084_ gnd vdd FILL
XFILL_2__2375_ gnd vdd FILL
XFILL_8__2833_ gnd vdd FILL
XFILL_0__3060_ gnd vdd FILL
XFILL_8__2764_ gnd vdd FILL
XFILL_0__2011_ gnd vdd FILL
XFILL_5__2986_ gnd vdd FILL
XFILL_8__1715_ gnd vdd FILL
XFILL_5__1937_ gnd vdd FILL
XFILL_8__2695_ gnd vdd FILL
X_2570_ _2570_/A _2570_/B _2570_/C _2571_/B vdd gnd OAI21X1
XFILL_5__1868_ gnd vdd FILL
XFILL_6__2400_ gnd vdd FILL
XFILL_0__2913_ gnd vdd FILL
XFILL_6__3380_ gnd vdd FILL
XFILL_5__1799_ gnd vdd FILL
XFILL_3__2622_ gnd vdd FILL
XFILL_2_BUFX2_insert2 gnd vdd FILL
XFILL_0__2844_ gnd vdd FILL
XFILL_5__3538_ gnd vdd FILL
XFILL_6__2331_ gnd vdd FILL
X_3122_ _3139_/A _3126_/B _3122_/C _3336_/D vdd gnd OAI21X1
XFILL_5__3469_ gnd vdd FILL
XFILL_6__2262_ gnd vdd FILL
XFILL_3__2553_ gnd vdd FILL
XFILL_3__2484_ gnd vdd FILL
XFILL_0__2775_ gnd vdd FILL
XFILL_8__3178_ gnd vdd FILL
X_3053_ _3317_/Q _3090_/A _3054_/C vdd gnd NAND2X1
XFILL_6__2193_ gnd vdd FILL
XFILL_0__1726_ gnd vdd FILL
XFILL_8__2129_ gnd vdd FILL
X_2004_ _3302_/Q _2005_/B vdd gnd INVX1
XFILL_3__3105_ gnd vdd FILL
XFILL_6_BUFX2_insert60 gnd vdd FILL
XFILL_6_BUFX2_insert71 gnd vdd FILL
XFILL_6_BUFX2_insert93 gnd vdd FILL
XFILL_6_BUFX2_insert82 gnd vdd FILL
XFILL_3__3036_ gnd vdd FILL
XFILL_1__2120_ gnd vdd FILL
X_2906_ _2906_/A _2906_/B _3285_/Q _2907_/C vdd gnd OAI21X1
XFILL_1__2051_ gnd vdd FILL
XFILL_6__1977_ gnd vdd FILL
XFILL_0__2209_ gnd vdd FILL
X_2837_ _2837_/A _2919_/B _2837_/C _2862_/A _3270_/D vdd gnd AOI22X1
XFILL_4__2800_ gnd vdd FILL
XFILL_0__3189_ gnd vdd FILL
XFILL_4__2731_ gnd vdd FILL
X_2768_ _2768_/A _2768_/B _2769_/B vdd gnd NAND2X1
XFILL_1__2953_ gnd vdd FILL
X_1719_ _2602_/A _1888_/B _2123_/B _2700_/B vdd gnd NAND3X1
XFILL_7__2440_ gnd vdd FILL
X_2699_ _2726_/C _2699_/B _3043_/A _2704_/C vdd gnd AOI21X1
XFILL_7__2371_ gnd vdd FILL
XFILL_1__1904_ gnd vdd FILL
XFILL_4__2662_ gnd vdd FILL
XFILL_1__2884_ gnd vdd FILL
XFILL_6__2529_ gnd vdd FILL
XFILL_4__2593_ gnd vdd FILL
XFILL_1__1835_ gnd vdd FILL
XFILL_1__1766_ gnd vdd FILL
XFILL_1__3505_ gnd vdd FILL
XFILL_4__3214_ gnd vdd FILL
XFILL_1__3436_ gnd vdd FILL
XFILL_1__1697_ gnd vdd FILL
XFILL_5_BUFX2_insert6 gnd vdd FILL
XFILL184650x58650 gnd vdd FILL
XFILL_4__3145_ gnd vdd FILL
XFILL_2__2160_ gnd vdd FILL
XFILL_4__3076_ gnd vdd FILL
XFILL_1__3367_ gnd vdd FILL
XFILL_4__2027_ gnd vdd FILL
XFILL_1__2318_ gnd vdd FILL
XFILL_2__2091_ gnd vdd FILL
XFILL_1__2249_ gnd vdd FILL
XFILL_5__2840_ gnd vdd FILL
XFILL_5__2771_ gnd vdd FILL
XFILL_4__2929_ gnd vdd FILL
XFILL_2__2993_ gnd vdd FILL
XFILL_7__2707_ gnd vdd FILL
XFILL_5__1722_ gnd vdd FILL
XFILL_8__2480_ gnd vdd FILL
XFILL_7__2638_ gnd vdd FILL
XFILL_2__1944_ gnd vdd FILL
XFILL_7__2569_ gnd vdd FILL
XFILL_2__1875_ gnd vdd FILL
XFILL_8__3101_ gnd vdd FILL
XFILL181950x101550 gnd vdd FILL
XFILL_2__3545_ gnd vdd FILL
XFILL_8__3032_ gnd vdd FILL
XFILL_0__2560_ gnd vdd FILL
XFILL_2__3476_ gnd vdd FILL
XFILL_5__2205_ gnd vdd FILL
XFILL_5__3185_ gnd vdd FILL
XFILL_2__2427_ gnd vdd FILL
XFILL_0__2491_ gnd vdd FILL
XFILL_5__2136_ gnd vdd FILL
XFILL_2__2358_ gnd vdd FILL
XFILL_5__2067_ gnd vdd FILL
XFILL_0__3112_ gnd vdd FILL
XFILL_6__2880_ gnd vdd FILL
XFILL_8__2816_ gnd vdd FILL
XFILL_6__1900_ gnd vdd FILL
XFILL_2__2289_ gnd vdd FILL
XFILL_0__3043_ gnd vdd FILL
XFILL_6__1831_ gnd vdd FILL
XFILL_8__2747_ gnd vdd FILL
XFILL_6__3501_ gnd vdd FILL
XFILL_5__2969_ gnd vdd FILL
XFILL_8__2678_ gnd vdd FILL
XFILL_6__1762_ gnd vdd FILL
X_2622_ _3241_/Q _2778_/A _2629_/C vdd gnd NAND2X1
XFILL_3__1984_ gnd vdd FILL
XFILL_6__1693_ gnd vdd FILL
X_2553_ _3252_/Q _2751_/A vdd gnd INVX1
XFILL_6__3432_ gnd vdd FILL
X_2484_ _2484_/A _2519_/C _2484_/C _3207_/B vdd gnd AOI21X1
XFILL_6__2314_ gnd vdd FILL
XFILL_3__3585_ gnd vdd FILL
XFILL_3__2605_ gnd vdd FILL
XFILL_0__2827_ gnd vdd FILL
XFILL_3__2536_ gnd vdd FILL
X_3105_ _3111_/A _3107_/B _3329_/Q _3106_/C vdd gnd OAI21X1
XFILL_6__2245_ gnd vdd FILL
XFILL_0__2758_ gnd vdd FILL
X_3036_ _3569_/Q _3085_/B _3056_/B _3042_/B vdd gnd OAI21X1
XFILL_0__1709_ gnd vdd FILL
XFILL_3__2467_ gnd vdd FILL
XFILL_6__2176_ gnd vdd FILL
XFILL_3__2398_ gnd vdd FILL
XFILL_0__2689_ gnd vdd FILL
XFILL_1__3221_ gnd vdd FILL
XFILL_7__1940_ gnd vdd FILL
XFILL_1__3152_ gnd vdd FILL
XFILL_7__1871_ gnd vdd FILL
XFILL_9__2856_ gnd vdd FILL
XFILL_1__2103_ gnd vdd FILL
XFILL_3__3019_ gnd vdd FILL
XFILL_1__3083_ gnd vdd FILL
XFILL_1__2034_ gnd vdd FILL
XFILL_7__3541_ gnd vdd FILL
XFILL_7__3472_ gnd vdd FILL
XFILL_7__2423_ gnd vdd FILL
XFILL_4__2714_ gnd vdd FILL
XFILL_1__2936_ gnd vdd FILL
XFILL_4__2645_ gnd vdd FILL
XFILL_1__2867_ gnd vdd FILL
XFILL_7__2354_ gnd vdd FILL
XFILL_2_BUFX2_insert80 gnd vdd FILL
XFILL_2_BUFX2_insert91 gnd vdd FILL
XFILL_4__2576_ gnd vdd FILL
XFILL_7__2285_ gnd vdd FILL
XFILL_1__1818_ gnd vdd FILL
XFILL_1__2798_ gnd vdd FILL
XFILL_1__1749_ gnd vdd FILL
XFILL_4__3128_ gnd vdd FILL
XFILL_1__3419_ gnd vdd FILL
XFILL_8__1980_ gnd vdd FILL
XFILL_2__2212_ gnd vdd FILL
XFILL_2__3192_ gnd vdd FILL
XFILL_2__2143_ gnd vdd FILL
XFILL_4__3059_ gnd vdd FILL
XFILL_2__2074_ gnd vdd FILL
XFILL_5__2823_ gnd vdd FILL
XFILL_8__3581_ gnd vdd FILL
XFILL_8__2601_ gnd vdd FILL
XFILL_8__2532_ gnd vdd FILL
XFILL_2_CLKBUF1_insert38 gnd vdd FILL
XFILL_8__2463_ gnd vdd FILL
XFILL_5__2754_ gnd vdd FILL
XFILL_2__2976_ gnd vdd FILL
XFILL_5__1705_ gnd vdd FILL
XFILL_5__2685_ gnd vdd FILL
XFILL_2__1927_ gnd vdd FILL
XFILL_0__1991_ gnd vdd FILL
XFILL_8__2394_ gnd vdd FILL
XFILL_2__1858_ gnd vdd FILL
XFILL_8__3015_ gnd vdd FILL
XFILL_3__3370_ gnd vdd FILL
XFILL_0__2612_ gnd vdd FILL
XFILL_2__1789_ gnd vdd FILL
XFILL_0_CLKBUF1_insert31 gnd vdd FILL
XFILL_2__3528_ gnd vdd FILL
XFILL_6__2030_ gnd vdd FILL
XFILL_3__2321_ gnd vdd FILL
XFILL_0__3592_ gnd vdd FILL
XFILL_2__3459_ gnd vdd FILL
XFILL_3__2252_ gnd vdd FILL
XFILL_0__2543_ gnd vdd FILL
XFILL_0__2474_ gnd vdd FILL
XFILL_5__3168_ gnd vdd FILL
XFILL_5__3099_ gnd vdd FILL
XFILL_3__2183_ gnd vdd FILL
XFILL_5__2119_ gnd vdd FILL
XFILL_6__2932_ gnd vdd FILL
X_1984_ _2993_/A _1984_/B _2771_/C _1985_/C vdd gnd OAI21X1
XFILL_6__2863_ gnd vdd FILL
XFILL_6__2794_ gnd vdd FILL
XFILL_0__3026_ gnd vdd FILL
XFILL_6__1814_ gnd vdd FILL
X_2605_ _2692_/A _2670_/B _2605_/C _2685_/B vdd gnd OAI21X1
XFILL_6__1745_ gnd vdd FILL
XFILL_3__1967_ gnd vdd FILL
X_3585_ _3585_/A AB[14] vdd gnd BUFX2
X_2536_ _2715_/A _2574_/B _2536_/C _3581_/A vdd gnd OAI21X1
XFILL_6__3415_ gnd vdd FILL
XFILL_3__1898_ gnd vdd FILL
X_2467_ _2621_/B _2574_/B _2467_/C _2468_/C vdd gnd OAI21X1
XFILL_4__2430_ gnd vdd FILL
XFILL_1__2721_ gnd vdd FILL
XFILL_1__2652_ gnd vdd FILL
XFILL_4__2361_ gnd vdd FILL
X_2398_ _2398_/A _2398_/B _2398_/C _3597_/A vdd gnd NAND3X1
XFILL_7__2070_ gnd vdd FILL
XFILL_3__3499_ gnd vdd FILL
XFILL_6__2228_ gnd vdd FILL
XFILL_1__2583_ gnd vdd FILL
XFILL_3__2519_ gnd vdd FILL
XFILL_4__2292_ gnd vdd FILL
X_3019_ _3019_/A _3019_/B _3019_/C _3313_/D vdd gnd OAI21X1
XFILL_6__2159_ gnd vdd FILL
XFILL_1__3204_ gnd vdd FILL
XFILL_7__2972_ gnd vdd FILL
XFILL_1__3135_ gnd vdd FILL
XFILL_7__1923_ gnd vdd FILL
XFILL_1__3066_ gnd vdd FILL
XFILL_7__1854_ gnd vdd FILL
XFILL_1__2017_ gnd vdd FILL
XFILL_7__1785_ gnd vdd FILL
XFILL_7__3524_ gnd vdd FILL
XFILL_2__2830_ gnd vdd FILL
XFILL_7__3455_ gnd vdd FILL
XFILL_2__2761_ gnd vdd FILL
XFILL_1__2919_ gnd vdd FILL
XFILL_7__3386_ gnd vdd FILL
XFILL_5__2470_ gnd vdd FILL
XFILL_2__1712_ gnd vdd FILL
XFILL_7__2406_ gnd vdd FILL
XFILL_7__2337_ gnd vdd FILL
XFILL_2__2692_ gnd vdd FILL
XFILL_4__2628_ gnd vdd FILL
XFILL_4__2559_ gnd vdd FILL
XFILL_7_BUFX2_insert26 gnd vdd FILL
XFILL_7__2268_ gnd vdd FILL
XFILL_7_BUFX2_insert15 gnd vdd FILL
XFILL_7_BUFX2_insert59 gnd vdd FILL
XFILL_7_BUFX2_insert48 gnd vdd FILL
XFILL_5__3022_ gnd vdd FILL
XFILL_7__2199_ gnd vdd FILL
XFILL_8__1963_ gnd vdd FILL
XFILL_2__3175_ gnd vdd FILL
XFILL_0__2190_ gnd vdd FILL
XFILL_2__2126_ gnd vdd FILL
XFILL_8__1894_ gnd vdd FILL
XFILL_2__2057_ gnd vdd FILL
XFILL_3__2870_ gnd vdd FILL
XFILL_5__2806_ gnd vdd FILL
XFILL_8__3564_ gnd vdd FILL
XFILL183450x101550 gnd vdd FILL
XFILL_8__3495_ gnd vdd FILL
XFILL_3__1821_ gnd vdd FILL
XFILL_8__2515_ gnd vdd FILL
X_3370_ _3578_/Q _3568_/Q _3372_/A vdd gnd XOR2X1
XFILL_2__2959_ gnd vdd FILL
XFILL_8__2446_ gnd vdd FILL
XFILL_3__1752_ gnd vdd FILL
XFILL_5__2737_ gnd vdd FILL
XFILL_0__1974_ gnd vdd FILL
X_2321_ _2321_/A _2321_/B _2321_/C _2324_/B vdd gnd NOR3X1
XFILL_8__2377_ gnd vdd FILL
XFILL_5__2668_ gnd vdd FILL
X_2252_ _2932_/B _2252_/B _2274_/C _2306_/C vdd gnd AOI21X1
XFILL_5__2599_ gnd vdd FILL
XFILL_6__3200_ gnd vdd FILL
XFILL_6__3131_ gnd vdd FILL
XFILL_3__3422_ gnd vdd FILL
X_2183_ _2307_/B _2305_/A _2184_/C vdd gnd OR2X2
XFILL_6__3062_ gnd vdd FILL
XFILL_3__2304_ gnd vdd FILL
XFILL_6__2013_ gnd vdd FILL
XFILL_0__2526_ gnd vdd FILL
XFILL_3__2235_ gnd vdd FILL
XFILL_3__2166_ gnd vdd FILL
XFILL_0__2457_ gnd vdd FILL
XFILL_0__2388_ gnd vdd FILL
XFILL_6__2915_ gnd vdd FILL
XFILL_3__2097_ gnd vdd FILL
X_1967_ _3321_/Q _3029_/B _1968_/B vdd gnd NAND2X1
XFILL_6__2846_ gnd vdd FILL
XFILL_4__1930_ gnd vdd FILL
XFILL_0__3009_ gnd vdd FILL
X_1898_ _1898_/A _1898_/B _1902_/C vdd gnd NOR2X1
XFILL_4__1861_ gnd vdd FILL
XFILL_4__3600_ gnd vdd FILL
XFILL_6__2777_ gnd vdd FILL
XFILL_4__3531_ gnd vdd FILL
X_3568_ _3568_/D vdd _3578_/R _3577_/CLK _3568_/Q vdd gnd DFFSR
XFILL_3__2999_ gnd vdd FILL
XFILL_4__1792_ gnd vdd FILL
XFILL_6__1728_ gnd vdd FILL
X_2519_ _3356_/Q _2538_/B _2519_/C _2523_/B vdd gnd AOI21X1
XFILL_4__3462_ gnd vdd FILL
X_3499_ _3524_/A _3499_/B _3502_/A vdd gnd NAND2X1
XFILL_7__3171_ gnd vdd FILL
XFILL_1__2704_ gnd vdd FILL
XFILL_4__3393_ gnd vdd FILL
XFILL_7__2122_ gnd vdd FILL
XFILL_4__2413_ gnd vdd FILL
XFILL_4__2344_ gnd vdd FILL
XFILL_1__2635_ gnd vdd FILL
XFILL_7__2053_ gnd vdd FILL
XFILL_1__2566_ gnd vdd FILL
XFILL_4__2275_ gnd vdd FILL
XFILL_1__2497_ gnd vdd FILL
XFILL_7__2955_ gnd vdd FILL
XFILL_1__3118_ gnd vdd FILL
XFILL_7__1906_ gnd vdd FILL
XFILL_5__1970_ gnd vdd FILL
XFILL_7__2886_ gnd vdd FILL
XFILL_1__3049_ gnd vdd FILL
XFILL_7__1837_ gnd vdd FILL
XFILL_7__1768_ gnd vdd FILL
XFILL_7__3507_ gnd vdd FILL
XFILL_2__2813_ gnd vdd FILL
XFILL_8__2300_ gnd vdd FILL
XFILL_7__1699_ gnd vdd FILL
XFILL_7__3438_ gnd vdd FILL
XFILL_8__2231_ gnd vdd FILL
XFILL_5__2522_ gnd vdd FILL
XFILL_5__2453_ gnd vdd FILL
XFILL_2__2744_ gnd vdd FILL
XFILL_8__2162_ gnd vdd FILL
XFILL_7__3369_ gnd vdd FILL
XFILL_2__2675_ gnd vdd FILL
XFILL_5__2384_ gnd vdd FILL
XFILL_0__1690_ gnd vdd FILL
XFILL_8__2093_ gnd vdd FILL
XFILL_0__2311_ gnd vdd FILL
XFILL_5__3005_ gnd vdd FILL
XFILL_3__2020_ gnd vdd FILL
XFILL_8__2995_ gnd vdd FILL
XFILL_2__3227_ gnd vdd FILL
X_2870_ _2887_/A _2870_/B _2871_/D vdd gnd NAND2X1
XFILL_8__1946_ gnd vdd FILL
XFILL183750x105450 gnd vdd FILL
XFILL_0__2242_ gnd vdd FILL
XFILL183450x74250 gnd vdd FILL
XFILL_2__3158_ gnd vdd FILL
X_1821_ _2627_/A _3189_/C _2985_/A _1831_/D _3442_/A vdd gnd OAI22X1
XFILL_0__2173_ gnd vdd FILL
XFILL_2__2109_ gnd vdd FILL
XFILL_2__3089_ gnd vdd FILL
XFILL_8__1877_ gnd vdd FILL
XFILL_6__2700_ gnd vdd FILL
XFILL_3__2922_ gnd vdd FILL
X_1752_ _2594_/A _2594_/B _3166_/D vdd gnd NOR2X1
XFILL_3_BUFX2_insert13 gnd vdd FILL
XFILL_8__3547_ gnd vdd FILL
XFILL_3__2853_ gnd vdd FILL
XFILL_3_BUFX2_insert24 gnd vdd FILL
XFILL_9__2340_ gnd vdd FILL
XFILL_3_BUFX2_insert46 gnd vdd FILL
XFILL_6__2631_ gnd vdd FILL
XFILL_3_BUFX2_insert57 gnd vdd FILL
X_3422_ _3453_/B _3428_/A _3425_/B vdd gnd AND2X2
XFILL_3_BUFX2_insert79 gnd vdd FILL
XFILL_3_BUFX2_insert68 gnd vdd FILL
XFILL_3__1804_ gnd vdd FILL
XFILL_6__2562_ gnd vdd FILL
XFILL_8__3478_ gnd vdd FILL
XFILL_3__2784_ gnd vdd FILL
XFILL_6__2493_ gnd vdd FILL
X_3353_ _3353_/D vdd _3353_/R _3578_/CLK _3353_/Q vdd gnd DFFSR
XFILL_3__1735_ gnd vdd FILL
XFILL_8__2429_ gnd vdd FILL
XFILL_0__1957_ gnd vdd FILL
X_3284_ _3284_/D vdd _3313_/R _3284_/CLK _3284_/Q vdd gnd DFFSR
X_2304_ _2304_/A _2304_/B _2304_/C _2326_/B vdd gnd NAND3X1
XFILL_3__3405_ gnd vdd FILL
X_2235_ _2786_/A _3163_/A _2235_/C _2245_/A vdd gnd NAND3X1
XFILL_0__1888_ gnd vdd FILL
XFILL_6__3114_ gnd vdd FILL
X_2166_ _2298_/A _3077_/C _2166_/C _2298_/D _2335_/B vdd gnd AOI22X1
XFILL_1__2420_ gnd vdd FILL
XFILL_6__3045_ gnd vdd FILL
XFILL_0__3558_ gnd vdd FILL
XFILL_1__2351_ gnd vdd FILL
X_2097_ _2349_/A _2097_/B _2098_/A vdd gnd NOR2X1
XFILL_4__2060_ gnd vdd FILL
XFILL_0__3489_ gnd vdd FILL
XFILL_1__2282_ gnd vdd FILL
XFILL_3__2218_ gnd vdd FILL
XFILL_0__2509_ gnd vdd FILL
XFILL_3__3198_ gnd vdd FILL
XFILL_3__2149_ gnd vdd FILL
XFILL_7__2740_ gnd vdd FILL
XFILL_4__2962_ gnd vdd FILL
X_2999_ _3011_/B _2999_/B _3269_/Q _2999_/D _3005_/A vdd gnd OAI22X1
XFILL_9__3587_ gnd vdd FILL
XFILL_4__1913_ gnd vdd FILL
XFILL_7__2671_ gnd vdd FILL
XFILL_6__2829_ gnd vdd FILL
XFILL_4__2893_ gnd vdd FILL
XFILL_4__1844_ gnd vdd FILL
XFILL_4__1775_ gnd vdd FILL
XFILL_4__3514_ gnd vdd FILL
XFILL_1__1997_ gnd vdd FILL
XFILL_4__3445_ gnd vdd FILL
XFILL_7__3223_ gnd vdd FILL
XFILL_2__2460_ gnd vdd FILL
XFILL_7__3154_ gnd vdd FILL
XFILL_4__3376_ gnd vdd FILL
XFILL_7__3085_ gnd vdd FILL
XFILL_1__2618_ gnd vdd FILL
XFILL_7__2105_ gnd vdd FILL
XFILL_7__2036_ gnd vdd FILL
XFILL_4__2327_ gnd vdd FILL
XFILL_1__3598_ gnd vdd FILL
XFILL_2__2391_ gnd vdd FILL
XFILL_4__2258_ gnd vdd FILL
XFILL_1__2549_ gnd vdd FILL
XFILL_4__2189_ gnd vdd FILL
XFILL_2__3012_ gnd vdd FILL
XFILL_8__1800_ gnd vdd FILL
XFILL_7_CLKBUF1_insert38 gnd vdd FILL
XFILL_8__2780_ gnd vdd FILL
XFILL_7__2938_ gnd vdd FILL
XFILL_8__1731_ gnd vdd FILL
XFILL_7__2869_ gnd vdd FILL
XFILL_5__1953_ gnd vdd FILL
XFILL_8__3401_ gnd vdd FILL
XFILL_5__1884_ gnd vdd FILL
XFILL_5_CLKBUF1_insert31 gnd vdd FILL
XFILL_5__3554_ gnd vdd FILL
XFILL_0__2860_ gnd vdd FILL
XFILL_5__2505_ gnd vdd FILL
XFILL_5__3485_ gnd vdd FILL
XFILL_0__2791_ gnd vdd FILL
XFILL_8__2214_ gnd vdd FILL
XFILL_8__3194_ gnd vdd FILL
XFILL_2__2727_ gnd vdd FILL
XFILL_0__1811_ gnd vdd FILL
XFILL_8__2145_ gnd vdd FILL
XFILL_0__1742_ gnd vdd FILL
XFILL_5__2436_ gnd vdd FILL
X_2020_ _2845_/A _2261_/B vdd gnd INVX1
XFILL_5__2367_ gnd vdd FILL
XFILL_2__2658_ gnd vdd FILL
XFILL_0__3412_ gnd vdd FILL
XFILL_8__2076_ gnd vdd FILL
XFILL_2__2589_ gnd vdd FILL
XFILL_3__3121_ gnd vdd FILL
XFILL183750x117150 gnd vdd FILL
XFILL_5__2298_ gnd vdd FILL
XFILL_3__3052_ gnd vdd FILL
XFILL_9__1840_ gnd vdd FILL
X_2922_ _2922_/A _2922_/B _2922_/C _2923_/B vdd gnd OAI21X1
XFILL_3__2003_ gnd vdd FILL
XFILL_8__2978_ gnd vdd FILL
XFILL_0__2225_ gnd vdd FILL
X_2853_ _2853_/A _2909_/C _2855_/C vdd gnd NAND2X1
XFILL_8__1929_ gnd vdd FILL
XFILL_6__1993_ gnd vdd FILL
X_2784_ _2910_/B _2933_/A vdd gnd INVX2
XFILL_0__2156_ gnd vdd FILL
X_1804_ _2602_/B _2091_/B _2701_/B _1805_/C vdd gnd OAI21X1
XFILL_0__2087_ gnd vdd FILL
X_1735_ _3233_/Q _1762_/B vdd gnd INVX1
XFILL_3__2905_ gnd vdd FILL
XFILL_1__1920_ gnd vdd FILL
XFILL_6__2614_ gnd vdd FILL
XFILL_3__2836_ gnd vdd FILL
XFILL_6__3594_ gnd vdd FILL
X_3405_ _3453_/B _3411_/A _3408_/B vdd gnd AND2X2
XFILL_1__1851_ gnd vdd FILL
XFILL_6__2545_ gnd vdd FILL
XFILL_3__2767_ gnd vdd FILL
X_3336_ _3336_/D vdd _3347_/R _3576_/CLK _3336_/Q vdd gnd DFFSR
XFILL_0__2989_ gnd vdd FILL
XFILL_6__2476_ gnd vdd FILL
XFILL_3__1718_ gnd vdd FILL
XFILL_1__1782_ gnd vdd FILL
XFILL_1__3521_ gnd vdd FILL
XFILL_3__2698_ gnd vdd FILL
X_3267_ _3267_/D vdd _3313_/R _3284_/CLK _3267_/Q vdd gnd DFFSR
XFILL_4__3230_ gnd vdd FILL
XFILL_1__3452_ gnd vdd FILL
X_2218_ _2299_/A _3183_/B _2367_/B vdd gnd NOR2X1
X_3198_ _3214_/A _3214_/B _3198_/Y vdd gnd NOR2X1
XFILL_4__3161_ gnd vdd FILL
XFILL_4__2112_ gnd vdd FILL
XFILL_1__3383_ gnd vdd FILL
XFILL_1__2403_ gnd vdd FILL
X_2149_ _2278_/A _3177_/B _2150_/C vdd gnd NAND2X1
XFILL_6__3028_ gnd vdd FILL
XFILL_4__3092_ gnd vdd FILL
XFILL_1__2334_ gnd vdd FILL
XFILL_4__2043_ gnd vdd FILL
XFILL_1__2265_ gnd vdd FILL
XFILL_1__2196_ gnd vdd FILL
XFILL_7__2723_ gnd vdd FILL
XFILL_4__2945_ gnd vdd FILL
XFILL_7__2654_ gnd vdd FILL
XFILL_4__2876_ gnd vdd FILL
XFILL_2__1960_ gnd vdd FILL
XFILL_4__1827_ gnd vdd FILL
XFILL_2__1891_ gnd vdd FILL
XFILL_7__2585_ gnd vdd FILL
XFILL_2__3561_ gnd vdd FILL
XFILL_4__1758_ gnd vdd FILL
XFILL_4__1689_ gnd vdd FILL
XFILL_7__3206_ gnd vdd FILL
XFILL_2__2512_ gnd vdd FILL
XFILL_2__3492_ gnd vdd FILL
XFILL_4__3428_ gnd vdd FILL
XFILL_5__2221_ gnd vdd FILL
XFILL_7__3137_ gnd vdd FILL
XFILL_5__2152_ gnd vdd FILL
XFILL_2__2443_ gnd vdd FILL
XFILL_7__3068_ gnd vdd FILL
XFILL_2__2374_ gnd vdd FILL
XFILL_5__2083_ gnd vdd FILL
XFILL_8__2901_ gnd vdd FILL
XFILL_7__2019_ gnd vdd FILL
XFILL_8__2832_ gnd vdd FILL
XFILL_8__2763_ gnd vdd FILL
XFILL_0__2010_ gnd vdd FILL
XFILL_5__2985_ gnd vdd FILL
XFILL_8__1714_ gnd vdd FILL
XFILL_5__1936_ gnd vdd FILL
XFILL_8__2694_ gnd vdd FILL
XFILL_5__1867_ gnd vdd FILL
XFILL_0__2912_ gnd vdd FILL
XFILL_3__2621_ gnd vdd FILL
XFILL_2_BUFX2_insert3 gnd vdd FILL
XFILL_5__1798_ gnd vdd FILL
XFILL_0__2843_ gnd vdd FILL
XFILL_5__3537_ gnd vdd FILL
XFILL_6__2330_ gnd vdd FILL
X_3121_ _3121_/A _3125_/B _3336_/Q _3122_/C vdd gnd OAI21X1
XFILL_5__3468_ gnd vdd FILL
XFILL_6__2261_ gnd vdd FILL
XFILL_3__2552_ gnd vdd FILL
XFILL_5__2419_ gnd vdd FILL
XFILL_3__2483_ gnd vdd FILL
XFILL_0__2774_ gnd vdd FILL
XFILL_8__3177_ gnd vdd FILL
XFILL_5__3399_ gnd vdd FILL
X_3052_ _3292_/D _3077_/C _3052_/C _3052_/D _3133_/A vdd gnd AOI22X1
XFILL_8__2128_ gnd vdd FILL
XFILL_6__2192_ gnd vdd FILL
XFILL_0__1725_ gnd vdd FILL
X_2003_ _2249_/A _2932_/A _2824_/A vdd gnd NAND2X1
XFILL_8__2059_ gnd vdd FILL
XFILL_3__3104_ gnd vdd FILL
XFILL_6_BUFX2_insert61 gnd vdd FILL
XFILL_6_BUFX2_insert50 gnd vdd FILL
XFILL_6_BUFX2_insert72 gnd vdd FILL
XFILL_6_BUFX2_insert94 gnd vdd FILL
XFILL_3__3035_ gnd vdd FILL
XFILL_6_BUFX2_insert83 gnd vdd FILL
X_2905_ _2905_/A _2907_/B vdd gnd INVX1
XFILL_1__2050_ gnd vdd FILL
XFILL_6__1976_ gnd vdd FILL
X_2836_ _2860_/A _2865_/D _2919_/B _2862_/A vdd gnd AOI21X1
XFILL_0__2208_ gnd vdd FILL
XFILL_0__3188_ gnd vdd FILL
XFILL_0__2139_ gnd vdd FILL
XFILL_4__2730_ gnd vdd FILL
X_2767_ _2767_/A _2767_/B _2767_/C _2769_/A vdd gnd NAND3X1
XFILL_1__2952_ gnd vdd FILL
X_1718_ _3233_/Q _1756_/A _1888_/B vdd gnd NOR2X1
X_2698_ _2733_/B _2706_/A vdd gnd INVX1
XFILL_4__2661_ gnd vdd FILL
XFILL_1__2883_ gnd vdd FILL
XFILL_7__2370_ gnd vdd FILL
XFILL_1__1903_ gnd vdd FILL
XFILL_3__2819_ gnd vdd FILL
XFILL_6__2528_ gnd vdd FILL
XFILL_1__1834_ gnd vdd FILL
XFILL_4__2592_ gnd vdd FILL
XFILL_9__2237_ gnd vdd FILL
X_3319_ _3319_/D vdd _3353_/R _3577_/CLK _3319_/Q vdd gnd DFFSR
XFILL_6__2459_ gnd vdd FILL
XFILL_1__1765_ gnd vdd FILL
XFILL_1__3504_ gnd vdd FILL
XFILL_1__1696_ gnd vdd FILL
XFILL_4__3213_ gnd vdd FILL
XFILL_1__3435_ gnd vdd FILL
XFILL_5_BUFX2_insert7 gnd vdd FILL
XFILL_4__3144_ gnd vdd FILL
XFILL_4__3075_ gnd vdd FILL
XFILL_1__3366_ gnd vdd FILL
XFILL_4__2026_ gnd vdd FILL
XFILL_1__2317_ gnd vdd FILL
XFILL_2__2090_ gnd vdd FILL
XFILL_1__2248_ gnd vdd FILL
XFILL_1__2179_ gnd vdd FILL
XFILL_7__2706_ gnd vdd FILL
XFILL_5__2770_ gnd vdd FILL
XFILL_4__2928_ gnd vdd FILL
XFILL_2__2992_ gnd vdd FILL
XFILL_5__1721_ gnd vdd FILL
XFILL_7__2637_ gnd vdd FILL
XFILL_2__1943_ gnd vdd FILL
XFILL_4__2859_ gnd vdd FILL
XFILL_7__2568_ gnd vdd FILL
XFILL_2__1874_ gnd vdd FILL
XFILL_8__3100_ gnd vdd FILL
XFILL_7__2499_ gnd vdd FILL
XFILL_2__3544_ gnd vdd FILL
XFILL_8__3031_ gnd vdd FILL
XFILL_2__3475_ gnd vdd FILL
XFILL_5__2204_ gnd vdd FILL
XFILL_2__2426_ gnd vdd FILL
XFILL_0__2490_ gnd vdd FILL
XFILL_5__3184_ gnd vdd FILL
XFILL_5__2135_ gnd vdd FILL
XFILL_5__2066_ gnd vdd FILL
XFILL_2__2357_ gnd vdd FILL
XFILL_2__2288_ gnd vdd FILL
XFILL_0__3111_ gnd vdd FILL
XFILL_8__2815_ gnd vdd FILL
XFILL_0__3042_ gnd vdd FILL
XFILL_6__1830_ gnd vdd FILL
XFILL_8__2746_ gnd vdd FILL
XFILL_6__3500_ gnd vdd FILL
XFILL_5__2968_ gnd vdd FILL
XFILL_6__1761_ gnd vdd FILL
X_2621_ _2767_/A _2621_/B _2621_/C _2621_/D _3240_/D vdd gnd OAI22X1
XFILL_8__2677_ gnd vdd FILL
XFILL_3__1983_ gnd vdd FILL
XFILL_5__2899_ gnd vdd FILL
XFILL_5__1919_ gnd vdd FILL
XFILL_6__1692_ gnd vdd FILL
X_2552_ _2744_/B _2574_/B _2552_/C _3583_/A vdd gnd OAI21X1
XFILL_6__3431_ gnd vdd FILL
X_2483_ _2641_/B _2574_/B _2483_/C _2484_/C vdd gnd OAI21X1
XFILL_6__2313_ gnd vdd FILL
XFILL_3__3584_ gnd vdd FILL
XFILL_3__2604_ gnd vdd FILL
XFILL_0__2826_ gnd vdd FILL
XFILL_3__2535_ gnd vdd FILL
XFILL_8__3229_ gnd vdd FILL
X_3104_ _3139_/A _3108_/B _3104_/C _3328_/D vdd gnd OAI21X1
XFILL_6__2244_ gnd vdd FILL
XFILL_0__2757_ gnd vdd FILL
X_3035_ _3339_/Q _3035_/B _3085_/B vdd gnd NAND2X1
XFILL_0__1708_ gnd vdd FILL
XFILL_3__2466_ gnd vdd FILL
XFILL_6__2175_ gnd vdd FILL
XFILL_3__2397_ gnd vdd FILL
XFILL_0__2688_ gnd vdd FILL
XFILL_1__3220_ gnd vdd FILL
XFILL_1__3151_ gnd vdd FILL
XFILL_1__3082_ gnd vdd FILL
XFILL_7__1870_ gnd vdd FILL
XFILL_3__3018_ gnd vdd FILL
XFILL_1__2102_ gnd vdd FILL
XFILL_1__2033_ gnd vdd FILL
XFILL_9__1737_ gnd vdd FILL
X_2819_ _2932_/B _2920_/A _2927_/B vdd gnd NOR2X1
XFILL_6__1959_ gnd vdd FILL
XFILL_7__3540_ gnd vdd FILL
XFILL_7__3471_ gnd vdd FILL
XFILL_7__2422_ gnd vdd FILL
XFILL_4__2713_ gnd vdd FILL
XFILL_1__2935_ gnd vdd FILL
XFILL_4__2644_ gnd vdd FILL
XFILL_1__2866_ gnd vdd FILL
XFILL_7__2353_ gnd vdd FILL
XFILL_2_BUFX2_insert81 gnd vdd FILL
XFILL_2_BUFX2_insert70 gnd vdd FILL
XFILL_2_BUFX2_insert92 gnd vdd FILL
XFILL_1__2797_ gnd vdd FILL
XFILL_4__2575_ gnd vdd FILL
XFILL_7__2284_ gnd vdd FILL
XFILL_1__1817_ gnd vdd FILL
XFILL_1__1748_ gnd vdd FILL
XFILL_4__3127_ gnd vdd FILL
XFILL_1__3418_ gnd vdd FILL
XFILL_2__2211_ gnd vdd FILL
XFILL_2__3191_ gnd vdd FILL
XFILL_2__2142_ gnd vdd FILL
XFILL_4__3058_ gnd vdd FILL
XFILL_2__2073_ gnd vdd FILL
XFILL_8__2600_ gnd vdd FILL
XFILL_4__2009_ gnd vdd FILL
XFILL_7__1999_ gnd vdd FILL
XFILL_5__2822_ gnd vdd FILL
XFILL_8__3580_ gnd vdd FILL
XFILL_8__2531_ gnd vdd FILL
XFILL_2_CLKBUF1_insert28 gnd vdd FILL
XFILL_8__2462_ gnd vdd FILL
XFILL_5__2753_ gnd vdd FILL
XFILL_2__2975_ gnd vdd FILL
XFILL_5__1704_ gnd vdd FILL
XFILL_5__2684_ gnd vdd FILL
XFILL_2__1926_ gnd vdd FILL
XFILL_8__2393_ gnd vdd FILL
XFILL_0__1990_ gnd vdd FILL
XFILL_2__1857_ gnd vdd FILL
XFILL_8__3014_ gnd vdd FILL
XFILL_0_CLKBUF1_insert32 gnd vdd FILL
XFILL_0__3591_ gnd vdd FILL
XFILL_3__2320_ gnd vdd FILL
XFILL_0__2611_ gnd vdd FILL
XFILL_2__1788_ gnd vdd FILL
XFILL_2__3527_ gnd vdd FILL
XFILL_0__2542_ gnd vdd FILL
XFILL_2__3458_ gnd vdd FILL
XFILL_3__2251_ gnd vdd FILL
XFILL_2__3389_ gnd vdd FILL
XFILL_3__2182_ gnd vdd FILL
XFILL_0__2473_ gnd vdd FILL
XFILL_5__3167_ gnd vdd FILL
XFILL_2__2409_ gnd vdd FILL
XFILL_5__3098_ gnd vdd FILL
XFILL_5__2118_ gnd vdd FILL
XFILL_6__2931_ gnd vdd FILL
XFILL_5__2049_ gnd vdd FILL
X_1983_ _2571_/A _2771_/C vdd gnd INVX1
XFILL_6__2862_ gnd vdd FILL
XFILL_6__2793_ gnd vdd FILL
XFILL_0__3025_ gnd vdd FILL
XFILL_8__2729_ gnd vdd FILL
XFILL_6__1813_ gnd vdd FILL
XFILL_6__1744_ gnd vdd FILL
X_2604_ _2604_/A _2605_/C vdd gnd INVX1
XFILL_3__1966_ gnd vdd FILL
X_3584_ _3584_/A AB[13] vdd gnd BUFX2
XFILL_6__3414_ gnd vdd FILL
X_2535_ _2565_/A _3292_/D _2535_/C _2536_/C vdd gnd AOI21X1
X_2466_ _2466_/A _2466_/B _2467_/C vdd gnd AND2X2
XFILL_3__1897_ gnd vdd FILL
XFILL_1__2720_ gnd vdd FILL
XFILL_1__2651_ gnd vdd FILL
XFILL_4__2360_ gnd vdd FILL
XFILL_0__2809_ gnd vdd FILL
X_2397_ _3572_/Q _2427_/B _2397_/C _2398_/B vdd gnd AOI21X1
XFILL_3__3498_ gnd vdd FILL
XFILL_6__2227_ gnd vdd FILL
XFILL_3__2518_ gnd vdd FILL
XFILL_1__2582_ gnd vdd FILL
XFILL_4__2291_ gnd vdd FILL
XFILL_3__2449_ gnd vdd FILL
X_3018_ _3313_/Q _3019_/A _3019_/C vdd gnd NAND2X1
XFILL_6__2158_ gnd vdd FILL
XFILL_7__2971_ gnd vdd FILL
XFILL_6__2089_ gnd vdd FILL
XFILL_1__3203_ gnd vdd FILL
XFILL_1__3134_ gnd vdd FILL
XFILL_7__1922_ gnd vdd FILL
XFILL_1__3065_ gnd vdd FILL
XFILL_7__1853_ gnd vdd FILL
XFILL_1__2016_ gnd vdd FILL
XFILL_7__1784_ gnd vdd FILL
XFILL_7__3523_ gnd vdd FILL
XFILL_7__3454_ gnd vdd FILL
XFILL_2__2760_ gnd vdd FILL
XFILL_1__2918_ gnd vdd FILL
XFILL_7__3385_ gnd vdd FILL
XFILL_7__2405_ gnd vdd FILL
XFILL_2__1711_ gnd vdd FILL
XFILL_2__2691_ gnd vdd FILL
XFILL_7__2336_ gnd vdd FILL
XFILL_4__2627_ gnd vdd FILL
XFILL_1__2849_ gnd vdd FILL
XFILL_4__2558_ gnd vdd FILL
XFILL_7__2267_ gnd vdd FILL
XFILL_7_BUFX2_insert27 gnd vdd FILL
XFILL_7_BUFX2_insert16 gnd vdd FILL
XFILL_7_BUFX2_insert49 gnd vdd FILL
XFILL_4__2489_ gnd vdd FILL
XFILL_5__3021_ gnd vdd FILL
XFILL_7__2198_ gnd vdd FILL
XFILL_8__1962_ gnd vdd FILL
XFILL_2__3174_ gnd vdd FILL
XFILL_2__2125_ gnd vdd FILL
XFILL_8__1893_ gnd vdd FILL
XFILL_2__2056_ gnd vdd FILL
XFILL_8__3563_ gnd vdd FILL
XFILL_5__2805_ gnd vdd FILL
XFILL_8__2514_ gnd vdd FILL
XFILL_8__3494_ gnd vdd FILL
XFILL_3__1820_ gnd vdd FILL
XFILL_5__2736_ gnd vdd FILL
XFILL_2__2958_ gnd vdd FILL
XFILL_3__1751_ gnd vdd FILL
XFILL_8__2445_ gnd vdd FILL
XFILL_0__1973_ gnd vdd FILL
X_2320_ _2332_/B _2320_/B _2320_/C _2321_/A vdd gnd NAND3X1
XFILL_8__2376_ gnd vdd FILL
XFILL_5__2667_ gnd vdd FILL
XFILL_2__1909_ gnd vdd FILL
XFILL_2__2889_ gnd vdd FILL
X_2251_ _2823_/B _2902_/A _2928_/B _2274_/C vdd gnd OAI21X1
XFILL_5__2598_ gnd vdd FILL
XFILL_6__3130_ gnd vdd FILL
XFILL_3__3421_ gnd vdd FILL
X_2182_ _2311_/A _2853_/A _2307_/B vdd gnd NAND2X1
XFILL_6__3061_ gnd vdd FILL
XFILL_3__2303_ gnd vdd FILL
XFILL_6__2012_ gnd vdd FILL
XFILL_0__2525_ gnd vdd FILL
XFILL_5__3219_ gnd vdd FILL
XFILL_3__2234_ gnd vdd FILL
XFILL_0__2456_ gnd vdd FILL
XFILL_3__2165_ gnd vdd FILL
XFILL_0__2387_ gnd vdd FILL
XFILL_3__2096_ gnd vdd FILL
XFILL_6__2914_ gnd vdd FILL
X_1966_ _3337_/Q _3110_/A _3127_/B _3346_/Q _1968_/C vdd gnd AOI22X1
XFILL_6__2845_ gnd vdd FILL
XFILL_4__1860_ gnd vdd FILL
XFILL_0__3008_ gnd vdd FILL
X_1897_ _3188_/A _3185_/A _1898_/B vdd gnd NAND2X1
XFILL_6__2776_ gnd vdd FILL
X_3567_ _3567_/D vdd _3578_/R _3576_/CLK _3567_/Q vdd gnd DFFSR
XFILL_4__3530_ gnd vdd FILL
XFILL_3__2998_ gnd vdd FILL
XFILL_4__1791_ gnd vdd FILL
XFILL_6__1727_ gnd vdd FILL
XFILL_3__1949_ gnd vdd FILL
X_2518_ _2697_/B _2574_/B _3216_/A vdd gnd NOR2X1
X_3498_ _3498_/A _3548_/B _3498_/C _3499_/B vdd gnd NAND3X1
XFILL_9__3106_ gnd vdd FILL
XFILL_4__3461_ gnd vdd FILL
XFILL_1__2703_ gnd vdd FILL
XFILL_7__3170_ gnd vdd FILL
XFILL_4__3392_ gnd vdd FILL
XFILL_4__2412_ gnd vdd FILL
XFILL_7__2121_ gnd vdd FILL
X_2449_ _2717_/B _2449_/B _2449_/C _2563_/A vdd gnd NAND3X1
XFILL_4__2343_ gnd vdd FILL
XFILL_1__2634_ gnd vdd FILL
XFILL_7__2052_ gnd vdd FILL
XFILL_1__2565_ gnd vdd FILL
XFILL_4__2274_ gnd vdd FILL
XFILL_1__2496_ gnd vdd FILL
XFILL_7__2954_ gnd vdd FILL
XFILL_1__3117_ gnd vdd FILL
XFILL_7__2885_ gnd vdd FILL
XFILL_7__1905_ gnd vdd FILL
XFILL_1__3048_ gnd vdd FILL
XFILL_7__1836_ gnd vdd FILL
XFILL_7__1767_ gnd vdd FILL
XFILL_2__2812_ gnd vdd FILL
XFILL_7__3506_ gnd vdd FILL
XFILL_4__1989_ gnd vdd FILL
XFILL_7__1698_ gnd vdd FILL
XFILL_7__3437_ gnd vdd FILL
XFILL_5__2521_ gnd vdd FILL
XFILL_8__2230_ gnd vdd FILL
XFILL_5__2452_ gnd vdd FILL
XFILL_2__2743_ gnd vdd FILL
XFILL_8__2161_ gnd vdd FILL
XFILL_7__3368_ gnd vdd FILL
XFILL_2__2674_ gnd vdd FILL
XFILL_5__2383_ gnd vdd FILL
XFILL_7__2319_ gnd vdd FILL
XFILL_8__2092_ gnd vdd FILL
XFILL_0__2310_ gnd vdd FILL
XFILL_5__3004_ gnd vdd FILL
XFILL_8__2994_ gnd vdd FILL
XFILL_2__3226_ gnd vdd FILL
XFILL_0__2241_ gnd vdd FILL
XFILL_8__1945_ gnd vdd FILL
XFILL_2__3157_ gnd vdd FILL
XFILL_0__2172_ gnd vdd FILL
X_1820_ _3241_/Q _2627_/A vdd gnd INVX1
XFILL_2__2108_ gnd vdd FILL
XFILL_8__1876_ gnd vdd FILL
XFILL_2__3088_ gnd vdd FILL
XFILL_3__2921_ gnd vdd FILL
XFILL_2__2039_ gnd vdd FILL
X_1751_ _1751_/A _1751_/B _1751_/C _1778_/A vdd gnd OAI21X1
XFILL_6__2630_ gnd vdd FILL
XFILL_8__3546_ gnd vdd FILL
XFILL_3__2852_ gnd vdd FILL
XFILL_3_BUFX2_insert25 gnd vdd FILL
XFILL_3_BUFX2_insert47 gnd vdd FILL
XFILL_3_BUFX2_insert14 gnd vdd FILL
XFILL_8__3477_ gnd vdd FILL
XFILL_3_BUFX2_insert58 gnd vdd FILL
X_3421_ _3521_/A _3421_/B _3426_/C vdd gnd NAND2X1
XFILL_3__1803_ gnd vdd FILL
XFILL_6__2561_ gnd vdd FILL
XFILL_3_BUFX2_insert69 gnd vdd FILL
XFILL_3__2783_ gnd vdd FILL
XFILL_8__2428_ gnd vdd FILL
XFILL_6__2492_ gnd vdd FILL
X_3352_ _3352_/D vdd _3355_/R _3355_/CLK _3352_/Q vdd gnd DFFSR
XFILL_5__2719_ gnd vdd FILL
X_2303_ _2303_/A _2303_/B _2304_/B vdd gnd NOR2X1
XFILL_3__1734_ gnd vdd FILL
XFILL_0__1956_ gnd vdd FILL
XFILL_8__2359_ gnd vdd FILL
X_3283_ _3283_/D vdd _3289_/R _3307_/CLK _3283_/Q vdd gnd DFFSR
XFILL_3__3404_ gnd vdd FILL
XFILL_0__1887_ gnd vdd FILL
X_2234_ _2441_/C _2234_/B _2234_/C _2246_/B vdd gnd NAND3X1
XFILL_6__3113_ gnd vdd FILL
X_2165_ _2792_/C _2312_/A _2166_/C vdd gnd NOR2X1
XFILL_6__3044_ gnd vdd FILL
XFILL_1__2350_ gnd vdd FILL
XFILL_0__3557_ gnd vdd FILL
X_2096_ _2294_/A _3158_/A _2096_/C _2097_/B vdd gnd OAI21X1
XFILL_0__3488_ gnd vdd FILL
XFILL_3__2217_ gnd vdd FILL
XFILL_1__2281_ gnd vdd FILL
XFILL_0__2508_ gnd vdd FILL
XFILL_3__3197_ gnd vdd FILL
XFILL_0__2439_ gnd vdd FILL
XFILL_3__2148_ gnd vdd FILL
XFILL_3__2079_ gnd vdd FILL
XFILL_4__2961_ gnd vdd FILL
X_2998_ _2998_/A _2998_/B _2998_/C _3311_/D vdd gnd OAI21X1
X_1949_ _3319_/Q _3029_/B _1950_/B vdd gnd NAND2X1
XFILL_4__1912_ gnd vdd FILL
XFILL_7__2670_ gnd vdd FILL
XFILL_6__2828_ gnd vdd FILL
XFILL_4__2892_ gnd vdd FILL
XFILL_4__1843_ gnd vdd FILL
XFILL_6__2759_ gnd vdd FILL
XFILL_4__1774_ gnd vdd FILL
XFILL_4__3513_ gnd vdd FILL
XFILL_9__2399_ gnd vdd FILL
XFILL_7__3222_ gnd vdd FILL
XFILL_1__1996_ gnd vdd FILL
XFILL_4__3444_ gnd vdd FILL
XFILL_7__3153_ gnd vdd FILL
XFILL_7__2104_ gnd vdd FILL
XFILL_4__3375_ gnd vdd FILL
XFILL_7__3084_ gnd vdd FILL
XFILL_1__2617_ gnd vdd FILL
XFILL_7__2035_ gnd vdd FILL
XFILL_4__2326_ gnd vdd FILL
XFILL_2__2390_ gnd vdd FILL
XFILL_1__3597_ gnd vdd FILL
XFILL_4__2257_ gnd vdd FILL
XFILL_1__2548_ gnd vdd FILL
XFILL_1__2479_ gnd vdd FILL
XFILL_4__2188_ gnd vdd FILL
XFILL_2__3011_ gnd vdd FILL
XFILL_7_CLKBUF1_insert28 gnd vdd FILL
XFILL_8__1730_ gnd vdd FILL
XFILL_7__2937_ gnd vdd FILL
XFILL_5__1952_ gnd vdd FILL
XFILL_7__2868_ gnd vdd FILL
XFILL_8__3400_ gnd vdd FILL
XFILL_7__2799_ gnd vdd FILL
XFILL_7__1819_ gnd vdd FILL
XFILL_5__1883_ gnd vdd FILL
XFILL_5_CLKBUF1_insert32 gnd vdd FILL
XFILL_5__3553_ gnd vdd FILL
XFILL_5__2504_ gnd vdd FILL
XFILL_5__3484_ gnd vdd FILL
XFILL_8__2213_ gnd vdd FILL
XFILL_0__2790_ gnd vdd FILL
XFILL_2__2726_ gnd vdd FILL
XFILL_8__3193_ gnd vdd FILL
XFILL_0__1810_ gnd vdd FILL
XFILL_8__2144_ gnd vdd FILL
XFILL_0__1741_ gnd vdd FILL
XFILL_5__2435_ gnd vdd FILL
XFILL_5__2366_ gnd vdd FILL
XFILL_2__2657_ gnd vdd FILL
XFILL_0__3411_ gnd vdd FILL
XFILL_8__2075_ gnd vdd FILL
XFILL_2__2588_ gnd vdd FILL
XFILL_3__3120_ gnd vdd FILL
XFILL_5__2297_ gnd vdd FILL
XFILL_3__3051_ gnd vdd FILL
X_2921_ _2921_/A _2932_/C _2935_/A _2922_/C vdd gnd AOI21X1
XFILL_3__2002_ gnd vdd FILL
XFILL_2__3209_ gnd vdd FILL
XFILL_8__2977_ gnd vdd FILL
XFILL_0__2224_ gnd vdd FILL
X_2852_ _2894_/A _2880_/A _2909_/C vdd gnd NOR2X1
XFILL_8__1928_ gnd vdd FILL
XFILL_6__1992_ gnd vdd FILL
XFILL_8__1859_ gnd vdd FILL
X_2783_ _3257_/Q _2786_/B vdd gnd INVX1
XFILL_0__2155_ gnd vdd FILL
X_1803_ _2442_/B _1803_/B _2091_/B vdd gnd NOR2X1
XFILL_3__2904_ gnd vdd FILL
XFILL_0__2086_ gnd vdd FILL
X_1734_ _2379_/A _1734_/Y vdd gnd INVX8
XFILL_8__3529_ gnd vdd FILL
XFILL_6__3593_ gnd vdd FILL
XFILL_6__2613_ gnd vdd FILL
XFILL_3__2835_ gnd vdd FILL
X_3404_ _3521_/A _3404_/B _3409_/C vdd gnd NAND2X1
XFILL_6__2544_ gnd vdd FILL
XFILL_3__2766_ gnd vdd FILL
XFILL_1__1850_ gnd vdd FILL
X_3335_ _3335_/D vdd _3345_/R _3576_/CLK _3335_/Q vdd gnd DFFSR
XFILL_0__2988_ gnd vdd FILL
XFILL_6__2475_ gnd vdd FILL
XFILL_3__1717_ gnd vdd FILL
XFILL_1__1781_ gnd vdd FILL
XFILL_0__1939_ gnd vdd FILL
XFILL_1__3520_ gnd vdd FILL
X_3266_ _3266_/D vdd _3282_/R _3313_/CLK _3266_/Q vdd gnd DFFSR
XFILL_3__2697_ gnd vdd FILL
X_2217_ _2885_/B _2932_/B _2797_/B vdd gnd NOR2X1
XFILL_1__3451_ gnd vdd FILL
X_3197_ _3197_/A _3197_/B _3197_/C _3214_/B vdd gnd OAI21X1
XFILL_4__3160_ gnd vdd FILL
XFILL_1__3382_ gnd vdd FILL
XFILL_1__2402_ gnd vdd FILL
X_2148_ _2717_/C _3177_/B vdd gnd INVX2
XFILL_4__2111_ gnd vdd FILL
X_2079_ _2915_/C _2931_/A _2902_/A vdd gnd NAND2X1
XFILL_4__3091_ gnd vdd FILL
XFILL_6__3027_ gnd vdd FILL
XFILL_1__2333_ gnd vdd FILL
XFILL_4__2042_ gnd vdd FILL
XFILL_1__2264_ gnd vdd FILL
XFILL_1__2195_ gnd vdd FILL
XFILL_9__1899_ gnd vdd FILL
XFILL_7__2722_ gnd vdd FILL
XFILL_4__2944_ gnd vdd FILL
XFILL_7__2653_ gnd vdd FILL
XFILL_4__2875_ gnd vdd FILL
XFILL_7__2584_ gnd vdd FILL
XFILL_2__1890_ gnd vdd FILL
XFILL_4__1826_ gnd vdd FILL
XFILL_2__3560_ gnd vdd FILL
XFILL_4__1757_ gnd vdd FILL
XFILL_1__1979_ gnd vdd FILL
XFILL_7__3205_ gnd vdd FILL
XFILL_2__2511_ gnd vdd FILL
XFILL_4__1688_ gnd vdd FILL
XFILL_2__3491_ gnd vdd FILL
XFILL_7__3136_ gnd vdd FILL
XFILL_4__3427_ gnd vdd FILL
XFILL_5__2220_ gnd vdd FILL
XFILL_5__2151_ gnd vdd FILL
XFILL_2__2442_ gnd vdd FILL
XFILL_4__2309_ gnd vdd FILL
XFILL_7__3067_ gnd vdd FILL
XFILL_2__2373_ gnd vdd FILL
XFILL_8__2900_ gnd vdd FILL
XFILL_7__2018_ gnd vdd FILL
XFILL_5__2082_ gnd vdd FILL
XFILL_8__2831_ gnd vdd FILL
XFILL_8__2762_ gnd vdd FILL
XFILL_5__2984_ gnd vdd FILL
XFILL_8__2693_ gnd vdd FILL
XFILL_8__1713_ gnd vdd FILL
XFILL_5__1935_ gnd vdd FILL
XFILL_5__1866_ gnd vdd FILL
XFILL_0__2911_ gnd vdd FILL
XFILL_3__2620_ gnd vdd FILL
XFILL_2_BUFX2_insert4 gnd vdd FILL
XFILL_5__1797_ gnd vdd FILL
XFILL_0__2842_ gnd vdd FILL
XFILL_5__3536_ gnd vdd FILL
X_3120_ _3137_/A _3126_/B _3120_/C _3335_/D vdd gnd OAI21X1
XFILL_5__3467_ gnd vdd FILL
XFILL_6__2260_ gnd vdd FILL
XFILL_3__2551_ gnd vdd FILL
XFILL_5__2418_ gnd vdd FILL
XFILL_3__2482_ gnd vdd FILL
XFILL_2__2709_ gnd vdd FILL
XFILL_0__2773_ gnd vdd FILL
XFILL_8__3176_ gnd vdd FILL
XFILL_5__3398_ gnd vdd FILL
XFILL_6__2191_ gnd vdd FILL
X_3051_ _3077_/C _3055_/A _3052_/C vdd gnd NOR2X1
XFILL_0__1724_ gnd vdd FILL
XFILL_8__2127_ gnd vdd FILL
X_2002_ _2025_/A _3290_/D _2002_/C _2932_/A vdd gnd OAI21X1
XFILL_5__2349_ gnd vdd FILL
XFILL_8__2058_ gnd vdd FILL
XFILL_3__3103_ gnd vdd FILL
XFILL_6_BUFX2_insert51 gnd vdd FILL
XFILL_6_BUFX2_insert62 gnd vdd FILL
XFILL_6_BUFX2_insert40 gnd vdd FILL
XFILL_6_BUFX2_insert95 gnd vdd FILL
XFILL_6_BUFX2_insert84 gnd vdd FILL
XFILL_3__3034_ gnd vdd FILL
XFILL_6_BUFX2_insert73 gnd vdd FILL
X_2904_ _2928_/B _2926_/B _2913_/C _2905_/A vdd gnd OAI21X1
X_2835_ _2835_/A _2835_/B _2860_/A vdd gnd NOR2X1
XFILL_6__1975_ gnd vdd FILL
XFILL_0__2207_ gnd vdd FILL
XFILL_0__3187_ gnd vdd FILL
XFILL_0__2138_ gnd vdd FILL
X_2766_ _2766_/A _2766_/B _2766_/C _2767_/C vdd gnd OAI21X1
XFILL_1__2951_ gnd vdd FILL
XFILL_0__2069_ gnd vdd FILL
X_1717_ _3234_/Q _1756_/A vdd gnd INVX1
X_2697_ _2767_/A _2697_/B _2697_/C _3247_/D vdd gnd OAI21X1
XFILL_4__2660_ gnd vdd FILL
XFILL_3__2818_ gnd vdd FILL
XFILL_1__2882_ gnd vdd FILL
XFILL_1__1902_ gnd vdd FILL
XFILL_6__2527_ gnd vdd FILL
XFILL_4__2591_ gnd vdd FILL
XFILL_1__1833_ gnd vdd FILL
X_3318_ _3318_/D vdd _3347_/R _3573_/CLK _3318_/Q vdd gnd DFFSR
XFILL_6__2458_ gnd vdd FILL
XFILL_3__2749_ gnd vdd FILL
XFILL_1__1764_ gnd vdd FILL
XFILL_1__3503_ gnd vdd FILL
XFILL_1__1695_ gnd vdd FILL
XFILL_6__2389_ gnd vdd FILL
XFILL_4__3212_ gnd vdd FILL
X_3249_ _3249_/D vdd _3291_/R _3362_/CLK _3249_/Q vdd gnd DFFSR
XFILL_1__3434_ gnd vdd FILL
XFILL_4__3143_ gnd vdd FILL
XFILL_5_BUFX2_insert8 gnd vdd FILL
XFILL_4__3074_ gnd vdd FILL
XFILL_1__3365_ gnd vdd FILL
XFILL_4__2025_ gnd vdd FILL
XFILL_1__2316_ gnd vdd FILL
XFILL_1__2247_ gnd vdd FILL
XFILL_1__2178_ gnd vdd FILL
XFILL_7__2705_ gnd vdd FILL
XFILL_4__2927_ gnd vdd FILL
XFILL_2__2991_ gnd vdd FILL
XFILL_5__1720_ gnd vdd FILL
XFILL_2__1942_ gnd vdd FILL
XFILL_7__2636_ gnd vdd FILL
XFILL_4__2858_ gnd vdd FILL
XFILL_7__2567_ gnd vdd FILL
XFILL_2__1873_ gnd vdd FILL
XFILL_4__2789_ gnd vdd FILL
XFILL_4__1809_ gnd vdd FILL
XFILL_7__2498_ gnd vdd FILL
XFILL_8__3030_ gnd vdd FILL
XFILL_2__3543_ gnd vdd FILL
XFILL_2__3474_ gnd vdd FILL
XFILL_5__2203_ gnd vdd FILL
XFILL_7__3119_ gnd vdd FILL
XFILL_2__2425_ gnd vdd FILL
XFILL_5__3183_ gnd vdd FILL
XFILL_5__2134_ gnd vdd FILL
XFILL_5__2065_ gnd vdd FILL
XFILL_2__2356_ gnd vdd FILL
XFILL182850x101550 gnd vdd FILL
XFILL_2__2287_ gnd vdd FILL
XFILL_0__3110_ gnd vdd FILL
XFILL_8__2814_ gnd vdd FILL
XFILL_0__3041_ gnd vdd FILL
XFILL_8__2745_ gnd vdd FILL
XFILL_6__1760_ gnd vdd FILL
XFILL_5__2967_ gnd vdd FILL
X_2620_ _2767_/A _2630_/A _2621_/D vdd gnd NAND2X1
XFILL_5__1918_ gnd vdd FILL
XFILL_3__1982_ gnd vdd FILL
XFILL_8__2676_ gnd vdd FILL
XFILL_5__2898_ gnd vdd FILL
XFILL_6__1691_ gnd vdd FILL
X_2551_ _2551_/A _2552_/C vdd gnd INVX1
XFILL_6__3430_ gnd vdd FILL
X_2482_ _2482_/A _3573_/Q _2482_/C _2483_/C vdd gnd AOI21X1
XFILL_5__1849_ gnd vdd FILL
XFILL_5__3519_ gnd vdd FILL
XFILL_6__2312_ gnd vdd FILL
XFILL_3__3583_ gnd vdd FILL
XFILL_3__2603_ gnd vdd FILL
XFILL_0__2825_ gnd vdd FILL
XFILL_3__2534_ gnd vdd FILL
XFILL_8__3228_ gnd vdd FILL
X_3103_ _3125_/A _3107_/B _3328_/Q _3104_/C vdd gnd OAI21X1
XFILL_6__2243_ gnd vdd FILL
XFILL_0__2756_ gnd vdd FILL
XFILL_8__3159_ gnd vdd FILL
X_3034_ _3339_/Q _3278_/Q _3569_/Q _3056_/B vdd gnd NAND3X1
XFILL_0__1707_ gnd vdd FILL
XFILL_6__2174_ gnd vdd FILL
XFILL_3__2465_ gnd vdd FILL
XFILL_3__2396_ gnd vdd FILL
XFILL_0__2687_ gnd vdd FILL
XFILL_1__3150_ gnd vdd FILL
XFILL_1__3081_ gnd vdd FILL
XFILL_3__3017_ gnd vdd FILL
XFILL182550x74250 gnd vdd FILL
XFILL_1__2101_ gnd vdd FILL
XFILL_1__2032_ gnd vdd FILL
XFILL_6__1958_ gnd vdd FILL
X_2818_ _2933_/A _2931_/B _2920_/A vdd gnd NAND2X1
XFILL_7__3470_ gnd vdd FILL
XFILL_6__1889_ gnd vdd FILL
XFILL_4__2712_ gnd vdd FILL
X_2749_ _2749_/A _2749_/B _2750_/C vdd gnd OR2X2
XFILL_1__2934_ gnd vdd FILL
XFILL_7__2421_ gnd vdd FILL
XFILL_6__3559_ gnd vdd FILL
XFILL_7__2352_ gnd vdd FILL
XFILL_4__2643_ gnd vdd FILL
XFILL_1__2865_ gnd vdd FILL
XFILL_2_BUFX2_insert60 gnd vdd FILL
XFILL_4__2574_ gnd vdd FILL
XFILL_2_BUFX2_insert71 gnd vdd FILL
XFILL_2_BUFX2_insert93 gnd vdd FILL
XFILL_1__2796_ gnd vdd FILL
XFILL_2_BUFX2_insert82 gnd vdd FILL
XFILL_1__1816_ gnd vdd FILL
XFILL_7__2283_ gnd vdd FILL
XFILL_1__1747_ gnd vdd FILL
XFILL_4__3126_ gnd vdd FILL
XFILL_1__3417_ gnd vdd FILL
XFILL_2__2210_ gnd vdd FILL
XFILL_2__3190_ gnd vdd FILL
XFILL_2__2141_ gnd vdd FILL
XFILL_4__3057_ gnd vdd FILL
XFILL_2__2072_ gnd vdd FILL
XFILL_4__2008_ gnd vdd FILL
XFILL_7__1998_ gnd vdd FILL
XFILL_5__2821_ gnd vdd FILL
XFILL_8__2530_ gnd vdd FILL
XFILL_2_CLKBUF1_insert29 gnd vdd FILL
XFILL_8__2461_ gnd vdd FILL
XFILL_5__2752_ gnd vdd FILL
XFILL_2__2974_ gnd vdd FILL
XFILL_5__1703_ gnd vdd FILL
XFILL_5__2683_ gnd vdd FILL
XFILL_7__2619_ gnd vdd FILL
XFILL_7__3599_ gnd vdd FILL
XFILL_8__2392_ gnd vdd FILL
XFILL_2__1925_ gnd vdd FILL
XFILL_2__1856_ gnd vdd FILL
XFILL_2__3526_ gnd vdd FILL
XFILL_0_CLKBUF1_insert33 gnd vdd FILL
XFILL_8__3013_ gnd vdd FILL
XFILL_0__3590_ gnd vdd FILL
XFILL_0__2610_ gnd vdd FILL
XFILL_2__1787_ gnd vdd FILL
XFILL_0__2541_ gnd vdd FILL
XFILL_3__2250_ gnd vdd FILL
XFILL_2__3457_ gnd vdd FILL
XFILL_5__3166_ gnd vdd FILL
XFILL_2__3388_ gnd vdd FILL
XFILL_3__2181_ gnd vdd FILL
XFILL_5__2117_ gnd vdd FILL
XFILL_0__2472_ gnd vdd FILL
XFILL_2__2408_ gnd vdd FILL
XFILL_5__3097_ gnd vdd FILL
XFILL_2__2339_ gnd vdd FILL
XFILL_6__2930_ gnd vdd FILL
XFILL_5__2048_ gnd vdd FILL
XFILL_6__2861_ gnd vdd FILL
X_1982_ _3232_/A _2700_/B _2571_/A vdd gnd NOR2X1
XFILL_6__1812_ gnd vdd FILL
XFILL_6__2792_ gnd vdd FILL
XFILL_0__3024_ gnd vdd FILL
XFILL_8__2728_ gnd vdd FILL
XFILL_6__1743_ gnd vdd FILL
X_3583_ _3583_/A AB[12] vdd gnd BUFX2
X_2603_ _2781_/A _2958_/B _2746_/B _2604_/A vdd gnd OAI21X1
XFILL_8__2659_ gnd vdd FILL
XFILL_3__1965_ gnd vdd FILL
X_2534_ _3221_/A _2572_/B _2534_/C _2535_/C vdd gnd OAI21X1
XFILL_6__3413_ gnd vdd FILL
XFILL_3__1896_ gnd vdd FILL
X_2465_ _3291_/D _2502_/B _2502_/C _3349_/Q _2466_/B vdd gnd AOI22X1
X_2396_ _2627_/A _2426_/B _2396_/C _2397_/C vdd gnd OAI21X1
XFILL_1__2650_ gnd vdd FILL
XFILL_0__2808_ gnd vdd FILL
XFILL_3__3566_ gnd vdd FILL
XFILL_3__3497_ gnd vdd FILL
XFILL_6__2226_ gnd vdd FILL
XFILL_4__2290_ gnd vdd FILL
XFILL_3__2517_ gnd vdd FILL
XFILL_1__2581_ gnd vdd FILL
XFILL_0__2739_ gnd vdd FILL
XFILL_3__2448_ gnd vdd FILL
X_3017_ _3017_/A _3017_/B _3017_/C _3019_/B vdd gnd OAI21X1
XFILL_6__2157_ gnd vdd FILL
XFILL_7__2970_ gnd vdd FILL
XFILL_6__2088_ gnd vdd FILL
XFILL_3__2379_ gnd vdd FILL
XFILL_1__3202_ gnd vdd FILL
XFILL_1__3133_ gnd vdd FILL
XFILL_7__1921_ gnd vdd FILL
XFILL_1__3064_ gnd vdd FILL
XFILL_7__1852_ gnd vdd FILL
XFILL_1__2015_ gnd vdd FILL
XFILL_7__1783_ gnd vdd FILL
XFILL_7__3522_ gnd vdd FILL
XFILL_7__3453_ gnd vdd FILL
XFILL_7__2404_ gnd vdd FILL
XFILL_1__2917_ gnd vdd FILL
XFILL_7__3384_ gnd vdd FILL
XFILL_2__1710_ gnd vdd FILL
XFILL_2__2690_ gnd vdd FILL
XFILL_4__2626_ gnd vdd FILL
XFILL_1__2848_ gnd vdd FILL
XFILL_7__2335_ gnd vdd FILL
XFILL_7__2266_ gnd vdd FILL
XFILL_4__2557_ gnd vdd FILL
XFILL_7_BUFX2_insert17 gnd vdd FILL
XFILL_4__2488_ gnd vdd FILL
XFILL_1__2779_ gnd vdd FILL
XFILL_7__2197_ gnd vdd FILL
XFILL_7_BUFX2_insert39 gnd vdd FILL
XFILL_5__3020_ gnd vdd FILL
XFILL_8__1961_ gnd vdd FILL
XFILL_4__3109_ gnd vdd FILL
XFILL_2__3173_ gnd vdd FILL
XFILL_2__2124_ gnd vdd FILL
XFILL_8__1892_ gnd vdd FILL
XFILL_2__2055_ gnd vdd FILL
XFILL_8__3562_ gnd vdd FILL
XFILL_5__2804_ gnd vdd FILL
XFILL_8__2513_ gnd vdd FILL
XFILL_8__3493_ gnd vdd FILL
XFILL_5__2735_ gnd vdd FILL
XFILL_2__2957_ gnd vdd FILL
XFILL_3__1750_ gnd vdd FILL
XFILL_8__2444_ gnd vdd FILL
XFILL_0__1972_ gnd vdd FILL
XFILL_8__2375_ gnd vdd FILL
XFILL_5__2666_ gnd vdd FILL
XFILL_2__1908_ gnd vdd FILL
X_2250_ _2921_/A _2931_/A _2928_/B vdd gnd NAND2X1
XFILL_3__3420_ gnd vdd FILL
XFILL_2__2888_ gnd vdd FILL
XFILL_5__2597_ gnd vdd FILL
XFILL_2__1839_ gnd vdd FILL
X_2181_ _2824_/A _2268_/B _2853_/A vdd gnd NOR2X1
XFILL_6__3060_ gnd vdd FILL
XFILL_6__2011_ gnd vdd FILL
XFILL_2__3509_ gnd vdd FILL
XFILL184350x101550 gnd vdd FILL
XFILL_3__2302_ gnd vdd FILL
XFILL_5__3218_ gnd vdd FILL
XFILL_0__2524_ gnd vdd FILL
XFILL_3__2233_ gnd vdd FILL
XFILL_0__2455_ gnd vdd FILL
XFILL_5__3149_ gnd vdd FILL
XFILL_3__2164_ gnd vdd FILL
XFILL_0__2386_ gnd vdd FILL
XFILL_3__2095_ gnd vdd FILL
XFILL_6__2913_ gnd vdd FILL
X_1965_ _3329_/Q _3092_/A _1968_/A vdd gnd NAND2X1
XFILL_6__2844_ gnd vdd FILL
XFILL_0__3007_ gnd vdd FILL
X_1896_ _2872_/B _2288_/B _3185_/A vdd gnd NOR2X1
XFILL_6__2775_ gnd vdd FILL
XFILL_3__2997_ gnd vdd FILL
XFILL_6__1726_ gnd vdd FILL
XFILL_4__1790_ gnd vdd FILL
XFILL_3__1948_ gnd vdd FILL
X_3566_ _3566_/A _3566_/B _3566_/C _3578_/D vdd gnd OAI21X1
X_3497_ _3497_/A _3497_/B _3497_/C _3498_/C vdd gnd NAND3X1
X_2517_ _3247_/Q _2697_/B vdd gnd INVX1
XFILL_3__1879_ gnd vdd FILL
XFILL_4__3460_ gnd vdd FILL
XFILL_1__2702_ gnd vdd FILL
X_2448_ _3024_/A _2448_/B _2448_/C _2538_/B vdd gnd OAI21X1
XFILL_4__3391_ gnd vdd FILL
XFILL_7__2120_ gnd vdd FILL
XFILL_4__2411_ gnd vdd FILL
XFILL_3__3549_ gnd vdd FILL
XFILL_4__2342_ gnd vdd FILL
XFILL_1__2633_ gnd vdd FILL
X_2379_ _2379_/A _3149_/C _2409_/C vdd gnd NAND2X1
XFILL_7__2051_ gnd vdd FILL
XFILL_1__2564_ gnd vdd FILL
XFILL_4__2273_ gnd vdd FILL
XFILL_6__2209_ gnd vdd FILL
XFILL_6__3189_ gnd vdd FILL
XFILL_1__2495_ gnd vdd FILL
XFILL_7__2953_ gnd vdd FILL
XFILL_7__2884_ gnd vdd FILL
XFILL_1__3116_ gnd vdd FILL
XFILL_7__1904_ gnd vdd FILL
XFILL_1__3047_ gnd vdd FILL
XFILL_7__1835_ gnd vdd FILL
XFILL_7__1766_ gnd vdd FILL
XFILL184350x70350 gnd vdd FILL
XFILL_2__2811_ gnd vdd FILL
XFILL_7__3505_ gnd vdd FILL
XFILL_7__1697_ gnd vdd FILL
XFILL_4__1988_ gnd vdd FILL
XFILL_5__2520_ gnd vdd FILL
XFILL_7__3436_ gnd vdd FILL
XFILL_2__2742_ gnd vdd FILL
XFILL_8__2160_ gnd vdd FILL
XFILL_7__3367_ gnd vdd FILL
XFILL_5__2451_ gnd vdd FILL
XFILL_7__2318_ gnd vdd FILL
XFILL_5__2382_ gnd vdd FILL
XFILL_4__3589_ gnd vdd FILL
XFILL_4__2609_ gnd vdd FILL
XFILL_2__2673_ gnd vdd FILL
XFILL_8__2091_ gnd vdd FILL
XFILL_7__2249_ gnd vdd FILL
XFILL_5__3003_ gnd vdd FILL
XFILL_8__2993_ gnd vdd FILL
XFILL_2__3225_ gnd vdd FILL
XFILL_0__2240_ gnd vdd FILL
XFILL_2__3156_ gnd vdd FILL
XFILL_8__1944_ gnd vdd FILL
XFILL_8__1875_ gnd vdd FILL
XFILL_0__2171_ gnd vdd FILL
XFILL_2__2107_ gnd vdd FILL
XFILL_2__3087_ gnd vdd FILL
X_1750_ _1750_/A _1750_/B _1751_/C vdd gnd NOR2X1
XFILL_3__2920_ gnd vdd FILL
XFILL_2__2038_ gnd vdd FILL
XFILL_8__3545_ gnd vdd FILL
XFILL_3_BUFX2_insert26 gnd vdd FILL
XFILL_3__2851_ gnd vdd FILL
XFILL_3_BUFX2_insert15 gnd vdd FILL
XFILL_8__3476_ gnd vdd FILL
XFILL_3_BUFX2_insert59 gnd vdd FILL
XFILL_3_BUFX2_insert48 gnd vdd FILL
X_3420_ _3420_/A _3428_/B _3420_/C _3508_/B vdd gnd OAI21X1
XFILL_6__2560_ gnd vdd FILL
XFILL_3__1802_ gnd vdd FILL
XFILL_8__2427_ gnd vdd FILL
XFILL_6__2491_ gnd vdd FILL
XFILL_5__2718_ gnd vdd FILL
XFILL_3__2782_ gnd vdd FILL
X_3351_ _3351_/D vdd _3362_/R _3355_/CLK _3351_/Q vdd gnd DFFSR
XFILL184350x113250 gnd vdd FILL
XFILL184650x105450 gnd vdd FILL
X_2302_ _2345_/A _2327_/B _2302_/C _2303_/B vdd gnd NAND3X1
XFILL_3__1733_ gnd vdd FILL
XFILL_5__2649_ gnd vdd FILL
XFILL184050x121050 gnd vdd FILL
X_3282_ _3282_/D vdd _3282_/R _3284_/CLK _3282_/Q vdd gnd DFFSR
XFILL_8__2358_ gnd vdd FILL
XFILL_0__1955_ gnd vdd FILL
XFILL_6__3112_ gnd vdd FILL
XFILL_3__3403_ gnd vdd FILL
XFILL_0__1886_ gnd vdd FILL
X_2233_ _3148_/B _2233_/B _2234_/C vdd gnd NOR2X1
XFILL_8__2289_ gnd vdd FILL
X_2164_ _2823_/B _2823_/C _2792_/C vdd gnd NAND2X1
XFILL_6__3043_ gnd vdd FILL
XFILL_0__3556_ gnd vdd FILL
XFILL_0__2507_ gnd vdd FILL
X_2095_ _2294_/A _2872_/B _2096_/C vdd gnd NAND2X1
XFILL_0__3487_ gnd vdd FILL
XFILL_3__2216_ gnd vdd FILL
XFILL_1__2280_ gnd vdd FILL
XFILL_3__3196_ gnd vdd FILL
XFILL_3__2147_ gnd vdd FILL
XFILL_0__2438_ gnd vdd FILL
XFILL_0__2369_ gnd vdd FILL
XFILL_3__2078_ gnd vdd FILL
XFILL_4__2960_ gnd vdd FILL
X_2997_ _3311_/Q _2998_/A _2998_/C vdd gnd NAND2X1
XFILL_4__2891_ gnd vdd FILL
X_1948_ _3335_/Q _3110_/A _3127_/B _3344_/Q _1950_/C vdd gnd AOI22X1
XFILL_4__1911_ gnd vdd FILL
XFILL_9__2605_ gnd vdd FILL
X_1879_ _1879_/A _1879_/B _1879_/C _3110_/A vdd gnd AOI21X1
XFILL_6__2827_ gnd vdd FILL
XFILL_4__1842_ gnd vdd FILL
XFILL_6__2758_ gnd vdd FILL
XFILL_6__1709_ gnd vdd FILL
XFILL_6__2689_ gnd vdd FILL
XFILL_4__1773_ gnd vdd FILL
X_3549_ _3572_/Q _3550_/A _3550_/C vdd gnd NAND2X1
XFILL_4__3512_ gnd vdd FILL
XFILL_7__3221_ gnd vdd FILL
XFILL_1__1995_ gnd vdd FILL
XFILL_4__3443_ gnd vdd FILL
XFILL_7__3152_ gnd vdd FILL
XFILL_4__3374_ gnd vdd FILL
XFILL_7__3083_ gnd vdd FILL
XFILL_1__2616_ gnd vdd FILL
XFILL_7__2103_ gnd vdd FILL
XFILL_7__2034_ gnd vdd FILL
XFILL_4__2325_ gnd vdd FILL
XFILL_1__3596_ gnd vdd FILL
XFILL_4__2256_ gnd vdd FILL
XFILL_1__2547_ gnd vdd FILL
XFILL_1__2478_ gnd vdd FILL
XFILL_2__3010_ gnd vdd FILL
XFILL_4__2187_ gnd vdd FILL
XFILL_7__2936_ gnd vdd FILL
XFILL_7_CLKBUF1_insert29 gnd vdd FILL
XFILL_5__1951_ gnd vdd FILL
XFILL184350x82050 gnd vdd FILL
XFILL_7__2867_ gnd vdd FILL
XFILL_7__2798_ gnd vdd FILL
XFILL_5__1882_ gnd vdd FILL
XFILL_7__1818_ gnd vdd FILL
XFILL_7__1749_ gnd vdd FILL
XFILL_5__3552_ gnd vdd FILL
XFILL_5_CLKBUF1_insert33 gnd vdd FILL
XFILL_5__3483_ gnd vdd FILL
XFILL_5__2503_ gnd vdd FILL
XFILL_8__2212_ gnd vdd FILL
XFILL_7__3419_ gnd vdd FILL
XFILL_2__2725_ gnd vdd FILL
XFILL_8__3192_ gnd vdd FILL
XFILL_5__2434_ gnd vdd FILL
XFILL_8__2143_ gnd vdd FILL
XFILL_0__1740_ gnd vdd FILL
XFILL_2__2656_ gnd vdd FILL
XFILL_8__2074_ gnd vdd FILL
XFILL_5__2365_ gnd vdd FILL
XFILL_0__3410_ gnd vdd FILL
XFILL_5__2296_ gnd vdd FILL
XFILL_2__2587_ gnd vdd FILL
XFILL_3__3050_ gnd vdd FILL
X_2920_ _2920_/A _2932_/C vdd gnd INVX1
XFILL_3__2001_ gnd vdd FILL
XFILL_2__3208_ gnd vdd FILL
XFILL_8__2976_ gnd vdd FILL
XFILL_6__1991_ gnd vdd FILL
XFILL_0__2223_ gnd vdd FILL
X_2851_ _2851_/A _2880_/A vdd gnd INVX1
XFILL_2__3139_ gnd vdd FILL
XFILL_8__1927_ gnd vdd FILL
XFILL_0__2154_ gnd vdd FILL
XFILL_8__1858_ gnd vdd FILL
X_2782_ _3256_/Q _2782_/B _2782_/C _3256_/D vdd gnd OAI21X1
X_1802_ _2058_/B _2602_/B _1885_/A vdd gnd NAND2X1
XFILL_3__2903_ gnd vdd FILL
XFILL_0__2085_ gnd vdd FILL
XFILL184650x117150 gnd vdd FILL
X_1733_ _3237_/Q _3166_/C _1733_/Y vdd gnd NOR2X1
XFILL_8__3528_ gnd vdd FILL
XFILL_6__3592_ gnd vdd FILL
XFILL_6__2612_ gnd vdd FILL
XFILL_8__1789_ gnd vdd FILL
XFILL_3__2834_ gnd vdd FILL
X_3403_ _3403_/A _3428_/B _3403_/C _3518_/B vdd gnd OAI21X1
XFILL_6__2543_ gnd vdd FILL
XFILL_8__3459_ gnd vdd FILL
XFILL_9__2252_ gnd vdd FILL
XFILL_3__2765_ gnd vdd FILL
X_3334_ _3334_/D vdd _3347_/R _3573_/CLK _3334_/Q vdd gnd DFFSR
XFILL_0__2987_ gnd vdd FILL
XFILL_1__1780_ gnd vdd FILL
XFILL_6__2474_ gnd vdd FILL
XFILL_3__1716_ gnd vdd FILL
XFILL_0__1938_ gnd vdd FILL
X_3265_ _3265_/D vdd _3282_/R _3284_/CLK _3265_/Q vdd gnd DFFSR
XFILL_3__2696_ gnd vdd FILL
XFILL_1__3450_ gnd vdd FILL
X_2216_ _2922_/A _2843_/C _2268_/B _2247_/B vdd gnd OAI21X1
XFILL_0__1869_ gnd vdd FILL
XFILL_1__2401_ gnd vdd FILL
X_3196_ _3196_/A _3196_/B _3196_/C _3196_/D _3197_/B vdd gnd AOI22X1
XFILL_4__3090_ gnd vdd FILL
XFILL_1__3381_ gnd vdd FILL
XFILL_6__3026_ gnd vdd FILL
X_2147_ _2341_/A _3077_/C _2147_/C _2330_/A vdd gnd OAI21X1
XFILL_4__2110_ gnd vdd FILL
X_2078_ _2824_/A _2915_/C vdd gnd INVX1
XFILL_4__2041_ gnd vdd FILL
XFILL_0__3539_ gnd vdd FILL
XFILL_1__2332_ gnd vdd FILL
XFILL_1__2263_ gnd vdd FILL
XFILL_3__3179_ gnd vdd FILL
XFILL_1__2194_ gnd vdd FILL
XFILL_4__2943_ gnd vdd FILL
XFILL_7__2721_ gnd vdd FILL
XFILL_7__2652_ gnd vdd FILL
XFILL_4__2874_ gnd vdd FILL
XFILL_7__2583_ gnd vdd FILL
XFILL_4__1825_ gnd vdd FILL
XFILL_4__1756_ gnd vdd FILL
XFILL_1__1978_ gnd vdd FILL
XFILL_7__3204_ gnd vdd FILL
XFILL_2__2510_ gnd vdd FILL
XFILL_7__3135_ gnd vdd FILL
XFILL_2__3490_ gnd vdd FILL
XFILL_4__3426_ gnd vdd FILL
XFILL_5__2150_ gnd vdd FILL
XFILL_2__2441_ gnd vdd FILL
XFILL_2__2372_ gnd vdd FILL
XFILL_7__3066_ gnd vdd FILL
XFILL_4__2308_ gnd vdd FILL
XFILL_1__3579_ gnd vdd FILL
XFILL_7__2017_ gnd vdd FILL
XFILL_5__2081_ gnd vdd FILL
XFILL_8__2830_ gnd vdd FILL
XFILL_4__2239_ gnd vdd FILL
XFILL_8__2761_ gnd vdd FILL
XFILL_7__2919_ gnd vdd FILL
XFILL_5__2983_ gnd vdd FILL
XFILL_8__1712_ gnd vdd FILL
XFILL_8__2692_ gnd vdd FILL
XFILL_5__1934_ gnd vdd FILL
XFILL_5__1865_ gnd vdd FILL
XFILL_0__2910_ gnd vdd FILL
XFILL_2_BUFX2_insert5 gnd vdd FILL
XFILL_5__1796_ gnd vdd FILL
XFILL_0__2841_ gnd vdd FILL
XFILL_5__3535_ gnd vdd FILL
XFILL_3__2550_ gnd vdd FILL
XFILL_5__3466_ gnd vdd FILL
XFILL_2__2708_ gnd vdd FILL
XFILL_8__3175_ gnd vdd FILL
XFILL_0__2772_ gnd vdd FILL
XFILL_5__3397_ gnd vdd FILL
X_3050_ _3050_/A _3050_/B _3055_/A vdd gnd NOR2X1
XFILL_6__2190_ gnd vdd FILL
XFILL_5__2417_ gnd vdd FILL
XFILL_8__2126_ gnd vdd FILL
XFILL_3__2481_ gnd vdd FILL
XFILL_0__1723_ gnd vdd FILL
X_2001_ _2001_/A _2025_/A _2702_/B _2002_/C vdd gnd AOI21X1
XFILL_5__2348_ gnd vdd FILL
XFILL_2__2639_ gnd vdd FILL
XFILL_8__2057_ gnd vdd FILL
XFILL_3__3102_ gnd vdd FILL
XFILL_5__2279_ gnd vdd FILL
XFILL_9__2870_ gnd vdd FILL
XFILL_6_BUFX2_insert63 gnd vdd FILL
XFILL_6_BUFX2_insert52 gnd vdd FILL
XFILL_6_BUFX2_insert41 gnd vdd FILL
XFILL_6_BUFX2_insert96 gnd vdd FILL
XFILL_3__3033_ gnd vdd FILL
XFILL_6_BUFX2_insert85 gnd vdd FILL
XFILL_6_BUFX2_insert74 gnd vdd FILL
X_2903_ _2915_/C _2903_/B _2903_/C _2913_/C vdd gnd AOI21X1
XFILL_8__2959_ gnd vdd FILL
X_2834_ _2870_/B _2865_/D vdd gnd INVX1
XFILL_0__2206_ gnd vdd FILL
XFILL_6__1974_ gnd vdd FILL
XFILL_0__3186_ gnd vdd FILL
XFILL_0__2137_ gnd vdd FILL
X_2765_ _2775_/A _2775_/C _2766_/C vdd gnd NAND2X1
XFILL_1__2950_ gnd vdd FILL
XFILL_0__2068_ gnd vdd FILL
X_2696_ _2696_/A _2696_/B _2767_/A _2697_/C vdd gnd OAI21X1
X_1716_ _3238_/Q _3237_/Q _1716_/Y vdd gnd NOR2X1
XFILL_3__2817_ gnd vdd FILL
XFILL_1__2881_ gnd vdd FILL
XFILL_1__1901_ gnd vdd FILL
XFILL_1__1832_ gnd vdd FILL
XFILL_4__2590_ gnd vdd FILL
XFILL_6__2526_ gnd vdd FILL
X_3317_ _3317_/D vdd _3345_/R _3576_/CLK _3317_/Q vdd gnd DFFSR
XFILL_6__2457_ gnd vdd FILL
XFILL_3__2748_ gnd vdd FILL
XFILL_1__3502_ gnd vdd FILL
XFILL_1__1763_ gnd vdd FILL
XFILL_3__2679_ gnd vdd FILL
XFILL_6__2388_ gnd vdd FILL
XFILL_1__1694_ gnd vdd FILL
XFILL_4__3211_ gnd vdd FILL
X_3248_ _3248_/D vdd _3291_/R _3362_/CLK _3248_/Q vdd gnd DFFSR
XFILL_4__3142_ gnd vdd FILL
XFILL_1__3433_ gnd vdd FILL
X_3179_ _3179_/A _3179_/B _3179_/C _3186_/C vdd gnd NAND3X1
XFILL_1__3364_ gnd vdd FILL
XFILL_5_BUFX2_insert9 gnd vdd FILL
XFILL_6__3009_ gnd vdd FILL
XFILL_1__2315_ gnd vdd FILL
XFILL_4__3073_ gnd vdd FILL
XFILL_4__2024_ gnd vdd FILL
XFILL_1__2246_ gnd vdd FILL
XFILL_1__2177_ gnd vdd FILL
XFILL_7__2704_ gnd vdd FILL
XFILL_4__2926_ gnd vdd FILL
XFILL_2__2990_ gnd vdd FILL
XFILL_2__1941_ gnd vdd FILL
XFILL_7__2635_ gnd vdd FILL
XFILL_2__1872_ gnd vdd FILL
XFILL_4__2857_ gnd vdd FILL
XFILL_7__2566_ gnd vdd FILL
XFILL_4__2788_ gnd vdd FILL
XFILL_7__2497_ gnd vdd FILL
XFILL_4__1808_ gnd vdd FILL
XFILL_4__1739_ gnd vdd FILL
XFILL_2__3542_ gnd vdd FILL
XFILL_2__3473_ gnd vdd FILL
XFILL_4__3409_ gnd vdd FILL
XFILL_5__2202_ gnd vdd FILL
XFILL_7__3118_ gnd vdd FILL
XFILL_2__2424_ gnd vdd FILL
XFILL_5__3182_ gnd vdd FILL
XFILL_7__3049_ gnd vdd FILL
XFILL_5__2133_ gnd vdd FILL
XFILL_5__2064_ gnd vdd FILL
XFILL_2__2355_ gnd vdd FILL
XFILL_2__2286_ gnd vdd FILL
XFILL_8__2813_ gnd vdd FILL
XFILL_0__3040_ gnd vdd FILL
XFILL_8__2744_ gnd vdd FILL
XFILL_5__2966_ gnd vdd FILL
XFILL_5__1917_ gnd vdd FILL
XFILL_3__1981_ gnd vdd FILL
XFILL_8__2675_ gnd vdd FILL
XFILL_5__2897_ gnd vdd FILL
XFILL_6__1690_ gnd vdd FILL
X_2550_ _3226_/A _2572_/B _2550_/C _2551_/A vdd gnd OAI21X1
X_2481_ _2948_/A _2510_/B _2632_/A _2510_/D _2482_/C vdd gnd OAI22X1
XFILL_5__1848_ gnd vdd FILL
XFILL_3__2602_ gnd vdd FILL
XFILL_5__1779_ gnd vdd FILL
XFILL_0__2824_ gnd vdd FILL
XFILL_5__3518_ gnd vdd FILL
XFILL_6__2311_ gnd vdd FILL
XFILL_3__3582_ gnd vdd FILL
XFILL_6__2242_ gnd vdd FILL
XFILL_3__2533_ gnd vdd FILL
XFILL_8__3227_ gnd vdd FILL
X_3102_ _3137_/A _3108_/B _3102_/C _3327_/D vdd gnd OAI21X1
XFILL_5__3449_ gnd vdd FILL
XFILL_3__2464_ gnd vdd FILL
XFILL_0__2755_ gnd vdd FILL
XFILL_8__3158_ gnd vdd FILL
X_3033_ _3090_/A _3129_/A _3033_/C _3315_/D vdd gnd OAI21X1
XFILL_6__2173_ gnd vdd FILL
XFILL_0__1706_ gnd vdd FILL
XFILL_0__2686_ gnd vdd FILL
XFILL_8__2109_ gnd vdd FILL
XFILL_8__3089_ gnd vdd FILL
XFILL_3__2395_ gnd vdd FILL
XFILL_1__3080_ gnd vdd FILL
XFILL_3__3016_ gnd vdd FILL
XFILL_1__2100_ gnd vdd FILL
XFILL_1__2031_ gnd vdd FILL
XFILL_6__1957_ gnd vdd FILL
X_2817_ _2933_/B _2857_/A _2931_/B vdd gnd NOR2X1
XFILL_0__3169_ gnd vdd FILL
XFILL_6__1888_ gnd vdd FILL
XFILL_4__2711_ gnd vdd FILL
X_2748_ _3228_/A _2748_/B _2748_/C _2749_/A vdd gnd OAI21X1
XFILL_1__2933_ gnd vdd FILL
XFILL_7__2420_ gnd vdd FILL
XFILL_6__3558_ gnd vdd FILL
XFILL_7__2351_ gnd vdd FILL
XFILL_4__2642_ gnd vdd FILL
X_2679_ _3570_/Q _2701_/B _3166_/D _2681_/B vdd gnd NAND3X1
XFILL_2_BUFX2_insert61 gnd vdd FILL
XFILL_2_BUFX2_insert50 gnd vdd FILL
XFILL_1__2864_ gnd vdd FILL
XFILL_6__2509_ gnd vdd FILL
XFILL_4__2573_ gnd vdd FILL
XFILL_2_BUFX2_insert72 gnd vdd FILL
XFILL_6__3489_ gnd vdd FILL
XFILL_2_BUFX2_insert94 gnd vdd FILL
XFILL_1__2795_ gnd vdd FILL
XFILL_2_BUFX2_insert83 gnd vdd FILL
XFILL_7__2282_ gnd vdd FILL
XFILL_1__1815_ gnd vdd FILL
XFILL_9__2149_ gnd vdd FILL
XFILL_1__1746_ gnd vdd FILL
XFILL_1__3416_ gnd vdd FILL
XFILL_4__3125_ gnd vdd FILL
XFILL_4__3056_ gnd vdd FILL
XFILL_2__2140_ gnd vdd FILL
XFILL_2__2071_ gnd vdd FILL
XFILL_4__2007_ gnd vdd FILL
XFILL_1__2229_ gnd vdd FILL
XFILL_5__2820_ gnd vdd FILL
XFILL_7__1997_ gnd vdd FILL
XFILL_2__2973_ gnd vdd FILL
XFILL_8__2460_ gnd vdd FILL
XFILL_5__2751_ gnd vdd FILL
XFILL_4__2909_ gnd vdd FILL
XFILL_8__2391_ gnd vdd FILL
XFILL_5__1702_ gnd vdd FILL
XFILL_5__2682_ gnd vdd FILL
XFILL_7__2618_ gnd vdd FILL
XFILL_2__1924_ gnd vdd FILL
XFILL_7__3598_ gnd vdd FILL
XFILL_2__1855_ gnd vdd FILL
XFILL_7__2549_ gnd vdd FILL
XFILL_2__1786_ gnd vdd FILL
XFILL_0_CLKBUF1_insert34 gnd vdd FILL
XFILL_2__3525_ gnd vdd FILL
XFILL_8__3012_ gnd vdd FILL
XFILL_0__2540_ gnd vdd FILL
XFILL_2__3456_ gnd vdd FILL
XFILL_5__3165_ gnd vdd FILL
XFILL_3__2180_ gnd vdd FILL
XFILL_2__3387_ gnd vdd FILL
XFILL_5__2116_ gnd vdd FILL
XFILL_0__2471_ gnd vdd FILL
XFILL_2__2407_ gnd vdd FILL
XFILL_5__3096_ gnd vdd FILL
XFILL_2__2338_ gnd vdd FILL
XFILL182250x148350 gnd vdd FILL
XFILL_5__2047_ gnd vdd FILL
XFILL_6__2860_ gnd vdd FILL
XFILL_2__2269_ gnd vdd FILL
X_1981_ _3363_/Q _3232_/A vdd gnd INVX1
XFILL_0__3023_ gnd vdd FILL
XFILL_6__1811_ gnd vdd FILL
XFILL_6__2791_ gnd vdd FILL
XFILL_8__2727_ gnd vdd FILL
XFILL_5__2949_ gnd vdd FILL
XFILL_6__1742_ gnd vdd FILL
X_2602_ _2602_/A _2602_/B _2889_/C _2746_/B vdd gnd NAND3X1
X_3582_ _3582_/A AB[11] vdd gnd BUFX2
XFILL_8__2658_ gnd vdd FILL
XFILL_3__1964_ gnd vdd FILL
X_2533_ _3358_/Q _2691_/A _2563_/A _3572_/Q _2534_/C vdd gnd AOI22X1
XFILL_6__3412_ gnd vdd FILL
XFILL_8__2589_ gnd vdd FILL
XFILL_3__1895_ gnd vdd FILL
X_2464_ _2508_/B _2511_/A _3571_/Q _2466_/A vdd gnd OAI21X1
XFILL_3__3565_ gnd vdd FILL
X_2395_ _3310_/Q _2425_/B _2396_/C vdd gnd NAND2X1
XFILL_1__2580_ gnd vdd FILL
XFILL_0__2807_ gnd vdd FILL
XFILL_3__3496_ gnd vdd FILL
XFILL_3__2516_ gnd vdd FILL
XFILL_6__2225_ gnd vdd FILL
XFILL_0__2738_ gnd vdd FILL
XFILL_6__2156_ gnd vdd FILL
XFILL_3__2447_ gnd vdd FILL
X_3016_ _3016_/A _3017_/A _3017_/C vdd gnd NAND2X1
XFILL_3__2378_ gnd vdd FILL
XFILL_0__2669_ gnd vdd FILL
XFILL_6__2087_ gnd vdd FILL
XFILL_1__3201_ gnd vdd FILL
XFILL_1__3132_ gnd vdd FILL
XFILL_7__1920_ gnd vdd FILL
XFILL_7__1851_ gnd vdd FILL
XFILL_9__2767_ gnd vdd FILL
XFILL_1__3063_ gnd vdd FILL
XFILL_6__2989_ gnd vdd FILL
XFILL_1__2014_ gnd vdd FILL
XFILL_7__1782_ gnd vdd FILL
XFILL_7__3521_ gnd vdd FILL
XFILL_7__3452_ gnd vdd FILL
XFILL_7__2403_ gnd vdd FILL
XFILL_1__2916_ gnd vdd FILL
XFILL_7__3383_ gnd vdd FILL
XFILL_4__2625_ gnd vdd FILL
XFILL_1__2847_ gnd vdd FILL
XFILL_7__2334_ gnd vdd FILL
XFILL_7__2265_ gnd vdd FILL
XFILL_4__2556_ gnd vdd FILL
XFILL_7_BUFX2_insert18 gnd vdd FILL
XFILL_4__2487_ gnd vdd FILL
XFILL_1__2778_ gnd vdd FILL
XFILL_7__2196_ gnd vdd FILL
XFILL_1__1729_ gnd vdd FILL
XFILL_8__1960_ gnd vdd FILL
XFILL_2__3172_ gnd vdd FILL
XFILL_4__3108_ gnd vdd FILL
XFILL_2__2123_ gnd vdd FILL
XFILL_4__3039_ gnd vdd FILL
XFILL_8__1891_ gnd vdd FILL
XFILL_2__2054_ gnd vdd FILL
XFILL_8__3561_ gnd vdd FILL
XFILL_5__2803_ gnd vdd FILL
XFILL_8__2512_ gnd vdd FILL
XFILL_8__3492_ gnd vdd FILL
XFILL_5__2734_ gnd vdd FILL
XFILL_2__2956_ gnd vdd FILL
XFILL_7_BUFX2_insert0 gnd vdd FILL
XFILL_8__2443_ gnd vdd FILL
XFILL_2__2887_ gnd vdd FILL
XFILL_8__2374_ gnd vdd FILL
XFILL_2__1907_ gnd vdd FILL
XFILL_0__1971_ gnd vdd FILL
XFILL_5__2665_ gnd vdd FILL
XFILL_5__2596_ gnd vdd FILL
X_2180_ _2864_/A _2915_/A _2268_/B vdd gnd NAND2X1
XFILL_2__1838_ gnd vdd FILL
XFILL_2__1769_ gnd vdd FILL
XFILL_6__2010_ gnd vdd FILL
XFILL_2__3508_ gnd vdd FILL
XFILL_3__2301_ gnd vdd FILL
XFILL_5__3217_ gnd vdd FILL
XFILL_2__3439_ gnd vdd FILL
XFILL_3__2232_ gnd vdd FILL
XFILL_0__2523_ gnd vdd FILL
XFILL_0__2454_ gnd vdd FILL
XFILL_5__3148_ gnd vdd FILL
XFILL_3__2163_ gnd vdd FILL
XFILL_5__3079_ gnd vdd FILL
XFILL_6__2912_ gnd vdd FILL
XFILL_0__2385_ gnd vdd FILL
XFILL_3__2094_ gnd vdd FILL
X_1964_ _1986_/A _2416_/B _1964_/C _3413_/B vdd gnd OAI21X1
XFILL_6__2843_ gnd vdd FILL
XFILL_0__3006_ gnd vdd FILL
XFILL_6__2774_ gnd vdd FILL
X_1895_ _1895_/A _2288_/B vdd gnd INVX1
XFILL_3__2996_ gnd vdd FILL
XFILL_6__1725_ gnd vdd FILL
XFILL_3__1947_ gnd vdd FILL
X_3565_ _3565_/A _3566_/A _3566_/C vdd gnd NAND2X1
X_3496_ _3526_/B _3526_/A _3498_/A vdd gnd NAND2X1
X_2516_ _3215_/B _3592_/A vdd gnd INVX1
XFILL_3__1878_ gnd vdd FILL
X_2447_ _2508_/B _2511_/A _2457_/A vdd gnd NOR2X1
XFILL_1__2701_ gnd vdd FILL
XFILL_4__3390_ gnd vdd FILL
XFILL_1__2632_ gnd vdd FILL
XFILL_4__2410_ gnd vdd FILL
XFILL_3__3548_ gnd vdd FILL
XFILL_4__2341_ gnd vdd FILL
X_2378_ _2872_/B _3077_/C _3247_/Q _2386_/A vdd gnd OAI21X1
XFILL_7__2050_ gnd vdd FILL
XFILL_4__2272_ gnd vdd FILL
XFILL_1__2563_ gnd vdd FILL
XFILL_3__3479_ gnd vdd FILL
XFILL_6__2208_ gnd vdd FILL
XFILL_1__2494_ gnd vdd FILL
XFILL_6__3188_ gnd vdd FILL
XFILL_6__2139_ gnd vdd FILL
XFILL_7__2952_ gnd vdd FILL
XFILL_7__2883_ gnd vdd FILL
XFILL_1__3115_ gnd vdd FILL
XFILL_7__1903_ gnd vdd FILL
XFILL_1__3046_ gnd vdd FILL
XFILL_7__1834_ gnd vdd FILL
XFILL184650x54750 gnd vdd FILL
XFILL_7__3504_ gnd vdd FILL
XFILL_7__1765_ gnd vdd FILL
XFILL_2__2810_ gnd vdd FILL
XFILL_7__1696_ gnd vdd FILL
XFILL_4__1987_ gnd vdd FILL
XFILL_7__3435_ gnd vdd FILL
XFILL_2__2741_ gnd vdd FILL
XFILL_7__3366_ gnd vdd FILL
XFILL_5__2450_ gnd vdd FILL
XFILL_7__2317_ gnd vdd FILL
XFILL_5__2381_ gnd vdd FILL
XFILL_4__3588_ gnd vdd FILL
XFILL_2__2672_ gnd vdd FILL
XFILL_4__2608_ gnd vdd FILL
XFILL_8__2090_ gnd vdd FILL
XFILL_4__2539_ gnd vdd FILL
XFILL_7__2248_ gnd vdd FILL
XFILL_7__2179_ gnd vdd FILL
XFILL_5__3002_ gnd vdd FILL
XFILL_2__3224_ gnd vdd FILL
XFILL_8__2992_ gnd vdd FILL
XFILL_2__3155_ gnd vdd FILL
XFILL_8__1943_ gnd vdd FILL
XFILL_8__1874_ gnd vdd FILL
XFILL_0__2170_ gnd vdd FILL
XFILL_2__3086_ gnd vdd FILL
XFILL_2__2106_ gnd vdd FILL
XFILL_2__2037_ gnd vdd FILL
XFILL_3__2850_ gnd vdd FILL
XFILL_8__3544_ gnd vdd FILL
XFILL_3_BUFX2_insert27 gnd vdd FILL
XFILL_3_BUFX2_insert16 gnd vdd FILL
XFILL_8__3475_ gnd vdd FILL
XFILL_3_BUFX2_insert49 gnd vdd FILL
XFILL_3__2781_ gnd vdd FILL
XFILL_3__1801_ gnd vdd FILL
XFILL_8__2426_ gnd vdd FILL
X_3350_ _3350_/D vdd _3355_/R _3578_/CLK _3350_/Q vdd gnd DFFSR
XFILL_6__2490_ gnd vdd FILL
XFILL_5__2717_ gnd vdd FILL
XFILL_2__2939_ gnd vdd FILL
X_2301_ _2314_/A _2305_/A _2302_/C vdd gnd OR2X2
XFILL_0__1954_ gnd vdd FILL
XFILL_3__1732_ gnd vdd FILL
XFILL_5__2648_ gnd vdd FILL
X_3281_ _3281_/D vdd _3289_/R _3307_/CLK _3281_/Q vdd gnd DFFSR
XFILL_8__2357_ gnd vdd FILL
XFILL_6__3111_ gnd vdd FILL
XFILL_5__2579_ gnd vdd FILL
XFILL_3__3402_ gnd vdd FILL
XFILL_8__2288_ gnd vdd FILL
XFILL_0__1885_ gnd vdd FILL
X_2232_ _3173_/B _2781_/A _2586_/B _2233_/B vdd gnd OAI21X1
X_2163_ _2910_/B _2857_/A _2823_/C vdd gnd NOR2X1
XFILL_0__3555_ gnd vdd FILL
XFILL_6__3042_ gnd vdd FILL
XFILL_0__2506_ gnd vdd FILL
X_2094_ _2293_/A _3183_/C _2094_/C _2349_/A vdd gnd OAI21X1
XFILL_0__3486_ gnd vdd FILL
XFILL_3__2215_ gnd vdd FILL
XFILL_3__3195_ gnd vdd FILL
XFILL_3__2146_ gnd vdd FILL
XFILL_0__2437_ gnd vdd FILL
XFILL_0__2368_ gnd vdd FILL
X_2996_ _3011_/B _2996_/B _2996_/C _2998_/B vdd gnd OAI21X1
XFILL_3__2077_ gnd vdd FILL
XFILL_4__2890_ gnd vdd FILL
X_1947_ _3327_/Q _3092_/A _1950_/A vdd gnd NAND2X1
XFILL_6__2826_ gnd vdd FILL
XFILL_0__2299_ gnd vdd FILL
XFILL_4__1910_ gnd vdd FILL
X_1878_ _1878_/A _1878_/B _3092_/A vdd gnd NOR2X1
XFILL_4__1841_ gnd vdd FILL
XFILL_6__2757_ gnd vdd FILL
X_3548_ _3550_/A _3548_/B _3548_/C _3571_/D vdd gnd OAI21X1
XFILL_3__2979_ gnd vdd FILL
XFILL_4__1772_ gnd vdd FILL
XFILL_6__1708_ gnd vdd FILL
XFILL_6__2688_ gnd vdd FILL
XFILL_4__3511_ gnd vdd FILL
XFILL_1__1994_ gnd vdd FILL
XFILL_7__3220_ gnd vdd FILL
X_3479_ _3479_/A _3480_/B vdd gnd INVX1
XFILL_4__3442_ gnd vdd FILL
XFILL_7__3151_ gnd vdd FILL
XFILL_7__3082_ gnd vdd FILL
XFILL_4__3373_ gnd vdd FILL
XFILL_1__3595_ gnd vdd FILL
XFILL_7__2102_ gnd vdd FILL
XFILL_1__2615_ gnd vdd FILL
XFILL_7__2033_ gnd vdd FILL
XFILL_4__2324_ gnd vdd FILL
XFILL_1__2546_ gnd vdd FILL
XFILL_4__2255_ gnd vdd FILL
XFILL_4__2186_ gnd vdd FILL
XFILL_1__2477_ gnd vdd FILL
XFILL_7__2935_ gnd vdd FILL
XFILL181650x74250 gnd vdd FILL
XFILL_5__1950_ gnd vdd FILL
XFILL_7__2866_ gnd vdd FILL
XFILL_1__3029_ gnd vdd FILL
XFILL_5__1881_ gnd vdd FILL
XFILL_7__2797_ gnd vdd FILL
XFILL_7__1817_ gnd vdd FILL
XFILL_7__1748_ gnd vdd FILL
XFILL_5__3551_ gnd vdd FILL
XFILL_5_CLKBUF1_insert34 gnd vdd FILL
XFILL_5__3482_ gnd vdd FILL
XFILL_7__3418_ gnd vdd FILL
XFILL_8__2211_ gnd vdd FILL
XFILL_5__2502_ gnd vdd FILL
XFILL_2__2724_ gnd vdd FILL
XFILL_8__3191_ gnd vdd FILL
XFILL_5__2433_ gnd vdd FILL
XFILL_8__2142_ gnd vdd FILL
XFILL_2__2655_ gnd vdd FILL
XFILL_8__2073_ gnd vdd FILL
XFILL_5__2364_ gnd vdd FILL
XFILL_5__2295_ gnd vdd FILL
XFILL_2__2586_ gnd vdd FILL
XFILL_3__2000_ gnd vdd FILL
XFILL_8__2975_ gnd vdd FILL
XFILL_2__3207_ gnd vdd FILL
X_2850_ _2850_/A _2916_/C vdd gnd INVX1
XFILL_2__3138_ gnd vdd FILL
XFILL_8__1926_ gnd vdd FILL
XFILL_6__1990_ gnd vdd FILL
XFILL_0__2222_ gnd vdd FILL
XFILL_0__2153_ gnd vdd FILL
X_1801_ _1858_/B _1891_/A _2602_/B vdd gnd AND2X2
XFILL_8__1857_ gnd vdd FILL
XFILL_2__3069_ gnd vdd FILL
X_2781_ _2781_/A _2781_/B _3256_/Q _2782_/C vdd gnd OAI21X1
XFILL_3__2902_ gnd vdd FILL
XFILL_0__2084_ gnd vdd FILL
X_1732_ _2444_/C _2700_/B _1751_/B vdd gnd AND2X2
XFILL_8__1788_ gnd vdd FILL
XFILL_8__3527_ gnd vdd FILL
XFILL_6__3591_ gnd vdd FILL
XFILL_6__2611_ gnd vdd FILL
XFILL_3__2833_ gnd vdd FILL
X_3402_ _3442_/B _3403_/A _3466_/B _3403_/C vdd gnd OAI21X1
XFILL_6__2542_ gnd vdd FILL
XFILL_8__3458_ gnd vdd FILL
XFILL_3__2764_ gnd vdd FILL
X_3333_ _3333_/D vdd _3345_/R _3576_/CLK _3333_/Q vdd gnd DFFSR
XFILL_8__3389_ gnd vdd FILL
XFILL_0__2986_ gnd vdd FILL
XFILL_6__2473_ gnd vdd FILL
XFILL_3__1715_ gnd vdd FILL
XFILL_8__2409_ gnd vdd FILL
X_3264_ _3264_/D vdd _3282_/R _3313_/CLK _3264_/Q vdd gnd DFFSR
XFILL_0__1937_ gnd vdd FILL
XFILL_3__2695_ gnd vdd FILL
XFILL_0__1868_ gnd vdd FILL
X_2215_ _2933_/C _2843_/C vdd gnd INVX1
XFILL_1__2400_ gnd vdd FILL
X_3195_ _3195_/A _3195_/B _3196_/B vdd gnd AND2X2
XFILL_1__3380_ gnd vdd FILL
X_2146_ _2276_/A _2781_/B _2341_/A _2147_/C vdd gnd OAI21X1
XFILL_0__1799_ gnd vdd FILL
XFILL_6__3025_ gnd vdd FILL
XFILL_4__2040_ gnd vdd FILL
XFILL_0__3538_ gnd vdd FILL
X_2077_ _2077_/A _2318_/B _2077_/C _2282_/A vdd gnd NAND3X1
XFILL_1__2331_ gnd vdd FILL
XFILL_0__3469_ gnd vdd FILL
XFILL_1__2262_ gnd vdd FILL
XFILL_3__3178_ gnd vdd FILL
XFILL_1__2193_ gnd vdd FILL
XFILL_7__2720_ gnd vdd FILL
XFILL_3__2129_ gnd vdd FILL
XFILL_4__2942_ gnd vdd FILL
X_2979_ _2979_/A _2979_/B _2979_/C _3309_/D vdd gnd OAI21X1
XFILL_7__2651_ gnd vdd FILL
XFILL_6__2809_ gnd vdd FILL
XFILL_4__2873_ gnd vdd FILL
XFILL_7__2582_ gnd vdd FILL
XFILL_4__1824_ gnd vdd FILL
XFILL_4__1755_ gnd vdd FILL
XFILL_1__1977_ gnd vdd FILL
XFILL_7__3203_ gnd vdd FILL
XFILL_7__3134_ gnd vdd FILL
XFILL_4__3425_ gnd vdd FILL
XFILL_2__2440_ gnd vdd FILL
XFILL_2__2371_ gnd vdd FILL
XFILL_5__2080_ gnd vdd FILL
XFILL_7__3065_ gnd vdd FILL
XFILL_4__2307_ gnd vdd FILL
XFILL184650x78150 gnd vdd FILL
XFILL_7__2016_ gnd vdd FILL
XFILL_1__2529_ gnd vdd FILL
XFILL_4__2238_ gnd vdd FILL
XFILL_4__2169_ gnd vdd FILL
XFILL_8__2760_ gnd vdd FILL
XFILL_7__2918_ gnd vdd FILL
XFILL_5__2982_ gnd vdd FILL
XFILL_8__1711_ gnd vdd FILL
XFILL_8__2691_ gnd vdd FILL
XFILL_7__2849_ gnd vdd FILL
XFILL_5__1933_ gnd vdd FILL
XFILL_5__1864_ gnd vdd FILL
XFILL_5__3603_ gnd vdd FILL
XFILL_5__3534_ gnd vdd FILL
XFILL_5__1795_ gnd vdd FILL
XFILL_0__2840_ gnd vdd FILL
XFILL_2_BUFX2_insert6 gnd vdd FILL
XFILL_5__3465_ gnd vdd FILL
XFILL_2__2707_ gnd vdd FILL
XFILL_0__2771_ gnd vdd FILL
XFILL_8__3174_ gnd vdd FILL
XFILL_5__3396_ gnd vdd FILL
XFILL_5__2416_ gnd vdd FILL
XFILL_8__2125_ gnd vdd FILL
XFILL_0__1722_ gnd vdd FILL
XFILL_3__2480_ gnd vdd FILL
X_2000_ _3299_/Q _2001_/A vdd gnd INVX1
XFILL_5__2347_ gnd vdd FILL
XFILL_2__2638_ gnd vdd FILL
XFILL_8__2056_ gnd vdd FILL
XFILL_2__2569_ gnd vdd FILL
XFILL_6_BUFX2_insert20 gnd vdd FILL
XFILL_3__3101_ gnd vdd FILL
XFILL_5__2278_ gnd vdd FILL
XFILL_3__3032_ gnd vdd FILL
XFILL_6_BUFX2_insert42 gnd vdd FILL
XFILL_6_BUFX2_insert53 gnd vdd FILL
XFILL_6_BUFX2_insert97 gnd vdd FILL
X_2902_ _2902_/A _2917_/B _2916_/C _2903_/C vdd gnd OAI21X1
XFILL_6_BUFX2_insert64 gnd vdd FILL
XFILL_6_BUFX2_insert75 gnd vdd FILL
XFILL_6_BUFX2_insert86 gnd vdd FILL
XFILL_0__2205_ gnd vdd FILL
XFILL_8__2958_ gnd vdd FILL
XFILL_9__1751_ gnd vdd FILL
X_2833_ _2833_/A _2837_/C vdd gnd INVX1
XFILL_8__2889_ gnd vdd FILL
XFILL_6__1973_ gnd vdd FILL
XFILL_0__3185_ gnd vdd FILL
XFILL_8__1909_ gnd vdd FILL
XFILL_0__2136_ gnd vdd FILL
X_2764_ _2775_/A _2774_/A _2775_/C _2767_/B vdd gnd NAND3X1
XFILL_0__2067_ gnd vdd FILL
X_1715_ _2594_/B _2123_/B vdd gnd INVX1
X_2695_ _2708_/A _2708_/B _2721_/B _2696_/A vdd gnd AOI21X1
XFILL_1__2880_ gnd vdd FILL
XFILL_3__2816_ gnd vdd FILL
XFILL_1__1900_ gnd vdd FILL
XFILL_1__1831_ gnd vdd FILL
XFILL_6__2525_ gnd vdd FILL
X_3316_ _3316_/D vdd _3345_/R _3577_/CLK _3316_/Q vdd gnd DFFSR
XFILL_6__2456_ gnd vdd FILL
XFILL_1__1762_ gnd vdd FILL
XFILL_3__2747_ gnd vdd FILL
XFILL_1__3501_ gnd vdd FILL
XFILL_0__2969_ gnd vdd FILL
XFILL_3__2678_ gnd vdd FILL
XFILL_6__2387_ gnd vdd FILL
XFILL_4__3210_ gnd vdd FILL
XFILL_1__1693_ gnd vdd FILL
X_3247_ _3247_/D vdd _3291_/R _3362_/CLK _3247_/Q vdd gnd DFFSR
XFILL_4__3141_ gnd vdd FILL
XFILL_1__3432_ gnd vdd FILL
X_3178_ _3185_/B _3178_/B _3179_/B vdd gnd AND2X2
X_2129_ _3197_/C _2759_/A _2129_/C _2331_/A vdd gnd OAI21X1
XFILL_6__3008_ gnd vdd FILL
XFILL_4__3072_ gnd vdd FILL
XFILL_1__2314_ gnd vdd FILL
XFILL_4__2023_ gnd vdd FILL
XFILL_1__2245_ gnd vdd FILL
XFILL_1__2176_ gnd vdd FILL
XFILL_7__2703_ gnd vdd FILL
XFILL_4__2925_ gnd vdd FILL
XFILL_7__2634_ gnd vdd FILL
XFILL_2__1940_ gnd vdd FILL
XFILL_4__2856_ gnd vdd FILL
XFILL_2__1871_ gnd vdd FILL
XFILL_4__1807_ gnd vdd FILL
XFILL_7__2565_ gnd vdd FILL
XFILL_4__2787_ gnd vdd FILL
XFILL_7__2496_ gnd vdd FILL
XFILL_4__1738_ gnd vdd FILL
XFILL_2__3541_ gnd vdd FILL
XFILL_2__3472_ gnd vdd FILL
XFILL_4__3408_ gnd vdd FILL
XFILL_5__2201_ gnd vdd FILL
XFILL_7__3117_ gnd vdd FILL
XFILL_2__2423_ gnd vdd FILL
XFILL_5__3181_ gnd vdd FILL
XFILL_2__2354_ gnd vdd FILL
XFILL_7__3048_ gnd vdd FILL
XFILL_5__2132_ gnd vdd FILL
XFILL_5__2063_ gnd vdd FILL
XFILL_2__2285_ gnd vdd FILL
XFILL_8__2812_ gnd vdd FILL
XFILL_8__2743_ gnd vdd FILL
XFILL_5__2965_ gnd vdd FILL
XFILL_5__1916_ gnd vdd FILL
XFILL_3__1980_ gnd vdd FILL
XFILL_8__2674_ gnd vdd FILL
XFILL_5__2896_ gnd vdd FILL
XFILL183750x101550 gnd vdd FILL
XFILL_5__1847_ gnd vdd FILL
X_2480_ _3351_/Q _2632_/A vdd gnd INVX1
XFILL_5__1778_ gnd vdd FILL
XFILL_3__2601_ gnd vdd FILL
XFILL_5__3517_ gnd vdd FILL
XFILL_0__2823_ gnd vdd FILL
XFILL_6__2310_ gnd vdd FILL
XFILL_3__3581_ gnd vdd FILL
XFILL_8__3226_ gnd vdd FILL
X_3101_ _3115_/A _3107_/B _3327_/Q _3102_/C vdd gnd OAI21X1
XFILL_5__3448_ gnd vdd FILL
XFILL_6__2241_ gnd vdd FILL
XFILL_3__2532_ gnd vdd FILL
XFILL_3__2463_ gnd vdd FILL
XFILL_0__2754_ gnd vdd FILL
XFILL_8__3157_ gnd vdd FILL
X_3032_ _3315_/Q _3090_/A _3033_/C vdd gnd NAND2X1
XFILL_5__3379_ gnd vdd FILL
XFILL_8__3088_ gnd vdd FILL
XFILL_6__2172_ gnd vdd FILL
XFILL_0__1705_ gnd vdd FILL
XFILL_0__2685_ gnd vdd FILL
XFILL_8__2108_ gnd vdd FILL
XFILL_8__2039_ gnd vdd FILL
XFILL_3__2394_ gnd vdd FILL
XFILL_3__3015_ gnd vdd FILL
XFILL_1__2030_ gnd vdd FILL
XFILL_6__1956_ gnd vdd FILL
X_2816_ _2906_/A _2888_/B _3268_/Q _2821_/C vdd gnd OAI21X1
XFILL_0__3168_ gnd vdd FILL
XFILL_0__2119_ gnd vdd FILL
XFILL_0__3099_ gnd vdd FILL
XFILL_6__1887_ gnd vdd FILL
XFILL_4__2710_ gnd vdd FILL
X_2747_ _3575_/Q _2770_/B _3177_/B _2748_/C vdd gnd AOI21X1
XFILL_1__2932_ gnd vdd FILL
X_2678_ _3217_/A _2700_/B _2697_/B _2746_/B _2682_/A vdd gnd OAI22X1
XFILL_6__3557_ gnd vdd FILL
XFILL_7__2350_ gnd vdd FILL
XFILL_4__2641_ gnd vdd FILL
XFILL_1__2863_ gnd vdd FILL
XFILL_2_BUFX2_insert51 gnd vdd FILL
XFILL_2_BUFX2_insert62 gnd vdd FILL
XFILL_2_BUFX2_insert40 gnd vdd FILL
XFILL_4__2572_ gnd vdd FILL
XFILL_6__2508_ gnd vdd FILL
XFILL_6__3488_ gnd vdd FILL
XFILL_2_BUFX2_insert95 gnd vdd FILL
XFILL_2_BUFX2_insert84 gnd vdd FILL
XFILL_1__2794_ gnd vdd FILL
XFILL_2_BUFX2_insert73 gnd vdd FILL
XFILL_7__2281_ gnd vdd FILL
XFILL_1__1814_ gnd vdd FILL
XFILL_1__1745_ gnd vdd FILL
XFILL_6__2439_ gnd vdd FILL
XFILL_1__3415_ gnd vdd FILL
XFILL_4__3124_ gnd vdd FILL
XFILL_4__3055_ gnd vdd FILL
XFILL_4__2006_ gnd vdd FILL
XFILL_2__2070_ gnd vdd FILL
XFILL_1__2228_ gnd vdd FILL
XFILL_7__1996_ gnd vdd FILL
XFILL_1__2159_ gnd vdd FILL
XFILL_5__2750_ gnd vdd FILL
XFILL_4__2908_ gnd vdd FILL
XFILL_2__2972_ gnd vdd FILL
XFILL_5__1701_ gnd vdd FILL
XFILL_8__2390_ gnd vdd FILL
XFILL_7__3597_ gnd vdd FILL
XFILL_2__1923_ gnd vdd FILL
XFILL_5__2681_ gnd vdd FILL
XFILL_7__2617_ gnd vdd FILL
XFILL_4__2839_ gnd vdd FILL
XFILL_7__2548_ gnd vdd FILL
XFILL_2__1854_ gnd vdd FILL
XFILL_7__2479_ gnd vdd FILL
XFILL_2__1785_ gnd vdd FILL
XFILL_0_CLKBUF1_insert35 gnd vdd FILL
XFILL_2__3524_ gnd vdd FILL
XFILL_8__3011_ gnd vdd FILL
XFILL_2__3455_ gnd vdd FILL
XFILL_0__2470_ gnd vdd FILL
XFILL_5__3164_ gnd vdd FILL
XFILL_2__3386_ gnd vdd FILL
XFILL_5__2115_ gnd vdd FILL
XFILL_2__2406_ gnd vdd FILL
XFILL_5__3095_ gnd vdd FILL
XFILL_2__2337_ gnd vdd FILL
X_1980_ _2515_/A _1986_/B vdd gnd INVX1
XFILL_5__2046_ gnd vdd FILL
XFILL_2__2268_ gnd vdd FILL
XFILL_0__3022_ gnd vdd FILL
XFILL_6__1810_ gnd vdd FILL
XFILL_2__2199_ gnd vdd FILL
XFILL_6__2790_ gnd vdd FILL
XFILL_8__2726_ gnd vdd FILL
XFILL_5__2948_ gnd vdd FILL
X_3581_ _3581_/A AB[10] vdd gnd BUFX2
X_2601_ _2601_/A _2601_/B _2601_/C _2612_/C vdd gnd AOI21X1
XFILL_8__2657_ gnd vdd FILL
XFILL_6__1741_ gnd vdd FILL
XFILL_5__2879_ gnd vdd FILL
XFILL_3__1963_ gnd vdd FILL
X_2532_ _3358_/Q _3221_/A vdd gnd INVX1
XFILL_9__3120_ gnd vdd FILL
XFILL_6__3411_ gnd vdd FILL
XFILL_8__2588_ gnd vdd FILL
XFILL_3__1894_ gnd vdd FILL
X_2463_ _3201_/B _3579_/A vdd gnd INVX1
XFILL_3__3564_ gnd vdd FILL
X_2394_ _2872_/B _3077_/C _3249_/Q _2398_/A vdd gnd OAI21X1
XFILL_0__2806_ gnd vdd FILL
XFILL_9__2002_ gnd vdd FILL
XFILL_8__3209_ gnd vdd FILL
XFILL_3__2515_ gnd vdd FILL
XFILL_3__3495_ gnd vdd FILL
XFILL_6__2224_ gnd vdd FILL
XFILL_0__2737_ gnd vdd FILL
X_3015_ _3015_/A _3015_/B _3015_/C _3017_/B vdd gnd OAI21X1
XFILL_6__2155_ gnd vdd FILL
XFILL_3__2446_ gnd vdd FILL
XFILL_3__2377_ gnd vdd FILL
XFILL_0__2668_ gnd vdd FILL
XFILL_6__2086_ gnd vdd FILL
XFILL_0__2599_ gnd vdd FILL
XFILL_1__3200_ gnd vdd FILL
XFILL_1__3131_ gnd vdd FILL
XFILL_1__3062_ gnd vdd FILL
XFILL_7__1850_ gnd vdd FILL
XFILL_1__2013_ gnd vdd FILL
XFILL_6__2988_ gnd vdd FILL
XFILL_7__1781_ gnd vdd FILL
XFILL_6__1939_ gnd vdd FILL
XFILL_7__3520_ gnd vdd FILL
XFILL_7__3451_ gnd vdd FILL
XFILL_7__2402_ gnd vdd FILL
XFILL_1__2915_ gnd vdd FILL
XFILL_7__3382_ gnd vdd FILL
XFILL_4__2624_ gnd vdd FILL
XFILL_1__2846_ gnd vdd FILL
XFILL_7__2333_ gnd vdd FILL
XFILL_7__2264_ gnd vdd FILL
XFILL_4__2555_ gnd vdd FILL
XFILL_4__2486_ gnd vdd FILL
XFILL_1__2777_ gnd vdd FILL
XFILL_7_BUFX2_insert19 gnd vdd FILL
XFILL_7__2195_ gnd vdd FILL
XFILL_1__1728_ gnd vdd FILL
XFILL182250x7950 gnd vdd FILL
XFILL_4__3107_ gnd vdd FILL
XFILL_2__3171_ gnd vdd FILL
XFILL_2__2122_ gnd vdd FILL
XFILL_4__3038_ gnd vdd FILL
XFILL_8__1890_ gnd vdd FILL
XFILL_2__2053_ gnd vdd FILL
XFILL_7__1979_ gnd vdd FILL
XFILL_8__3560_ gnd vdd FILL
XFILL_5__2802_ gnd vdd FILL
XFILL_8__3491_ gnd vdd FILL
XFILL_8__2511_ gnd vdd FILL
XFILL_5__2733_ gnd vdd FILL
XFILL_8__2442_ gnd vdd FILL
XFILL_2__2955_ gnd vdd FILL
XFILL_7_BUFX2_insert1 gnd vdd FILL
XFILL_5__2664_ gnd vdd FILL
XFILL_2__2886_ gnd vdd FILL
XFILL_8__2373_ gnd vdd FILL
XFILL_0__1970_ gnd vdd FILL
XFILL_2__1906_ gnd vdd FILL
XFILL_5__2595_ gnd vdd FILL
XFILL_2__1837_ gnd vdd FILL
XFILL_2__1768_ gnd vdd FILL
XFILL_2__3507_ gnd vdd FILL
XFILL_3__2300_ gnd vdd FILL
XFILL_5__3216_ gnd vdd FILL
XFILL_2__1699_ gnd vdd FILL
XFILL_2__3438_ gnd vdd FILL
XFILL_3__2231_ gnd vdd FILL
XFILL_0__2522_ gnd vdd FILL
XFILL_0__2453_ gnd vdd FILL
XFILL_5__3147_ gnd vdd FILL
XFILL_3__2162_ gnd vdd FILL
XFILL_5__3078_ gnd vdd FILL
XFILL_0__2384_ gnd vdd FILL
XFILL_2__3369_ gnd vdd FILL
XFILL_6__2911_ gnd vdd FILL
XFILL_5__2029_ gnd vdd FILL
XFILL_3__2093_ gnd vdd FILL
X_1963_ _1985_/A _3575_/Q _1963_/C _1964_/C vdd gnd AOI21X1
XFILL_9__2620_ gnd vdd FILL
XFILL_6__2842_ gnd vdd FILL
X_1894_ _3189_/B _3146_/A _1895_/A vdd gnd NAND2X1
XFILL_0__3005_ gnd vdd FILL
XFILL_8__2709_ gnd vdd FILL
XFILL_6__2773_ gnd vdd FILL
XFILL_3__2995_ gnd vdd FILL
XFILL_6__1724_ gnd vdd FILL
XFILL_3__1946_ gnd vdd FILL
X_3564_ _3578_/Q _3566_/B vdd gnd INVX1
X_3495_ _3495_/A _3497_/C _3548_/B vdd gnd NAND2X1
X_2515_ _2515_/A _2519_/C _2515_/C _3215_/B vdd gnd AOI21X1
XFILL_3__1877_ gnd vdd FILL
X_2446_ _2966_/A _2446_/B _2541_/B _2511_/A vdd gnd OAI21X1
XFILL_1__2700_ gnd vdd FILL
XFILL_1__2631_ gnd vdd FILL
XFILL_3__3547_ gnd vdd FILL
XFILL_4__2340_ gnd vdd FILL
X_2377_ _2423_/A _2462_/A _2386_/C vdd gnd NAND2X1
XFILL_3__3478_ gnd vdd FILL
XFILL_4__2271_ gnd vdd FILL
XFILL_6__2207_ gnd vdd FILL
XFILL_1__2562_ gnd vdd FILL
XFILL_1__2493_ gnd vdd FILL
XFILL_6__3187_ gnd vdd FILL
XFILL_3__2429_ gnd vdd FILL
XFILL_6__2138_ gnd vdd FILL
XFILL_7__2951_ gnd vdd FILL
XFILL_6__2069_ gnd vdd FILL
XFILL_7__1902_ gnd vdd FILL
XFILL_1__3114_ gnd vdd FILL
XFILL_7__2882_ gnd vdd FILL
XFILL_1__3045_ gnd vdd FILL
XFILL_7__1833_ gnd vdd FILL
XFILL_7__1764_ gnd vdd FILL
XFILL_7__3503_ gnd vdd FILL
XFILL_4__1986_ gnd vdd FILL
XFILL_7__1695_ gnd vdd FILL
XFILL_7__3434_ gnd vdd FILL
XFILL_2__2740_ gnd vdd FILL
XFILL_7__3365_ gnd vdd FILL
XFILL_4__3587_ gnd vdd FILL
XFILL_5__2380_ gnd vdd FILL
XFILL_7__2316_ gnd vdd FILL
XFILL_4__2607_ gnd vdd FILL
XFILL_2__2671_ gnd vdd FILL
XFILL_1__2829_ gnd vdd FILL
XFILL_4__2538_ gnd vdd FILL
XFILL_7__2247_ gnd vdd FILL
XFILL_5__3001_ gnd vdd FILL
XFILL_4__2469_ gnd vdd FILL
XFILL_7__2178_ gnd vdd FILL
XFILL_2__3223_ gnd vdd FILL
XFILL_8__2991_ gnd vdd FILL
XFILL_8__1942_ gnd vdd FILL
XFILL_2__3154_ gnd vdd FILL
XFILL_8__1873_ gnd vdd FILL
XFILL_2__3085_ gnd vdd FILL
XFILL_2__2105_ gnd vdd FILL
XFILL_2__2036_ gnd vdd FILL
XFILL_8__3543_ gnd vdd FILL
XFILL_3_BUFX2_insert17 gnd vdd FILL
XFILL_8__3474_ gnd vdd FILL
XFILL_5__2716_ gnd vdd FILL
XFILL_3_BUFX2_insert39 gnd vdd FILL
XFILL_3__2780_ gnd vdd FILL
XFILL_3__1800_ gnd vdd FILL
XFILL_8__2425_ gnd vdd FILL
XFILL_2__2938_ gnd vdd FILL
XFILL_3__1731_ gnd vdd FILL
X_3280_ _3280_/D vdd _3282_/R _3284_/CLK _3280_/Q vdd gnd DFFSR
XFILL_8__2356_ gnd vdd FILL
XFILL_0__1953_ gnd vdd FILL
X_2300_ _2341_/A _3017_/A _2300_/C _2345_/A vdd gnd OAI21X1
XFILL_5__2647_ gnd vdd FILL
XFILL_5__2578_ gnd vdd FILL
XFILL_2__2869_ gnd vdd FILL
X_2231_ _3166_/C _3166_/D _2586_/B vdd gnd NAND2X1
XFILL_6__3110_ gnd vdd FILL
XFILL_3__3401_ gnd vdd FILL
XFILL_8__2287_ gnd vdd FILL
XFILL_0__1884_ gnd vdd FILL
X_2162_ _2889_/C _2889_/A _2910_/B vdd gnd NAND2X1
XFILL_0__3554_ gnd vdd FILL
XFILL_6__3041_ gnd vdd FILL
X_2093_ _2293_/A _2229_/A _2094_/C vdd gnd NAND2X1
XFILL_0__2505_ gnd vdd FILL
XFILL_0__3485_ gnd vdd FILL
XFILL_3__2214_ gnd vdd FILL
XFILL_3__3194_ gnd vdd FILL
XFILL_3__2145_ gnd vdd FILL
XFILL_0__2436_ gnd vdd FILL
XFILL_0__2367_ gnd vdd FILL
XFILL_0__2298_ gnd vdd FILL
X_2995_ _2995_/A _3011_/B _2995_/C _2996_/C vdd gnd OAI21X1
XFILL_3__2076_ gnd vdd FILL
XFILL_6__2825_ gnd vdd FILL
X_1946_ _1986_/A _1946_/B _1946_/C _3434_/A vdd gnd OAI21X1
X_1877_ _3315_/Q _3029_/B _1881_/B vdd gnd NAND2X1
XFILL_4__1840_ gnd vdd FILL
XFILL_6__2756_ gnd vdd FILL
X_3547_ _3571_/Q _3550_/A _3548_/C vdd gnd NAND2X1
XFILL_4__3510_ gnd vdd FILL
XFILL_3__2978_ gnd vdd FILL
XFILL_4__1771_ gnd vdd FILL
XFILL_6__1707_ gnd vdd FILL
XFILL_6__2687_ gnd vdd FILL
XFILL_3__1929_ gnd vdd FILL
XFILL_1__1993_ gnd vdd FILL
X_3478_ _3514_/A _3482_/B _3479_/A vdd gnd NAND2X1
XFILL_4__3441_ gnd vdd FILL
XFILL_7__3150_ gnd vdd FILL
XFILL_4__3372_ gnd vdd FILL
XFILL_7__2101_ gnd vdd FILL
X_2429_ _2429_/A _2431_/A vdd gnd INVX1
XFILL_7__3081_ gnd vdd FILL
XFILL_9__3017_ gnd vdd FILL
XFILL_4__2323_ gnd vdd FILL
XFILL_1__3594_ gnd vdd FILL
XFILL_1__2614_ gnd vdd FILL
XFILL_7__2032_ gnd vdd FILL
XFILL_1__2545_ gnd vdd FILL
XFILL_4__2254_ gnd vdd FILL
XFILL_4__2185_ gnd vdd FILL
XFILL_1__2476_ gnd vdd FILL
XFILL_7__2934_ gnd vdd FILL
XFILL_7__2865_ gnd vdd FILL
XFILL_5__1880_ gnd vdd FILL
XFILL_7__1816_ gnd vdd FILL
XFILL_1__3028_ gnd vdd FILL
XFILL_7__2796_ gnd vdd FILL
XFILL_7__1747_ gnd vdd FILL
XFILL_5_CLKBUF1_insert35 gnd vdd FILL
XFILL_5__3550_ gnd vdd FILL
XFILL_4__1969_ gnd vdd FILL
XFILL_5__3481_ gnd vdd FILL
XFILL_7__3417_ gnd vdd FILL
XFILL_8__2210_ gnd vdd FILL
XFILL_5__2501_ gnd vdd FILL
XFILL_2__2723_ gnd vdd FILL
XFILL_5__2432_ gnd vdd FILL
XFILL_8__3190_ gnd vdd FILL
XFILL_8__2141_ gnd vdd FILL
XFILL_2__2654_ gnd vdd FILL
XFILL_8__2072_ gnd vdd FILL
XFILL_5__2363_ gnd vdd FILL
XFILL_2__2585_ gnd vdd FILL
XFILL_5__2294_ gnd vdd FILL
XFILL_8__2974_ gnd vdd FILL
XFILL184050x4050 gnd vdd FILL
XFILL_2__3206_ gnd vdd FILL
XFILL_2__3137_ gnd vdd FILL
XFILL_8__1925_ gnd vdd FILL
XFILL_0__2221_ gnd vdd FILL
XFILL_0__2152_ gnd vdd FILL
X_1800_ _3148_/B _3182_/C vdd gnd INVX1
XFILL_2__3068_ gnd vdd FILL
XFILL_8__1856_ gnd vdd FILL
X_2780_ NMI _2780_/B _2782_/B vdd gnd NAND2X1
XFILL_0__2083_ gnd vdd FILL
XFILL_3__2901_ gnd vdd FILL
XFILL_2__2019_ gnd vdd FILL
X_1731_ _2063_/B _2279_/A _2444_/C vdd gnd NOR2X1
XFILL_6__2610_ gnd vdd FILL
XFILL_8__1787_ gnd vdd FILL
XFILL_8__3526_ gnd vdd FILL
XFILL_3__2832_ gnd vdd FILL
XFILL_6__3590_ gnd vdd FILL
X_3401_ _3514_/B _3466_/B vdd gnd INVX2
XFILL_8__3457_ gnd vdd FILL
XFILL_6__2541_ gnd vdd FILL
X_3332_ _3332_/D vdd _3347_/R _3576_/CLK _3332_/Q vdd gnd DFFSR
XFILL_6__2472_ gnd vdd FILL
XFILL_3__2763_ gnd vdd FILL
XFILL_8__3388_ gnd vdd FILL
XFILL_0__2985_ gnd vdd FILL
XFILL_3__2694_ gnd vdd FILL
XFILL_3__1714_ gnd vdd FILL
XFILL_8__2408_ gnd vdd FILL
X_3263_ _3263_/D vdd _3289_/R _3313_/CLK _3263_/Q vdd gnd DFFSR
XFILL_0__1936_ gnd vdd FILL
XFILL_8__2339_ gnd vdd FILL
XFILL_0__1867_ gnd vdd FILL
X_2214_ _2298_/A _3177_/A _2214_/C _2298_/D _2327_/A vdd gnd AOI22X1
X_3194_ _3194_/A _3194_/B _3194_/C _3195_/A vdd gnd OAI21X1
X_2145_ _3088_/S _3077_/C vdd gnd INVX4
XFILL_6__3024_ gnd vdd FILL
XFILL_0__1798_ gnd vdd FILL
XFILL_0__3537_ gnd vdd FILL
X_2076_ _2318_/C _2318_/A _2077_/C vdd gnd AND2X2
XFILL_1__2330_ gnd vdd FILL
XFILL_0__3468_ gnd vdd FILL
XFILL_1__2261_ gnd vdd FILL
XFILL_0__2419_ gnd vdd FILL
XFILL_1__2192_ gnd vdd FILL
XFILL_3__3177_ gnd vdd FILL
XFILL_0__3399_ gnd vdd FILL
XFILL_3__2128_ gnd vdd FILL
XFILL_4__2941_ gnd vdd FILL
X_2978_ _3293_/D _2978_/B _3017_/A _2979_/B vdd gnd MUX2X1
XFILL_3__2059_ gnd vdd FILL
X_1929_ _3333_/Q _3110_/A _3127_/B _3342_/Q _1931_/C vdd gnd AOI22X1
XFILL_7__2650_ gnd vdd FILL
XFILL_6__2808_ gnd vdd FILL
XFILL_4__2872_ gnd vdd FILL
XFILL_9__2517_ gnd vdd FILL
XFILL_7__2581_ gnd vdd FILL
XFILL_4__1823_ gnd vdd FILL
XFILL_6__2739_ gnd vdd FILL
XFILL_4__1754_ gnd vdd FILL
XFILL_1__1976_ gnd vdd FILL
XFILL_7__3202_ gnd vdd FILL
XFILL_4__3424_ gnd vdd FILL
XFILL_7__3133_ gnd vdd FILL
XFILL_7__3064_ gnd vdd FILL
XFILL_2__2370_ gnd vdd FILL
XFILL_4__2306_ gnd vdd FILL
XFILL_7__2015_ gnd vdd FILL
XFILL_4__2237_ gnd vdd FILL
XFILL_1__2528_ gnd vdd FILL
XFILL_1__2459_ gnd vdd FILL
XFILL_4__2168_ gnd vdd FILL
XFILL_5__2981_ gnd vdd FILL
XFILL_8__1710_ gnd vdd FILL
XFILL_4__2099_ gnd vdd FILL
XFILL_7__2917_ gnd vdd FILL
XFILL_5__1932_ gnd vdd FILL
XFILL_8__2690_ gnd vdd FILL
XFILL_7__2848_ gnd vdd FILL
XFILL_5__1863_ gnd vdd FILL
XFILL_7__2779_ gnd vdd FILL
XFILL_5__3602_ gnd vdd FILL
XFILL_5__1794_ gnd vdd FILL
XFILL_5__3533_ gnd vdd FILL
XFILL_2_BUFX2_insert7 gnd vdd FILL
XFILL_5__3464_ gnd vdd FILL
XFILL_2__2706_ gnd vdd FILL
XFILL_0__2770_ gnd vdd FILL
XFILL_8__3173_ gnd vdd FILL
XFILL_5__3395_ gnd vdd FILL
XFILL_5__2415_ gnd vdd FILL
XFILL_8__2124_ gnd vdd FILL
XFILL_0__1721_ gnd vdd FILL
XFILL181650x148350 gnd vdd FILL
XFILL_5__2346_ gnd vdd FILL
XFILL_2__2637_ gnd vdd FILL
XFILL_8__2055_ gnd vdd FILL
XFILL_2__2568_ gnd vdd FILL
XFILL_3__3100_ gnd vdd FILL
XFILL_6_BUFX2_insert21 gnd vdd FILL
XFILL_6_BUFX2_insert10 gnd vdd FILL
XFILL_5__2277_ gnd vdd FILL
XFILL_3__3031_ gnd vdd FILL
XFILL_2__2499_ gnd vdd FILL
XFILL_6_BUFX2_insert43 gnd vdd FILL
XFILL_6_BUFX2_insert54 gnd vdd FILL
X_2901_ _2901_/A _2933_/A _2917_/B vdd gnd OR2X2
XFILL_6_BUFX2_insert87 gnd vdd FILL
XFILL_6_BUFX2_insert65 gnd vdd FILL
XFILL_6_BUFX2_insert76 gnd vdd FILL
XFILL_8__2957_ gnd vdd FILL
XFILL_0__2204_ gnd vdd FILL
X_2832_ _2910_/B _2832_/B _2832_/C _2833_/A vdd gnd OAI21X1
XFILL_8__2888_ gnd vdd FILL
XFILL_6__1972_ gnd vdd FILL
XFILL_0__3184_ gnd vdd FILL
XFILL_8__1908_ gnd vdd FILL
XFILL_8__1839_ gnd vdd FILL
XFILL_0__2135_ gnd vdd FILL
X_2763_ _2766_/B _2766_/A _2774_/A vdd gnd NOR2X1
XFILL_0__2066_ gnd vdd FILL
X_1714_ _3235_/Q _1793_/B _2594_/B vdd gnd NAND2X1
X_2694_ _2741_/B _2741_/C _2721_/B vdd gnd NOR2X1
XFILL_8__3509_ gnd vdd FILL
XFILL_3__2815_ gnd vdd FILL
XFILL_6__2524_ gnd vdd FILL
XFILL_3__2746_ gnd vdd FILL
XFILL_1__1830_ gnd vdd FILL
XFILL_9__2164_ gnd vdd FILL
X_3315_ _3315_/D vdd _3353_/R _3577_/CLK _3315_/Q vdd gnd DFFSR
XFILL_0__2968_ gnd vdd FILL
XFILL_6__2455_ gnd vdd FILL
XFILL_1__1761_ gnd vdd FILL
XFILL_1__3500_ gnd vdd FILL
XFILL_0__1919_ gnd vdd FILL
XFILL_6__2386_ gnd vdd FILL
XFILL_3__2677_ gnd vdd FILL
X_3246_ _3246_/D vdd _3362_/R _3362_/CLK _3246_/Q vdd gnd DFFSR
XFILL_0__2899_ gnd vdd FILL
XFILL_1__1692_ gnd vdd FILL
XFILL_4__3140_ gnd vdd FILL
XFILL_1__3431_ gnd vdd FILL
X_3177_ _3177_/A _3177_/B _3185_/B vdd gnd NOR2X1
X_2128_ _2594_/A _2594_/B _3147_/A _2759_/A vdd gnd NOR3X1
XFILL_6__3007_ gnd vdd FILL
XFILL_1__2313_ gnd vdd FILL
XFILL_4__3071_ gnd vdd FILL
X_2059_ _3160_/C _3190_/B _3160_/B _2060_/B vdd gnd OAI21X1
XFILL_4__2022_ gnd vdd FILL
XFILL_3__3229_ gnd vdd FILL
XFILL_1__2244_ gnd vdd FILL
XFILL_1__2175_ gnd vdd FILL
XFILL_7__2702_ gnd vdd FILL
XFILL_4__2924_ gnd vdd FILL
XFILL_7__2633_ gnd vdd FILL
XFILL_4__2855_ gnd vdd FILL
XFILL_2__1870_ gnd vdd FILL
XFILL_7__2564_ gnd vdd FILL
XFILL_4__1806_ gnd vdd FILL
XFILL_4__2786_ gnd vdd FILL
XFILL_7__2495_ gnd vdd FILL
XFILL_2__3540_ gnd vdd FILL
XFILL_4__1737_ gnd vdd FILL
XFILL_1__1959_ gnd vdd FILL
XFILL_2__3471_ gnd vdd FILL
XFILL_7__3116_ gnd vdd FILL
XFILL_4__3407_ gnd vdd FILL
XFILL_5__2200_ gnd vdd FILL
XFILL_5__3180_ gnd vdd FILL
XFILL_2__2422_ gnd vdd FILL
XFILL_5__2131_ gnd vdd FILL
XFILL_7__3047_ gnd vdd FILL
XFILL_2__2353_ gnd vdd FILL
XFILL_5__2062_ gnd vdd FILL
XFILL_2__2284_ gnd vdd FILL
XFILL_8__2811_ gnd vdd FILL
XFILL_8__2742_ gnd vdd FILL
XFILL_5__2964_ gnd vdd FILL
XFILL_8__2673_ gnd vdd FILL
XFILL_5__2895_ gnd vdd FILL
XFILL_5__1915_ gnd vdd FILL
XFILL_5__1846_ gnd vdd FILL
XFILL_5__1777_ gnd vdd FILL
XFILL_3__2600_ gnd vdd FILL
XFILL_5__3516_ gnd vdd FILL
XFILL_2__1999_ gnd vdd FILL
XFILL_0__2822_ gnd vdd FILL
XFILL_3__3580_ gnd vdd FILL
XFILL_8__3225_ gnd vdd FILL
X_3100_ _3135_/A _3108_/B _3100_/C _3326_/D vdd gnd OAI21X1
XFILL_5__3447_ gnd vdd FILL
XFILL_6__2240_ gnd vdd FILL
XFILL_3__2531_ gnd vdd FILL
XFILL_3__2462_ gnd vdd FILL
XFILL_0__2753_ gnd vdd FILL
XFILL_8__3156_ gnd vdd FILL
XFILL_5__3378_ gnd vdd FILL
X_3031_ _3290_/D _3088_/S _3031_/C _3129_/A vdd gnd OAI21X1
XFILL_6__2171_ gnd vdd FILL
XFILL_8__3087_ gnd vdd FILL
XFILL_0__1704_ gnd vdd FILL
XFILL_8__2107_ gnd vdd FILL
XFILL_0__2684_ gnd vdd FILL
XFILL_8__2038_ gnd vdd FILL
XFILL_3__2393_ gnd vdd FILL
XFILL_5__2329_ gnd vdd FILL
XFILL_3__3014_ gnd vdd FILL
XFILL_9__2782_ gnd vdd FILL
X_2815_ _2815_/A _2815_/B _2815_/C _3267_/D vdd gnd OAI21X1
XFILL_6__1955_ gnd vdd FILL
XFILL_0__3167_ gnd vdd FILL
XFILL_0__2118_ gnd vdd FILL
XFILL_0__3098_ gnd vdd FILL
XFILL_6__1886_ gnd vdd FILL
X_2746_ _2751_/A _2746_/B _2746_/C _2749_/B vdd gnd OAI21X1
XFILL_1__2931_ gnd vdd FILL
XFILL_0__2049_ gnd vdd FILL
X_2677_ _2726_/C _2699_/B _3016_/A _2682_/C vdd gnd AOI21X1
XFILL_4__2640_ gnd vdd FILL
XFILL_1__2862_ gnd vdd FILL
XFILL_6__3556_ gnd vdd FILL
XFILL_6__3487_ gnd vdd FILL
XFILL_2_BUFX2_insert63 gnd vdd FILL
XFILL_7__2280_ gnd vdd FILL
XFILL_6__2507_ gnd vdd FILL
XFILL_2_BUFX2_insert52 gnd vdd FILL
XFILL_4__2571_ gnd vdd FILL
XFILL_1__1813_ gnd vdd FILL
XFILL_2_BUFX2_insert41 gnd vdd FILL
XFILL_2_BUFX2_insert96 gnd vdd FILL
XFILL_2_BUFX2_insert85 gnd vdd FILL
XFILL_2_BUFX2_insert74 gnd vdd FILL
XFILL_1__2793_ gnd vdd FILL
XFILL_3__2729_ gnd vdd FILL
XFILL_6__2438_ gnd vdd FILL
XFILL_1__1744_ gnd vdd FILL
XFILL_6__2369_ gnd vdd FILL
X_3229_ _3585_/A _3230_/B _3230_/C vdd gnd NAND2X1
XFILL_1__3414_ gnd vdd FILL
XFILL_4__3123_ gnd vdd FILL
XFILL_4__3054_ gnd vdd FILL
XFILL_4__2005_ gnd vdd FILL
XFILL_1__2227_ gnd vdd FILL
XFILL_7__1995_ gnd vdd FILL
XFILL_1__2158_ gnd vdd FILL
XFILL_4__2907_ gnd vdd FILL
XFILL_5__1700_ gnd vdd FILL
XFILL_2__2971_ gnd vdd FILL
XFILL_1__2089_ gnd vdd FILL
XFILL_7__3596_ gnd vdd FILL
XFILL_2__1922_ gnd vdd FILL
XFILL_5__2680_ gnd vdd FILL
XFILL_7__2616_ gnd vdd FILL
XFILL_4__2838_ gnd vdd FILL
XFILL_7__2547_ gnd vdd FILL
XFILL_2__1853_ gnd vdd FILL
XFILL_4__2769_ gnd vdd FILL
XFILL_8__3010_ gnd vdd FILL
XFILL_7__2478_ gnd vdd FILL
XFILL_2__1784_ gnd vdd FILL
XFILL_2__3523_ gnd vdd FILL
XFILL_0_CLKBUF1_insert36 gnd vdd FILL
XFILL_5__3232_ gnd vdd FILL
XFILL_2__3454_ gnd vdd FILL
XFILL_2__2405_ gnd vdd FILL
XFILL_5__3163_ gnd vdd FILL
XFILL_5__3094_ gnd vdd FILL
XFILL_2__3385_ gnd vdd FILL
XFILL_5__2114_ gnd vdd FILL
XFILL_5__2045_ gnd vdd FILL
XFILL_2__2336_ gnd vdd FILL
XFILL_2__2267_ gnd vdd FILL
XFILL_0__3021_ gnd vdd FILL
XFILL_2__2198_ gnd vdd FILL
XFILL_8__2725_ gnd vdd FILL
XFILL_6__1740_ gnd vdd FILL
XFILL_5__2947_ gnd vdd FILL
XFILL_3__1962_ gnd vdd FILL
X_3580_ _3580_/A AB[1] vdd gnd BUFX2
X_2600_ _2612_/B _2756_/B _2601_/B vdd gnd NAND2X1
XFILL_8__2656_ gnd vdd FILL
XFILL_5__2878_ gnd vdd FILL
X_2531_ _3249_/Q _2715_/A vdd gnd INVX1
XFILL_6__3410_ gnd vdd FILL
XFILL_5__1829_ gnd vdd FILL
XFILL_8__2587_ gnd vdd FILL
XFILL_3__1893_ gnd vdd FILL
XFILL183150x148350 gnd vdd FILL
X_2462_ _2462_/A _2519_/C _2462_/C _3201_/B vdd gnd AOI21X1
XFILL_3__3563_ gnd vdd FILL
X_2393_ _2423_/A _2474_/A _2398_/C vdd gnd NAND2X1
XFILL_0__2805_ gnd vdd FILL
XFILL_8__3208_ gnd vdd FILL
XFILL_3__2514_ gnd vdd FILL
XFILL_3__3494_ gnd vdd FILL
XFILL_8__3139_ gnd vdd FILL
XFILL_0__2736_ gnd vdd FILL
XFILL_6__2223_ gnd vdd FILL
X_3014_ _3568_/Q _3015_/A _3015_/C vdd gnd NAND2X1
XFILL_6__2154_ gnd vdd FILL
XFILL_3__2445_ gnd vdd FILL
XFILL_3__2376_ gnd vdd FILL
XFILL_0__2667_ gnd vdd FILL
XFILL_6__2085_ gnd vdd FILL
XFILL_0__2598_ gnd vdd FILL
XFILL_1__3130_ gnd vdd FILL
XFILL_1__3061_ gnd vdd FILL
XFILL_1__2012_ gnd vdd FILL
XFILL_0__3219_ gnd vdd FILL
XFILL_6__2987_ gnd vdd FILL
XFILL_7__1780_ gnd vdd FILL
XFILL_6__1938_ gnd vdd FILL
XFILL_7__3450_ gnd vdd FILL
XFILL_6__1869_ gnd vdd FILL
X_2729_ _3293_/D _2772_/B _2729_/C _2730_/C vdd gnd AOI21X1
XFILL_1__2914_ gnd vdd FILL
XFILL_7__3381_ gnd vdd FILL
XFILL_7__2401_ gnd vdd FILL
XFILL_7__2332_ gnd vdd FILL
XFILL_4__2623_ gnd vdd FILL
XFILL_1__2845_ gnd vdd FILL
XFILL_6__3539_ gnd vdd FILL
XFILL_4__2554_ gnd vdd FILL
XFILL_7__2263_ gnd vdd FILL
XFILL_1__2776_ gnd vdd FILL
XFILL_7__2194_ gnd vdd FILL
XFILL_4__2485_ gnd vdd FILL
XFILL_1__1727_ gnd vdd FILL
XFILL_9__3179_ gnd vdd FILL
XFILL_4__3106_ gnd vdd FILL
XFILL_2__3170_ gnd vdd FILL
XFILL_2__2121_ gnd vdd FILL
XFILL_4__3037_ gnd vdd FILL
XFILL_2__2052_ gnd vdd FILL
XFILL_7__1978_ gnd vdd FILL
XFILL_5__2801_ gnd vdd FILL
XFILL_8__3490_ gnd vdd FILL
XFILL_8__2510_ gnd vdd FILL
XFILL_5__2732_ gnd vdd FILL
XFILL_8__2441_ gnd vdd FILL
XFILL_2__2954_ gnd vdd FILL
XFILL_7_BUFX2_insert2 gnd vdd FILL
XFILL_5__2663_ gnd vdd FILL
XFILL_8__2372_ gnd vdd FILL
XFILL_2__2885_ gnd vdd FILL
XFILL_7__3579_ gnd vdd FILL
XFILL_2__1905_ gnd vdd FILL
XFILL_2__1836_ gnd vdd FILL
XFILL_5__2594_ gnd vdd FILL
XFILL_2__1767_ gnd vdd FILL
XFILL_2__3506_ gnd vdd FILL
XFILL_5__3215_ gnd vdd FILL
XFILL_0__2521_ gnd vdd FILL
XFILL_2__1698_ gnd vdd FILL
XFILL_2__3437_ gnd vdd FILL
XFILL_5__3146_ gnd vdd FILL
XFILL_3__2230_ gnd vdd FILL
XFILL_3__2161_ gnd vdd FILL
XFILL_2__3368_ gnd vdd FILL
XFILL_0__2452_ gnd vdd FILL
XFILL_5__3077_ gnd vdd FILL
XFILL_0__2383_ gnd vdd FILL
XFILL_2__2319_ gnd vdd FILL
XFILL_6__2910_ gnd vdd FILL
XFILL_5__2028_ gnd vdd FILL
XFILL_3__2092_ gnd vdd FILL
X_1962_ _2952_/A _1984_/B _2746_/C _1963_/C vdd gnd OAI21X1
XFILL_6__2841_ gnd vdd FILL
X_1893_ _3182_/B _3146_/A vdd gnd INVX2
XFILL_0__3004_ gnd vdd FILL
XFILL_8__2708_ gnd vdd FILL
XFILL_6__2772_ gnd vdd FILL
XFILL_3__2994_ gnd vdd FILL
XFILL_6__1723_ gnd vdd FILL
X_3563_ _3563_/A _3566_/A _3563_/C _3577_/D vdd gnd OAI21X1
XFILL_3__1945_ gnd vdd FILL
XFILL_8__2639_ gnd vdd FILL
X_3494_ _3494_/A _3494_/B _3495_/A vdd gnd NAND2X1
XFILL_3__1876_ gnd vdd FILL
X_2514_ _2676_/B _2574_/B _2514_/C _2515_/C vdd gnd OAI21X1
X_2445_ _2569_/A _2569_/B _2541_/B vdd gnd NOR2X1
XFILL_1__2630_ gnd vdd FILL
XFILL_3__3546_ gnd vdd FILL
X_2376_ _2376_/A _2423_/A _3603_/A vdd gnd NAND2X1
XFILL_3__3477_ gnd vdd FILL
XFILL_4__2270_ gnd vdd FILL
XFILL_6__2206_ gnd vdd FILL
XFILL_1__2561_ gnd vdd FILL
XFILL_3__2428_ gnd vdd FILL
XFILL_1__2492_ gnd vdd FILL
XFILL_0__2719_ gnd vdd FILL
XFILL_6__3186_ gnd vdd FILL
XFILL_6__2137_ gnd vdd FILL
XFILL_3__2359_ gnd vdd FILL
XFILL_7__2950_ gnd vdd FILL
XFILL_6__2068_ gnd vdd FILL
XFILL_1__3113_ gnd vdd FILL
XFILL_7__1901_ gnd vdd FILL
XFILL_7__2881_ gnd vdd FILL
XFILL_1__3044_ gnd vdd FILL
XFILL_7__1832_ gnd vdd FILL
XFILL_7__1763_ gnd vdd FILL
XFILL_7__3502_ gnd vdd FILL
XFILL_4__1985_ gnd vdd FILL
XFILL_9__2679_ gnd vdd FILL
XFILL_7__1694_ gnd vdd FILL
XFILL_7__3433_ gnd vdd FILL
XFILL_7__3364_ gnd vdd FILL
XFILL_2__2670_ gnd vdd FILL
XFILL_1__2828_ gnd vdd FILL
XFILL_7__2315_ gnd vdd FILL
XFILL_4__3586_ gnd vdd FILL
XFILL_4__2606_ gnd vdd FILL
XFILL_7__2246_ gnd vdd FILL
XFILL_4__2537_ gnd vdd FILL
XFILL_4__2468_ gnd vdd FILL
XFILL_1__2759_ gnd vdd FILL
XFILL_5__3000_ gnd vdd FILL
XFILL_7__2177_ gnd vdd FILL
XFILL_4__2399_ gnd vdd FILL
XFILL_2__3222_ gnd vdd FILL
XFILL_8__2990_ gnd vdd FILL
XFILL_8__1941_ gnd vdd FILL
XFILL_2__3153_ gnd vdd FILL
XFILL_2__2104_ gnd vdd FILL
XFILL_8__1872_ gnd vdd FILL
XFILL_2__3084_ gnd vdd FILL
XFILL_2__2035_ gnd vdd FILL
XFILL_8__3542_ gnd vdd FILL
XFILL_3_BUFX2_insert18 gnd vdd FILL
XFILL_8__3473_ gnd vdd FILL
XFILL_5__2715_ gnd vdd FILL
XFILL_8__2424_ gnd vdd FILL
XFILL_3__1730_ gnd vdd FILL
XFILL_2__2937_ gnd vdd FILL
XFILL_8__2355_ gnd vdd FILL
XFILL_0__1952_ gnd vdd FILL
XFILL_5__2646_ gnd vdd FILL
XFILL_2__2868_ gnd vdd FILL
XFILL_3__3400_ gnd vdd FILL
XFILL_5__2577_ gnd vdd FILL
X_2230_ _3149_/C _3146_/A _3160_/A _2234_/B vdd gnd OAI21X1
XFILL_2__2799_ gnd vdd FILL
XFILL_2__1819_ gnd vdd FILL
XFILL_8__2286_ gnd vdd FILL
XFILL_0__1883_ gnd vdd FILL
X_2161_ _2161_/A _2161_/B _2889_/C _2823_/B vdd gnd OAI21X1
XFILL_6__3040_ gnd vdd FILL
XFILL_0__3553_ gnd vdd FILL
X_2092_ _2292_/B _3189_/A _2229_/A vdd gnd NOR2X1
XFILL_0__3484_ gnd vdd FILL
XFILL_3__2213_ gnd vdd FILL
XFILL_0__2504_ gnd vdd FILL
XFILL_5__3129_ gnd vdd FILL
XFILL_3__3193_ gnd vdd FILL
XFILL_0__2435_ gnd vdd FILL
XFILL_3__2144_ gnd vdd FILL
X_2994_ _3577_/Q _2995_/C vdd gnd INVX1
XFILL_3__2075_ gnd vdd FILL
XFILL_0__2366_ gnd vdd FILL
XFILL_0__2297_ gnd vdd FILL
X_1945_ _1985_/A _3573_/Q _1945_/C _1946_/C vdd gnd AOI21X1
XFILL_6__2824_ gnd vdd FILL
X_1876_ _1879_/B _1879_/A _1878_/A _3029_/B vdd gnd AOI21X1
XFILL_4__1770_ gnd vdd FILL
XFILL_6__2755_ gnd vdd FILL
X_3546_ _3546_/A _3546_/B _3546_/C _3570_/D vdd gnd OAI21X1
XFILL_3__2977_ gnd vdd FILL
XFILL_1__1992_ gnd vdd FILL
XFILL_6__1706_ gnd vdd FILL
XFILL_6__2686_ gnd vdd FILL
XFILL_3__1928_ gnd vdd FILL
XFILL_3__1859_ gnd vdd FILL
X_3477_ _3482_/B _3482_/A _3480_/C vdd gnd NAND2X1
XFILL_4__3440_ gnd vdd FILL
XFILL_4__3371_ gnd vdd FILL
X_2428_ _2428_/A _2428_/B _2428_/C _3602_/A vdd gnd NAND3X1
XFILL_7__2100_ gnd vdd FILL
X_2359_ _2837_/A _2579_/B _2361_/C _3468_/S vdd gnd OAI21X1
XFILL_7__3080_ gnd vdd FILL
XFILL_3__3529_ gnd vdd FILL
XFILL_4__2322_ gnd vdd FILL
XFILL_1__3593_ gnd vdd FILL
XFILL_1__2613_ gnd vdd FILL
XFILL_7__2031_ gnd vdd FILL
XFILL_1__2544_ gnd vdd FILL
XFILL_4__2253_ gnd vdd FILL
XFILL_6__3169_ gnd vdd FILL
XFILL_1__2475_ gnd vdd FILL
XFILL_4__2184_ gnd vdd FILL
XFILL_7__2933_ gnd vdd FILL
XFILL_7__2864_ gnd vdd FILL
XFILL_1__3027_ gnd vdd FILL
XFILL_7__1815_ gnd vdd FILL
XFILL_7__2795_ gnd vdd FILL
XFILL_7__1746_ gnd vdd FILL
XFILL_4__1968_ gnd vdd FILL
XFILL_5_CLKBUF1_insert36 gnd vdd FILL
XFILL_5__3480_ gnd vdd FILL
XFILL_7__3416_ gnd vdd FILL
XFILL_4__1899_ gnd vdd FILL
XFILL_5__2500_ gnd vdd FILL
XFILL_2__2722_ gnd vdd FILL
XFILL_8__2140_ gnd vdd FILL
XFILL_5__2431_ gnd vdd FILL
XFILL_5__2362_ gnd vdd FILL
XFILL_2__2653_ gnd vdd FILL
XFILL_8__2071_ gnd vdd FILL
XFILL_2__2584_ gnd vdd FILL
XFILL_7__2229_ gnd vdd FILL
XFILL_5__2293_ gnd vdd FILL
XFILL_8__2973_ gnd vdd FILL
XFILL_2__3205_ gnd vdd FILL
XFILL_2__3136_ gnd vdd FILL
XFILL_0__2220_ gnd vdd FILL
XFILL_8__1924_ gnd vdd FILL
XFILL_0__2151_ gnd vdd FILL
XFILL_2__3067_ gnd vdd FILL
XFILL_8__1855_ gnd vdd FILL
XFILL_3__2900_ gnd vdd FILL
XFILL_2__2018_ gnd vdd FILL
XFILL_0__2082_ gnd vdd FILL
X_1730_ _2453_/A _3147_/B _2063_/B vdd gnd NOR2X1
XFILL_8__1786_ gnd vdd FILL
XFILL_8__3525_ gnd vdd FILL
XFILL_3__2831_ gnd vdd FILL
XFILL_8__3456_ gnd vdd FILL
X_3400_ _3514_/B _3514_/A _3428_/B vdd gnd NAND2X1
XFILL_6__2540_ gnd vdd FILL
X_3331_ _3331_/D vdd _3346_/R _3346_/CLK _3331_/Q vdd gnd DFFSR
XFILL_6__2471_ gnd vdd FILL
XFILL_3__2762_ gnd vdd FILL
XFILL_8__2407_ gnd vdd FILL
XFILL_8__3387_ gnd vdd FILL
XFILL_0__2984_ gnd vdd FILL
XFILL_3__2693_ gnd vdd FILL
XFILL_3__1713_ gnd vdd FILL
XFILL_5__2629_ gnd vdd FILL
X_3262_ _3262_/D vdd _3289_/R _3307_/CLK _3262_/Q vdd gnd DFFSR
XFILL_8__2338_ gnd vdd FILL
XFILL_0__1935_ gnd vdd FILL
XFILL_0__1866_ gnd vdd FILL
XFILL_8__2269_ gnd vdd FILL
X_2213_ _2932_/B _2896_/B _2214_/C vdd gnd NOR2X1
X_3193_ _3193_/A _3193_/B _3196_/C vdd gnd NOR2X1
X_2144_ _2332_/B _2144_/B _2330_/B _2156_/A vdd gnd NAND3X1
XFILL_6__3023_ gnd vdd FILL
XFILL_0__3536_ gnd vdd FILL
XFILL_0__1797_ gnd vdd FILL
X_2075_ _2075_/A _2075_/B _2075_/C _2318_/C vdd gnd AOI21X1
XFILL_0__3467_ gnd vdd FILL
XFILL_1__2260_ gnd vdd FILL
XFILL_3__3176_ gnd vdd FILL
XFILL_0__3398_ gnd vdd FILL
XFILL_1__2191_ gnd vdd FILL
XFILL_0__2418_ gnd vdd FILL
XFILL_3__2127_ gnd vdd FILL
XFILL_0__2349_ gnd vdd FILL
XFILL_4__2940_ gnd vdd FILL
X_2977_ _3260_/Q _3264_/Q _2977_/C _2978_/B vdd gnd OAI21X1
XFILL_3__2058_ gnd vdd FILL
X_1928_ _3325_/Q _3092_/A _1931_/A vdd gnd NAND2X1
X_1859_ _2924_/A _2906_/B _1862_/B _1871_/A vdd gnd OAI21X1
XFILL_7__2580_ gnd vdd FILL
XFILL_6__2807_ gnd vdd FILL
XFILL_4__2871_ gnd vdd FILL
XFILL_6__2738_ gnd vdd FILL
XFILL_4__1822_ gnd vdd FILL
XFILL_4__1753_ gnd vdd FILL
X_3529_ _3555_/A _3555_/B _3529_/C _3531_/B vdd gnd OAI21X1
XFILL_1__1975_ gnd vdd FILL
XFILL_6__2669_ gnd vdd FILL
XFILL_7__3201_ gnd vdd FILL
XFILL_4__3423_ gnd vdd FILL
XFILL_7__3132_ gnd vdd FILL
XFILL_7__3063_ gnd vdd FILL
XFILL_7__2014_ gnd vdd FILL
XFILL_4__2305_ gnd vdd FILL
XFILL_4__2236_ gnd vdd FILL
XFILL_1__2527_ gnd vdd FILL
XFILL_1__2458_ gnd vdd FILL
XFILL_4__2167_ gnd vdd FILL
XFILL_7__2916_ gnd vdd FILL
XFILL_5__2980_ gnd vdd FILL
XFILL_1__2389_ gnd vdd FILL
XFILL_4__2098_ gnd vdd FILL
XFILL_5__1931_ gnd vdd FILL
XFILL_7__2847_ gnd vdd FILL
XFILL_5__1862_ gnd vdd FILL
XFILL_7__2778_ gnd vdd FILL
XFILL_5__3601_ gnd vdd FILL
XFILL_7__1729_ gnd vdd FILL
XFILL_5__1793_ gnd vdd FILL
XFILL_5__3532_ gnd vdd FILL
XFILL_2_BUFX2_insert8 gnd vdd FILL
XFILL_5__3463_ gnd vdd FILL
XFILL_2__2705_ gnd vdd FILL
XFILL_8__3172_ gnd vdd FILL
XFILL_5__3394_ gnd vdd FILL
XFILL_5__2414_ gnd vdd FILL
XFILL_0__1720_ gnd vdd FILL
XFILL_8__2123_ gnd vdd FILL
XFILL_5__2345_ gnd vdd FILL
XFILL_2__2636_ gnd vdd FILL
XFILL_8__2054_ gnd vdd FILL
XFILL_5__2276_ gnd vdd FILL
XFILL_2__2567_ gnd vdd FILL
XFILL_2__2498_ gnd vdd FILL
XFILL_6_BUFX2_insert11 gnd vdd FILL
XFILL_6_BUFX2_insert22 gnd vdd FILL
XFILL_3__3030_ gnd vdd FILL
XFILL_6_BUFX2_insert44 gnd vdd FILL
X_2900_ _2900_/A _2900_/B _2908_/A _2903_/B vdd gnd OAI21X1
XFILL_6_BUFX2_insert88 gnd vdd FILL
XFILL_6_BUFX2_insert66 gnd vdd FILL
XFILL_6_BUFX2_insert55 gnd vdd FILL
XFILL_6_BUFX2_insert77 gnd vdd FILL
XFILL_8__2956_ gnd vdd FILL
XFILL_0__2203_ gnd vdd FILL
X_2831_ _2870_/B _2835_/B _2832_/C vdd gnd NOR2X1
XFILL_2__3119_ gnd vdd FILL
XFILL_8__2887_ gnd vdd FILL
XFILL_8__1907_ gnd vdd FILL
XFILL_0__3183_ gnd vdd FILL
XFILL_6__1971_ gnd vdd FILL
XFILL_8__1838_ gnd vdd FILL
XFILL_0__2134_ gnd vdd FILL
X_2762_ _2762_/A _2762_/B _2762_/C _2766_/B vdd gnd NAND3X1
XFILL_0__2065_ gnd vdd FILL
X_1713_ _3236_/Q _1793_/B vdd gnd INVX1
XFILL_8__3508_ gnd vdd FILL
XFILL_8__1769_ gnd vdd FILL
X_2693_ _3247_/Q _2725_/D _2725_/C _2708_/B vdd gnd NAND3X1
XFILL_3__2814_ gnd vdd FILL
XFILL_6__2523_ gnd vdd FILL
XFILL_8__3439_ gnd vdd FILL
XFILL_3__2745_ gnd vdd FILL
XFILL_1__1760_ gnd vdd FILL
XFILL_0__2967_ gnd vdd FILL
X_3314_ _3314_/D vdd _3362_/R _3578_/CLK _3314_/Q vdd gnd DFFSR
XFILL_6__2454_ gnd vdd FILL
XFILL_0__1918_ gnd vdd FILL
XFILL_6__2385_ gnd vdd FILL
XFILL_3__2676_ gnd vdd FILL
X_3245_ _3245_/D vdd _3362_/R _3362_/CLK _3245_/Q vdd gnd DFFSR
XFILL_1__3430_ gnd vdd FILL
XFILL_0__2898_ gnd vdd FILL
XFILL_1__1691_ gnd vdd FILL
XFILL_0__1849_ gnd vdd FILL
X_3176_ _3176_/A _3176_/B _3176_/C _3197_/A vdd gnd NAND3X1
XFILL_4__3070_ gnd vdd FILL
X_2127_ _3147_/A _2446_/B _3197_/C _2129_/C vdd gnd OAI21X1
XFILL_4__2021_ gnd vdd FILL
XFILL_0__3519_ gnd vdd FILL
XFILL_6__3006_ gnd vdd FILL
XFILL_1__2312_ gnd vdd FILL
X_2058_ _3160_/A _2058_/B _3166_/A _2060_/A vdd gnd OAI21X1
XFILL_1__2243_ gnd vdd FILL
XFILL_3__3228_ gnd vdd FILL
XFILL_3__3159_ gnd vdd FILL
XFILL_1__2174_ gnd vdd FILL
XFILL_7__2701_ gnd vdd FILL
XFILL_4__2923_ gnd vdd FILL
XFILL_7__2632_ gnd vdd FILL
XFILL_4__2854_ gnd vdd FILL
XFILL_4__1805_ gnd vdd FILL
XFILL_7__2563_ gnd vdd FILL
XFILL_4__2785_ gnd vdd FILL
XFILL_7__2494_ gnd vdd FILL
XFILL_4__1736_ gnd vdd FILL
XFILL_1__1958_ gnd vdd FILL
XFILL_2__3470_ gnd vdd FILL
XFILL_7__3115_ gnd vdd FILL
XFILL_4__3406_ gnd vdd FILL
XFILL_1__1889_ gnd vdd FILL
XFILL_2__2421_ gnd vdd FILL
XFILL_5__2130_ gnd vdd FILL
XFILL_1__3559_ gnd vdd FILL
XFILL_7__3046_ gnd vdd FILL
XFILL_2__2352_ gnd vdd FILL
XFILL_5__2061_ gnd vdd FILL
XFILL_8__2810_ gnd vdd FILL
XFILL_2__2283_ gnd vdd FILL
XFILL_4__2219_ gnd vdd FILL
XFILL_4__3199_ gnd vdd FILL
XFILL_8__2741_ gnd vdd FILL
XFILL_5__2963_ gnd vdd FILL
XFILL_8__2672_ gnd vdd FILL
XFILL_5__2894_ gnd vdd FILL
XFILL_5__1914_ gnd vdd FILL
XFILL_5__1845_ gnd vdd FILL
XFILL_5__1776_ gnd vdd FILL
XFILL_5__3515_ gnd vdd FILL
XFILL_2__1998_ gnd vdd FILL
XFILL_0__2821_ gnd vdd FILL
XFILL_8__3224_ gnd vdd FILL
XFILL_5__3446_ gnd vdd FILL
XFILL_3__2530_ gnd vdd FILL
XFILL_0__2752_ gnd vdd FILL
XFILL_6__2170_ gnd vdd FILL
XFILL_0__1703_ gnd vdd FILL
XFILL_3__2461_ gnd vdd FILL
XFILL_8__3155_ gnd vdd FILL
XFILL_5__3377_ gnd vdd FILL
XFILL_8__3086_ gnd vdd FILL
XFILL_3__2392_ gnd vdd FILL
X_3030_ _3165_/A _3063_/B _3030_/C _3031_/C vdd gnd OAI21X1
XFILL_0__2683_ gnd vdd FILL
XFILL_2__2619_ gnd vdd FILL
XFILL_8__2106_ gnd vdd FILL
XFILL_8__2037_ gnd vdd FILL
XFILL_5__2328_ gnd vdd FILL
XFILL_2__3599_ gnd vdd FILL
XFILL_5__2259_ gnd vdd FILL
XFILL184650x101550 gnd vdd FILL
XFILL_3__3013_ gnd vdd FILL
XFILL_8__2939_ gnd vdd FILL
X_2814_ _2814_/A _3006_/B _3267_/Q _2815_/C vdd gnd OAI21X1
XFILL_6__1954_ gnd vdd FILL
XFILL_0__3166_ gnd vdd FILL
XFILL_0__2117_ gnd vdd FILL
XFILL_0__3097_ gnd vdd FILL
XFILL_6__1885_ gnd vdd FILL
X_2745_ _3252_/Q _2778_/A _2754_/C vdd gnd NAND2X1
XFILL_1__2930_ gnd vdd FILL
X_2676_ _3197_/C _2676_/B _2676_/C _3246_/D vdd gnd OAI21X1
XFILL_0__2048_ gnd vdd FILL
XFILL_2_BUFX2_insert20 gnd vdd FILL
XFILL_1__2861_ gnd vdd FILL
XFILL_6__3555_ gnd vdd FILL
XFILL_6__3486_ gnd vdd FILL
XFILL_6__2506_ gnd vdd FILL
XFILL_2_BUFX2_insert42 gnd vdd FILL
XFILL_2_BUFX2_insert53 gnd vdd FILL
XFILL_4__2570_ gnd vdd FILL
XFILL_1__1812_ gnd vdd FILL
XFILL_2_BUFX2_insert97 gnd vdd FILL
XFILL_2_BUFX2_insert64 gnd vdd FILL
XFILL_1__2792_ gnd vdd FILL
XFILL_2_BUFX2_insert75 gnd vdd FILL
XFILL_3__2728_ gnd vdd FILL
XFILL_2_BUFX2_insert86 gnd vdd FILL
XFILL_6__2437_ gnd vdd FILL
XFILL_1__1743_ gnd vdd FILL
XFILL_3__2659_ gnd vdd FILL
XFILL_6__2368_ gnd vdd FILL
X_3228_ _3228_/A _3228_/B _3228_/C _3361_/D vdd gnd OAI21X1
XFILL_1__3413_ gnd vdd FILL
XFILL_6__2299_ gnd vdd FILL
X_3159_ _3159_/A _3159_/B _3169_/C vdd gnd NOR2X1
XFILL_4__3122_ gnd vdd FILL
XFILL_4__3053_ gnd vdd FILL
XFILL_4__2004_ gnd vdd FILL
XFILL_7__1994_ gnd vdd FILL
XFILL_1__2226_ gnd vdd FILL
XFILL_1__2157_ gnd vdd FILL
XFILL_4__2906_ gnd vdd FILL
XFILL_2__2970_ gnd vdd FILL
XFILL_1__2088_ gnd vdd FILL
XFILL_2__1921_ gnd vdd FILL
XFILL_7__3595_ gnd vdd FILL
XFILL_7__2615_ gnd vdd FILL
XFILL_4__2837_ gnd vdd FILL
XFILL_7__2546_ gnd vdd FILL
XFILL_2__1852_ gnd vdd FILL
XFILL_4__2768_ gnd vdd FILL
XFILL_4__1719_ gnd vdd FILL
XFILL_2__1783_ gnd vdd FILL
XFILL_7__2477_ gnd vdd FILL
XFILL_0_CLKBUF1_insert37 gnd vdd FILL
XFILL_2__3522_ gnd vdd FILL
XFILL_5__3231_ gnd vdd FILL
XFILL_4__2699_ gnd vdd FILL
XFILL_2__3453_ gnd vdd FILL
XFILL_2__2404_ gnd vdd FILL
XFILL_5__3162_ gnd vdd FILL
XFILL_7__3029_ gnd vdd FILL
XFILL_5__3093_ gnd vdd FILL
XFILL_2__3384_ gnd vdd FILL
XFILL_5__2113_ gnd vdd FILL
XFILL_5__2044_ gnd vdd FILL
XFILL_2__2335_ gnd vdd FILL
XFILL_2__2266_ gnd vdd FILL
XFILL_2__2197_ gnd vdd FILL
XFILL_0__3020_ gnd vdd FILL
XFILL_8__2724_ gnd vdd FILL
XFILL_5__2946_ gnd vdd FILL
XFILL_3__1961_ gnd vdd FILL
XFILL_8__2655_ gnd vdd FILL
XFILL_5__2877_ gnd vdd FILL
X_2530_ _2711_/B _2574_/B _2530_/C _3594_/A vdd gnd OAI21X1
XFILL_8__2586_ gnd vdd FILL
X_2461_ _2612_/B _2574_/B _2461_/C _2462_/C vdd gnd OAI21X1
XFILL_3__1892_ gnd vdd FILL
XFILL_5__1828_ gnd vdd FILL
XFILL_5__1759_ gnd vdd FILL
XFILL_3__3562_ gnd vdd FILL
X_2392_ _2392_/A _2392_/B _2392_/C _3596_/A vdd gnd NAND3X1
XFILL_0__2804_ gnd vdd FILL
XFILL184650x113250 gnd vdd FILL
XFILL_8__3207_ gnd vdd FILL
XFILL_3__2513_ gnd vdd FILL
XFILL_3__3493_ gnd vdd FILL
XFILL_8__3138_ gnd vdd FILL
XFILL_5__3429_ gnd vdd FILL
XFILL184350x121050 gnd vdd FILL
XFILL_6__2222_ gnd vdd FILL
XFILL_0__2735_ gnd vdd FILL
X_3013_ _3260_/Q _3570_/Q _3013_/C _3015_/B vdd gnd AOI21X1
XFILL_6__2153_ gnd vdd FILL
XFILL_0__2666_ gnd vdd FILL
XFILL_3__2444_ gnd vdd FILL
XFILL_6__2084_ gnd vdd FILL
XFILL_8__3069_ gnd vdd FILL
XFILL_3__2375_ gnd vdd FILL
XFILL_0__2597_ gnd vdd FILL
XFILL_1__3060_ gnd vdd FILL
XFILL_1__2011_ gnd vdd FILL
XFILL_0__3218_ gnd vdd FILL
XFILL_6__2986_ gnd vdd FILL
XFILL_6__1937_ gnd vdd FILL
XFILL_0__3149_ gnd vdd FILL
XFILL_6__1868_ gnd vdd FILL
X_2728_ _2728_/A _2728_/B _2728_/C _2729_/C vdd gnd NAND3X1
XFILL_1__2913_ gnd vdd FILL
XFILL_7__3380_ gnd vdd FILL
XFILL_7__2400_ gnd vdd FILL
XFILL_6__3538_ gnd vdd FILL
XFILL_7__2331_ gnd vdd FILL
XFILL_6__1799_ gnd vdd FILL
XFILL_4__2622_ gnd vdd FILL
X_2659_ _2675_/A _2659_/B _2659_/C _2659_/D _3244_/D vdd gnd OAI22X1
XFILL_1__2844_ gnd vdd FILL
XFILL_4__2553_ gnd vdd FILL
XFILL_6__3469_ gnd vdd FILL
XFILL_7__2262_ gnd vdd FILL
XFILL_1__2775_ gnd vdd FILL
XFILL_7__2193_ gnd vdd FILL
XFILL_4__2484_ gnd vdd FILL
XFILL_1__1726_ gnd vdd FILL
XFILL_4__3105_ gnd vdd FILL
XFILL_2__2120_ gnd vdd FILL
XFILL_4__3036_ gnd vdd FILL
XFILL_2__2051_ gnd vdd FILL
XFILL_7__1977_ gnd vdd FILL
XFILL_5__2800_ gnd vdd FILL
XFILL_1__2209_ gnd vdd FILL
XFILL_1__3189_ gnd vdd FILL
XFILL_5__2731_ gnd vdd FILL
XFILL_8__2440_ gnd vdd FILL
XFILL_2__2953_ gnd vdd FILL
XFILL_5__2662_ gnd vdd FILL
XFILL_2__2884_ gnd vdd FILL
XFILL_8__2371_ gnd vdd FILL
XFILL_7_BUFX2_insert3 gnd vdd FILL
XFILL_2__1904_ gnd vdd FILL
XFILL_7__2529_ gnd vdd FILL
XFILL_5__2593_ gnd vdd FILL
XFILL_2__1835_ gnd vdd FILL
XFILL_2__3505_ gnd vdd FILL
XFILL_2__1766_ gnd vdd FILL
XFILL_2__1697_ gnd vdd FILL
XFILL_5__3214_ gnd vdd FILL
XFILL_0__2520_ gnd vdd FILL
XFILL_2__3436_ gnd vdd FILL
XFILL_5__3145_ gnd vdd FILL
XFILL_3__2160_ gnd vdd FILL
XFILL_2__3367_ gnd vdd FILL
XFILL_0__2451_ gnd vdd FILL
XFILL_5__3076_ gnd vdd FILL
XFILL_2__2318_ gnd vdd FILL
XFILL_0__2382_ gnd vdd FILL
XFILL_5__2027_ gnd vdd FILL
XFILL_3__2091_ gnd vdd FILL
XFILL_6__2840_ gnd vdd FILL
XFILL_2__2249_ gnd vdd FILL
X_1961_ _3361_/Q _2691_/A _2746_/C vdd gnd NAND2X1
XFILL_0__3003_ gnd vdd FILL
X_1892_ _2108_/A _3145_/B _2872_/B vdd gnd NOR2X1
XFILL_8__2707_ gnd vdd FILL
XFILL_6__2771_ gnd vdd FILL
XFILL_5__2929_ gnd vdd FILL
X_3562_ _3566_/A _3562_/B _3563_/C vdd gnd NAND2X1
XFILL_3__2993_ gnd vdd FILL
XFILL_6__1722_ gnd vdd FILL
XFILL_8__2638_ gnd vdd FILL
X_2513_ _2513_/A _2514_/C vdd gnd INVX1
XFILL_3__1944_ gnd vdd FILL
XFILL_3__1875_ gnd vdd FILL
X_3493_ _3493_/A _3493_/B _3497_/A _3494_/B vdd gnd OAI21X1
XFILL_8__2569_ gnd vdd FILL
X_2444_ _2444_/A _2444_/B _2444_/C _2569_/B vdd gnd NAND3X1
XFILL_9__3032_ gnd vdd FILL
X_2375_ _2375_/A _2375_/B _3283_/Q _2376_/A vdd gnd OAI21X1
XFILL_3__3545_ gnd vdd FILL
XFILL_1__2560_ gnd vdd FILL
XFILL_3__3476_ gnd vdd FILL
XFILL_6__2205_ gnd vdd FILL
XFILL_3__2427_ gnd vdd FILL
XFILL_1__2491_ gnd vdd FILL
XFILL_0__2718_ gnd vdd FILL
XFILL_6__3185_ gnd vdd FILL
XFILL_6__2136_ gnd vdd FILL
XFILL_0__2649_ gnd vdd FILL
XFILL_3__2358_ gnd vdd FILL
XFILL_6__2067_ gnd vdd FILL
XFILL_1__3112_ gnd vdd FILL
XFILL_7__1900_ gnd vdd FILL
XFILL_3__2289_ gnd vdd FILL
XFILL_7__2880_ gnd vdd FILL
XFILL_1__3043_ gnd vdd FILL
XFILL_7__1831_ gnd vdd FILL
XFILL_5_BUFX2_insert90 gnd vdd FILL
XFILL_6__2969_ gnd vdd FILL
XFILL_7__1762_ gnd vdd FILL
XFILL_7__3501_ gnd vdd FILL
XFILL_4__1984_ gnd vdd FILL
XFILL_7__3432_ gnd vdd FILL
XFILL_7__1693_ gnd vdd FILL
XFILL_4__2605_ gnd vdd FILL
XFILL_1__2827_ gnd vdd FILL
XFILL_7__2314_ gnd vdd FILL
XFILL_4__3585_ gnd vdd FILL
XFILL_7__2245_ gnd vdd FILL
XFILL_4__2536_ gnd vdd FILL
XFILL_4__2467_ gnd vdd FILL
XFILL_1__2758_ gnd vdd FILL
XFILL_1__1709_ gnd vdd FILL
XFILL_7__2176_ gnd vdd FILL
XFILL_1__2689_ gnd vdd FILL
XFILL_4__2398_ gnd vdd FILL
XFILL_2__3221_ gnd vdd FILL
XFILL_8__1940_ gnd vdd FILL
XFILL_2__3152_ gnd vdd FILL
XFILL_8__1871_ gnd vdd FILL
XFILL_4__3019_ gnd vdd FILL
XFILL_2__3083_ gnd vdd FILL
XFILL_2__2103_ gnd vdd FILL
XFILL_2__2034_ gnd vdd FILL
XFILL_8__3541_ gnd vdd FILL
XFILL_3_BUFX2_insert19 gnd vdd FILL
XFILL_8__3472_ gnd vdd FILL
XFILL_5__2714_ gnd vdd FILL
XFILL_2__2936_ gnd vdd FILL
XFILL_8__2423_ gnd vdd FILL
XFILL_8__2354_ gnd vdd FILL
XFILL_0__1951_ gnd vdd FILL
XFILL_5__2645_ gnd vdd FILL
XFILL_2__2867_ gnd vdd FILL
XFILL_5__2576_ gnd vdd FILL
XFILL_0__1882_ gnd vdd FILL
XFILL_2__2798_ gnd vdd FILL
XFILL_8__2285_ gnd vdd FILL
XFILL_2__1818_ gnd vdd FILL
X_2160_ _2270_/A _2312_/A vdd gnd INVX1
XFILL_2__1749_ gnd vdd FILL
XFILL_0__3552_ gnd vdd FILL
X_2091_ _2432_/A _2091_/B _3183_/C vdd gnd NAND2X1
XFILL_0__3483_ gnd vdd FILL
XFILL_2__3419_ gnd vdd FILL
XFILL_0__2503_ gnd vdd FILL
XFILL_3__2212_ gnd vdd FILL
XFILL_5__3128_ gnd vdd FILL
XFILL_3__3192_ gnd vdd FILL
XFILL_0__2434_ gnd vdd FILL
XFILL_5__3059_ gnd vdd FILL
XFILL_3__2143_ gnd vdd FILL
X_2993_ _2993_/A _2993_/B _2993_/C _2996_/B vdd gnd OAI21X1
XFILL_3__2074_ gnd vdd FILL
XFILL_0__2365_ gnd vdd FILL
XFILL_0__2296_ gnd vdd FILL
X_1944_ _2948_/A _1984_/B _2728_/B _1945_/C vdd gnd OAI21X1
XFILL_6__2823_ gnd vdd FILL
XFILL_9__2532_ gnd vdd FILL
X_1875_ _1875_/A _3285_/Q _1879_/B vdd gnd OR2X2
XFILL_6__2754_ gnd vdd FILL
XFILL_3__2976_ gnd vdd FILL
XFILL_6__1705_ gnd vdd FILL
X_3545_ _3545_/A _3545_/B _3566_/A _3546_/B vdd gnd OAI21X1
XFILL_3__1927_ gnd vdd FILL
XFILL_1__1991_ gnd vdd FILL
XFILL_6__2685_ gnd vdd FILL
X_3476_ _3476_/A _3494_/A _3497_/A _3526_/A vdd gnd OAI21X1
X_2427_ _3577_/Q _2427_/B _2427_/C _2428_/B vdd gnd AOI21X1
XFILL_3__1858_ gnd vdd FILL
XFILL_4__3370_ gnd vdd FILL
XFILL_3__1789_ gnd vdd FILL
XFILL_3__3528_ gnd vdd FILL
X_2358_ _2968_/A _2444_/B _2579_/B _2361_/C vdd gnd NAND3X1
XFILL_4__2321_ gnd vdd FILL
XFILL_1__3592_ gnd vdd FILL
XFILL_1__2612_ gnd vdd FILL
XFILL_7__2030_ gnd vdd FILL
XFILL_1__2543_ gnd vdd FILL
X_2289_ _2438_/A _2289_/B _2293_/A _2290_/A vdd gnd MUX2X1
XFILL_3__3459_ gnd vdd FILL
XFILL_4__2252_ gnd vdd FILL
XFILL_6__3168_ gnd vdd FILL
XFILL_4__2183_ gnd vdd FILL
XFILL_6__2119_ gnd vdd FILL
XFILL_1__2474_ gnd vdd FILL
XFILL_6__3099_ gnd vdd FILL
XFILL_7__2932_ gnd vdd FILL
XFILL_7__2863_ gnd vdd FILL
XFILL_1__3026_ gnd vdd FILL
XFILL_7__1814_ gnd vdd FILL
XFILL_7__2794_ gnd vdd FILL
XFILL_7__1745_ gnd vdd FILL
XFILL_5_CLKBUF1_insert37 gnd vdd FILL
XFILL_4__1967_ gnd vdd FILL
XFILL_7__3415_ gnd vdd FILL
XFILL_4__1898_ gnd vdd FILL
XFILL_2__2721_ gnd vdd FILL
XFILL_5__2430_ gnd vdd FILL
XFILL_5__2361_ gnd vdd FILL
XFILL_2__2652_ gnd vdd FILL
XFILL_8__2070_ gnd vdd FILL
XFILL_2__2583_ gnd vdd FILL
XFILL_4__2519_ gnd vdd FILL
XFILL_4__3499_ gnd vdd FILL
XFILL_7__2228_ gnd vdd FILL
XFILL_3_CLKBUF1_insert30 gnd vdd FILL
XFILL_5__2292_ gnd vdd FILL
XFILL_7__2159_ gnd vdd FILL
XFILL_8__2972_ gnd vdd FILL
XFILL_2__3204_ gnd vdd FILL
XFILL_2__3135_ gnd vdd FILL
XFILL_8__1923_ gnd vdd FILL
XFILL_8__1854_ gnd vdd FILL
XFILL_0__2150_ gnd vdd FILL
XFILL_0__2081_ gnd vdd FILL
XFILL_2__3066_ gnd vdd FILL
XFILL_2__2017_ gnd vdd FILL
XFILL_8__1785_ gnd vdd FILL
XFILL_3__2830_ gnd vdd FILL
XFILL_8__3524_ gnd vdd FILL
XFILL_8__3455_ gnd vdd FILL
X_3330_ _3330_/D vdd _3347_/R _3576_/CLK _3330_/Q vdd gnd DFFSR
XFILL_6__2470_ gnd vdd FILL
XFILL_3__2761_ gnd vdd FILL
XFILL_8__2406_ gnd vdd FILL
XFILL_2__2919_ gnd vdd FILL
XFILL_8__3386_ gnd vdd FILL
XFILL_0__2983_ gnd vdd FILL
XFILL_3__1712_ gnd vdd FILL
XFILL_3__2692_ gnd vdd FILL
XFILL_5__2628_ gnd vdd FILL
X_3261_ _3261_/D vdd _3313_/R _3313_/CLK _3261_/Q vdd gnd DFFSR
XFILL_8__2337_ gnd vdd FILL
XFILL_0__1934_ gnd vdd FILL
XFILL_0__1865_ gnd vdd FILL
XFILL_8__2268_ gnd vdd FILL
X_2212_ _2212_/A _3183_/B _3177_/A vdd gnd NOR2X1
XFILL_5__2559_ gnd vdd FILL
X_3192_ _3192_/A _3192_/B _3192_/C _3193_/B vdd gnd NAND3X1
X_2143_ _2342_/A _3171_/B _2143_/C _2330_/B vdd gnd OAI21X1
XFILL_0__3535_ gnd vdd FILL
XFILL_6__3022_ gnd vdd FILL
XFILL_0__1796_ gnd vdd FILL
XFILL_8__2199_ gnd vdd FILL
X_2074_ _2074_/A _2074_/B _2075_/C vdd gnd OR2X2
XFILL_0__3466_ gnd vdd FILL
XFILL_3__3175_ gnd vdd FILL
XFILL_0__3397_ gnd vdd FILL
XFILL_1__2190_ gnd vdd FILL
XFILL_0__2417_ gnd vdd FILL
XFILL_3__2126_ gnd vdd FILL
XFILL_0__2348_ gnd vdd FILL
X_2976_ _3260_/Q _3573_/Q _2977_/C vdd gnd NAND2X1
XFILL_3__2057_ gnd vdd FILL
XFILL_4__2870_ gnd vdd FILL
XFILL_6__2806_ gnd vdd FILL
X_1927_ _1986_/A _1927_/B _1927_/C _3460_/B vdd gnd OAI21X1
XFILL_0__2279_ gnd vdd FILL
XFILL_4__1821_ gnd vdd FILL
X_1858_ _1891_/A _1858_/B _2602_/A _1858_/Y vdd gnd NAND3X1
XFILL_6__2737_ gnd vdd FILL
XFILL_3__2959_ gnd vdd FILL
XFILL_4__1752_ gnd vdd FILL
X_1789_ _1846_/B _3161_/B vdd gnd INVX1
XFILL_6__2668_ gnd vdd FILL
X_3528_ _3528_/A _3528_/B _3528_/C _3555_/B vdd gnd AOI21X1
XFILL_1__1974_ gnd vdd FILL
XFILL_7__3200_ gnd vdd FILL
X_3459_ _3459_/A _3459_/B _3461_/B vdd gnd NAND2X1
XFILL_4__3422_ gnd vdd FILL
XFILL_6__2599_ gnd vdd FILL
XFILL_7__3131_ gnd vdd FILL
XFILL_7__3062_ gnd vdd FILL
XFILL_7__2013_ gnd vdd FILL
XFILL_4__2304_ gnd vdd FILL
XFILL_4__2235_ gnd vdd FILL
XFILL_1__2526_ gnd vdd FILL
XFILL_1__2457_ gnd vdd FILL
XFILL_4__2166_ gnd vdd FILL
XFILL_7__2915_ gnd vdd FILL
XFILL_1__2388_ gnd vdd FILL
XFILL_4__2097_ gnd vdd FILL
XFILL_5__1930_ gnd vdd FILL
XFILL_7__2846_ gnd vdd FILL
XFILL_1__3009_ gnd vdd FILL
XFILL_5__3600_ gnd vdd FILL
XFILL_5__1861_ gnd vdd FILL
XFILL_7__2777_ gnd vdd FILL
XFILL_4__2999_ gnd vdd FILL
XFILL_5__1792_ gnd vdd FILL
XFILL_7__1728_ gnd vdd FILL
XFILL_5__3531_ gnd vdd FILL
XFILL182850x7950 gnd vdd FILL
XFILL_5__3462_ gnd vdd FILL
XFILL_2_BUFX2_insert9 gnd vdd FILL
XFILL_8__3171_ gnd vdd FILL
XFILL_2__2704_ gnd vdd FILL
XFILL_5__2413_ gnd vdd FILL
XFILL_5__3393_ gnd vdd FILL
XFILL_8__2122_ gnd vdd FILL
XFILL_2__2635_ gnd vdd FILL
XFILL_5__2344_ gnd vdd FILL
XFILL_8__2053_ gnd vdd FILL
XFILL_5__2275_ gnd vdd FILL
XFILL_2__2566_ gnd vdd FILL
XFILL_2__2497_ gnd vdd FILL
XFILL_6_BUFX2_insert12 gnd vdd FILL
XFILL_6_BUFX2_insert23 gnd vdd FILL
XFILL_6_BUFX2_insert45 gnd vdd FILL
XFILL_6_BUFX2_insert56 gnd vdd FILL
XFILL_6_BUFX2_insert78 gnd vdd FILL
XFILL_6_BUFX2_insert67 gnd vdd FILL
X_2830_ _2887_/B _2911_/A _2870_/B vdd gnd NOR2X1
XFILL_8__2955_ gnd vdd FILL
XFILL_0__2202_ gnd vdd FILL
XFILL_0__3182_ gnd vdd FILL
XFILL_6__1970_ gnd vdd FILL
XFILL_6_BUFX2_insert89 gnd vdd FILL
XFILL_2__3118_ gnd vdd FILL
XFILL182550x148350 gnd vdd FILL
XFILL_8__2886_ gnd vdd FILL
XFILL_0__2133_ gnd vdd FILL
XFILL_8__1906_ gnd vdd FILL
XFILL_2__3049_ gnd vdd FILL
X_2761_ _3576_/Q _2770_/B _2770_/C _3362_/Q _2762_/B vdd gnd AOI22X1
XFILL_8__1837_ gnd vdd FILL
XFILL_8__1768_ gnd vdd FILL
XFILL_0__2064_ gnd vdd FILL
X_1712_ _3568_/Q _1751_/A vdd gnd INVX1
X_2692_ _2692_/A _2725_/D vdd gnd INVX1
XFILL_8__3507_ gnd vdd FILL
XFILL_3__2813_ gnd vdd FILL
XFILL_8__1699_ gnd vdd FILL
XFILL_6__2522_ gnd vdd FILL
XFILL_8__3438_ gnd vdd FILL
XFILL_3__2744_ gnd vdd FILL
X_3313_ _3313_/D vdd _3313_/R _3313_/CLK _3313_/Q vdd gnd DFFSR
XFILL_0__2966_ gnd vdd FILL
XFILL_8__3369_ gnd vdd FILL
XFILL_6__2453_ gnd vdd FILL
XFILL_0__1917_ gnd vdd FILL
XFILL_6__2384_ gnd vdd FILL
XFILL_3__2675_ gnd vdd FILL
X_3244_ _3244_/D vdd _3362_/R _3355_/CLK _3244_/Q vdd gnd DFFSR
XFILL_0__2897_ gnd vdd FILL
XFILL_1__1690_ gnd vdd FILL
XFILL_0__1848_ gnd vdd FILL
X_3175_ _3175_/A _3175_/B _3176_/C vdd gnd AND2X2
XFILL_6__3005_ gnd vdd FILL
X_2126_ _2278_/A _3017_/A _2126_/C _2348_/B vdd gnd OAI21X1
XFILL_0__1779_ gnd vdd FILL
XFILL_4__2020_ gnd vdd FILL
XFILL_0__3518_ gnd vdd FILL
XFILL_1__2311_ gnd vdd FILL
XFILL_3__3227_ gnd vdd FILL
X_2057_ _2057_/A _2442_/A _3166_/A vdd gnd NOR2X1
XFILL_0__3449_ gnd vdd FILL
XFILL_1__2242_ gnd vdd FILL
XFILL_3__3158_ gnd vdd FILL
XFILL_3__3089_ gnd vdd FILL
XFILL_1__2173_ gnd vdd FILL
XFILL_7__2700_ gnd vdd FILL
XFILL_3__2109_ gnd vdd FILL
XFILL_4__2922_ gnd vdd FILL
X_2959_ _2999_/B _2981_/A vdd gnd INVX1
XFILL_7__2631_ gnd vdd FILL
XFILL_4__2853_ gnd vdd FILL
XFILL_7__2562_ gnd vdd FILL
XFILL_4__2784_ gnd vdd FILL
XFILL_4__1804_ gnd vdd FILL
XFILL_7__2493_ gnd vdd FILL
XFILL_4__1735_ gnd vdd FILL
XFILL_9__2429_ gnd vdd FILL
XFILL_1__1957_ gnd vdd FILL
XFILL_7__3114_ gnd vdd FILL
XFILL_4__3405_ gnd vdd FILL
XFILL_1__1888_ gnd vdd FILL
XFILL_2__2420_ gnd vdd FILL
XFILL_1__3558_ gnd vdd FILL
XFILL_7__3045_ gnd vdd FILL
XFILL_2__2351_ gnd vdd FILL
XFILL184350x85950 gnd vdd FILL
XFILL_1__2509_ gnd vdd FILL
XFILL_5__2060_ gnd vdd FILL
XFILL_1__3489_ gnd vdd FILL
XFILL_2__2282_ gnd vdd FILL
XFILL_4__2218_ gnd vdd FILL
XFILL_4__3198_ gnd vdd FILL
XFILL_4__2149_ gnd vdd FILL
XFILL_8__2740_ gnd vdd FILL
XFILL_5__2962_ gnd vdd FILL
XFILL_8__2671_ gnd vdd FILL
XFILL_7__2829_ gnd vdd FILL
XFILL_5__2893_ gnd vdd FILL
XFILL_5__1913_ gnd vdd FILL
XFILL_5__1844_ gnd vdd FILL
XFILL_5__3514_ gnd vdd FILL
XFILL_5__1775_ gnd vdd FILL
XFILL_0__2820_ gnd vdd FILL
XFILL_8__3223_ gnd vdd FILL
XFILL_2__1997_ gnd vdd FILL
XFILL_5__3445_ gnd vdd FILL
XFILL_0__2751_ gnd vdd FILL
XFILL_8__3154_ gnd vdd FILL
XFILL_5__3376_ gnd vdd FILL
XFILL_0__1702_ gnd vdd FILL
XFILL_3__2460_ gnd vdd FILL
XFILL_8__2105_ gnd vdd FILL
XFILL_5__2327_ gnd vdd FILL
XFILL_8__3085_ gnd vdd FILL
XFILL_2__3598_ gnd vdd FILL
XFILL_3__2391_ gnd vdd FILL
XFILL_0__2682_ gnd vdd FILL
XFILL_2__2618_ gnd vdd FILL
XFILL_8__2036_ gnd vdd FILL
XFILL_2__2549_ gnd vdd FILL
XFILL_5__2258_ gnd vdd FILL
XFILL_5__2189_ gnd vdd FILL
XFILL_3__3012_ gnd vdd FILL
XFILL_8__2938_ gnd vdd FILL
X_2813_ _2980_/A _2898_/B _2813_/C _2815_/A _3266_/D vdd gnd OAI22X1
XFILL_6__1953_ gnd vdd FILL
XFILL_0__3165_ gnd vdd FILL
XFILL_8__2869_ gnd vdd FILL
XFILL_0__3096_ gnd vdd FILL
XFILL_0__2116_ gnd vdd FILL
XFILL_6__1884_ gnd vdd FILL
X_2744_ _3197_/C _2744_/B _2744_/C _3251_/D vdd gnd OAI21X1
XFILL_0__2047_ gnd vdd FILL
X_2675_ _2675_/A _2733_/B _2675_/C _2676_/C vdd gnd NAND3X1
XFILL_1__2860_ gnd vdd FILL
XFILL_6__3554_ gnd vdd FILL
XFILL_2_BUFX2_insert10 gnd vdd FILL
XFILL_6__3485_ gnd vdd FILL
XFILL_2_BUFX2_insert21 gnd vdd FILL
XFILL_6__2505_ gnd vdd FILL
XFILL_2_BUFX2_insert43 gnd vdd FILL
XFILL_2_BUFX2_insert54 gnd vdd FILL
XFILL_1__1811_ gnd vdd FILL
XFILL_1__2791_ gnd vdd FILL
XFILL_2_BUFX2_insert87 gnd vdd FILL
XFILL_2_BUFX2_insert65 gnd vdd FILL
XFILL_9__3194_ gnd vdd FILL
XFILL_3__2727_ gnd vdd FILL
XFILL_2_BUFX2_insert76 gnd vdd FILL
XFILL_6__2436_ gnd vdd FILL
XFILL_0__2949_ gnd vdd FILL
XFILL_1__1742_ gnd vdd FILL
XFILL_3__2658_ gnd vdd FILL
XFILL_6__2367_ gnd vdd FILL
X_3227_ _3584_/A _3227_/B _3228_/C vdd gnd NAND2X1
XFILL_4__3121_ gnd vdd FILL
XFILL_1__3412_ gnd vdd FILL
XFILL_6__2298_ gnd vdd FILL
XFILL_3__2589_ gnd vdd FILL
X_3158_ _3158_/A _3158_/B _3158_/C _3159_/B vdd gnd NAND3X1
X_2109_ _2221_/A _3182_/B _2294_/A _2110_/C vdd gnd OAI21X1
X_3089_ _3322_/Q _3090_/A _3090_/C vdd gnd NAND2X1
XFILL_4__3052_ gnd vdd FILL
XFILL_4__2003_ gnd vdd FILL
XFILL_7__1993_ gnd vdd FILL
XFILL_1__2225_ gnd vdd FILL
XFILL_1__2156_ gnd vdd FILL
XFILL_4__2905_ gnd vdd FILL
XFILL_1__2087_ gnd vdd FILL
XFILL_7__2614_ gnd vdd FILL
XFILL_4__2836_ gnd vdd FILL
XFILL_2__1920_ gnd vdd FILL
XFILL184650x62550 gnd vdd FILL
XFILL_7__3594_ gnd vdd FILL
XFILL_8_CLKBUF1_insert30 gnd vdd FILL
XFILL_2__1851_ gnd vdd FILL
XFILL_7__2545_ gnd vdd FILL
XFILL_7__2476_ gnd vdd FILL
XFILL_4__2767_ gnd vdd FILL
XFILL_1__2989_ gnd vdd FILL
XFILL_4__1718_ gnd vdd FILL
XFILL_4__2698_ gnd vdd FILL
XFILL_2__1782_ gnd vdd FILL
XFILL_2__3521_ gnd vdd FILL
XFILL_5__3230_ gnd vdd FILL
XFILL_2__3452_ gnd vdd FILL
XFILL_0_CLKBUF1_insert38 gnd vdd FILL
XFILL184350x97650 gnd vdd FILL
XFILL_2__2403_ gnd vdd FILL
XFILL_5__3161_ gnd vdd FILL
XFILL_5__2112_ gnd vdd FILL
XFILL_7__3028_ gnd vdd FILL
XFILL_5__3092_ gnd vdd FILL
XFILL_2__3383_ gnd vdd FILL
XFILL_5__2043_ gnd vdd FILL
XFILL_2__2334_ gnd vdd FILL
XFILL_2__2265_ gnd vdd FILL
XFILL_2__2196_ gnd vdd FILL
XFILL_8__2723_ gnd vdd FILL
XFILL_5__2945_ gnd vdd FILL
XFILL_3__1960_ gnd vdd FILL
XFILL_8__2654_ gnd vdd FILL
XFILL_5__2876_ gnd vdd FILL
XFILL_8__2585_ gnd vdd FILL
XFILL_5__1827_ gnd vdd FILL
X_2460_ _2460_/A _2460_/B _2461_/C vdd gnd AND2X2
XFILL_3__1891_ gnd vdd FILL
XFILL_5__1758_ gnd vdd FILL
XFILL_0__2803_ gnd vdd FILL
XFILL_3__3561_ gnd vdd FILL
X_2391_ _3571_/Q _2427_/B _2391_/C _2392_/B vdd gnd AOI21X1
XFILL184650x4050 gnd vdd FILL
XFILL_3__3492_ gnd vdd FILL
XFILL_5__3428_ gnd vdd FILL
XFILL_5__1689_ gnd vdd FILL
XFILL_8__3206_ gnd vdd FILL
XFILL_6__2221_ gnd vdd FILL
XFILL_3__2512_ gnd vdd FILL
XFILL_8__3137_ gnd vdd FILL
XFILL_0__2734_ gnd vdd FILL
XFILL_3__2443_ gnd vdd FILL
X_3012_ _3012_/A _3012_/B _3019_/A vdd gnd AND2X2
XFILL_8__3068_ gnd vdd FILL
XFILL_6__2152_ gnd vdd FILL
XFILL_0__2665_ gnd vdd FILL
XFILL_6__2083_ gnd vdd FILL
XFILL_8__2019_ gnd vdd FILL
XFILL_3__2374_ gnd vdd FILL
XFILL184050x148350 gnd vdd FILL
XFILL_0__2596_ gnd vdd FILL
XFILL_4_BUFX2_insert0 gnd vdd FILL
XFILL_1__2010_ gnd vdd FILL
XFILL_6__2985_ gnd vdd FILL
XFILL_0__3217_ gnd vdd FILL
XFILL_6__1936_ gnd vdd FILL
XFILL_9__2694_ gnd vdd FILL
XFILL_0__3148_ gnd vdd FILL
XFILL_6__1867_ gnd vdd FILL
XFILL_0__3079_ gnd vdd FILL
X_2727_ _3573_/Q _2770_/B _2770_/C _3359_/Q _2728_/C vdd gnd AOI22X1
XFILL_1__2912_ gnd vdd FILL
XFILL_6__1798_ gnd vdd FILL
XFILL_6__3537_ gnd vdd FILL
XFILL_7__2330_ gnd vdd FILL
XFILL_4__2621_ gnd vdd FILL
X_2658_ _2660_/A _2741_/C _2675_/A _2659_/C vdd gnd OAI21X1
XFILL_1__2843_ gnd vdd FILL
XFILL_4__2552_ gnd vdd FILL
X_2589_ _2589_/A _3166_/B _3166_/A _2589_/D _2726_/C vdd gnd OAI22X1
XFILL_6__3468_ gnd vdd FILL
XFILL_7__2261_ gnd vdd FILL
XFILL_1__2774_ gnd vdd FILL
XFILL_6__3399_ gnd vdd FILL
XFILL_6__2419_ gnd vdd FILL
XFILL_4__2483_ gnd vdd FILL
XFILL_7__2192_ gnd vdd FILL
XFILL_1__1725_ gnd vdd FILL
XFILL_4__3104_ gnd vdd FILL
XFILL184050x27450 gnd vdd FILL
XFILL_4__3035_ gnd vdd FILL
XFILL_2__2050_ gnd vdd FILL
XFILL_1__2208_ gnd vdd FILL
XFILL_7__1976_ gnd vdd FILL
XFILL184650x74250 gnd vdd FILL
XFILL_1__3188_ gnd vdd FILL
XFILL_1__2139_ gnd vdd FILL
XFILL_5__2730_ gnd vdd FILL
XFILL_2__2952_ gnd vdd FILL
XFILL_8__2370_ gnd vdd FILL
XFILL_2__1903_ gnd vdd FILL
XFILL_5__2661_ gnd vdd FILL
XFILL_4__2819_ gnd vdd FILL
XFILL_2__2883_ gnd vdd FILL
XFILL_5__2592_ gnd vdd FILL
XFILL_7_BUFX2_insert4 gnd vdd FILL
XFILL_7__2528_ gnd vdd FILL
XFILL_2__1834_ gnd vdd FILL
XFILL_7__2459_ gnd vdd FILL
XFILL_2__1765_ gnd vdd FILL
XFILL_2__3504_ gnd vdd FILL
XFILL_2__1696_ gnd vdd FILL
XFILL_5__3213_ gnd vdd FILL
XFILL_2__3435_ gnd vdd FILL
XFILL_5__3144_ gnd vdd FILL
XFILL_2__3366_ gnd vdd FILL
XFILL_0__2450_ gnd vdd FILL
XFILL_5__3075_ gnd vdd FILL
XFILL_2__2317_ gnd vdd FILL
XFILL_0__2381_ gnd vdd FILL
XFILL_5__2026_ gnd vdd FILL
XFILL_3__2090_ gnd vdd FILL
XFILL_2__2248_ gnd vdd FILL
X_1960_ _2499_/A _2416_/B vdd gnd INVX1
XFILL_2__2179_ gnd vdd FILL
XFILL_0__3002_ gnd vdd FILL
X_1891_ _1891_/A _1891_/B _3145_/B vdd gnd NAND2X1
XFILL_8__2706_ gnd vdd FILL
XFILL_6__2770_ gnd vdd FILL
XFILL_5__2928_ gnd vdd FILL
X_3561_ _3577_/Q _3563_/A vdd gnd INVX1
XFILL_3__2992_ gnd vdd FILL
XFILL_6__1721_ gnd vdd FILL
XFILL_8__2637_ gnd vdd FILL
XFILL_5__2859_ gnd vdd FILL
XFILL_3__1943_ gnd vdd FILL
X_2512_ _2512_/A _2512_/B _2513_/A vdd gnd NAND2X1
X_3492_ _3492_/A _3492_/B _3497_/C vdd gnd NAND2X1
XFILL_3__1874_ gnd vdd FILL
XFILL_8__2568_ gnd vdd FILL
XFILL_8__2499_ gnd vdd FILL
X_2443_ _3166_/B _2589_/D _2444_/A vdd gnd NAND2X1
XFILL_3__3544_ gnd vdd FILL
X_2374_ _2453_/A _2430_/B _2374_/C _2375_/B vdd gnd OAI21X1
XFILL_3__3475_ gnd vdd FILL
XFILL_6__2204_ gnd vdd FILL
XFILL_6__3184_ gnd vdd FILL
XFILL_0__2717_ gnd vdd FILL
XFILL_3__2426_ gnd vdd FILL
XFILL_1__2490_ gnd vdd FILL
XFILL_6__2135_ gnd vdd FILL
XFILL_0__2648_ gnd vdd FILL
XFILL_3__2357_ gnd vdd FILL
XFILL_0__2579_ gnd vdd FILL
XFILL_6__2066_ gnd vdd FILL
XFILL_1__3111_ gnd vdd FILL
XFILL_3__2288_ gnd vdd FILL
XFILL_7__1830_ gnd vdd FILL
XFILL_1__3042_ gnd vdd FILL
XFILL_5_BUFX2_insert80 gnd vdd FILL
XFILL_5_BUFX2_insert91 gnd vdd FILL
XFILL_6__2968_ gnd vdd FILL
XFILL_7__1761_ gnd vdd FILL
XFILL_7__3500_ gnd vdd FILL
XFILL_6__1919_ gnd vdd FILL
XFILL_7__1692_ gnd vdd FILL
XFILL_4__1983_ gnd vdd FILL
XFILL_6__2899_ gnd vdd FILL
XFILL_7__3431_ gnd vdd FILL
XFILL_4__2604_ gnd vdd FILL
XFILL_7__2313_ gnd vdd FILL
XFILL_1__2826_ gnd vdd FILL
XFILL_4__3584_ gnd vdd FILL
XFILL_7__2244_ gnd vdd FILL
XFILL_4__2535_ gnd vdd FILL
XFILL_4__2466_ gnd vdd FILL
XFILL_1__2757_ gnd vdd FILL
XFILL_1__1708_ gnd vdd FILL
XFILL_7__2175_ gnd vdd FILL
XFILL_1__2688_ gnd vdd FILL
XFILL_4__2397_ gnd vdd FILL
XFILL_2__3220_ gnd vdd FILL
XFILL_2__3151_ gnd vdd FILL
XFILL_2__2102_ gnd vdd FILL
XFILL_2__3082_ gnd vdd FILL
XFILL_8__1870_ gnd vdd FILL
XFILL_4__3018_ gnd vdd FILL
XFILL_2__2033_ gnd vdd FILL
XFILL_7__1959_ gnd vdd FILL
XFILL_8__3540_ gnd vdd FILL
XFILL_8__3471_ gnd vdd FILL
XFILL_5__2713_ gnd vdd FILL
XFILL_2__2935_ gnd vdd FILL
XFILL_8__2422_ gnd vdd FILL
XFILL_5__2644_ gnd vdd FILL
XFILL_2__2866_ gnd vdd FILL
XFILL_0__1950_ gnd vdd FILL
XFILL_8__2353_ gnd vdd FILL
XFILL_0__1881_ gnd vdd FILL
XFILL_5__2575_ gnd vdd FILL
XFILL_8__2284_ gnd vdd FILL
XFILL_2__1817_ gnd vdd FILL
XFILL_2__2797_ gnd vdd FILL
XFILL_2__1748_ gnd vdd FILL
XFILL_0__3551_ gnd vdd FILL
X_2090_ _2298_/A _3144_/C _2090_/C _2332_/A vdd gnd OAI21X1
XFILL_0__3482_ gnd vdd FILL
XFILL_2__3418_ gnd vdd FILL
XFILL_3__2211_ gnd vdd FILL
XFILL_0__2502_ gnd vdd FILL
XFILL_5__3127_ gnd vdd FILL
XFILL_3__3191_ gnd vdd FILL
XFILL_0__2433_ gnd vdd FILL
XFILL_5__3058_ gnd vdd FILL
XFILL_3__2142_ gnd vdd FILL
X_2992_ _2992_/A _3577_/Q _2993_/B _2993_/C vdd gnd OAI21X1
XFILL_3__2073_ gnd vdd FILL
XFILL_0__2364_ gnd vdd FILL
XFILL_5__2009_ gnd vdd FILL
XFILL_0__2295_ gnd vdd FILL
X_1943_ _3359_/Q _2691_/A _2728_/B vdd gnd NAND2X1
XFILL_8__1999_ gnd vdd FILL
XFILL_6__2822_ gnd vdd FILL
X_1874_ _1875_/A _1874_/B _1874_/C _1879_/A vdd gnd NAND3X1
XFILL_6__2753_ gnd vdd FILL
XFILL_3__2975_ gnd vdd FILL
XFILL_6__1704_ gnd vdd FILL
X_3544_ _3544_/A _3544_/B _3544_/C _3545_/B vdd gnd OAI21X1
XFILL_3__1926_ gnd vdd FILL
XFILL_1__1990_ gnd vdd FILL
XFILL_6__2684_ gnd vdd FILL
X_3475_ _3493_/B _3493_/A _3476_/A vdd gnd NOR2X1
XFILL_3__1857_ gnd vdd FILL
X_2426_ _2676_/B _2426_/B _2426_/C _2427_/C vdd gnd OAI21X1
XFILL_1__2611_ gnd vdd FILL
XFILL_3__1788_ gnd vdd FILL
XFILL_3__3527_ gnd vdd FILL
XFILL_1__3591_ gnd vdd FILL
XFILL_4__2320_ gnd vdd FILL
X_2357_ _2357_/A _2444_/B vdd gnd INVX1
XFILL_3__3458_ gnd vdd FILL
XFILL_4__2251_ gnd vdd FILL
X_2288_ _2298_/A _2288_/B _2288_/C _2797_/B _2344_/A vdd gnd AOI22X1
XFILL_1__2542_ gnd vdd FILL
XFILL_1__2473_ gnd vdd FILL
XFILL_6__3167_ gnd vdd FILL
XFILL_3__2409_ gnd vdd FILL
XFILL_6__3098_ gnd vdd FILL
XFILL_3__3389_ gnd vdd FILL
XFILL_4__2182_ gnd vdd FILL
XFILL_6__2118_ gnd vdd FILL
XFILL_6__2049_ gnd vdd FILL
XFILL_7__2931_ gnd vdd FILL
XFILL_7__2862_ gnd vdd FILL
XFILL_1__3025_ gnd vdd FILL
XFILL_7__1813_ gnd vdd FILL
XFILL_7__2793_ gnd vdd FILL
XFILL_4__1966_ gnd vdd FILL
XFILL_7__1744_ gnd vdd FILL
XFILL_5_CLKBUF1_insert38 gnd vdd FILL
XFILL_7__3414_ gnd vdd FILL
XFILL_4__1897_ gnd vdd FILL
XFILL_2__2720_ gnd vdd FILL
XFILL_5__2360_ gnd vdd FILL
XFILL_2__2651_ gnd vdd FILL
XFILL_1__2809_ gnd vdd FILL
XFILL_4__2518_ gnd vdd FILL
XFILL_2__2582_ gnd vdd FILL
XFILL_4__3498_ gnd vdd FILL
XFILL_7__2227_ gnd vdd FILL
XFILL_3_CLKBUF1_insert31 gnd vdd FILL
XFILL_5__2291_ gnd vdd FILL
XFILL_7__2158_ gnd vdd FILL
XFILL_4__2449_ gnd vdd FILL
XFILL_2__3203_ gnd vdd FILL
XFILL_8__2971_ gnd vdd FILL
XFILL_7__2089_ gnd vdd FILL
XFILL_2__3134_ gnd vdd FILL
XFILL_8__1922_ gnd vdd FILL
XFILL_2__3065_ gnd vdd FILL
XFILL_8__1853_ gnd vdd FILL
XFILL_0__2080_ gnd vdd FILL
XFILL_2__2016_ gnd vdd FILL
XFILL_8__1784_ gnd vdd FILL
XFILL_8__3523_ gnd vdd FILL
XFILL_8__3454_ gnd vdd FILL
XFILL_3__2760_ gnd vdd FILL
XFILL_0__2982_ gnd vdd FILL
XFILL_8__2405_ gnd vdd FILL
XFILL_3__1711_ gnd vdd FILL
XFILL_2__2918_ gnd vdd FILL
XFILL_8__3385_ gnd vdd FILL
XFILL_3__2691_ gnd vdd FILL
XFILL_0__1933_ gnd vdd FILL
XFILL_5__2627_ gnd vdd FILL
XFILL_2__2849_ gnd vdd FILL
X_3260_ _3260_/D vdd _3282_/R _3284_/CLK _3260_/Q vdd gnd DFFSR
XFILL_8__2336_ gnd vdd FILL
XFILL_5__2558_ gnd vdd FILL
XFILL_8__2267_ gnd vdd FILL
X_2211_ _2328_/A _2323_/A _2283_/B _2304_/A vdd gnd NOR3X1
XFILL_0__1864_ gnd vdd FILL
X_3191_ _3191_/A _3194_/C _3192_/C vdd gnd NOR2X1
XFILL_5__2489_ gnd vdd FILL
X_2142_ _2212_/A _3183_/B _2342_/A _2143_/C vdd gnd OAI21X1
XFILL_0__3603_ gnd vdd FILL
XFILL_8__2198_ gnd vdd FILL
XFILL_0__1795_ gnd vdd FILL
XFILL_0__3534_ gnd vdd FILL
X_2073_ _2073_/A _2073_/B _2329_/B _2074_/B vdd gnd NAND3X1
XFILL_6__3021_ gnd vdd FILL
XFILL_0__3465_ gnd vdd FILL
XFILL_3__3174_ gnd vdd FILL
XFILL_0__3396_ gnd vdd FILL
XFILL_0__2416_ gnd vdd FILL
XFILL_3__2125_ gnd vdd FILL
XFILL_0__2347_ gnd vdd FILL
X_2975_ _3309_/Q _2979_/A _2979_/C vdd gnd NAND2X1
XFILL_3__2056_ gnd vdd FILL
XFILL_6__2805_ gnd vdd FILL
X_1926_ _1985_/A _3571_/Q _1926_/C _1927_/C vdd gnd AOI21X1
XFILL_0__2278_ gnd vdd FILL
X_1857_ _3288_/Q _2924_/A vdd gnd INVX1
XFILL_4__1820_ gnd vdd FILL
XFILL_6__2736_ gnd vdd FILL
X_3527_ _3550_/B _3548_/B _3537_/C _3528_/A vdd gnd AOI21X1
XFILL_3__2958_ gnd vdd FILL
XFILL_4__1751_ gnd vdd FILL
XFILL_6__2667_ gnd vdd FILL
X_1788_ _1788_/A _3194_/A _1796_/A vdd gnd OR2X2
XFILL_3__2889_ gnd vdd FILL
XFILL_1__1973_ gnd vdd FILL
XFILL_3__1909_ gnd vdd FILL
XFILL_7__3130_ gnd vdd FILL
X_3458_ _3468_/S _3468_/B _3471_/B _3459_/B vdd gnd OAI21X1
XFILL_4__3421_ gnd vdd FILL
XFILL_6__2598_ gnd vdd FILL
X_3389_ _3519_/A _3485_/A _3519_/B _3391_/B vdd gnd AOI21X1
X_2409_ _3024_/A _2448_/B _2409_/C _2413_/A vdd gnd OAI21X1
XFILL_7__3061_ gnd vdd FILL
XFILL_4__2303_ gnd vdd FILL
XFILL_7__2012_ gnd vdd FILL
XFILL_1__2525_ gnd vdd FILL
XFILL_6__3219_ gnd vdd FILL
XFILL_4__2234_ gnd vdd FILL
XFILL_4__2165_ gnd vdd FILL
XFILL_1__2456_ gnd vdd FILL
XFILL_1__2387_ gnd vdd FILL
XFILL_7__2914_ gnd vdd FILL
XFILL_4__2096_ gnd vdd FILL
XFILL_5__1860_ gnd vdd FILL
XFILL_7__2845_ gnd vdd FILL
XFILL_1__3008_ gnd vdd FILL
XFILL_7__2776_ gnd vdd FILL
XFILL_4__2998_ gnd vdd FILL
XFILL_5__1791_ gnd vdd FILL
XFILL_7__1727_ gnd vdd FILL
XFILL_5__3530_ gnd vdd FILL
XFILL_4__1949_ gnd vdd FILL
XFILL_5__3461_ gnd vdd FILL
XFILL_5__2412_ gnd vdd FILL
XFILL_2__2703_ gnd vdd FILL
XFILL_8__3170_ gnd vdd FILL
XFILL_5__3392_ gnd vdd FILL
XFILL_8__2121_ gnd vdd FILL
XFILL_2__2634_ gnd vdd FILL
XFILL_5__2343_ gnd vdd FILL
XFILL_8__2052_ gnd vdd FILL
XFILL_5__2274_ gnd vdd FILL
XFILL_2__2565_ gnd vdd FILL
XFILL_2__2496_ gnd vdd FILL
XFILL_6_BUFX2_insert24 gnd vdd FILL
XFILL_6_BUFX2_insert13 gnd vdd FILL
XFILL_6_BUFX2_insert57 gnd vdd FILL
XFILL_8__2954_ gnd vdd FILL
XFILL_6_BUFX2_insert79 gnd vdd FILL
XFILL_6_BUFX2_insert68 gnd vdd FILL
XFILL_6_BUFX2_insert46 gnd vdd FILL
XFILL_2__3117_ gnd vdd FILL
XFILL_0__2201_ gnd vdd FILL
XFILL_0__3181_ gnd vdd FILL
XFILL_8__1905_ gnd vdd FILL
XFILL_8__2885_ gnd vdd FILL
XFILL_0__2132_ gnd vdd FILL
XFILL_2__3048_ gnd vdd FILL
XFILL_8__1836_ gnd vdd FILL
X_2760_ _3177_/B _2760_/B _2762_/C vdd gnd NOR2X1
XFILL_8__1767_ gnd vdd FILL
XFILL_0__2063_ gnd vdd FILL
X_1711_ _2993_/A _3297_/D vdd gnd INVX1
X_2691_ _2691_/A _2759_/A _2759_/B _2725_/C vdd gnd NOR3X1
XFILL_8__3506_ gnd vdd FILL
XFILL_5__1989_ gnd vdd FILL
XFILL_3__2812_ gnd vdd FILL
XFILL_6__2521_ gnd vdd FILL
XFILL_8__1698_ gnd vdd FILL
XFILL_8__3437_ gnd vdd FILL
XFILL_6__2452_ gnd vdd FILL
XFILL_3__2743_ gnd vdd FILL
XFILL_0__2965_ gnd vdd FILL
X_3312_ _3312_/D vdd _3313_/R _3578_/CLK _3312_/Q vdd gnd DFFSR
XFILL_8__3368_ gnd vdd FILL
XFILL_3__2674_ gnd vdd FILL
XFILL_0__2896_ gnd vdd FILL
XFILL_0__1916_ gnd vdd FILL
XFILL_6__2383_ gnd vdd FILL
XFILL_8__2319_ gnd vdd FILL
X_3243_ _3243_/D vdd _3355_/R _3355_/CLK _3243_/Q vdd gnd DFFSR
XFILL_0__1847_ gnd vdd FILL
X_3174_ _3174_/A _3174_/B _3175_/A vdd gnd NOR2X1
XFILL_6__3004_ gnd vdd FILL
X_2125_ _2299_/A _2446_/B _2278_/A _2126_/C vdd gnd OAI21X1
XFILL_0__1778_ gnd vdd FILL
XFILL_0__3517_ gnd vdd FILL
XFILL_1__2310_ gnd vdd FILL
X_2056_ _3011_/B _3003_/S vdd gnd INVX1
XFILL_3__3226_ gnd vdd FILL
XFILL_0__3448_ gnd vdd FILL
XFILL_1__2241_ gnd vdd FILL
XFILL_3__3157_ gnd vdd FILL
XFILL_0__3379_ gnd vdd FILL
XFILL_3__3088_ gnd vdd FILL
XFILL_1__2172_ gnd vdd FILL
XFILL183450x7950 gnd vdd FILL
XFILL_3__2108_ gnd vdd FILL
XFILL_4__2921_ gnd vdd FILL
XFILL_3__2039_ gnd vdd FILL
X_2958_ _2958_/A _2958_/B _2968_/A _2999_/B vdd gnd OAI21X1
XFILL_9__3546_ gnd vdd FILL
XFILL_7__2630_ gnd vdd FILL
X_1909_ _2435_/B _1910_/B vdd gnd INVX1
XFILL_4__2852_ gnd vdd FILL
X_2889_ _2889_/A _2889_/B _2889_/C _2891_/C vdd gnd OAI21X1
XFILL_7__2561_ gnd vdd FILL
XFILL_4__2783_ gnd vdd FILL
XFILL_4__1803_ gnd vdd FILL
XFILL_6__2719_ gnd vdd FILL
XFILL_7__2492_ gnd vdd FILL
XFILL_4__1734_ gnd vdd FILL
XFILL_1__1956_ gnd vdd FILL
XFILL_7__3113_ gnd vdd FILL
XFILL_4__3404_ gnd vdd FILL
XFILL_1__1887_ gnd vdd FILL
XFILL_1__3557_ gnd vdd FILL
XFILL_7__3044_ gnd vdd FILL
XFILL_2__2350_ gnd vdd FILL
XFILL_1__3488_ gnd vdd FILL
XFILL_4__2217_ gnd vdd FILL
XFILL_2__2281_ gnd vdd FILL
XFILL_1__2508_ gnd vdd FILL
XFILL_4__3197_ gnd vdd FILL
XFILL_1__2439_ gnd vdd FILL
XFILL_4__2148_ gnd vdd FILL
XFILL_4__2079_ gnd vdd FILL
XFILL_5__2961_ gnd vdd FILL
XFILL_8__2670_ gnd vdd FILL
XFILL_7__2828_ gnd vdd FILL
XFILL_5__2892_ gnd vdd FILL
XFILL_5__1912_ gnd vdd FILL
XFILL_5__1843_ gnd vdd FILL
XFILL_5__1774_ gnd vdd FILL
XFILL_7__2759_ gnd vdd FILL
XFILL_5__3513_ gnd vdd FILL
XFILL_2__1996_ gnd vdd FILL
XFILL_8__3222_ gnd vdd FILL
XFILL_5__3444_ gnd vdd FILL
XFILL_8__3153_ gnd vdd FILL
XFILL_0__2750_ gnd vdd FILL
XFILL_8__2104_ gnd vdd FILL
XFILL_5__3375_ gnd vdd FILL
XFILL_0__1701_ gnd vdd FILL
XFILL_8__3084_ gnd vdd FILL
XFILL_5__2326_ gnd vdd FILL
XFILL_3__2390_ gnd vdd FILL
XFILL_2__3597_ gnd vdd FILL
XFILL_0__2681_ gnd vdd FILL
XFILL_2__2617_ gnd vdd FILL
XFILL_8__2035_ gnd vdd FILL
XFILL_2__2548_ gnd vdd FILL
XFILL_5__2257_ gnd vdd FILL
XFILL_5__2188_ gnd vdd FILL
XFILL_3__3011_ gnd vdd FILL
XFILL_2__2479_ gnd vdd FILL
XFILL_8__2937_ gnd vdd FILL
XFILL_8__2868_ gnd vdd FILL
X_2812_ _2859_/A _2881_/A _2815_/A vdd gnd NAND2X1
XFILL_6__1952_ gnd vdd FILL
XFILL_0__3164_ gnd vdd FILL
XFILL_0__3095_ gnd vdd FILL
XFILL_8__1819_ gnd vdd FILL
XFILL_0__2115_ gnd vdd FILL
XFILL_6__1883_ gnd vdd FILL
X_2743_ _3197_/C _2743_/B _2744_/C vdd gnd NAND2X1
XFILL_8__2799_ gnd vdd FILL
XFILL_0__2046_ gnd vdd FILL
X_2674_ _2674_/A _2674_/B _2674_/C _2733_/B vdd gnd NAND3X1
XFILL_6__3553_ gnd vdd FILL
XFILL_2_BUFX2_insert11 gnd vdd FILL
XFILL_6__3484_ gnd vdd FILL
XFILL_1__2790_ gnd vdd FILL
XFILL_2_BUFX2_insert22 gnd vdd FILL
XFILL_6__2504_ gnd vdd FILL
XFILL_2_BUFX2_insert44 gnd vdd FILL
XFILL_1__1810_ gnd vdd FILL
XFILL_0__2948_ gnd vdd FILL
XFILL_2_BUFX2_insert88 gnd vdd FILL
XFILL_2_BUFX2_insert66 gnd vdd FILL
XFILL_2_BUFX2_insert55 gnd vdd FILL
XFILL_3__2726_ gnd vdd FILL
XFILL_1__1741_ gnd vdd FILL
XFILL_6__2435_ gnd vdd FILL
XFILL_2_BUFX2_insert77 gnd vdd FILL
XFILL_3__2657_ gnd vdd FILL
XFILL_0__2879_ gnd vdd FILL
XFILL_9__2075_ gnd vdd FILL
XFILL_6__2366_ gnd vdd FILL
X_3226_ _3226_/A _3232_/B _3226_/C _3360_/D vdd gnd OAI21X1
XFILL_3__2588_ gnd vdd FILL
XFILL_4__3120_ gnd vdd FILL
XFILL_1__3411_ gnd vdd FILL
XFILL_6__2297_ gnd vdd FILL
X_3157_ _3157_/A _3157_/B _3157_/C _3158_/C vdd gnd AOI21X1
X_2108_ _2108_/A _3156_/B _2357_/A vdd gnd NOR2X1
XFILL_4__3051_ gnd vdd FILL
X_3088_ _3088_/A _3297_/D _3088_/S _3143_/A vdd gnd MUX2X1
X_2039_ _2932_/A _2039_/B _2933_/C vdd gnd NOR2X1
XFILL_4__2002_ gnd vdd FILL
XFILL_3__3209_ gnd vdd FILL
XFILL_9__1928_ gnd vdd FILL
XFILL_7__1992_ gnd vdd FILL
XFILL_1__2224_ gnd vdd FILL
XFILL_1__2155_ gnd vdd FILL
XFILL_4__2904_ gnd vdd FILL
XFILL_1__2086_ gnd vdd FILL
XFILL_7__2613_ gnd vdd FILL
XFILL_4__2835_ gnd vdd FILL
XFILL_7__3593_ gnd vdd FILL
XFILL_7__2544_ gnd vdd FILL
XFILL_2__1850_ gnd vdd FILL
XFILL_7__2475_ gnd vdd FILL
XFILL_4__2766_ gnd vdd FILL
XFILL_8_CLKBUF1_insert31 gnd vdd FILL
XFILL_2__3520_ gnd vdd FILL
XFILL_1__2988_ gnd vdd FILL
XFILL_4__1717_ gnd vdd FILL
XFILL_4__2697_ gnd vdd FILL
XFILL_2__1781_ gnd vdd FILL
XFILL_0_CLKBUF1_insert28 gnd vdd FILL
XFILL_1__1939_ gnd vdd FILL
XFILL_2__3451_ gnd vdd FILL
XFILL_5__3160_ gnd vdd FILL
XFILL_2__3382_ gnd vdd FILL
XFILL_2__2402_ gnd vdd FILL
XFILL_5__2111_ gnd vdd FILL
XFILL_5__3091_ gnd vdd FILL
XFILL_7__3027_ gnd vdd FILL
XFILL_2__2333_ gnd vdd FILL
XFILL_5__2042_ gnd vdd FILL
XFILL_2__2264_ gnd vdd FILL
XFILL_2__2195_ gnd vdd FILL
XFILL_8__2722_ gnd vdd FILL
XFILL_5__2944_ gnd vdd FILL
XFILL181350x140550 gnd vdd FILL
XFILL_8__2653_ gnd vdd FILL
XFILL_5__2875_ gnd vdd FILL
XFILL_8__2584_ gnd vdd FILL
XFILL_3__1890_ gnd vdd FILL
XFILL_5__1826_ gnd vdd FILL
XFILL_5__1757_ gnd vdd FILL
XFILL_2__1979_ gnd vdd FILL
XFILL_3__3560_ gnd vdd FILL
XFILL_0__2802_ gnd vdd FILL
X_2390_ _2621_/B _2426_/B _2390_/C _2391_/C vdd gnd OAI21X1
XFILL_8__3205_ gnd vdd FILL
XFILL_3__3491_ gnd vdd FILL
XFILL_5__3427_ gnd vdd FILL
XFILL_9_BUFX2_insert83 gnd vdd FILL
XFILL_6__2220_ gnd vdd FILL
XFILL_3__2511_ gnd vdd FILL
XFILL_5__1688_ gnd vdd FILL
XFILL_8__3136_ gnd vdd FILL
XFILL_0__2733_ gnd vdd FILL
XFILL_3__2442_ gnd vdd FILL
XFILL_8__3067_ gnd vdd FILL
X_3011_ _3277_/Q _3011_/B _3017_/A _3012_/A vdd gnd AOI21X1
XFILL_6__2151_ gnd vdd FILL
XFILL_0__2664_ gnd vdd FILL
XFILL_9__2900_ gnd vdd FILL
XFILL_8__2018_ gnd vdd FILL
XFILL_5__2309_ gnd vdd FILL
XFILL_6__2082_ gnd vdd FILL
XFILL_3__2373_ gnd vdd FILL
XFILL_0__2595_ gnd vdd FILL
XFILL_6__2984_ gnd vdd FILL
XFILL_0__3216_ gnd vdd FILL
XFILL_4_BUFX2_insert1 gnd vdd FILL
XFILL_6__1935_ gnd vdd FILL
XFILL_0__3147_ gnd vdd FILL
XFILL_6__1866_ gnd vdd FILL
XFILL_0__3078_ gnd vdd FILL
X_2726_ _3147_/A _2958_/B _2726_/C _2772_/B vdd gnd OAI21X1
XFILL_1__2911_ gnd vdd FILL
XFILL_0__2029_ gnd vdd FILL
X_2657_ _2687_/A _2660_/A vdd gnd INVX1
XFILL_6__1797_ gnd vdd FILL
XFILL_1__2842_ gnd vdd FILL
XFILL_6__3536_ gnd vdd FILL
XFILL_4__2620_ gnd vdd FILL
XFILL_4__2551_ gnd vdd FILL
X_2588_ _2609_/B _2609_/A _2601_/C vdd gnd NAND2X1
XFILL_6__3467_ gnd vdd FILL
XFILL_7__2260_ gnd vdd FILL
XFILL_4__2482_ gnd vdd FILL
XFILL_3__2709_ gnd vdd FILL
XFILL_1__2773_ gnd vdd FILL
XFILL_6__3398_ gnd vdd FILL
XFILL_7__2191_ gnd vdd FILL
XFILL_6__2418_ gnd vdd FILL
XFILL_1__1724_ gnd vdd FILL
X_3209_ _3215_/A _3209_/B _3209_/C _3352_/D vdd gnd OAI21X1
XFILL_6__2349_ gnd vdd FILL
XFILL_4__3103_ gnd vdd FILL
XFILL_4__3034_ gnd vdd FILL
XFILL_1__2207_ gnd vdd FILL
XFILL_7__1975_ gnd vdd FILL
XFILL_1__3187_ gnd vdd FILL
XFILL_1__2138_ gnd vdd FILL
XFILL_2__2951_ gnd vdd FILL
XFILL_1__2069_ gnd vdd FILL
XFILL_2__1902_ gnd vdd FILL
XFILL_5__2660_ gnd vdd FILL
XFILL_4__2818_ gnd vdd FILL
XFILL_2__2882_ gnd vdd FILL
XFILL_7_BUFX2_insert5 gnd vdd FILL
XFILL_7__2527_ gnd vdd FILL
XFILL_5__2591_ gnd vdd FILL
XFILL_4__2749_ gnd vdd FILL
XFILL_2__1833_ gnd vdd FILL
XFILL_7__2458_ gnd vdd FILL
XFILL_2__1764_ gnd vdd FILL
XFILL_2__3503_ gnd vdd FILL
XFILL_7__2389_ gnd vdd FILL
XFILL_2__1695_ gnd vdd FILL
XFILL_5__3212_ gnd vdd FILL
XFILL_5__3143_ gnd vdd FILL
XFILL_2__3434_ gnd vdd FILL
XFILL_5__3074_ gnd vdd FILL
XFILL_2__3365_ gnd vdd FILL
XFILL_5__2025_ gnd vdd FILL
XFILL_0__2380_ gnd vdd FILL
XFILL_2__2316_ gnd vdd FILL
XFILL_2__2247_ gnd vdd FILL
XFILL_0__3001_ gnd vdd FILL
X_1890_ _2432_/A _2058_/B _3152_/C _3188_/A vdd gnd OAI21X1
XFILL_2__2178_ gnd vdd FILL
XFILL_8__2705_ gnd vdd FILL
XFILL_5__2927_ gnd vdd FILL
X_3560_ _3560_/A _3560_/B _3560_/C _3576_/D vdd gnd OAI21X1
XFILL_3__2991_ gnd vdd FILL
XFILL_6__1720_ gnd vdd FILL
XFILL_8__2636_ gnd vdd FILL
XFILL_5__2858_ gnd vdd FILL
XFILL_3__1942_ gnd vdd FILL
X_2511_ _2511_/A _3577_/Q _2511_/C _2512_/B vdd gnd AOI21X1
X_3491_ _3491_/A _3491_/B _3493_/A _3492_/A vdd gnd MUX2X1
XFILL_3__1873_ gnd vdd FILL
XFILL_5__1809_ gnd vdd FILL
XFILL_8__2567_ gnd vdd FILL
XFILL_5__2789_ gnd vdd FILL
XFILL_8__2498_ gnd vdd FILL
X_2442_ _2442_/A _2442_/B _2589_/D vdd gnd NOR2X1
XFILL_3__3543_ gnd vdd FILL
X_2373_ _3011_/B _2373_/B _2423_/A vdd gnd NOR2X1
XFILL_3__3474_ gnd vdd FILL
XFILL_8__3119_ gnd vdd FILL
XFILL_6__2203_ gnd vdd FILL
XFILL_0__2716_ gnd vdd FILL
XFILL_6__3183_ gnd vdd FILL
XFILL_3__2425_ gnd vdd FILL
XFILL_6__2134_ gnd vdd FILL
XFILL_3__2356_ gnd vdd FILL
XFILL_0__2647_ gnd vdd FILL
XFILL_0__2578_ gnd vdd FILL
XFILL_6__2065_ gnd vdd FILL
XFILL_1__3110_ gnd vdd FILL
XFILL_3__2287_ gnd vdd FILL
XFILL_1__3041_ gnd vdd FILL
XFILL_5_BUFX2_insert70 gnd vdd FILL
XFILL_5_BUFX2_insert92 gnd vdd FILL
XFILL_7__1760_ gnd vdd FILL
XFILL_6__2967_ gnd vdd FILL
XFILL_5_BUFX2_insert81 gnd vdd FILL
XFILL_6__1918_ gnd vdd FILL
XFILL_6__2898_ gnd vdd FILL
XFILL_7__1691_ gnd vdd FILL
XFILL_4__1982_ gnd vdd FILL
XFILL_7__3430_ gnd vdd FILL
X_2709_ _2732_/C _2724_/A vdd gnd INVX1
XFILL_6__1849_ gnd vdd FILL
XFILL_4__2603_ gnd vdd FILL
XFILL_1__2825_ gnd vdd FILL
XFILL_6__3519_ gnd vdd FILL
XFILL_7__2312_ gnd vdd FILL
XFILL_4__3583_ gnd vdd FILL
XFILL_7__2243_ gnd vdd FILL
XFILL_4__2534_ gnd vdd FILL
XFILL_4__2465_ gnd vdd FILL
XFILL_1__2756_ gnd vdd FILL
XFILL_4__2396_ gnd vdd FILL
XFILL_1__1707_ gnd vdd FILL
XFILL_7__2174_ gnd vdd FILL
XFILL_1__2687_ gnd vdd FILL
XFILL_2__3150_ gnd vdd FILL
XFILL_2__2101_ gnd vdd FILL
XFILL_2__3081_ gnd vdd FILL
XFILL_4__3017_ gnd vdd FILL
XFILL_2__2032_ gnd vdd FILL
XFILL_7__1958_ gnd vdd FILL
XFILL_8__3470_ gnd vdd FILL
XFILL_7__1889_ gnd vdd FILL
XFILL_8__2421_ gnd vdd FILL
XFILL_5__2712_ gnd vdd FILL
XFILL_2__2934_ gnd vdd FILL
XFILL_5__2643_ gnd vdd FILL
XFILL_7__3559_ gnd vdd FILL
XFILL_2__2865_ gnd vdd FILL
XFILL_8__2352_ gnd vdd FILL
XFILL_0__1880_ gnd vdd FILL
XFILL_2__1816_ gnd vdd FILL
XFILL_8__2283_ gnd vdd FILL
XFILL_5__2574_ gnd vdd FILL
XFILL_2__2796_ gnd vdd FILL
XFILL_0__3550_ gnd vdd FILL
XFILL_2__1747_ gnd vdd FILL
XFILL_0__2501_ gnd vdd FILL
XFILL_0__3481_ gnd vdd FILL
XFILL181950x148350 gnd vdd FILL
XFILL_2__3417_ gnd vdd FILL
XFILL_3__2210_ gnd vdd FILL
XFILL_3__3190_ gnd vdd FILL
XFILL_5__3126_ gnd vdd FILL
XFILL_3__2141_ gnd vdd FILL
XFILL_0__2432_ gnd vdd FILL
XFILL_5__3057_ gnd vdd FILL
XFILL_0__2363_ gnd vdd FILL
X_2991_ _3011_/B _2991_/B _2999_/D _2998_/A vdd gnd OAI21X1
XFILL_3__2072_ gnd vdd FILL
XFILL_5__2008_ gnd vdd FILL
XFILL_8__1998_ gnd vdd FILL
X_1942_ _2484_/A _1946_/B vdd gnd INVX1
XFILL_0__2294_ gnd vdd FILL
X_1873_ _1873_/A _1873_/B _1874_/C vdd gnd AND2X2
XFILL_6__2821_ gnd vdd FILL
XFILL_6__2752_ gnd vdd FILL
XFILL_3__2974_ gnd vdd FILL
XFILL_6__1703_ gnd vdd FILL
X_3543_ _3544_/C _3543_/B _3543_/C _3546_/A vdd gnd AOI21X1
XFILL_8__3599_ gnd vdd FILL
XFILL_3__1925_ gnd vdd FILL
XFILL_6__2683_ gnd vdd FILL
XFILL_8__2619_ gnd vdd FILL
X_3474_ _3544_/A _3474_/B _3543_/B _3543_/C _3494_/A vdd gnd AOI22X1
X_2425_ _3311_/Q _2425_/B _2426_/C vdd gnd NAND2X1
XFILL_3__1856_ gnd vdd FILL
XFILL_1__2610_ gnd vdd FILL
XFILL_3__1787_ gnd vdd FILL
XFILL_3__3526_ gnd vdd FILL
X_2356_ _2356_/A _2579_/B vdd gnd INVX2
XFILL_1__3590_ gnd vdd FILL
XFILL_4__2250_ gnd vdd FILL
XFILL_3__3457_ gnd vdd FILL
X_2287_ _2326_/A _2287_/B _3235_/D vdd gnd OR2X2
XFILL_1__2541_ gnd vdd FILL
XFILL_1__2472_ gnd vdd FILL
XFILL_6__3166_ gnd vdd FILL
XFILL_3__2408_ gnd vdd FILL
XFILL_3__3388_ gnd vdd FILL
XFILL_4__2181_ gnd vdd FILL
XFILL_6__3097_ gnd vdd FILL
XFILL_6__2117_ gnd vdd FILL
XFILL_7__2930_ gnd vdd FILL
XFILL_3__2339_ gnd vdd FILL
XFILL_6__2048_ gnd vdd FILL
XFILL_7__2861_ gnd vdd FILL
XFILL_7__2792_ gnd vdd FILL
XFILL_1__3024_ gnd vdd FILL
XFILL_7__1812_ gnd vdd FILL
XFILL_7__1743_ gnd vdd FILL
XFILL_4__1965_ gnd vdd FILL
XFILL_5_CLKBUF1_insert28 gnd vdd FILL
XFILL_7__3413_ gnd vdd FILL
XFILL_4__1896_ gnd vdd FILL
XFILL_4__3566_ gnd vdd FILL
XFILL_2__2650_ gnd vdd FILL
XFILL_1__2808_ gnd vdd FILL
XFILL_5__2290_ gnd vdd FILL
XFILL_4__2517_ gnd vdd FILL
XFILL_2__2581_ gnd vdd FILL
XFILL_4__3497_ gnd vdd FILL
XFILL_3_CLKBUF1_insert32 gnd vdd FILL
XFILL_7__2226_ gnd vdd FILL
XFILL_1__2739_ gnd vdd FILL
XFILL_1_BUFX2_insert90 gnd vdd FILL
XFILL_7__2157_ gnd vdd FILL
XFILL_4__2448_ gnd vdd FILL
XFILL_4__2379_ gnd vdd FILL
XFILL_2__3202_ gnd vdd FILL
XFILL_8__2970_ gnd vdd FILL
XFILL_7__2088_ gnd vdd FILL
XFILL_2__3133_ gnd vdd FILL
XFILL_8__1921_ gnd vdd FILL
XFILL_2__3064_ gnd vdd FILL
XFILL_8__1852_ gnd vdd FILL
XFILL_2__2015_ gnd vdd FILL
XFILL_8__3522_ gnd vdd FILL
XFILL_8__1783_ gnd vdd FILL
XFILL_8__3453_ gnd vdd FILL
XFILL_2__2917_ gnd vdd FILL
XFILL_8__3384_ gnd vdd FILL
XFILL_0__2981_ gnd vdd FILL
XFILL_8__2404_ gnd vdd FILL
XFILL_3__1710_ gnd vdd FILL
XFILL_0__1932_ gnd vdd FILL
XFILL_8__2335_ gnd vdd FILL
XFILL_3__2690_ gnd vdd FILL
XFILL_5__2626_ gnd vdd FILL
XFILL_2__2848_ gnd vdd FILL
X_2210_ _2210_/A _2322_/A _2283_/B vdd gnd NAND2X1
XFILL_5__2557_ gnd vdd FILL
XFILL_8__2266_ gnd vdd FILL
XFILL_0__1863_ gnd vdd FILL
XFILL_2__2779_ gnd vdd FILL
X_3190_ _3194_/B _3190_/B _3194_/C vdd gnd OR2X2
XFILL_8__2197_ gnd vdd FILL
XFILL_0__3602_ gnd vdd FILL
XFILL_5__2488_ gnd vdd FILL
X_2141_ _3158_/B _3171_/B vdd gnd INVX1
XFILL_0__1794_ gnd vdd FILL
XFILL_0__3533_ gnd vdd FILL
X_2072_ _2242_/A _2072_/B _2073_/A vdd gnd NAND2X1
XFILL_6__3020_ gnd vdd FILL
XFILL_0__3464_ gnd vdd FILL
XFILL_5__3109_ gnd vdd FILL
XFILL_0__2415_ gnd vdd FILL
XFILL_3__3173_ gnd vdd FILL
XFILL_0__3395_ gnd vdd FILL
XFILL_3__2124_ gnd vdd FILL
X_2974_ _3006_/B _2974_/B _2999_/B _2979_/A vdd gnd OAI21X1
XFILL_0__2346_ gnd vdd FILL
XFILL_3__2055_ gnd vdd FILL
X_1925_ _3043_/A _1984_/B _1925_/C _1926_/C vdd gnd OAI21X1
XFILL_0__2277_ gnd vdd FILL
XFILL_6__2804_ gnd vdd FILL
X_1856_ _1856_/A _1856_/B _1860_/A vdd gnd NOR2X1
XFILL_6__2735_ gnd vdd FILL
X_1787_ _2292_/B _3156_/B _2199_/B _1788_/A vdd gnd OAI21X1
X_3526_ _3526_/A _3526_/B _3550_/B vdd gnd XOR2X1
XFILL_3__2957_ gnd vdd FILL
XFILL_4__1750_ gnd vdd FILL
XFILL_6__2666_ gnd vdd FILL
XFILL_3__2888_ gnd vdd FILL
XFILL_1__1972_ gnd vdd FILL
XFILL_3__1908_ gnd vdd FILL
X_3457_ _3521_/B _3471_/B vdd gnd INVX1
XFILL_4__3420_ gnd vdd FILL
XFILL_3__1839_ gnd vdd FILL
XFILL_6__2597_ gnd vdd FILL
X_3388_ _3514_/B _3514_/A _3485_/A vdd gnd NOR2X1
X_2408_ _2966_/A _3145_/B _3088_/S _2413_/D vdd gnd OAI21X1
XFILL_3__3509_ gnd vdd FILL
XFILL_7__3060_ gnd vdd FILL
X_2339_ _2339_/A _2339_/B _2339_/C _2353_/B vdd gnd NAND3X1
XFILL_4__2302_ gnd vdd FILL
XFILL_7__2011_ gnd vdd FILL
XFILL_1__2524_ gnd vdd FILL
XFILL_6__3218_ gnd vdd FILL
XFILL_4__2233_ gnd vdd FILL
XFILL_6__3149_ gnd vdd FILL
XFILL_4__2164_ gnd vdd FILL
XFILL_1__2455_ gnd vdd FILL
XFILL_1__2386_ gnd vdd FILL
XFILL_7__2913_ gnd vdd FILL
XFILL_4__2095_ gnd vdd FILL
XFILL_7__2844_ gnd vdd FILL
XFILL_1__3007_ gnd vdd FILL
XFILL_7__2775_ gnd vdd FILL
XFILL_4__2997_ gnd vdd FILL
XFILL_7__1726_ gnd vdd FILL
XFILL_5__1790_ gnd vdd FILL
XFILL_4__1948_ gnd vdd FILL
XFILL_4__1879_ gnd vdd FILL
XFILL_5__3460_ gnd vdd FILL
XFILL_2__2702_ gnd vdd FILL
XFILL_5__2411_ gnd vdd FILL
XFILL_5__3391_ gnd vdd FILL
XFILL_8__2120_ gnd vdd FILL
XFILL_2__2633_ gnd vdd FILL
XFILL_4__3549_ gnd vdd FILL
XFILL_8__2051_ gnd vdd FILL
XFILL_5__2342_ gnd vdd FILL
XFILL_5__2273_ gnd vdd FILL
XFILL_7__2209_ gnd vdd FILL
XFILL_2__2564_ gnd vdd FILL
XFILL_2__2495_ gnd vdd FILL
XFILL_7__3189_ gnd vdd FILL
XFILL_6_BUFX2_insert25 gnd vdd FILL
XFILL_6_BUFX2_insert14 gnd vdd FILL
XFILL_6_BUFX2_insert58 gnd vdd FILL
XFILL_8__2953_ gnd vdd FILL
XFILL_6_BUFX2_insert47 gnd vdd FILL
XFILL_6_BUFX2_insert69 gnd vdd FILL
XFILL_2__3116_ gnd vdd FILL
XFILL_0__2200_ gnd vdd FILL
XFILL_0__3180_ gnd vdd FILL
XFILL_8__1904_ gnd vdd FILL
XFILL_8__2884_ gnd vdd FILL
XFILL_0__2131_ gnd vdd FILL
XFILL_2__3047_ gnd vdd FILL
XFILL183750x74250 gnd vdd FILL
XFILL_8__1835_ gnd vdd FILL
XFILL_0__2062_ gnd vdd FILL
XFILL_8__1766_ gnd vdd FILL
X_1710_ DI[7] _3297_/Q _3197_/C _2993_/A vdd gnd MUX2X1
X_2690_ _3024_/A _3147_/A _3189_/A _3173_/B _2759_/B vdd gnd AOI22X1
XFILL_3__2811_ gnd vdd FILL
XFILL_8__3505_ gnd vdd FILL
XFILL_5__1988_ gnd vdd FILL
XFILL_8__3436_ gnd vdd FILL
XFILL_8__1697_ gnd vdd FILL
XFILL_6__2520_ gnd vdd FILL
X_3311_ _3311_/D vdd _3353_/R _3313_/CLK _3311_/Q vdd gnd DFFSR
XFILL_6__2451_ gnd vdd FILL
XFILL_3__2742_ gnd vdd FILL
XFILL_0__2964_ gnd vdd FILL
XFILL_8__3367_ gnd vdd FILL
XFILL_5__2609_ gnd vdd FILL
XFILL_3__2673_ gnd vdd FILL
XFILL183450x148350 gnd vdd FILL
XFILL_0__2895_ gnd vdd FILL
XFILL_8__2318_ gnd vdd FILL
XFILL_6__2382_ gnd vdd FILL
XFILL_0__1915_ gnd vdd FILL
XFILL_5__3589_ gnd vdd FILL
X_3242_ _3242_/D vdd _3291_/R _3355_/CLK _3242_/Q vdd gnd DFFSR
XFILL_8__2249_ gnd vdd FILL
XFILL_0__1846_ gnd vdd FILL
X_3173_ _3237_/Q _3173_/B _3173_/C _3174_/B vdd gnd OAI21X1
X_2124_ _2430_/A _2958_/B _3017_/A vdd gnd NOR2X1
XFILL_6__3003_ gnd vdd FILL
XFILL_0__1777_ gnd vdd FILL
XFILL_0__3516_ gnd vdd FILL
X_2055_ _2958_/A _2448_/B _3011_/B vdd gnd NOR2X1
XFILL_3__3225_ gnd vdd FILL
XFILL_0__3447_ gnd vdd FILL
XFILL_1__2240_ gnd vdd FILL
XFILL_1__2171_ gnd vdd FILL
XFILL_3__3156_ gnd vdd FILL
XFILL_0__3378_ gnd vdd FILL
XFILL_3__3087_ gnd vdd FILL
XFILL_3__2107_ gnd vdd FILL
XFILL_4__2920_ gnd vdd FILL
XFILL_3__2038_ gnd vdd FILL
X_2957_ _2957_/A _2957_/B _2957_/C _3307_/D vdd gnd OAI21X1
XFILL_0__2329_ gnd vdd FILL
X_2888_ _2906_/A _2888_/B _3283_/Q _2892_/C vdd gnd OAI21X1
X_1908_ _3024_/A _2446_/B _2717_/C _2435_/B vdd gnd OAI21X1
XFILL_4__2851_ gnd vdd FILL
X_1839_ _1861_/B _1843_/B vdd gnd INVX1
XFILL_7__2560_ gnd vdd FILL
XFILL_6__2718_ gnd vdd FILL
XFILL_4__2782_ gnd vdd FILL
XFILL_4__1802_ gnd vdd FILL
XFILL_7__2491_ gnd vdd FILL
XFILL_4__1733_ gnd vdd FILL
X_3509_ _3514_/A _3514_/B _3509_/C _3510_/A vdd gnd OAI21X1
XFILL_1__1955_ gnd vdd FILL
XFILL_6__2649_ gnd vdd FILL
XFILL_4__3403_ gnd vdd FILL
XFILL_7__3112_ gnd vdd FILL
XFILL_1__1886_ gnd vdd FILL
XFILL_7__3043_ gnd vdd FILL
XFILL_1__3556_ gnd vdd FILL
XFILL_1__3487_ gnd vdd FILL
XFILL_4__2216_ gnd vdd FILL
XFILL_2__2280_ gnd vdd FILL
XFILL_1__2507_ gnd vdd FILL
XFILL_4__3196_ gnd vdd FILL
XFILL_1__2438_ gnd vdd FILL
XFILL_4__2147_ gnd vdd FILL
XFILL_4__2078_ gnd vdd FILL
XFILL_5__2960_ gnd vdd FILL
XFILL_1__2369_ gnd vdd FILL
XFILL_5__1911_ gnd vdd FILL
XFILL_5__2891_ gnd vdd FILL
XFILL_7__2827_ gnd vdd FILL
XFILL_5__1842_ gnd vdd FILL
XFILL_7__2758_ gnd vdd FILL
XFILL_7__1709_ gnd vdd FILL
XFILL_5__1773_ gnd vdd FILL
XFILL_5__3512_ gnd vdd FILL
XFILL_7__2689_ gnd vdd FILL
XFILL_2__1995_ gnd vdd FILL
XFILL_8__3221_ gnd vdd FILL
XFILL_5__3443_ gnd vdd FILL
XFILL_8__3152_ gnd vdd FILL
XFILL_5__3374_ gnd vdd FILL
XFILL_0__1700_ gnd vdd FILL
XFILL_0__2680_ gnd vdd FILL
XFILL_8__2103_ gnd vdd FILL
XFILL_8__3083_ gnd vdd FILL
XFILL_5__2325_ gnd vdd FILL
XFILL_2__3596_ gnd vdd FILL
XFILL184050x7950 gnd vdd FILL
XFILL_2__2616_ gnd vdd FILL
XFILL_8__2034_ gnd vdd FILL
XFILL_2__2547_ gnd vdd FILL
XFILL_5__2256_ gnd vdd FILL
XFILL_3__3010_ gnd vdd FILL
XFILL_5__2187_ gnd vdd FILL
XFILL_2__2478_ gnd vdd FILL
XFILL_0__3232_ gnd vdd FILL
XFILL_8__2936_ gnd vdd FILL
XFILL_8__2867_ gnd vdd FILL
X_2811_ _2811_/A _2859_/A vdd gnd INVX1
XFILL_6__1951_ gnd vdd FILL
XFILL_0__3163_ gnd vdd FILL
XFILL_0__3094_ gnd vdd FILL
XFILL_0__2114_ gnd vdd FILL
XFILL_6__1882_ gnd vdd FILL
XFILL_8__1818_ gnd vdd FILL
X_2742_ _2775_/C _2752_/A _2743_/B vdd gnd XOR2X1
XFILL_8__2798_ gnd vdd FILL
XFILL_0__2045_ gnd vdd FILL
XFILL_6__3552_ gnd vdd FILL
XFILL_8__1749_ gnd vdd FILL
X_2673_ _2673_/A _2673_/B _2675_/C vdd gnd NAND2X1
XFILL_6__2503_ gnd vdd FILL
XFILL_6__3483_ gnd vdd FILL
XFILL_2_BUFX2_insert23 gnd vdd FILL
XFILL_8__3419_ gnd vdd FILL
XFILL_2_BUFX2_insert12 gnd vdd FILL
XFILL_3__2725_ gnd vdd FILL
XFILL_2_BUFX2_insert45 gnd vdd FILL
XFILL_0__2947_ gnd vdd FILL
XFILL_2_BUFX2_insert56 gnd vdd FILL
XFILL_2_BUFX2_insert78 gnd vdd FILL
XFILL_1__1740_ gnd vdd FILL
XFILL_2_BUFX2_insert67 gnd vdd FILL
XFILL_6__2434_ gnd vdd FILL
XFILL_6__2365_ gnd vdd FILL
X_3225_ _3583_/A _3232_/B _3226_/C vdd gnd NAND2X1
XFILL_3__2656_ gnd vdd FILL
XFILL_2_BUFX2_insert89 gnd vdd FILL
XFILL_0__2878_ gnd vdd FILL
XFILL_3__2587_ gnd vdd FILL
XFILL_1__3410_ gnd vdd FILL
XFILL_6__2296_ gnd vdd FILL
XFILL_0__1829_ gnd vdd FILL
X_3156_ _3165_/A _3156_/B _3156_/C _3159_/A vdd gnd OAI21X1
X_3087_ _3087_/A _3087_/B _3088_/A vdd gnd XOR2X1
X_2107_ _2349_/B _2107_/B _2332_/C vdd gnd NOR2X1
X_2038_ _2249_/A _2039_/B vdd gnd INVX1
XFILL_4__3050_ gnd vdd FILL
XFILL_4__2001_ gnd vdd FILL
XFILL_3__3208_ gnd vdd FILL
XFILL_3__3139_ gnd vdd FILL
XFILL_7__1991_ gnd vdd FILL
XFILL_1__2223_ gnd vdd FILL
XFILL_1__2154_ gnd vdd FILL
XFILL_1__2085_ gnd vdd FILL
XFILL_4__2903_ gnd vdd FILL
XFILL_7__2612_ gnd vdd FILL
XFILL_4__2834_ gnd vdd FILL
XFILL_7__3592_ gnd vdd FILL
XFILL_7__2543_ gnd vdd FILL
XFILL_8_CLKBUF1_insert32 gnd vdd FILL
XFILL_7__2474_ gnd vdd FILL
XFILL_4__2765_ gnd vdd FILL
XFILL_1__2987_ gnd vdd FILL
XFILL_2__1780_ gnd vdd FILL
XFILL_4__2696_ gnd vdd FILL
XFILL_4__1716_ gnd vdd FILL
XFILL_1__1938_ gnd vdd FILL
XFILL_2__3450_ gnd vdd FILL
XFILL_1__1869_ gnd vdd FILL
XFILL_0_CLKBUF1_insert29 gnd vdd FILL
XFILL_2__3381_ gnd vdd FILL
XFILL_2__2401_ gnd vdd FILL
XFILL_5__2110_ gnd vdd FILL
XFILL_5__3090_ gnd vdd FILL
XFILL_1__3539_ gnd vdd FILL
XFILL_7__3026_ gnd vdd FILL
XFILL_2__2332_ gnd vdd FILL
XFILL_5__2041_ gnd vdd FILL
XFILL_2__2263_ gnd vdd FILL
XFILL_4__3179_ gnd vdd FILL
XFILL_2__2194_ gnd vdd FILL
XFILL_8__2721_ gnd vdd FILL
XFILL_5__2943_ gnd vdd FILL
XFILL_8__2652_ gnd vdd FILL
XFILL_5__2874_ gnd vdd FILL
XFILL_5__1825_ gnd vdd FILL
XFILL_8__2583_ gnd vdd FILL
XFILL_5__1756_ gnd vdd FILL
XFILL_2__1978_ gnd vdd FILL
XFILL_0__2801_ gnd vdd FILL
XFILL_8__3204_ gnd vdd FILL
XFILL_3__3490_ gnd vdd FILL
XFILL_5__3426_ gnd vdd FILL
XFILL_3__2510_ gnd vdd FILL
XFILL_8__3135_ gnd vdd FILL
XFILL_0__2732_ gnd vdd FILL
XFILL_3__2441_ gnd vdd FILL
XFILL_8__3066_ gnd vdd FILL
X_3010_ _3015_/A _3010_/B _3010_/C _3012_/B vdd gnd OAI21X1
XFILL_6__2150_ gnd vdd FILL
XFILL_0__2663_ gnd vdd FILL
XFILL_3__2372_ gnd vdd FILL
XFILL_8__2017_ gnd vdd FILL
XFILL_6__2081_ gnd vdd FILL
XFILL_5__2308_ gnd vdd FILL
XFILL_2__3579_ gnd vdd FILL
XFILL_5__2239_ gnd vdd FILL
XFILL_0__2594_ gnd vdd FILL
XFILL_8__2919_ gnd vdd FILL
XFILL_6__2983_ gnd vdd FILL
XFILL_0__3215_ gnd vdd FILL
XFILL_4_BUFX2_insert2 gnd vdd FILL
XFILL_6__1934_ gnd vdd FILL
XFILL_0__3146_ gnd vdd FILL
XFILL_6__1865_ gnd vdd FILL
XFILL_0__3077_ gnd vdd FILL
X_2725_ _2993_/B _2889_/C _2725_/C _2725_/D _2773_/B vdd gnd AOI22X1
XFILL_1__2910_ gnd vdd FILL
XFILL_0__2028_ gnd vdd FILL
XFILL_6__1796_ gnd vdd FILL
X_2656_ _2656_/A _2656_/B _2656_/C _2656_/D _2687_/A vdd gnd AOI22X1
XFILL_1__2841_ gnd vdd FILL
XFILL_6__3535_ gnd vdd FILL
XFILL_6__3466_ gnd vdd FILL
X_2587_ _2587_/A _2587_/B _2609_/B vdd gnd NOR2X1
XFILL_4__2550_ gnd vdd FILL
XFILL_6__2417_ gnd vdd FILL
XFILL_4__2481_ gnd vdd FILL
XFILL_3__2708_ gnd vdd FILL
XFILL_1__2772_ gnd vdd FILL
XFILL_6__3397_ gnd vdd FILL
XFILL_7__2190_ gnd vdd FILL
XFILL_1__1723_ gnd vdd FILL
XFILL_3__2639_ gnd vdd FILL
XFILL_6__2348_ gnd vdd FILL
X_3208_ _3214_/A _3214_/B _3352_/Q _3209_/C vdd gnd OAI21X1
X_3139_ _3139_/A _3143_/B _3139_/C _3345_/D vdd gnd OAI21X1
XFILL_6__2279_ gnd vdd FILL
XFILL_4__3102_ gnd vdd FILL
XFILL_4__3033_ gnd vdd FILL
XFILL_1__2206_ gnd vdd FILL
XFILL_9__2959_ gnd vdd FILL
XFILL_7__1974_ gnd vdd FILL
XFILL_1__3186_ gnd vdd FILL
XFILL_1__2137_ gnd vdd FILL
XFILL_2__2950_ gnd vdd FILL
XFILL_1__2068_ gnd vdd FILL
XFILL_2__1901_ gnd vdd FILL
XFILL_4__2817_ gnd vdd FILL
XFILL_2__2881_ gnd vdd FILL
XFILL_7_BUFX2_insert6 gnd vdd FILL
XFILL_5__2590_ gnd vdd FILL
XFILL_7__2526_ gnd vdd FILL
XFILL_2__1832_ gnd vdd FILL
XFILL_4__2748_ gnd vdd FILL
XFILL_7__2457_ gnd vdd FILL
XFILL_2__1763_ gnd vdd FILL
XFILL_2__3502_ gnd vdd FILL
XFILL_7__2388_ gnd vdd FILL
XFILL_5__3211_ gnd vdd FILL
XFILL_4__2679_ gnd vdd FILL
XFILL_2__3433_ gnd vdd FILL
XFILL_2__1694_ gnd vdd FILL
XFILL_5__3142_ gnd vdd FILL
XFILL_7__3009_ gnd vdd FILL
XFILL_5__3073_ gnd vdd FILL
XFILL_2__3364_ gnd vdd FILL
XFILL_5__2024_ gnd vdd FILL
XFILL_2__2315_ gnd vdd FILL
XFILL_2__2246_ gnd vdd FILL
XFILL_0__3000_ gnd vdd FILL
XFILL_2__2177_ gnd vdd FILL
XFILL_5__2926_ gnd vdd FILL
XFILL_3__2990_ gnd vdd FILL
XFILL_8__2704_ gnd vdd FILL
XFILL_3__1941_ gnd vdd FILL
XFILL_8__2635_ gnd vdd FILL
X_3490_ _3514_/A _3514_/B _3491_/B _3491_/A vdd gnd OAI21X1
XFILL_5__2857_ gnd vdd FILL
X_2510_ _2993_/A _2510_/B _2669_/A _2510_/D _2511_/C vdd gnd OAI22X1
XFILL_8__2566_ gnd vdd FILL
XFILL_3__1872_ gnd vdd FILL
XFILL_5__2788_ gnd vdd FILL
XFILL_5__1808_ gnd vdd FILL
X_2441_ _2699_/B _2441_/B _2441_/C _2569_/A vdd gnd NAND3X1
XFILL_8__2497_ gnd vdd FILL
XFILL_5__1739_ gnd vdd FILL
XFILL_3__3542_ gnd vdd FILL
X_2372_ _2863_/A _2579_/B _3442_/B vdd gnd NOR2X1
XFILL_8__3118_ gnd vdd FILL
XFILL_3__3473_ gnd vdd FILL
XFILL_5__3409_ gnd vdd FILL
XFILL_6__2202_ gnd vdd FILL
XFILL_0__2715_ gnd vdd FILL
XFILL_6__3182_ gnd vdd FILL
XFILL_3__2424_ gnd vdd FILL
XFILL_6__2133_ gnd vdd FILL
XFILL_8__3049_ gnd vdd FILL
XFILL_3__2355_ gnd vdd FILL
XFILL_0__2646_ gnd vdd FILL
XFILL_0__2577_ gnd vdd FILL
XFILL_6__2064_ gnd vdd FILL
XFILL_3__2286_ gnd vdd FILL
XFILL_1__3040_ gnd vdd FILL
XFILL_5_BUFX2_insert60 gnd vdd FILL
XFILL_5_BUFX2_insert71 gnd vdd FILL
XFILL_5_BUFX2_insert93 gnd vdd FILL
XFILL_5_BUFX2_insert82 gnd vdd FILL
XFILL_6__2966_ gnd vdd FILL
XFILL_0__3129_ gnd vdd FILL
XFILL_6__1917_ gnd vdd FILL
XFILL_6__2897_ gnd vdd FILL
XFILL_7__1690_ gnd vdd FILL
XFILL_4__1981_ gnd vdd FILL
X_2708_ _2708_/A _2708_/B _2708_/C _2708_/D _2732_/C vdd gnd AOI22X1
XFILL_6__1848_ gnd vdd FILL
XFILL_6__3518_ gnd vdd FILL
XFILL_7__2311_ gnd vdd FILL
XFILL_4__2602_ gnd vdd FILL
XFILL_4__3582_ gnd vdd FILL
X_2639_ _2639_/A _2639_/B _2639_/C _2741_/C vdd gnd NAND3X1
XFILL_6__1779_ gnd vdd FILL
XFILL_1__2824_ gnd vdd FILL
XFILL_4__2533_ gnd vdd FILL
XFILL_6__3449_ gnd vdd FILL
XFILL_7__2242_ gnd vdd FILL
XFILL_1__2755_ gnd vdd FILL
XFILL_7__2173_ gnd vdd FILL
XFILL_1__1706_ gnd vdd FILL
XFILL_4__2464_ gnd vdd FILL
XFILL_4__2395_ gnd vdd FILL
XFILL_1__2686_ gnd vdd FILL
XFILL_2__2100_ gnd vdd FILL
XFILL_2__3080_ gnd vdd FILL
XFILL_4__3016_ gnd vdd FILL
XFILL_2__2031_ gnd vdd FILL
XFILL_7__1957_ gnd vdd FILL
XFILL_1__3169_ gnd vdd FILL
XFILL_7__1888_ gnd vdd FILL
XFILL_8__2420_ gnd vdd FILL
XFILL_5__2711_ gnd vdd FILL
XFILL_2__2933_ gnd vdd FILL
XFILL_5__2642_ gnd vdd FILL
XFILL_7__3558_ gnd vdd FILL
XFILL_2__2864_ gnd vdd FILL
XFILL_8__2351_ gnd vdd FILL
XFILL_7__3489_ gnd vdd FILL
XFILL_8__2282_ gnd vdd FILL
XFILL_7__2509_ gnd vdd FILL
XFILL_5__2573_ gnd vdd FILL
XFILL_2__1815_ gnd vdd FILL
XFILL_2__2795_ gnd vdd FILL
XFILL_2__1746_ gnd vdd FILL
XFILL_0__2500_ gnd vdd FILL
XFILL_0__3480_ gnd vdd FILL
XFILL_5__3125_ gnd vdd FILL
XFILL_2__3416_ gnd vdd FILL
XFILL_3__2140_ gnd vdd FILL
XFILL_0__2431_ gnd vdd FILL
XFILL_0__2362_ gnd vdd FILL
XFILL_5__3056_ gnd vdd FILL
X_2990_ _3023_/A _3092_/A _2990_/C _2999_/D vdd gnd OAI21X1
XFILL_3__2071_ gnd vdd FILL
XFILL_5__2007_ gnd vdd FILL
X_1941_ _1941_/A _1941_/B _1941_/C _2484_/A vdd gnd NAND3X1
XFILL_6__2820_ gnd vdd FILL
XFILL_8__1997_ gnd vdd FILL
XFILL_2__2229_ gnd vdd FILL
XFILL_0__2293_ gnd vdd FILL
X_1872_ _2913_/A _1875_/A _1872_/C _1878_/A vdd gnd OAI21X1
XFILL_6__2751_ gnd vdd FILL
XFILL_5__2909_ gnd vdd FILL
XFILL_3__2973_ gnd vdd FILL
XFILL_6__1702_ gnd vdd FILL
XFILL_6__2682_ gnd vdd FILL
X_3542_ _3570_/Q _3550_/A _3546_/C vdd gnd NAND2X1
XFILL_8__3598_ gnd vdd FILL
XFILL_8__2618_ gnd vdd FILL
XFILL_3__1924_ gnd vdd FILL
X_3473_ _3473_/A _3473_/B _3473_/C _3543_/B vdd gnd NAND3X1
XFILL_3__1855_ gnd vdd FILL
XFILL_8__2549_ gnd vdd FILL
X_2424_ _2872_/B _3077_/C _3254_/Q _2428_/A vdd gnd OAI21X1
X_2355_ _3173_/B _2966_/A _2448_/C _2356_/A vdd gnd OAI21X1
XFILL_3__1786_ gnd vdd FILL
XFILL_3__3525_ gnd vdd FILL
XFILL_3__3456_ gnd vdd FILL
X_2286_ _2286_/A _2286_/B _2286_/C _2287_/B vdd gnd NAND3X1
XFILL_1__2540_ gnd vdd FILL
XFILL_1__2471_ gnd vdd FILL
XFILL_6__3165_ gnd vdd FILL
XFILL_3__2407_ gnd vdd FILL
XFILL_4__2180_ gnd vdd FILL
XFILL_6__3096_ gnd vdd FILL
XFILL_3__3387_ gnd vdd FILL
XFILL_6__2116_ gnd vdd FILL
XFILL_0__2629_ gnd vdd FILL
XFILL_3__2338_ gnd vdd FILL
XFILL_6__2047_ gnd vdd FILL
XFILL_3__2269_ gnd vdd FILL
XFILL_7__2860_ gnd vdd FILL
XFILL_1__3023_ gnd vdd FILL
XFILL_7__2791_ gnd vdd FILL
XFILL_7__1811_ gnd vdd FILL
XFILL_6__2949_ gnd vdd FILL
XFILL_7__1742_ gnd vdd FILL
XFILL_4__1964_ gnd vdd FILL
XFILL_7__3412_ gnd vdd FILL
XFILL_5_CLKBUF1_insert29 gnd vdd FILL
XFILL_4__1895_ gnd vdd FILL
XFILL_1__2807_ gnd vdd FILL
XFILL_4__3565_ gnd vdd FILL
XFILL_4__3496_ gnd vdd FILL
XFILL_2__2580_ gnd vdd FILL
XFILL_4__2516_ gnd vdd FILL
XFILL_7__2225_ gnd vdd FILL
XFILL_3_CLKBUF1_insert33 gnd vdd FILL
XFILL_4__2447_ gnd vdd FILL
XFILL_1__2738_ gnd vdd FILL
XFILL_1_BUFX2_insert91 gnd vdd FILL
XFILL_1_BUFX2_insert80 gnd vdd FILL
XFILL_7__2156_ gnd vdd FILL
XFILL_1__2669_ gnd vdd FILL
XFILL_7__2087_ gnd vdd FILL
XFILL_4__2378_ gnd vdd FILL
XFILL_2__3201_ gnd vdd FILL
XFILL_2__3132_ gnd vdd FILL
XFILL_8__1920_ gnd vdd FILL
XFILL_8__1851_ gnd vdd FILL
XFILL_2__3063_ gnd vdd FILL
XFILL_2__2014_ gnd vdd FILL
XFILL_8__1782_ gnd vdd FILL
XFILL_7__2989_ gnd vdd FILL
XFILL_8__3521_ gnd vdd FILL
XFILL_8__3452_ gnd vdd FILL
XFILL_2__2916_ gnd vdd FILL
XFILL_8__3383_ gnd vdd FILL
XFILL_0__2980_ gnd vdd FILL
XFILL_8__2403_ gnd vdd FILL
XFILL_0__1931_ gnd vdd FILL
XFILL_8__2334_ gnd vdd FILL
XFILL_5__2625_ gnd vdd FILL
XFILL_2__2847_ gnd vdd FILL
XFILL_5__2556_ gnd vdd FILL
XFILL_0__1862_ gnd vdd FILL
XFILL_8__2265_ gnd vdd FILL
XFILL_0__3601_ gnd vdd FILL
XFILL_2__2778_ gnd vdd FILL
XFILL_8__2196_ gnd vdd FILL
X_2140_ _2342_/A _2433_/A _2140_/C _2332_/B vdd gnd OAI21X1
XFILL_5__2487_ gnd vdd FILL
XFILL_2__1729_ gnd vdd FILL
XFILL_0__1793_ gnd vdd FILL
XFILL_0__3532_ gnd vdd FILL
X_2071_ _2347_/A _2347_/B _2073_/B vdd gnd NAND2X1
XFILL_0__3463_ gnd vdd FILL
XFILL_5__3108_ gnd vdd FILL
XFILL_0__2414_ gnd vdd FILL
XFILL_3__3172_ gnd vdd FILL
XFILL_5__3039_ gnd vdd FILL
XFILL_0__3394_ gnd vdd FILL
XFILL_3__2123_ gnd vdd FILL
X_2973_ _2973_/A _2973_/B _2974_/B vdd gnd NAND2X1
XFILL_3__2054_ gnd vdd FILL
XFILL_0__2345_ gnd vdd FILL
XFILL_0__2276_ gnd vdd FILL
X_1924_ _2527_/C _1925_/C vdd gnd INVX1
XFILL_6__2803_ gnd vdd FILL
XFILL_9__3561_ gnd vdd FILL
X_1855_ _2966_/A _2966_/B _1862_/B _1856_/B vdd gnd OAI21X1
XFILL_6__2734_ gnd vdd FILL
XFILL_3__2956_ gnd vdd FILL
XFILL_9__2443_ gnd vdd FILL
X_1786_ _3160_/A _3160_/C _2199_/B vdd gnd NAND2X1
X_3525_ _3525_/A _3525_/B _3528_/B vdd gnd XOR2X1
XFILL_3__1907_ gnd vdd FILL
XFILL_1__1971_ gnd vdd FILL
XFILL_6__2665_ gnd vdd FILL
XFILL_3__2887_ gnd vdd FILL
XFILL_6__2596_ gnd vdd FILL
X_3456_ _3484_/B _3468_/B vdd gnd INVX1
XFILL_3__1838_ gnd vdd FILL
X_3387_ _3514_/B _3387_/B _3387_/C _3519_/B vdd gnd AOI21X1
XFILL_3__1769_ gnd vdd FILL
X_2407_ _2407_/A _3243_/Q _2407_/C _2411_/A vdd gnd AOI21X1
XFILL_3__3508_ gnd vdd FILL
XFILL_4__2301_ gnd vdd FILL
X_2338_ _2338_/A _2338_/B _2339_/A vdd gnd AND2X2
X_2269_ _2269_/A _2269_/B _2269_/C _2853_/A _2314_/A vdd gnd AOI22X1
XFILL_7__2010_ gnd vdd FILL
XFILL_6__3217_ gnd vdd FILL
XFILL_1__2523_ gnd vdd FILL
XFILL_3__3439_ gnd vdd FILL
XFILL_6__3148_ gnd vdd FILL
XFILL_4__2232_ gnd vdd FILL
XFILL_4__2163_ gnd vdd FILL
XFILL_1__2454_ gnd vdd FILL
XFILL_6__3079_ gnd vdd FILL
XFILL_1__2385_ gnd vdd FILL
XFILL_7__2912_ gnd vdd FILL
XFILL_4__2094_ gnd vdd FILL
XFILL_7__2843_ gnd vdd FILL
XFILL_1__3006_ gnd vdd FILL
XFILL_7__2774_ gnd vdd FILL
XFILL_4__2996_ gnd vdd FILL
XFILL_7__1725_ gnd vdd FILL
XFILL_4__1947_ gnd vdd FILL
XFILL_4__1878_ gnd vdd FILL
XFILL_2__2701_ gnd vdd FILL
XFILL_5__3390_ gnd vdd FILL
XFILL_5__2410_ gnd vdd FILL
XFILL_4__3548_ gnd vdd FILL
XFILL_5__2341_ gnd vdd FILL
XFILL_2__2632_ gnd vdd FILL
XFILL_8__2050_ gnd vdd FILL
XFILL_2__2563_ gnd vdd FILL
XFILL_4__3479_ gnd vdd FILL
XFILL_5__2272_ gnd vdd FILL
XFILL_7__2208_ gnd vdd FILL
XFILL_7__3188_ gnd vdd FILL
XFILL_7__2139_ gnd vdd FILL
XFILL_2__2494_ gnd vdd FILL
XFILL_6_BUFX2_insert26 gnd vdd FILL
XFILL_6_BUFX2_insert15 gnd vdd FILL
XFILL_6_BUFX2_insert59 gnd vdd FILL
XFILL_8__2952_ gnd vdd FILL
XFILL_6_BUFX2_insert48 gnd vdd FILL
XFILL_2__3115_ gnd vdd FILL
XFILL_8__1903_ gnd vdd FILL
XFILL_8__2883_ gnd vdd FILL
XFILL_0__2130_ gnd vdd FILL
XFILL_2__3046_ gnd vdd FILL
XFILL_8__1834_ gnd vdd FILL
XFILL_0__2061_ gnd vdd FILL
XFILL_8__1765_ gnd vdd FILL
XFILL_8__3504_ gnd vdd FILL
XFILL_3__2810_ gnd vdd FILL
XFILL_8__1696_ gnd vdd FILL
XFILL_5__1987_ gnd vdd FILL
XFILL_8__3435_ gnd vdd FILL
X_3310_ _3310_/D vdd _3313_/R _3578_/CLK _3310_/Q vdd gnd DFFSR
XFILL_6__2450_ gnd vdd FILL
XFILL_3__2741_ gnd vdd FILL
XFILL_0__2963_ gnd vdd FILL
XFILL_8__3366_ gnd vdd FILL
XFILL_3__2672_ gnd vdd FILL
XFILL_5__2608_ gnd vdd FILL
XFILL_0__2894_ gnd vdd FILL
XFILL_8__2317_ gnd vdd FILL
XFILL_6__2381_ gnd vdd FILL
XFILL_9__2090_ gnd vdd FILL
XFILL_0__1914_ gnd vdd FILL
XFILL_5__3588_ gnd vdd FILL
X_3241_ _3241_/D vdd _3291_/R _3355_/CLK _3241_/Q vdd gnd DFFSR
XFILL_8__2248_ gnd vdd FILL
XFILL_0__1845_ gnd vdd FILL
X_3172_ _3172_/A _3172_/B _3175_/B vdd gnd AND2X2
XFILL_5__2539_ gnd vdd FILL
XFILL184650x121050 gnd vdd FILL
X_2123_ _2123_/A _2123_/B _2958_/B vdd gnd NAND2X1
XFILL_0__3515_ gnd vdd FILL
XFILL_8__2179_ gnd vdd FILL
XFILL_6__3002_ gnd vdd FILL
XFILL_0__1776_ gnd vdd FILL
X_2054_ _2075_/A _2115_/B vdd gnd INVX1
XFILL_3__3224_ gnd vdd FILL
XFILL_0__3446_ gnd vdd FILL
XFILL_3__3155_ gnd vdd FILL
XFILL_9__1943_ gnd vdd FILL
XFILL_0__3377_ gnd vdd FILL
XFILL_1__2170_ gnd vdd FILL
XFILL_3__2106_ gnd vdd FILL
XFILL_3__3086_ gnd vdd FILL
XFILL_0__2328_ gnd vdd FILL
XFILL_3__2037_ gnd vdd FILL
X_2956_ _2993_/A _2956_/B _2956_/C _3306_/D vdd gnd OAI21X1
XFILL_4__2850_ gnd vdd FILL
X_2887_ _2887_/A _2887_/B _2892_/A vdd gnd NAND2X1
XFILL_0__2259_ gnd vdd FILL
X_1907_ _2701_/B _3152_/C _1907_/Y vdd gnd NAND2X1
X_1838_ _3192_/A _2199_/B _3088_/S _1861_/B vdd gnd NAND3X1
XFILL_4__1801_ gnd vdd FILL
XFILL_7__2490_ gnd vdd FILL
XFILL_4__2781_ gnd vdd FILL
XFILL_6__2717_ gnd vdd FILL
XFILL_3__2939_ gnd vdd FILL
X_1769_ _3281_/Q _1769_/B _3007_/C _1770_/B vdd gnd OAI21X1
XFILL_4__1732_ gnd vdd FILL
X_3508_ _3508_/A _3508_/B _3554_/B _3554_/A _3532_/B vdd gnd AOI22X1
XFILL_1__1954_ gnd vdd FILL
XFILL_6__2648_ gnd vdd FILL
XFILL_6__2579_ gnd vdd FILL
XFILL_4__3402_ gnd vdd FILL
X_3439_ _3468_/S _3439_/B _3449_/A _3440_/B vdd gnd OAI21X1
XFILL_1__1885_ gnd vdd FILL
XFILL_7__3111_ gnd vdd FILL
XFILL_7__3042_ gnd vdd FILL
XFILL_1__3555_ gnd vdd FILL
XFILL_1__3486_ gnd vdd FILL
XFILL_4__2215_ gnd vdd FILL
XFILL_1__2506_ gnd vdd FILL
XFILL_4__3195_ gnd vdd FILL
XFILL_1__2437_ gnd vdd FILL
XFILL_4__2146_ gnd vdd FILL
XFILL_4__2077_ gnd vdd FILL
XFILL_1__2368_ gnd vdd FILL
XFILL_1__2299_ gnd vdd FILL
XFILL_5__1910_ gnd vdd FILL
XFILL_5__2890_ gnd vdd FILL
XFILL_7__2826_ gnd vdd FILL
XFILL_7__2757_ gnd vdd FILL
XFILL_5__1841_ gnd vdd FILL
XFILL_4__2979_ gnd vdd FILL
XFILL_5__1772_ gnd vdd FILL
XFILL_7__1708_ gnd vdd FILL
XFILL_5__3511_ gnd vdd FILL
XFILL_2__1994_ gnd vdd FILL
XFILL_7__2688_ gnd vdd FILL
XFILL_5__3442_ gnd vdd FILL
XFILL_8__3220_ gnd vdd FILL
XFILL_8__3151_ gnd vdd FILL
XFILL_8__3082_ gnd vdd FILL
XFILL_5__3373_ gnd vdd FILL
XFILL_8__2102_ gnd vdd FILL
XFILL_2__2615_ gnd vdd FILL
XFILL_8__2033_ gnd vdd FILL
XFILL_5__2324_ gnd vdd FILL
XFILL_2__3595_ gnd vdd FILL
XFILL_5__2255_ gnd vdd FILL
XFILL_2__2546_ gnd vdd FILL
XFILL_2__2477_ gnd vdd FILL
XFILL_5__2186_ gnd vdd FILL
XFILL_0__3231_ gnd vdd FILL
XFILL_8__2935_ gnd vdd FILL
XFILL_8__2866_ gnd vdd FILL
XFILL_6__1950_ gnd vdd FILL
X_2810_ _3266_/Q _2980_/A vdd gnd INVX1
XFILL_0__3162_ gnd vdd FILL
XFILL_2__3029_ gnd vdd FILL
XFILL_0__3093_ gnd vdd FILL
XFILL_6__1881_ gnd vdd FILL
XFILL_0__2113_ gnd vdd FILL
X_2741_ _2741_/A _2741_/B _2741_/C _2775_/C vdd gnd NOR3X1
XFILL_8__1817_ gnd vdd FILL
XFILL_0__2044_ gnd vdd FILL
XFILL_8__2797_ gnd vdd FILL
XFILL_6__3551_ gnd vdd FILL
XFILL_8__1748_ gnd vdd FILL
X_2672_ _2674_/B _2673_/A vdd gnd INVX1
XFILL_6__2502_ gnd vdd FILL
XFILL_6__3482_ gnd vdd FILL
XFILL_8__3418_ gnd vdd FILL
XFILL_2_BUFX2_insert24 gnd vdd FILL
XFILL_3__2724_ gnd vdd FILL
XFILL_2_BUFX2_insert13 gnd vdd FILL
XFILL_2_BUFX2_insert57 gnd vdd FILL
XFILL_0__2946_ gnd vdd FILL
XFILL_2_BUFX2_insert79 gnd vdd FILL
XFILL_2_BUFX2_insert68 gnd vdd FILL
XFILL_2_BUFX2_insert46 gnd vdd FILL
XFILL_6__2433_ gnd vdd FILL
XFILL_6__2364_ gnd vdd FILL
X_3224_ _3224_/A _3230_/B _3224_/C _3359_/D vdd gnd OAI21X1
XFILL_3__2655_ gnd vdd FILL
.ends

