magic
tech scmos
magscale 1 3
timestamp 1725342160
<< nwell >>
rect 0 0 270 270
<< diffusion >>
rect 41 231 229 249
rect 21 41 39 229
rect 87 87 183 183
rect 231 41 249 229
rect 41 21 229 39
<< psubstratepdiff >>
rect 85 183 185 185
rect 85 87 87 183
rect 183 87 185 183
rect 85 85 185 87
<< nsubstratendiff >>
rect 20 249 250 250
rect 20 231 41 249
rect 229 231 250 249
rect 20 230 250 231
rect 20 229 40 230
rect 20 41 21 229
rect 39 41 40 229
rect 230 229 250 230
rect 20 40 40 41
rect 230 41 231 229
rect 249 41 250 229
rect 230 40 250 41
rect 20 39 250 40
rect 20 21 41 39
rect 229 21 250 39
rect 20 20 250 21
<< metal1 >>
rect 20 230 250 250
rect 20 40 40 230
rect 85 85 185 185
rect 230 40 250 230
rect 20 20 250 40
<< end >>
