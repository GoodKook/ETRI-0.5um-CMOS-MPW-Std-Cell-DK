/* Verilog module written by vlogFanout (qflow) */
/* With clock tree generation and fanout reduction */
/* and gate resizing */

module fir_pe(
    input [5:0] Cin,
    input Rdy,
    output Vld,
    input [3:0] Xin,
    output [3:0] Xout,
    input [3:0] Yin,
    output [3:0] Yout,
    input clk
);

wire [15:0] y ;
wire _588_ ;
wire _168_ ;
wire _60_ ;
wire _397_ ;
wire _703_ ;
wire _19_ ;
wire _512_ ;
wire [4:0] LoadCtl ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire _453_ ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire _54_ ;
wire _603_ ;
wire _412_ ;
wire _92_ ;
wire _641_ ;
wire _221_ ;
wire _450_ ;
wire _506_ ;
wire _735_ ;
wire _315_ ;
wire _544_ ;
wire _124_ ;
wire _353_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire _391_ ;
wire _447_ ;
wire _676_ ;
wire _256_ ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire _600_ ;
wire Rdy ;
wire _197_ ;
wire _7_ ;
wire _503_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _541_ ;
wire _121_ ;
wire _350_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire _444_ ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire [7:0] XinHL ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire _45_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _441_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _535_ ;
wire _115_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire _438_ ;
wire _191_ ;
wire _667_ ;
wire _247_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire clk_bF$buf5 ;
wire clk_bF$buf6 ;
wire clk_bF$buf7 ;
wire _285_ ;
wire _1_ ;
wire _42_ ;
wire _379_ ;
wire _188_ ;
wire _400_ ;
wire _80_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire _341_ ;
wire clk ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire [3:0] _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _376_ ;
wire _185_ ;
wire _699_ ;
wire _279_ ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire _74_ ;
wire _623_ ;
wire _203_ ;
wire _432_ ;
wire _661_ ;
wire _241_ ;
wire Cin_1_bF$buf0 ;
wire Cin_1_bF$buf1 ;
wire Cin_1_bF$buf2 ;
wire Cin_1_bF$buf3 ;
wire _717_ ;
wire _470_ ;
wire _526_ ;
wire _106_ ;
wire _755_ ;
wire _335_ ;
wire _564_ ;
wire _144_ ;
wire _373_ ;
wire _429_ ;
wire _182_ ;
wire LoadCtl_0_bF$buf0 ;
wire LoadCtl_0_bF$buf1 ;
wire LoadCtl_0_bF$buf2 ;
wire LoadCtl_0_bF$buf3 ;
wire LoadCtl_0_bF$buf4 ;
wire _658_ ;
wire _238_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _71_ ;
wire _620_ ;
wire _200_ ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire _617_ ;
wire _370_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _464_ ;
wire _693_ ;
wire _273_ ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _367_ ;
wire _596_ ;
wire _176_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire _65_ ;
wire _614_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _461_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire _555_ ;
wire _135_ ;
wire _364_ ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire _458_ ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire _24_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire _420_ ;
wire _705_ ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _361_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _646_ ;
wire _226_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _358_ ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire _702_ ;
wire _299_ ;
wire _18_ ;
wire _511_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire _605_ ;
wire _414_ ;
wire _94_ ;
wire _643_ ;
wire _223_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire _355_ ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _449_ ;
wire _678_ ;
wire _258_ ;
wire _487_ ;
wire _296_ ;
wire _15_ ;
wire _53_ ;
wire _602_ ;
wire _199_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _505_ ;
wire _734_ ;
wire _314_ ;
wire _543_ ;
wire _123_ ;
wire _352_ ;
wire _408_ ;
wire _88_ ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _446_ ;
wire [3:0] Yin ;
wire _675_ ;
wire _255_ ;
wire _484_ ;
wire _293_ ;
wire _12_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire _405_ ;
wire _85_ ;
wire [3:0] Yin0 ;
wire [3:0] Yin1 ;
wire [3:0] Yin2 ;
wire [3:0] Yin3 ;
wire _634_ ;
wire _214_ ;
wire _443_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _346_ ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire _478_ ;
wire _287_ ;
wire _3_ ;
wire _44_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _440_ ;
wire _725_ ;
wire _305_ ;
wire [3:0] XinH ;
wire _534_ ;
wire _114_ ;
wire _343_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire _475_ ;
wire _284_ ;
wire _0_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _378_ ;
wire _187_ ;
wire [3:0] Yout ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire _340_ ;
wire _76_ ;
wire _625_ ;
wire _205_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire _375_ ;
wire _184_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _35_ ;
wire [3:0] Xout ;
wire _73_ ;
wire _622_ ;
wire _202_ ;
wire _431_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire _619_ ;
wire _372_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire _32_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _70_ ;
wire LoadCtl_4_bF$buf0 ;
wire LoadCtl_4_bF$buf1 ;
wire LoadCtl_4_bF$buf2 ;
wire LoadCtl_4_bF$buf3 ;
wire LoadCtl_4_bF$buf4 ;
wire LoadCtl_4_bF$buf5 ;
wire LoadCtl_4_bF$buf6 ;
wire LoadCtl_4_bF$buf7 ;
wire _713_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire _751_ ;
wire _331_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire _616_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire _463_ ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire _366_ ;
wire _595_ ;
wire _175_ ;
wire _689_ ;
wire _269_ ;
wire _498_ ;
wire _710_ ;
wire _26_ ;
wire Cin_0_bF$buf0 ;
wire Cin_0_bF$buf1 ;
wire Cin_0_bF$buf2 ;
wire Cin_0_bF$buf3 ;
wire _64_ ;
wire _613_ ;
wire _422_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _460_ ;
wire _516_ ;
wire _745_ ;
wire _325_ ;
wire _554_ ;
wire _134_ ;
wire _363_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire Vld ;
wire _648_ ;
wire _228_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire _495_ ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire _61_ ;
wire _398_ ;
wire _610_ ;
wire _704_ ;
wire _513_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _360_ ;
wire _416_ ;
wire _96_ ;
wire [5:0] Cin ;
wire _645_ ;
wire _225_ ;
wire _454_ ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire _489_ ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire _55_ ;
wire _604_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _736_ ;
wire _316_ ;
wire _545_ ;
wire _125_ ;
wire _354_ ;
wire _583_ ;
wire _163_ ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _448_ ;
wire _677_ ;
wire _257_ ;
wire _486_ ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire _351_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _470__bF$buf0 ;
wire _470__bF$buf1 ;
wire _470__bF$buf2 ;
wire _470__bF$buf3 ;
wire _470__bF$buf4 ;
wire _636_ ;
wire _216_ ;
wire _445_ ;
wire _674_ ;
wire _254_ ;
wire _483_ ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _442_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _536_ ;
wire _116_ ;
wire _345_ ;
wire _574_ ;
wire _154_ ;
wire _383_ ;
wire _439_ ;
wire _192_ ;
wire _668_ ;
wire _248_ ;
wire _477_ ;
wire _286_ ;
wire _2_ ;
wire _43_ ;
wire _189_ ;
wire _401_ ;
wire _81_ ;
wire _630_ ;
wire _210_ ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire _342_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _436_ ;
wire [3:0] Xin ;
wire _665_ ;
wire _245_ ;
wire _474_ ;
wire _283_ ;
wire [3:0] _759_ ;
wire _339_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _377_ ;
wire _186_ ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire _75_ ;
wire _624_ ;
wire _204_ ;
wire _433_ ;
wire [13:0] mul ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _374_ ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire _34_ ;
wire _72_ ;
wire _621_ ;
wire _201_ ;
wire _430_ ;
wire _715_ ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _371_ ;
wire [15:0] rYin ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _368_ ;
wire _597_ ;
wire _177_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire _66_ ;
wire _615_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _462_ ;
wire _518_ ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire _556_ ;
wire _136_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire _459_ ;
wire _688_ ;
wire _268_ ;
wire _497_ ;
wire _25_ ;
wire _63_ ;
wire _612_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _362_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _456_ ;
wire _685_ ;
wire _265_ ;
wire _494_ ;
wire _22_ ;
wire _359_ ;

BUFX2 BUFX2_insert33 (
    .A(Cin[1]),
    .Y(Cin_1_bF$buf0)
);

BUFX2 BUFX2_insert32 (
    .A(Cin[1]),
    .Y(Cin_1_bF$buf1)
);

BUFX2 BUFX2_insert31 (
    .A(Cin[1]),
    .Y(Cin_1_bF$buf2)
);

BUFX2 BUFX2_insert30 (
    .A(Cin[1]),
    .Y(Cin_1_bF$buf3)
);

BUFX2 BUFX2_insert29 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf0)
);

BUFX2 BUFX2_insert28 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf1)
);

BUFX2 BUFX2_insert27 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf2)
);

BUFX2 BUFX2_insert26 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf3)
);

BUFX2 BUFX2_insert25 (
    .A(LoadCtl[0]),
    .Y(LoadCtl_0_bF$buf4)
);

BUFX2 BUFX2_insert24 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf0)
);

BUFX2 BUFX2_insert23 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf1)
);

BUFX2 BUFX2_insert22 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf2)
);

BUFX2 BUFX2_insert21 (
    .A(Cin[0]),
    .Y(Cin_0_bF$buf3)
);

BUFX2 BUFX2_insert20 (
    .A(_470_),
    .Y(_470__bF$buf0)
);

BUFX2 BUFX2_insert19 (
    .A(_470_),
    .Y(_470__bF$buf1)
);

BUFX2 BUFX2_insert18 (
    .A(_470_),
    .Y(_470__bF$buf2)
);

BUFX2 BUFX2_insert17 (
    .A(_470_),
    .Y(_470__bF$buf3)
);

BUFX2 BUFX2_insert16 (
    .A(_470_),
    .Y(_470__bF$buf4)
);

CLKBUF1 CLKBUF1_insert15 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert14 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert13 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert12 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert11 (
    .A(clk),
    .Y(clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert10 (
    .A(clk),
    .Y(clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert9 (
    .A(clk),
    .Y(clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert8 (
    .A(clk),
    .Y(clk_bF$buf7)
);

BUFX2 BUFX2_insert7 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf0)
);

BUFX2 BUFX2_insert6 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf1)
);

BUFX2 BUFX2_insert5 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf2)
);

BUFX2 BUFX2_insert4 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf3)
);

BUFX2 BUFX2_insert3 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf4)
);

BUFX2 BUFX2_insert2 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf5)
);

BUFX2 BUFX2_insert1 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf6)
);

BUFX2 BUFX2_insert0 (
    .A(LoadCtl[4]),
    .Y(LoadCtl_4_bF$buf7)
);

NAND2X1 _1000_ (
    .A(_221_),
    .B(_228_),
    .Y(_277_)
);

OR2X2 _1001_ (
    .A(_277_),
    .B(_276_),
    .Y(_278_)
);

AOI22X1 _1002_ (
    .A(_272_),
    .B(_275_),
    .C(_221_),
    .D(_228_),
    .Y(_279_)
);

INVX1 _1003_ (
    .A(_279_),
    .Y(_280_)
);

NAND3X1 _1004_ (
    .A(LoadCtl_4_bF$buf7),
    .B(_280_),
    .C(_278_),
    .Y(_281_)
);

OAI21X1 _1005_ (
    .A(_230_),
    .B(LoadCtl_4_bF$buf6),
    .C(_281_),
    .Y(_25_)
);

INVX1 _1006_ (
    .A(mul[6]),
    .Y(_282_)
);

AOI21X1 _1007_ (
    .A(_263_),
    .B(_267_),
    .C(_269_),
    .Y(_283_)
);

OAI21X1 _1008_ (
    .A(_232_),
    .B(_283_),
    .C(_273_),
    .Y(_284_)
);

NAND2X1 _1009_ (
    .A(XinHL[2]),
    .B(Cin[4]),
    .Y(_285_)
);

OAI21X1 _1010_ (
    .A(_213_),
    .B(_285_),
    .C(_245_),
    .Y(_286_)
);

INVX1 _1011_ (
    .A(_286_),
    .Y(_287_)
);

INVX1 _1012_ (
    .A(_265_),
    .Y(_288_)
);

AOI21X1 _1013_ (
    .A(_264_),
    .B(_266_),
    .C(_288_),
    .Y(_289_)
);

NAND2X1 _1014_ (
    .A(XinHL[1]),
    .B(Cin[5]),
    .Y(_290_)
);

AND2X2 _1015_ (
    .A(XinHL[3]),
    .B(Cin[3]),
    .Y(_291_)
);

OAI21X1 _1016_ (
    .A(_176_),
    .B(_212_),
    .C(_291_),
    .Y(_292_)
);

AND2X2 _1017_ (
    .A(XinHL[2]),
    .B(Cin[4]),
    .Y(_293_)
);

OAI21X1 _1018_ (
    .A(_178_),
    .B(_239_),
    .C(_293_),
    .Y(_294_)
);

NAND3X1 _1019_ (
    .A(_290_),
    .B(_292_),
    .C(_294_),
    .Y(_295_)
);

INVX1 _1020_ (
    .A(_290_),
    .Y(_296_)
);

NAND2X1 _1021_ (
    .A(_293_),
    .B(_291_),
    .Y(_297_)
);

OAI21X1 _1022_ (
    .A(_178_),
    .B(_239_),
    .C(_285_),
    .Y(_298_)
);

NAND3X1 _1023_ (
    .A(_298_),
    .B(_296_),
    .C(_297_),
    .Y(_299_)
);

NAND2X1 _1024_ (
    .A(_299_),
    .B(_295_),
    .Y(_300_)
);

NOR2X1 _1025_ (
    .A(_203_),
    .B(_251_),
    .Y(_301_)
);

AOI21X1 _1026_ (
    .A(_254_),
    .B(_256_),
    .C(_301_),
    .Y(_302_)
);

NAND2X1 _1027_ (
    .A(XinH[0]),
    .B(Cin[2]),
    .Y(_303_)
);

AND2X2 _1028_ (
    .A(XinH[2]),
    .B(Cin_0_bF$buf3),
    .Y(_304_)
);

OAI21X1 _1029_ (
    .A(_91_),
    .B(_141_),
    .C(_304_),
    .Y(_305_)
);

NAND2X1 _1030_ (
    .A(XinH[2]),
    .B(Cin_0_bF$buf2),
    .Y(_306_)
);

NAND3X1 _1031_ (
    .A(XinH[1]),
    .B(Cin_1_bF$buf3),
    .C(_306_),
    .Y(_307_)
);

NAND3X1 _1032_ (
    .A(_303_),
    .B(_307_),
    .C(_305_),
    .Y(_308_)
);

INVX1 _1033_ (
    .A(_303_),
    .Y(_309_)
);

AND2X2 _1034_ (
    .A(XinH[2]),
    .B(Cin_1_bF$buf2),
    .Y(_310_)
);

NAND2X1 _1035_ (
    .A(_249_),
    .B(_310_),
    .Y(_311_)
);

OAI21X1 _1036_ (
    .A(_91_),
    .B(_141_),
    .C(_306_),
    .Y(_312_)
);

NAND3X1 _1037_ (
    .A(_312_),
    .B(_309_),
    .C(_311_),
    .Y(_313_)
);

NAND3X1 _1038_ (
    .A(_308_),
    .B(_313_),
    .C(_302_),
    .Y(_314_)
);

AOI22X1 _1039_ (
    .A(XinH[0]),
    .B(Cin_1_bF$buf1),
    .C(XinH[1]),
    .D(Cin_0_bF$buf1),
    .Y(_315_)
);

OAI21X1 _1040_ (
    .A(_248_),
    .B(_315_),
    .C(_255_),
    .Y(_316_)
);

AOI21X1 _1041_ (
    .A(_311_),
    .B(_312_),
    .C(_309_),
    .Y(_317_)
);

AOI21X1 _1042_ (
    .A(_305_),
    .B(_307_),
    .C(_303_),
    .Y(_318_)
);

OAI21X1 _1043_ (
    .A(_317_),
    .B(_318_),
    .C(_316_),
    .Y(_319_)
);

NAND3X1 _1044_ (
    .A(_300_),
    .B(_314_),
    .C(_319_),
    .Y(_320_)
);

AND2X2 _1045_ (
    .A(_295_),
    .B(_299_),
    .Y(_321_)
);

NAND3X1 _1046_ (
    .A(_316_),
    .B(_313_),
    .C(_308_),
    .Y(_322_)
);

OAI21X1 _1047_ (
    .A(_317_),
    .B(_318_),
    .C(_302_),
    .Y(_323_)
);

NAND3X1 _1048_ (
    .A(_322_),
    .B(_321_),
    .C(_323_),
    .Y(_324_)
);

NAND3X1 _1049_ (
    .A(_320_),
    .B(_324_),
    .C(_289_),
    .Y(_325_)
);

AOI21X1 _1050_ (
    .A(_253_),
    .B(_257_),
    .C(_259_),
    .Y(_326_)
);

OAI21X1 _1051_ (
    .A(_246_),
    .B(_326_),
    .C(_265_),
    .Y(_327_)
);

AOI21X1 _1052_ (
    .A(_323_),
    .B(_322_),
    .C(_321_),
    .Y(_328_)
);

AOI21X1 _1053_ (
    .A(_319_),
    .B(_314_),
    .C(_300_),
    .Y(_329_)
);

OAI21X1 _1054_ (
    .A(_328_),
    .B(_329_),
    .C(_327_),
    .Y(_330_)
);

NAND3X1 _1055_ (
    .A(_287_),
    .B(_330_),
    .C(_325_),
    .Y(_331_)
);

NAND3X1 _1056_ (
    .A(_320_),
    .B(_324_),
    .C(_327_),
    .Y(_332_)
);

OAI21X1 _1057_ (
    .A(_328_),
    .B(_329_),
    .C(_289_),
    .Y(_333_)
);

NAND3X1 _1058_ (
    .A(_286_),
    .B(_332_),
    .C(_333_),
    .Y(_334_)
);

NAND3X1 _1059_ (
    .A(_334_),
    .B(_284_),
    .C(_331_),
    .Y(_335_)
);

INVX1 _1060_ (
    .A(_273_),
    .Y(_336_)
);

AOI21X1 _1061_ (
    .A(_233_),
    .B(_274_),
    .C(_336_),
    .Y(_337_)
);

AOI21X1 _1062_ (
    .A(_333_),
    .B(_332_),
    .C(_286_),
    .Y(_338_)
);

AOI21X1 _1063_ (
    .A(_325_),
    .B(_330_),
    .C(_287_),
    .Y(_339_)
);

OAI21X1 _1064_ (
    .A(_338_),
    .B(_339_),
    .C(_337_),
    .Y(_340_)
);

AND2X2 _1065_ (
    .A(_340_),
    .B(_335_),
    .Y(_341_)
);

NOR2X1 _1066_ (
    .A(_279_),
    .B(_341_),
    .Y(_342_)
);

INVX1 _1067_ (
    .A(_341_),
    .Y(_343_)
);

OAI21X1 _1068_ (
    .A(_280_),
    .B(_343_),
    .C(LoadCtl_4_bF$buf5),
    .Y(_344_)
);

OAI22X1 _1069_ (
    .A(_282_),
    .B(LoadCtl_4_bF$buf4),
    .C(_342_),
    .D(_344_),
    .Y(_26_)
);

INVX1 _1070_ (
    .A(mul[7]),
    .Y(_345_)
);

NAND3X1 _1071_ (
    .A(_335_),
    .B(_279_),
    .C(_340_),
    .Y(_346_)
);

AOI21X1 _1072_ (
    .A(_324_),
    .B(_320_),
    .C(_327_),
    .Y(_347_)
);

OAI21X1 _1073_ (
    .A(_287_),
    .B(_347_),
    .C(_332_),
    .Y(_348_)
);

NAND2X1 _1074_ (
    .A(_297_),
    .B(_299_),
    .Y(_349_)
);

AOI21X1 _1075_ (
    .A(_308_),
    .B(_313_),
    .C(_316_),
    .Y(_350_)
);

OAI21X1 _1076_ (
    .A(_300_),
    .B(_350_),
    .C(_322_),
    .Y(_351_)
);

NAND2X1 _1077_ (
    .A(XinHL[2]),
    .B(Cin[5]),
    .Y(_352_)
);

AND2X2 _1078_ (
    .A(XinH[0]),
    .B(Cin[3]),
    .Y(_353_)
);

OAI21X1 _1079_ (
    .A(_178_),
    .B(_212_),
    .C(_353_),
    .Y(_354_)
);

AND2X2 _1080_ (
    .A(XinHL[3]),
    .B(Cin[4]),
    .Y(_355_)
);

OAI21X1 _1081_ (
    .A(_89_),
    .B(_239_),
    .C(_355_),
    .Y(_356_)
);

NAND3X1 _1082_ (
    .A(_352_),
    .B(_354_),
    .C(_356_),
    .Y(_357_)
);

INVX1 _1083_ (
    .A(_352_),
    .Y(_358_)
);

NAND2X1 _1084_ (
    .A(_355_),
    .B(_353_),
    .Y(_359_)
);

NAND2X1 _1085_ (
    .A(XinH[0]),
    .B(Cin[3]),
    .Y(_360_)
);

OAI21X1 _1086_ (
    .A(_178_),
    .B(_212_),
    .C(_360_),
    .Y(_361_)
);

NAND3X1 _1087_ (
    .A(_361_),
    .B(_358_),
    .C(_359_),
    .Y(_362_)
);

NAND2X1 _1088_ (
    .A(_362_),
    .B(_357_),
    .Y(_363_)
);

AOI22X1 _1089_ (
    .A(_249_),
    .B(_310_),
    .C(_312_),
    .D(_309_),
    .Y(_364_)
);

NAND2X1 _1090_ (
    .A(XinH[1]),
    .B(Cin[2]),
    .Y(_365_)
);

AND2X2 _1091_ (
    .A(XinH[3]),
    .B(Cin_0_bF$buf0),
    .Y(_366_)
);

OAI21X1 _1092_ (
    .A(_93_),
    .B(_141_),
    .C(_366_),
    .Y(_367_)
);

OAI21X1 _1093_ (
    .A(_95_),
    .B(_179_),
    .C(_310_),
    .Y(_368_)
);

NAND3X1 _1094_ (
    .A(_365_),
    .B(_367_),
    .C(_368_),
    .Y(_369_)
);

INVX1 _1095_ (
    .A(_365_),
    .Y(_370_)
);

NAND2X1 _1096_ (
    .A(_310_),
    .B(_366_),
    .Y(_371_)
);

AOI22X1 _1097_ (
    .A(XinH[2]),
    .B(Cin_1_bF$buf0),
    .C(XinH[3]),
    .D(Cin_0_bF$buf3),
    .Y(_372_)
);

INVX1 _1098_ (
    .A(_372_),
    .Y(_373_)
);

NAND3X1 _1099_ (
    .A(_370_),
    .B(_373_),
    .C(_371_),
    .Y(_374_)
);

NAND3X1 _1100_ (
    .A(_374_),
    .B(_364_),
    .C(_369_),
    .Y(_375_)
);

AOI22X1 _1101_ (
    .A(XinH[1]),
    .B(Cin_1_bF$buf3),
    .C(XinH[2]),
    .D(Cin_0_bF$buf2),
    .Y(_376_)
);

OAI21X1 _1102_ (
    .A(_303_),
    .B(_376_),
    .C(_311_),
    .Y(_377_)
);

AOI21X1 _1103_ (
    .A(_371_),
    .B(_373_),
    .C(_370_),
    .Y(_378_)
);

AOI21X1 _1104_ (
    .A(_367_),
    .B(_368_),
    .C(_365_),
    .Y(_379_)
);

OAI21X1 _1105_ (
    .A(_378_),
    .B(_379_),
    .C(_377_),
    .Y(_380_)
);

NAND3X1 _1106_ (
    .A(_363_),
    .B(_375_),
    .C(_380_),
    .Y(_381_)
);

AND2X2 _1107_ (
    .A(_357_),
    .B(_362_),
    .Y(_382_)
);

NAND3X1 _1108_ (
    .A(_377_),
    .B(_374_),
    .C(_369_),
    .Y(_383_)
);

OAI21X1 _1109_ (
    .A(_378_),
    .B(_379_),
    .C(_364_),
    .Y(_384_)
);

NAND3X1 _1110_ (
    .A(_383_),
    .B(_382_),
    .C(_384_),
    .Y(_385_)
);

NAND3X1 _1111_ (
    .A(_351_),
    .B(_381_),
    .C(_385_),
    .Y(_386_)
);

INVX1 _1112_ (
    .A(_322_),
    .Y(_387_)
);

AOI21X1 _1113_ (
    .A(_321_),
    .B(_323_),
    .C(_387_),
    .Y(_388_)
);

AOI21X1 _1114_ (
    .A(_384_),
    .B(_383_),
    .C(_382_),
    .Y(_389_)
);

AOI21X1 _1115_ (
    .A(_380_),
    .B(_375_),
    .C(_363_),
    .Y(_390_)
);

OAI21X1 _1116_ (
    .A(_389_),
    .B(_390_),
    .C(_388_),
    .Y(_391_)
);

NAND3X1 _1117_ (
    .A(_349_),
    .B(_386_),
    .C(_391_),
    .Y(_392_)
);

INVX1 _1118_ (
    .A(_349_),
    .Y(_393_)
);

NAND3X1 _1119_ (
    .A(_381_),
    .B(_385_),
    .C(_388_),
    .Y(_394_)
);

OAI21X1 _1120_ (
    .A(_389_),
    .B(_390_),
    .C(_351_),
    .Y(_395_)
);

NAND3X1 _1121_ (
    .A(_393_),
    .B(_395_),
    .C(_394_),
    .Y(_396_)
);

AOI21X1 _1122_ (
    .A(_396_),
    .B(_392_),
    .C(_348_),
    .Y(_397_)
);

NAND3X1 _1123_ (
    .A(_349_),
    .B(_395_),
    .C(_394_),
    .Y(_398_)
);

NAND3X1 _1124_ (
    .A(_393_),
    .B(_386_),
    .C(_391_),
    .Y(_399_)
);

AOI22X1 _1125_ (
    .A(_334_),
    .B(_332_),
    .C(_398_),
    .D(_399_),
    .Y(_400_)
);

NOR2X1 _1126_ (
    .A(_397_),
    .B(_400_),
    .Y(_401_)
);

AOI21X1 _1127_ (
    .A(_346_),
    .B(_335_),
    .C(_401_),
    .Y(_402_)
);

OAI21X1 _1128_ (
    .A(_280_),
    .B(_343_),
    .C(_335_),
    .Y(_403_)
);

INVX1 _1129_ (
    .A(_348_),
    .Y(_404_)
);

NAND3X1 _1130_ (
    .A(_398_),
    .B(_399_),
    .C(_404_),
    .Y(_405_)
);

NAND3X1 _1131_ (
    .A(_348_),
    .B(_392_),
    .C(_396_),
    .Y(_406_)
);

NAND2X1 _1132_ (
    .A(_406_),
    .B(_405_),
    .Y(_407_)
);

NOR2X1 _1133_ (
    .A(_407_),
    .B(_403_),
    .Y(_408_)
);

OAI21X1 _1134_ (
    .A(_402_),
    .B(_408_),
    .C(LoadCtl_4_bF$buf3),
    .Y(_409_)
);

OAI21X1 _1135_ (
    .A(_345_),
    .B(LoadCtl_4_bF$buf2),
    .C(_409_),
    .Y(_27_)
);

INVX1 _1136_ (
    .A(mul[8]),
    .Y(_410_)
);

NAND2X1 _1137_ (
    .A(_406_),
    .B(_335_),
    .Y(_411_)
);

NAND2X1 _1138_ (
    .A(_405_),
    .B(_411_),
    .Y(_412_)
);

OAI21X1 _1139_ (
    .A(_407_),
    .B(_346_),
    .C(_412_),
    .Y(_413_)
);

AOI21X1 _1140_ (
    .A(_381_),
    .B(_385_),
    .C(_351_),
    .Y(_414_)
);

OAI21X1 _1141_ (
    .A(_393_),
    .B(_414_),
    .C(_386_),
    .Y(_415_)
);

NAND2X1 _1142_ (
    .A(_359_),
    .B(_362_),
    .Y(_416_)
);

INVX1 _1143_ (
    .A(_416_),
    .Y(_417_)
);

INVX1 _1144_ (
    .A(_383_),
    .Y(_418_)
);

AOI21X1 _1145_ (
    .A(_382_),
    .B(_384_),
    .C(_418_),
    .Y(_419_)
);

INVX2 _1146_ (
    .A(Cin[5]),
    .Y(_420_)
);

NOR2X1 _1147_ (
    .A(_178_),
    .B(_420_),
    .Y(_421_)
);

AND2X2 _1148_ (
    .A(XinH[1]),
    .B(Cin[3]),
    .Y(_422_)
);

NAND3X1 _1149_ (
    .A(XinH[0]),
    .B(Cin[4]),
    .C(_422_),
    .Y(_423_)
);

AOI22X1 _1150_ (
    .A(XinH[0]),
    .B(Cin[4]),
    .C(XinH[1]),
    .D(Cin[3]),
    .Y(_424_)
);

INVX1 _1151_ (
    .A(_424_),
    .Y(_425_)
);

NAND3X1 _1152_ (
    .A(_425_),
    .B(_421_),
    .C(_423_),
    .Y(_426_)
);

NAND2X1 _1153_ (
    .A(XinH[1]),
    .B(Cin[4]),
    .Y(_427_)
);

NOR2X1 _1154_ (
    .A(_360_),
    .B(_427_),
    .Y(_428_)
);

OAI22X1 _1155_ (
    .A(_178_),
    .B(_420_),
    .C(_424_),
    .D(_428_),
    .Y(_429_)
);

NAND2X1 _1156_ (
    .A(_426_),
    .B(_429_),
    .Y(_430_)
);

AND2X2 _1157_ (
    .A(XinH[3]),
    .B(Cin_1_bF$buf2),
    .Y(_431_)
);

AOI22X1 _1158_ (
    .A(_304_),
    .B(_431_),
    .C(_373_),
    .D(_370_),
    .Y(_432_)
);

NAND2X1 _1159_ (
    .A(XinH[2]),
    .B(Cin_1_bF$buf1),
    .Y(_433_)
);

NAND2X1 _1160_ (
    .A(XinH[3]),
    .B(Cin[2]),
    .Y(_434_)
);

AOI22X1 _1161_ (
    .A(XinH[2]),
    .B(Cin[2]),
    .C(XinH[3]),
    .D(Cin_1_bF$buf0),
    .Y(_435_)
);

INVX1 _1162_ (
    .A(_435_),
    .Y(_436_)
);

OAI21X1 _1163_ (
    .A(_433_),
    .B(_434_),
    .C(_436_),
    .Y(_437_)
);

NOR2X1 _1164_ (
    .A(_437_),
    .B(_432_),
    .Y(_438_)
);

OAI21X1 _1165_ (
    .A(_365_),
    .B(_372_),
    .C(_371_),
    .Y(_439_)
);

INVX1 _1166_ (
    .A(_434_),
    .Y(_440_)
);

AOI21X1 _1167_ (
    .A(_440_),
    .B(_310_),
    .C(_435_),
    .Y(_441_)
);

NOR2X1 _1168_ (
    .A(_441_),
    .B(_439_),
    .Y(_442_)
);

OAI21X1 _1169_ (
    .A(_442_),
    .B(_438_),
    .C(_430_),
    .Y(_443_)
);

AND2X2 _1170_ (
    .A(_429_),
    .B(_426_),
    .Y(_444_)
);

NAND2X1 _1171_ (
    .A(_441_),
    .B(_432_),
    .Y(_445_)
);

NAND2X1 _1172_ (
    .A(_437_),
    .B(_439_),
    .Y(_446_)
);

NAND2X1 _1173_ (
    .A(_446_),
    .B(_445_),
    .Y(_447_)
);

NAND2X1 _1174_ (
    .A(_444_),
    .B(_447_),
    .Y(_448_)
);

NAND3X1 _1175_ (
    .A(_443_),
    .B(_448_),
    .C(_419_),
    .Y(_449_)
);

AOI21X1 _1176_ (
    .A(_369_),
    .B(_374_),
    .C(_377_),
    .Y(_450_)
);

OAI21X1 _1177_ (
    .A(_363_),
    .B(_450_),
    .C(_383_),
    .Y(_451_)
);

NOR2X1 _1178_ (
    .A(_444_),
    .B(_447_),
    .Y(_452_)
);

AOI21X1 _1179_ (
    .A(_445_),
    .B(_446_),
    .C(_430_),
    .Y(_453_)
);

OAI21X1 _1180_ (
    .A(_453_),
    .B(_452_),
    .C(_451_),
    .Y(_454_)
);

NAND3X1 _1181_ (
    .A(_417_),
    .B(_449_),
    .C(_454_),
    .Y(_455_)
);

NAND3X1 _1182_ (
    .A(_451_),
    .B(_443_),
    .C(_448_),
    .Y(_456_)
);

OAI21X1 _1183_ (
    .A(_453_),
    .B(_452_),
    .C(_419_),
    .Y(_457_)
);

NAND3X1 _1184_ (
    .A(_416_),
    .B(_456_),
    .C(_457_),
    .Y(_458_)
);

NAND3X1 _1185_ (
    .A(_415_),
    .B(_458_),
    .C(_455_),
    .Y(_459_)
);

INVX1 _1186_ (
    .A(_415_),
    .Y(_460_)
);

AOI21X1 _1187_ (
    .A(_457_),
    .B(_456_),
    .C(_416_),
    .Y(_461_)
);

AOI21X1 _1188_ (
    .A(_454_),
    .B(_449_),
    .C(_417_),
    .Y(_462_)
);

OAI21X1 _1189_ (
    .A(_461_),
    .B(_462_),
    .C(_460_),
    .Y(_463_)
);

NAND2X1 _1190_ (
    .A(_459_),
    .B(_463_),
    .Y(_464_)
);

INVX1 _1191_ (
    .A(_464_),
    .Y(_465_)
);

NOR2X1 _1192_ (
    .A(_465_),
    .B(_413_),
    .Y(_466_)
);

INVX1 _1193_ (
    .A(_413_),
    .Y(_467_)
);

OAI21X1 _1194_ (
    .A(_464_),
    .B(_467_),
    .C(LoadCtl_4_bF$buf1),
    .Y(_468_)
);

OAI22X1 _1195_ (
    .A(_410_),
    .B(LoadCtl_4_bF$buf0),
    .C(_466_),
    .D(_468_),
    .Y(_28_)
);

INVX1 _1196_ (
    .A(mul[9]),
    .Y(_469_)
);

INVX8 _1197_ (
    .A(LoadCtl_4_bF$buf7),
    .Y(_470_)
);

INVX1 _1198_ (
    .A(_459_),
    .Y(_471_)
);

AOI21X1 _1199_ (
    .A(_413_),
    .B(_465_),
    .C(_471_),
    .Y(_472_)
);

AOI21X1 _1200_ (
    .A(_448_),
    .B(_443_),
    .C(_451_),
    .Y(_473_)
);

OAI21X1 _1201_ (
    .A(_417_),
    .B(_473_),
    .C(_456_),
    .Y(_474_)
);

AOI21X1 _1202_ (
    .A(_421_),
    .B(_425_),
    .C(_428_),
    .Y(_475_)
);

INVX1 _1203_ (
    .A(_475_),
    .Y(_476_)
);

NAND2X1 _1204_ (
    .A(_441_),
    .B(_439_),
    .Y(_477_)
);

OAI21X1 _1205_ (
    .A(_430_),
    .B(_442_),
    .C(_477_),
    .Y(_478_)
);

NOR2X1 _1206_ (
    .A(_89_),
    .B(_420_),
    .Y(_479_)
);

NAND2X1 _1207_ (
    .A(XinH[2]),
    .B(Cin[4]),
    .Y(_480_)
);

INVX1 _1208_ (
    .A(_480_),
    .Y(_481_)
);

NAND2X1 _1209_ (
    .A(_422_),
    .B(_481_),
    .Y(_482_)
);

OAI21X1 _1210_ (
    .A(_93_),
    .B(_239_),
    .C(_427_),
    .Y(_483_)
);

NAND3X1 _1211_ (
    .A(_483_),
    .B(_479_),
    .C(_482_),
    .Y(_484_)
);

NAND2X1 _1212_ (
    .A(XinH[1]),
    .B(Cin[3]),
    .Y(_485_)
);

OAI21X1 _1213_ (
    .A(_485_),
    .B(_480_),
    .C(_483_),
    .Y(_486_)
);

OAI21X1 _1214_ (
    .A(_89_),
    .B(_420_),
    .C(_486_),
    .Y(_487_)
);

NAND2X1 _1215_ (
    .A(_484_),
    .B(_487_),
    .Y(_488_)
);

OAI21X1 _1216_ (
    .A(_310_),
    .B(_434_),
    .C(_488_),
    .Y(_489_)
);

OAI21X1 _1217_ (
    .A(_93_),
    .B(_141_),
    .C(_440_),
    .Y(_490_)
);

INVX1 _1218_ (
    .A(_490_),
    .Y(_491_)
);

NAND3X1 _1219_ (
    .A(_484_),
    .B(_491_),
    .C(_487_),
    .Y(_492_)
);

NAND3X1 _1220_ (
    .A(_478_),
    .B(_492_),
    .C(_489_),
    .Y(_493_)
);

NAND2X1 _1221_ (
    .A(_437_),
    .B(_432_),
    .Y(_494_)
);

AOI21X1 _1222_ (
    .A(_444_),
    .B(_494_),
    .C(_438_),
    .Y(_495_)
);

AOI21X1 _1223_ (
    .A(_487_),
    .B(_484_),
    .C(_491_),
    .Y(_496_)
);

INVX1 _1224_ (
    .A(_492_),
    .Y(_497_)
);

OAI21X1 _1225_ (
    .A(_496_),
    .B(_497_),
    .C(_495_),
    .Y(_498_)
);

NAND3X1 _1226_ (
    .A(_476_),
    .B(_493_),
    .C(_498_),
    .Y(_499_)
);

NAND3X1 _1227_ (
    .A(_489_),
    .B(_492_),
    .C(_495_),
    .Y(_500_)
);

OAI21X1 _1228_ (
    .A(_496_),
    .B(_497_),
    .C(_478_),
    .Y(_501_)
);

NAND3X1 _1229_ (
    .A(_475_),
    .B(_501_),
    .C(_500_),
    .Y(_502_)
);

AOI21X1 _1230_ (
    .A(_499_),
    .B(_502_),
    .C(_474_),
    .Y(_503_)
);

NAND3X1 _1231_ (
    .A(_476_),
    .B(_501_),
    .C(_500_),
    .Y(_504_)
);

NAND3X1 _1232_ (
    .A(_475_),
    .B(_493_),
    .C(_498_),
    .Y(_505_)
);

AOI22X1 _1233_ (
    .A(_504_),
    .B(_505_),
    .C(_458_),
    .D(_456_),
    .Y(_506_)
);

NOR2X1 _1234_ (
    .A(_503_),
    .B(_506_),
    .Y(_507_)
);

OR2X2 _1235_ (
    .A(_472_),
    .B(_507_),
    .Y(_508_)
);

AOI21X1 _1236_ (
    .A(_472_),
    .B(_507_),
    .C(_470__bF$buf4),
    .Y(_509_)
);

AOI22X1 _1237_ (
    .A(_469_),
    .B(_470__bF$buf3),
    .C(_508_),
    .D(_509_),
    .Y(_29_)
);

INVX1 _1238_ (
    .A(mul[10]),
    .Y(_510_)
);

NAND2X1 _1239_ (
    .A(_499_),
    .B(_502_),
    .Y(_511_)
);

NAND3X1 _1240_ (
    .A(_456_),
    .B(_458_),
    .C(_511_),
    .Y(_512_)
);

NAND3X1 _1241_ (
    .A(_499_),
    .B(_502_),
    .C(_474_),
    .Y(_513_)
);

NAND2X1 _1242_ (
    .A(_513_),
    .B(_512_),
    .Y(_514_)
);

NOR2X1 _1243_ (
    .A(_514_),
    .B(_464_),
    .Y(_515_)
);

OAI21X1 _1244_ (
    .A(_459_),
    .B(_503_),
    .C(_513_),
    .Y(_516_)
);

AOI21X1 _1245_ (
    .A(_413_),
    .B(_515_),
    .C(_516_),
    .Y(_517_)
);

NAND2X1 _1246_ (
    .A(_493_),
    .B(_499_),
    .Y(_518_)
);

OAI21X1 _1247_ (
    .A(_485_),
    .B(_480_),
    .C(_484_),
    .Y(_519_)
);

INVX1 _1248_ (
    .A(_519_),
    .Y(_520_)
);

NAND2X1 _1249_ (
    .A(_310_),
    .B(_440_),
    .Y(_521_)
);

NAND2X1 _1250_ (
    .A(XinH[1]),
    .B(Cin[5]),
    .Y(_522_)
);

NAND2X1 _1251_ (
    .A(XinH[2]),
    .B(Cin[3]),
    .Y(_523_)
);

OAI21X1 _1252_ (
    .A(_95_),
    .B(_239_),
    .C(_480_),
    .Y(_524_)
);

NAND2X1 _1253_ (
    .A(XinH[3]),
    .B(Cin[4]),
    .Y(_525_)
);

OAI21X1 _1254_ (
    .A(_523_),
    .B(_525_),
    .C(_524_),
    .Y(_526_)
);

OR2X2 _1255_ (
    .A(_526_),
    .B(_522_),
    .Y(_527_)
);

OAI21X1 _1256_ (
    .A(_91_),
    .B(_420_),
    .C(_526_),
    .Y(_528_)
);

NAND2X1 _1257_ (
    .A(_528_),
    .B(_527_),
    .Y(_529_)
);

AOI21X1 _1258_ (
    .A(_521_),
    .B(_492_),
    .C(_529_),
    .Y(_530_)
);

NAND3X1 _1259_ (
    .A(_521_),
    .B(_492_),
    .C(_529_),
    .Y(_531_)
);

INVX1 _1260_ (
    .A(_531_),
    .Y(_532_)
);

OAI21X1 _1261_ (
    .A(_530_),
    .B(_532_),
    .C(_520_),
    .Y(_533_)
);

INVX1 _1262_ (
    .A(_530_),
    .Y(_534_)
);

NAND3X1 _1263_ (
    .A(_519_),
    .B(_531_),
    .C(_534_),
    .Y(_535_)
);

NAND3X1 _1264_ (
    .A(_533_),
    .B(_535_),
    .C(_518_),
    .Y(_536_)
);

NAND2X1 _1265_ (
    .A(_533_),
    .B(_535_),
    .Y(_537_)
);

NAND3X1 _1266_ (
    .A(_493_),
    .B(_499_),
    .C(_537_),
    .Y(_538_)
);

NAND2X1 _1267_ (
    .A(_536_),
    .B(_538_),
    .Y(_539_)
);

NAND2X1 _1268_ (
    .A(_539_),
    .B(_517_),
    .Y(_540_)
);

NAND3X1 _1269_ (
    .A(_279_),
    .B(_401_),
    .C(_341_),
    .Y(_541_)
);

NAND3X1 _1270_ (
    .A(_459_),
    .B(_463_),
    .C(_507_),
    .Y(_542_)
);

AOI21X1 _1271_ (
    .A(_541_),
    .B(_412_),
    .C(_542_),
    .Y(_543_)
);

INVX1 _1272_ (
    .A(_539_),
    .Y(_544_)
);

OAI21X1 _1273_ (
    .A(_516_),
    .B(_543_),
    .C(_544_),
    .Y(_545_)
);

NAND3X1 _1274_ (
    .A(LoadCtl_4_bF$buf6),
    .B(_540_),
    .C(_545_),
    .Y(_546_)
);

OAI21X1 _1275_ (
    .A(_510_),
    .B(LoadCtl_4_bF$buf5),
    .C(_546_),
    .Y(_30_)
);

NAND2X1 _1276_ (
    .A(mul[11]),
    .B(_470__bF$buf2),
    .Y(_547_)
);

AOI21X1 _1277_ (
    .A(_519_),
    .B(_531_),
    .C(_530_),
    .Y(_548_)
);

OAI21X1 _1278_ (
    .A(_523_),
    .B(_525_),
    .C(_527_),
    .Y(_549_)
);

OAI21X1 _1279_ (
    .A(_93_),
    .B(_420_),
    .C(_525_),
    .Y(_550_)
);

NOR2X1 _1280_ (
    .A(_95_),
    .B(_420_),
    .Y(_551_)
);

NAND2X1 _1281_ (
    .A(_481_),
    .B(_551_),
    .Y(_552_)
);

AND2X2 _1282_ (
    .A(_552_),
    .B(_550_),
    .Y(_553_)
);

OR2X2 _1283_ (
    .A(_549_),
    .B(_553_),
    .Y(_554_)
);

NAND2X1 _1284_ (
    .A(_553_),
    .B(_549_),
    .Y(_555_)
);

NAND2X1 _1285_ (
    .A(_555_),
    .B(_554_),
    .Y(_556_)
);

NOR2X1 _1286_ (
    .A(_548_),
    .B(_556_),
    .Y(_557_)
);

AND2X2 _1287_ (
    .A(_556_),
    .B(_548_),
    .Y(_558_)
);

NOR2X1 _1288_ (
    .A(_557_),
    .B(_558_),
    .Y(_559_)
);

INVX1 _1289_ (
    .A(_559_),
    .Y(_560_)
);

NAND3X1 _1290_ (
    .A(_536_),
    .B(_560_),
    .C(_545_),
    .Y(_561_)
);

OAI21X1 _1291_ (
    .A(_539_),
    .B(_517_),
    .C(_536_),
    .Y(_562_)
);

NAND2X1 _1292_ (
    .A(_559_),
    .B(_562_),
    .Y(_563_)
);

NAND3X1 _1293_ (
    .A(LoadCtl_4_bF$buf4),
    .B(_563_),
    .C(_561_),
    .Y(_564_)
);

NAND2X1 _1294_ (
    .A(_547_),
    .B(_564_),
    .Y(_31_)
);

INVX1 _1295_ (
    .A(mul[12]),
    .Y(_565_)
);

NAND3X1 _1296_ (
    .A(_536_),
    .B(_538_),
    .C(_559_),
    .Y(_566_)
);

NOR2X1 _1297_ (
    .A(_566_),
    .B(_542_),
    .Y(_567_)
);

INVX1 _1298_ (
    .A(_516_),
    .Y(_568_)
);

NOR2X1 _1299_ (
    .A(_558_),
    .B(_536_),
    .Y(_569_)
);

NOR2X1 _1300_ (
    .A(_557_),
    .B(_569_),
    .Y(_570_)
);

OAI21X1 _1301_ (
    .A(_566_),
    .B(_568_),
    .C(_570_),
    .Y(_571_)
);

AOI21X1 _1302_ (
    .A(_567_),
    .B(_413_),
    .C(_571_),
    .Y(_572_)
);

INVX1 _1303_ (
    .A(_555_),
    .Y(_573_)
);

NAND3X1 _1304_ (
    .A(_551_),
    .B(_552_),
    .C(_573_),
    .Y(_574_)
);

INVX1 _1305_ (
    .A(_551_),
    .Y(_575_)
);

OAI21X1 _1306_ (
    .A(_481_),
    .B(_575_),
    .C(_555_),
    .Y(_576_)
);

NAND2X1 _1307_ (
    .A(_576_),
    .B(_574_),
    .Y(_577_)
);

NAND2X1 _1308_ (
    .A(_577_),
    .B(_572_),
    .Y(_578_)
);

INVX1 _1309_ (
    .A(_578_),
    .Y(_579_)
);

OAI21X1 _1310_ (
    .A(_577_),
    .B(_572_),
    .C(LoadCtl_4_bF$buf3),
    .Y(_580_)
);

OAI22X1 _1311_ (
    .A(_565_),
    .B(LoadCtl_4_bF$buf2),
    .C(_580_),
    .D(_579_),
    .Y(_32_)
);

INVX1 _1312_ (
    .A(mul[13]),
    .Y(_581_)
);

OR2X2 _1313_ (
    .A(_572_),
    .B(_577_),
    .Y(_582_)
);

INVX1 _1314_ (
    .A(_574_),
    .Y(_583_)
);

OAI21X1 _1315_ (
    .A(_480_),
    .B(_575_),
    .C(LoadCtl_4_bF$buf1),
    .Y(_584_)
);

NOR2X1 _1316_ (
    .A(_584_),
    .B(_583_),
    .Y(_585_)
);

AOI22X1 _1317_ (
    .A(_581_),
    .B(_470__bF$buf1),
    .C(_582_),
    .D(_585_),
    .Y(_33_)
);

NOR2X1 _1318_ (
    .A(_101_),
    .B(_133_),
    .Y(_586_)
);

INVX1 _1319_ (
    .A(_586_),
    .Y(_587_)
);

NAND2X1 _1320_ (
    .A(_101_),
    .B(_133_),
    .Y(_588_)
);

NAND2X1 _1321_ (
    .A(_588_),
    .B(_587_),
    .Y(_589_)
);

NAND2X1 _1322_ (
    .A(y[0]),
    .B(_470__bF$buf0),
    .Y(_590_)
);

OAI21X1 _1323_ (
    .A(_470__bF$buf4),
    .B(_589_),
    .C(_590_),
    .Y(_34_)
);

NOR2X1 _1324_ (
    .A(_103_),
    .B(_135_),
    .Y(_591_)
);

NOR2X1 _1325_ (
    .A(rYin[1]),
    .B(mul[1]),
    .Y(_592_)
);

NOR2X1 _1326_ (
    .A(_592_),
    .B(_591_),
    .Y(_593_)
);

NAND2X1 _1327_ (
    .A(_586_),
    .B(_593_),
    .Y(_594_)
);

OAI21X1 _1328_ (
    .A(_591_),
    .B(_592_),
    .C(_587_),
    .Y(_595_)
);

NAND2X1 _1329_ (
    .A(_595_),
    .B(_594_),
    .Y(_596_)
);

NAND2X1 _1330_ (
    .A(y[1]),
    .B(_470__bF$buf3),
    .Y(_597_)
);

OAI21X1 _1331_ (
    .A(_470__bF$buf2),
    .B(_596_),
    .C(_597_),
    .Y(_35_)
);

OAI21X1 _1332_ (
    .A(_103_),
    .B(_135_),
    .C(_594_),
    .Y(_598_)
);

NOR2X1 _1333_ (
    .A(rYin[2]),
    .B(mul[2]),
    .Y(_599_)
);

NOR2X1 _1334_ (
    .A(_105_),
    .B(_144_),
    .Y(_600_)
);

NOR2X1 _1335_ (
    .A(_599_),
    .B(_600_),
    .Y(_601_)
);

NAND2X1 _1336_ (
    .A(_601_),
    .B(_598_),
    .Y(_602_)
);

OR2X2 _1337_ (
    .A(_598_),
    .B(_601_),
    .Y(_603_)
);

NAND2X1 _1338_ (
    .A(_602_),
    .B(_603_),
    .Y(_604_)
);

NAND2X1 _1339_ (
    .A(y[2]),
    .B(_470__bF$buf1),
    .Y(_605_)
);

OAI21X1 _1340_ (
    .A(_470__bF$buf0),
    .B(_604_),
    .C(_605_),
    .Y(_36_)
);

AOI21X1 _1341_ (
    .A(_598_),
    .B(_601_),
    .C(_600_),
    .Y(_606_)
);

NOR2X1 _1342_ (
    .A(rYin[3]),
    .B(mul[3]),
    .Y(_607_)
);

NOR2X1 _1343_ (
    .A(_107_),
    .B(_160_),
    .Y(_608_)
);

OAI21X1 _1344_ (
    .A(_607_),
    .B(_608_),
    .C(_606_),
    .Y(_609_)
);

INVX1 _1345_ (
    .A(_606_),
    .Y(_610_)
);

INVX1 _1346_ (
    .A(_607_),
    .Y(_611_)
);

INVX1 _1347_ (
    .A(_608_),
    .Y(_612_)
);

NAND3X1 _1348_ (
    .A(_611_),
    .B(_612_),
    .C(_610_),
    .Y(_613_)
);

NAND2X1 _1349_ (
    .A(_609_),
    .B(_613_),
    .Y(_614_)
);

NAND2X1 _1350_ (
    .A(y[3]),
    .B(_470__bF$buf4),
    .Y(_615_)
);

OAI21X1 _1351_ (
    .A(_470__bF$buf3),
    .B(_614_),
    .C(_615_),
    .Y(_37_)
);

NAND2X1 _1352_ (
    .A(y[4]),
    .B(_470__bF$buf2),
    .Y(_616_)
);

NOR2X1 _1353_ (
    .A(rYin[4]),
    .B(mul[4]),
    .Y(_617_)
);

NOR2X1 _1354_ (
    .A(_109_),
    .B(_191_),
    .Y(_618_)
);

OAI21X1 _1355_ (
    .A(_607_),
    .B(_606_),
    .C(_612_),
    .Y(_619_)
);

INVX1 _1356_ (
    .A(_619_),
    .Y(_620_)
);

OAI21X1 _1357_ (
    .A(_617_),
    .B(_618_),
    .C(_620_),
    .Y(_621_)
);

NOR2X1 _1358_ (
    .A(_617_),
    .B(_618_),
    .Y(_622_)
);

NAND2X1 _1359_ (
    .A(_622_),
    .B(_619_),
    .Y(_623_)
);

NAND2X1 _1360_ (
    .A(_623_),
    .B(_621_),
    .Y(_624_)
);

OAI21X1 _1361_ (
    .A(_470__bF$buf1),
    .B(_624_),
    .C(_616_),
    .Y(_38_)
);

INVX1 _1362_ (
    .A(y[5]),
    .Y(_625_)
);

AOI21X1 _1363_ (
    .A(_619_),
    .B(_622_),
    .C(_618_),
    .Y(_626_)
);

NOR2X1 _1364_ (
    .A(rYin[5]),
    .B(mul[5]),
    .Y(_627_)
);

NOR2X1 _1365_ (
    .A(_111_),
    .B(_230_),
    .Y(_628_)
);

NOR2X1 _1366_ (
    .A(_627_),
    .B(_628_),
    .Y(_629_)
);

AND2X2 _1367_ (
    .A(_626_),
    .B(_629_),
    .Y(_630_)
);

NOR2X1 _1368_ (
    .A(_629_),
    .B(_626_),
    .Y(_631_)
);

OAI21X1 _1369_ (
    .A(_631_),
    .B(_630_),
    .C(LoadCtl_4_bF$buf0),
    .Y(_632_)
);

OAI21X1 _1370_ (
    .A(_625_),
    .B(LoadCtl_4_bF$buf7),
    .C(_632_),
    .Y(_39_)
);

NAND2X1 _1371_ (
    .A(y[6]),
    .B(_470__bF$buf0),
    .Y(_633_)
);

NAND2X1 _1372_ (
    .A(_618_),
    .B(_629_),
    .Y(_634_)
);

OAI21X1 _1373_ (
    .A(_111_),
    .B(_230_),
    .C(_634_),
    .Y(_635_)
);

AND2X2 _1374_ (
    .A(_622_),
    .B(_629_),
    .Y(_636_)
);

AOI21X1 _1375_ (
    .A(_619_),
    .B(_636_),
    .C(_635_),
    .Y(_637_)
);

NOR2X1 _1376_ (
    .A(rYin[6]),
    .B(mul[6]),
    .Y(_638_)
);

NOR2X1 _1377_ (
    .A(_113_),
    .B(_282_),
    .Y(_639_)
);

NOR2X1 _1378_ (
    .A(_638_),
    .B(_639_),
    .Y(_640_)
);

INVX1 _1379_ (
    .A(_640_),
    .Y(_641_)
);

AND2X2 _1380_ (
    .A(_637_),
    .B(_641_),
    .Y(_642_)
);

OAI21X1 _1381_ (
    .A(_641_),
    .B(_637_),
    .C(LoadCtl_4_bF$buf6),
    .Y(_643_)
);

OAI21X1 _1382_ (
    .A(_643_),
    .B(_642_),
    .C(_633_),
    .Y(_40_)
);

INVX1 _1383_ (
    .A(_639_),
    .Y(_644_)
);

OAI21X1 _1384_ (
    .A(_638_),
    .B(_637_),
    .C(_644_),
    .Y(_645_)
);

NOR2X1 _1385_ (
    .A(rYin[7]),
    .B(mul[7]),
    .Y(_646_)
);

NOR2X1 _1386_ (
    .A(_115_),
    .B(_345_),
    .Y(_647_)
);

NOR2X1 _1387_ (
    .A(_646_),
    .B(_647_),
    .Y(_648_)
);

OR2X2 _1388_ (
    .A(_645_),
    .B(_648_),
    .Y(_649_)
);

NAND2X1 _1389_ (
    .A(_648_),
    .B(_645_),
    .Y(_650_)
);

NAND2X1 _1390_ (
    .A(_650_),
    .B(_649_),
    .Y(_651_)
);

NAND2X1 _1391_ (
    .A(y[7]),
    .B(_470__bF$buf4),
    .Y(_652_)
);

OAI21X1 _1392_ (
    .A(_470__bF$buf3),
    .B(_651_),
    .C(_652_),
    .Y(_41_)
);

NAND2X1 _1393_ (
    .A(y[8]),
    .B(_470__bF$buf2),
    .Y(_653_)
);

INVX1 _1394_ (
    .A(_647_),
    .Y(_654_)
);

OAI21X1 _1395_ (
    .A(_646_),
    .B(_644_),
    .C(_654_),
    .Y(_655_)
);

AND2X2 _1396_ (
    .A(_640_),
    .B(_648_),
    .Y(_656_)
);

AOI21X1 _1397_ (
    .A(_635_),
    .B(_656_),
    .C(_655_),
    .Y(_657_)
);

NAND3X1 _1398_ (
    .A(_636_),
    .B(_656_),
    .C(_619_),
    .Y(_658_)
);

AND2X2 _1399_ (
    .A(_658_),
    .B(_657_),
    .Y(_659_)
);

INVX1 _1400_ (
    .A(_659_),
    .Y(_660_)
);

NOR2X1 _1401_ (
    .A(rYin[8]),
    .B(mul[8]),
    .Y(_661_)
);

NOR2X1 _1402_ (
    .A(_117_),
    .B(_410_),
    .Y(_662_)
);

NOR2X1 _1403_ (
    .A(_661_),
    .B(_662_),
    .Y(_663_)
);

NOR2X1 _1404_ (
    .A(_663_),
    .B(_660_),
    .Y(_664_)
);

INVX1 _1405_ (
    .A(_663_),
    .Y(_665_)
);

OAI21X1 _1406_ (
    .A(_665_),
    .B(_659_),
    .C(LoadCtl_4_bF$buf5),
    .Y(_666_)
);

OAI21X1 _1407_ (
    .A(_666_),
    .B(_664_),
    .C(_653_),
    .Y(_42_)
);

AOI21X1 _1408_ (
    .A(_660_),
    .B(_663_),
    .C(_662_),
    .Y(_667_)
);

NOR2X1 _1409_ (
    .A(rYin[9]),
    .B(mul[9]),
    .Y(_668_)
);

NOR2X1 _1410_ (
    .A(_119_),
    .B(_469_),
    .Y(_669_)
);

NOR2X1 _1411_ (
    .A(_668_),
    .B(_669_),
    .Y(_670_)
);

AND2X2 _1412_ (
    .A(_667_),
    .B(_670_),
    .Y(_671_)
);

NOR2X1 _1413_ (
    .A(_670_),
    .B(_667_),
    .Y(_672_)
);

OAI21X1 _1414_ (
    .A(_672_),
    .B(_671_),
    .C(LoadCtl_4_bF$buf4),
    .Y(_673_)
);

OAI21X1 _1415_ (
    .A(_78_),
    .B(LoadCtl_4_bF$buf3),
    .C(_673_),
    .Y(_43_)
);

NAND2X1 _1416_ (
    .A(y[10]),
    .B(_470__bF$buf1),
    .Y(_674_)
);

AND2X2 _1417_ (
    .A(_663_),
    .B(_670_),
    .Y(_675_)
);

OAI21X1 _1418_ (
    .A(rYin[9]),
    .B(mul[9]),
    .C(_662_),
    .Y(_676_)
);

OAI21X1 _1419_ (
    .A(_119_),
    .B(_469_),
    .C(_676_),
    .Y(_677_)
);

AOI21X1 _1420_ (
    .A(_660_),
    .B(_675_),
    .C(_677_),
    .Y(_678_)
);

NOR2X1 _1421_ (
    .A(rYin[10]),
    .B(mul[10]),
    .Y(_679_)
);

NOR2X1 _1422_ (
    .A(_121_),
    .B(_510_),
    .Y(_680_)
);

NOR2X1 _1423_ (
    .A(_679_),
    .B(_680_),
    .Y(_681_)
);

INVX1 _1424_ (
    .A(_681_),
    .Y(_682_)
);

AND2X2 _1425_ (
    .A(_678_),
    .B(_682_),
    .Y(_683_)
);

OAI21X1 _1426_ (
    .A(_682_),
    .B(_678_),
    .C(LoadCtl_4_bF$buf2),
    .Y(_684_)
);

OAI21X1 _1427_ (
    .A(_684_),
    .B(_683_),
    .C(_674_),
    .Y(_44_)
);

INVX1 _1428_ (
    .A(_680_),
    .Y(_685_)
);

OAI21X1 _1429_ (
    .A(_679_),
    .B(_678_),
    .C(_685_),
    .Y(_686_)
);

NOR2X1 _1430_ (
    .A(rYin[11]),
    .B(mul[11]),
    .Y(_687_)
);

NAND2X1 _1431_ (
    .A(rYin[11]),
    .B(mul[11]),
    .Y(_688_)
);

INVX1 _1432_ (
    .A(_688_),
    .Y(_689_)
);

NOR2X1 _1433_ (
    .A(_687_),
    .B(_689_),
    .Y(_690_)
);

INVX1 _1434_ (
    .A(_690_),
    .Y(_691_)
);

OR2X2 _1435_ (
    .A(_686_),
    .B(_691_),
    .Y(_692_)
);

AOI21X1 _1436_ (
    .A(_686_),
    .B(_691_),
    .C(_470__bF$buf0),
    .Y(_693_)
);

AOI22X1 _1437_ (
    .A(_85_),
    .B(_470__bF$buf4),
    .C(_692_),
    .D(_693_),
    .Y(_45_)
);

NAND2X1 _1438_ (
    .A(y[12]),
    .B(_470__bF$buf3),
    .Y(_694_)
);

AOI21X1 _1439_ (
    .A(_690_),
    .B(_680_),
    .C(_689_),
    .Y(_695_)
);

NOR2X1 _1440_ (
    .A(_691_),
    .B(_682_),
    .Y(_696_)
);

NAND2X1 _1441_ (
    .A(_677_),
    .B(_696_),
    .Y(_697_)
);

NAND2X1 _1442_ (
    .A(_695_),
    .B(_697_),
    .Y(_698_)
);

NAND2X1 _1443_ (
    .A(_675_),
    .B(_696_),
    .Y(_699_)
);

NOR2X1 _1444_ (
    .A(_699_),
    .B(_659_),
    .Y(_700_)
);

OR2X2 _1445_ (
    .A(_700_),
    .B(_698_),
    .Y(_701_)
);

NOR2X1 _1446_ (
    .A(rYin[12]),
    .B(mul[12]),
    .Y(_702_)
);

NOR2X1 _1447_ (
    .A(_125_),
    .B(_565_),
    .Y(_703_)
);

NOR2X1 _1448_ (
    .A(_702_),
    .B(_703_),
    .Y(_704_)
);

NOR2X1 _1449_ (
    .A(_704_),
    .B(_701_),
    .Y(_705_)
);

NOR2X1 _1450_ (
    .A(_698_),
    .B(_700_),
    .Y(_706_)
);

INVX1 _1451_ (
    .A(_704_),
    .Y(_707_)
);

OAI21X1 _1452_ (
    .A(_707_),
    .B(_706_),
    .C(LoadCtl_4_bF$buf1),
    .Y(_708_)
);

OAI21X1 _1453_ (
    .A(_708_),
    .B(_705_),
    .C(_694_),
    .Y(_46_)
);

INVX1 _1454_ (
    .A(y[13]),
    .Y(_709_)
);

INVX1 _1455_ (
    .A(_703_),
    .Y(_710_)
);

OAI21X1 _1456_ (
    .A(_702_),
    .B(_706_),
    .C(_710_),
    .Y(_711_)
);

NOR2X1 _1457_ (
    .A(rYin[13]),
    .B(mul[13]),
    .Y(_712_)
);

NOR2X1 _1458_ (
    .A(_127_),
    .B(_581_),
    .Y(_713_)
);

NOR2X1 _1459_ (
    .A(_712_),
    .B(_713_),
    .Y(_714_)
);

INVX1 _1460_ (
    .A(_714_),
    .Y(_715_)
);

OR2X2 _1461_ (
    .A(_711_),
    .B(_715_),
    .Y(_716_)
);

AOI21X1 _1462_ (
    .A(_711_),
    .B(_715_),
    .C(_470__bF$buf2),
    .Y(_717_)
);

AOI22X1 _1463_ (
    .A(_709_),
    .B(_470__bF$buf1),
    .C(_716_),
    .D(_717_),
    .Y(_47_)
);

NAND2X1 _1464_ (
    .A(y[14]),
    .B(_470__bF$buf0),
    .Y(_718_)
);

AOI21X1 _1465_ (
    .A(_714_),
    .B(_703_),
    .C(_713_),
    .Y(_719_)
);

NOR2X1 _1466_ (
    .A(_707_),
    .B(_715_),
    .Y(_720_)
);

INVX1 _1467_ (
    .A(_720_),
    .Y(_721_)
);

OAI21X1 _1468_ (
    .A(_721_),
    .B(_706_),
    .C(_719_),
    .Y(_722_)
);

NOR2X1 _1469_ (
    .A(rYin[14]),
    .B(_722_),
    .Y(_723_)
);

INVX1 _1470_ (
    .A(_719_),
    .Y(_724_)
);

AOI21X1 _1471_ (
    .A(_701_),
    .B(_720_),
    .C(_724_),
    .Y(_725_)
);

OAI21X1 _1472_ (
    .A(_129_),
    .B(_725_),
    .C(LoadCtl_4_bF$buf0),
    .Y(_726_)
);

OAI21X1 _1473_ (
    .A(_723_),
    .B(_726_),
    .C(_718_),
    .Y(_48_)
);

NAND2X1 _1474_ (
    .A(y[15]),
    .B(_470__bF$buf4),
    .Y(_727_)
);

NAND3X1 _1475_ (
    .A(rYin[14]),
    .B(rYin[15]),
    .C(_722_),
    .Y(_728_)
);

OAI21X1 _1476_ (
    .A(_129_),
    .B(_725_),
    .C(_131_),
    .Y(_729_)
);

NAND2X1 _1477_ (
    .A(_728_),
    .B(_729_),
    .Y(_730_)
);

OAI21X1 _1478_ (
    .A(_470__bF$buf3),
    .B(_730_),
    .C(_727_),
    .Y(_49_)
);

INVX1 _1479_ (
    .A(Yin[0]),
    .Y(_731_)
);

NAND3X1 _1480_ (
    .A(LoadCtl[3]),
    .B(_71_),
    .C(_72_),
    .Y(_732_)
);

NAND2X1 _1481_ (
    .A(Yin3[0]),
    .B(_732_),
    .Y(_733_)
);

OAI21X1 _1482_ (
    .A(_731_),
    .B(_732_),
    .C(_733_),
    .Y(_50_)
);

INVX1 _1483_ (
    .A(Yin[1]),
    .Y(_734_)
);

NAND2X1 _1484_ (
    .A(Yin3[1]),
    .B(_732_),
    .Y(_735_)
);

OAI21X1 _1485_ (
    .A(_734_),
    .B(_732_),
    .C(_735_),
    .Y(_51_)
);

INVX1 _1486_ (
    .A(Yin[2]),
    .Y(_736_)
);

NAND2X1 _1487_ (
    .A(Yin3[2]),
    .B(_732_),
    .Y(_737_)
);

OAI21X1 _1488_ (
    .A(_736_),
    .B(_732_),
    .C(_737_),
    .Y(_52_)
);

INVX1 _1489_ (
    .A(Yin[3]),
    .Y(_738_)
);

NAND2X1 _1490_ (
    .A(Yin3[3]),
    .B(_732_),
    .Y(_739_)
);

OAI21X1 _1491_ (
    .A(_738_),
    .B(_732_),
    .C(_739_),
    .Y(_53_)
);

NOR2X1 _1492_ (
    .A(_71_),
    .B(_77_),
    .Y(_740_)
);

NOR2X1 _1493_ (
    .A(Yin2[0]),
    .B(_740_),
    .Y(_741_)
);

AOI21X1 _1494_ (
    .A(_731_),
    .B(_740_),
    .C(_741_),
    .Y(_54_)
);

NOR2X1 _1495_ (
    .A(Yin2[1]),
    .B(_740_),
    .Y(_742_)
);

AOI21X1 _1496_ (
    .A(_734_),
    .B(_740_),
    .C(_742_),
    .Y(_55_)
);

NOR2X1 _1497_ (
    .A(Yin2[2]),
    .B(_740_),
    .Y(_743_)
);

AOI21X1 _1498_ (
    .A(_736_),
    .B(_740_),
    .C(_743_),
    .Y(_56_)
);

NOR2X1 _1499_ (
    .A(Yin2[3]),
    .B(_740_),
    .Y(_744_)
);

AOI21X1 _1500_ (
    .A(_738_),
    .B(_740_),
    .C(_744_),
    .Y(_57_)
);

INVX1 _1501_ (
    .A(_75_),
    .Y(_745_)
);

OAI21X1 _1502_ (
    .A(LoadCtl_0_bF$buf4),
    .B(_74_),
    .C(Yin1[0]),
    .Y(_746_)
);

OAI21X1 _1503_ (
    .A(_731_),
    .B(_745_),
    .C(_746_),
    .Y(_58_)
);

OAI21X1 _1504_ (
    .A(LoadCtl_0_bF$buf3),
    .B(_74_),
    .C(Yin1[1]),
    .Y(_747_)
);

OAI21X1 _1505_ (
    .A(_734_),
    .B(_745_),
    .C(_747_),
    .Y(_59_)
);

OAI21X1 _1506_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_74_),
    .C(Yin1[2]),
    .Y(_748_)
);

OAI21X1 _1507_ (
    .A(_736_),
    .B(_745_),
    .C(_748_),
    .Y(_60_)
);

OAI21X1 _1508_ (
    .A(LoadCtl_0_bF$buf1),
    .B(_74_),
    .C(Yin1[3]),
    .Y(_749_)
);

OAI21X1 _1509_ (
    .A(_738_),
    .B(_745_),
    .C(_749_),
    .Y(_61_)
);

NOR2X1 _1510_ (
    .A(LoadCtl_0_bF$buf0),
    .B(Yin0[0]),
    .Y(_750_)
);

AOI21X1 _1511_ (
    .A(LoadCtl_0_bF$buf4),
    .B(_731_),
    .C(_750_),
    .Y(_62_)
);

NOR2X1 _1512_ (
    .A(LoadCtl_0_bF$buf3),
    .B(Yin0[1]),
    .Y(_751_)
);

AOI21X1 _1513_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_734_),
    .C(_751_),
    .Y(_63_)
);

NOR2X1 _1514_ (
    .A(LoadCtl_0_bF$buf1),
    .B(Yin0[2]),
    .Y(_752_)
);

AOI21X1 _1515_ (
    .A(LoadCtl_0_bF$buf0),
    .B(_736_),
    .C(_752_),
    .Y(_64_)
);

NOR2X1 _1516_ (
    .A(LoadCtl_0_bF$buf4),
    .B(Yin0[3]),
    .Y(_753_)
);

AOI21X1 _1517_ (
    .A(LoadCtl_0_bF$buf3),
    .B(_738_),
    .C(_753_),
    .Y(_65_)
);

NAND2X1 _1518_ (
    .A(LoadCtl_0_bF$buf2),
    .B(Xin[0]),
    .Y(_754_)
);

OAI21X1 _1519_ (
    .A(LoadCtl_0_bF$buf1),
    .B(_140_),
    .C(_754_),
    .Y(_66_)
);

NAND2X1 _1520_ (
    .A(LoadCtl_0_bF$buf0),
    .B(Xin[1]),
    .Y(_755_)
);

OAI21X1 _1521_ (
    .A(LoadCtl_0_bF$buf4),
    .B(_236_),
    .C(_755_),
    .Y(_67_)
);

NAND2X1 _1522_ (
    .A(LoadCtl_0_bF$buf3),
    .B(Xin[2]),
    .Y(_756_)
);

OAI21X1 _1523_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_176_),
    .C(_756_),
    .Y(_68_)
);

NAND2X1 _1524_ (
    .A(LoadCtl_0_bF$buf1),
    .B(Xin[3]),
    .Y(_757_)
);

OAI21X1 _1525_ (
    .A(LoadCtl_0_bF$buf0),
    .B(_178_),
    .C(_757_),
    .Y(_69_)
);

DFFPOSX1 _1526_ (
    .CLK(clk_bF$buf7),
    .D(_0_),
    .Q(XinH[0])
);

DFFPOSX1 _1527_ (
    .CLK(clk_bF$buf6),
    .D(_1_),
    .Q(XinH[1])
);

DFFPOSX1 _1528_ (
    .CLK(clk_bF$buf5),
    .D(_2_),
    .Q(XinH[2])
);

DFFPOSX1 _1529_ (
    .CLK(clk_bF$buf4),
    .D(_3_),
    .Q(XinH[3])
);

DFFPOSX1 _1530_ (
    .CLK(clk_bF$buf3),
    .D(_4_),
    .Q(rYin[0])
);

DFFPOSX1 _1531_ (
    .CLK(clk_bF$buf2),
    .D(_5_),
    .Q(rYin[1])
);

DFFPOSX1 _1532_ (
    .CLK(clk_bF$buf1),
    .D(_6_),
    .Q(rYin[2])
);

DFFPOSX1 _1533_ (
    .CLK(clk_bF$buf0),
    .D(_7_),
    .Q(rYin[3])
);

DFFPOSX1 _1534_ (
    .CLK(clk_bF$buf7),
    .D(_8_),
    .Q(rYin[4])
);

DFFPOSX1 _1535_ (
    .CLK(clk_bF$buf6),
    .D(_9_),
    .Q(rYin[5])
);

DFFPOSX1 _1536_ (
    .CLK(clk_bF$buf5),
    .D(_10_),
    .Q(rYin[6])
);

DFFPOSX1 _1537_ (
    .CLK(clk_bF$buf4),
    .D(_11_),
    .Q(rYin[7])
);

DFFPOSX1 _1538_ (
    .CLK(clk_bF$buf3),
    .D(_12_),
    .Q(rYin[8])
);

DFFPOSX1 _1539_ (
    .CLK(clk_bF$buf2),
    .D(_13_),
    .Q(rYin[9])
);

DFFPOSX1 _1540_ (
    .CLK(clk_bF$buf1),
    .D(_14_),
    .Q(rYin[10])
);

DFFPOSX1 _1541_ (
    .CLK(clk_bF$buf0),
    .D(_15_),
    .Q(rYin[11])
);

DFFPOSX1 _1542_ (
    .CLK(clk_bF$buf7),
    .D(_16_),
    .Q(rYin[12])
);

DFFPOSX1 _1543_ (
    .CLK(clk_bF$buf6),
    .D(_17_),
    .Q(rYin[13])
);

DFFPOSX1 _1544_ (
    .CLK(clk_bF$buf5),
    .D(_18_),
    .Q(rYin[14])
);

DFFPOSX1 _1545_ (
    .CLK(clk_bF$buf4),
    .D(_19_),
    .Q(rYin[15])
);

DFFPOSX1 _1546_ (
    .CLK(clk_bF$buf3),
    .D(_20_),
    .Q(mul[0])
);

DFFPOSX1 _1547_ (
    .CLK(clk_bF$buf2),
    .D(_21_),
    .Q(mul[1])
);

DFFPOSX1 _1548_ (
    .CLK(clk_bF$buf1),
    .D(_22_),
    .Q(mul[2])
);

DFFPOSX1 _1549_ (
    .CLK(clk_bF$buf0),
    .D(_23_),
    .Q(mul[3])
);

DFFPOSX1 _1550_ (
    .CLK(clk_bF$buf7),
    .D(_24_),
    .Q(mul[4])
);

DFFPOSX1 _1551_ (
    .CLK(clk_bF$buf6),
    .D(_25_),
    .Q(mul[5])
);

DFFPOSX1 _1552_ (
    .CLK(clk_bF$buf5),
    .D(_26_),
    .Q(mul[6])
);

DFFPOSX1 _1553_ (
    .CLK(clk_bF$buf4),
    .D(_27_),
    .Q(mul[7])
);

DFFPOSX1 _1554_ (
    .CLK(clk_bF$buf3),
    .D(_28_),
    .Q(mul[8])
);

DFFPOSX1 _1555_ (
    .CLK(clk_bF$buf2),
    .D(_29_),
    .Q(mul[9])
);

DFFPOSX1 _1556_ (
    .CLK(clk_bF$buf1),
    .D(_30_),
    .Q(mul[10])
);

DFFPOSX1 _1557_ (
    .CLK(clk_bF$buf0),
    .D(_31_),
    .Q(mul[11])
);

DFFPOSX1 _1558_ (
    .CLK(clk_bF$buf7),
    .D(_32_),
    .Q(mul[12])
);

DFFPOSX1 _1559_ (
    .CLK(clk_bF$buf6),
    .D(_33_),
    .Q(mul[13])
);

DFFPOSX1 _1560_ (
    .CLK(clk_bF$buf5),
    .D(_34_),
    .Q(y[0])
);

DFFPOSX1 _1561_ (
    .CLK(clk_bF$buf4),
    .D(_35_),
    .Q(y[1])
);

DFFPOSX1 _1562_ (
    .CLK(clk_bF$buf3),
    .D(_36_),
    .Q(y[2])
);

DFFPOSX1 _1563_ (
    .CLK(clk_bF$buf2),
    .D(_37_),
    .Q(y[3])
);

DFFPOSX1 _1564_ (
    .CLK(clk_bF$buf1),
    .D(_38_),
    .Q(y[4])
);

DFFPOSX1 _1565_ (
    .CLK(clk_bF$buf0),
    .D(_39_),
    .Q(y[5])
);

DFFPOSX1 _1566_ (
    .CLK(clk_bF$buf7),
    .D(_40_),
    .Q(y[6])
);

DFFPOSX1 _1567_ (
    .CLK(clk_bF$buf6),
    .D(_41_),
    .Q(y[7])
);

DFFPOSX1 _1568_ (
    .CLK(clk_bF$buf5),
    .D(_42_),
    .Q(y[8])
);

DFFPOSX1 _1569_ (
    .CLK(clk_bF$buf4),
    .D(_43_),
    .Q(y[9])
);

DFFPOSX1 _1570_ (
    .CLK(clk_bF$buf3),
    .D(_44_),
    .Q(y[10])
);

DFFPOSX1 _1571_ (
    .CLK(clk_bF$buf2),
    .D(_45_),
    .Q(y[11])
);

DFFPOSX1 _1572_ (
    .CLK(clk_bF$buf1),
    .D(_46_),
    .Q(y[12])
);

DFFPOSX1 _1573_ (
    .CLK(clk_bF$buf0),
    .D(_47_),
    .Q(y[13])
);

DFFPOSX1 _1574_ (
    .CLK(clk_bF$buf7),
    .D(_48_),
    .Q(y[14])
);

DFFPOSX1 _1575_ (
    .CLK(clk_bF$buf6),
    .D(_49_),
    .Q(y[15])
);

DFFPOSX1 _1576_ (
    .CLK(clk_bF$buf5),
    .D(_50_),
    .Q(Yin3[0])
);

DFFPOSX1 _1577_ (
    .CLK(clk_bF$buf4),
    .D(_51_),
    .Q(Yin3[1])
);

DFFPOSX1 _1578_ (
    .CLK(clk_bF$buf3),
    .D(_52_),
    .Q(Yin3[2])
);

DFFPOSX1 _1579_ (
    .CLK(clk_bF$buf2),
    .D(_53_),
    .Q(Yin3[3])
);

DFFPOSX1 _1580_ (
    .CLK(clk_bF$buf1),
    .D(_54_),
    .Q(Yin2[0])
);

DFFPOSX1 _1581_ (
    .CLK(clk_bF$buf0),
    .D(_55_),
    .Q(Yin2[1])
);

DFFPOSX1 _1582_ (
    .CLK(clk_bF$buf7),
    .D(_56_),
    .Q(Yin2[2])
);

DFFPOSX1 _1583_ (
    .CLK(clk_bF$buf6),
    .D(_57_),
    .Q(Yin2[3])
);

DFFPOSX1 _1584_ (
    .CLK(clk_bF$buf5),
    .D(_58_),
    .Q(Yin1[0])
);

DFFPOSX1 _1585_ (
    .CLK(clk_bF$buf4),
    .D(_59_),
    .Q(Yin1[1])
);

DFFPOSX1 _1586_ (
    .CLK(clk_bF$buf3),
    .D(_60_),
    .Q(Yin1[2])
);

DFFPOSX1 _1587_ (
    .CLK(clk_bF$buf2),
    .D(_61_),
    .Q(Yin1[3])
);

DFFPOSX1 _1588_ (
    .CLK(clk_bF$buf1),
    .D(_62_),
    .Q(Yin0[0])
);

DFFPOSX1 _1589_ (
    .CLK(clk_bF$buf0),
    .D(_63_),
    .Q(Yin0[1])
);

DFFPOSX1 _1590_ (
    .CLK(clk_bF$buf7),
    .D(_64_),
    .Q(Yin0[2])
);

DFFPOSX1 _1591_ (
    .CLK(clk_bF$buf6),
    .D(_65_),
    .Q(Yin0[3])
);

DFFPOSX1 _1592_ (
    .CLK(clk_bF$buf5),
    .D(_66_),
    .Q(XinHL[0])
);

DFFPOSX1 _1593_ (
    .CLK(clk_bF$buf4),
    .D(_67_),
    .Q(XinHL[1])
);

DFFPOSX1 _1594_ (
    .CLK(clk_bF$buf3),
    .D(_68_),
    .Q(XinHL[2])
);

DFFPOSX1 _1595_ (
    .CLK(clk_bF$buf2),
    .D(_69_),
    .Q(XinHL[3])
);

DFFPOSX1 _1596_ (
    .CLK(clk_bF$buf1),
    .D(Rdy),
    .Q(LoadCtl[0])
);

DFFPOSX1 _1597_ (
    .CLK(clk_bF$buf0),
    .D(LoadCtl_0_bF$buf4),
    .Q(LoadCtl[1])
);

DFFPOSX1 _1598_ (
    .CLK(clk_bF$buf7),
    .D(LoadCtl[1]),
    .Q(LoadCtl[2])
);

DFFPOSX1 _1599_ (
    .CLK(clk_bF$buf6),
    .D(LoadCtl[2]),
    .Q(LoadCtl[3])
);

DFFPOSX1 _1600_ (
    .CLK(clk_bF$buf5),
    .D(LoadCtl[3]),
    .Q(LoadCtl[4])
);

BUFX2 _1601_ (
    .A(LoadCtl_4_bF$buf7),
    .Y(Vld)
);

BUFX2 _1602_ (
    .A(_758_[0]),
    .Y(Xout[0])
);

BUFX2 _1603_ (
    .A(_758_[1]),
    .Y(Xout[1])
);

BUFX2 _1604_ (
    .A(_758_[2]),
    .Y(Xout[2])
);

BUFX2 _1605_ (
    .A(_758_[3]),
    .Y(Xout[3])
);

BUFX2 _1606_ (
    .A(_759_[0]),
    .Y(Yout[0])
);

BUFX2 _1607_ (
    .A(_759_[1]),
    .Y(Yout[1])
);

BUFX2 _1608_ (
    .A(_759_[2]),
    .Y(Yout[2])
);

BUFX2 _1609_ (
    .A(_759_[3]),
    .Y(Yout[3])
);

NOR2X1 _760_ (
    .A(LoadCtl[2]),
    .B(y[12]),
    .Y(_70_)
);

INVX1 _761_ (
    .A(LoadCtl[2]),
    .Y(_71_)
);

NOR2X1 _762_ (
    .A(LoadCtl[1]),
    .B(LoadCtl_0_bF$buf3),
    .Y(_72_)
);

OAI21X1 _763_ (
    .A(_71_),
    .B(y[8]),
    .C(_72_),
    .Y(_73_)
);

INVX2 _764_ (
    .A(LoadCtl[1]),
    .Y(_74_)
);

NOR2X1 _765_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_74_),
    .Y(_75_)
);

AOI22X1 _766_ (
    .A(LoadCtl_0_bF$buf1),
    .B(y[0]),
    .C(_75_),
    .D(y[4]),
    .Y(_76_)
);

OAI21X1 _767_ (
    .A(_70_),
    .B(_73_),
    .C(_76_),
    .Y(_759_[0])
);

INVX1 _768_ (
    .A(_72_),
    .Y(_77_)
);

INVX1 _769_ (
    .A(y[9]),
    .Y(_78_)
);

NAND2X1 _770_ (
    .A(LoadCtl[2]),
    .B(_78_),
    .Y(_79_)
);

OAI21X1 _771_ (
    .A(LoadCtl[2]),
    .B(y[13]),
    .C(_79_),
    .Y(_80_)
);

AOI22X1 _772_ (
    .A(LoadCtl_0_bF$buf0),
    .B(y[1]),
    .C(_75_),
    .D(y[5]),
    .Y(_81_)
);

OAI21X1 _773_ (
    .A(_77_),
    .B(_80_),
    .C(_81_),
    .Y(_759_[1])
);

NOR2X1 _774_ (
    .A(LoadCtl[2]),
    .B(y[14]),
    .Y(_82_)
);

OAI21X1 _775_ (
    .A(_71_),
    .B(y[10]),
    .C(_72_),
    .Y(_83_)
);

AOI22X1 _776_ (
    .A(LoadCtl_0_bF$buf4),
    .B(y[2]),
    .C(_75_),
    .D(y[6]),
    .Y(_84_)
);

OAI21X1 _777_ (
    .A(_82_),
    .B(_83_),
    .C(_84_),
    .Y(_759_[2])
);

INVX1 _778_ (
    .A(y[11]),
    .Y(_85_)
);

NAND2X1 _779_ (
    .A(LoadCtl[2]),
    .B(_85_),
    .Y(_86_)
);

OAI21X1 _780_ (
    .A(LoadCtl[2]),
    .B(y[15]),
    .C(_86_),
    .Y(_87_)
);

AOI22X1 _781_ (
    .A(LoadCtl_0_bF$buf3),
    .B(y[3]),
    .C(_75_),
    .D(y[7]),
    .Y(_88_)
);

OAI21X1 _782_ (
    .A(_77_),
    .B(_87_),
    .C(_88_),
    .Y(_759_[3])
);

INVX2 _783_ (
    .A(XinH[0]),
    .Y(_89_)
);

NAND2X1 _784_ (
    .A(LoadCtl_0_bF$buf2),
    .B(XinHL[0]),
    .Y(_90_)
);

OAI21X1 _785_ (
    .A(LoadCtl_0_bF$buf1),
    .B(_89_),
    .C(_90_),
    .Y(_758_[0])
);

INVX2 _786_ (
    .A(XinH[1]),
    .Y(_91_)
);

NAND2X1 _787_ (
    .A(LoadCtl_0_bF$buf0),
    .B(XinHL[1]),
    .Y(_92_)
);

OAI21X1 _788_ (
    .A(LoadCtl_0_bF$buf4),
    .B(_91_),
    .C(_92_),
    .Y(_758_[1])
);

INVX2 _789_ (
    .A(XinH[2]),
    .Y(_93_)
);

NAND2X1 _790_ (
    .A(LoadCtl_0_bF$buf3),
    .B(XinHL[2]),
    .Y(_94_)
);

OAI21X1 _791_ (
    .A(LoadCtl_0_bF$buf2),
    .B(_93_),
    .C(_94_),
    .Y(_758_[2])
);

INVX2 _792_ (
    .A(XinH[3]),
    .Y(_95_)
);

NAND2X1 _793_ (
    .A(LoadCtl_0_bF$buf1),
    .B(XinHL[3]),
    .Y(_96_)
);

OAI21X1 _794_ (
    .A(LoadCtl_0_bF$buf0),
    .B(_95_),
    .C(_96_),
    .Y(_758_[3])
);

NAND2X1 _795_ (
    .A(Xin[0]),
    .B(_75_),
    .Y(_97_)
);

OAI21X1 _796_ (
    .A(_89_),
    .B(_75_),
    .C(_97_),
    .Y(_0_)
);

NAND2X1 _797_ (
    .A(Xin[1]),
    .B(_75_),
    .Y(_98_)
);

OAI21X1 _798_ (
    .A(_91_),
    .B(_75_),
    .C(_98_),
    .Y(_1_)
);

NAND2X1 _799_ (
    .A(Xin[2]),
    .B(_75_),
    .Y(_99_)
);

OAI21X1 _800_ (
    .A(_93_),
    .B(_75_),
    .C(_99_),
    .Y(_2_)
);

NAND2X1 _801_ (
    .A(Xin[3]),
    .B(_75_),
    .Y(_100_)
);

OAI21X1 _802_ (
    .A(_95_),
    .B(_75_),
    .C(_100_),
    .Y(_3_)
);

INVX1 _803_ (
    .A(rYin[0]),
    .Y(_101_)
);

NAND2X1 _804_ (
    .A(Yin0[0]),
    .B(LoadCtl_4_bF$buf6),
    .Y(_102_)
);

OAI21X1 _805_ (
    .A(LoadCtl_4_bF$buf5),
    .B(_101_),
    .C(_102_),
    .Y(_4_)
);

INVX1 _806_ (
    .A(rYin[1]),
    .Y(_103_)
);

NAND2X1 _807_ (
    .A(LoadCtl_4_bF$buf4),
    .B(Yin0[1]),
    .Y(_104_)
);

OAI21X1 _808_ (
    .A(LoadCtl_4_bF$buf3),
    .B(_103_),
    .C(_104_),
    .Y(_5_)
);

INVX1 _809_ (
    .A(rYin[2]),
    .Y(_105_)
);

NAND2X1 _810_ (
    .A(LoadCtl_4_bF$buf2),
    .B(Yin0[2]),
    .Y(_106_)
);

OAI21X1 _811_ (
    .A(LoadCtl_4_bF$buf1),
    .B(_105_),
    .C(_106_),
    .Y(_6_)
);

INVX1 _812_ (
    .A(rYin[3]),
    .Y(_107_)
);

NAND2X1 _813_ (
    .A(LoadCtl_4_bF$buf0),
    .B(Yin0[3]),
    .Y(_108_)
);

OAI21X1 _814_ (
    .A(LoadCtl_4_bF$buf7),
    .B(_107_),
    .C(_108_),
    .Y(_7_)
);

INVX1 _815_ (
    .A(rYin[4]),
    .Y(_109_)
);

NAND2X1 _816_ (
    .A(LoadCtl_4_bF$buf6),
    .B(Yin1[0]),
    .Y(_110_)
);

OAI21X1 _817_ (
    .A(LoadCtl_4_bF$buf5),
    .B(_109_),
    .C(_110_),
    .Y(_8_)
);

INVX1 _818_ (
    .A(rYin[5]),
    .Y(_111_)
);

NAND2X1 _819_ (
    .A(LoadCtl_4_bF$buf4),
    .B(Yin1[1]),
    .Y(_112_)
);

OAI21X1 _820_ (
    .A(LoadCtl_4_bF$buf3),
    .B(_111_),
    .C(_112_),
    .Y(_9_)
);

INVX1 _821_ (
    .A(rYin[6]),
    .Y(_113_)
);

NAND2X1 _822_ (
    .A(LoadCtl_4_bF$buf2),
    .B(Yin1[2]),
    .Y(_114_)
);

OAI21X1 _823_ (
    .A(LoadCtl_4_bF$buf1),
    .B(_113_),
    .C(_114_),
    .Y(_10_)
);

INVX1 _824_ (
    .A(rYin[7]),
    .Y(_115_)
);

NAND2X1 _825_ (
    .A(LoadCtl_4_bF$buf0),
    .B(Yin1[3]),
    .Y(_116_)
);

OAI21X1 _826_ (
    .A(LoadCtl_4_bF$buf7),
    .B(_115_),
    .C(_116_),
    .Y(_11_)
);

INVX1 _827_ (
    .A(rYin[8]),
    .Y(_117_)
);

NAND2X1 _828_ (
    .A(LoadCtl_4_bF$buf6),
    .B(Yin2[0]),
    .Y(_118_)
);

OAI21X1 _829_ (
    .A(LoadCtl_4_bF$buf5),
    .B(_117_),
    .C(_118_),
    .Y(_12_)
);

INVX1 _830_ (
    .A(rYin[9]),
    .Y(_119_)
);

NAND2X1 _831_ (
    .A(LoadCtl_4_bF$buf4),
    .B(Yin2[1]),
    .Y(_120_)
);

OAI21X1 _832_ (
    .A(LoadCtl_4_bF$buf3),
    .B(_119_),
    .C(_120_),
    .Y(_13_)
);

INVX1 _833_ (
    .A(rYin[10]),
    .Y(_121_)
);

NAND2X1 _834_ (
    .A(LoadCtl_4_bF$buf2),
    .B(Yin2[2]),
    .Y(_122_)
);

OAI21X1 _835_ (
    .A(LoadCtl_4_bF$buf1),
    .B(_121_),
    .C(_122_),
    .Y(_14_)
);

INVX1 _836_ (
    .A(rYin[11]),
    .Y(_123_)
);

NAND2X1 _837_ (
    .A(LoadCtl_4_bF$buf0),
    .B(Yin2[3]),
    .Y(_124_)
);

OAI21X1 _838_ (
    .A(LoadCtl_4_bF$buf7),
    .B(_123_),
    .C(_124_),
    .Y(_15_)
);

INVX1 _839_ (
    .A(rYin[12]),
    .Y(_125_)
);

NAND2X1 _840_ (
    .A(LoadCtl_4_bF$buf6),
    .B(Yin3[0]),
    .Y(_126_)
);

OAI21X1 _841_ (
    .A(LoadCtl_4_bF$buf5),
    .B(_125_),
    .C(_126_),
    .Y(_16_)
);

INVX1 _842_ (
    .A(rYin[13]),
    .Y(_127_)
);

NAND2X1 _843_ (
    .A(LoadCtl_4_bF$buf4),
    .B(Yin3[1]),
    .Y(_128_)
);

OAI21X1 _844_ (
    .A(LoadCtl_4_bF$buf3),
    .B(_127_),
    .C(_128_),
    .Y(_17_)
);

INVX1 _845_ (
    .A(rYin[14]),
    .Y(_129_)
);

NAND2X1 _846_ (
    .A(LoadCtl_4_bF$buf2),
    .B(Yin3[2]),
    .Y(_130_)
);

OAI21X1 _847_ (
    .A(LoadCtl_4_bF$buf1),
    .B(_129_),
    .C(_130_),
    .Y(_18_)
);

INVX1 _848_ (
    .A(rYin[15]),
    .Y(_131_)
);

NAND2X1 _849_ (
    .A(LoadCtl_4_bF$buf0),
    .B(Yin3[3]),
    .Y(_132_)
);

OAI21X1 _850_ (
    .A(LoadCtl_4_bF$buf7),
    .B(_131_),
    .C(_132_),
    .Y(_19_)
);

INVX1 _851_ (
    .A(mul[0]),
    .Y(_133_)
);

NAND3X1 _852_ (
    .A(XinHL[0]),
    .B(Cin_0_bF$buf1),
    .C(LoadCtl_4_bF$buf6),
    .Y(_134_)
);

OAI21X1 _853_ (
    .A(_133_),
    .B(LoadCtl_4_bF$buf5),
    .C(_134_),
    .Y(_20_)
);

INVX1 _854_ (
    .A(mul[1]),
    .Y(_135_)
);

NAND2X1 _855_ (
    .A(XinHL[0]),
    .B(Cin_1_bF$buf3),
    .Y(_136_)
);

NAND2X1 _856_ (
    .A(XinHL[1]),
    .B(Cin_0_bF$buf0),
    .Y(_137_)
);

NOR2X1 _857_ (
    .A(_136_),
    .B(_137_),
    .Y(_138_)
);

INVX1 _858_ (
    .A(_138_),
    .Y(_139_)
);

INVX1 _859_ (
    .A(XinHL[0]),
    .Y(_140_)
);

INVX2 _860_ (
    .A(Cin_1_bF$buf2),
    .Y(_141_)
);

OAI21X1 _861_ (
    .A(_140_),
    .B(_141_),
    .C(_137_),
    .Y(_142_)
);

NAND3X1 _862_ (
    .A(LoadCtl_4_bF$buf4),
    .B(_142_),
    .C(_139_),
    .Y(_143_)
);

OAI21X1 _863_ (
    .A(_135_),
    .B(LoadCtl_4_bF$buf3),
    .C(_143_),
    .Y(_21_)
);

INVX1 _864_ (
    .A(mul[2]),
    .Y(_144_)
);

NAND2X1 _865_ (
    .A(XinHL[0]),
    .B(Cin[2]),
    .Y(_145_)
);

NAND2X1 _866_ (
    .A(XinHL[2]),
    .B(Cin_1_bF$buf1),
    .Y(_146_)
);

NOR2X1 _867_ (
    .A(_137_),
    .B(_146_),
    .Y(_147_)
);

AOI22X1 _868_ (
    .A(XinHL[1]),
    .B(Cin_1_bF$buf0),
    .C(XinHL[2]),
    .D(Cin_0_bF$buf3),
    .Y(_148_)
);

OAI21X1 _869_ (
    .A(_148_),
    .B(_147_),
    .C(_145_),
    .Y(_149_)
);

INVX1 _870_ (
    .A(_145_),
    .Y(_150_)
);

AND2X2 _871_ (
    .A(XinHL[2]),
    .B(Cin_1_bF$buf3),
    .Y(_151_)
);

NAND3X1 _872_ (
    .A(XinHL[1]),
    .B(Cin_0_bF$buf2),
    .C(_151_),
    .Y(_152_)
);

INVX1 _873_ (
    .A(_148_),
    .Y(_153_)
);

NAND3X1 _874_ (
    .A(_150_),
    .B(_153_),
    .C(_152_),
    .Y(_154_)
);

NAND3X1 _875_ (
    .A(_138_),
    .B(_154_),
    .C(_149_),
    .Y(_155_)
);

INVX1 _876_ (
    .A(_155_),
    .Y(_156_)
);

AOI21X1 _877_ (
    .A(_149_),
    .B(_154_),
    .C(_138_),
    .Y(_157_)
);

NOR2X1 _878_ (
    .A(_157_),
    .B(_156_),
    .Y(_158_)
);

NAND2X1 _879_ (
    .A(LoadCtl_4_bF$buf2),
    .B(_158_),
    .Y(_159_)
);

OAI21X1 _880_ (
    .A(_144_),
    .B(LoadCtl_4_bF$buf1),
    .C(_159_),
    .Y(_22_)
);

INVX1 _881_ (
    .A(mul[3]),
    .Y(_160_)
);

NAND2X1 _882_ (
    .A(XinHL[0]),
    .B(Cin[3]),
    .Y(_161_)
);

AOI21X1 _883_ (
    .A(_150_),
    .B(_153_),
    .C(_147_),
    .Y(_162_)
);

NAND2X1 _884_ (
    .A(XinHL[1]),
    .B(Cin[2]),
    .Y(_163_)
);

NAND2X1 _885_ (
    .A(XinHL[3]),
    .B(Cin_0_bF$buf1),
    .Y(_164_)
);

NOR2X1 _886_ (
    .A(_146_),
    .B(_164_),
    .Y(_165_)
);

AOI22X1 _887_ (
    .A(XinHL[2]),
    .B(Cin_1_bF$buf2),
    .C(XinHL[3]),
    .D(Cin_0_bF$buf0),
    .Y(_166_)
);

OAI21X1 _888_ (
    .A(_166_),
    .B(_165_),
    .C(_163_),
    .Y(_167_)
);

INVX1 _889_ (
    .A(_163_),
    .Y(_168_)
);

AND2X2 _890_ (
    .A(XinHL[3]),
    .B(Cin_0_bF$buf3),
    .Y(_169_)
);

NAND2X1 _891_ (
    .A(_151_),
    .B(_169_),
    .Y(_170_)
);

INVX1 _892_ (
    .A(_166_),
    .Y(_171_)
);

NAND3X1 _893_ (
    .A(_168_),
    .B(_171_),
    .C(_170_),
    .Y(_172_)
);

NAND3X1 _894_ (
    .A(_172_),
    .B(_167_),
    .C(_162_),
    .Y(_173_)
);

OAI21X1 _895_ (
    .A(_145_),
    .B(_148_),
    .C(_152_),
    .Y(_174_)
);

AOI21X1 _896_ (
    .A(_170_),
    .B(_171_),
    .C(_168_),
    .Y(_175_)
);

INVX2 _897_ (
    .A(XinHL[2]),
    .Y(_176_)
);

OAI21X1 _898_ (
    .A(_176_),
    .B(_141_),
    .C(_169_),
    .Y(_177_)
);

INVX2 _899_ (
    .A(XinHL[3]),
    .Y(_178_)
);

INVX1 _900_ (
    .A(Cin_0_bF$buf2),
    .Y(_179_)
);

OAI21X1 _901_ (
    .A(_178_),
    .B(_179_),
    .C(_151_),
    .Y(_180_)
);

AOI21X1 _902_ (
    .A(_177_),
    .B(_180_),
    .C(_163_),
    .Y(_181_)
);

OAI21X1 _903_ (
    .A(_175_),
    .B(_181_),
    .C(_174_),
    .Y(_182_)
);

NAND3X1 _904_ (
    .A(_161_),
    .B(_173_),
    .C(_182_),
    .Y(_183_)
);

INVX1 _905_ (
    .A(_161_),
    .Y(_184_)
);

NAND3X1 _906_ (
    .A(_174_),
    .B(_172_),
    .C(_167_),
    .Y(_185_)
);

OAI21X1 _907_ (
    .A(_175_),
    .B(_181_),
    .C(_162_),
    .Y(_186_)
);

NAND3X1 _908_ (
    .A(_184_),
    .B(_185_),
    .C(_186_),
    .Y(_187_)
);

AOI21X1 _909_ (
    .A(_183_),
    .B(_187_),
    .C(_156_),
    .Y(_188_)
);

NAND3X1 _910_ (
    .A(_156_),
    .B(_183_),
    .C(_187_),
    .Y(_189_)
);

NAND2X1 _911_ (
    .A(LoadCtl_4_bF$buf0),
    .B(_189_),
    .Y(_190_)
);

OAI22X1 _912_ (
    .A(_160_),
    .B(LoadCtl_4_bF$buf7),
    .C(_188_),
    .D(_190_),
    .Y(_23_)
);

INVX1 _913_ (
    .A(mul[4]),
    .Y(_191_)
);

INVX1 _914_ (
    .A(_189_),
    .Y(_192_)
);

AOI21X1 _915_ (
    .A(_167_),
    .B(_172_),
    .C(_174_),
    .Y(_193_)
);

OAI21X1 _916_ (
    .A(_161_),
    .B(_193_),
    .C(_185_),
    .Y(_194_)
);

OAI21X1 _917_ (
    .A(_163_),
    .B(_166_),
    .C(_170_),
    .Y(_195_)
);

AND2X2 _918_ (
    .A(XinH[0]),
    .B(Cin_1_bF$buf1),
    .Y(_196_)
);

NAND2X1 _919_ (
    .A(_169_),
    .B(_196_),
    .Y(_197_)
);

AOI22X1 _920_ (
    .A(XinH[0]),
    .B(Cin_0_bF$buf1),
    .C(XinHL[3]),
    .D(Cin_1_bF$buf0),
    .Y(_198_)
);

INVX1 _921_ (
    .A(_198_),
    .Y(_199_)
);

NAND2X1 _922_ (
    .A(XinHL[2]),
    .B(Cin[2]),
    .Y(_200_)
);

INVX1 _923_ (
    .A(_200_),
    .Y(_201_)
);

NAND3X1 _924_ (
    .A(_201_),
    .B(_199_),
    .C(_197_),
    .Y(_202_)
);

NAND2X1 _925_ (
    .A(XinH[0]),
    .B(Cin_1_bF$buf3),
    .Y(_203_)
);

NOR2X1 _926_ (
    .A(_164_),
    .B(_203_),
    .Y(_204_)
);

OAI21X1 _927_ (
    .A(_198_),
    .B(_204_),
    .C(_200_),
    .Y(_205_)
);

AOI21X1 _928_ (
    .A(_205_),
    .B(_202_),
    .C(_195_),
    .Y(_206_)
);

AOI21X1 _929_ (
    .A(_168_),
    .B(_171_),
    .C(_165_),
    .Y(_207_)
);

NAND3X1 _930_ (
    .A(_200_),
    .B(_199_),
    .C(_197_),
    .Y(_208_)
);

OAI21X1 _931_ (
    .A(_198_),
    .B(_204_),
    .C(_201_),
    .Y(_209_)
);

AOI21X1 _932_ (
    .A(_209_),
    .B(_208_),
    .C(_207_),
    .Y(_210_)
);

NAND2X1 _933_ (
    .A(XinHL[1]),
    .B(Cin[4]),
    .Y(_211_)
);

INVX2 _934_ (
    .A(Cin[4]),
    .Y(_212_)
);

NAND2X1 _935_ (
    .A(XinHL[1]),
    .B(Cin[3]),
    .Y(_213_)
);

OAI21X1 _936_ (
    .A(_140_),
    .B(_212_),
    .C(_213_),
    .Y(_214_)
);

OAI21X1 _937_ (
    .A(_161_),
    .B(_211_),
    .C(_214_),
    .Y(_215_)
);

OAI21X1 _938_ (
    .A(_206_),
    .B(_210_),
    .C(_215_),
    .Y(_216_)
);

NAND3X1 _939_ (
    .A(_208_),
    .B(_209_),
    .C(_207_),
    .Y(_217_)
);

NAND3X1 _940_ (
    .A(_195_),
    .B(_202_),
    .C(_205_),
    .Y(_218_)
);

INVX1 _941_ (
    .A(_215_),
    .Y(_219_)
);

NAND3X1 _942_ (
    .A(_219_),
    .B(_218_),
    .C(_217_),
    .Y(_220_)
);

NAND3X1 _943_ (
    .A(_220_),
    .B(_194_),
    .C(_216_),
    .Y(_221_)
);

INVX1 _944_ (
    .A(_185_),
    .Y(_222_)
);

AOI21X1 _945_ (
    .A(_184_),
    .B(_186_),
    .C(_222_),
    .Y(_223_)
);

AOI21X1 _946_ (
    .A(_217_),
    .B(_218_),
    .C(_219_),
    .Y(_224_)
);

INVX1 _947_ (
    .A(_220_),
    .Y(_225_)
);

OAI21X1 _948_ (
    .A(_224_),
    .B(_225_),
    .C(_223_),
    .Y(_226_)
);

AOI21X1 _949_ (
    .A(_221_),
    .B(_226_),
    .C(_192_),
    .Y(_227_)
);

NAND3X1 _950_ (
    .A(_221_),
    .B(_226_),
    .C(_192_),
    .Y(_228_)
);

NAND2X1 _951_ (
    .A(LoadCtl_4_bF$buf6),
    .B(_228_),
    .Y(_229_)
);

OAI22X1 _952_ (
    .A(_191_),
    .B(LoadCtl_4_bF$buf5),
    .C(_227_),
    .D(_229_),
    .Y(_24_)
);

INVX1 _953_ (
    .A(mul[5]),
    .Y(_230_)
);

AND2X2 _954_ (
    .A(XinHL[1]),
    .B(Cin[4]),
    .Y(_231_)
);

NAND2X1 _955_ (
    .A(_231_),
    .B(_184_),
    .Y(_232_)
);

INVX1 _956_ (
    .A(_232_),
    .Y(_233_)
);

AOI21X1 _957_ (
    .A(_217_),
    .B(_219_),
    .C(_210_),
    .Y(_234_)
);

NAND2X1 _958_ (
    .A(XinHL[0]),
    .B(Cin[5]),
    .Y(_235_)
);

INVX1 _959_ (
    .A(XinHL[1]),
    .Y(_236_)
);

AND2X2 _960_ (
    .A(XinHL[2]),
    .B(Cin[3]),
    .Y(_237_)
);

OAI21X1 _961_ (
    .A(_236_),
    .B(_212_),
    .C(_237_),
    .Y(_238_)
);

INVX2 _962_ (
    .A(Cin[3]),
    .Y(_239_)
);

OAI21X1 _963_ (
    .A(_176_),
    .B(_239_),
    .C(_231_),
    .Y(_240_)
);

NAND3X1 _964_ (
    .A(_235_),
    .B(_238_),
    .C(_240_),
    .Y(_241_)
);

INVX1 _965_ (
    .A(_235_),
    .Y(_242_)
);

NAND2X1 _966_ (
    .A(_231_),
    .B(_237_),
    .Y(_243_)
);

OAI21X1 _967_ (
    .A(_176_),
    .B(_239_),
    .C(_211_),
    .Y(_244_)
);

NAND3X1 _968_ (
    .A(_244_),
    .B(_242_),
    .C(_243_),
    .Y(_245_)
);

NAND2X1 _969_ (
    .A(_245_),
    .B(_241_),
    .Y(_246_)
);

AOI21X1 _970_ (
    .A(_199_),
    .B(_201_),
    .C(_204_),
    .Y(_247_)
);

NAND2X1 _971_ (
    .A(XinHL[3]),
    .B(Cin[2]),
    .Y(_248_)
);

AND2X2 _972_ (
    .A(XinH[1]),
    .B(Cin_0_bF$buf0),
    .Y(_249_)
);

NAND2X1 _973_ (
    .A(_203_),
    .B(_249_),
    .Y(_250_)
);

NAND2X1 _974_ (
    .A(XinH[1]),
    .B(Cin_0_bF$buf3),
    .Y(_251_)
);

NAND2X1 _975_ (
    .A(_251_),
    .B(_196_),
    .Y(_252_)
);

NAND3X1 _976_ (
    .A(_248_),
    .B(_250_),
    .C(_252_),
    .Y(_253_)
);

INVX1 _977_ (
    .A(_248_),
    .Y(_254_)
);

NAND2X1 _978_ (
    .A(_196_),
    .B(_249_),
    .Y(_255_)
);

OAI21X1 _979_ (
    .A(_91_),
    .B(_179_),
    .C(_203_),
    .Y(_256_)
);

NAND3X1 _980_ (
    .A(_256_),
    .B(_254_),
    .C(_255_),
    .Y(_257_)
);

NAND3X1 _981_ (
    .A(_253_),
    .B(_257_),
    .C(_247_),
    .Y(_258_)
);

OAI21X1 _982_ (
    .A(_198_),
    .B(_200_),
    .C(_197_),
    .Y(_259_)
);

AOI21X1 _983_ (
    .A(_255_),
    .B(_256_),
    .C(_254_),
    .Y(_260_)
);

AOI21X1 _984_ (
    .A(_250_),
    .B(_252_),
    .C(_248_),
    .Y(_261_)
);

OAI21X1 _985_ (
    .A(_261_),
    .B(_260_),
    .C(_259_),
    .Y(_262_)
);

NAND3X1 _986_ (
    .A(_246_),
    .B(_258_),
    .C(_262_),
    .Y(_263_)
);

AND2X2 _987_ (
    .A(_241_),
    .B(_245_),
    .Y(_264_)
);

NAND3X1 _988_ (
    .A(_259_),
    .B(_257_),
    .C(_253_),
    .Y(_265_)
);

OAI21X1 _989_ (
    .A(_261_),
    .B(_260_),
    .C(_247_),
    .Y(_266_)
);

NAND3X1 _990_ (
    .A(_265_),
    .B(_264_),
    .C(_266_),
    .Y(_267_)
);

NAND3X1 _991_ (
    .A(_263_),
    .B(_267_),
    .C(_234_),
    .Y(_268_)
);

OAI21X1 _992_ (
    .A(_215_),
    .B(_206_),
    .C(_218_),
    .Y(_269_)
);

NAND2X1 _993_ (
    .A(_263_),
    .B(_267_),
    .Y(_270_)
);

NAND2X1 _994_ (
    .A(_269_),
    .B(_270_),
    .Y(_271_)
);

NAND3X1 _995_ (
    .A(_233_),
    .B(_268_),
    .C(_271_),
    .Y(_272_)
);

NAND3X1 _996_ (
    .A(_263_),
    .B(_267_),
    .C(_269_),
    .Y(_273_)
);

NAND2X1 _997_ (
    .A(_234_),
    .B(_270_),
    .Y(_274_)
);

NAND3X1 _998_ (
    .A(_232_),
    .B(_273_),
    .C(_274_),
    .Y(_275_)
);

NAND2X1 _999_ (
    .A(_272_),
    .B(_275_),
    .Y(_276_)
);

endmodule
