magic
tech scmos
magscale 1 2
timestamp 1771034318
<< metal1 >>
rect -62 12002 30 12018
rect -62 11538 -2 12002
rect 3887 11897 3933 11903
rect 5427 11837 5473 11843
rect 11527 11837 11593 11843
rect 12222 11778 12282 12018
rect 12190 11762 12282 11778
rect 6307 11697 6333 11703
rect 6887 11677 6933 11683
rect 6347 11617 6413 11623
rect 11387 11597 11413 11603
rect -62 11522 30 11538
rect -62 11058 -2 11522
rect 9947 11497 9993 11503
rect 10667 11437 10773 11443
rect 9157 11383 9163 11433
rect 9147 11377 9163 11383
rect 3407 11357 3513 11363
rect 10847 11357 10933 11363
rect 12222 11298 12282 11762
rect 12190 11282 12282 11298
rect 2447 11217 2473 11223
rect 3447 11217 3473 11223
rect 9987 11217 10073 11223
rect 10147 11217 10273 11223
rect 3367 11197 3393 11203
rect 8507 11197 8533 11203
rect -62 11042 30 11058
rect -62 10578 -2 11042
rect 3367 10957 3433 10963
rect 5947 10877 6013 10883
rect 12222 10818 12282 11282
rect 12190 10802 12282 10818
rect 1887 10677 1953 10683
rect -62 10562 30 10578
rect -62 10098 -2 10562
rect 7947 10497 8053 10503
rect 8147 10497 8253 10503
rect 7947 10417 8033 10423
rect 11707 10417 11793 10423
rect 7767 10397 7873 10403
rect 9947 10377 10053 10383
rect 12222 10338 12282 10802
rect 12190 10322 12282 10338
rect 1567 10257 1633 10263
rect 7127 10257 7153 10263
rect 9607 10257 9613 10263
rect 9627 10257 9673 10263
rect 10387 10257 10403 10263
rect 10397 10167 10403 10257
rect 10587 10237 10693 10243
rect -62 10082 30 10098
rect -62 9618 -2 10082
rect 9647 10057 9673 10063
rect 12222 9858 12282 10322
rect 12190 9842 12282 9858
rect 1807 9797 1893 9803
rect 5007 9717 5093 9723
rect -62 9602 30 9618
rect -62 9138 -2 9602
rect 10287 9517 10393 9523
rect 11147 9437 11173 9443
rect 11127 9397 11153 9403
rect 12222 9378 12282 9842
rect 12190 9362 12282 9378
rect 10267 9317 10293 9323
rect 367 9297 453 9303
rect 8007 9297 8053 9303
rect 7927 9277 7943 9283
rect 7937 9203 7943 9277
rect 7927 9197 7943 9203
rect -62 9122 30 9138
rect -62 8658 -2 9122
rect 297 9103 303 9123
rect 267 9097 303 9103
rect 10727 9097 10793 9103
rect 11257 9037 11353 9043
rect 11257 9027 11263 9037
rect 11077 8963 11083 8973
rect 11067 8957 11083 8963
rect 11287 8917 11313 8923
rect 12222 8898 12282 9362
rect 12190 8882 12282 8898
rect 11727 8857 11753 8863
rect 6247 8837 6293 8843
rect 9747 8837 9793 8843
rect 8507 8817 8553 8823
rect 2857 8803 2863 8813
rect 2747 8797 2863 8803
rect 1887 8677 1943 8683
rect -62 8642 30 8658
rect 1937 8657 1943 8677
rect -62 8178 -2 8642
rect 4867 8537 4913 8543
rect 7327 8497 7393 8503
rect 4267 8477 4393 8483
rect 4667 8477 4753 8483
rect 5107 8477 5173 8483
rect 6167 8477 6213 8483
rect 7887 8477 7973 8483
rect 7767 8457 7813 8463
rect 7907 8457 7973 8463
rect 12222 8418 12282 8882
rect 12190 8402 12282 8418
rect 9087 8377 9113 8383
rect 4207 8337 4233 8343
rect 8907 8337 8993 8343
rect 9607 8337 9713 8343
rect 10127 8337 10233 8343
rect 11347 8337 11373 8343
rect 11987 8337 12053 8343
rect 7747 8317 7813 8323
rect 6537 8263 6543 8313
rect 6537 8257 6553 8263
rect 8947 8257 8993 8263
rect 4567 8237 4673 8243
rect -62 8162 30 8178
rect -62 7698 -2 8162
rect 8707 8097 8773 8103
rect 3947 8077 4013 8083
rect 8407 8077 8453 8083
rect 8507 8077 8573 8083
rect 1387 8057 1413 8063
rect 2727 8037 2793 8043
rect 7607 8017 7713 8023
rect 8147 7997 8213 8003
rect 12222 7938 12282 8402
rect 12190 7922 12282 7938
rect 467 7857 493 7863
rect 2567 7857 2653 7863
rect 4667 7857 4713 7863
rect 9147 7857 9193 7863
rect 2667 7797 2713 7803
rect 8767 7757 8873 7763
rect -62 7682 30 7698
rect -62 7218 -2 7682
rect 5627 7617 5693 7623
rect 1687 7537 1733 7543
rect 2227 7537 2333 7543
rect 11267 7537 11353 7543
rect 11747 7537 11813 7543
rect 4867 7517 4913 7523
rect 8727 7497 8773 7503
rect 3367 7477 3393 7483
rect 12222 7458 12282 7922
rect 12190 7442 12282 7458
rect 3807 7417 3853 7423
rect 6807 7397 6893 7403
rect 10447 7377 10533 7383
rect 7787 7357 7853 7363
rect 6687 7317 6753 7323
rect 4187 7257 4233 7263
rect -62 7202 30 7218
rect -62 6738 -2 7202
rect 5807 7157 5833 7163
rect 4947 7097 4973 7103
rect 6377 7103 6383 7113
rect 6377 7097 6453 7103
rect 5877 7083 5883 7093
rect 5867 7077 5883 7083
rect 5687 7057 5713 7063
rect 10547 7057 10593 7063
rect 4407 6997 4493 7003
rect 12222 6978 12282 7442
rect 12190 6962 12282 6978
rect 1927 6917 1953 6923
rect 3887 6917 3933 6923
rect 3307 6897 3333 6903
rect 5407 6897 5513 6903
rect 5627 6857 5643 6863
rect 2487 6837 2513 6843
rect 4607 6837 4693 6843
rect 5637 6843 5643 6857
rect 6807 6857 6853 6863
rect 5637 6837 5733 6843
rect 7507 6837 7553 6843
rect 4847 6817 4893 6823
rect -62 6722 30 6738
rect -62 6258 -2 6722
rect 877 6703 883 6723
rect 787 6697 883 6703
rect 6247 6697 6313 6703
rect 4807 6617 4863 6623
rect 2487 6577 2573 6583
rect 3387 6577 3413 6583
rect 4127 6557 4253 6563
rect 4567 6557 4633 6563
rect 4857 6563 4863 6617
rect 8007 6597 8033 6603
rect 6587 6577 6693 6583
rect 4857 6557 4873 6563
rect 5167 6557 5283 6563
rect 5277 6547 5283 6557
rect 12222 6498 12282 6962
rect 12190 6482 12282 6498
rect 3367 6457 3413 6463
rect 4287 6457 4373 6463
rect 7447 6457 7473 6463
rect 2847 6437 2913 6443
rect 3367 6417 3453 6423
rect 4467 6417 4553 6423
rect 4927 6417 4953 6423
rect 5247 6417 5253 6423
rect 5267 6417 5273 6423
rect 5767 6417 5783 6423
rect 5777 6347 5783 6417
rect 6377 6417 6393 6423
rect 6377 6403 6383 6417
rect 6827 6417 6933 6423
rect 6267 6397 6383 6403
rect 2307 6277 2393 6283
rect -62 6242 30 6258
rect -62 5778 -2 6242
rect 6057 6177 6073 6183
rect 4187 6137 4343 6143
rect 4337 6103 4343 6137
rect 5247 6137 5343 6143
rect 4337 6097 4353 6103
rect 3267 6077 3373 6083
rect 5017 6083 5023 6133
rect 5337 6103 5343 6137
rect 5787 6137 5903 6143
rect 5337 6097 5353 6103
rect 5007 6077 5023 6083
rect 5427 6077 5453 6083
rect 4027 6057 4113 6063
rect 5437 6063 5443 6077
rect 5657 6083 5663 6113
rect 5897 6087 5903 6137
rect 6057 6103 6063 6177
rect 6467 6157 6533 6163
rect 7377 6137 7413 6143
rect 6007 6097 6063 6103
rect 6647 6097 6773 6103
rect 7377 6103 7383 6137
rect 9687 6137 9753 6143
rect 7267 6097 7383 6103
rect 5627 6077 5663 6083
rect 5437 6057 5513 6063
rect 12222 6018 12282 6482
rect 12190 6002 12282 6018
rect 6407 5937 6423 5943
rect 4407 5917 4513 5923
rect 6417 5907 6423 5937
rect 10167 5937 10273 5943
rect 10147 5917 10193 5923
rect 6717 5903 6723 5913
rect 6707 5897 6723 5903
rect 5477 5863 5483 5893
rect 5477 5857 5493 5863
rect -62 5762 30 5778
rect -62 5298 -2 5762
rect 7367 5697 7393 5703
rect 9427 5617 9453 5623
rect 5587 5597 5653 5603
rect 2547 5557 2613 5563
rect 12222 5538 12282 6002
rect 12190 5522 12282 5538
rect 7787 5457 7813 5463
rect 4927 5437 4993 5443
rect 10227 5437 10333 5443
rect 5987 5397 6013 5403
rect 6367 5397 6453 5403
rect 7407 5377 7513 5383
rect -62 5282 30 5298
rect -62 4818 -2 5282
rect 637 5197 653 5203
rect 637 5147 643 5197
rect 6167 5197 6213 5203
rect 8327 5117 8433 5123
rect 12222 5058 12282 5522
rect 12190 5042 12282 5058
rect 1107 4977 1123 4983
rect 1117 4947 1123 4977
rect -62 4802 30 4818
rect -62 4338 -2 4802
rect 8297 4783 8303 4803
rect 8247 4777 8303 4783
rect 5787 4717 5853 4723
rect 8447 4717 8493 4723
rect 12222 4578 12282 5042
rect 12190 4562 12282 4578
rect 2387 4497 2493 4503
rect 1507 4477 1613 4483
rect 4047 4437 4133 4443
rect 6667 4397 6713 4403
rect -62 4322 30 4338
rect -62 3858 -2 4322
rect 7127 4157 7213 4163
rect 12222 4098 12282 4562
rect 12190 4082 12282 4098
rect 11407 3997 11473 4003
rect 5047 3957 5133 3963
rect -62 3842 30 3858
rect -62 3378 -2 3842
rect 9947 3677 9953 3683
rect 9967 3677 10053 3683
rect 3347 3657 3393 3663
rect 12222 3618 12282 4082
rect 12190 3602 12282 3618
rect 5137 3537 5153 3543
rect 947 3517 973 3523
rect 987 3517 1013 3523
rect 5137 3507 5143 3537
rect 10067 3477 10173 3483
rect -62 3362 30 3378
rect -62 2898 -2 3362
rect 9327 3257 9433 3263
rect 12222 3138 12282 3602
rect 12190 3122 12282 3138
rect 10027 3057 10113 3063
rect 10607 3057 10673 3063
rect 307 2917 323 2923
rect -62 2882 30 2898
rect 317 2897 323 2917
rect 4527 2917 4603 2923
rect 4597 2897 4603 2917
rect -62 2418 -2 2882
rect 11687 2857 11713 2863
rect 7387 2717 7413 2723
rect 7447 2717 7493 2723
rect 9027 2697 9053 2703
rect 12222 2658 12282 3122
rect 12190 2642 12282 2658
rect 8867 2597 8933 2603
rect 11207 2577 11273 2583
rect 11477 2577 11493 2583
rect 11367 2557 11383 2563
rect 6607 2517 6713 2523
rect 10567 2517 10633 2523
rect 11377 2523 11383 2557
rect 11477 2547 11483 2577
rect 11377 2517 11413 2523
rect 9087 2497 9193 2503
rect -62 2402 30 2418
rect -62 1938 -2 2402
rect 9327 2337 9393 2343
rect 8547 2297 8633 2303
rect 10507 2297 10593 2303
rect 347 2277 433 2283
rect 6167 2257 6293 2263
rect 8867 2257 8893 2263
rect 12222 2178 12282 2642
rect 12190 2162 12282 2178
rect 6567 2097 6653 2103
rect 7987 2097 8033 2103
rect 8147 2057 8213 2063
rect 9787 2037 9853 2043
rect -62 1922 30 1938
rect -62 1458 -2 1922
rect 8227 1897 8293 1903
rect 7007 1857 7093 1863
rect 5237 1763 5243 1793
rect 9367 1777 9393 1783
rect 11327 1777 11413 1783
rect 5227 1757 5243 1763
rect 7087 1757 7113 1763
rect 9787 1757 9813 1763
rect 7867 1717 7893 1723
rect 11367 1717 11393 1723
rect 12222 1698 12282 2162
rect 12190 1682 12282 1698
rect 6967 1657 7013 1663
rect 8277 1657 8333 1663
rect 8277 1647 8283 1657
rect 6847 1617 6873 1623
rect 7207 1617 7233 1623
rect 8487 1617 8573 1623
rect 6467 1537 6493 1543
rect 7737 1517 7813 1523
rect 7737 1507 7743 1517
rect -62 1442 30 1458
rect -62 978 -2 1442
rect 6767 1277 6793 1283
rect 7897 1283 7903 1353
rect 7927 1337 8013 1343
rect 7917 1297 7953 1303
rect 7917 1287 7923 1297
rect 7847 1277 7903 1283
rect 12222 1218 12282 1682
rect 12190 1202 12282 1218
rect 10027 1137 10043 1143
rect 3167 1117 3273 1123
rect 9607 1117 9623 1123
rect 9617 1043 9623 1117
rect 9807 1117 9933 1123
rect 10037 1107 10043 1137
rect 9607 1037 9623 1043
rect -62 962 30 978
rect -62 498 -2 962
rect 407 857 473 863
rect 2447 857 2573 863
rect 8847 837 8893 843
rect 5227 817 5253 823
rect 12222 738 12282 1202
rect 12190 722 12282 738
rect 6747 637 6773 643
rect 8687 637 8733 643
rect 10947 637 11033 643
rect 7427 597 7453 603
rect -62 482 30 498
rect -62 18 -2 482
rect 4247 337 4273 343
rect 8727 337 8753 343
rect 12222 258 12282 722
rect 12190 242 12282 258
rect 5887 117 5933 123
rect -62 2 30 18
rect 12222 2 12282 242
<< m2contact >>
rect 9493 12013 9507 12027
rect 10033 12013 10047 12027
rect 3873 11893 3887 11907
rect 3933 11893 3947 11907
rect 5413 11833 5427 11847
rect 5473 11833 5487 11847
rect 11513 11833 11527 11847
rect 11593 11833 11607 11847
rect 6293 11693 6307 11707
rect 6333 11693 6347 11707
rect 6873 11673 6887 11687
rect 6933 11673 6947 11687
rect 6333 11613 6347 11627
rect 6413 11613 6427 11627
rect 11373 11593 11387 11607
rect 11413 11593 11427 11607
rect 6473 11513 6487 11527
rect 7113 11513 7127 11527
rect 11613 11513 11627 11527
rect 11753 11513 11767 11527
rect 9933 11493 9947 11507
rect 9993 11493 10007 11507
rect 9153 11433 9167 11447
rect 10653 11433 10667 11447
rect 10773 11433 10787 11447
rect 9133 11373 9147 11387
rect 3393 11353 3407 11367
rect 3513 11353 3527 11367
rect 10833 11353 10847 11367
rect 10933 11353 10947 11367
rect 2433 11213 2447 11227
rect 2473 11213 2487 11227
rect 3433 11213 3447 11227
rect 3473 11213 3487 11227
rect 9973 11213 9987 11227
rect 10073 11213 10087 11227
rect 10133 11213 10147 11227
rect 10273 11213 10287 11227
rect 3353 11193 3367 11207
rect 3393 11193 3407 11207
rect 8493 11193 8507 11207
rect 8533 11193 8547 11207
rect 73 11033 87 11047
rect 6293 11033 6307 11047
rect 7513 11033 7527 11047
rect 11333 11033 11347 11047
rect 3353 10953 3367 10967
rect 3433 10953 3447 10967
rect 5933 10873 5947 10887
rect 6013 10873 6027 10887
rect 1873 10673 1887 10687
rect 1953 10673 1967 10687
rect 73 10553 87 10567
rect 393 10553 407 10567
rect 1633 10553 1647 10567
rect 2033 10553 2047 10567
rect 3613 10553 3627 10567
rect 4833 10553 4847 10567
rect 5893 10553 5907 10567
rect 6033 10553 6047 10567
rect 6673 10553 6687 10567
rect 7273 10553 7287 10567
rect 11713 10553 11727 10567
rect 7933 10493 7947 10507
rect 8053 10493 8067 10507
rect 8133 10493 8147 10507
rect 8253 10493 8267 10507
rect 7933 10413 7947 10427
rect 8033 10413 8047 10427
rect 11693 10413 11707 10427
rect 11793 10413 11807 10427
rect 7753 10393 7767 10407
rect 7873 10393 7887 10407
rect 9933 10373 9947 10387
rect 10053 10373 10067 10387
rect 1553 10253 1567 10267
rect 1633 10253 1647 10267
rect 7113 10253 7127 10267
rect 7153 10253 7167 10267
rect 9593 10253 9607 10267
rect 9613 10253 9627 10267
rect 9673 10253 9687 10267
rect 10373 10253 10387 10267
rect 10573 10233 10587 10247
rect 10693 10233 10707 10247
rect 10393 10153 10407 10167
rect 753 10093 767 10107
rect 5393 10093 5407 10107
rect 6873 10093 6887 10107
rect 2533 10073 2547 10087
rect 2633 10073 2647 10087
rect 3653 10073 3667 10087
rect 4673 10073 4687 10087
rect 4913 10073 4927 10087
rect 5573 10073 5587 10087
rect 6553 10073 6567 10087
rect 9633 10053 9647 10067
rect 9673 10053 9687 10067
rect 1793 9793 1807 9807
rect 1893 9793 1907 9807
rect 4993 9713 5007 9727
rect 5093 9713 5107 9727
rect 3753 9613 3767 9627
rect 953 9593 967 9607
rect 2293 9593 2307 9607
rect 3033 9593 3047 9607
rect 3213 9593 3227 9607
rect 4593 9593 4607 9607
rect 5573 9593 5587 9607
rect 10273 9513 10287 9527
rect 10393 9513 10407 9527
rect 11133 9433 11147 9447
rect 11173 9433 11187 9447
rect 11113 9393 11127 9407
rect 11153 9393 11167 9407
rect 10253 9313 10267 9327
rect 10293 9313 10307 9327
rect 353 9293 367 9307
rect 453 9293 467 9307
rect 7993 9293 8007 9307
rect 8053 9293 8067 9307
rect 7913 9273 7927 9287
rect 7913 9193 7927 9207
rect 253 9093 267 9107
rect 2913 9113 2927 9127
rect 3613 9113 3627 9127
rect 4133 9113 4147 9127
rect 4353 9113 4367 9127
rect 10713 9093 10727 9107
rect 10793 9093 10807 9107
rect 11353 9033 11367 9047
rect 11253 9013 11267 9027
rect 11073 8973 11087 8987
rect 11053 8953 11067 8967
rect 11273 8913 11287 8927
rect 11313 8913 11327 8927
rect 11713 8853 11727 8867
rect 11753 8853 11767 8867
rect 6233 8833 6247 8847
rect 6293 8833 6307 8847
rect 9733 8833 9747 8847
rect 9793 8833 9807 8847
rect 2853 8813 2867 8827
rect 8493 8813 8507 8827
rect 8553 8813 8567 8827
rect 2733 8793 2747 8807
rect 1873 8673 1887 8687
rect 4733 8633 4747 8647
rect 4853 8533 4867 8547
rect 4913 8533 4927 8547
rect 7313 8493 7327 8507
rect 7393 8493 7407 8507
rect 4253 8473 4267 8487
rect 4393 8473 4407 8487
rect 4653 8473 4667 8487
rect 4753 8473 4767 8487
rect 5093 8473 5107 8487
rect 5173 8473 5187 8487
rect 6153 8473 6167 8487
rect 6213 8473 6227 8487
rect 7873 8473 7887 8487
rect 7973 8473 7987 8487
rect 7753 8453 7767 8467
rect 7813 8453 7827 8467
rect 7893 8453 7907 8467
rect 7973 8453 7987 8467
rect 9073 8373 9087 8387
rect 9113 8373 9127 8387
rect 4193 8333 4207 8347
rect 4233 8333 4247 8347
rect 8893 8333 8907 8347
rect 8993 8333 9007 8347
rect 9593 8333 9607 8347
rect 9713 8333 9727 8347
rect 10113 8333 10127 8347
rect 10233 8333 10247 8347
rect 11333 8333 11347 8347
rect 11373 8333 11387 8347
rect 11973 8333 11987 8347
rect 12053 8333 12067 8347
rect 6533 8313 6547 8327
rect 7733 8313 7747 8327
rect 7813 8313 7827 8327
rect 6553 8253 6567 8267
rect 8933 8253 8947 8267
rect 8993 8253 9007 8267
rect 4553 8233 4567 8247
rect 4673 8233 4687 8247
rect 3553 8153 3567 8167
rect 4933 8153 4947 8167
rect 5513 8153 5527 8167
rect 8693 8093 8707 8107
rect 8773 8093 8787 8107
rect 3933 8073 3947 8087
rect 4013 8073 4027 8087
rect 8393 8073 8407 8087
rect 8453 8073 8467 8087
rect 8493 8073 8507 8087
rect 8573 8073 8587 8087
rect 1373 8053 1387 8067
rect 1413 8053 1427 8067
rect 2713 8033 2727 8047
rect 2793 8033 2807 8047
rect 7593 8013 7607 8027
rect 7713 8013 7727 8027
rect 8133 7993 8147 8007
rect 8213 7993 8227 8007
rect 453 7853 467 7867
rect 493 7853 507 7867
rect 2553 7853 2567 7867
rect 2653 7853 2667 7867
rect 4653 7853 4667 7867
rect 4713 7853 4727 7867
rect 9133 7853 9147 7867
rect 9193 7853 9207 7867
rect 2653 7793 2667 7807
rect 2713 7793 2727 7807
rect 8753 7753 8767 7767
rect 8873 7753 8887 7767
rect 433 7673 447 7687
rect 773 7673 787 7687
rect 3773 7673 3787 7687
rect 6093 7673 6107 7687
rect 5613 7613 5627 7627
rect 5693 7613 5707 7627
rect 1673 7533 1687 7547
rect 1733 7533 1747 7547
rect 2213 7533 2227 7547
rect 2333 7533 2347 7547
rect 11253 7533 11267 7547
rect 11353 7533 11367 7547
rect 11733 7533 11747 7547
rect 11813 7533 11827 7547
rect 4853 7513 4867 7527
rect 4913 7513 4927 7527
rect 8713 7493 8727 7507
rect 8773 7493 8787 7507
rect 3353 7473 3367 7487
rect 3393 7473 3407 7487
rect 3793 7413 3807 7427
rect 3853 7413 3867 7427
rect 6793 7393 6807 7407
rect 6893 7393 6907 7407
rect 10433 7373 10447 7387
rect 10533 7373 10547 7387
rect 7773 7353 7787 7367
rect 7853 7353 7867 7367
rect 6673 7313 6687 7327
rect 6753 7313 6767 7327
rect 4173 7253 4187 7267
rect 4233 7253 4247 7267
rect 7513 7213 7527 7227
rect 633 7193 647 7207
rect 1033 7193 1047 7207
rect 1393 7193 1407 7207
rect 1993 7193 2007 7207
rect 6593 7193 6607 7207
rect 5793 7153 5807 7167
rect 5833 7153 5847 7167
rect 6373 7113 6387 7127
rect 4933 7093 4947 7107
rect 4973 7093 4987 7107
rect 5873 7093 5887 7107
rect 6453 7093 6467 7107
rect 5853 7073 5867 7087
rect 5673 7053 5687 7067
rect 5713 7053 5727 7067
rect 10533 7053 10547 7067
rect 10593 7053 10607 7067
rect 4393 6993 4407 7007
rect 4493 6993 4507 7007
rect 1913 6913 1927 6927
rect 1953 6913 1967 6927
rect 3873 6913 3887 6927
rect 3933 6913 3947 6927
rect 3293 6893 3307 6907
rect 3333 6893 3347 6907
rect 5393 6893 5407 6907
rect 5513 6893 5527 6907
rect 5613 6853 5627 6867
rect 2473 6833 2487 6847
rect 2513 6833 2527 6847
rect 4593 6833 4607 6847
rect 4693 6833 4707 6847
rect 6793 6853 6807 6867
rect 6853 6853 6867 6867
rect 5733 6833 5747 6847
rect 7493 6833 7507 6847
rect 7553 6833 7567 6847
rect 4833 6813 4847 6827
rect 4893 6813 4907 6827
rect 773 6693 787 6707
rect 3373 6713 3387 6727
rect 8033 6713 8047 6727
rect 6233 6693 6247 6707
rect 6313 6693 6327 6707
rect 4793 6613 4807 6627
rect 2473 6573 2487 6587
rect 2573 6573 2587 6587
rect 3373 6573 3387 6587
rect 3413 6573 3427 6587
rect 4113 6553 4127 6567
rect 4253 6553 4267 6567
rect 4553 6553 4567 6567
rect 4633 6553 4647 6567
rect 7993 6593 8007 6607
rect 8033 6593 8047 6607
rect 6573 6573 6587 6587
rect 6693 6573 6707 6587
rect 4873 6553 4887 6567
rect 5153 6553 5167 6567
rect 5273 6533 5287 6547
rect 3353 6453 3367 6467
rect 3413 6453 3427 6467
rect 4273 6453 4287 6467
rect 4373 6453 4387 6467
rect 7433 6453 7447 6467
rect 7473 6453 7487 6467
rect 2833 6433 2847 6447
rect 2913 6433 2927 6447
rect 3353 6413 3367 6427
rect 3453 6413 3467 6427
rect 4453 6413 4467 6427
rect 4553 6413 4567 6427
rect 4913 6413 4927 6427
rect 4953 6413 4967 6427
rect 5233 6413 5247 6427
rect 5253 6413 5267 6427
rect 5273 6413 5287 6427
rect 5753 6413 5767 6427
rect 6253 6393 6267 6407
rect 6393 6413 6407 6427
rect 6813 6413 6827 6427
rect 6933 6413 6947 6427
rect 5773 6333 5787 6347
rect 2293 6273 2307 6287
rect 2393 6273 2407 6287
rect 2393 6253 2407 6267
rect 973 6233 987 6247
rect 1853 6233 1867 6247
rect 1913 6233 1927 6247
rect 2933 6233 2947 6247
rect 8753 6233 8767 6247
rect 4173 6133 4187 6147
rect 5013 6133 5027 6147
rect 5233 6133 5247 6147
rect 4353 6093 4367 6107
rect 3253 6073 3267 6087
rect 3373 6073 3387 6087
rect 4993 6073 5007 6087
rect 5773 6133 5787 6147
rect 5653 6113 5667 6127
rect 5353 6093 5367 6107
rect 5413 6073 5427 6087
rect 4013 6053 4027 6067
rect 4113 6053 4127 6067
rect 5453 6073 5467 6087
rect 5613 6073 5627 6087
rect 5993 6093 6007 6107
rect 6073 6173 6087 6187
rect 6453 6153 6467 6167
rect 6533 6153 6547 6167
rect 6633 6093 6647 6107
rect 6773 6093 6787 6107
rect 7253 6093 7267 6107
rect 7413 6133 7427 6147
rect 9673 6133 9687 6147
rect 9753 6133 9767 6147
rect 5893 6073 5907 6087
rect 5513 6053 5527 6067
rect 6393 5933 6407 5947
rect 4393 5913 4407 5927
rect 4513 5913 4527 5927
rect 10153 5933 10167 5947
rect 10273 5933 10287 5947
rect 6713 5913 6727 5927
rect 10133 5913 10147 5927
rect 10193 5913 10207 5927
rect 5473 5893 5487 5907
rect 6413 5893 6427 5907
rect 6693 5893 6707 5907
rect 5493 5853 5507 5867
rect 293 5773 307 5787
rect 8493 5753 8507 5767
rect 7353 5693 7367 5707
rect 7393 5693 7407 5707
rect 9413 5613 9427 5627
rect 9453 5613 9467 5627
rect 5573 5593 5587 5607
rect 5653 5593 5667 5607
rect 2533 5553 2547 5567
rect 2613 5553 2627 5567
rect 7773 5453 7787 5467
rect 7813 5453 7827 5467
rect 4913 5433 4927 5447
rect 4993 5433 5007 5447
rect 10213 5433 10227 5447
rect 10333 5433 10347 5447
rect 5973 5393 5987 5407
rect 6013 5393 6027 5407
rect 6353 5393 6367 5407
rect 6453 5393 6467 5407
rect 7393 5373 7407 5387
rect 7513 5373 7527 5387
rect 7893 5293 7907 5307
rect 433 5273 447 5287
rect 633 5273 647 5287
rect 1213 5273 1227 5287
rect 1413 5273 1427 5287
rect 2253 5273 2267 5287
rect 3353 5273 3367 5287
rect 653 5193 667 5207
rect 6153 5193 6167 5207
rect 6213 5193 6227 5207
rect 633 5133 647 5147
rect 8313 5113 8327 5127
rect 8433 5113 8447 5127
rect 1093 4973 1107 4987
rect 1113 4933 1127 4947
rect 7413 4813 7427 4827
rect 2073 4793 2087 4807
rect 3053 4793 3067 4807
rect 8093 4793 8107 4807
rect 8233 4773 8247 4787
rect 8813 4793 8827 4807
rect 8833 4793 8847 4807
rect 9533 4793 9547 4807
rect 5773 4713 5787 4727
rect 5853 4713 5867 4727
rect 8433 4713 8447 4727
rect 8493 4713 8507 4727
rect 2373 4493 2387 4507
rect 2493 4493 2507 4507
rect 1493 4473 1507 4487
rect 1613 4473 1627 4487
rect 4033 4433 4047 4447
rect 4133 4433 4147 4447
rect 6653 4393 6667 4407
rect 6713 4393 6727 4407
rect 73 4313 87 4327
rect 93 4313 107 4327
rect 453 4313 467 4327
rect 1113 4313 1127 4327
rect 1673 4313 1687 4327
rect 2913 4313 2927 4327
rect 3573 4313 3587 4327
rect 4233 4313 4247 4327
rect 4313 4313 4327 4327
rect 5153 4313 5167 4327
rect 8213 4313 8227 4327
rect 9873 4313 9887 4327
rect 10053 4313 10067 4327
rect 7113 4153 7127 4167
rect 7213 4153 7227 4167
rect 11393 3993 11407 4007
rect 11473 3993 11487 4007
rect 5033 3953 5047 3967
rect 5133 3953 5147 3967
rect 73 3833 87 3847
rect 873 3833 887 3847
rect 1473 3833 1487 3847
rect 2133 3833 2147 3847
rect 2353 3833 2367 3847
rect 3173 3833 3187 3847
rect 3633 3833 3647 3847
rect 4113 3833 4127 3847
rect 4753 3833 4767 3847
rect 8833 3833 8847 3847
rect 9933 3673 9947 3687
rect 9953 3673 9967 3687
rect 10053 3673 10067 3687
rect 3333 3653 3347 3667
rect 3393 3653 3407 3667
rect 933 3513 947 3527
rect 973 3513 987 3527
rect 1013 3513 1027 3527
rect 5153 3533 5167 3547
rect 5133 3493 5147 3507
rect 10053 3473 10067 3487
rect 10173 3473 10187 3487
rect 793 3373 807 3387
rect 1053 3353 1067 3367
rect 1893 3353 1907 3367
rect 5773 3353 5787 3367
rect 6993 3353 7007 3367
rect 7713 3353 7727 3367
rect 9313 3253 9327 3267
rect 9433 3253 9447 3267
rect 10013 3053 10027 3067
rect 10113 3053 10127 3067
rect 10593 3053 10607 3067
rect 10673 3053 10687 3067
rect 293 2913 307 2927
rect 4513 2913 4527 2927
rect 1153 2893 1167 2907
rect 493 2873 507 2887
rect 513 2873 527 2887
rect 2773 2873 2787 2887
rect 2953 2873 2967 2887
rect 4873 2873 4887 2887
rect 5273 2873 5287 2887
rect 5313 2873 5327 2887
rect 5433 2873 5447 2887
rect 11673 2853 11687 2867
rect 11713 2853 11727 2867
rect 7373 2713 7387 2727
rect 7413 2713 7427 2727
rect 7433 2713 7447 2727
rect 7493 2713 7507 2727
rect 9013 2693 9027 2707
rect 9053 2693 9067 2707
rect 8853 2593 8867 2607
rect 8933 2593 8947 2607
rect 11193 2573 11207 2587
rect 11273 2573 11287 2587
rect 11353 2553 11367 2567
rect 6593 2513 6607 2527
rect 6713 2513 6727 2527
rect 10553 2513 10567 2527
rect 10633 2513 10647 2527
rect 11493 2573 11507 2587
rect 11473 2533 11487 2547
rect 11413 2513 11427 2527
rect 9073 2493 9087 2507
rect 9193 2493 9207 2507
rect 1193 2393 1207 2407
rect 1693 2393 1707 2407
rect 3033 2393 3047 2407
rect 3993 2393 4007 2407
rect 4973 2393 4987 2407
rect 9313 2333 9327 2347
rect 9393 2333 9407 2347
rect 8533 2293 8547 2307
rect 8633 2293 8647 2307
rect 10493 2293 10507 2307
rect 10593 2293 10607 2307
rect 333 2273 347 2287
rect 433 2273 447 2287
rect 6153 2253 6167 2267
rect 6293 2253 6307 2267
rect 8853 2253 8867 2267
rect 8893 2253 8907 2267
rect 6553 2093 6567 2107
rect 6653 2093 6667 2107
rect 7973 2093 7987 2107
rect 8033 2093 8047 2107
rect 8133 2053 8147 2067
rect 8213 2053 8227 2067
rect 9773 2033 9787 2047
rect 9853 2033 9867 2047
rect 2373 1933 2387 1947
rect 253 1913 267 1927
rect 1573 1913 1587 1927
rect 2913 1913 2927 1927
rect 2933 1913 2947 1927
rect 8213 1893 8227 1907
rect 8293 1893 8307 1907
rect 6993 1853 7007 1867
rect 7093 1853 7107 1867
rect 5233 1793 5247 1807
rect 5213 1753 5227 1767
rect 9353 1773 9367 1787
rect 9393 1773 9407 1787
rect 11313 1773 11327 1787
rect 11413 1773 11427 1787
rect 7073 1753 7087 1767
rect 7113 1753 7127 1767
rect 9773 1753 9787 1767
rect 9813 1753 9827 1767
rect 7853 1713 7867 1727
rect 7893 1713 7907 1727
rect 11353 1713 11367 1727
rect 11393 1713 11407 1727
rect 6953 1653 6967 1667
rect 7013 1653 7027 1667
rect 8333 1653 8347 1667
rect 8273 1633 8287 1647
rect 6833 1613 6847 1627
rect 6873 1613 6887 1627
rect 7193 1613 7207 1627
rect 7233 1613 7247 1627
rect 8473 1613 8487 1627
rect 8573 1613 8587 1627
rect 6453 1533 6467 1547
rect 6493 1533 6507 1547
rect 7813 1513 7827 1527
rect 7733 1493 7747 1507
rect 493 1433 507 1447
rect 793 1433 807 1447
rect 7893 1353 7907 1367
rect 6753 1273 6767 1287
rect 6793 1273 6807 1287
rect 7833 1273 7847 1287
rect 7913 1333 7927 1347
rect 8013 1333 8027 1347
rect 7953 1293 7967 1307
rect 7913 1273 7927 1287
rect 10013 1133 10027 1147
rect 3153 1113 3167 1127
rect 3273 1113 3287 1127
rect 9593 1113 9607 1127
rect 9593 1033 9607 1047
rect 9793 1113 9807 1127
rect 9933 1113 9947 1127
rect 10033 1093 10047 1107
rect 1473 953 1487 967
rect 1553 953 1567 967
rect 393 853 407 867
rect 473 853 487 867
rect 2433 853 2447 867
rect 2573 853 2587 867
rect 8833 833 8847 847
rect 8893 833 8907 847
rect 5213 813 5227 827
rect 5253 813 5267 827
rect 6733 633 6747 647
rect 6773 633 6787 647
rect 8673 633 8687 647
rect 8733 633 8747 647
rect 10933 633 10947 647
rect 11033 633 11047 647
rect 7413 593 7427 607
rect 7453 593 7467 607
rect 113 493 127 507
rect 673 473 687 487
rect 753 473 767 487
rect 953 473 967 487
rect 1713 473 1727 487
rect 2553 473 2567 487
rect 4233 333 4247 347
rect 4273 333 4287 347
rect 8713 333 8727 347
rect 8753 333 8767 347
rect 5873 113 5887 127
rect 5933 113 5947 127
<< metal2 >>
rect 1256 12023 1263 12063
rect 5996 12027 6003 12063
rect 1236 12016 1263 12023
rect 196 11876 203 11913
rect 96 11676 103 11853
rect 256 11847 263 11873
rect 296 11863 303 11893
rect 296 11856 323 11863
rect 176 11827 183 11843
rect 316 11687 323 11856
rect 356 11827 363 11853
rect 156 11383 163 11653
rect 136 11376 163 11383
rect 216 11376 223 11413
rect 136 11207 143 11376
rect 356 11367 363 11813
rect 496 11663 503 12013
rect 736 11876 743 11913
rect 716 11727 723 11863
rect 756 11847 763 11863
rect 796 11847 803 11893
rect 636 11676 643 11693
rect 776 11683 783 11813
rect 796 11687 803 11833
rect 756 11676 783 11683
rect 496 11656 523 11663
rect 796 11423 803 11673
rect 796 11416 823 11423
rect 636 11383 643 11413
rect 576 11367 583 11383
rect 616 11376 643 11383
rect 776 11367 783 11403
rect 816 11387 823 11416
rect 96 11196 123 11203
rect 76 10696 83 11033
rect 116 10903 123 11196
rect 156 10916 163 11213
rect 216 11187 223 11203
rect 416 11203 423 11353
rect 396 11196 423 11203
rect 196 10916 203 11073
rect 236 10907 243 11193
rect 376 10936 383 10973
rect 416 10947 423 11196
rect 816 11203 823 11373
rect 796 11196 823 11203
rect 116 10896 143 10903
rect 176 10736 203 10743
rect 36 10676 63 10683
rect 56 10487 63 10676
rect 56 10203 63 10473
rect 76 10216 83 10553
rect 176 10547 183 10736
rect 376 10727 383 10893
rect 416 10887 423 10933
rect 556 10916 563 10933
rect 596 10927 603 11163
rect 776 11087 783 11183
rect 736 10916 743 10933
rect 376 10696 383 10713
rect 116 10467 123 10533
rect 156 10456 183 10463
rect 176 10407 183 10456
rect 276 10423 283 10453
rect 396 10447 403 10553
rect 276 10416 303 10423
rect 336 10347 343 10423
rect 376 10407 383 10423
rect 196 10256 203 10333
rect 36 10196 63 10203
rect 36 9983 43 10196
rect 36 9976 63 9983
rect 56 9947 63 9976
rect 396 9963 403 10213
rect 416 10207 423 10873
rect 536 10867 543 10903
rect 576 10887 583 10903
rect 576 10716 583 10853
rect 436 10487 443 10513
rect 436 10456 443 10473
rect 456 10467 463 10703
rect 436 10007 443 10393
rect 496 10227 503 10713
rect 716 10707 723 10873
rect 776 10507 783 11073
rect 816 10927 823 11196
rect 836 10487 843 11393
rect 876 11263 883 11913
rect 1096 11896 1123 11903
rect 916 11763 923 11843
rect 936 11827 943 11863
rect 896 11756 923 11763
rect 896 11667 903 11756
rect 956 11696 963 11853
rect 1116 11827 1123 11896
rect 916 11676 923 11693
rect 1156 11656 1163 11873
rect 976 11367 983 11403
rect 996 11387 1003 11433
rect 876 11256 903 11263
rect 796 10443 803 10453
rect 776 10436 803 10443
rect 456 9983 463 10223
rect 456 9976 483 9983
rect 376 9956 403 9963
rect 196 9783 203 9923
rect 176 9776 203 9783
rect 156 9756 163 9773
rect 76 9647 83 9753
rect 16 2987 23 6413
rect 36 6116 63 6123
rect 56 5867 63 6116
rect 36 5127 43 5423
rect 76 4647 83 9633
rect 176 9467 183 9776
rect 336 9756 343 9773
rect 216 9496 223 9593
rect 116 9283 123 9453
rect 156 9307 163 9463
rect 96 9276 123 9283
rect 96 6927 103 9276
rect 136 9043 143 9243
rect 116 9036 143 9043
rect 116 8987 123 9036
rect 176 9027 183 9243
rect 256 9107 263 9483
rect 356 9307 363 9773
rect 376 9756 383 9933
rect 396 9767 403 9956
rect 436 9956 463 9963
rect 436 9587 443 9956
rect 476 9927 483 9976
rect 576 9787 583 10033
rect 596 9987 603 10403
rect 796 10236 803 10313
rect 836 10247 843 10433
rect 676 10203 683 10233
rect 616 10067 623 10203
rect 656 10196 683 10203
rect 736 10096 753 10103
rect 616 9956 623 9993
rect 636 9847 643 9913
rect 516 9756 543 9763
rect 576 9756 583 9773
rect 516 9607 523 9756
rect 596 9487 603 9753
rect 616 9747 623 9763
rect 656 9747 663 10053
rect 736 9967 743 10096
rect 696 9767 703 9813
rect 756 9747 763 9943
rect 776 9916 803 9923
rect 796 9727 803 9916
rect 816 9747 823 10223
rect 636 9476 663 9483
rect 376 9287 383 9443
rect 656 9387 663 9476
rect 396 9247 403 9293
rect 136 8963 143 9003
rect 136 8956 163 8963
rect 156 8827 163 8956
rect 236 8927 243 8993
rect 136 8747 143 8783
rect 236 8567 243 8913
rect 256 8767 263 9013
rect 356 8947 363 8963
rect 116 8536 123 8553
rect 156 8467 163 8533
rect 176 8427 183 8523
rect 276 8507 283 8813
rect 356 8776 363 8933
rect 116 8316 143 8323
rect 116 7847 123 8316
rect 136 8056 143 8073
rect 216 8047 223 8453
rect 236 8067 243 8413
rect 316 8327 323 8333
rect 316 8283 323 8313
rect 356 8296 363 8313
rect 316 8276 343 8283
rect 156 7847 163 8043
rect 116 7816 123 7833
rect 176 7707 183 7803
rect 156 7556 163 7613
rect 116 7356 143 7363
rect 116 7327 123 7356
rect 216 7363 223 7693
rect 236 7527 243 7793
rect 196 7356 223 7363
rect 176 7323 183 7353
rect 216 7347 223 7356
rect 156 7316 183 7323
rect 156 7107 163 7316
rect 256 7307 263 8073
rect 336 8047 343 8073
rect 396 8067 403 9053
rect 416 8007 423 8353
rect 396 7887 403 7993
rect 396 7836 403 7873
rect 367 7816 383 7823
rect 376 7567 383 7816
rect 436 7687 443 8043
rect 456 7867 463 9293
rect 556 9276 563 9293
rect 656 9276 683 9283
rect 716 9276 723 9313
rect 776 9307 783 9463
rect 836 9307 843 9483
rect 876 9367 883 10473
rect 896 9347 903 11256
rect 936 11196 943 11233
rect 996 11196 1023 11203
rect 1016 11147 1023 11196
rect 916 10907 923 10923
rect 956 10916 963 10973
rect 996 10903 1003 10913
rect 1016 10907 1023 11133
rect 1076 11007 1083 11653
rect 1116 11416 1143 11423
rect 1176 11416 1203 11423
rect 1116 11367 1123 11416
rect 1196 11387 1203 11416
rect 1116 11207 1123 11353
rect 1096 10943 1103 11153
rect 1176 11147 1183 11163
rect 1076 10936 1103 10943
rect 1136 10936 1143 11053
rect 1216 11027 1223 12013
rect 1236 11847 1243 12016
rect 1436 11896 1463 11903
rect 976 10896 1003 10903
rect 976 10707 983 10896
rect 1036 10807 1043 10933
rect 976 10447 983 10693
rect 1016 10467 1023 10703
rect 1036 10447 1043 10793
rect 1016 10283 1023 10403
rect 1016 10276 1043 10283
rect 936 9963 943 10213
rect 976 9983 983 10193
rect 976 9976 1003 9983
rect 996 9967 1003 9976
rect 936 9956 963 9963
rect 916 9787 923 9953
rect 1036 9947 1043 10276
rect 1056 10227 1063 10423
rect 1076 10267 1083 10936
rect 1156 10927 1163 10953
rect 1176 10703 1183 11013
rect 1156 10696 1183 10703
rect 1176 10487 1183 10696
rect 1176 10443 1183 10453
rect 1116 10436 1143 10443
rect 1176 10436 1203 10443
rect 976 9887 983 9943
rect 1096 9927 1103 10433
rect 1136 10307 1143 10436
rect 1196 10287 1203 10436
rect 1176 10236 1183 10253
rect 1156 10207 1163 10223
rect 1136 9956 1163 9963
rect 1136 9947 1143 9956
rect 996 9787 1003 9793
rect 1116 9756 1123 9873
rect 1156 9756 1163 9813
rect 1176 9767 1183 9923
rect 1216 9887 1223 10993
rect 1236 10767 1243 11193
rect 1256 11187 1263 11773
rect 1276 11647 1283 11673
rect 1336 11656 1343 11693
rect 1276 11187 1283 11633
rect 1356 11623 1363 11633
rect 1336 11616 1363 11623
rect 1336 11387 1343 11616
rect 1316 11227 1323 11373
rect 1356 11347 1363 11383
rect 1356 11176 1363 11213
rect 1276 10936 1283 11133
rect 1316 10716 1323 10733
rect 1376 10347 1383 10403
rect 1336 10256 1343 10293
rect 1296 9963 1303 9993
rect 1396 9967 1403 11873
rect 1456 11427 1463 11896
rect 1476 11827 1483 11863
rect 1476 11447 1483 11813
rect 1516 11676 1523 11933
rect 1676 11863 1683 11933
rect 1856 11876 1883 11883
rect 1656 11856 1683 11863
rect 1556 11676 1583 11683
rect 1516 11383 1523 11413
rect 1496 11376 1523 11383
rect 1536 11347 1543 11383
rect 1576 11367 1583 11676
rect 1596 11667 1603 11713
rect 1616 11347 1623 11853
rect 1696 11656 1703 11713
rect 1516 11196 1523 11273
rect 1556 11196 1563 11313
rect 1476 11087 1483 11193
rect 1476 10916 1483 11013
rect 1436 10716 1443 10733
rect 1516 10327 1523 10753
rect 1536 10456 1543 10513
rect 1516 10243 1523 10313
rect 1496 10236 1523 10243
rect 1496 10203 1503 10236
rect 1536 10216 1543 10313
rect 1556 10267 1563 10933
rect 1496 10196 1523 10203
rect 1296 9956 1323 9963
rect 976 9727 983 9743
rect 956 9447 963 9593
rect 976 9476 983 9573
rect 536 9247 543 9263
rect 516 8943 523 8983
rect 536 8967 543 9033
rect 496 8936 523 8943
rect 496 8787 503 8936
rect 556 8796 563 8813
rect 476 8467 483 8523
rect 576 8487 583 8773
rect 596 8507 603 9233
rect 656 9027 663 9276
rect 736 9267 743 9293
rect 916 9276 923 9293
rect 696 9047 703 9263
rect 896 9027 903 9263
rect 656 8947 663 8983
rect 696 8927 703 8983
rect 796 8816 803 8833
rect 636 8367 643 8793
rect 716 8536 743 8543
rect 636 8316 643 8353
rect 476 7827 483 7853
rect 336 7547 343 7563
rect 356 7467 363 7543
rect 396 7527 403 7533
rect 176 6907 183 7053
rect 176 6856 183 6893
rect 196 6847 203 7073
rect 276 7067 283 7333
rect 336 7087 343 7293
rect 296 7056 323 7063
rect 116 6596 123 6843
rect 156 6596 163 6613
rect 136 6447 143 6563
rect 176 6396 183 6413
rect 296 6396 303 7056
rect 356 7047 363 7063
rect 336 6867 343 6873
rect 376 6856 403 6863
rect 316 6427 323 6843
rect 396 6647 403 6856
rect 416 6623 423 7613
rect 407 6616 423 6623
rect 396 6596 403 6613
rect 376 6507 383 6583
rect 416 6567 423 6583
rect 116 5647 123 6123
rect 296 5927 303 6083
rect 316 5947 323 6393
rect 176 5867 183 5883
rect 416 5787 423 6123
rect 436 5927 443 6613
rect 456 6167 463 7573
rect 476 6887 483 7793
rect 496 7587 503 7853
rect 536 7807 543 8303
rect 656 8267 663 8513
rect 696 8147 703 8493
rect 736 8427 743 8536
rect 756 8307 763 8813
rect 776 8796 783 8813
rect 836 8487 843 9013
rect 856 8847 863 9003
rect 876 8967 883 8983
rect 916 8887 923 8983
rect 936 8927 943 8993
rect 876 8767 883 8793
rect 916 8787 923 8873
rect 936 8796 943 8913
rect 996 8776 1003 8973
rect 776 8287 783 8433
rect 796 8316 803 8413
rect 1016 8347 1023 9733
rect 1276 9727 1283 9953
rect 1296 9707 1303 9956
rect 1336 9927 1343 9943
rect 1336 9607 1343 9913
rect 1376 9867 1383 9943
rect 1416 9767 1423 9953
rect 1436 9883 1443 10193
rect 1516 9907 1523 9943
rect 1436 9876 1463 9883
rect 1376 9707 1383 9723
rect 1056 9503 1063 9593
rect 1056 9496 1083 9503
rect 1036 8627 1043 9333
rect 1076 9067 1083 9496
rect 1096 9447 1103 9483
rect 1116 9296 1123 9373
rect 1096 9247 1103 9263
rect 1076 9047 1083 9053
rect 1056 8967 1063 8983
rect 1056 8547 1063 8813
rect 1076 8807 1083 8963
rect 1096 8547 1103 8973
rect 1116 8503 1123 8773
rect 856 8316 883 8323
rect 876 8247 883 8316
rect 1016 8247 1023 8283
rect 576 7807 583 7873
rect 616 7847 623 7873
rect 676 7836 683 7853
rect 616 7816 623 7833
rect 596 7587 603 7813
rect 656 7807 663 7823
rect 696 7803 703 8053
rect 736 7927 743 8043
rect 816 8036 843 8043
rect 776 7867 783 7973
rect 836 7907 843 8036
rect 756 7816 783 7823
rect 696 7796 723 7803
rect 496 7523 503 7553
rect 496 7516 523 7523
rect 656 7407 663 7793
rect 716 7647 723 7796
rect 776 7687 783 7816
rect 676 7527 683 7563
rect 576 7356 583 7373
rect 676 7367 683 7513
rect 556 7327 563 7343
rect 596 7127 603 7343
rect 636 7207 643 7333
rect 536 7047 543 7063
rect 516 7003 523 7043
rect 536 7027 543 7033
rect 516 6996 543 7003
rect 536 6856 543 6996
rect 676 6987 683 7353
rect 516 6723 523 6843
rect 556 6836 563 6893
rect 496 6716 523 6723
rect 496 6587 503 6716
rect 516 6587 523 6653
rect 536 6547 543 6813
rect 576 6547 583 6563
rect 496 6383 503 6433
rect 536 6416 543 6533
rect 496 6376 523 6383
rect 536 6143 543 6353
rect 527 6136 543 6143
rect 536 5967 543 6136
rect 476 5936 503 5943
rect 436 5887 443 5913
rect 476 5867 483 5936
rect 307 5776 313 5783
rect 136 5636 143 5653
rect 316 5647 323 5773
rect 536 5747 543 5953
rect 576 5907 583 6513
rect 656 6383 663 6893
rect 696 6876 703 6913
rect 716 6847 723 7393
rect 796 7327 803 7633
rect 856 7447 863 8133
rect 876 7507 883 7813
rect 1036 7727 1043 8033
rect 1056 8027 1063 8503
rect 1096 8496 1123 8503
rect 1096 8007 1103 8033
rect 1056 7823 1063 7913
rect 1096 7827 1103 7993
rect 1056 7816 1083 7823
rect 936 7556 943 7713
rect 1076 7683 1083 7816
rect 1056 7676 1083 7683
rect 916 7507 923 7543
rect 956 7527 963 7543
rect 756 7076 763 7093
rect 736 6876 743 6973
rect 796 6867 803 7063
rect 696 6547 703 6633
rect 716 6567 723 6583
rect 696 6416 703 6533
rect 716 6387 723 6553
rect 656 6376 683 6383
rect 776 6376 783 6693
rect 656 5927 663 6153
rect 836 6123 843 6253
rect 836 6116 863 6123
rect 336 5656 343 5733
rect 116 5416 123 5633
rect 296 5456 323 5463
rect 316 5207 323 5456
rect 256 5167 263 5193
rect 296 5156 303 5173
rect 176 4956 183 5053
rect 116 4683 123 4933
rect 116 4676 143 4683
rect 176 4676 183 4893
rect 156 4627 163 4663
rect 296 4663 303 4913
rect 336 4907 343 4923
rect 296 4656 323 4663
rect 76 4456 103 4463
rect 56 3967 63 4433
rect 96 4327 103 4456
rect 76 3976 83 4313
rect 176 4307 183 4633
rect 196 4496 203 4613
rect 336 4427 343 4643
rect 36 3956 53 3963
rect 56 3483 63 3953
rect 76 3496 83 3833
rect 36 3476 63 3483
rect 36 3267 43 3476
rect 16 2247 23 2973
rect 76 2927 83 3243
rect 96 2847 103 4293
rect 176 3907 183 4183
rect 196 4016 203 4113
rect 296 4087 303 4293
rect 336 4196 343 4353
rect 356 4287 363 4653
rect 396 4463 403 5613
rect 416 5416 443 5423
rect 436 5287 443 5416
rect 476 5403 483 5733
rect 496 5587 503 5603
rect 456 5396 483 5403
rect 636 5303 643 5653
rect 656 5443 663 5853
rect 676 5683 683 6083
rect 696 5916 703 5953
rect 676 5676 703 5683
rect 676 5627 683 5643
rect 696 5447 703 5676
rect 656 5436 683 5443
rect 616 5296 643 5303
rect 456 5176 483 5183
rect 456 5147 463 5176
rect 376 4456 403 4463
rect 376 4367 383 4413
rect 396 4307 403 4456
rect 316 4127 323 4183
rect 396 4167 403 4273
rect 356 3847 363 4153
rect 376 4007 383 4073
rect 376 3976 383 3993
rect 316 3707 323 3723
rect 116 3027 123 3053
rect 136 3036 143 3153
rect 176 3087 183 3703
rect 396 3703 403 3833
rect 336 3627 343 3703
rect 376 3696 403 3703
rect 416 3667 423 3713
rect 196 3536 203 3613
rect 436 3543 443 5053
rect 456 4927 463 5133
rect 476 4956 483 5113
rect 456 4867 463 4913
rect 456 4187 463 4313
rect 476 4163 483 4913
rect 496 4507 503 4943
rect 536 4927 543 4943
rect 536 4467 543 4633
rect 576 4567 583 5173
rect 596 4527 603 5173
rect 596 4476 603 4513
rect 576 4447 583 4473
rect 476 4156 503 4163
rect 416 3536 443 3543
rect 396 3247 403 3493
rect 376 3236 393 3243
rect 196 3167 203 3203
rect 196 3063 203 3133
rect 176 3056 203 3063
rect 36 2347 43 2833
rect 176 2567 183 2743
rect 196 2736 223 2743
rect 36 1587 43 2333
rect 196 2327 203 2736
rect 256 2543 263 3093
rect 287 2916 293 2923
rect 316 2743 323 3073
rect 336 3047 343 3113
rect 296 2587 303 2743
rect 316 2736 343 2743
rect 296 2547 303 2573
rect 396 2567 403 2873
rect 416 2567 423 3536
rect 436 3243 443 3513
rect 476 3507 483 3993
rect 496 3987 503 4156
rect 516 3807 523 3953
rect 536 3747 543 4233
rect 576 4216 583 4433
rect 616 4247 623 5296
rect 636 5167 643 5273
rect 656 5207 663 5213
rect 676 5183 683 5436
rect 716 5187 723 5913
rect 656 5176 683 5183
rect 636 5127 643 5133
rect 656 4307 663 5176
rect 676 5107 683 5143
rect 676 4967 683 5033
rect 716 4956 723 4973
rect 676 4696 683 4953
rect 696 4907 703 4943
rect 696 4667 703 4683
rect 616 4187 623 4203
rect 556 3976 563 4173
rect 716 4087 723 4293
rect 736 4207 743 5873
rect 756 5636 783 5643
rect 776 5607 783 5636
rect 836 5627 843 6116
rect 856 5667 863 5893
rect 836 5467 843 5613
rect 756 5176 763 5293
rect 776 5087 783 5393
rect 796 5207 803 5423
rect 856 5423 863 5633
rect 876 5627 883 7213
rect 936 7076 943 7093
rect 936 6903 943 6953
rect 916 6896 943 6903
rect 936 6867 943 6896
rect 976 6587 983 7653
rect 996 7576 1003 7633
rect 996 7336 1003 7493
rect 1036 7207 1043 7563
rect 1056 7507 1063 7676
rect 1116 7663 1123 8333
rect 1136 8167 1143 9353
rect 1156 9267 1163 9293
rect 1156 8787 1163 9253
rect 1176 8967 1183 9273
rect 1196 9247 1203 9573
rect 1436 9487 1443 9813
rect 1216 9287 1223 9443
rect 1276 9087 1283 9243
rect 1236 8847 1243 8983
rect 1276 8967 1283 8983
rect 1296 8943 1303 9253
rect 1276 8936 1303 8943
rect 1176 8796 1183 8813
rect 1236 8787 1243 8833
rect 1176 8323 1183 8533
rect 1236 8516 1243 8553
rect 1276 8516 1283 8936
rect 1316 8647 1323 9373
rect 1376 8987 1383 9453
rect 1436 9447 1443 9473
rect 1456 9347 1463 9876
rect 1436 9256 1443 9313
rect 1496 9276 1503 9293
rect 1516 9003 1523 9873
rect 1536 9367 1543 9953
rect 1576 9903 1583 10973
rect 1596 10307 1603 11333
rect 1676 11176 1683 11363
rect 1696 11347 1703 11383
rect 1696 11207 1703 11213
rect 1616 10903 1623 11093
rect 1656 11027 1663 11173
rect 1696 11156 1703 11193
rect 1756 11047 1763 11193
rect 1776 11167 1783 11193
rect 1696 10903 1703 10993
rect 1796 10987 1803 11863
rect 1876 11703 1883 11876
rect 1876 11696 1903 11703
rect 1856 11676 1883 11683
rect 1856 11607 1863 11676
rect 1876 11427 1883 11433
rect 1916 11383 1923 11573
rect 1836 11367 1843 11383
rect 1896 11376 1923 11383
rect 1836 11067 1843 11313
rect 1856 11176 1883 11183
rect 1856 11147 1863 11176
rect 1896 11156 1903 11253
rect 1616 10896 1643 10903
rect 1676 10896 1703 10903
rect 1616 10887 1623 10896
rect 1636 10716 1643 10753
rect 1696 10716 1703 10853
rect 1636 10447 1643 10553
rect 1676 10423 1683 10673
rect 1676 10416 1703 10423
rect 1596 10207 1603 10253
rect 1596 9967 1603 10193
rect 1556 9896 1583 9903
rect 1556 9707 1563 9896
rect 1616 9843 1623 10293
rect 1676 10267 1683 10416
rect 1636 9927 1643 10253
rect 1716 10236 1723 10333
rect 1736 10307 1743 10423
rect 1756 10236 1763 10973
rect 1836 10943 1843 11053
rect 1956 10963 1963 11693
rect 1976 11427 1983 11813
rect 1996 11487 2003 11883
rect 2036 11876 2043 11893
rect 2156 11876 2183 11883
rect 2056 11787 2063 11863
rect 2016 11676 2043 11683
rect 2096 11676 2123 11683
rect 2016 11667 2023 11676
rect 1996 11067 2003 11473
rect 2076 11447 2083 11633
rect 2116 11467 2123 11676
rect 2076 11416 2083 11433
rect 2096 11156 2103 11293
rect 2116 11287 2123 11453
rect 2136 11387 2143 11713
rect 2156 11647 2163 11876
rect 2256 11863 2263 11913
rect 2236 11856 2263 11863
rect 2376 11896 2403 11903
rect 2196 11827 2203 11843
rect 2376 11827 2383 11896
rect 2567 11896 2583 11903
rect 2616 11896 2623 11913
rect 2936 11896 2943 11913
rect 3816 11907 3823 11913
rect 3616 11896 3643 11903
rect 3676 11896 3693 11903
rect 2176 11627 2183 11693
rect 2276 11667 2283 11673
rect 2256 11627 2263 11643
rect 2116 11176 2123 11193
rect 2156 11187 2163 11233
rect 1936 10956 1963 10963
rect 1836 10936 1863 10943
rect 1816 10916 1843 10923
rect 1836 10907 1843 10916
rect 1816 10687 1823 10733
rect 1856 10716 1863 10936
rect 1596 9836 1623 9843
rect 1596 9787 1603 9836
rect 1636 9827 1643 9833
rect 1596 9756 1603 9773
rect 1636 9756 1643 9813
rect 1616 9727 1623 9743
rect 1496 8996 1523 9003
rect 1396 8927 1403 8983
rect 1436 8887 1443 8983
rect 1196 8347 1203 8513
rect 1216 8467 1223 8503
rect 1216 8407 1223 8453
rect 1256 8447 1263 8503
rect 1296 8487 1303 8503
rect 1176 8316 1203 8323
rect 1236 8316 1243 8333
rect 1216 8267 1223 8303
rect 1176 8036 1183 8053
rect 1156 7967 1163 8023
rect 1216 7667 1223 8253
rect 1256 7867 1263 8273
rect 1276 7827 1283 8333
rect 1356 8267 1363 8533
rect 1376 8316 1383 8783
rect 1356 7887 1363 7953
rect 1296 7836 1303 7873
rect 1356 7836 1363 7873
rect 1116 7656 1143 7663
rect 1096 7343 1103 7393
rect 1076 7336 1103 7343
rect 1136 7123 1143 7656
rect 1156 7367 1163 7523
rect 1136 7116 1163 7123
rect 1056 7007 1063 7033
rect 1056 6896 1063 6993
rect 1076 6983 1083 7063
rect 1136 7047 1143 7083
rect 1136 6987 1143 7033
rect 1076 6976 1103 6983
rect 1096 6876 1103 6976
rect 1016 6863 1023 6873
rect 1016 6856 1043 6863
rect 1156 6767 1163 7116
rect 956 6527 963 6583
rect 1156 6583 1163 6633
rect 1096 6567 1103 6583
rect 1136 6576 1163 6583
rect 1116 6547 1123 6563
rect 896 6416 903 6493
rect 1176 6383 1183 6413
rect 1056 6376 1083 6383
rect 1156 6376 1183 6383
rect 1056 6267 1063 6376
rect 896 5907 903 6213
rect 976 6127 983 6233
rect 936 6116 963 6123
rect 836 5416 863 5423
rect 816 5127 823 5413
rect 836 4936 863 4943
rect 836 4727 843 4936
rect 876 4916 883 5073
rect 896 4987 903 5653
rect 956 5603 963 6116
rect 976 5987 983 6113
rect 1036 5967 1043 6133
rect 1136 6047 1143 6103
rect 1036 5883 1043 5953
rect 1096 5896 1103 5973
rect 1036 5876 1063 5883
rect 1036 5687 1043 5876
rect 936 5596 963 5603
rect 916 5167 923 5453
rect 936 5403 943 5596
rect 1036 5403 1043 5673
rect 1116 5636 1143 5643
rect 1056 5483 1063 5613
rect 1096 5567 1103 5623
rect 1056 5476 1083 5483
rect 936 5396 963 5403
rect 996 5387 1003 5403
rect 1036 5396 1063 5403
rect 1036 5307 1043 5396
rect 1076 5223 1083 5476
rect 1056 5216 1083 5223
rect 916 5007 923 5123
rect 936 4923 943 5053
rect 1056 4967 1063 5216
rect 1076 4976 1093 4983
rect 1116 4967 1123 5613
rect 1136 5607 1143 5636
rect 1136 5507 1143 5593
rect 1196 5487 1203 7433
rect 1236 7336 1243 7453
rect 1296 7356 1303 7513
rect 1336 7507 1343 7563
rect 1376 7363 1383 8053
rect 1396 7927 1403 8073
rect 1416 8067 1423 8593
rect 1436 8507 1443 8813
rect 1496 8587 1503 8996
rect 1516 8543 1523 8973
rect 1536 8847 1543 9253
rect 1556 9107 1563 9293
rect 1576 9127 1583 9593
rect 1656 9587 1663 10233
rect 1796 10087 1803 10413
rect 1676 9907 1683 9953
rect 1816 9947 1823 10673
rect 1696 9927 1703 9943
rect 1736 9916 1763 9923
rect 1616 9303 1623 9473
rect 1636 9447 1643 9463
rect 1596 9296 1623 9303
rect 1596 9027 1603 9296
rect 1556 8956 1583 8963
rect 1556 8927 1563 8956
rect 1536 8796 1543 8833
rect 1576 8796 1583 8933
rect 1596 8807 1603 8983
rect 1596 8776 1623 8783
rect 1516 8536 1543 8543
rect 1456 8487 1463 8523
rect 1536 8503 1543 8536
rect 1556 8527 1563 8773
rect 1516 8496 1543 8503
rect 1456 8447 1463 8473
rect 1556 8343 1563 8513
rect 1576 8387 1583 8573
rect 1616 8567 1623 8776
rect 1636 8587 1643 8633
rect 1656 8607 1663 9533
rect 1716 9456 1723 9473
rect 1676 9007 1683 9433
rect 1696 8747 1703 9333
rect 1716 8763 1723 9293
rect 1736 9187 1743 9733
rect 1756 9167 1763 9916
rect 1796 9807 1803 9853
rect 1796 9776 1803 9793
rect 1776 9727 1783 9743
rect 1836 9547 1843 10473
rect 1856 10227 1863 10413
rect 1856 9907 1863 9973
rect 1856 9447 1863 9793
rect 1876 9687 1883 10673
rect 1896 10456 1903 10693
rect 1916 10687 1923 10703
rect 1936 10323 1943 10956
rect 1956 10936 1983 10943
rect 2016 10936 2023 10973
rect 1956 10887 1963 10936
rect 1996 10747 2003 10913
rect 1956 10687 1963 10733
rect 1916 10316 1943 10323
rect 1916 10236 1923 10316
rect 1936 10256 1943 10293
rect 1956 10247 1963 10313
rect 1976 10203 1983 10513
rect 1976 10196 1993 10203
rect 1896 9927 1903 9963
rect 1936 9956 1943 10053
rect 1916 9907 1923 9943
rect 1936 9847 1943 9913
rect 1896 9567 1903 9793
rect 1936 9756 1943 9833
rect 1956 9776 1963 9793
rect 1976 9756 2003 9763
rect 1996 9647 2003 9756
rect 1896 9476 1903 9493
rect 1936 9476 1963 9483
rect 1856 9296 1883 9303
rect 1876 9227 1883 9296
rect 1956 9107 1963 9476
rect 1976 9287 1983 9573
rect 1996 9447 2003 9493
rect 2016 9327 2023 10493
rect 2036 10216 2043 10553
rect 2056 10267 2063 10453
rect 2096 10436 2103 11113
rect 2136 10923 2143 11053
rect 2196 10947 2203 11593
rect 2296 11547 2303 11643
rect 2316 11387 2323 11653
rect 2216 11327 2223 11383
rect 2236 11327 2243 11363
rect 2136 10916 2163 10923
rect 2236 10903 2243 11273
rect 2256 11127 2263 11193
rect 2276 11023 2283 11313
rect 2336 11227 2343 11793
rect 2376 11267 2383 11813
rect 2556 11767 2563 11893
rect 2396 11676 2423 11683
rect 2396 11607 2403 11676
rect 2396 11416 2403 11453
rect 2436 11447 2443 11663
rect 2476 11656 2503 11663
rect 2496 11507 2503 11656
rect 2596 11647 2603 11883
rect 2756 11847 2763 11863
rect 2616 11676 2623 11753
rect 2776 11707 2783 11843
rect 2796 11747 2803 11863
rect 2696 11676 2703 11693
rect 2676 11627 2683 11663
rect 2447 11416 2463 11423
rect 2396 11267 2403 11353
rect 2316 11167 2323 11183
rect 2356 11167 2363 11183
rect 2416 11127 2423 11373
rect 2436 11187 2443 11213
rect 2316 11107 2323 11113
rect 2276 11016 2303 11023
rect 2136 10436 2143 10453
rect 2116 10367 2123 10423
rect 2156 10363 2163 10423
rect 2176 10407 2183 10903
rect 2216 10896 2243 10903
rect 2276 10716 2283 10753
rect 2296 10707 2303 11016
rect 2316 10903 2323 11093
rect 2456 11007 2463 11416
rect 2476 11227 2483 11413
rect 2496 11203 2503 11493
rect 2516 11247 2523 11453
rect 2576 11407 2583 11433
rect 2476 11196 2503 11203
rect 2476 10947 2483 11196
rect 2556 11196 2563 11233
rect 2576 11187 2583 11213
rect 2636 10987 2643 11433
rect 2656 11327 2663 11593
rect 2696 11407 2703 11633
rect 2676 11307 2683 11353
rect 2676 11216 2683 11273
rect 2696 11196 2703 11393
rect 2716 11307 2723 11673
rect 2756 11383 2763 11473
rect 2836 11396 2843 11413
rect 2756 11376 2783 11383
rect 2736 11363 2743 11373
rect 2736 11356 2823 11363
rect 2796 11247 2803 11333
rect 2356 10916 2363 10933
rect 2316 10896 2343 10903
rect 2376 10887 2383 10903
rect 2396 10847 2403 10923
rect 2476 10887 2483 10933
rect 2456 10736 2463 10873
rect 2596 10807 2603 10873
rect 2396 10716 2423 10723
rect 2276 10423 2283 10593
rect 2356 10467 2363 10633
rect 2396 10607 2403 10716
rect 2496 10703 2503 10773
rect 2596 10716 2603 10793
rect 2636 10743 2643 10973
rect 2616 10736 2643 10743
rect 2656 10723 2663 10933
rect 2716 10927 2723 11133
rect 2736 11067 2743 11183
rect 2776 10923 2783 11013
rect 2756 10916 2783 10923
rect 2636 10716 2663 10723
rect 2436 10687 2443 10703
rect 2476 10696 2503 10703
rect 2516 10683 2523 10713
rect 2496 10676 2523 10683
rect 2356 10436 2363 10453
rect 2276 10416 2303 10423
rect 2136 10356 2163 10363
rect 2136 9967 2143 10356
rect 2156 10256 2163 10333
rect 2296 10167 2303 10393
rect 2336 10347 2343 10423
rect 2036 9487 2043 9753
rect 2076 9743 2083 9933
rect 2116 9887 2123 9923
rect 2076 9736 2103 9743
rect 2036 9463 2043 9473
rect 2036 9456 2063 9463
rect 2016 9276 2023 9293
rect 1996 9227 2003 9263
rect 2036 9256 2043 9273
rect 2136 9147 2143 9813
rect 2176 9756 2203 9763
rect 2196 9647 2203 9756
rect 2216 9723 2223 9993
rect 2256 9976 2263 10113
rect 2296 9976 2303 10053
rect 2276 9883 2283 9963
rect 2256 9876 2283 9883
rect 2256 9747 2263 9876
rect 2316 9823 2323 10313
rect 2336 10216 2343 10273
rect 2296 9816 2323 9823
rect 2296 9767 2303 9816
rect 2276 9736 2303 9743
rect 2216 9716 2243 9723
rect 2236 9463 2243 9673
rect 2276 9507 2283 9693
rect 2296 9607 2303 9736
rect 2276 9476 2283 9493
rect 2236 9456 2263 9463
rect 1736 9027 1743 9053
rect 1776 9016 1783 9073
rect 1756 8867 1763 9003
rect 1796 8827 1803 9093
rect 1836 9016 1843 9033
rect 1756 8767 1763 8783
rect 1796 8776 1803 8813
rect 1716 8756 1743 8763
rect 1596 8507 1603 8553
rect 1536 8336 1563 8343
rect 1416 7567 1423 8033
rect 1456 7847 1463 8313
rect 1536 8187 1543 8336
rect 1616 8343 1623 8553
rect 1636 8523 1643 8573
rect 1636 8516 1663 8523
rect 1616 8336 1643 8343
rect 1596 8316 1603 8333
rect 1636 8316 1643 8336
rect 1576 8287 1583 8303
rect 1656 8103 1663 8373
rect 1636 8096 1663 8103
rect 1496 8036 1503 8053
rect 1496 7836 1503 7873
rect 1536 7836 1543 7853
rect 1576 7836 1583 8013
rect 1516 7807 1523 7823
rect 1556 7667 1563 7823
rect 1556 7567 1563 7653
rect 1576 7556 1603 7563
rect 1536 7523 1543 7553
rect 1596 7527 1603 7556
rect 1536 7516 1563 7523
rect 1356 7356 1383 7363
rect 1476 7376 1503 7383
rect 1336 7167 1343 7313
rect 1356 7103 1363 7356
rect 1376 7336 1403 7343
rect 1396 7207 1403 7336
rect 1356 7096 1383 7103
rect 1296 7067 1303 7083
rect 1336 7076 1343 7093
rect 1356 7047 1363 7063
rect 1216 6587 1223 6853
rect 1236 6103 1243 6873
rect 1316 6847 1323 7033
rect 1296 6836 1313 6843
rect 1256 6827 1263 6833
rect 1356 6583 1363 6973
rect 1296 6363 1303 6583
rect 1336 6576 1363 6583
rect 1376 6387 1383 7096
rect 1296 6356 1323 6363
rect 1216 6096 1243 6103
rect 1216 5936 1223 6096
rect 1316 6083 1323 6356
rect 1376 6227 1383 6373
rect 1396 6367 1403 7153
rect 1476 7123 1483 7376
rect 1636 7307 1643 8096
rect 1456 7116 1483 7123
rect 1456 7067 1463 7116
rect 1476 7007 1483 7083
rect 1496 7027 1503 7063
rect 1456 6807 1463 6843
rect 1456 6567 1463 6793
rect 1476 6596 1483 6613
rect 1316 6076 1343 6083
rect 1516 5987 1523 6123
rect 1396 5907 1403 5973
rect 1516 5927 1523 5973
rect 1376 5656 1383 5673
rect 1276 5567 1283 5643
rect 1316 5636 1323 5653
rect 1296 5587 1303 5623
rect 1336 5527 1343 5623
rect 1376 5527 1383 5553
rect 1196 5456 1223 5463
rect 1196 5183 1203 5456
rect 1216 5287 1223 5413
rect 1196 5176 1223 5183
rect 1176 5156 1203 5163
rect 1196 4967 1203 5156
rect 1216 5147 1223 5176
rect 1236 5027 1243 5293
rect 1376 5207 1383 5513
rect 1396 5416 1403 5633
rect 1416 5287 1423 5643
rect 1436 5227 1443 5733
rect 1516 5647 1523 5913
rect 1536 5827 1543 6413
rect 1556 5747 1563 7233
rect 1656 7227 1663 8073
rect 1676 7547 1683 8413
rect 1696 8307 1703 8473
rect 1716 8367 1723 8503
rect 1736 8427 1743 8756
rect 1756 8347 1763 8513
rect 1816 8487 1823 8853
rect 1836 8516 1843 8533
rect 1856 8527 1863 9073
rect 1876 8687 1883 9003
rect 1856 8467 1863 8483
rect 1736 8287 1743 8313
rect 1756 8307 1763 8333
rect 1776 8316 1783 8353
rect 1836 8296 1863 8303
rect 1696 8056 1703 8133
rect 1736 8056 1743 8093
rect 1716 7903 1723 8043
rect 1756 7907 1763 8153
rect 1796 8067 1803 8293
rect 1716 7896 1743 7903
rect 1696 7887 1703 7893
rect 1696 7856 1703 7873
rect 1736 7787 1743 7896
rect 1776 7647 1783 7993
rect 1816 7987 1823 8273
rect 1836 8007 1843 8133
rect 1796 7583 1803 7873
rect 1816 7827 1823 7933
rect 1796 7576 1823 7583
rect 1776 7556 1783 7573
rect 1676 7427 1683 7493
rect 1676 7336 1683 7413
rect 1716 7067 1723 7093
rect 1656 7047 1663 7053
rect 1576 6876 1583 7033
rect 1676 6967 1683 7043
rect 1656 6876 1663 6893
rect 1596 6747 1603 6863
rect 1576 6243 1583 6413
rect 1596 6267 1603 6733
rect 1696 6596 1703 6613
rect 1616 6487 1623 6593
rect 1676 6507 1683 6563
rect 1576 6236 1603 6243
rect 1596 6116 1603 6236
rect 1636 5947 1643 6253
rect 1676 6147 1683 6493
rect 1636 5916 1643 5933
rect 1476 5367 1483 5423
rect 1296 5007 1303 5193
rect 1336 5156 1343 5193
rect 1316 5127 1323 5143
rect 916 4916 943 4923
rect 776 4463 783 4693
rect 836 4647 843 4683
rect 816 4496 823 4613
rect 776 4456 803 4463
rect 796 4447 803 4456
rect 856 4427 863 4703
rect 896 4696 903 4713
rect 876 4467 883 4683
rect 956 4483 963 4553
rect 936 4476 963 4483
rect 456 3487 463 3503
rect 436 3236 463 3243
rect 436 3047 443 3236
rect 496 3107 503 3733
rect 516 3487 523 3723
rect 556 3716 563 3913
rect 576 3587 583 3703
rect 656 3647 663 4073
rect 856 3976 863 3993
rect 716 3736 723 3773
rect 616 3516 623 3533
rect 656 3516 663 3613
rect 736 3547 743 3723
rect 756 3567 763 3743
rect 876 3707 883 3833
rect 896 3727 903 4453
rect 916 4007 923 4203
rect 936 4147 943 4476
rect 996 4247 1003 4873
rect 1016 4627 1023 4953
rect 1116 4907 1123 4933
rect 1136 4907 1143 4953
rect 1076 4696 1083 4733
rect 1236 4707 1243 4973
rect 1256 4956 1263 4993
rect 1296 4976 1303 4993
rect 1356 4947 1363 4973
rect 1316 4927 1323 4943
rect 1056 4583 1063 4683
rect 1236 4676 1243 4693
rect 1276 4667 1283 4683
rect 1056 4576 1083 4583
rect 1016 4507 1023 4533
rect 1016 4476 1023 4493
rect 956 3787 963 4233
rect 996 4196 1003 4213
rect 976 3827 983 4193
rect 996 3947 1003 4133
rect 636 3487 643 3503
rect 816 3496 823 3533
rect 876 3523 883 3653
rect 876 3516 903 3523
rect 856 3427 863 3503
rect 896 3447 903 3516
rect 787 3376 793 3383
rect 576 3243 583 3373
rect 556 3236 583 3243
rect 556 3036 563 3173
rect 896 3147 903 3433
rect 916 3207 923 3513
rect 936 3236 943 3513
rect 896 3047 903 3133
rect 456 3007 463 3033
rect 496 2887 503 3013
rect 516 2747 523 2873
rect 596 2787 603 3003
rect 956 2803 963 3633
rect 976 3527 983 3723
rect 996 3127 1003 3933
rect 1016 3807 1023 3873
rect 1016 3736 1023 3793
rect 1036 3727 1043 3993
rect 1056 3767 1063 4413
rect 1076 4267 1083 4576
rect 1116 4507 1123 4573
rect 1216 4523 1223 4663
rect 1256 4587 1263 4663
rect 1316 4567 1323 4913
rect 1196 4516 1223 4523
rect 1096 4456 1123 4463
rect 1116 4327 1123 4456
rect 1076 4187 1083 4253
rect 1196 4247 1203 4516
rect 1376 4267 1383 5113
rect 1396 4547 1403 5213
rect 1476 5187 1483 5353
rect 1536 5207 1543 5603
rect 1616 5416 1623 5493
rect 1656 5416 1663 5433
rect 1696 5407 1703 6333
rect 1556 5176 1583 5183
rect 1436 4967 1443 5133
rect 1576 5127 1583 5176
rect 1596 5127 1603 5393
rect 1676 5347 1683 5403
rect 1476 4956 1503 4963
rect 1496 4927 1503 4956
rect 1436 4727 1443 4893
rect 1436 4676 1443 4713
rect 1536 4703 1543 5013
rect 1556 4747 1563 5093
rect 1576 5027 1583 5113
rect 1616 4956 1623 4993
rect 1656 4956 1663 5193
rect 1716 5156 1723 5213
rect 1736 5187 1743 7533
rect 1796 7527 1803 7543
rect 1776 7343 1783 7373
rect 1796 7347 1803 7513
rect 1756 7336 1783 7343
rect 1756 6427 1763 7093
rect 1796 6967 1803 7333
rect 1816 7227 1823 7576
rect 1836 7247 1843 7953
rect 1856 7887 1863 8296
rect 1896 8287 1903 8773
rect 1936 8767 1943 8873
rect 1996 8796 2003 8963
rect 2156 8843 2163 9393
rect 2176 9287 2183 9413
rect 2256 9307 2263 9456
rect 2256 9276 2283 9283
rect 2136 8836 2163 8843
rect 2036 8796 2043 8813
rect 1916 8287 1923 8513
rect 1936 8327 1943 8493
rect 1956 8483 1963 8733
rect 1976 8547 1983 8783
rect 1956 8476 1983 8483
rect 1916 8067 1923 8273
rect 1936 8127 1943 8313
rect 1876 8027 1883 8043
rect 1916 8036 1923 8053
rect 1896 7867 1903 8023
rect 1956 7867 1963 8053
rect 1976 7827 1983 8476
rect 1996 8316 2003 8473
rect 2016 8467 2023 8503
rect 2016 8267 2023 8283
rect 2016 8127 2023 8253
rect 1996 8027 2003 8113
rect 1856 7347 1863 7813
rect 1876 7247 1883 7793
rect 1896 7187 1903 7823
rect 1996 7567 2003 7913
rect 2016 7507 2023 8093
rect 2036 7967 2043 8493
rect 2056 8316 2083 8323
rect 2056 8023 2063 8233
rect 2076 8147 2083 8316
rect 2096 8036 2103 8113
rect 2116 8047 2123 8113
rect 2136 8063 2143 8836
rect 2196 8783 2203 9093
rect 2176 8776 2203 8783
rect 2176 8523 2183 8776
rect 2156 8516 2183 8523
rect 2156 8083 2163 8516
rect 2216 8507 2223 9233
rect 2236 8507 2243 9113
rect 2276 8927 2283 9276
rect 2176 8367 2183 8473
rect 2236 8323 2243 8373
rect 2216 8316 2243 8323
rect 2236 8287 2243 8316
rect 2156 8076 2183 8083
rect 2136 8056 2163 8063
rect 2056 8016 2083 8023
rect 1936 7387 1943 7453
rect 1896 7063 1903 7153
rect 1916 7067 1923 7343
rect 1876 7056 1903 7063
rect 1816 6876 1823 6933
rect 1916 6927 1923 7053
rect 1856 6876 1883 6883
rect 1876 6847 1883 6876
rect 1776 6327 1783 6383
rect 1796 6187 1803 6613
rect 1836 6596 1843 6613
rect 1816 6487 1823 6583
rect 1816 6327 1823 6473
rect 1856 6376 1883 6383
rect 1816 6287 1823 6313
rect 1836 6187 1843 6353
rect 1856 6247 1863 6376
rect 1756 6136 1763 6173
rect 1776 5883 1783 6123
rect 1816 6107 1823 6173
rect 1816 5896 1823 5973
rect 1776 5876 1803 5883
rect 1756 5167 1763 5633
rect 1836 5627 1843 5873
rect 1796 5147 1803 5453
rect 1816 5367 1823 5403
rect 1856 5387 1863 5403
rect 1876 5387 1883 5883
rect 1896 5607 1903 6913
rect 1916 6807 1923 6873
rect 1936 6567 1943 7293
rect 1956 6987 1963 7493
rect 1996 7336 2023 7343
rect 1996 7207 2003 7336
rect 2036 7147 2043 7853
rect 2056 7727 2063 7953
rect 2076 7816 2083 7913
rect 2096 7836 2103 7993
rect 2116 7927 2123 8003
rect 2116 7807 2123 7823
rect 2136 7556 2143 7773
rect 2156 7627 2163 8056
rect 2176 7707 2183 8076
rect 2256 8007 2263 8833
rect 2296 8783 2303 8993
rect 2316 8947 2323 9493
rect 2336 8887 2343 9313
rect 2356 8827 2363 9633
rect 2376 9507 2383 10053
rect 2396 9776 2403 10353
rect 2436 10223 2443 10393
rect 2476 10387 2483 10433
rect 2416 10216 2443 10223
rect 2476 10007 2483 10193
rect 2496 9947 2503 10676
rect 2636 10256 2643 10413
rect 2656 10327 2663 10716
rect 2696 10707 2703 10903
rect 2736 10827 2743 10903
rect 2796 10787 2803 11233
rect 2876 11227 2883 11753
rect 2916 11547 2923 11893
rect 2956 11847 2963 11883
rect 3136 11876 3163 11883
rect 3156 11867 3163 11876
rect 3116 11807 3123 11863
rect 2916 11347 2923 11533
rect 2936 11407 2943 11653
rect 2956 11427 2963 11653
rect 2996 11643 3003 11733
rect 3076 11656 3083 11713
rect 2996 11636 3023 11643
rect 3016 11487 3023 11636
rect 3036 11423 3043 11533
rect 3016 11416 3043 11423
rect 3016 11396 3023 11416
rect 3056 11407 3063 11473
rect 3156 11447 3163 11853
rect 3256 11747 3263 11863
rect 3196 11643 3203 11713
rect 3196 11636 3223 11643
rect 3256 11587 3263 11633
rect 3276 11563 3283 11843
rect 3456 11767 3463 11863
rect 3376 11676 3403 11683
rect 3316 11667 3323 11673
rect 3256 11556 3283 11563
rect 3136 11416 3183 11423
rect 2856 11196 2883 11203
rect 2836 10943 2843 11193
rect 2856 10963 2863 11196
rect 2936 11176 2943 11393
rect 3056 11383 3063 11393
rect 3036 11376 3063 11383
rect 2856 10956 2883 10963
rect 2836 10936 2863 10943
rect 2856 10727 2863 10936
rect 2876 10907 2883 10956
rect 2916 10927 2923 10933
rect 2876 10787 2883 10893
rect 2896 10887 2903 10903
rect 2956 10867 2963 10923
rect 2976 10907 2983 10973
rect 2776 10696 2803 10703
rect 2756 10423 2763 10693
rect 2776 10467 2783 10696
rect 2836 10667 2843 10703
rect 2876 10683 2883 10733
rect 2896 10687 2903 10713
rect 2976 10696 2983 10713
rect 2856 10676 2883 10683
rect 2676 10387 2683 10423
rect 2736 10416 2763 10423
rect 2856 10423 2863 10676
rect 2996 10676 3003 11293
rect 3016 10707 3023 11053
rect 2936 10436 2943 10453
rect 2856 10416 2883 10423
rect 2516 10216 2543 10223
rect 2536 10087 2543 10216
rect 2796 10083 2803 10273
rect 2816 10216 2823 10273
rect 2916 10223 2923 10253
rect 2956 10227 2963 10423
rect 2896 10216 2923 10223
rect 2796 10076 2823 10083
rect 2576 9956 2583 10053
rect 2636 9967 2643 10073
rect 2676 9976 2683 9993
rect 2536 9943 2543 9953
rect 2616 9947 2623 9963
rect 2536 9936 2563 9943
rect 2596 9907 2603 9943
rect 2396 9483 2403 9733
rect 2396 9476 2423 9483
rect 2456 9476 2463 9493
rect 2436 9387 2443 9463
rect 2376 8996 2383 9353
rect 2456 9287 2463 9433
rect 2476 9347 2483 9463
rect 2536 9347 2543 9473
rect 2476 9296 2503 9303
rect 2496 9227 2503 9296
rect 2496 9087 2503 9213
rect 2476 8947 2483 8993
rect 2536 8987 2543 9333
rect 2556 8983 2563 9773
rect 2636 9743 2643 9873
rect 2696 9743 2703 9913
rect 2776 9747 2783 9873
rect 2636 9736 2663 9743
rect 2696 9736 2723 9743
rect 2656 9467 2663 9736
rect 2716 9367 2723 9736
rect 2816 9743 2823 10076
rect 2996 9927 3003 10613
rect 3056 10307 3063 11213
rect 3116 11196 3123 11353
rect 3136 11307 3143 11416
rect 3176 11396 3183 11416
rect 3156 11347 3163 11373
rect 3136 11287 3143 11293
rect 3156 11196 3163 11233
rect 3076 11176 3103 11183
rect 3076 11147 3083 11176
rect 3136 11127 3143 11183
rect 3196 11167 3203 11383
rect 3076 10667 3083 11053
rect 3096 10887 3103 10903
rect 3116 10456 3123 10873
rect 3136 10627 3143 10733
rect 3096 10227 3103 10433
rect 3016 9947 3023 9963
rect 2976 9776 2983 9893
rect 3016 9887 3023 9933
rect 2796 9736 2823 9743
rect 2776 9483 2783 9733
rect 2776 9476 2803 9483
rect 2916 9476 2923 9533
rect 2776 9296 2783 9373
rect 2796 9287 2803 9476
rect 2596 9256 2603 9273
rect 2896 9256 2923 9263
rect 2556 8976 2583 8983
rect 2296 8776 2323 8783
rect 2296 8283 2303 8333
rect 2316 8307 2323 8776
rect 2376 8516 2383 8533
rect 2416 8527 2423 8933
rect 2496 8776 2503 8973
rect 2556 8796 2583 8803
rect 2336 8283 2343 8473
rect 2356 8447 2363 8503
rect 2396 8387 2403 8483
rect 2416 8316 2443 8323
rect 2296 8276 2323 8283
rect 2336 8276 2363 8283
rect 2216 7607 2223 7913
rect 2216 7547 2223 7593
rect 2116 7527 2123 7543
rect 2156 7523 2163 7543
rect 2136 7516 2163 7523
rect 2136 7376 2143 7516
rect 2196 7507 2203 7543
rect 2236 7447 2243 7993
rect 2276 7887 2283 8043
rect 2316 8036 2323 8276
rect 2356 8247 2363 8276
rect 2356 8023 2363 8233
rect 2396 8147 2403 8303
rect 2436 8267 2443 8316
rect 2456 8227 2463 8773
rect 2576 8747 2583 8796
rect 2336 8016 2363 8023
rect 2316 7803 2323 7873
rect 2336 7836 2343 7853
rect 2296 7796 2323 7803
rect 2296 7627 2303 7796
rect 2396 7787 2403 8133
rect 2416 8047 2423 8173
rect 2456 8107 2463 8173
rect 2496 8167 2503 8513
rect 2596 8503 2603 8933
rect 2616 8787 2623 8983
rect 2576 8496 2603 8503
rect 2516 8207 2523 8493
rect 2596 8447 2603 8496
rect 2616 8387 2623 8773
rect 2596 8316 2603 8333
rect 2576 8287 2583 8303
rect 2516 8056 2523 8093
rect 2416 7827 2423 8033
rect 2516 7836 2523 7973
rect 2556 7867 2563 8213
rect 2416 7723 2423 7813
rect 2496 7807 2503 7823
rect 2416 7716 2443 7723
rect 2336 7547 2343 7563
rect 2376 7556 2383 7573
rect 2296 7427 2303 7493
rect 2296 7343 2303 7413
rect 2296 7336 2323 7343
rect 2076 7076 2083 7153
rect 2116 7063 2123 7113
rect 2056 7007 2063 7063
rect 2096 7056 2123 7063
rect 1956 6463 1963 6913
rect 1996 6856 2003 6873
rect 2036 6847 2043 6933
rect 1996 6607 2003 6793
rect 2036 6607 2043 6613
rect 2096 6603 2103 6773
rect 2076 6596 2103 6603
rect 2016 6547 2023 6583
rect 2056 6507 2063 6583
rect 2136 6467 2143 7333
rect 2236 7096 2243 7133
rect 2256 7047 2263 7083
rect 2196 6856 2203 6893
rect 2236 6867 2243 6913
rect 2176 6827 2183 6843
rect 2276 6747 2283 6873
rect 2196 6587 2203 6633
rect 2236 6596 2243 6633
rect 2296 6627 2303 7336
rect 2216 6567 2223 6583
rect 1956 6456 1983 6463
rect 1976 6267 1983 6456
rect 1996 6416 2003 6433
rect 2156 6343 2163 6533
rect 2156 6336 2183 6343
rect 2176 6327 2183 6336
rect 1916 5896 1923 6233
rect 1996 5987 2003 6113
rect 1936 5607 1943 5623
rect 2016 5507 2023 6253
rect 2176 6116 2183 6313
rect 2216 6227 2223 6553
rect 2276 6547 2283 6603
rect 2116 6087 2123 6103
rect 2156 6027 2163 6103
rect 2036 5936 2043 6013
rect 2196 5887 2203 6103
rect 2216 5927 2223 5993
rect 2216 5896 2223 5913
rect 2236 5787 2243 6453
rect 2276 6383 2283 6413
rect 2296 6387 2303 6613
rect 2256 6376 2283 6383
rect 2276 5667 2283 6133
rect 2296 6127 2303 6273
rect 2316 5903 2323 6473
rect 2336 6347 2343 7473
rect 2396 7383 2403 7533
rect 2376 7376 2403 7383
rect 2356 6876 2363 7033
rect 2376 6987 2383 7376
rect 2436 7167 2443 7716
rect 2456 7547 2463 7793
rect 2536 7787 2543 7823
rect 2496 7627 2503 7673
rect 2556 7627 2563 7653
rect 2476 7167 2483 7573
rect 2496 7523 2503 7613
rect 2576 7527 2583 8273
rect 2596 8067 2603 8213
rect 2596 7567 2603 8053
rect 2496 7516 2523 7523
rect 2416 7096 2423 7133
rect 2456 7096 2483 7103
rect 2396 6876 2403 6893
rect 2436 6876 2443 7083
rect 2376 6807 2383 6863
rect 2416 6787 2423 6863
rect 2476 6847 2483 7096
rect 2396 6687 2403 6753
rect 2376 6587 2383 6653
rect 2396 6583 2403 6673
rect 2436 6596 2443 6633
rect 2476 6587 2483 6603
rect 2396 6576 2423 6583
rect 2436 6396 2443 6433
rect 2396 6376 2423 6383
rect 2396 6287 2403 6376
rect 2456 6267 2463 6383
rect 2336 6147 2343 6253
rect 2396 6127 2403 6253
rect 2496 6223 2503 7433
rect 2516 7347 2523 7516
rect 2576 7407 2583 7433
rect 2576 7376 2583 7393
rect 2536 7343 2543 7373
rect 2536 7336 2563 7343
rect 2536 7127 2543 7336
rect 2616 7327 2623 8153
rect 2636 8056 2643 9133
rect 2916 9127 2923 9256
rect 2956 9087 2963 9093
rect 2976 9087 2983 9293
rect 2996 9127 3003 9233
rect 2776 8996 2783 9073
rect 2956 9016 2963 9073
rect 2656 8427 2663 8953
rect 2716 8796 2733 8803
rect 2716 8776 2723 8796
rect 2696 8507 2703 8613
rect 2656 8267 2663 8313
rect 2656 8127 2663 8153
rect 2676 8087 2683 8453
rect 2696 8087 2703 8293
rect 2716 8047 2723 8733
rect 2736 8347 2743 8503
rect 2756 8443 2763 8483
rect 2756 8436 2783 8443
rect 2736 8227 2743 8333
rect 2736 8047 2743 8113
rect 2656 7867 2663 8013
rect 2696 7856 2703 7873
rect 2636 7747 2643 7853
rect 2656 7807 2663 7853
rect 2716 7807 2723 7823
rect 2636 7707 2643 7713
rect 2516 6487 2523 6833
rect 2536 6587 2543 7113
rect 2476 6216 2503 6223
rect 2416 6136 2423 6173
rect 2436 6103 2443 6133
rect 2416 6096 2443 6103
rect 2296 5896 2323 5903
rect 2356 5707 2363 5933
rect 2396 5867 2403 5913
rect 2396 5747 2403 5853
rect 2416 5847 2423 6096
rect 2476 5947 2483 6216
rect 2556 6063 2563 7313
rect 2576 7063 2583 7153
rect 2596 7107 2603 7273
rect 2616 7076 2623 7133
rect 2576 7056 2603 7063
rect 2596 6907 2603 7056
rect 2636 7027 2643 7693
rect 2656 7087 2663 7553
rect 2676 7307 2683 7543
rect 2756 7487 2763 8353
rect 2776 8316 2783 8436
rect 2796 8367 2803 8983
rect 2976 8927 2983 9003
rect 3016 8967 3023 9433
rect 3036 9256 3043 9593
rect 3076 9547 3083 10213
rect 3116 9483 3123 10393
rect 3156 10247 3163 10913
rect 3176 10907 3183 11093
rect 3196 10927 3203 11113
rect 3216 10867 3223 11373
rect 3196 10716 3203 10793
rect 3236 10767 3243 11333
rect 3256 10907 3263 11556
rect 3316 11407 3323 11653
rect 3376 11507 3383 11676
rect 3436 11627 3443 11633
rect 3436 11503 3443 11613
rect 3456 11527 3463 11693
rect 3476 11627 3483 11843
rect 3496 11787 3503 11863
rect 3616 11827 3623 11896
rect 3947 11896 3963 11903
rect 3996 11896 4023 11903
rect 3436 11496 3463 11503
rect 3316 11323 3323 11393
rect 3336 11343 3343 11413
rect 3376 11396 3403 11403
rect 3396 11367 3403 11396
rect 3336 11336 3363 11343
rect 3316 11316 3343 11323
rect 3316 11176 3323 11193
rect 3276 10767 3283 11133
rect 3296 10747 3303 11163
rect 3336 11156 3343 11316
rect 3356 11207 3363 11336
rect 3356 11176 3363 11193
rect 3376 10967 3383 11353
rect 3396 11307 3403 11353
rect 3436 11267 3443 11293
rect 3436 11207 3443 11213
rect 3456 11203 3463 11496
rect 3496 11387 3503 11773
rect 3576 11656 3583 11753
rect 3536 11487 3543 11533
rect 3536 11396 3543 11473
rect 3556 11467 3563 11643
rect 3596 11587 3603 11643
rect 3556 11427 3563 11453
rect 3596 11403 3603 11533
rect 3576 11396 3603 11403
rect 3516 11367 3523 11383
rect 3487 11216 3503 11223
rect 3456 11196 3483 11203
rect 3396 11147 3403 11193
rect 3436 10967 3443 11193
rect 3316 10936 3323 10953
rect 3356 10936 3363 10953
rect 3236 10716 3243 10733
rect 3256 10647 3263 10703
rect 3296 10687 3303 10713
rect 3316 10663 3323 10893
rect 3336 10847 3343 10913
rect 3376 10887 3383 10953
rect 3456 10847 3463 11196
rect 3556 11067 3563 11383
rect 3576 10903 3583 11153
rect 3616 11107 3623 11553
rect 3636 11267 3643 11653
rect 3656 11487 3663 11883
rect 3636 11207 3643 11253
rect 3696 11207 3703 11893
rect 3796 11867 3803 11883
rect 3756 11676 3763 11753
rect 3796 11676 3823 11683
rect 3816 11567 3823 11676
rect 3876 11647 3883 11893
rect 3976 11687 3983 11883
rect 3916 11547 3923 11653
rect 3996 11643 4003 11773
rect 4016 11687 4023 11896
rect 4176 11896 4203 11903
rect 4196 11847 4203 11896
rect 4136 11696 4143 11773
rect 4296 11707 4303 11713
rect 4156 11676 4183 11683
rect 3936 11547 3943 11643
rect 3976 11636 4003 11643
rect 3736 11247 3743 11273
rect 3636 10987 3643 11193
rect 3716 11156 3723 11213
rect 3736 11176 3743 11233
rect 3296 10656 3323 10663
rect 3176 10007 3183 10473
rect 3296 10456 3303 10656
rect 3276 10423 3283 10443
rect 3276 10416 3303 10423
rect 3216 10236 3243 10243
rect 3256 10236 3263 10293
rect 3236 10207 3243 10236
rect 3236 10067 3243 10193
rect 3136 9976 3163 9983
rect 3136 9863 3143 9976
rect 3136 9856 3163 9863
rect 3156 9723 3163 9856
rect 3136 9716 3163 9723
rect 3176 9723 3183 9993
rect 3196 9763 3203 9963
rect 3216 9787 3223 9953
rect 3296 9867 3303 10416
rect 3316 10027 3323 10233
rect 3376 10187 3383 10733
rect 3436 10716 3443 10733
rect 3416 10687 3423 10703
rect 3456 10696 3463 10713
rect 3476 10467 3483 10713
rect 3396 10236 3403 10313
rect 3456 10267 3463 10443
rect 3496 10436 3503 10903
rect 3556 10896 3583 10903
rect 3476 10343 3483 10423
rect 3476 10336 3503 10343
rect 3456 10207 3463 10223
rect 3496 10203 3503 10336
rect 3536 10307 3543 10733
rect 3476 10196 3503 10203
rect 3456 9867 3463 10013
rect 3476 9927 3483 10196
rect 3556 10047 3563 10353
rect 3496 9947 3503 9963
rect 3536 9887 3543 9933
rect 3196 9756 3223 9763
rect 3216 9747 3223 9756
rect 3176 9716 3203 9723
rect 3136 9587 3143 9716
rect 3216 9607 3223 9733
rect 3116 9476 3143 9483
rect 2856 8807 2863 8813
rect 2836 8767 2843 8793
rect 2816 8343 2823 8553
rect 2856 8507 2863 8633
rect 2796 8336 2823 8343
rect 2776 7787 2783 8213
rect 2796 8067 2803 8293
rect 2836 8083 2843 8373
rect 2856 8227 2863 8493
rect 2876 8227 2883 8813
rect 2916 8567 2923 8753
rect 2996 8627 3003 8793
rect 3056 8667 3063 9453
rect 3076 9427 3083 9463
rect 3236 9387 3243 9473
rect 3256 9367 3263 9773
rect 3336 9743 3343 9853
rect 3356 9776 3363 9853
rect 3336 9736 3363 9743
rect 3536 9736 3543 9873
rect 3316 9476 3323 9493
rect 3356 9487 3363 9736
rect 3376 9527 3383 9573
rect 3096 8987 3103 9013
rect 3076 8796 3083 8813
rect 3116 8796 3123 9113
rect 3136 8996 3143 9353
rect 3296 9347 3303 9463
rect 3156 9296 3163 9333
rect 3176 8996 3183 9113
rect 2996 8527 3003 8613
rect 2976 8487 2983 8523
rect 2936 8183 2943 8433
rect 2996 8316 3003 8433
rect 2936 8176 2963 8183
rect 2816 8076 2843 8083
rect 2756 7356 2763 7393
rect 2776 7347 2783 7373
rect 2696 7327 2703 7343
rect 2796 7167 2803 8033
rect 2816 7827 2823 8076
rect 2856 7967 2863 8043
rect 2816 7347 2823 7813
rect 2816 7327 2823 7333
rect 2616 6876 2623 6913
rect 2636 6856 2643 6913
rect 2576 6587 2583 6713
rect 2596 6607 2603 6853
rect 2656 6647 2663 7073
rect 2696 6603 2703 6853
rect 2676 6596 2703 6603
rect 2656 6567 2663 6583
rect 2596 6427 2603 6433
rect 2676 6367 2683 6573
rect 2716 6527 2723 7153
rect 2736 7023 2743 7053
rect 2776 7047 2783 7063
rect 2796 7047 2803 7083
rect 2836 7067 2843 7893
rect 2856 7667 2863 7873
rect 2876 7867 2883 8063
rect 2896 7856 2903 7993
rect 2916 7887 2923 8073
rect 2916 7787 2923 7823
rect 2956 7787 2963 8176
rect 2736 7016 2763 7023
rect 2736 6087 2743 6413
rect 2756 6163 2763 7016
rect 2796 6487 2803 6753
rect 2836 6616 2843 6633
rect 2876 6623 2883 7773
rect 2936 7387 2943 7773
rect 2976 7743 2983 8193
rect 2996 8023 3003 8213
rect 3016 8047 3023 8473
rect 3036 8327 3043 8513
rect 3096 8483 3103 8733
rect 3156 8587 3163 8953
rect 3196 8787 3203 8793
rect 3236 8787 3243 9173
rect 3316 8827 3323 9333
rect 3336 9256 3343 9273
rect 3376 9247 3383 9513
rect 3516 9476 3523 9493
rect 3376 8983 3383 9173
rect 3356 8947 3363 8983
rect 3376 8976 3403 8983
rect 3416 8947 3423 9263
rect 3316 8796 3343 8803
rect 3116 8507 3123 8523
rect 3136 8483 3143 8503
rect 3096 8476 3143 8483
rect 3176 8447 3183 8503
rect 3196 8487 3203 8773
rect 3336 8687 3343 8796
rect 3336 8503 3343 8673
rect 3136 8147 3143 8283
rect 3176 8276 3183 8373
rect 3196 8296 3203 8473
rect 3296 8287 3303 8333
rect 3156 8167 3163 8213
rect 3316 8167 3323 8503
rect 3336 8496 3363 8503
rect 3336 8316 3343 8393
rect 3416 8347 3423 8873
rect 3436 8847 3443 9453
rect 3496 9327 3503 9463
rect 3536 9247 3543 9463
rect 3556 9347 3563 10033
rect 3576 9987 3583 10693
rect 3616 10447 3623 10553
rect 3636 10463 3643 10773
rect 3656 10747 3663 11093
rect 3676 10987 3683 11113
rect 3676 10936 3683 10973
rect 3716 10936 3743 10943
rect 3696 10887 3703 10923
rect 3736 10847 3743 10936
rect 3656 10716 3663 10733
rect 3636 10456 3663 10463
rect 3656 10436 3663 10456
rect 3676 10407 3683 10423
rect 3696 10307 3703 10443
rect 3636 10236 3643 10253
rect 3676 10236 3683 10253
rect 3596 10216 3623 10223
rect 3596 9963 3603 10216
rect 3576 9956 3603 9963
rect 3596 9943 3603 9956
rect 3596 9936 3623 9943
rect 3576 9496 3583 9513
rect 3596 9447 3603 9913
rect 3616 9867 3623 9936
rect 3616 9727 3623 9743
rect 3616 9527 3623 9693
rect 3636 9487 3643 10173
rect 3656 9967 3663 10073
rect 3676 9587 3683 9973
rect 3696 9627 3703 10233
rect 3716 9807 3723 10833
rect 3736 9983 3743 10753
rect 3756 10527 3763 11213
rect 3776 10907 3783 11473
rect 3836 11163 3843 11413
rect 3876 11347 3883 11393
rect 3916 11347 3923 11363
rect 3936 11347 3943 11383
rect 3956 11367 3963 11533
rect 3936 11327 3943 11333
rect 3836 11156 3863 11163
rect 3896 11147 3903 11163
rect 3896 11127 3903 11133
rect 3916 11087 3923 11193
rect 3756 10456 3763 10473
rect 3776 10327 3783 10893
rect 3836 10867 3843 10933
rect 3796 10716 3803 10793
rect 3836 10736 3843 10853
rect 3876 10847 3883 10853
rect 3876 10703 3883 10833
rect 3816 10647 3823 10703
rect 3856 10696 3883 10703
rect 3916 10667 3923 11073
rect 3996 10903 4003 11493
rect 4076 11287 4083 11673
rect 4176 11567 4183 11676
rect 4356 11667 4363 11863
rect 4256 11656 4283 11663
rect 4256 11607 4263 11656
rect 4096 11396 4103 11453
rect 4076 11176 4083 11213
rect 4116 11163 4123 11433
rect 4136 11287 4143 11383
rect 4176 11367 4183 11553
rect 4256 11507 4263 11593
rect 4276 11423 4283 11533
rect 4296 11527 4303 11653
rect 4316 11587 4323 11663
rect 4356 11647 4363 11653
rect 4376 11647 4383 11673
rect 4316 11427 4323 11573
rect 4356 11487 4363 11493
rect 4256 11416 4283 11423
rect 4236 11387 4243 11413
rect 4156 11287 4163 11363
rect 4136 11203 4143 11273
rect 4156 11227 4163 11273
rect 4136 11196 4163 11203
rect 4056 11027 4063 11163
rect 4096 11156 4123 11163
rect 4076 10903 4083 11073
rect 4136 10927 4143 11173
rect 3996 10896 4023 10903
rect 4056 10896 4083 10903
rect 4036 10867 4043 10883
rect 4116 10787 4123 10913
rect 4156 10887 4163 11196
rect 4176 11187 4183 11293
rect 4196 11196 4223 11203
rect 4256 11196 4263 11416
rect 4296 11307 4303 11363
rect 4316 11267 4323 11383
rect 4196 11047 4203 11196
rect 4336 11187 4343 11453
rect 4356 11207 4363 11473
rect 4396 11207 4403 11853
rect 4516 11807 4523 11843
rect 4576 11807 4583 11873
rect 4496 11696 4503 11773
rect 4236 10867 4243 10903
rect 3996 10736 4003 10753
rect 4116 10707 4123 10773
rect 4256 10727 4263 10923
rect 3976 10667 3983 10703
rect 4176 10683 4183 10713
rect 4176 10676 4203 10683
rect 3816 10427 3823 10633
rect 3936 10247 3943 10253
rect 3976 10236 3983 10293
rect 4096 10287 4103 10443
rect 4156 10436 4183 10443
rect 4156 10307 4163 10436
rect 4156 10267 4163 10293
rect 3736 9976 3763 9983
rect 3716 9647 3723 9773
rect 3756 9763 3763 9976
rect 3796 9947 3803 10213
rect 3816 9976 3843 9983
rect 3776 9827 3783 9943
rect 3776 9767 3783 9793
rect 3736 9756 3763 9763
rect 3736 9487 3743 9756
rect 3816 9756 3823 9773
rect 3756 9627 3763 9733
rect 3836 9707 3843 9976
rect 3876 9927 3883 10233
rect 3996 10216 4003 10253
rect 4176 10236 4183 10253
rect 4156 10007 4163 10213
rect 4156 9887 4163 9963
rect 3916 9747 3923 9773
rect 3856 9707 3863 9723
rect 3616 9267 3623 9483
rect 3636 9296 3643 9313
rect 3816 9256 3823 9273
rect 3476 9227 3483 9233
rect 3616 9127 3623 9253
rect 3516 9003 3523 9053
rect 3516 8996 3543 9003
rect 3436 8796 3443 8833
rect 3516 8796 3543 8803
rect 3536 8787 3543 8796
rect 3456 8727 3463 8783
rect 3476 8523 3483 8553
rect 3476 8516 3503 8523
rect 3536 8516 3543 8733
rect 3556 8547 3563 8983
rect 3596 8967 3603 8983
rect 3576 8956 3593 8963
rect 3576 8503 3583 8956
rect 3036 8036 3043 8053
rect 3076 8036 3103 8043
rect 2996 8016 3023 8023
rect 2976 7736 3003 7743
rect 2956 7527 2963 7553
rect 2996 7427 3003 7736
rect 3016 7523 3023 8016
rect 3076 8003 3083 8036
rect 3056 7996 3083 8003
rect 3076 7787 3083 7873
rect 3156 7867 3163 8133
rect 3116 7836 3123 7853
rect 3096 7816 3103 7833
rect 3036 7543 3043 7593
rect 3116 7556 3143 7563
rect 3036 7536 3063 7543
rect 3016 7516 3043 7523
rect 2936 7356 2983 7363
rect 2896 6827 2903 7213
rect 2976 7127 2983 7356
rect 2996 7347 3003 7393
rect 2936 7063 2943 7093
rect 2976 7076 2983 7093
rect 3036 7083 3043 7516
rect 3096 7403 3103 7513
rect 3076 7396 3103 7403
rect 3016 7076 3043 7083
rect 2936 7056 2963 7063
rect 3036 7043 3043 7076
rect 2996 7027 3003 7043
rect 3016 7036 3043 7043
rect 2936 6876 2943 7013
rect 2976 6876 2983 6893
rect 2856 6616 2883 6623
rect 2816 6547 2823 6583
rect 2796 6416 2803 6473
rect 2836 6447 2843 6513
rect 2856 6443 2863 6616
rect 2916 6603 2923 6853
rect 2916 6596 2943 6603
rect 2876 6487 2883 6583
rect 2936 6547 2943 6596
rect 2956 6587 2963 6863
rect 2996 6856 3003 6873
rect 2856 6436 2883 6443
rect 2776 6327 2783 6383
rect 2776 6247 2783 6313
rect 2756 6156 2783 6163
rect 2556 6056 2583 6063
rect 2436 5916 2443 5933
rect 2276 5636 2283 5653
rect 1976 5416 2003 5423
rect 1776 5047 1783 5143
rect 1676 4936 1683 4953
rect 1836 4936 1843 5153
rect 1856 5107 1863 5373
rect 1976 5347 1983 5416
rect 2036 5416 2043 5453
rect 2016 5396 2023 5413
rect 2076 5403 2083 5533
rect 2056 5396 2083 5403
rect 1936 5127 1943 5143
rect 1896 4956 1923 4963
rect 1516 4696 1543 4703
rect 1476 4676 1503 4683
rect 1416 4627 1423 4663
rect 1396 4456 1403 4473
rect 1056 3707 1063 3723
rect 1076 3643 1083 4173
rect 1116 4023 1123 4233
rect 1156 4196 1163 4233
rect 1376 4216 1383 4253
rect 1176 4167 1183 4183
rect 1116 4016 1143 4023
rect 1096 3996 1103 4013
rect 1216 3987 1223 4013
rect 1316 3996 1343 4003
rect 1156 3947 1163 3983
rect 1336 3947 1343 3996
rect 1176 3667 1183 3683
rect 1076 3636 1103 3643
rect 1036 3516 1043 3533
rect 1076 3516 1083 3573
rect 1016 3496 1023 3513
rect 1056 3387 1063 3503
rect 1056 3247 1063 3353
rect 936 2796 963 2803
rect 656 2747 663 2763
rect 756 2723 763 2753
rect 576 2707 583 2723
rect 756 2716 783 2723
rect 436 2556 443 2573
rect 636 2567 643 2633
rect 936 2627 943 2796
rect 976 2763 983 3013
rect 1076 2787 1083 3273
rect 1096 3267 1103 3636
rect 1216 3496 1223 3553
rect 1256 3483 1263 3593
rect 1336 3496 1343 3673
rect 1376 3667 1383 4013
rect 1396 3607 1403 4253
rect 1416 3727 1423 4453
rect 1436 3987 1443 4533
rect 1496 4487 1503 4676
rect 1496 4463 1503 4473
rect 1476 4456 1503 4463
rect 1516 4447 1523 4696
rect 1556 4267 1563 4733
rect 1576 4327 1583 4683
rect 1596 4387 1603 4933
rect 1876 4807 1883 4943
rect 1916 4667 1923 4956
rect 1916 4627 1923 4653
rect 1616 4456 1623 4473
rect 1636 4447 1643 4573
rect 1656 4467 1663 4593
rect 1936 4587 1943 5113
rect 1956 5107 1963 5123
rect 1956 5007 1963 5093
rect 1976 4867 1983 4953
rect 1996 4907 2003 5373
rect 2096 5227 2103 5613
rect 2136 5587 2143 5603
rect 2296 5527 2303 5623
rect 2036 5147 2043 5173
rect 2176 5147 2183 5473
rect 2227 5436 2243 5443
rect 2196 5187 2203 5423
rect 2096 5127 2103 5143
rect 2156 5047 2163 5143
rect 2016 4956 2043 4963
rect 2016 4807 2023 4956
rect 2056 4927 2063 4943
rect 1956 4676 1963 4733
rect 2056 4567 2063 4913
rect 2076 4807 2083 4933
rect 2156 4927 2163 5033
rect 2096 4907 2103 4923
rect 1676 4423 1683 4443
rect 1656 4416 1683 4423
rect 1456 4107 1463 4233
rect 1556 4216 1563 4253
rect 1456 3996 1463 4093
rect 1496 3996 1503 4013
rect 1476 3867 1483 3983
rect 1516 3976 1523 4033
rect 1596 3847 1603 4373
rect 1656 4207 1663 4416
rect 1696 4323 1703 4453
rect 1736 4347 1743 4443
rect 1687 4316 1703 4323
rect 1676 4187 1683 4313
rect 1756 4216 1763 4313
rect 1736 4027 1743 4203
rect 1696 3996 1703 4013
rect 1796 4007 1803 4553
rect 2076 4547 2083 4673
rect 2116 4627 2123 4683
rect 2156 4676 2163 4693
rect 2136 4647 2143 4663
rect 1896 4496 1903 4513
rect 2076 4487 2083 4533
rect 2076 4456 2083 4473
rect 1816 4223 1823 4333
rect 1816 4216 1843 4223
rect 1676 3967 1683 3973
rect 1436 3716 1443 3773
rect 1476 3687 1483 3833
rect 1596 3716 1603 3833
rect 1636 3707 1643 3723
rect 1576 3667 1583 3703
rect 1616 3607 1623 3703
rect 1456 3536 1463 3593
rect 1616 3496 1643 3503
rect 1236 3476 1263 3483
rect 1156 3263 1163 3473
rect 1176 3287 1183 3453
rect 1256 3347 1263 3476
rect 1296 3467 1303 3483
rect 1136 3256 1163 3263
rect 1176 3256 1183 3273
rect 1116 3227 1123 3243
rect 1156 3027 1163 3256
rect 1176 3016 1183 3213
rect 1236 3067 1243 3253
rect 1516 3227 1523 3243
rect 1196 3036 1203 3053
rect 1236 3036 1243 3053
rect 1336 3047 1343 3203
rect 1356 3036 1403 3043
rect 1436 3036 1443 3053
rect 1356 3007 1363 3036
rect 1456 3027 1463 3133
rect 1516 3107 1523 3213
rect 1087 2776 1103 2783
rect 956 2756 983 2763
rect 1036 2756 1063 2763
rect 956 2667 963 2756
rect 1056 2687 1063 2756
rect 256 2536 283 2543
rect 276 2347 283 2536
rect 136 2296 143 2313
rect 156 1807 163 2283
rect 196 1783 203 2233
rect 276 2067 283 2333
rect 316 2276 333 2283
rect 396 2107 403 2293
rect 256 1943 263 2063
rect 396 2056 403 2093
rect 416 2047 423 2313
rect 516 2307 523 2563
rect 676 2556 683 2573
rect 636 2276 663 2283
rect 436 2056 443 2273
rect 636 2267 643 2276
rect 476 2067 483 2263
rect 676 2243 683 2293
rect 756 2247 763 2563
rect 816 2267 823 2563
rect 896 2556 903 2573
rect 936 2556 943 2613
rect 956 2587 963 2653
rect 1076 2527 1083 2773
rect 1156 2763 1163 2893
rect 1136 2756 1163 2763
rect 1236 2723 1243 2993
rect 1516 2867 1523 3093
rect 1536 3003 1543 3253
rect 1616 3227 1623 3496
rect 1656 3147 1663 3653
rect 1696 3407 1703 3813
rect 1716 3787 1723 3973
rect 1776 3807 1783 3953
rect 1736 3503 1743 3553
rect 1776 3527 1783 3793
rect 1796 3787 1803 3993
rect 1816 3743 1823 3913
rect 1836 3887 1843 4216
rect 2136 4203 2143 4533
rect 2176 4487 2183 4663
rect 2216 4247 2223 4693
rect 2236 4607 2243 5436
rect 2256 5287 2263 5413
rect 2276 5387 2283 5393
rect 2316 5156 2323 5193
rect 2336 5087 2343 5143
rect 2296 4683 2303 4733
rect 2296 4676 2313 4683
rect 2356 4676 2363 4713
rect 2336 4627 2343 4663
rect 2336 4476 2343 4513
rect 2316 4387 2323 4463
rect 2356 4456 2363 4513
rect 2376 4507 2383 4653
rect 2416 4647 2423 5833
rect 2456 5727 2463 5903
rect 2496 5896 2503 5913
rect 2447 5656 2463 5663
rect 2436 5627 2443 5653
rect 2536 5567 2543 5993
rect 2436 5456 2443 5513
rect 2436 4943 2443 5413
rect 2576 5387 2583 6056
rect 2756 6007 2763 6123
rect 2756 5947 2763 5993
rect 2616 5647 2623 5893
rect 2636 5667 2643 5673
rect 2676 5667 2683 5883
rect 2436 4936 2463 4943
rect 2376 4423 2383 4493
rect 2356 4416 2383 4423
rect 1856 4187 1863 4203
rect 2136 4196 2163 4203
rect 1916 3996 1923 4033
rect 1956 4007 1963 4133
rect 2156 4016 2163 4033
rect 1816 3736 1843 3743
rect 1796 3567 1803 3723
rect 1836 3716 1843 3736
rect 1876 3703 1883 3993
rect 1936 3927 1943 3983
rect 1936 3827 1943 3913
rect 1996 3887 2003 3963
rect 2136 3847 2143 3973
rect 2196 3827 2203 3873
rect 1856 3696 1883 3703
rect 1856 3587 1863 3696
rect 1936 3647 1943 3773
rect 1976 3736 2003 3743
rect 1976 3707 1983 3736
rect 1936 3627 1943 3633
rect 1796 3527 1803 3553
rect 1836 3516 1863 3523
rect 1896 3516 1903 3533
rect 1936 3516 1943 3613
rect 1776 3507 1783 3513
rect 1716 3496 1743 3503
rect 1616 3003 1623 3053
rect 1536 2996 1563 3003
rect 1596 2996 1623 3003
rect 1536 2843 1543 2996
rect 1516 2836 1543 2843
rect 1236 2716 1263 2723
rect 1396 2707 1403 2733
rect 1436 2667 1443 2763
rect 1516 2756 1523 2836
rect 1556 2667 1563 2853
rect 1696 2727 1703 3393
rect 1836 3247 1843 3516
rect 2056 3507 2063 3723
rect 2076 3496 2083 3693
rect 2116 3496 2123 3533
rect 2156 3483 2163 3773
rect 2196 3716 2203 3813
rect 2176 3587 2183 3703
rect 2216 3667 2223 3703
rect 2136 3476 2163 3483
rect 1756 3127 1763 3223
rect 1776 3067 1783 3203
rect 1796 3056 1803 3133
rect 1836 3023 1843 3113
rect 1816 3016 1843 3023
rect 1896 3016 1903 3353
rect 1956 3256 1963 3333
rect 1976 3247 1983 3473
rect 2116 3427 2123 3453
rect 1996 3267 2003 3273
rect 1996 3007 2003 3253
rect 2116 3236 2123 3413
rect 2176 3243 2183 3513
rect 2156 3236 2183 3243
rect 2016 3056 2023 3153
rect 2096 3147 2103 3223
rect 2136 3167 2143 3223
rect 2196 3016 2203 3093
rect 1976 2747 1983 2893
rect 1716 2687 1723 2743
rect 1936 2727 1943 2743
rect 1736 2707 1743 2723
rect 1936 2687 1943 2713
rect 2056 2707 2063 2713
rect 2076 2667 2083 2743
rect 1176 2576 1183 2593
rect 1136 2543 1143 2573
rect 1136 2536 1163 2543
rect 1556 2536 1563 2653
rect 1656 2543 1663 2653
rect 1836 2576 1863 2583
rect 1836 2547 1843 2576
rect 1636 2536 1663 2543
rect 1716 2536 1743 2543
rect 1196 2407 1203 2533
rect 856 2296 883 2303
rect 856 2267 863 2296
rect 836 2247 843 2263
rect 256 1936 283 1943
rect 176 1776 203 1783
rect 156 1667 163 1763
rect 156 1547 163 1583
rect 256 1576 263 1913
rect 276 1587 283 1936
rect 356 1767 363 1823
rect 376 1667 383 1803
rect 456 1747 463 2043
rect 496 1807 503 2243
rect 656 2236 683 2243
rect 596 2076 603 2093
rect 656 2076 663 2236
rect 576 1783 583 2073
rect 696 1823 703 2093
rect 856 2087 863 2253
rect 996 2047 1003 2063
rect 796 1827 803 2043
rect 676 1816 703 1823
rect 556 1776 583 1783
rect 536 1727 543 1763
rect 356 1616 383 1623
rect 216 1547 223 1563
rect 36 1336 43 1433
rect 96 1323 103 1533
rect 76 1316 103 1323
rect 136 1116 143 1153
rect 176 1147 183 1313
rect 356 1307 363 1616
rect 376 1363 383 1573
rect 596 1567 603 1813
rect 676 1787 683 1816
rect 1096 1823 1103 2263
rect 1296 2247 1303 2263
rect 1136 2027 1143 2093
rect 1196 2087 1203 2233
rect 1236 2047 1243 2093
rect 1016 1816 1043 1823
rect 1076 1816 1103 1823
rect 1256 1816 1263 2093
rect 1316 2043 1323 2293
rect 1436 2276 1443 2333
rect 1316 2036 1343 2043
rect 1416 2027 1423 2083
rect 1516 2083 1523 2113
rect 1556 2083 1563 2493
rect 1696 2443 1703 2523
rect 1676 2436 1703 2443
rect 1576 2276 1583 2293
rect 1496 2076 1523 2083
rect 1536 2076 1563 2083
rect 716 1787 723 1803
rect 796 1647 803 1813
rect 856 1767 863 1793
rect 896 1663 903 1733
rect 916 1707 923 1783
rect 1016 1767 1023 1816
rect 896 1656 923 1663
rect 656 1583 663 1613
rect 916 1596 923 1656
rect 636 1576 663 1583
rect 487 1436 493 1443
rect 376 1356 403 1363
rect 396 1323 403 1356
rect 616 1327 623 1573
rect 376 1316 403 1323
rect 456 1316 483 1323
rect 196 1167 203 1283
rect 96 647 103 1093
rect 196 843 203 1093
rect 196 836 223 843
rect 96 367 103 633
rect 136 616 143 823
rect 156 636 163 653
rect 176 587 183 623
rect 216 587 223 836
rect 236 807 243 1133
rect 396 867 403 1316
rect 476 1107 483 1316
rect 476 1083 483 1093
rect 476 1076 503 1083
rect 536 1067 543 1083
rect 596 1067 603 1303
rect 676 1287 683 1303
rect 696 1127 703 1313
rect 716 1096 723 1313
rect 796 1307 803 1433
rect 896 1367 903 1533
rect 896 1336 903 1353
rect 836 1316 883 1323
rect 876 1287 883 1316
rect 936 1307 943 1323
rect 736 1087 743 1093
rect 256 667 263 853
rect 336 807 343 823
rect 127 496 143 503
rect 136 367 143 496
rect 107 356 123 363
rect 156 356 163 373
rect 176 156 183 553
rect 276 387 283 673
rect 316 623 323 713
rect 376 687 383 823
rect 396 807 403 833
rect 476 787 483 853
rect 356 656 383 663
rect 316 616 343 623
rect 376 567 383 656
rect 396 567 403 623
rect 476 616 483 773
rect 496 687 503 1053
rect 696 1047 703 1083
rect 536 836 543 1033
rect 756 836 763 853
rect 796 836 803 1113
rect 856 1107 863 1283
rect 876 1116 883 1273
rect 916 1127 923 1273
rect 956 1107 963 1553
rect 1036 1347 1043 1613
rect 1056 1387 1063 1803
rect 1216 1783 1223 1793
rect 1216 1776 1243 1783
rect 1296 1767 1303 1783
rect 1396 1763 1403 2013
rect 1436 1796 1463 1803
rect 1396 1756 1423 1763
rect 1076 1607 1083 1713
rect 1456 1667 1463 1796
rect 1076 1563 1083 1593
rect 1276 1576 1283 1593
rect 1316 1576 1323 1653
rect 1476 1616 1483 2073
rect 1076 1556 1103 1563
rect 1336 1487 1343 1563
rect 1056 1143 1063 1283
rect 1236 1147 1243 1323
rect 1316 1316 1343 1323
rect 1336 1167 1343 1316
rect 1056 1136 1083 1143
rect 1036 1116 1043 1133
rect 1076 1116 1083 1136
rect 856 1067 863 1093
rect 516 807 523 823
rect 556 767 563 823
rect 596 727 603 823
rect 856 807 863 1053
rect 936 856 943 953
rect 996 847 1003 1113
rect 1056 1087 1063 1103
rect 1096 1087 1103 1103
rect 1016 836 1023 1053
rect 656 656 663 753
rect 756 616 783 623
rect 756 487 763 616
rect 216 376 243 383
rect 236 127 243 376
rect 376 187 383 323
rect 256 176 283 183
rect 256 27 263 176
rect 476 156 483 173
rect 496 136 503 233
rect 516 147 523 393
rect 636 356 643 373
rect 676 267 683 473
rect 796 356 803 573
rect 856 387 863 753
rect 856 363 863 373
rect 836 356 863 363
rect 876 347 883 673
rect 896 367 903 773
rect 956 636 983 643
rect 1016 636 1023 673
rect 1036 667 1043 853
rect 1076 667 1083 953
rect 1116 843 1123 1033
rect 1216 967 1223 1113
rect 1236 1047 1243 1133
rect 1256 1096 1283 1103
rect 1256 1067 1263 1096
rect 1436 1047 1443 1353
rect 1456 1167 1463 1213
rect 1456 1136 1463 1153
rect 1516 1147 1523 2076
rect 1556 1783 1563 2076
rect 1656 1967 1663 2043
rect 1676 1967 1683 2436
rect 1716 2403 1723 2536
rect 2016 2536 2043 2543
rect 1707 2396 1723 2403
rect 1696 2056 1703 2393
rect 1876 2276 1883 2313
rect 2016 2307 2023 2536
rect 1816 2096 1823 2273
rect 1996 2067 2003 2293
rect 1576 1807 1583 1913
rect 1676 1816 1683 1953
rect 1816 1867 1823 2053
rect 1556 1776 1583 1783
rect 1556 1316 1563 1473
rect 1536 1247 1543 1303
rect 1536 1127 1543 1233
rect 1576 1187 1583 1776
rect 1596 1627 1603 1783
rect 1616 1567 1623 1633
rect 1636 1623 1643 1783
rect 1816 1763 1823 1813
rect 2036 1803 2043 2053
rect 2076 1927 2083 2063
rect 2096 1847 2103 2753
rect 2176 2727 2183 2993
rect 2216 2747 2223 3533
rect 2236 3027 2243 3493
rect 2216 2607 2223 2733
rect 2136 2543 2143 2573
rect 2116 2536 2143 2543
rect 2016 1796 2043 1803
rect 2036 1787 2043 1796
rect 1816 1756 1843 1763
rect 1636 1616 1663 1623
rect 1656 1547 1663 1616
rect 1816 1563 1823 1613
rect 1856 1576 1863 1693
rect 1816 1556 1843 1563
rect 1876 1547 1883 1563
rect 1956 1347 1963 1593
rect 2016 1576 2023 1633
rect 2036 1556 2043 1653
rect 2116 1647 2123 2053
rect 2136 1927 2143 2243
rect 2156 1827 2163 2273
rect 2236 2247 2243 2933
rect 2256 2887 2263 3833
rect 2276 3516 2283 3573
rect 2316 3547 2323 4213
rect 2356 4147 2363 4416
rect 2376 4207 2383 4273
rect 2416 4227 2423 4613
rect 2436 4207 2443 4793
rect 2456 4547 2463 4936
rect 2516 4867 2523 4943
rect 2476 4667 2483 4713
rect 2456 4147 2463 4183
rect 2436 3983 2443 4013
rect 2416 3976 2443 3983
rect 2476 3847 2483 4633
rect 2516 4587 2523 4703
rect 2536 4607 2543 4683
rect 2496 4476 2503 4493
rect 2536 4476 2543 4513
rect 2356 3687 2363 3833
rect 2396 3716 2403 3793
rect 2296 3467 2303 3503
rect 2356 3467 2363 3533
rect 2296 3387 2303 3453
rect 2376 3243 2383 3703
rect 2396 3267 2403 3483
rect 2376 3236 2403 3243
rect 2376 3223 2383 3236
rect 2316 3127 2323 3223
rect 2356 3216 2383 3223
rect 2316 3027 2323 3113
rect 2336 2967 2343 3203
rect 2416 3187 2423 3613
rect 2436 3496 2443 3673
rect 2456 3647 2463 3703
rect 2496 3627 2503 4353
rect 2516 4207 2523 4463
rect 2516 3887 2523 4193
rect 2416 3056 2423 3173
rect 2416 3016 2443 3023
rect 2336 2687 2343 2743
rect 2296 2543 2303 2553
rect 2276 2536 2303 2543
rect 2356 2327 2363 2453
rect 2356 2276 2363 2313
rect 2196 2096 2223 2103
rect 2196 1807 2203 2096
rect 2276 2063 2283 2263
rect 2236 2056 2283 2063
rect 2356 2047 2363 2073
rect 2136 1776 2163 1783
rect 2136 1627 2143 1776
rect 2056 1576 2063 1593
rect 1736 1336 1763 1343
rect 1736 1287 1743 1336
rect 1996 1336 2023 1343
rect 2016 1327 2023 1336
rect 1776 1207 1783 1323
rect 1816 1267 1823 1323
rect 1976 1307 1983 1323
rect 2076 1187 2083 1563
rect 2136 1336 2163 1343
rect 2096 1303 2103 1333
rect 2136 1327 2143 1336
rect 2096 1296 2123 1303
rect 2136 1287 2143 1313
rect 2176 1267 2183 1303
rect 1676 1136 1703 1143
rect 1476 1087 1483 1103
rect 1556 1096 1583 1103
rect 1536 1047 1543 1083
rect 1436 863 1443 1033
rect 1556 967 1563 1096
rect 1416 856 1443 863
rect 1096 836 1123 843
rect 1096 787 1103 836
rect 956 587 963 636
rect 1036 627 1043 653
rect 1176 643 1183 733
rect 1276 647 1283 803
rect 1296 747 1303 853
rect 1156 636 1183 643
rect 1176 603 1183 636
rect 1316 616 1323 653
rect 1376 647 1383 673
rect 1416 663 1423 856
rect 1476 847 1483 953
rect 1396 656 1423 663
rect 1156 596 1183 603
rect 596 136 603 253
rect 716 176 723 293
rect 816 247 823 343
rect 896 147 903 353
rect 956 287 963 473
rect 976 183 983 323
rect 956 176 983 183
rect 956 27 963 176
rect 996 143 1003 313
rect 976 136 1003 143
rect 1056 123 1063 593
rect 1156 407 1163 596
rect 1356 587 1363 623
rect 1396 607 1403 656
rect 1407 596 1423 603
rect 1156 356 1163 393
rect 1396 367 1403 573
rect 1196 347 1203 363
rect 1176 307 1183 343
rect 1356 327 1363 363
rect 1436 347 1443 633
rect 1456 616 1463 833
rect 1556 427 1563 833
rect 1576 656 1583 813
rect 1596 787 1603 843
rect 1636 836 1643 853
rect 1676 827 1683 1136
rect 1656 727 1663 823
rect 1716 567 1723 713
rect 1556 367 1563 413
rect 1716 367 1723 473
rect 1536 327 1543 333
rect 1356 287 1363 313
rect 1076 136 1083 273
rect 1596 247 1603 363
rect 1596 147 1603 233
rect 1616 136 1623 333
rect 1736 227 1743 853
rect 1756 627 1763 933
rect 1796 847 1803 993
rect 1856 947 1863 1133
rect 1876 1096 1883 1133
rect 1836 836 1863 843
rect 1776 807 1783 823
rect 1776 647 1783 793
rect 1816 787 1823 823
rect 1856 787 1863 836
rect 1856 623 1863 773
rect 1976 636 1983 1173
rect 2076 1116 2103 1123
rect 2056 867 2063 1113
rect 2036 836 2043 853
rect 2076 807 2083 1116
rect 2156 1107 2163 1133
rect 2116 1007 2123 1103
rect 2196 923 2203 1793
rect 2276 1747 2283 1783
rect 2216 1627 2223 1633
rect 2216 1596 2223 1613
rect 2256 1596 2283 1603
rect 2276 1547 2283 1596
rect 2276 1367 2283 1533
rect 2276 1307 2283 1353
rect 2356 1327 2363 2033
rect 2376 1987 2383 2753
rect 2416 2267 2423 3016
rect 2456 2707 2463 3453
rect 2536 3367 2543 4253
rect 2556 3647 2563 4413
rect 2596 4267 2603 5513
rect 2616 5467 2623 5553
rect 2616 5447 2623 5453
rect 2616 5416 2623 5433
rect 2616 4427 2623 5213
rect 2636 4407 2643 5653
rect 2736 5623 2743 5653
rect 2656 5616 2683 5623
rect 2716 5616 2743 5623
rect 2656 5567 2663 5616
rect 2676 5423 2683 5573
rect 2676 5416 2703 5423
rect 2676 5147 2683 5163
rect 2716 5156 2723 5253
rect 2756 5143 2763 5793
rect 2776 5487 2783 6156
rect 2796 5727 2803 6353
rect 2696 5127 2703 5143
rect 2736 5136 2763 5143
rect 2756 5047 2763 5136
rect 2656 4956 2663 5013
rect 2696 4956 2703 4973
rect 2676 4907 2683 4943
rect 2736 4927 2743 5013
rect 2676 4487 2683 4893
rect 2716 4687 2723 4703
rect 2756 4696 2763 5013
rect 2716 4483 2723 4553
rect 2736 4503 2743 4683
rect 2776 4627 2783 5473
rect 2796 5427 2803 5713
rect 2816 5527 2823 6153
rect 2836 6116 2843 6433
rect 2856 5936 2863 6093
rect 2876 6087 2883 6436
rect 2916 6416 2923 6433
rect 2896 6063 2903 6313
rect 2956 6307 2963 6553
rect 2876 6056 2903 6063
rect 2856 5807 2863 5893
rect 2876 5647 2883 6056
rect 2916 5907 2923 6133
rect 2936 5896 2943 6233
rect 2896 5876 2923 5883
rect 2816 5436 2823 5493
rect 2796 5207 2803 5413
rect 2896 5287 2903 5623
rect 2916 5407 2923 5876
rect 2936 5387 2943 5433
rect 2896 5176 2903 5193
rect 2816 4907 2823 4973
rect 2916 4927 2923 5373
rect 2936 5127 2943 5143
rect 2736 4496 2763 4503
rect 2696 4476 2723 4483
rect 2756 4476 2763 4496
rect 2636 4207 2643 4373
rect 2696 4347 2703 4476
rect 2776 4443 2783 4463
rect 2836 4447 2843 4893
rect 2856 4867 2863 4923
rect 2896 4883 2903 4913
rect 2876 4876 2903 4883
rect 2856 4587 2863 4693
rect 2776 4436 2803 4443
rect 2596 4176 2623 4183
rect 2596 4167 2603 4176
rect 2656 4167 2663 4183
rect 2576 3996 2583 4033
rect 2616 4016 2623 4153
rect 2656 3987 2663 4033
rect 2636 3947 2643 3983
rect 2676 3843 2683 4193
rect 2656 3836 2683 3843
rect 2616 3667 2623 3723
rect 2656 3716 2663 3836
rect 2636 3667 2643 3703
rect 2676 3687 2683 3703
rect 2556 3536 2563 3573
rect 2696 3487 2703 4233
rect 2716 3783 2723 4433
rect 2736 3807 2743 4193
rect 2756 4187 2763 4333
rect 2796 4207 2803 4436
rect 2836 4196 2843 4273
rect 2856 4227 2863 4573
rect 2776 4163 2783 4183
rect 2756 4156 2783 4163
rect 2756 4027 2763 4156
rect 2816 4127 2823 4183
rect 2776 4016 2783 4033
rect 2756 3996 2763 4013
rect 2796 4007 2803 4093
rect 2776 3967 2783 3973
rect 2716 3776 2743 3783
rect 2716 3567 2723 3673
rect 2736 3627 2743 3776
rect 2776 3723 2783 3953
rect 2836 3947 2843 3993
rect 2876 3927 2883 4876
rect 2896 4696 2903 4853
rect 2936 4703 2943 4993
rect 2956 4907 2963 6293
rect 2976 6147 2983 6733
rect 2996 6127 3003 6573
rect 3016 6567 3023 7036
rect 3056 6867 3063 7353
rect 3076 7227 3083 7396
rect 3116 7376 3123 7393
rect 3136 7387 3143 7556
rect 3176 7507 3183 8043
rect 3196 7607 3203 8073
rect 3356 8047 3363 8303
rect 3396 8207 3403 8303
rect 3216 7707 3223 8033
rect 3376 7927 3383 8153
rect 3416 8147 3423 8333
rect 3456 8187 3463 8493
rect 3516 8483 3523 8503
rect 3556 8496 3583 8503
rect 3516 8476 3543 8483
rect 3516 8316 3523 8433
rect 3536 8367 3543 8476
rect 3496 8287 3503 8313
rect 3576 8296 3583 8313
rect 3536 8187 3543 8293
rect 3236 7847 3243 7893
rect 3256 7807 3263 7853
rect 3316 7807 3323 7823
rect 3096 7367 3103 7373
rect 3136 7356 3163 7363
rect 3156 7327 3163 7356
rect 3076 7027 3083 7213
rect 3076 6787 3083 6993
rect 3116 6747 3123 7153
rect 3136 6847 3143 7173
rect 3196 7167 3203 7573
rect 3236 7556 3243 7773
rect 3256 7587 3263 7793
rect 3216 7307 3223 7543
rect 3176 7067 3183 7083
rect 3176 6747 3183 6843
rect 3236 6707 3243 7513
rect 3276 7487 3283 7563
rect 3296 7463 3303 7593
rect 3316 7567 3323 7693
rect 3336 7527 3343 7833
rect 3376 7767 3383 7823
rect 3356 7627 3363 7693
rect 3356 7487 3363 7593
rect 3276 7456 3303 7463
rect 3256 7087 3263 7113
rect 3016 6327 3023 6553
rect 3036 6407 3043 6513
rect 3056 6387 3063 6433
rect 3116 6396 3123 6413
rect 3096 6347 3103 6383
rect 3136 6376 3143 6393
rect 3096 6267 3103 6333
rect 3036 6107 3043 6123
rect 2976 6087 2983 6103
rect 3016 6007 3023 6033
rect 3036 5807 3043 6053
rect 3056 6047 3063 6113
rect 3156 6067 3163 6433
rect 3176 6267 3183 6563
rect 3196 6167 3203 6693
rect 3276 6447 3283 7456
rect 3336 7376 3343 7413
rect 3356 7187 3363 7343
rect 3296 7067 3303 7133
rect 3376 7087 3383 7613
rect 3396 7547 3403 7893
rect 3416 7576 3423 7773
rect 3436 7607 3443 7913
rect 3456 7767 3463 8173
rect 3547 8156 3553 8163
rect 3516 8056 3523 8153
rect 3596 8147 3603 8793
rect 3656 8523 3663 8693
rect 3676 8607 3683 8763
rect 3696 8707 3703 8773
rect 3716 8747 3723 8993
rect 3756 8947 3763 8963
rect 3756 8867 3763 8933
rect 3816 8847 3823 8993
rect 3856 8963 3863 9353
rect 3876 9047 3883 9473
rect 3916 9287 3923 9483
rect 3936 9027 3943 9633
rect 3996 9607 4003 9753
rect 4196 9736 4203 9873
rect 3956 9147 3963 9573
rect 3956 9007 3963 9133
rect 3856 8956 3883 8963
rect 3656 8516 3683 8523
rect 3716 8287 3723 8523
rect 3756 8487 3763 8813
rect 3816 8796 3823 8833
rect 3876 8827 3883 8956
rect 3776 8607 3783 8793
rect 3876 8787 3883 8793
rect 3836 8727 3843 8783
rect 3736 8296 3763 8303
rect 3756 8207 3763 8296
rect 3756 8187 3763 8193
rect 3736 8167 3743 8173
rect 3476 7927 3483 8043
rect 3496 7847 3503 7973
rect 3476 7816 3503 7823
rect 3396 7127 3403 7473
rect 3416 7087 3423 7353
rect 3296 6647 3303 6893
rect 3316 6623 3323 7073
rect 3436 7063 3443 7533
rect 3476 7507 3483 7816
rect 3516 7807 3523 7953
rect 3536 7787 3543 8133
rect 3636 8023 3643 8053
rect 3716 8023 3723 8133
rect 3636 8016 3663 8023
rect 3696 8016 3723 8023
rect 3656 7967 3663 8016
rect 3676 7856 3683 7973
rect 3736 7907 3743 8153
rect 3756 7987 3763 8173
rect 3776 7867 3783 8273
rect 3796 8203 3803 8493
rect 3856 8483 3863 8533
rect 3896 8516 3923 8523
rect 3916 8507 3923 8516
rect 3856 8476 3883 8483
rect 3816 8227 3823 8333
rect 3796 8196 3823 8203
rect 3776 7816 3803 7823
rect 3776 7687 3783 7816
rect 3816 7783 3823 8196
rect 3836 7987 3843 8433
rect 3887 8316 3903 8323
rect 3936 8316 3943 8393
rect 3956 8367 3963 8813
rect 3976 8767 3983 9553
rect 3996 9476 4023 9483
rect 4156 9476 4163 9493
rect 4016 9367 4023 9476
rect 4136 9407 4143 9463
rect 4176 9447 4183 9463
rect 4216 9447 4223 10293
rect 4236 10187 4243 10213
rect 4236 9956 4243 10173
rect 4256 9947 4263 10233
rect 4256 9667 4263 9813
rect 4016 9296 4043 9303
rect 4016 9267 4023 9296
rect 4056 9247 4063 9263
rect 4136 9256 4163 9263
rect 4116 9227 4123 9243
rect 4016 9003 4023 9033
rect 4016 8996 4043 9003
rect 4016 8796 4043 8803
rect 4036 8687 4043 8796
rect 4116 8767 4123 9213
rect 4136 9127 4143 9256
rect 4256 9187 4263 9653
rect 4276 9527 4283 9743
rect 4296 9507 4303 10973
rect 4316 10456 4323 10653
rect 4356 10467 4363 11013
rect 4376 10947 4383 11193
rect 4396 11087 4403 11173
rect 4416 11027 4423 11553
rect 4436 11387 4443 11693
rect 4476 11567 4483 11663
rect 4516 11647 4523 11663
rect 4476 11403 4483 11553
rect 4456 11396 4483 11403
rect 4536 11383 4543 11553
rect 4556 11467 4563 11793
rect 4716 11767 4723 11843
rect 4756 11827 4763 11913
rect 5076 11896 5103 11903
rect 5136 11896 5143 11913
rect 4896 11876 4903 11893
rect 4596 11607 4603 11753
rect 4576 11507 4583 11593
rect 4516 11376 4543 11383
rect 4496 11163 4503 11233
rect 4616 11216 4623 11653
rect 4716 11567 4723 11643
rect 4736 11383 4743 11433
rect 4656 11183 4663 11233
rect 4636 11176 4663 11183
rect 4436 11147 4443 11163
rect 4476 11156 4503 11163
rect 4676 11147 4683 11383
rect 4716 11376 4743 11383
rect 4756 11367 4763 11813
rect 4876 11807 4883 11863
rect 4876 11656 4883 11753
rect 4896 11636 4903 11693
rect 4956 11687 4963 11863
rect 4976 11787 4983 11893
rect 5076 11847 5083 11896
rect 5256 11876 5283 11883
rect 5076 11767 5083 11833
rect 5116 11827 5123 11873
rect 5236 11807 5243 11873
rect 5256 11827 5263 11876
rect 5456 11847 5463 11893
rect 5487 11836 5503 11843
rect 4916 11656 4923 11673
rect 4936 11627 4943 11643
rect 4976 11627 4983 11713
rect 5116 11656 5123 11673
rect 5096 11627 5103 11643
rect 4816 11383 4823 11413
rect 4816 11376 4843 11383
rect 4796 11196 4803 11333
rect 4856 11307 4863 11363
rect 4436 11087 4443 11133
rect 4376 10903 4383 10913
rect 4376 10896 4403 10903
rect 4456 10903 4463 11033
rect 4476 11007 4483 11073
rect 4447 10896 4463 10903
rect 4416 10847 4423 10883
rect 4476 10727 4483 10993
rect 4516 10867 4523 10953
rect 4476 10463 4483 10713
rect 4536 10683 4543 11073
rect 4596 10887 4603 10903
rect 4596 10723 4603 10873
rect 4636 10867 4643 10903
rect 4596 10716 4623 10723
rect 4616 10683 4623 10716
rect 4536 10676 4563 10683
rect 4596 10676 4623 10683
rect 4476 10456 4503 10463
rect 4536 10456 4543 10676
rect 4636 10647 4643 10853
rect 4316 9927 4323 10233
rect 4336 10227 4343 10443
rect 4356 10216 4363 10253
rect 4416 10236 4423 10373
rect 4376 9956 4383 9993
rect 4396 9927 4403 9943
rect 4416 9767 4423 9933
rect 4456 9756 4463 9773
rect 4476 9767 4483 10456
rect 4516 10387 4523 10443
rect 4536 10236 4543 10333
rect 4576 10236 4583 10253
rect 4596 10216 4603 10233
rect 4636 10203 4643 10413
rect 4656 10407 4663 11053
rect 4756 10916 4783 10923
rect 4756 10883 4763 10916
rect 4936 10903 4943 11193
rect 4956 11043 4963 11333
rect 5016 11327 5023 11383
rect 5096 11367 5103 11613
rect 5136 11407 5143 11643
rect 4996 11187 5003 11213
rect 4976 11067 4983 11163
rect 5016 11156 5023 11253
rect 5036 11176 5043 11193
rect 4956 11036 4983 11043
rect 4976 10916 4983 11036
rect 5056 10927 5063 11193
rect 5076 10947 5083 11173
rect 5136 11127 5143 11393
rect 5216 11227 5223 11363
rect 5236 11347 5243 11383
rect 5256 11347 5263 11643
rect 5296 11507 5303 11643
rect 5156 11196 5183 11203
rect 5176 11127 5183 11196
rect 5216 11167 5223 11213
rect 5176 11107 5183 11113
rect 4936 10896 4963 10903
rect 4756 10876 4783 10883
rect 4756 10736 4763 10793
rect 4736 10716 4743 10733
rect 4776 10716 4783 10876
rect 5136 10883 5143 11053
rect 5316 11047 5323 11833
rect 5416 11707 5423 11833
rect 5516 11803 5523 11863
rect 5496 11796 5523 11803
rect 5656 11856 5683 11863
rect 5436 11707 5443 11733
rect 5496 11703 5503 11796
rect 5476 11696 5503 11703
rect 5436 11676 5443 11693
rect 5476 11676 5483 11696
rect 5516 11676 5523 11773
rect 5656 11687 5663 11856
rect 5696 11747 5703 11843
rect 5716 11787 5723 11863
rect 5336 11587 5343 11653
rect 5456 11507 5463 11663
rect 5636 11656 5663 11663
rect 5556 11627 5563 11653
rect 5596 11587 5603 11653
rect 5376 11347 5383 11383
rect 5416 11367 5423 11383
rect 5396 11327 5403 11363
rect 5356 11167 5363 11183
rect 5396 10903 5403 11313
rect 5436 11227 5443 11493
rect 5636 11467 5643 11656
rect 5716 11607 5723 11643
rect 5616 11416 5633 11423
rect 5496 11247 5503 11413
rect 4696 10423 4703 10713
rect 4676 10416 4703 10423
rect 4676 10367 4683 10416
rect 4676 10216 4703 10223
rect 4636 10196 4663 10203
rect 4596 9956 4603 10153
rect 4676 10087 4683 10216
rect 4716 9967 4723 10393
rect 4756 10347 4763 10693
rect 4796 10167 4803 10873
rect 4836 10847 4843 10883
rect 5136 10876 5183 10883
rect 5196 10787 5203 10903
rect 5336 10847 5343 10903
rect 5376 10896 5403 10903
rect 4956 10736 4983 10743
rect 4836 10696 4863 10703
rect 4816 10427 4823 10683
rect 4836 10567 4843 10696
rect 4856 10456 4863 10513
rect 4956 10407 4963 10736
rect 5256 10703 5263 10733
rect 5356 10707 5363 10883
rect 5156 10696 5183 10703
rect 5236 10696 5263 10703
rect 4376 9507 4383 9753
rect 4516 9747 4523 9953
rect 4616 9927 4623 9943
rect 4696 9776 4703 9913
rect 4796 9887 4803 9943
rect 4916 9927 4923 10073
rect 4976 9956 4983 10533
rect 5036 10427 5043 10473
rect 5116 10436 5123 10453
rect 5156 10423 5163 10653
rect 4996 10216 5003 10273
rect 5036 10207 5043 10413
rect 5056 10387 5063 10423
rect 5096 10407 5103 10423
rect 5136 10416 5163 10423
rect 5056 10367 5063 10373
rect 5136 10267 5143 10416
rect 5176 10287 5183 10696
rect 5336 10467 5343 10673
rect 5396 10667 5403 10703
rect 5476 10687 5483 11193
rect 5496 11187 5503 11233
rect 5576 11203 5583 11373
rect 5596 11367 5603 11403
rect 5636 11387 5643 11413
rect 5716 11387 5723 11493
rect 5776 11416 5783 11913
rect 5796 11427 5803 11933
rect 6016 11863 6023 11893
rect 5856 11787 5863 11863
rect 5876 11787 5883 11843
rect 5896 11807 5903 11863
rect 6016 11856 6043 11863
rect 6076 11807 6083 11863
rect 6096 11847 6103 11913
rect 6216 11876 6223 12013
rect 6696 11876 6723 11883
rect 6516 11827 6523 11863
rect 6556 11807 6563 11863
rect 6676 11827 6683 11843
rect 6716 11827 6723 11876
rect 5936 11647 5943 11673
rect 5856 11587 5863 11643
rect 5896 11627 5903 11643
rect 5936 11627 5943 11633
rect 5896 11587 5903 11613
rect 5896 11436 5963 11443
rect 5896 11407 5903 11436
rect 5956 11416 5963 11436
rect 5976 11407 5983 11793
rect 6216 11696 6293 11703
rect 6216 11687 6223 11696
rect 6236 11667 6243 11673
rect 6056 11487 6063 11663
rect 6096 11656 6123 11663
rect 5756 11387 5763 11403
rect 6056 11387 6063 11473
rect 6116 11447 6123 11656
rect 6236 11643 6243 11653
rect 6236 11636 6263 11643
rect 6296 11607 6303 11633
rect 6256 11416 6283 11423
rect 6316 11416 6323 11753
rect 6336 11627 6343 11693
rect 5756 11367 5763 11373
rect 6076 11363 6083 11413
rect 6116 11396 6143 11403
rect 6076 11356 6103 11363
rect 6136 11347 6143 11396
rect 5736 11267 5743 11333
rect 5576 11196 5603 11203
rect 5696 11196 5703 11213
rect 5736 11196 5743 11253
rect 5516 11176 5523 11193
rect 5536 10887 5543 11113
rect 5596 10987 5603 11196
rect 5756 11127 5763 11213
rect 5976 11196 6003 11203
rect 5916 11167 5923 11173
rect 5956 11167 5963 11183
rect 5796 10927 5803 10953
rect 5656 10847 5663 10903
rect 5696 10887 5703 10903
rect 5796 10883 5803 10913
rect 5856 10903 5863 10933
rect 5876 10916 5883 10973
rect 5956 10947 5963 11153
rect 5836 10896 5863 10903
rect 5936 10887 5943 10933
rect 5796 10876 5823 10883
rect 5956 10847 5963 10933
rect 5596 10683 5603 10833
rect 5656 10687 5663 10833
rect 5996 10787 6003 11196
rect 6096 11196 6103 11273
rect 6016 11107 6023 11193
rect 6156 11176 6163 11253
rect 6176 11087 6183 11273
rect 6016 10887 6023 10903
rect 6056 10847 6063 10903
rect 6096 10827 6103 10913
rect 6136 10767 6143 10833
rect 5756 10716 5763 10733
rect 5796 10716 5823 10723
rect 5776 10687 5783 10703
rect 5576 10676 5603 10683
rect 5656 10547 5663 10673
rect 5816 10667 5823 10716
rect 5876 10696 5903 10703
rect 5396 10456 5403 10473
rect 5336 10436 5343 10453
rect 5276 10347 5283 10423
rect 5316 10407 5323 10423
rect 5276 10327 5283 10333
rect 5436 10307 5443 10443
rect 5736 10387 5743 10443
rect 5236 10256 5243 10293
rect 5036 9976 5043 10193
rect 4956 9907 4963 9943
rect 4476 9736 4503 9743
rect 4316 9496 4343 9503
rect 4276 9296 4283 9453
rect 4296 9427 4303 9493
rect 4316 9367 4323 9496
rect 4496 9487 4503 9736
rect 4576 9736 4603 9743
rect 4876 9736 4883 9753
rect 4536 9707 4543 9723
rect 4516 9496 4523 9513
rect 4456 9256 4463 9273
rect 4276 9187 4283 9233
rect 4256 9023 4263 9173
rect 4256 9016 4283 9023
rect 4276 8983 4283 9016
rect 4036 8507 4043 8573
rect 4056 8536 4063 8573
rect 4096 8543 4103 8653
rect 4096 8536 4123 8543
rect 3976 8316 4003 8323
rect 3876 8267 3883 8313
rect 3856 8056 3863 8253
rect 3916 8207 3923 8303
rect 3956 8227 3963 8303
rect 3956 8147 3963 8213
rect 3936 8043 3943 8073
rect 3876 8027 3883 8043
rect 3916 8036 3943 8043
rect 3796 7776 3823 7783
rect 3456 7327 3463 7413
rect 3476 7356 3483 7453
rect 3536 7427 3543 7593
rect 3556 7347 3563 7553
rect 3496 7327 3503 7343
rect 3396 7047 3403 7063
rect 3416 7056 3443 7063
rect 3356 6927 3363 7013
rect 3336 6876 3343 6893
rect 3316 6616 3343 6623
rect 3356 6467 3363 6863
rect 3376 6607 3383 6713
rect 3296 6376 3303 6393
rect 3276 6347 3283 6363
rect 3316 6343 3323 6363
rect 3296 6336 3323 6343
rect 3176 6003 3183 6113
rect 3196 6027 3203 6123
rect 3216 6007 3223 6103
rect 3256 6087 3263 6103
rect 3276 6063 3283 6173
rect 3256 6056 3283 6063
rect 3176 5996 3203 6003
rect 3056 5936 3063 5973
rect 3196 5843 3203 5996
rect 3236 5896 3243 5933
rect 3196 5836 3223 5843
rect 2976 5347 2983 5793
rect 3056 5656 3063 5793
rect 3036 5623 3043 5643
rect 3016 5616 3043 5623
rect 3016 5367 3023 5616
rect 2936 4696 2963 4703
rect 2956 4587 2963 4696
rect 3016 4667 3023 5333
rect 3056 4936 3063 5353
rect 3076 5187 3083 5413
rect 3096 5176 3103 5213
rect 3116 4987 3123 5653
rect 3216 5643 3223 5836
rect 3196 5636 3223 5643
rect 3076 4956 3083 4973
rect 3116 4956 3123 4973
rect 3096 4927 3103 4943
rect 3056 4687 3063 4793
rect 3136 4767 3143 5073
rect 3116 4696 3143 4703
rect 3096 4667 3103 4683
rect 3136 4607 3143 4696
rect 3156 4607 3163 5633
rect 3176 4887 3183 5603
rect 3256 5587 3263 6056
rect 3256 5487 3263 5513
rect 3216 5436 3223 5453
rect 3256 5436 3263 5473
rect 3276 5427 3283 6033
rect 3296 5587 3303 6336
rect 3316 6327 3323 6336
rect 3336 5763 3343 6213
rect 3356 5887 3363 6413
rect 3376 6123 3383 6573
rect 3396 6227 3403 6813
rect 3416 6587 3423 7056
rect 3436 6807 3443 6913
rect 3456 6807 3463 7293
rect 3476 7227 3483 7273
rect 3476 6907 3483 7113
rect 3456 6607 3463 6633
rect 3476 6503 3483 6793
rect 3516 6667 3523 7213
rect 3576 7076 3583 7653
rect 3596 7543 3603 7573
rect 3676 7556 3703 7563
rect 3596 7536 3623 7543
rect 3616 7367 3623 7473
rect 3636 7267 3643 7473
rect 3576 6876 3583 7033
rect 3556 6663 3563 6863
rect 3596 6856 3603 6893
rect 3616 6823 3623 7153
rect 3636 6887 3643 7173
rect 3656 7167 3663 7513
rect 3696 7427 3703 7556
rect 3796 7427 3803 7776
rect 3836 7627 3843 7803
rect 3816 7547 3823 7563
rect 3856 7556 3863 7893
rect 3876 7627 3883 7913
rect 3896 7543 3903 7973
rect 3936 7847 3943 7893
rect 3956 7843 3963 7993
rect 3996 7863 4003 8316
rect 4016 8087 4023 8333
rect 4036 8027 4043 8473
rect 4056 8227 4063 8493
rect 4076 8467 4083 8523
rect 4076 8307 4083 8353
rect 4116 8336 4123 8536
rect 4156 8347 4163 8793
rect 4176 8647 4183 8933
rect 4196 8796 4203 8853
rect 4256 8803 4263 8983
rect 4276 8976 4303 8983
rect 4256 8796 4283 8803
rect 4216 8727 4223 8783
rect 4276 8503 4283 8796
rect 4216 8467 4223 8503
rect 4256 8496 4283 8503
rect 4236 8476 4253 8483
rect 4247 8336 4253 8343
rect 4196 8327 4203 8333
rect 4156 8316 4183 8323
rect 4096 8087 4103 8303
rect 4176 8227 4183 8316
rect 4216 8307 4223 8333
rect 4016 7987 4023 8013
rect 4056 7927 4063 8023
rect 4076 7887 4083 8033
rect 3996 7856 4023 7863
rect 3956 7836 3983 7843
rect 4016 7836 4023 7856
rect 3996 7807 4003 7823
rect 3736 7387 3743 7393
rect 3676 7167 3683 7373
rect 3716 7227 3723 7333
rect 3696 7067 3703 7133
rect 3596 6816 3623 6823
rect 3556 6656 3583 6663
rect 3456 6496 3483 6503
rect 3416 6167 3423 6453
rect 3456 6427 3463 6496
rect 3496 6487 3503 6583
rect 3556 6563 3563 6593
rect 3476 6463 3483 6473
rect 3516 6463 3523 6563
rect 3476 6456 3523 6463
rect 3536 6556 3563 6563
rect 3516 6403 3523 6433
rect 3436 6396 3463 6403
rect 3496 6396 3523 6403
rect 3436 6367 3443 6396
rect 3376 6116 3403 6123
rect 3436 6116 3443 6153
rect 3376 5767 3383 6073
rect 3396 5967 3403 6116
rect 3476 6103 3483 6353
rect 3416 6067 3423 6103
rect 3456 6096 3483 6103
rect 3396 5927 3403 5953
rect 3456 5947 3463 6096
rect 3516 5987 3523 6396
rect 3536 6367 3543 6556
rect 3556 6427 3563 6473
rect 3576 6447 3583 6656
rect 3496 5916 3503 5973
rect 3556 5907 3563 6333
rect 3576 6067 3583 6103
rect 3456 5896 3483 5903
rect 3316 5756 3343 5763
rect 3176 4696 3183 4713
rect 3196 4707 3203 5373
rect 3216 5047 3223 5353
rect 3236 5267 3243 5413
rect 3296 5187 3303 5393
rect 3316 5347 3323 5756
rect 3336 5656 3343 5733
rect 3396 5663 3403 5893
rect 3376 5656 3403 5663
rect 3396 5507 3403 5656
rect 3456 5647 3463 5896
rect 3516 5827 3523 5873
rect 3516 5656 3523 5813
rect 3556 5656 3563 5813
rect 3576 5807 3583 5993
rect 3596 5867 3603 6816
rect 3616 6387 3623 6433
rect 3636 6407 3643 6873
rect 3656 6827 3663 7053
rect 3656 6727 3663 6773
rect 3676 6596 3683 6713
rect 3696 6587 3703 6653
rect 3716 6607 3723 7193
rect 3756 7107 3763 7343
rect 3796 7207 3803 7353
rect 3796 7083 3803 7153
rect 3836 7127 3843 7543
rect 3876 7536 3903 7543
rect 3796 7076 3823 7083
rect 3816 6903 3823 7076
rect 3836 6907 3843 7073
rect 3796 6896 3823 6903
rect 3736 6876 3763 6883
rect 3736 6747 3743 6876
rect 3836 6867 3843 6893
rect 3756 6587 3763 6613
rect 3656 6547 3663 6563
rect 3656 6467 3663 6493
rect 3636 6307 3643 6363
rect 3676 6347 3683 6363
rect 3676 6307 3683 6333
rect 3696 6267 3703 6473
rect 3616 5807 3623 5973
rect 3656 5936 3663 5953
rect 3696 5883 3703 6193
rect 3716 5887 3723 6493
rect 3676 5876 3703 5883
rect 3336 5416 3363 5423
rect 3356 5287 3363 5416
rect 3436 5327 3443 5433
rect 3596 5387 3603 5573
rect 3276 5107 3283 5163
rect 3356 5083 3363 5173
rect 3436 5147 3443 5293
rect 3476 5167 3483 5173
rect 3447 5136 3463 5143
rect 3496 5127 3503 5143
rect 3336 5076 3363 5083
rect 3216 4947 3223 5033
rect 3236 4956 3243 4973
rect 3296 4936 3323 4943
rect 3316 4787 3323 4936
rect 3336 4727 3343 5076
rect 3416 4983 3423 5093
rect 3416 4976 3443 4983
rect 3416 4847 3423 4976
rect 3516 4867 3523 5153
rect 2936 4483 2943 4533
rect 2956 4496 2963 4513
rect 2916 4476 2943 4483
rect 2916 4443 2923 4476
rect 2996 4447 3003 4513
rect 2916 4436 2943 4443
rect 2896 4316 2913 4323
rect 2896 3976 2903 4316
rect 2936 4107 2943 4436
rect 2976 4163 2983 4393
rect 3056 4267 3063 4593
rect 3116 4496 3123 4533
rect 3156 4476 3163 4513
rect 3136 4447 3143 4463
rect 3236 4263 3243 4653
rect 3216 4256 3243 4263
rect 3216 4247 3223 4256
rect 3016 4196 3023 4233
rect 3056 4187 3063 4203
rect 3036 4163 3043 4183
rect 2976 4156 3003 4163
rect 2776 3716 2803 3723
rect 2736 3527 2743 3573
rect 2756 3503 2763 3593
rect 2736 3496 2763 3503
rect 2496 3243 2503 3333
rect 2476 3236 2503 3243
rect 2476 3107 2483 3236
rect 2596 3036 2603 3073
rect 2636 3056 2643 3113
rect 2656 3087 2663 3203
rect 2616 2967 2623 3023
rect 2676 2807 2683 3353
rect 2636 2776 2663 2783
rect 2476 2627 2483 2743
rect 2516 2736 2543 2743
rect 2496 2556 2503 2693
rect 2536 2647 2543 2736
rect 2636 2727 2643 2776
rect 2676 2747 2683 2763
rect 2636 2576 2643 2633
rect 2516 2467 2523 2543
rect 2496 2227 2503 2263
rect 2536 2256 2563 2263
rect 2436 2076 2463 2083
rect 2456 2007 2463 2076
rect 2476 2067 2483 2083
rect 2376 1807 2383 1933
rect 2396 1816 2403 1953
rect 2416 1667 2423 1973
rect 2396 1587 2403 1613
rect 2416 1596 2423 1633
rect 2456 1596 2463 1993
rect 2536 1687 2543 2213
rect 2556 2187 2563 2256
rect 2576 2247 2583 2553
rect 2696 2527 2703 2773
rect 2556 2076 2563 2113
rect 2696 2027 2703 2243
rect 2336 1116 2343 1253
rect 2176 916 2203 923
rect 2176 807 2183 916
rect 2276 867 2283 1103
rect 2316 847 2323 1103
rect 2336 836 2343 853
rect 2216 707 2223 803
rect 2356 787 2363 803
rect 2176 636 2203 643
rect 2216 636 2223 673
rect 1836 616 1863 623
rect 1756 356 1763 553
rect 1816 387 1823 593
rect 1636 156 1643 173
rect 1736 147 1743 213
rect 1047 116 1063 123
rect 296 -24 303 13
rect 996 -24 1003 13
rect 1776 -17 1783 323
rect 1756 -24 1783 -17
rect 1796 -17 1803 173
rect 1876 127 1883 373
rect 1956 187 1963 633
rect 2136 407 2143 613
rect 2136 363 2143 393
rect 2136 356 2163 363
rect 1976 207 1983 323
rect 1916 176 1943 183
rect 1796 -24 1823 -17
rect 1916 -24 1923 176
rect 1996 -24 2003 173
rect 2076 147 2083 213
rect 2136 156 2143 193
rect 2156 136 2163 293
rect 2116 -24 2123 13
rect 2196 -17 2203 636
rect 2256 27 2263 693
rect 2376 367 2383 653
rect 2416 623 2423 1373
rect 2436 867 2443 1373
rect 2436 847 2443 853
rect 2436 627 2443 833
rect 2456 827 2463 1333
rect 2476 1307 2483 1653
rect 2576 1316 2583 1373
rect 2496 1267 2503 1313
rect 2516 1147 2523 1303
rect 2616 1267 2623 1673
rect 2716 1627 2723 2573
rect 2736 2507 2743 3073
rect 2756 2067 2763 3496
rect 2796 3347 2803 3716
rect 2976 3667 2983 3683
rect 2996 3627 3003 4156
rect 3016 4156 3043 4163
rect 3016 4016 3023 4156
rect 3156 3947 3163 4233
rect 3216 4196 3223 4233
rect 3196 4147 3203 4183
rect 3276 4183 3283 4593
rect 3336 4547 3343 4643
rect 3476 4496 3483 4513
rect 3296 4456 3323 4463
rect 3256 4176 3283 4183
rect 3176 3863 3183 4133
rect 3216 3947 3223 4153
rect 3156 3856 3183 3863
rect 2836 3503 2843 3573
rect 2816 3496 2843 3503
rect 2776 2887 2783 3243
rect 2816 3087 2823 3093
rect 2816 3056 2823 3073
rect 2736 1787 2743 1803
rect 2776 1627 2783 2793
rect 2796 2767 2803 3023
rect 2836 2756 2843 3033
rect 2856 2907 2863 3333
rect 2876 2787 2883 3613
rect 2896 3127 2903 3293
rect 2836 2536 2843 2553
rect 2876 2523 2883 2673
rect 2856 2516 2883 2523
rect 2796 2087 2803 2493
rect 2916 2327 2923 2453
rect 2856 2276 2883 2283
rect 2916 2276 2923 2313
rect 2876 2167 2883 2276
rect 2936 2227 2943 3613
rect 2956 3516 2963 3553
rect 2976 3487 2983 3503
rect 3036 3307 3043 3553
rect 3056 3287 3063 3633
rect 2976 3127 2983 3243
rect 3056 3223 3063 3273
rect 2996 3187 3003 3223
rect 3036 3216 3063 3223
rect 2956 2927 2963 3023
rect 2956 2747 2963 2873
rect 2836 2076 2863 2083
rect 2636 1596 2643 1613
rect 2636 1296 2643 1353
rect 2476 1083 2483 1133
rect 2556 1096 2583 1103
rect 2476 1076 2503 1083
rect 2576 1007 2583 1096
rect 2476 847 2483 853
rect 2576 836 2583 853
rect 2396 616 2423 623
rect 2416 387 2423 616
rect 2476 587 2483 833
rect 2556 767 2563 803
rect 2636 687 2643 1253
rect 2516 587 2523 623
rect 2556 607 2563 613
rect 2436 356 2443 413
rect 2416 307 2423 343
rect 2456 327 2463 343
rect 2276 176 2303 183
rect 2276 27 2283 176
rect 2336 147 2343 213
rect 2496 156 2503 173
rect 2516 136 2523 333
rect 2556 267 2563 473
rect 2596 356 2603 413
rect 2656 407 2663 1153
rect 2576 327 2583 343
rect 2636 327 2643 363
rect 2176 -24 2203 -17
rect 2316 -24 2323 13
rect 2596 -24 2603 213
rect 2616 136 2623 253
rect 2676 227 2683 1593
rect 2696 1307 2703 1413
rect 2716 1167 2723 1303
rect 2756 1267 2763 1303
rect 2776 1103 2783 1583
rect 2756 1096 2783 1103
rect 2716 147 2723 1053
rect 2776 867 2783 1073
rect 2836 667 2843 1613
rect 2776 636 2783 653
rect 2816 636 2843 643
rect 2796 607 2803 623
rect 2796 387 2803 593
rect 2836 567 2843 636
rect 2756 363 2763 373
rect 2756 356 2783 363
rect 2796 267 2803 343
rect 2836 247 2843 343
rect 2856 247 2863 2076
rect 2916 2056 2943 2063
rect 2876 1787 2883 2053
rect 2896 1967 2903 2043
rect 2916 1927 2923 2056
rect 2896 1127 2903 1853
rect 2916 1627 2923 1793
rect 2936 1787 2943 1913
rect 2956 1827 2963 2313
rect 2976 2267 2983 3073
rect 2996 2847 3003 3013
rect 3056 3007 3063 3216
rect 3076 3027 3083 3833
rect 3116 3736 3143 3743
rect 3116 3687 3123 3736
rect 3116 3267 3123 3673
rect 3156 3516 3163 3856
rect 3176 3727 3183 3833
rect 3196 3547 3203 3933
rect 3236 3747 3243 3813
rect 3256 3667 3263 4176
rect 3296 3827 3303 4213
rect 3316 4007 3323 4456
rect 3356 3987 3363 4193
rect 3376 4187 3383 4253
rect 3456 4216 3483 4223
rect 3476 4207 3483 4216
rect 3436 4187 3443 4203
rect 3276 3587 3283 3723
rect 3176 3307 3183 3373
rect 3116 3207 3123 3233
rect 3136 3223 3143 3253
rect 3176 3236 3183 3293
rect 3236 3227 3243 3533
rect 3276 3507 3283 3573
rect 3136 3216 3163 3223
rect 3136 3016 3143 3113
rect 3336 3107 3343 3653
rect 3356 3267 3363 3913
rect 3376 3767 3383 4173
rect 3396 3667 3403 4133
rect 3416 3907 3423 4153
rect 3496 4147 3503 4693
rect 3536 4683 3543 5313
rect 3556 5167 3563 5313
rect 3596 5147 3603 5213
rect 3616 4956 3623 5793
rect 3636 5416 3643 5433
rect 3656 5407 3663 5633
rect 3636 5127 3643 5373
rect 3676 5327 3683 5876
rect 3736 5667 3743 6393
rect 3756 6103 3763 6453
rect 3776 6267 3783 6813
rect 3796 6403 3803 6713
rect 3816 6707 3823 6863
rect 3856 6827 3863 7413
rect 3876 7047 3883 7413
rect 3916 7356 3923 7753
rect 3956 7387 3963 7753
rect 3976 7607 3983 7793
rect 3996 7627 4003 7793
rect 4036 7556 4043 7773
rect 4076 7767 4083 7873
rect 4076 7556 4083 7613
rect 3976 7407 3983 7453
rect 3896 7023 3903 7253
rect 3936 7207 3943 7343
rect 3996 7283 4003 7373
rect 4016 7327 4023 7543
rect 4096 7487 4103 7553
rect 4116 7447 4123 7953
rect 3996 7276 4023 7283
rect 3996 7076 4003 7173
rect 3876 7016 3903 7023
rect 3876 6927 3883 7016
rect 3916 6883 3923 7053
rect 3936 7027 3943 7063
rect 3956 7036 3983 7043
rect 3956 7003 3963 7036
rect 3936 6996 3963 7003
rect 3936 6927 3943 6996
rect 4016 6887 4023 7276
rect 4036 7207 4043 7373
rect 4056 7323 4063 7433
rect 4136 7423 4143 8193
rect 4196 8007 4203 8033
rect 4156 7927 4163 7953
rect 4216 7847 4223 8253
rect 4236 8087 4243 8313
rect 4276 8143 4283 8496
rect 4316 8327 4323 8533
rect 4276 8136 4303 8143
rect 4236 8056 4243 8073
rect 4276 8056 4283 8113
rect 4176 7543 4183 7833
rect 4236 7767 4243 7803
rect 4256 7787 4263 8043
rect 4296 7867 4303 8136
rect 4236 7556 4243 7573
rect 4176 7536 4203 7543
rect 4176 7447 4183 7513
rect 4196 7487 4203 7536
rect 4296 7527 4303 7543
rect 4116 7416 4143 7423
rect 4116 7387 4123 7416
rect 4096 7336 4103 7353
rect 4136 7323 4143 7373
rect 4256 7356 4263 7513
rect 4296 7356 4303 7473
rect 4316 7387 4323 8073
rect 4336 7807 4343 8793
rect 4356 8776 4363 9113
rect 4536 9027 4543 9263
rect 4416 9003 4423 9013
rect 4416 8996 4443 9003
rect 4376 8567 4383 8993
rect 4436 8867 4443 8996
rect 4456 8963 4463 8983
rect 4456 8956 4483 8963
rect 4476 8816 4483 8956
rect 4496 8887 4503 8983
rect 4576 8967 4583 9673
rect 4596 9607 4603 9736
rect 4996 9727 5003 9933
rect 4616 8996 4623 9353
rect 4636 9327 4643 9513
rect 4676 9507 4683 9513
rect 4676 9463 4683 9493
rect 4716 9476 4723 9593
rect 4936 9496 4943 9513
rect 4676 9456 4703 9463
rect 4636 9247 4643 9313
rect 4416 8516 4423 8633
rect 4396 8487 4403 8503
rect 4436 8487 4443 8503
rect 4456 8487 4463 8513
rect 4336 7487 4343 7773
rect 4356 7567 4363 8293
rect 4516 8276 4523 8373
rect 4396 7856 4403 8273
rect 4556 8247 4563 8593
rect 4416 8036 4423 8113
rect 4556 8107 4563 8233
rect 4456 8036 4483 8043
rect 4456 8003 4463 8036
rect 4436 7996 4463 8003
rect 4376 7787 4383 7823
rect 4456 7807 4463 7996
rect 4516 7967 4523 8053
rect 4576 8043 4583 8313
rect 4596 8287 4603 8613
rect 4616 8516 4623 8553
rect 4636 8527 4643 8983
rect 4656 8783 4663 9273
rect 4676 9243 4683 9293
rect 4676 9236 4703 9243
rect 4696 9023 4703 9236
rect 4836 9027 4843 9493
rect 5056 9467 5063 10173
rect 5076 9927 5083 9963
rect 5116 9776 5123 9853
rect 5176 9827 5183 10253
rect 5196 10236 5223 10243
rect 5196 10187 5203 10236
rect 5276 10147 5283 10293
rect 5356 9963 5363 10273
rect 5396 10107 5403 10293
rect 5436 10236 5443 10253
rect 5656 10223 5663 10333
rect 5676 10256 5683 10293
rect 5456 10107 5463 10223
rect 5556 10216 5583 10223
rect 5656 10216 5683 10223
rect 5576 10087 5583 10216
rect 5356 9956 5383 9963
rect 5456 9956 5483 9963
rect 5196 9907 5203 9923
rect 5356 9867 5363 9956
rect 5476 9927 5483 9956
rect 5296 9767 5303 9853
rect 5156 9756 5183 9763
rect 5096 9727 5103 9743
rect 5076 9487 5083 9713
rect 5116 9527 5123 9613
rect 5116 9463 5123 9513
rect 5096 9456 5123 9463
rect 4876 9276 4883 9313
rect 4916 9247 4923 9263
rect 4676 9016 4703 9023
rect 4676 8996 4683 9016
rect 4896 9016 4903 9053
rect 4656 8776 4683 8783
rect 4636 8476 4653 8483
rect 4676 8327 4683 8776
rect 4736 8707 4743 8783
rect 4776 8747 4783 8753
rect 4716 8507 4723 8593
rect 4736 8467 4743 8633
rect 4776 8516 4783 8733
rect 4856 8547 4863 8773
rect 4936 8763 4943 9413
rect 5036 9243 5043 9253
rect 5036 9236 5063 9243
rect 5116 9227 5123 9253
rect 5116 8983 5123 9013
rect 5096 8976 5123 8983
rect 5136 8967 5143 9733
rect 5176 9047 5183 9756
rect 5216 9507 5223 9743
rect 5296 9736 5303 9753
rect 5216 9263 5223 9473
rect 5256 9296 5263 9313
rect 5276 9307 5283 9443
rect 5216 9256 5243 9263
rect 5236 9023 5243 9256
rect 5236 9016 5263 9023
rect 4876 8627 4883 8763
rect 4916 8756 4943 8763
rect 4956 8747 4963 8793
rect 4816 8507 4823 8523
rect 4916 8507 4923 8533
rect 4976 8516 4983 8553
rect 5016 8516 5023 8853
rect 5036 8816 5043 8893
rect 5056 8747 5063 8783
rect 4796 8483 4803 8503
rect 4816 8487 4823 8493
rect 4767 8476 4803 8483
rect 4796 8296 4803 8453
rect 4876 8447 4883 8473
rect 4896 8447 4903 8493
rect 4736 8283 4743 8293
rect 4676 8247 4683 8283
rect 4716 8276 4743 8283
rect 4556 8036 4583 8043
rect 4596 7807 4603 8093
rect 4756 8067 4763 8283
rect 4896 8147 4903 8413
rect 4916 8336 4923 8453
rect 4956 8427 4963 8503
rect 4996 8467 5003 8503
rect 5056 8467 5063 8613
rect 5056 8307 5063 8453
rect 4647 7856 4653 7863
rect 4376 7527 4383 7613
rect 4396 7587 4403 7793
rect 4056 7316 4083 7323
rect 4116 7316 4143 7323
rect 4116 7227 4123 7316
rect 4176 7267 4183 7333
rect 3916 6876 3943 6883
rect 3916 6727 3923 6876
rect 4016 6827 4023 6873
rect 3876 6596 3883 6633
rect 3816 6447 3823 6583
rect 3916 6567 3923 6613
rect 3796 6396 3823 6403
rect 3856 6396 3863 6473
rect 3836 6307 3843 6383
rect 3756 6096 3783 6103
rect 3756 5987 3763 6073
rect 3776 5847 3783 6053
rect 3796 5943 3803 6073
rect 3816 6067 3823 6103
rect 3856 5947 3863 6093
rect 3796 5936 3823 5943
rect 3796 5727 3803 5936
rect 3696 5187 3703 5633
rect 3716 5507 3723 5623
rect 3736 5447 3743 5603
rect 3756 5567 3763 5623
rect 3756 5427 3763 5553
rect 3656 5047 3663 5153
rect 3636 4976 3643 5033
rect 3516 4676 3543 4683
rect 3596 4676 3623 4683
rect 3616 4647 3623 4676
rect 3576 4456 3603 4463
rect 3576 4327 3583 4456
rect 3616 4227 3623 4573
rect 3656 4507 3663 4713
rect 3656 4443 3663 4493
rect 3636 4436 3663 4443
rect 3496 3963 3503 4013
rect 3436 3927 3443 3963
rect 3476 3956 3503 3963
rect 3416 3563 3423 3893
rect 3396 3556 3423 3563
rect 3396 3536 3403 3556
rect 3376 3467 3383 3503
rect 3367 3256 3383 3263
rect 3416 3256 3423 3413
rect 3356 3067 3363 3133
rect 3156 2807 3163 3003
rect 3296 2987 3303 3013
rect 3356 2996 3363 3053
rect 3376 3016 3403 3023
rect 3176 2783 3183 2913
rect 3156 2776 3183 2783
rect 3076 2756 3103 2763
rect 3056 2727 3063 2743
rect 3096 2607 3103 2756
rect 3136 2743 3143 2773
rect 3116 2736 3143 2743
rect 3156 2723 3163 2776
rect 3216 2747 3223 2763
rect 3136 2716 3163 2723
rect 2996 2523 3003 2573
rect 3036 2536 3043 2593
rect 2996 2516 3023 2523
rect 3016 2247 3023 2293
rect 3036 2287 3043 2393
rect 3056 2307 3063 2523
rect 3136 2507 3143 2716
rect 3156 2556 3183 2563
rect 3136 2303 3143 2493
rect 3116 2296 3143 2303
rect 3116 2267 3123 2296
rect 3036 1967 3043 2253
rect 3056 2187 3063 2263
rect 3096 2207 3103 2263
rect 3156 2227 3163 2556
rect 3236 2387 3243 2793
rect 3316 2787 3323 2993
rect 3396 2887 3403 3016
rect 3456 2947 3463 3873
rect 3556 3803 3563 4213
rect 3636 4187 3643 4203
rect 3576 3996 3603 4003
rect 3636 3996 3643 4033
rect 3576 3927 3583 3996
rect 3676 3987 3683 5113
rect 3756 5107 3763 5393
rect 3696 4027 3703 4213
rect 3716 4027 3723 4913
rect 3736 4807 3743 4973
rect 3776 4967 3783 5653
rect 3796 5127 3803 5253
rect 3816 5127 3823 5893
rect 3836 5827 3843 5903
rect 3856 5623 3863 5933
rect 3876 5887 3883 6213
rect 3896 5647 3903 6153
rect 3916 5907 3923 6533
rect 3936 6227 3943 6693
rect 3956 6283 3963 6593
rect 3976 6547 3983 6813
rect 4036 6747 4043 7033
rect 4056 6887 4063 7093
rect 4116 6863 4123 7083
rect 4136 7047 4143 7103
rect 4096 6856 4123 6863
rect 4016 6487 4023 6653
rect 4076 6623 4083 6693
rect 4096 6667 4103 6856
rect 4176 6836 4183 6893
rect 4196 6856 4203 7133
rect 4216 7047 4223 7353
rect 4276 7323 4283 7343
rect 4256 7316 4283 7323
rect 4116 6667 4123 6813
rect 4076 6616 4103 6623
rect 4096 6596 4103 6616
rect 4036 6563 4043 6583
rect 4076 6567 4083 6583
rect 4136 6583 4143 6733
rect 4127 6576 4143 6583
rect 4036 6556 4063 6563
rect 4036 6347 4043 6383
rect 3956 6276 3983 6283
rect 3936 5687 3943 5833
rect 3856 5616 3883 5623
rect 3856 5307 3863 5616
rect 3956 5507 3963 6253
rect 3976 6067 3983 6276
rect 3996 6167 4003 6253
rect 4036 6083 4043 6293
rect 4056 6187 4063 6556
rect 4016 6076 4043 6083
rect 4007 6056 4013 6063
rect 3916 5467 3923 5493
rect 3876 5436 3883 5453
rect 3836 5143 3843 5193
rect 3876 5156 3883 5193
rect 3916 5167 3923 5293
rect 3836 5136 3863 5143
rect 3796 4936 3803 5093
rect 3776 4903 3783 4923
rect 3776 4896 3803 4903
rect 3756 4676 3763 4713
rect 3616 3947 3623 3983
rect 3696 3983 3703 4013
rect 3696 3976 3723 3983
rect 3556 3796 3583 3803
rect 3496 3523 3503 3743
rect 3536 3736 3543 3753
rect 3516 3707 3523 3723
rect 3556 3587 3563 3673
rect 3496 3516 3523 3523
rect 3516 3496 3523 3516
rect 3496 3427 3503 3483
rect 3556 3467 3563 3573
rect 3576 3487 3583 3796
rect 3596 3467 3603 3483
rect 3536 3236 3563 3243
rect 3536 3207 3543 3236
rect 3476 3056 3503 3063
rect 3476 3007 3483 3056
rect 3336 2527 3343 2723
rect 3356 2576 3363 2593
rect 3476 2547 3483 2793
rect 3496 2567 3503 2953
rect 3516 2807 3523 2993
rect 3516 2707 3523 2763
rect 3536 2627 3543 3053
rect 3576 2987 3583 3153
rect 3556 2587 3563 2773
rect 3056 2096 3063 2153
rect 3196 2003 3203 2373
rect 3296 2067 3303 2243
rect 3436 2096 3443 2313
rect 3316 2027 3323 2063
rect 3196 1996 3223 2003
rect 3096 1816 3103 1953
rect 3216 1903 3223 1996
rect 3216 1896 3243 1903
rect 2996 1796 3023 1803
rect 3056 1796 3063 1813
rect 2976 1587 2983 1783
rect 3016 1767 3023 1796
rect 2956 1316 2983 1323
rect 2956 1096 2963 1316
rect 2996 1267 3003 1283
rect 2896 883 2903 1083
rect 2876 876 2903 883
rect 2876 627 2883 876
rect 2956 856 2983 863
rect 2976 847 2983 856
rect 2996 667 3003 1173
rect 3016 727 3023 1613
rect 3036 1547 3043 1783
rect 3076 1596 3083 1713
rect 3116 1596 3123 1833
rect 3136 1787 3143 1803
rect 3156 1596 3183 1603
rect 3036 907 3043 1093
rect 3036 867 3043 893
rect 3056 827 3063 1453
rect 3096 1387 3103 1583
rect 3136 1467 3143 1583
rect 3116 1307 3123 1353
rect 3176 1347 3183 1596
rect 3156 1316 3163 1333
rect 3196 1316 3203 1373
rect 3236 1367 3243 1896
rect 3256 1567 3263 1763
rect 3316 1547 3323 1583
rect 3136 1287 3143 1303
rect 3076 1116 3143 1123
rect 3076 1083 3083 1116
rect 3136 1107 3143 1116
rect 3156 1096 3163 1113
rect 3076 1076 3103 1083
rect 3176 1067 3183 1273
rect 3116 856 3123 1053
rect 3196 1027 3203 1073
rect 3236 1067 3243 1333
rect 3256 1307 3263 1353
rect 3276 1127 3283 1313
rect 3396 1287 3403 1853
rect 3416 1803 3423 2073
rect 3436 1867 3443 2013
rect 3416 1796 3443 1803
rect 3456 1623 3463 1793
rect 3496 1747 3503 2553
rect 3516 2247 3523 2573
rect 3556 2276 3563 2293
rect 3516 2007 3523 2083
rect 3496 1707 3503 1733
rect 3436 1616 3463 1623
rect 3376 1267 3383 1283
rect 3416 1263 3423 1613
rect 3436 1267 3443 1616
rect 3476 1287 3483 1303
rect 3396 1256 3423 1263
rect 3256 1096 3283 1103
rect 3256 1007 3263 1096
rect 3356 1083 3363 1153
rect 3336 1076 3363 1083
rect 3156 807 3163 863
rect 3176 827 3183 843
rect 3256 827 3263 993
rect 3316 856 3323 1053
rect 2936 603 2943 633
rect 3016 616 3023 673
rect 2936 596 2963 603
rect 2956 427 2963 573
rect 2896 27 2903 233
rect 2916 136 2923 393
rect 2936 367 2943 393
rect 2956 356 2963 413
rect 2996 356 3003 373
rect 3036 343 3043 773
rect 3136 636 3143 793
rect 3176 687 3183 813
rect 3156 636 3183 643
rect 3156 443 3163 636
rect 3016 336 3043 343
rect 3136 436 3163 443
rect 2976 287 2983 323
rect 3016 143 3023 313
rect 3136 207 3143 436
rect 3156 356 3163 413
rect 3196 387 3203 493
rect 3196 356 3203 373
rect 3236 367 3243 793
rect 3316 636 3343 643
rect 3216 327 3223 343
rect 2996 136 3023 143
rect 3116 176 3143 183
rect 2816 -24 2823 13
rect 3116 -24 3123 176
rect 3156 127 3163 143
rect 3176 -17 3183 193
rect 3316 167 3323 636
rect 3356 587 3363 863
rect 3376 827 3383 843
rect 3376 807 3383 813
rect 3396 783 3403 1256
rect 3476 1136 3483 1173
rect 3376 776 3403 783
rect 3376 636 3383 776
rect 3336 376 3363 383
rect 3336 263 3343 376
rect 3416 347 3423 1073
rect 3436 367 3443 593
rect 3336 256 3363 263
rect 3356 147 3363 256
rect 3336 116 3353 123
rect 3156 -24 3183 -17
rect 3336 -24 3343 93
rect 3436 -17 3443 173
rect 3456 27 3463 873
rect 3496 847 3503 893
rect 3516 887 3523 1303
rect 3556 1187 3563 2233
rect 3576 887 3583 2973
rect 3596 2756 3603 2773
rect 3596 2287 3603 2693
rect 3596 2087 3603 2273
rect 3616 1627 3623 3913
rect 3636 3496 3643 3833
rect 3736 3747 3743 4593
rect 3636 2227 3643 3253
rect 3656 3087 3663 3713
rect 3756 3707 3763 4473
rect 3796 4447 3803 4896
rect 3836 4607 3843 4893
rect 3856 4667 3863 4953
rect 3816 4476 3823 4493
rect 3796 4187 3803 4223
rect 3836 4216 3843 4473
rect 3876 4387 3883 5113
rect 3896 4967 3903 5123
rect 3936 4907 3943 5173
rect 3956 4923 3963 5153
rect 3976 4967 3983 5853
rect 4016 5827 4023 5883
rect 3996 5187 4003 5773
rect 4016 5607 4023 5733
rect 3956 4916 3983 4923
rect 4016 4907 4023 4923
rect 3936 4696 3963 4703
rect 3956 4687 3963 4696
rect 4036 4627 4043 5933
rect 4056 5867 4063 5993
rect 4056 5587 4063 5673
rect 4076 5647 4083 6473
rect 4116 6467 4123 6553
rect 4096 6327 4103 6433
rect 4096 6067 4103 6133
rect 4116 5683 4123 6053
rect 4136 5883 4143 6533
rect 4156 6207 4163 6813
rect 4216 6567 4223 6853
rect 4236 6827 4243 7253
rect 4256 6767 4263 7316
rect 4316 7307 4323 7343
rect 4236 6607 4243 6733
rect 4276 6596 4283 7273
rect 4356 7247 4363 7373
rect 4296 7063 4303 7113
rect 4316 7096 4323 7173
rect 4356 7107 4363 7193
rect 4296 7056 4323 7063
rect 4296 6727 4303 7033
rect 4316 6827 4323 7056
rect 4336 6876 4343 6913
rect 4176 6187 4183 6363
rect 4176 6147 4183 6173
rect 4216 6116 4223 6213
rect 4156 6067 4163 6103
rect 4236 6067 4243 6573
rect 4256 6567 4263 6583
rect 4256 6367 4263 6473
rect 4256 5967 4263 6113
rect 4276 6103 4283 6453
rect 4296 6127 4303 6553
rect 4316 6327 4323 6373
rect 4316 6107 4323 6133
rect 4276 6096 4303 6103
rect 4176 5936 4183 5953
rect 4196 5916 4223 5923
rect 4136 5876 4163 5883
rect 4107 5676 4123 5683
rect 4096 5656 4103 5673
rect 4156 5567 4163 5876
rect 4216 5807 4223 5916
rect 4236 5767 4243 5913
rect 4076 5436 4083 5453
rect 4096 5436 4123 5443
rect 4096 5287 4103 5436
rect 4076 5156 4083 5173
rect 4056 5107 4063 5143
rect 3936 4467 3943 4493
rect 3996 4456 4003 4493
rect 4016 4436 4033 4443
rect 3816 4127 3823 4203
rect 3976 4163 3983 4433
rect 4036 4163 4043 4313
rect 4056 4167 4063 4993
rect 4096 4747 4103 5273
rect 4116 4907 4123 5273
rect 4136 5147 4143 5393
rect 4196 5307 4203 5673
rect 4236 5407 4243 5753
rect 4276 5636 4283 5873
rect 4296 5603 4303 6096
rect 4336 6087 4343 6833
rect 4376 6823 4383 7333
rect 4396 7307 4403 7573
rect 4416 7543 4423 7693
rect 4496 7556 4503 7593
rect 4416 7536 4443 7543
rect 4416 7167 4423 7513
rect 4436 7267 4443 7513
rect 4496 7376 4503 7413
rect 4536 7356 4543 7573
rect 4456 7343 4463 7353
rect 4576 7347 4583 7673
rect 4596 7587 4603 7793
rect 4596 7543 4603 7573
rect 4596 7536 4623 7543
rect 4656 7467 4663 7543
rect 4636 7367 4643 7453
rect 4676 7443 4683 7933
rect 4716 7867 4723 7933
rect 4736 7856 4743 7913
rect 4756 7883 4763 8053
rect 4936 8047 4943 8153
rect 4756 7876 4783 7883
rect 4716 7836 4723 7853
rect 4756 7836 4763 7853
rect 4756 7547 4763 7693
rect 4776 7627 4783 7876
rect 4816 7787 4823 7833
rect 4796 7543 4803 7773
rect 4836 7687 4843 8033
rect 4856 7576 4863 7893
rect 4876 7836 4883 7913
rect 4956 7867 4963 8073
rect 4896 7807 4903 7823
rect 4936 7816 4963 7823
rect 4796 7536 4823 7543
rect 4656 7436 4683 7443
rect 4456 7336 4483 7343
rect 4396 6876 4403 6993
rect 4416 6927 4423 7153
rect 4356 6816 4383 6823
rect 4356 6567 4363 6816
rect 4376 6467 4383 6713
rect 4356 6267 4363 6453
rect 4396 6376 4403 6833
rect 4416 6387 4423 6893
rect 4436 6583 4443 6973
rect 4476 6867 4483 7336
rect 4516 7147 4523 7213
rect 4536 7096 4543 7313
rect 4576 7103 4583 7253
rect 4556 7096 4583 7103
rect 4496 6907 4503 6993
rect 4516 6843 4523 7063
rect 4536 6876 4543 6993
rect 4556 6903 4563 7096
rect 4596 7063 4603 7153
rect 4576 7056 4603 7063
rect 4556 6896 4583 6903
rect 4516 6836 4543 6843
rect 4436 6576 4463 6583
rect 4456 6367 4463 6413
rect 4376 6307 4383 6363
rect 4356 6167 4363 6253
rect 4356 6107 4363 6123
rect 4396 6116 4403 6153
rect 4316 5827 4323 6073
rect 4376 6067 4383 6103
rect 4416 6087 4423 6103
rect 4276 5596 4303 5603
rect 4256 5547 4263 5593
rect 4276 5456 4283 5596
rect 4256 5416 4283 5423
rect 4276 5163 4283 5416
rect 4296 5167 4303 5473
rect 4256 5156 4283 5163
rect 4136 4987 4143 5133
rect 4136 4956 4143 4973
rect 4176 4956 4183 4993
rect 4196 4936 4203 5113
rect 4136 4827 4143 4913
rect 4156 4687 4163 4933
rect 4216 4927 4223 4953
rect 4236 4907 4243 5143
rect 4076 4367 4083 4633
rect 4116 4627 4123 4663
rect 4096 4427 4103 4613
rect 4136 4467 4143 4653
rect 4176 4647 4183 4893
rect 4196 4667 4203 4693
rect 4156 4456 4163 4493
rect 4176 4476 4183 4533
rect 4216 4476 4223 4713
rect 4236 4507 4243 4853
rect 4256 4623 4263 4953
rect 4276 4947 4283 4993
rect 4296 4867 4303 5153
rect 4276 4636 4303 4643
rect 4256 4616 4283 4623
rect 4136 4447 4143 4453
rect 3976 4156 4003 4163
rect 4016 4156 4043 4163
rect 3776 3983 3783 3993
rect 3776 3976 3803 3983
rect 3696 3587 3703 3703
rect 3736 3696 3753 3703
rect 3776 3607 3783 3976
rect 3836 3927 3843 4113
rect 3976 4016 3983 4033
rect 3896 3627 3903 3683
rect 3936 3496 3943 3593
rect 3756 3256 3763 3273
rect 3776 3247 3783 3293
rect 3856 3256 3863 3273
rect 3896 3256 3923 3263
rect 3856 3036 3863 3053
rect 3896 3036 3903 3093
rect 3696 3016 3703 3033
rect 3716 2987 3723 3003
rect 3736 2776 3763 2783
rect 3736 2547 3743 2776
rect 3716 2527 3723 2543
rect 3776 2327 3783 2533
rect 3636 2107 3643 2193
rect 3636 2076 3643 2093
rect 3716 1827 3723 2263
rect 3656 1623 3663 1813
rect 3696 1647 3703 1763
rect 3656 1616 3683 1623
rect 3656 1567 3663 1583
rect 3676 1343 3683 1616
rect 3736 1583 3743 2313
rect 3756 2047 3763 2083
rect 3756 1787 3763 2033
rect 3756 1667 3763 1773
rect 3716 1576 3743 1583
rect 3656 1336 3683 1343
rect 3596 787 3603 1313
rect 3656 1147 3663 1336
rect 3736 1316 3743 1373
rect 3676 1167 3683 1303
rect 3776 1303 3783 1313
rect 3796 1307 3803 2213
rect 3816 2067 3823 2333
rect 3836 2107 3843 3033
rect 3876 2787 3883 2893
rect 3916 2607 3923 3256
rect 3936 3207 3943 3233
rect 3956 3187 3963 3733
rect 3976 3227 3983 3973
rect 3996 3147 4003 4156
rect 4176 4163 4183 4183
rect 4156 4156 4183 4163
rect 4096 3976 4123 3983
rect 4116 3847 4123 3976
rect 4156 3887 4163 4156
rect 4016 3427 4023 3503
rect 4036 3307 4043 3723
rect 4056 3667 4063 3703
rect 4096 3527 4103 3703
rect 4096 3287 4103 3513
rect 3976 2756 3983 2993
rect 4016 2967 4023 3213
rect 4076 3183 4083 3203
rect 4056 3176 4083 3183
rect 4036 3016 4043 3053
rect 4056 2996 4063 3176
rect 4096 3047 4103 3213
rect 3936 2687 3943 2743
rect 4116 2667 4123 3733
rect 4176 3543 4183 4013
rect 4216 3963 4223 4433
rect 4236 4347 4243 4473
rect 4236 3976 4243 4313
rect 4207 3956 4223 3963
rect 4256 3747 4263 4413
rect 4276 4147 4283 4616
rect 4296 4487 4303 4636
rect 4316 4487 4323 5413
rect 4336 4907 4343 6053
rect 4436 6027 4443 6173
rect 4356 5847 4363 5883
rect 4396 5876 4403 5913
rect 4456 5907 4463 6313
rect 4356 4936 4363 5753
rect 4476 5727 4483 6553
rect 4436 5656 4443 5673
rect 4376 5423 4383 5593
rect 4496 5427 4503 6583
rect 4516 6567 4523 6603
rect 4536 6543 4543 6836
rect 4556 6767 4563 6863
rect 4616 6847 4623 7193
rect 4656 7067 4663 7436
rect 4756 7356 4763 7533
rect 4696 7327 4703 7343
rect 4636 6867 4643 6873
rect 4556 6567 4563 6633
rect 4516 6536 4543 6543
rect 4516 6027 4523 6536
rect 4576 6487 4583 6733
rect 4596 6487 4603 6833
rect 4567 6416 4573 6423
rect 4616 6423 4623 6593
rect 4636 6583 4643 6853
rect 4676 6827 4683 7093
rect 4716 7076 4723 7273
rect 4776 7167 4783 7353
rect 4796 7127 4803 7473
rect 4756 7067 4763 7083
rect 4736 7047 4743 7063
rect 4696 6847 4703 6873
rect 4716 6847 4723 7013
rect 4756 6907 4763 6993
rect 4776 6907 4783 7073
rect 4796 6927 4803 7093
rect 4816 7027 4823 7536
rect 4836 7047 4843 7563
rect 4816 6876 4823 6913
rect 4856 6903 4863 7513
rect 4876 7323 4883 7513
rect 4896 7347 4903 7773
rect 4916 7527 4923 7793
rect 4936 7487 4943 7673
rect 4956 7607 4963 7816
rect 4976 7807 4983 8193
rect 4996 7567 5003 8093
rect 5076 8087 5083 8553
rect 5096 8487 5103 8513
rect 5096 8296 5103 8313
rect 5116 8247 5123 8533
rect 5096 8063 5103 8213
rect 5136 8207 5143 8893
rect 5156 8547 5163 9013
rect 5216 8927 5223 8963
rect 5176 8816 5203 8823
rect 5176 8707 5183 8816
rect 5236 8783 5243 8873
rect 5256 8807 5263 9016
rect 5216 8776 5243 8783
rect 5256 8567 5263 8793
rect 5156 8503 5163 8533
rect 5156 8496 5183 8503
rect 5187 8476 5203 8483
rect 5156 8107 5163 8413
rect 5176 8407 5183 8433
rect 5016 8056 5043 8063
rect 5076 8056 5103 8063
rect 5016 7927 5023 8056
rect 5056 8027 5063 8043
rect 5016 7807 5023 7833
rect 4916 7356 4923 7393
rect 4996 7356 5003 7433
rect 5036 7387 5043 7833
rect 5076 7787 5083 7853
rect 5116 7816 5123 7833
rect 5156 7816 5163 7853
rect 4936 7327 4943 7343
rect 4876 7316 4903 7323
rect 4836 6896 4863 6903
rect 4836 6847 4843 6896
rect 4676 6747 4683 6813
rect 4676 6607 4683 6653
rect 4716 6596 4723 6613
rect 4636 6576 4663 6583
rect 4636 6523 4643 6553
rect 4656 6547 4663 6576
rect 4736 6567 4743 6583
rect 4636 6516 4663 6523
rect 4616 6416 4643 6423
rect 4536 6387 4543 6413
rect 4596 6396 4603 6413
rect 4636 6396 4643 6416
rect 4656 6407 4663 6516
rect 4736 6487 4743 6513
rect 4576 6227 4583 6383
rect 4536 6167 4543 6193
rect 4576 6027 4583 6103
rect 4516 5847 4523 5913
rect 4376 5416 4403 5423
rect 4396 5047 4403 5143
rect 4416 5087 4423 5123
rect 4456 5087 4463 5153
rect 4496 5147 4503 5393
rect 4516 5007 4523 5173
rect 4536 5127 4543 5953
rect 4556 5896 4563 6013
rect 4576 5916 4583 5933
rect 4616 5927 4623 6113
rect 4596 5887 4603 5903
rect 4656 5767 4663 6373
rect 4676 6227 4683 6473
rect 4716 6307 4723 6393
rect 4736 6327 4743 6393
rect 4756 6387 4763 6833
rect 4776 6587 4783 6713
rect 4796 6627 4803 6833
rect 4816 6627 4823 6793
rect 4796 6567 4803 6593
rect 4816 6396 4823 6613
rect 4836 6563 4843 6813
rect 4856 6583 4863 6873
rect 4876 6707 4883 6913
rect 4896 6827 4903 7316
rect 4936 7107 4943 7173
rect 4956 7087 4963 7213
rect 4976 7187 4983 7333
rect 5056 7227 5063 7593
rect 4976 7083 4983 7093
rect 4976 7076 5003 7083
rect 4956 7027 4963 7043
rect 4996 6927 5003 7076
rect 4896 6647 4903 6793
rect 4996 6783 5003 6863
rect 4996 6776 5023 6783
rect 4936 6587 4943 6773
rect 4856 6576 4883 6583
rect 4916 6567 4923 6583
rect 4836 6556 4863 6563
rect 4696 5687 4703 6213
rect 4716 5823 4723 6153
rect 4736 6107 4743 6123
rect 4776 6116 4783 6153
rect 4816 6127 4823 6153
rect 4776 5916 4783 5993
rect 4796 5947 4803 6103
rect 4836 5963 4843 6513
rect 4856 5967 4863 6556
rect 4876 6207 4883 6553
rect 4896 6547 4903 6563
rect 4956 6427 4963 6773
rect 4976 6607 4983 6633
rect 4996 6607 5003 6693
rect 4996 6487 5003 6533
rect 4816 5956 4843 5963
rect 4816 5927 4823 5956
rect 4716 5816 4743 5823
rect 4616 5647 4623 5663
rect 4656 5656 4683 5663
rect 4596 5627 4603 5643
rect 4636 5567 4643 5643
rect 4676 5607 4683 5656
rect 4556 5143 4563 5453
rect 4616 5436 4623 5493
rect 4696 5436 4703 5513
rect 4616 5156 4623 5173
rect 4556 5136 4583 5143
rect 4536 5047 4543 5053
rect 4536 4976 4543 5033
rect 4556 5027 4563 5053
rect 4576 5007 4583 5136
rect 4656 5143 4663 5153
rect 4636 5136 4663 5143
rect 4676 5087 4683 5253
rect 4696 5147 4703 5313
rect 4716 5147 4723 5793
rect 4416 4956 4423 4973
rect 4336 4587 4343 4733
rect 4296 4456 4323 4463
rect 4316 4327 4323 4456
rect 4396 4167 4403 4893
rect 4436 4696 4443 4753
rect 4416 4496 4423 4613
rect 4276 3716 4303 3723
rect 4276 3683 4283 3716
rect 4256 3676 4283 3683
rect 4336 3627 4343 4133
rect 4416 4107 4423 4453
rect 4496 4203 4503 4373
rect 4496 4196 4523 4203
rect 4556 4196 4563 4253
rect 4576 4223 4583 4973
rect 4696 4863 4703 5013
rect 4716 4956 4723 5133
rect 4736 5027 4743 5816
rect 4756 5427 4763 5633
rect 4756 5407 4763 5413
rect 4776 5387 4783 5653
rect 4796 5647 4803 5893
rect 4816 5636 4823 5653
rect 4836 5647 4843 5933
rect 4876 5907 4883 6113
rect 4896 6107 4903 6373
rect 4916 6143 4923 6413
rect 4936 6267 4943 6413
rect 5016 6323 5023 6776
rect 5036 6487 5043 6913
rect 5056 6847 5063 6873
rect 5076 6827 5083 6873
rect 5096 6827 5103 7803
rect 5136 7796 5143 7813
rect 5136 7527 5143 7593
rect 5156 7587 5163 7673
rect 5176 7607 5183 8303
rect 5196 8127 5203 8476
rect 5196 8023 5203 8113
rect 5276 8107 5283 8913
rect 5236 8036 5243 8053
rect 5196 8016 5223 8023
rect 5256 8007 5263 8023
rect 5276 7807 5283 7913
rect 5296 7907 5303 9053
rect 5316 8787 5323 9813
rect 5336 9207 5343 9273
rect 5316 8296 5323 8313
rect 5336 8127 5343 9153
rect 5356 8907 5363 9313
rect 5396 8996 5403 9473
rect 5496 9467 5503 9913
rect 5576 9736 5603 9743
rect 5576 9607 5583 9736
rect 5656 9723 5663 10193
rect 5676 9887 5683 10216
rect 5836 10207 5843 10683
rect 5856 10387 5863 10693
rect 5896 10567 5903 10696
rect 5916 10407 5923 10433
rect 5936 10427 5943 10433
rect 5936 10383 5943 10413
rect 5916 10376 5943 10383
rect 5856 10287 5863 10373
rect 5856 10216 5863 10273
rect 5756 9976 5763 10133
rect 5796 9976 5823 9983
rect 5636 9716 5663 9723
rect 5476 9276 5483 9293
rect 5456 9187 5463 9233
rect 5516 9207 5523 9273
rect 5436 9047 5443 9173
rect 5456 9027 5463 9133
rect 5456 9003 5463 9013
rect 5436 8996 5463 9003
rect 5536 9003 5543 9273
rect 5616 9016 5623 9173
rect 5536 8996 5563 9003
rect 5576 8996 5603 9003
rect 5476 8547 5483 8793
rect 5436 8536 5463 8543
rect 5456 8447 5463 8536
rect 5516 8527 5523 8773
rect 5496 8336 5503 8413
rect 5536 8387 5543 8893
rect 5576 8887 5583 8996
rect 5596 8816 5603 8953
rect 5556 8536 5563 8553
rect 5596 8536 5623 8543
rect 5616 8323 5623 8536
rect 5596 8316 5623 8323
rect 5316 7836 5323 7953
rect 5356 7927 5363 8193
rect 5516 8167 5523 8293
rect 5376 7987 5383 8053
rect 5356 7836 5363 7913
rect 5376 7847 5383 7893
rect 5176 7547 5183 7563
rect 5156 7487 5163 7533
rect 5116 7347 5123 7473
rect 5216 7467 5223 7753
rect 5156 7356 5163 7453
rect 5136 7336 5143 7353
rect 5176 7323 5183 7343
rect 5156 7316 5183 7323
rect 5156 7247 5163 7316
rect 5116 7047 5123 7083
rect 5156 7076 5163 7233
rect 5176 6927 5183 7063
rect 5196 7027 5203 7133
rect 5216 6927 5223 7353
rect 5136 6876 5143 6893
rect 5176 6876 5183 6893
rect 5236 6883 5243 7713
rect 5336 7583 5343 7823
rect 5396 7587 5403 8093
rect 5416 7807 5423 8093
rect 5456 8027 5463 8043
rect 5476 7967 5483 8063
rect 5516 7907 5523 8133
rect 5576 8087 5583 8193
rect 5596 8063 5603 8316
rect 5616 8087 5623 8233
rect 5636 8083 5643 9533
rect 5676 9467 5683 9873
rect 5656 9407 5663 9463
rect 5656 9187 5663 9243
rect 5696 9227 5703 9243
rect 5716 8927 5723 9493
rect 5736 9287 5743 9953
rect 5776 9943 5783 9963
rect 5776 9936 5803 9943
rect 5796 9736 5803 9936
rect 5816 9827 5823 9976
rect 5816 9756 5823 9793
rect 5856 9756 5863 9913
rect 5916 9907 5923 10376
rect 5936 10107 5943 10173
rect 5936 9943 5943 10093
rect 6016 9943 6023 10473
rect 6036 10216 6043 10553
rect 6196 10447 6203 11393
rect 6256 11027 6263 11416
rect 6396 11383 6403 11693
rect 6436 11623 6443 11693
rect 6476 11676 6503 11683
rect 6496 11667 6503 11676
rect 6616 11656 6623 11693
rect 6427 11616 6443 11623
rect 6556 11547 6563 11633
rect 6676 11627 6683 11643
rect 6396 11376 6423 11383
rect 6296 11196 6303 11373
rect 6476 11363 6483 11513
rect 6436 11247 6443 11363
rect 6456 11356 6483 11363
rect 6456 11176 6463 11356
rect 6416 11147 6423 11163
rect 6296 10927 6303 11033
rect 6356 10943 6363 11133
rect 6336 10936 6363 10943
rect 6256 10847 6263 10903
rect 6276 10763 6283 10923
rect 6356 10827 6363 10936
rect 6276 10756 6303 10763
rect 6276 10703 6283 10733
rect 6256 10696 6283 10703
rect 6116 10327 6123 10423
rect 6156 10307 6163 10423
rect 6176 10407 6183 10443
rect 6296 10427 6303 10756
rect 6376 10467 6383 10673
rect 6416 10667 6423 10703
rect 6376 10436 6383 10453
rect 6316 10367 6323 10423
rect 6136 9963 6143 10273
rect 6036 9956 6063 9963
rect 6116 9956 6143 9963
rect 5936 9936 5963 9943
rect 5996 9936 6023 9943
rect 5956 9867 5963 9936
rect 5776 9227 5783 9593
rect 5836 9523 5843 9743
rect 5836 9516 5863 9523
rect 5856 9276 5863 9516
rect 5876 9507 5883 9793
rect 5896 9567 5903 9773
rect 5916 9523 5923 9733
rect 5896 9516 5923 9523
rect 5896 9487 5903 9516
rect 5756 8967 5763 8983
rect 5716 8796 5723 8913
rect 5776 8776 5783 8913
rect 5816 8827 5823 9003
rect 5656 8276 5683 8283
rect 5636 8076 5663 8083
rect 5656 8067 5663 8076
rect 5576 8056 5603 8063
rect 5616 8056 5643 8063
rect 5336 7576 5363 7583
rect 5356 7556 5363 7576
rect 5416 7556 5423 7793
rect 5256 7067 5263 7533
rect 5396 7387 5403 7543
rect 5296 7356 5323 7363
rect 5356 7356 5363 7373
rect 5276 7307 5283 7353
rect 5276 7147 5283 7293
rect 5276 6907 5283 7093
rect 5296 7047 5303 7356
rect 5336 7327 5343 7343
rect 5316 7067 5323 7083
rect 5356 7076 5363 7273
rect 5416 7227 5423 7333
rect 5396 7047 5403 7173
rect 5216 6876 5243 6883
rect 5116 6787 5123 6853
rect 5156 6843 5163 6863
rect 5156 6836 5183 6843
rect 5136 6823 5143 6833
rect 5136 6816 5163 6823
rect 5056 6603 5063 6713
rect 5056 6596 5083 6603
rect 5116 6596 5123 6693
rect 5156 6627 5163 6816
rect 5176 6807 5183 6836
rect 5156 6583 5163 6613
rect 5096 6567 5103 6583
rect 5136 6576 5163 6583
rect 5016 6316 5043 6323
rect 4916 6136 4943 6143
rect 4936 6127 4943 6136
rect 4976 6116 4983 6313
rect 5036 6267 5043 6316
rect 5016 6147 5023 6253
rect 4916 5987 4923 6103
rect 4956 6027 4963 6103
rect 4916 5967 4923 5973
rect 4796 5467 4803 5533
rect 4836 5463 4843 5633
rect 4816 5456 4843 5463
rect 4816 5443 4823 5456
rect 4796 5436 4823 5443
rect 4756 4983 4763 5193
rect 4796 5167 4803 5436
rect 4736 4976 4763 4983
rect 4756 4956 4783 4963
rect 4696 4856 4723 4863
rect 4636 4676 4643 4853
rect 4676 4623 4683 4753
rect 4656 4616 4683 4623
rect 4596 4456 4623 4463
rect 4616 4223 4623 4456
rect 4636 4247 4643 4493
rect 4576 4216 4603 4223
rect 4616 4216 4643 4223
rect 4536 4127 4543 4183
rect 4596 4183 4603 4216
rect 4636 4207 4643 4216
rect 4587 4176 4603 4183
rect 4356 3723 4363 3973
rect 4356 3716 4383 3723
rect 4376 3607 4383 3716
rect 4176 3536 4203 3543
rect 4396 3536 4403 3813
rect 4556 3667 4563 3683
rect 4196 3516 4203 3536
rect 4216 3496 4243 3503
rect 4236 3267 4243 3496
rect 4416 3247 4423 3593
rect 4516 3516 4523 3613
rect 4576 3547 4583 4093
rect 4616 3827 4623 3983
rect 4556 3516 4583 3523
rect 4396 3187 4403 3203
rect 4176 2807 4183 3053
rect 4256 2907 4263 3023
rect 4176 2747 4183 2793
rect 4296 2787 4303 2953
rect 4196 2776 4223 2783
rect 4196 2747 4203 2776
rect 3856 2267 3863 2573
rect 3916 2247 3923 2293
rect 3876 2127 3883 2173
rect 3876 2076 3883 2113
rect 3836 1796 3863 1803
rect 3836 1427 3843 1796
rect 3896 1763 3903 1773
rect 3876 1756 3903 1763
rect 3756 1296 3783 1303
rect 3876 1267 3883 1303
rect 3616 1027 3623 1073
rect 3616 867 3623 1013
rect 3696 883 3703 1083
rect 3676 876 3703 883
rect 3476 307 3483 573
rect 3556 527 3563 623
rect 3676 447 3683 876
rect 3716 863 3723 1133
rect 3696 856 3723 863
rect 3547 376 3563 383
rect 3596 376 3623 383
rect 3536 187 3543 373
rect 3616 343 3623 376
rect 3596 336 3623 343
rect 3536 127 3543 173
rect 3596 147 3603 336
rect 3616 176 3643 183
rect 3436 -24 3463 -17
rect 3496 -24 3503 13
rect 3616 -24 3623 176
rect 3696 -17 3703 856
rect 3756 843 3763 1113
rect 3896 1103 3903 1633
rect 3936 1627 3943 2653
rect 3956 2303 3963 2593
rect 4136 2576 4143 2713
rect 4316 2567 4323 2693
rect 4376 2587 4383 3133
rect 4396 3036 4403 3053
rect 4416 2987 4423 3023
rect 4456 3016 4483 3023
rect 4476 2967 4483 3016
rect 4496 3007 4503 3033
rect 4496 2943 4503 2993
rect 4476 2936 4503 2943
rect 4476 2756 4483 2936
rect 4516 2927 4523 3243
rect 4456 2727 4463 2743
rect 3996 2536 4023 2543
rect 4316 2536 4323 2553
rect 3976 2507 3983 2523
rect 3996 2407 4003 2536
rect 3956 2296 3983 2303
rect 3956 2207 3963 2273
rect 3916 1147 3923 1303
rect 3876 1096 3903 1103
rect 3916 1096 3923 1113
rect 3816 907 3823 1093
rect 3736 836 3763 843
rect 3816 836 3823 893
rect 3716 667 3723 823
rect 3736 803 3743 836
rect 3856 827 3863 1083
rect 3936 1047 3943 1613
rect 3736 796 3763 803
rect 3716 636 3723 653
rect 3756 647 3763 796
rect 3876 687 3883 873
rect 3876 636 3883 673
rect 3896 667 3903 853
rect 3916 636 3923 813
rect 3956 547 3963 1133
rect 3976 887 3983 2296
rect 4036 2283 4043 2493
rect 4036 2276 4063 2283
rect 4096 2276 4103 2293
rect 4276 2227 4283 2263
rect 4296 2247 4303 2283
rect 4416 2263 4423 2693
rect 4516 2623 4523 2753
rect 4556 2747 4563 3053
rect 4496 2616 4523 2623
rect 4496 2527 4503 2616
rect 4516 2576 4543 2583
rect 4516 2547 4523 2576
rect 4416 2256 4443 2263
rect 4476 2247 4483 2263
rect 4356 2076 4363 2213
rect 4396 2087 4403 2093
rect 4496 2087 4503 2283
rect 4516 2147 4523 2533
rect 4556 2527 4563 2543
rect 4536 2127 4543 2273
rect 3996 1796 4023 1803
rect 3996 1727 4003 1796
rect 4056 1763 4063 2033
rect 4296 1783 4303 2053
rect 4296 1776 4313 1783
rect 4036 1756 4063 1763
rect 3996 1596 4003 1693
rect 4176 1616 4183 1653
rect 4016 1596 4043 1603
rect 4016 1163 4023 1596
rect 4156 1327 4163 1613
rect 4336 1603 4343 1993
rect 4376 1783 4383 1933
rect 4356 1776 4383 1783
rect 4456 1776 4483 1783
rect 4456 1767 4463 1776
rect 4336 1596 4363 1603
rect 4396 1596 4403 1613
rect 4196 1347 4203 1583
rect 4456 1567 4463 1753
rect 4556 1667 4563 1773
rect 4556 1616 4563 1633
rect 4216 1336 4243 1343
rect 3996 1156 4023 1163
rect 3996 867 4003 1156
rect 4016 1136 4043 1143
rect 4016 1107 4023 1136
rect 4056 1116 4063 1213
rect 4116 1103 4123 1273
rect 4156 1127 4163 1313
rect 4216 1167 4223 1336
rect 4316 1323 4323 1553
rect 4456 1387 4463 1393
rect 4296 1316 4323 1323
rect 4396 1316 4423 1323
rect 4456 1316 4463 1373
rect 4536 1367 4543 1583
rect 4216 1136 4243 1143
rect 4096 1096 4123 1103
rect 3976 727 3983 803
rect 3716 376 3743 383
rect 3776 376 3803 383
rect 3716 187 3723 376
rect 3756 347 3763 363
rect 3796 227 3803 376
rect 3836 327 3843 353
rect 3856 347 3863 453
rect 3776 176 3803 183
rect 3776 27 3783 176
rect 3836 143 3843 213
rect 3816 136 3843 143
rect 3696 -24 3723 -17
rect 3816 -24 3823 13
rect 3876 -17 3883 533
rect 3956 356 3963 493
rect 3976 387 3983 653
rect 3996 347 4003 393
rect 4016 367 4023 873
rect 3976 327 3983 343
rect 3956 123 3963 173
rect 3996 136 4003 293
rect 3956 116 3983 123
rect 4036 -17 4043 853
rect 4156 836 4163 853
rect 4196 803 4203 1133
rect 4216 1067 4223 1136
rect 4176 796 4203 803
rect 4056 603 4063 793
rect 4096 616 4103 633
rect 4056 596 4083 603
rect 4116 596 4123 653
rect 4076 507 4083 596
rect 4096 367 4103 433
rect 4116 376 4123 453
rect 4176 407 4183 633
rect 4096 176 4123 183
rect 4096 27 4103 176
rect 4156 147 4163 383
rect 4196 363 4203 493
rect 4176 356 4203 363
rect 4216 287 4223 1033
rect 4256 887 4263 1093
rect 4256 827 4263 853
rect 4236 347 4243 713
rect 4276 683 4283 1153
rect 4276 676 4303 683
rect 4296 667 4303 676
rect 4296 636 4303 653
rect 4316 647 4323 843
rect 4396 503 4403 1316
rect 4476 1287 4483 1303
rect 4536 1047 4543 1133
rect 4476 856 4483 873
rect 4456 656 4463 673
rect 4436 607 4443 613
rect 4396 496 4423 503
rect 4416 427 4423 496
rect 4256 367 4263 393
rect 4276 363 4283 373
rect 4276 356 4303 363
rect 4276 156 4283 333
rect 4316 327 4323 383
rect 4356 376 4383 383
rect 4376 187 4383 376
rect 4396 347 4403 373
rect 4416 207 4423 413
rect 4496 383 4503 843
rect 4576 663 4583 3516
rect 4656 3147 4663 4616
rect 4696 4463 4703 4833
rect 4676 4456 4703 4463
rect 4676 3767 4683 4433
rect 4716 4267 4723 4856
rect 4776 4667 4783 4956
rect 4816 4727 4823 5133
rect 4836 4947 4843 5423
rect 4876 5416 4883 5453
rect 4836 4687 4843 4693
rect 4816 4647 4823 4663
rect 4736 4447 4743 4633
rect 4856 4463 4863 4653
rect 4836 4456 4863 4463
rect 4696 3987 4703 4193
rect 4716 3987 4723 4253
rect 4876 4207 4883 5373
rect 4896 5107 4903 5913
rect 4916 5447 4923 5953
rect 4936 5916 4943 5933
rect 4956 5887 4963 5903
rect 4996 5896 5003 6073
rect 5016 6067 5023 6113
rect 5036 6067 5043 6093
rect 5016 5767 5023 6013
rect 4916 4976 4923 5413
rect 4936 5287 4943 5753
rect 4996 5656 5023 5663
rect 4976 5623 4983 5643
rect 5016 5627 5023 5656
rect 4956 5616 4983 5623
rect 4956 5427 4963 5616
rect 5036 5487 5043 5893
rect 5056 5847 5063 6093
rect 5056 5607 5063 5733
rect 5076 5567 5083 6353
rect 5096 5987 5103 6473
rect 5116 6416 5123 6553
rect 5156 6387 5163 6553
rect 5176 6487 5183 6633
rect 5196 6407 5203 6713
rect 5216 6567 5223 6813
rect 5256 6727 5263 6893
rect 5276 6787 5283 6873
rect 5296 6627 5303 6873
rect 5316 6867 5323 6893
rect 5236 6427 5243 6593
rect 5256 6523 5263 6553
rect 5276 6547 5283 6553
rect 5296 6523 5303 6563
rect 5256 6516 5303 6523
rect 5336 6507 5343 7033
rect 5396 6747 5403 6893
rect 5356 6487 5363 6613
rect 5116 6376 5143 6383
rect 5116 6187 5123 6376
rect 5236 6367 5243 6393
rect 5116 6027 5123 6073
rect 5136 6047 5143 6253
rect 5236 6147 5243 6153
rect 5216 6116 5243 6123
rect 5196 6047 5203 6083
rect 5096 5707 5103 5973
rect 5136 5916 5143 5933
rect 4976 5387 4983 5433
rect 4956 5156 4963 5173
rect 4896 4163 4903 4633
rect 4916 4627 4923 4673
rect 4956 4667 4963 4773
rect 4976 4643 4983 4793
rect 4996 4727 5003 5433
rect 5036 5207 5043 5413
rect 5076 4987 5083 5453
rect 5096 5123 5103 5693
rect 5116 5687 5123 5913
rect 5196 5896 5203 5933
rect 5216 5863 5223 6013
rect 5196 5856 5223 5863
rect 5136 5636 5163 5643
rect 5136 5427 5143 5636
rect 5176 5587 5183 5603
rect 5196 5587 5203 5856
rect 5216 5647 5223 5693
rect 5236 5607 5243 6116
rect 5256 5647 5263 6413
rect 5276 6396 5283 6413
rect 5356 6396 5363 6473
rect 5336 6367 5343 6383
rect 5276 6047 5283 6353
rect 5276 5787 5283 6033
rect 5156 5267 5163 5513
rect 5176 5436 5203 5443
rect 5236 5436 5243 5473
rect 5256 5467 5263 5633
rect 5296 5487 5303 6133
rect 5316 6027 5323 6153
rect 5336 6047 5343 6333
rect 5376 6147 5383 6593
rect 5396 6307 5403 6473
rect 5396 6116 5403 6193
rect 5416 6187 5423 7213
rect 5436 6483 5443 7793
rect 5456 7187 5463 7533
rect 5456 7087 5463 7153
rect 5476 7067 5483 7893
rect 5536 7787 5543 7803
rect 5556 7703 5563 7873
rect 5576 7767 5583 8056
rect 5616 8047 5623 8056
rect 5616 8007 5623 8033
rect 5636 8016 5663 8023
rect 5596 7907 5603 7993
rect 5636 7987 5643 8016
rect 5676 8003 5683 8276
rect 5656 7996 5683 8003
rect 5596 7787 5603 7813
rect 5536 7696 5563 7703
rect 5536 7607 5543 7696
rect 5516 7307 5523 7573
rect 5536 7356 5543 7593
rect 5556 7576 5563 7673
rect 5596 7576 5603 7673
rect 5616 7627 5623 7913
rect 5636 7603 5643 7953
rect 5656 7627 5663 7996
rect 5676 7807 5683 7823
rect 5636 7596 5663 7603
rect 5576 7543 5583 7563
rect 5656 7547 5663 7596
rect 5576 7536 5603 7543
rect 5556 7247 5563 7343
rect 5596 7336 5603 7536
rect 5656 7467 5663 7513
rect 5616 7227 5623 7353
rect 5536 7076 5543 7213
rect 5456 6727 5463 6913
rect 5456 6596 5463 6613
rect 5476 6607 5483 6913
rect 5476 6547 5483 6563
rect 5456 6507 5463 6533
rect 5436 6476 5463 6483
rect 5436 6387 5443 6413
rect 5356 6027 5363 6093
rect 5416 6087 5423 6103
rect 5336 5916 5343 5993
rect 5376 5916 5383 5933
rect 5396 5847 5403 5913
rect 5376 5607 5383 5623
rect 5176 5403 5183 5436
rect 5176 5396 5203 5403
rect 5156 5156 5163 5193
rect 5196 5147 5203 5396
rect 5296 5367 5303 5453
rect 5316 5367 5323 5413
rect 5376 5403 5383 5593
rect 5396 5467 5403 5773
rect 5416 5527 5423 5993
rect 5436 5767 5443 6233
rect 5456 6087 5463 6476
rect 5476 5907 5483 6533
rect 5496 6396 5503 7053
rect 5516 6907 5523 7063
rect 5596 7043 5603 7113
rect 5556 7027 5563 7043
rect 5576 7036 5603 7043
rect 5556 6887 5563 7013
rect 5516 6427 5523 6773
rect 5536 6767 5543 6843
rect 5576 6836 5583 7036
rect 5616 6867 5623 7013
rect 5556 6627 5563 6813
rect 5616 6807 5623 6833
rect 5636 6807 5643 7453
rect 5676 7347 5683 7753
rect 5656 7227 5663 7333
rect 5696 7107 5703 7613
rect 5716 7563 5723 8713
rect 5816 8707 5823 8793
rect 5836 8747 5843 9263
rect 5876 9256 5883 9333
rect 5916 9307 5923 9473
rect 5936 8947 5943 9393
rect 5956 8947 5963 9813
rect 5976 9496 5983 9893
rect 6056 9787 6063 9956
rect 6296 9907 6303 9923
rect 6316 9883 6323 10293
rect 6336 10216 6343 10273
rect 6356 10267 6363 10423
rect 6396 10107 6403 10423
rect 6416 10307 6423 10653
rect 6436 10223 6443 10253
rect 6416 10216 6443 10223
rect 6456 9987 6463 10193
rect 6296 9876 6323 9883
rect 6076 9763 6083 9793
rect 6216 9767 6223 9853
rect 6056 9756 6083 9763
rect 6156 9756 6183 9763
rect 6016 9527 6023 9713
rect 6016 9496 6023 9513
rect 5996 9027 6003 9483
rect 6036 9427 6043 9743
rect 6156 9667 6163 9756
rect 6156 9547 6163 9653
rect 6016 9263 6023 9373
rect 6076 9276 6083 9313
rect 6016 9256 6043 9263
rect 6016 8996 6023 9053
rect 5976 8976 6003 8983
rect 5976 8927 5983 8976
rect 5996 8796 6003 8953
rect 6036 8847 6043 8983
rect 5756 8516 5783 8523
rect 5776 8507 5783 8516
rect 5736 8467 5743 8483
rect 5756 7687 5763 8433
rect 5796 8316 5803 8693
rect 5836 8447 5843 8733
rect 5896 8723 5903 8793
rect 5916 8776 5933 8783
rect 5916 8747 5923 8776
rect 5976 8747 5983 8783
rect 5896 8716 5923 8723
rect 5836 8316 5843 8353
rect 5776 8147 5783 8273
rect 5796 8047 5803 8273
rect 5816 8056 5823 8303
rect 5856 8296 5863 8313
rect 5876 8263 5883 8573
rect 5916 8516 5923 8716
rect 5956 8567 5963 8733
rect 5956 8516 5963 8553
rect 5936 8427 5943 8503
rect 5976 8407 5983 8503
rect 5876 8256 5903 8263
rect 5896 8043 5903 8256
rect 5876 8036 5903 8043
rect 5716 7556 5743 7563
rect 5776 7556 5783 8013
rect 5876 7947 5883 8036
rect 5916 7967 5923 8333
rect 5796 7583 5803 7933
rect 5936 7927 5943 8073
rect 5956 7987 5963 8373
rect 5976 7987 5983 8353
rect 5996 8296 6023 8303
rect 5996 8043 6003 8296
rect 6036 8227 6043 8813
rect 6056 8527 6063 8873
rect 6076 8607 6083 8973
rect 6076 8287 6083 8593
rect 6096 8483 6103 8773
rect 6116 8747 6123 9133
rect 6136 8983 6143 9173
rect 6156 9147 6163 9453
rect 6196 9427 6203 9463
rect 6176 9027 6183 9293
rect 6216 9276 6223 9433
rect 6236 9243 6243 9263
rect 6276 9256 6283 9293
rect 6236 9236 6263 9243
rect 6216 9087 6223 9213
rect 6136 8976 6163 8983
rect 6176 8947 6183 8963
rect 6196 8827 6203 8983
rect 6096 8476 6123 8483
rect 6116 8107 6123 8476
rect 5996 8036 6023 8043
rect 6036 8007 6043 8023
rect 5816 7816 5843 7823
rect 5796 7576 5823 7583
rect 5756 7447 5763 7543
rect 5816 7363 5823 7576
rect 5836 7507 5843 7816
rect 5856 7807 5863 7833
rect 5896 7547 5903 7573
rect 5796 7356 5823 7363
rect 5836 7167 5843 7353
rect 5756 7076 5763 7113
rect 5656 7047 5663 7073
rect 5796 7063 5803 7153
rect 5836 7107 5843 7133
rect 5856 7107 5863 7513
rect 5916 7376 5923 7693
rect 5976 7687 5983 7713
rect 5956 7663 5963 7673
rect 5956 7656 5983 7663
rect 5976 7587 5983 7656
rect 5936 7247 5943 7343
rect 5876 7107 5883 7173
rect 5536 6547 5543 6593
rect 5536 6396 5543 6433
rect 5516 6363 5523 6383
rect 5496 6356 5523 6363
rect 5456 5547 5463 5893
rect 5496 5883 5503 6356
rect 5576 6343 5583 6353
rect 5556 6336 5583 6343
rect 5516 6087 5523 6173
rect 5536 6116 5543 6213
rect 5556 6147 5563 6336
rect 5516 5927 5523 6053
rect 5576 5923 5583 6313
rect 5596 5967 5603 6583
rect 5636 6347 5643 6583
rect 5616 6107 5623 6193
rect 5556 5916 5583 5923
rect 5576 5907 5583 5916
rect 5476 5876 5503 5883
rect 5476 5727 5483 5876
rect 5496 5747 5503 5853
rect 5476 5647 5483 5713
rect 5476 5603 5483 5633
rect 5576 5627 5583 5753
rect 5536 5616 5563 5623
rect 5476 5596 5503 5603
rect 5456 5467 5463 5533
rect 5396 5436 5403 5453
rect 5476 5436 5483 5473
rect 5496 5427 5503 5596
rect 5416 5407 5423 5423
rect 5456 5407 5463 5413
rect 5376 5396 5403 5403
rect 5096 5116 5123 5123
rect 5116 4956 5123 5116
rect 5036 4867 5043 4953
rect 5136 4947 5143 5143
rect 5296 5143 5303 5213
rect 5316 5187 5323 5353
rect 5356 5247 5363 5333
rect 5376 5156 5383 5173
rect 5296 5136 5323 5143
rect 5096 4927 5103 4943
rect 4996 4643 5003 4683
rect 5056 4647 5063 4663
rect 4976 4636 5003 4643
rect 4876 4156 4903 4163
rect 4736 3536 4743 4133
rect 4976 4127 4983 4636
rect 4996 4476 5003 4613
rect 5036 4483 5043 4573
rect 5036 4476 5063 4483
rect 5016 4216 5043 4223
rect 4796 4016 4823 4023
rect 4816 3987 4823 4016
rect 4756 3727 4763 3833
rect 4816 3787 4823 3973
rect 4916 3847 4923 3983
rect 4596 3036 4623 3043
rect 4596 2787 4603 3036
rect 4616 2267 4623 2533
rect 4636 2267 4643 2573
rect 4656 2547 4663 2723
rect 4676 2347 4683 3493
rect 4696 3223 4703 3533
rect 4716 3387 4723 3503
rect 4836 3267 4843 3733
rect 4856 3716 4883 3723
rect 4696 3216 4723 3223
rect 4756 3107 4763 3223
rect 4856 3127 4863 3716
rect 4936 3687 4943 3993
rect 4976 3983 4983 4073
rect 4956 3976 4983 3983
rect 4996 3967 5003 4173
rect 5016 3747 5023 4216
rect 5036 3967 5043 4173
rect 5056 3867 5063 4476
rect 5076 3843 5083 4773
rect 5096 4187 5103 4853
rect 5156 4607 5163 4973
rect 5216 4827 5223 4953
rect 5156 4476 5163 4593
rect 5216 4456 5223 4493
rect 5136 4427 5143 4453
rect 5156 4207 5163 4313
rect 5176 4203 5183 4433
rect 5176 4196 5203 4203
rect 5236 4196 5243 5093
rect 5356 5087 5363 5123
rect 5296 4976 5303 5013
rect 5316 4847 5323 4943
rect 5396 4847 5403 5396
rect 5416 5347 5423 5393
rect 5416 4767 5423 5293
rect 5296 4667 5303 4693
rect 5256 4627 5263 4663
rect 5116 4016 5123 4153
rect 5216 4147 5223 4183
rect 5256 4127 5263 4183
rect 5256 4047 5263 4113
rect 5336 4027 5343 4713
rect 5416 4627 5423 4663
rect 5436 4603 5443 4953
rect 5456 4936 5463 5153
rect 5496 4987 5503 5413
rect 5516 5307 5523 5553
rect 5536 5187 5543 5593
rect 5496 4927 5503 4933
rect 5416 4596 5443 4603
rect 5356 4496 5363 4533
rect 5376 4427 5383 4463
rect 5376 4196 5383 4333
rect 5416 4196 5423 4596
rect 5536 4527 5543 4993
rect 5556 4663 5563 5616
rect 5576 4827 5583 5593
rect 5596 5167 5603 5913
rect 5616 5527 5623 6073
rect 5636 5463 5643 6273
rect 5656 6127 5663 6573
rect 5676 6563 5683 7053
rect 5696 6907 5703 7013
rect 5716 6896 5723 7053
rect 5736 6927 5743 7063
rect 5776 7056 5803 7063
rect 5756 6876 5763 6993
rect 5696 6827 5703 6863
rect 5696 6587 5703 6793
rect 5716 6643 5723 6853
rect 5736 6807 5743 6833
rect 5716 6636 5743 6643
rect 5676 6556 5703 6563
rect 5696 6363 5703 6556
rect 5716 6527 5723 6613
rect 5736 6376 5743 6636
rect 5756 6427 5763 6593
rect 5776 6487 5783 7033
rect 5796 7007 5803 7056
rect 5816 6603 5823 6913
rect 5836 6607 5843 7093
rect 5896 7076 5903 7093
rect 5936 7076 5943 7153
rect 5796 6596 5823 6603
rect 5696 6356 5723 6363
rect 5696 6123 5703 6293
rect 5716 6147 5723 6356
rect 5676 6116 5703 6123
rect 5736 6116 5743 6333
rect 5756 6127 5763 6153
rect 5776 6147 5783 6333
rect 5796 6167 5803 6596
rect 5816 6267 5823 6373
rect 5656 6087 5663 6093
rect 5656 5607 5663 6073
rect 5676 5867 5683 6116
rect 5676 5567 5683 5753
rect 5696 5547 5703 6093
rect 5716 5896 5723 6103
rect 5796 6067 5803 6133
rect 5796 5923 5803 6053
rect 5776 5916 5803 5923
rect 5756 5887 5763 5903
rect 5816 5887 5823 6253
rect 5736 5636 5743 5873
rect 5756 5647 5763 5773
rect 5776 5636 5783 5813
rect 5816 5627 5823 5733
rect 5756 5567 5763 5593
rect 5696 5487 5703 5533
rect 5616 5456 5643 5463
rect 5616 5436 5623 5456
rect 5676 5416 5683 5453
rect 5696 5367 5703 5413
rect 5716 5307 5723 5433
rect 5616 5143 5623 5293
rect 5656 5156 5663 5253
rect 5696 5187 5703 5193
rect 5696 5156 5703 5173
rect 5596 5136 5623 5143
rect 5596 4947 5603 5136
rect 5636 5107 5643 5143
rect 5616 4943 5623 5033
rect 5656 4976 5663 4993
rect 5696 4956 5723 4963
rect 5616 4936 5643 4943
rect 5616 4696 5623 4853
rect 5596 4667 5603 4683
rect 5556 4656 5583 4663
rect 5347 4016 5363 4023
rect 5156 3996 5183 4003
rect 5056 3836 5083 3843
rect 5016 3703 5023 3733
rect 5016 3696 5043 3703
rect 4896 3503 4903 3653
rect 4876 3496 4903 3503
rect 4896 3247 4903 3496
rect 4696 2567 4703 3053
rect 4756 3036 4783 3043
rect 4816 3036 4823 3073
rect 4716 2727 4723 3033
rect 4756 2987 4763 3036
rect 4756 2787 4763 2973
rect 4876 2887 4883 3243
rect 4896 3067 4903 3233
rect 4976 3203 4983 3513
rect 5056 3507 5063 3836
rect 5096 3767 5103 3983
rect 5136 3967 5143 3983
rect 5116 3723 5123 3953
rect 5116 3716 5143 3723
rect 5136 3523 5143 3716
rect 5176 3627 5183 3996
rect 5196 3667 5203 3723
rect 5167 3536 5183 3543
rect 5136 3516 5163 3523
rect 5196 3516 5203 3533
rect 5136 3487 5143 3493
rect 5216 3347 5223 4013
rect 5396 3983 5403 3993
rect 5336 3967 5343 3983
rect 5376 3976 5403 3983
rect 5436 3927 5443 4183
rect 5456 4167 5463 4513
rect 5556 4476 5563 4493
rect 5476 4007 5483 4473
rect 5576 4443 5583 4656
rect 5556 4436 5583 4443
rect 5516 4016 5523 4153
rect 5556 4143 5563 4436
rect 5556 4136 5583 4143
rect 5556 3996 5563 4013
rect 5576 3987 5583 4136
rect 5536 3747 5543 3773
rect 5256 3236 5263 3553
rect 5316 3503 5323 3613
rect 5376 3543 5383 3683
rect 5376 3536 5403 3543
rect 5396 3516 5403 3536
rect 5316 3496 5343 3503
rect 5496 3367 5503 3723
rect 5636 3647 5643 4013
rect 5636 3503 5643 3633
rect 5656 3567 5663 4813
rect 5716 4583 5723 4956
rect 5736 4907 5743 5453
rect 5736 4767 5743 4893
rect 5756 4827 5763 5513
rect 5776 5287 5783 5533
rect 5736 4696 5743 4753
rect 5776 4727 5783 5253
rect 5796 4967 5803 5513
rect 5816 5107 5823 5613
rect 5836 5467 5843 6563
rect 5856 5867 5863 7073
rect 5876 6867 5883 7073
rect 5896 6747 5903 7013
rect 5916 6907 5923 7043
rect 5976 6927 5983 7333
rect 5976 6876 5983 6913
rect 5956 6847 5963 6853
rect 5856 5787 5863 5833
rect 5876 5807 5883 6433
rect 5916 6416 5923 6533
rect 5896 6367 5903 6383
rect 5936 6367 5943 6813
rect 5996 6767 6003 7813
rect 6016 7547 6023 7973
rect 6076 7907 6083 7993
rect 6096 7907 6103 8053
rect 6096 7816 6123 7823
rect 6096 7687 6103 7816
rect 6136 7783 6143 8483
rect 6156 8263 6163 8473
rect 6176 8327 6183 8513
rect 6216 8487 6223 9073
rect 6236 8467 6243 8833
rect 6196 8316 6203 8333
rect 6236 8316 6243 8453
rect 6256 8367 6263 9236
rect 6296 8847 6303 9876
rect 6336 9756 6363 9763
rect 6336 9727 6343 9756
rect 6416 9736 6443 9743
rect 6316 9227 6323 9493
rect 6336 8783 6343 9713
rect 6436 9647 6443 9736
rect 6456 9707 6463 9753
rect 6476 9687 6483 11333
rect 6556 11147 6563 11533
rect 6576 11383 6583 11613
rect 6696 11587 6703 11633
rect 6716 11627 6723 11673
rect 6736 11627 6743 11713
rect 6756 11707 6763 11873
rect 6576 11376 6603 11383
rect 6656 11287 6663 11393
rect 6736 11027 6743 11373
rect 6756 11183 6763 11693
rect 6776 11387 6783 11553
rect 6796 11347 6803 11893
rect 6836 11863 6843 11913
rect 7516 11896 7543 11903
rect 6916 11876 6923 11893
rect 7136 11876 7143 11893
rect 6836 11856 6863 11863
rect 6896 11767 6903 11863
rect 6936 11847 6943 11863
rect 6836 11627 6843 11663
rect 6876 11656 6883 11673
rect 6896 11607 6903 11673
rect 6756 11176 6783 11183
rect 6676 10907 6683 10923
rect 6776 10907 6783 11176
rect 6836 11167 6843 11183
rect 6496 10847 6503 10883
rect 6776 10827 6783 10893
rect 6596 10727 6603 10813
rect 6576 10436 6603 10443
rect 6496 10187 6503 10433
rect 6516 10387 6523 10423
rect 6556 10407 6563 10423
rect 6516 10247 6523 10373
rect 6596 10227 6603 10436
rect 6576 10107 6583 10223
rect 6416 9503 6423 9573
rect 6396 9496 6423 9503
rect 6416 9467 6423 9496
rect 6436 9347 6443 9633
rect 6356 8947 6363 8973
rect 6376 8967 6383 9273
rect 6416 9023 6423 9313
rect 6456 9296 6463 9353
rect 6496 9267 6503 10073
rect 6556 9967 6563 10073
rect 6596 10023 6603 10213
rect 6576 10016 6603 10023
rect 6516 9447 6523 9893
rect 6536 9496 6543 9773
rect 6576 9756 6583 10016
rect 6616 10003 6623 10753
rect 6676 10696 6703 10703
rect 6596 9996 6623 10003
rect 6636 10003 6643 10453
rect 6656 10207 6663 10683
rect 6676 10567 6683 10696
rect 6716 10387 6723 10423
rect 6696 10236 6723 10243
rect 6716 10207 6723 10236
rect 6776 10227 6783 10443
rect 6796 10067 6803 11153
rect 6816 10736 6823 11093
rect 6856 10967 6863 11383
rect 6916 11023 6923 11353
rect 6936 11047 6943 11673
rect 7016 11663 7023 11873
rect 7156 11847 7163 11863
rect 6996 11656 7023 11663
rect 7056 11656 7063 11813
rect 7296 11787 7303 11863
rect 7336 11827 7343 11863
rect 7376 11847 7383 11863
rect 7376 11787 7383 11833
rect 7276 11696 7303 11703
rect 6996 11627 7003 11656
rect 6956 11367 6963 11393
rect 6996 11383 7003 11613
rect 7076 11487 7083 11643
rect 7116 11527 7123 11653
rect 6996 11376 7023 11383
rect 6916 11016 6943 11023
rect 6856 10867 6863 10953
rect 6896 10903 6903 10993
rect 6936 10916 6943 11016
rect 6976 10947 6983 11373
rect 7016 11196 7023 11213
rect 6996 11176 7003 11193
rect 7076 11187 7083 11413
rect 7136 11407 7143 11643
rect 6976 10916 7003 10923
rect 6896 10896 6923 10903
rect 6996 10883 7003 10916
rect 7016 10887 7023 10933
rect 7036 10907 7043 10973
rect 6956 10707 6963 10883
rect 6976 10876 7003 10883
rect 6976 10603 6983 10876
rect 6996 10696 7003 10813
rect 6976 10596 7003 10603
rect 6916 10423 6923 10433
rect 6996 10427 7003 10596
rect 6916 10416 6943 10423
rect 6976 10387 6983 10413
rect 7016 10407 7023 10873
rect 6896 10247 6903 10253
rect 6916 10236 6923 10293
rect 7036 10287 7043 10813
rect 6896 10216 6903 10233
rect 6636 9996 6663 10003
rect 6596 9963 6603 9996
rect 6596 9956 6623 9963
rect 6656 9956 6663 9996
rect 6636 9927 6643 9943
rect 6776 9756 6783 9773
rect 6576 9503 6583 9713
rect 6596 9667 6603 9743
rect 6636 9707 6643 9743
rect 6796 9727 6803 9743
rect 6576 9496 6603 9503
rect 6556 9427 6563 9483
rect 6596 9467 6603 9496
rect 6756 9447 6763 9463
rect 6776 9427 6783 9483
rect 6836 9447 6843 9473
rect 6616 9276 6623 9333
rect 6756 9276 6763 9313
rect 6796 9276 6803 9293
rect 6396 9016 6423 9023
rect 6396 8996 6403 9016
rect 6436 8983 6443 9013
rect 6416 8976 6443 8983
rect 6356 8827 6363 8853
rect 6356 8796 6363 8813
rect 6536 8807 6543 8893
rect 6407 8796 6423 8803
rect 6316 8776 6343 8783
rect 6316 8587 6323 8776
rect 6376 8647 6383 8773
rect 6416 8607 6423 8796
rect 6276 8483 6283 8553
rect 6276 8476 6303 8483
rect 6176 8296 6183 8313
rect 6256 8307 6263 8353
rect 6156 8256 6183 8263
rect 6156 8027 6163 8073
rect 6176 7827 6183 8256
rect 6116 7776 6143 7783
rect 6116 7663 6123 7776
rect 6096 7656 6123 7663
rect 6036 7463 6043 7653
rect 6016 7456 6043 7463
rect 6016 7127 6023 7456
rect 6016 6867 6023 6893
rect 5976 6596 5983 6753
rect 6016 6647 6023 6833
rect 6036 6583 6043 7373
rect 6056 7347 6063 7473
rect 6096 7467 6103 7656
rect 6156 7627 6163 7803
rect 6076 7356 6083 7453
rect 6116 7363 6123 7473
rect 6136 7447 6143 7543
rect 6196 7487 6203 8053
rect 6216 8007 6223 8023
rect 6216 7556 6223 7573
rect 6236 7427 6243 8003
rect 6256 7987 6263 8023
rect 6276 7523 6283 8133
rect 6336 8067 6343 8553
rect 6476 8516 6483 8793
rect 6516 8747 6523 8783
rect 6516 8507 6523 8523
rect 6456 8483 6463 8503
rect 6456 8476 6483 8483
rect 6356 8387 6363 8413
rect 6436 8316 6463 8323
rect 6416 8287 6423 8303
rect 6416 8147 6423 8273
rect 6456 8147 6463 8316
rect 6476 8187 6483 8476
rect 6496 8407 6503 8503
rect 6376 8047 6383 8133
rect 6456 8087 6463 8133
rect 6496 8067 6503 8313
rect 6296 7887 6303 7913
rect 6336 7836 6343 7853
rect 6316 7807 6323 7823
rect 6376 7787 6383 7833
rect 6396 7807 6403 8023
rect 6416 7887 6423 8013
rect 6436 8007 6443 8033
rect 6496 7816 6503 8053
rect 6516 7867 6523 8433
rect 6536 8327 6543 8333
rect 6556 8327 6563 8733
rect 6576 8567 6583 9193
rect 6736 9107 6743 9253
rect 6776 9167 6783 9263
rect 6836 9223 6843 9293
rect 6856 9267 6863 10053
rect 6876 9967 6883 10093
rect 7036 9963 7043 10273
rect 7056 10267 7063 11033
rect 7076 10747 7083 10913
rect 7096 10883 7103 11393
rect 7216 11383 7223 11413
rect 7276 11387 7283 11696
rect 7196 11376 7223 11383
rect 7156 11216 7183 11223
rect 7156 11167 7163 11216
rect 7316 11207 7323 11433
rect 7336 11416 7363 11423
rect 7336 11327 7343 11416
rect 7316 11163 7323 11193
rect 7356 11187 7363 11253
rect 7316 11156 7343 11163
rect 7376 11127 7383 11163
rect 7136 10916 7143 11053
rect 7396 10967 7403 11073
rect 7176 10916 7183 10953
rect 7216 10903 7223 10933
rect 7396 10916 7403 10953
rect 7096 10876 7123 10883
rect 7116 10727 7123 10876
rect 7156 10767 7163 10903
rect 7196 10896 7223 10903
rect 7236 10807 7243 10913
rect 7376 10887 7383 10903
rect 7416 10807 7423 10903
rect 7296 10736 7303 10753
rect 7076 10667 7083 10703
rect 7076 10487 7083 10653
rect 7076 10263 7083 10373
rect 7096 10287 7103 10693
rect 7116 10683 7123 10713
rect 7116 10676 7143 10683
rect 7136 10347 7143 10423
rect 7156 10267 7163 10733
rect 7276 10567 7283 10693
rect 7176 10416 7203 10423
rect 7076 10256 7103 10263
rect 7116 10236 7123 10253
rect 7156 10227 7163 10253
rect 7156 9987 7163 10213
rect 7036 9956 7063 9963
rect 6876 9487 6883 9733
rect 6956 9687 6963 9853
rect 6996 9776 7003 9793
rect 6976 9756 6983 9773
rect 7016 9756 7043 9763
rect 7036 9727 7043 9756
rect 7036 9647 7043 9713
rect 6976 9487 6983 9633
rect 6876 9367 6883 9473
rect 6996 9443 7003 9463
rect 6976 9436 7003 9443
rect 6976 9407 6983 9436
rect 6816 9216 6843 9223
rect 6636 9016 6643 9093
rect 6776 9027 6783 9153
rect 6816 9027 6823 9216
rect 6876 9187 6883 9353
rect 6936 9276 6963 9283
rect 6996 9276 7003 9293
rect 6936 9247 6943 9276
rect 6936 9227 6943 9233
rect 6676 8987 6683 9023
rect 6836 9016 6843 9113
rect 6856 8987 6863 9003
rect 6676 8796 6683 8953
rect 6636 8503 6643 8593
rect 6676 8516 6683 8633
rect 6636 8496 6663 8503
rect 6616 8327 6623 8373
rect 6736 8316 6743 8493
rect 6756 8447 6763 8833
rect 6776 8327 6783 8853
rect 6536 8027 6543 8293
rect 6556 8267 6563 8283
rect 6596 8247 6603 8283
rect 6536 7816 6543 8013
rect 6256 7516 6283 7523
rect 6096 7356 6123 7363
rect 6136 7356 6143 7373
rect 5956 6563 5963 6583
rect 5956 6556 5983 6563
rect 5936 6187 5943 6253
rect 5936 6116 5943 6173
rect 5896 5916 5903 6073
rect 5916 6067 5923 6103
rect 5936 5916 5943 5933
rect 5956 5927 5963 6453
rect 5976 6387 5983 6556
rect 5996 6547 6003 6583
rect 6016 6576 6043 6583
rect 5976 5903 5983 6353
rect 5996 6307 6003 6393
rect 5996 6027 6003 6093
rect 5956 5896 5983 5903
rect 5896 5847 5903 5873
rect 5896 5667 5903 5733
rect 5916 5647 5923 5873
rect 5976 5667 5983 5896
rect 5976 5623 5983 5653
rect 5896 5436 5903 5593
rect 5876 5407 5883 5423
rect 5916 5407 5923 5433
rect 5936 5427 5943 5623
rect 5956 5616 5983 5623
rect 5836 5187 5843 5353
rect 5836 4983 5843 5153
rect 5816 4976 5843 4983
rect 5776 4696 5803 4703
rect 5796 4647 5803 4696
rect 5816 4587 5823 4976
rect 5836 4867 5843 4953
rect 5856 4936 5863 5273
rect 5876 5176 5883 5213
rect 5916 5176 5943 5183
rect 5896 5127 5903 5163
rect 5916 5047 5923 5073
rect 5936 4987 5943 5176
rect 5916 4956 5943 4963
rect 5896 4867 5903 4943
rect 5696 4576 5723 4583
rect 5676 3983 5683 4193
rect 5696 4147 5703 4576
rect 5716 4527 5723 4533
rect 5716 4476 5723 4513
rect 5756 4476 5763 4573
rect 5716 4016 5723 4193
rect 5756 4167 5763 4213
rect 5776 4207 5783 4453
rect 5796 4227 5803 4493
rect 5756 3996 5783 4003
rect 5676 3976 5703 3983
rect 5776 3967 5783 3996
rect 5856 3987 5863 4713
rect 5936 4707 5943 4956
rect 5956 4927 5963 5616
rect 5996 5603 6003 5853
rect 5976 5596 6003 5603
rect 5976 5407 5983 5596
rect 6016 5567 6023 6576
rect 6056 6563 6063 7053
rect 6076 7027 6083 7153
rect 6036 6556 6063 6563
rect 6036 6416 6043 6556
rect 6056 6123 6063 6383
rect 6076 6187 6083 6793
rect 6096 6147 6103 7356
rect 6156 7076 6163 7233
rect 6176 7187 6183 7373
rect 6196 7327 6203 7343
rect 6196 7127 6203 7313
rect 6216 7247 6223 7293
rect 6176 7027 6183 7063
rect 6116 6787 6123 6843
rect 6156 6743 6163 6843
rect 6136 6736 6163 6743
rect 6116 6547 6123 6593
rect 6136 6307 6143 6736
rect 6176 6647 6183 6993
rect 6196 6827 6203 6853
rect 6236 6707 6243 7073
rect 6256 7007 6263 7516
rect 6296 7507 6303 7563
rect 6276 7336 6283 7493
rect 6256 6767 6263 6933
rect 6296 6896 6303 7413
rect 6456 7376 6463 7453
rect 6476 7447 6483 7523
rect 6576 7463 6583 8173
rect 6616 8083 6623 8313
rect 6796 8187 6803 8813
rect 6856 8627 6863 8973
rect 6816 8567 6823 8613
rect 6816 8287 6823 8513
rect 6836 8503 6843 8593
rect 6876 8527 6883 8753
rect 6836 8496 6863 8503
rect 6916 8467 6923 8523
rect 6596 8076 6623 8083
rect 6596 8067 6603 8076
rect 6636 8063 6643 8113
rect 6636 8056 6663 8063
rect 6616 8027 6623 8043
rect 6596 7807 6603 7833
rect 6556 7456 6583 7463
rect 6376 7107 6383 7113
rect 6436 7107 6443 7153
rect 6456 7107 6463 7153
rect 6496 7096 6503 7233
rect 6556 7187 6563 7456
rect 6596 7343 6603 7563
rect 6616 7363 6623 7613
rect 6636 7576 6643 7613
rect 6636 7387 6643 7413
rect 6616 7356 6643 7363
rect 6576 7336 6603 7343
rect 6596 7207 6603 7336
rect 6636 7323 6643 7356
rect 6616 7316 6643 7323
rect 6656 7303 6663 8056
rect 6676 7327 6683 7933
rect 6696 7836 6703 8053
rect 6756 8043 6763 8093
rect 6816 8047 6823 8113
rect 6756 8036 6783 8043
rect 6716 7807 6723 7823
rect 6756 7816 6763 8013
rect 6636 7296 6663 7303
rect 6536 7096 6543 7113
rect 6316 6907 6323 7063
rect 6336 6876 6343 6993
rect 6356 6927 6363 7063
rect 6276 6847 6283 6863
rect 6156 6487 6163 6553
rect 6176 6427 6183 6583
rect 6196 6547 6203 6563
rect 6196 6407 6203 6513
rect 6276 6427 6283 6833
rect 6236 6396 6243 6413
rect 6056 6116 6083 6123
rect 6116 6116 6123 6173
rect 6076 6096 6103 6103
rect 6036 5647 6043 5933
rect 6036 5587 6043 5613
rect 5996 5423 6003 5553
rect 6056 5527 6063 5913
rect 6076 5767 6083 6096
rect 6136 6027 6143 6103
rect 6136 5947 6143 5973
rect 6096 5916 6123 5923
rect 6156 5916 6163 6013
rect 6176 5987 6183 6253
rect 6196 5916 6203 6273
rect 6216 6207 6223 6383
rect 6256 6376 6263 6393
rect 6216 6107 6223 6133
rect 6096 5887 6103 5916
rect 5996 5416 6023 5423
rect 5976 5247 5983 5273
rect 5996 5247 6003 5416
rect 5976 4883 5983 5233
rect 6016 5027 6023 5393
rect 6076 5156 6083 5253
rect 6096 5183 6103 5753
rect 6136 5747 6143 5903
rect 6156 5827 6163 5873
rect 6176 5847 6183 5903
rect 6116 5656 6123 5733
rect 6116 5307 6123 5373
rect 6116 5183 6123 5193
rect 6096 5176 6123 5183
rect 6136 5183 6143 5493
rect 6156 5207 6163 5553
rect 6136 5176 6163 5183
rect 6116 5156 6123 5176
rect 6156 5143 6163 5176
rect 6036 4947 6043 5113
rect 6056 5087 6063 5133
rect 6096 5127 6103 5143
rect 6136 5136 6163 5143
rect 6096 4987 6103 5033
rect 6056 4956 6063 4973
rect 5976 4876 6003 4883
rect 5936 4687 5943 4693
rect 5976 4667 5983 4853
rect 5896 4476 5903 4613
rect 5936 4476 5943 4533
rect 5956 4467 5963 4573
rect 5916 4447 5923 4463
rect 5976 4216 5983 4493
rect 5996 4247 6003 4876
rect 5876 4187 5883 4213
rect 5996 4187 6003 4203
rect 5916 3947 5923 3983
rect 6016 3707 6023 4133
rect 5676 3647 5683 3703
rect 5696 3507 5703 3573
rect 5616 3496 5643 3503
rect 5716 3483 5723 3703
rect 5736 3516 5743 3553
rect 5756 3536 5763 3573
rect 5776 3516 5783 3533
rect 5696 3476 5723 3483
rect 5696 3427 5703 3476
rect 4976 3196 5003 3203
rect 4896 2967 4903 3023
rect 4796 2756 4813 2763
rect 4696 2536 4703 2553
rect 4656 2207 4663 2283
rect 4696 2276 4703 2473
rect 4716 2303 4723 2713
rect 4736 2687 4743 2753
rect 4816 2707 4823 2753
rect 4736 2487 4743 2673
rect 4916 2623 4923 3093
rect 5156 3056 5163 3073
rect 4976 3016 4983 3053
rect 5256 3016 5283 3023
rect 5256 3007 5263 3016
rect 4936 2756 4943 2773
rect 5016 2743 5023 2753
rect 4996 2736 5023 2743
rect 4956 2687 4963 2723
rect 4896 2616 4923 2623
rect 4896 2303 4903 2616
rect 4976 2536 5003 2543
rect 4976 2407 4983 2536
rect 5036 2507 5043 2523
rect 4716 2296 4743 2303
rect 4896 2296 4923 2303
rect 4736 2263 4743 2296
rect 4716 2256 4743 2263
rect 4656 2076 4683 2083
rect 4596 1327 4603 1593
rect 4676 1387 4683 2076
rect 4616 1336 4643 1343
rect 4616 1247 4623 1336
rect 4676 1147 4683 1343
rect 4696 1267 4703 1323
rect 4616 1116 4623 1133
rect 4596 1067 4603 1083
rect 4716 867 4723 1373
rect 4476 376 4503 383
rect 4556 656 4583 663
rect 4476 343 4483 376
rect 4476 336 4503 343
rect 4296 156 4323 163
rect 4136 127 4143 143
rect 3876 -24 3903 -17
rect 4016 -24 4043 -17
rect 4136 -24 4143 13
rect 4296 -24 4303 156
rect 4516 156 4523 273
rect 4436 -24 4443 153
rect 4556 -17 4563 656
rect 4596 643 4603 813
rect 4616 647 4623 853
rect 4576 636 4603 643
rect 4576 616 4583 636
rect 4616 616 4623 633
rect 4596 607 4603 613
rect 4636 347 4643 603
rect 4656 167 4663 853
rect 4696 707 4703 803
rect 4736 383 4743 2256
rect 4856 2247 4863 2263
rect 4836 2096 4843 2133
rect 4816 1823 4823 2063
rect 4876 2047 4883 2083
rect 4796 1816 4823 1823
rect 4796 1147 4803 1816
rect 4916 1787 4923 2296
rect 5056 2283 5063 2553
rect 5036 2276 5063 2283
rect 5136 2267 5143 2913
rect 5156 2776 5163 2793
rect 5176 2747 5183 2763
rect 5176 2327 5183 2593
rect 5196 2583 5203 2783
rect 5216 2607 5223 2763
rect 5196 2576 5223 2583
rect 5256 2507 5263 2993
rect 5316 2887 5323 3003
rect 5276 2847 5283 2873
rect 5336 2863 5343 3173
rect 5316 2856 5343 2863
rect 5276 2567 5283 2573
rect 5216 2276 5223 2293
rect 4956 2076 4963 2093
rect 4996 2076 5003 2113
rect 4976 1747 4983 1783
rect 4936 1603 4943 1613
rect 4936 1596 4963 1603
rect 5036 1596 5043 1653
rect 5056 1627 5063 2233
rect 5076 1596 5103 1603
rect 4876 1303 4883 1353
rect 4896 1327 4903 1573
rect 5096 1567 5103 1596
rect 4956 1347 4963 1553
rect 5056 1336 5063 1353
rect 4816 1123 4823 1303
rect 4856 1296 4883 1303
rect 4836 1207 4843 1283
rect 5036 1267 5043 1323
rect 5076 1307 5083 1333
rect 4796 1116 4823 1123
rect 4756 1083 4763 1113
rect 4796 1096 4803 1116
rect 4756 1076 4783 1083
rect 4816 1067 4823 1083
rect 4816 827 4823 1053
rect 4836 847 4843 1133
rect 4856 1067 4863 1133
rect 4856 856 4863 893
rect 4876 807 4883 843
rect 4796 596 4803 633
rect 4816 616 4823 693
rect 4896 407 4903 853
rect 4916 427 4923 653
rect 4736 376 4763 383
rect 4536 -24 4563 -17
rect 4616 -17 4623 153
rect 4696 123 4703 173
rect 4676 116 4703 123
rect 4756 27 4763 376
rect 4856 367 4863 373
rect 4916 347 4923 413
rect 4876 207 4883 343
rect 4936 327 4943 773
rect 4956 347 4963 1173
rect 4996 1116 5023 1123
rect 5076 1116 5083 1133
rect 4976 1087 4983 1103
rect 4996 1067 5003 1116
rect 5036 1087 5043 1093
rect 5036 827 5043 843
rect 4996 667 5003 793
rect 4976 636 4983 653
rect 5056 643 5063 813
rect 5076 787 5083 843
rect 5016 636 5043 643
rect 5056 636 5083 643
rect 5036 607 5043 636
rect 5016 376 5023 393
rect 5056 376 5083 383
rect 4796 176 4823 183
rect 4796 27 4803 176
rect 4996 156 5023 163
rect 5036 156 5043 333
rect 5076 327 5083 376
rect 5136 187 5143 1913
rect 5156 927 5163 2253
rect 5176 2076 5183 2233
rect 5216 2076 5223 2093
rect 5236 1807 5243 2313
rect 5276 2267 5283 2553
rect 5296 2287 5303 2553
rect 5216 1776 5243 1783
rect 5196 1756 5213 1763
rect 5236 1647 5243 1776
rect 5176 1603 5183 1633
rect 5176 1596 5203 1603
rect 5256 1367 5263 2253
rect 5276 1607 5283 1653
rect 5196 1187 5203 1353
rect 5276 1316 5283 1393
rect 5296 1343 5303 2083
rect 5316 1596 5323 2856
rect 5356 2847 5363 3243
rect 5656 3127 5663 3233
rect 5516 3056 5543 3063
rect 5416 3016 5443 3023
rect 5436 2887 5443 3016
rect 5396 2263 5403 2833
rect 5436 2743 5443 2853
rect 5516 2767 5523 3056
rect 5696 2983 5703 3413
rect 5736 3236 5743 3473
rect 5767 3356 5773 3363
rect 5836 3207 5843 3513
rect 5716 3016 5723 3113
rect 5816 3023 5823 3053
rect 5796 3016 5823 3023
rect 5696 2976 5723 2983
rect 5416 2736 5443 2743
rect 5416 2556 5423 2713
rect 5396 2256 5423 2263
rect 5416 2056 5443 2063
rect 5416 1987 5423 2056
rect 5476 2056 5483 2093
rect 5456 2036 5463 2053
rect 5516 2043 5523 2693
rect 5536 2047 5543 2733
rect 5556 2556 5563 2763
rect 5616 2627 5623 2743
rect 5596 2576 5603 2613
rect 5576 2263 5583 2493
rect 5556 2256 5583 2263
rect 5616 2083 5623 2543
rect 5676 2487 5683 2553
rect 5696 2287 5703 2933
rect 5676 2087 5683 2093
rect 5596 2076 5623 2083
rect 5496 2036 5523 2043
rect 5336 1783 5343 1813
rect 5416 1796 5443 1803
rect 5336 1776 5363 1783
rect 5296 1336 5323 1343
rect 5216 1287 5223 1303
rect 5256 1267 5263 1303
rect 5316 1287 5323 1336
rect 5156 636 5163 693
rect 5196 636 5203 1173
rect 5236 1136 5243 1253
rect 5256 1116 5283 1123
rect 5276 1067 5283 1116
rect 5216 827 5223 893
rect 5276 887 5283 1053
rect 5256 827 5263 863
rect 5296 856 5303 1273
rect 5336 1267 5343 1353
rect 5316 1047 5323 1123
rect 5276 347 5283 843
rect 5196 183 5203 323
rect 5176 176 5203 183
rect 5156 156 5163 173
rect 4836 127 4843 143
rect 4616 -24 4643 -17
rect 4676 -24 4683 13
rect 4836 -24 4843 13
rect 5016 -17 5023 156
rect 5176 -17 5183 176
rect 5296 167 5303 653
rect 5356 607 5363 1393
rect 5376 1147 5383 1613
rect 5396 1307 5403 1593
rect 5436 1443 5443 1796
rect 5456 1767 5463 1973
rect 5496 1787 5503 2036
rect 5596 1847 5603 2076
rect 5616 2056 5643 2063
rect 5616 1827 5623 2056
rect 5676 2056 5683 2073
rect 5656 2036 5663 2053
rect 5696 2027 5703 2043
rect 5596 1796 5603 1813
rect 5636 1787 5643 1833
rect 5476 1587 5483 1773
rect 5536 1607 5543 1633
rect 5576 1596 5583 1673
rect 5616 1667 5623 1783
rect 5676 1607 5683 1813
rect 5696 1767 5703 1793
rect 5716 1747 5723 2976
rect 5736 2727 5743 2743
rect 5776 2607 5783 2743
rect 5736 2467 5743 2593
rect 5816 2556 5843 2563
rect 5736 2327 5743 2453
rect 5776 2276 5783 2473
rect 5736 1847 5743 2253
rect 5756 2247 5763 2263
rect 5736 1687 5743 1833
rect 5796 1827 5803 2263
rect 5756 1783 5763 1813
rect 5816 1803 5823 2313
rect 5836 2307 5843 2556
rect 5836 2227 5843 2293
rect 5856 2267 5863 3673
rect 5896 3627 5903 3703
rect 5916 3696 5943 3703
rect 5896 3207 5903 3223
rect 5836 2087 5843 2193
rect 5876 2083 5883 2873
rect 5896 2527 5903 3193
rect 5916 2927 5923 3696
rect 6016 3503 6023 3693
rect 6036 3527 6043 4913
rect 6116 4907 6123 4943
rect 6116 4847 6123 4893
rect 6136 4847 6143 5136
rect 6096 4707 6103 4733
rect 6056 4476 6063 4633
rect 6116 4527 6123 4683
rect 6076 4496 6083 4513
rect 6116 4447 6123 4513
rect 6136 4447 6143 4473
rect 6116 4227 6123 4433
rect 6156 4427 6163 5073
rect 6176 4287 6183 5813
rect 6216 5463 6223 6093
rect 6236 5767 6243 6353
rect 6276 6287 6283 6373
rect 6256 6116 6263 6133
rect 6236 5667 6243 5753
rect 6256 5607 6263 6073
rect 6276 5607 6283 6053
rect 6296 6003 6303 6713
rect 6396 6707 6403 6733
rect 6316 6067 6323 6693
rect 6336 6087 6343 6633
rect 6356 6547 6363 6583
rect 6356 6367 6363 6533
rect 6376 6403 6383 6553
rect 6396 6507 6403 6573
rect 6416 6547 6423 6713
rect 6436 6567 6443 6853
rect 6456 6827 6463 7093
rect 6556 7007 6563 7093
rect 6476 6876 6503 6883
rect 6436 6507 6443 6553
rect 6407 6416 6423 6423
rect 6376 6396 6403 6403
rect 6296 5996 6323 6003
rect 6296 5907 6303 5973
rect 6316 5927 6323 5996
rect 6376 5947 6383 6373
rect 6456 6367 6463 6693
rect 6476 6447 6483 6876
rect 6516 6827 6523 6933
rect 6536 6927 6543 6933
rect 6536 6876 6543 6913
rect 6556 6807 6563 6913
rect 6576 6887 6583 7033
rect 6576 6847 6583 6873
rect 6536 6596 6543 6693
rect 6576 6587 6583 6603
rect 6396 6167 6403 6293
rect 6416 6167 6423 6193
rect 6436 6187 6443 6293
rect 6456 6167 6463 6353
rect 6396 5947 6403 6153
rect 6416 6136 6423 6153
rect 6456 6136 6463 6153
rect 6476 6127 6483 6153
rect 6416 5923 6423 5993
rect 6396 5916 6423 5923
rect 6336 5847 6343 5903
rect 6376 5747 6383 5903
rect 6416 5887 6423 5893
rect 6336 5636 6343 5653
rect 6196 5456 6223 5463
rect 6196 4547 6203 5456
rect 6216 4707 6223 5193
rect 6236 4947 6243 5593
rect 6316 5527 6323 5623
rect 6276 5436 6283 5473
rect 6316 5156 6323 5413
rect 6256 4787 6263 4943
rect 6296 4867 6303 5123
rect 6336 4927 6343 5593
rect 6356 5547 6363 5623
rect 6356 5407 6363 5513
rect 6376 5407 6383 5433
rect 6356 5147 6363 5213
rect 6396 5183 6403 5593
rect 6436 5507 6443 6093
rect 6456 5887 6463 5993
rect 6456 5567 6463 5873
rect 6476 5647 6483 6033
rect 6496 6007 6503 6393
rect 6516 6107 6523 6553
rect 6596 6547 6603 7173
rect 6616 6567 6623 7073
rect 6636 6843 6643 7296
rect 6696 7187 6703 7593
rect 6716 7227 6723 7373
rect 6656 6876 6663 6973
rect 6716 6907 6723 6973
rect 6736 6876 6743 7673
rect 6776 7556 6783 8036
rect 6836 7987 6843 8023
rect 6856 7807 6863 8333
rect 6796 7447 6803 7543
rect 6636 6836 6663 6843
rect 6636 6707 6643 6753
rect 6556 6347 6563 6513
rect 6596 6347 6603 6383
rect 6636 6323 6643 6673
rect 6656 6627 6663 6836
rect 6676 6767 6683 6863
rect 6656 6587 6663 6613
rect 6676 6607 6683 6753
rect 6616 6316 6643 6323
rect 6616 6287 6623 6316
rect 6596 6187 6603 6273
rect 6536 6047 6543 6153
rect 6556 6007 6563 6173
rect 6596 6116 6603 6173
rect 6656 6163 6663 6433
rect 6676 6427 6683 6593
rect 6696 6587 6703 6773
rect 6716 6707 6723 6863
rect 6756 6627 6763 7313
rect 6776 7287 6783 7343
rect 6776 6927 6783 7213
rect 6776 6807 6783 6893
rect 6796 6867 6803 7393
rect 6816 7223 6823 7753
rect 6876 7727 6883 8433
rect 6936 8347 6943 9133
rect 6956 8407 6963 8433
rect 6916 8316 6923 8333
rect 6956 8316 6963 8393
rect 6976 8247 6983 9263
rect 7016 9256 7023 9493
rect 7036 9387 7043 9473
rect 7076 9087 7083 9273
rect 6996 8767 7003 9013
rect 7056 8927 7063 8963
rect 7036 8776 7043 8813
rect 7076 8763 7083 8953
rect 7016 8707 7023 8763
rect 7056 8756 7083 8763
rect 7096 8503 7103 9273
rect 7116 8547 7123 9973
rect 7136 9956 7163 9963
rect 7156 9927 7163 9956
rect 7176 9807 7183 10273
rect 7196 10267 7203 10416
rect 7196 9776 7203 9813
rect 7176 9727 7183 9743
rect 7176 9667 7183 9713
rect 7216 9667 7223 10233
rect 7216 9607 7223 9653
rect 7136 9447 7143 9463
rect 7176 9387 7183 9443
rect 7136 8907 7143 9373
rect 7236 9247 7243 10273
rect 7276 10216 7283 10253
rect 7296 10236 7303 10433
rect 7316 10347 7323 10423
rect 7356 10367 7363 10413
rect 7456 10407 7463 11873
rect 7516 11767 7523 11896
rect 7576 11863 7583 11913
rect 7716 11896 7743 11903
rect 7556 11856 7583 11863
rect 7476 11656 7483 11693
rect 7516 11547 7523 11753
rect 7576 11663 7583 11693
rect 7556 11656 7583 11663
rect 7476 10696 7483 10813
rect 7336 10236 7343 10313
rect 7456 10236 7463 10313
rect 7476 10263 7483 10553
rect 7496 10287 7503 11433
rect 7576 11407 7583 11413
rect 7576 11196 7603 11203
rect 7596 11087 7603 11196
rect 7656 11163 7663 11893
rect 7716 11847 7723 11896
rect 7716 11827 7723 11833
rect 7756 11727 7763 11863
rect 7836 11676 7863 11683
rect 7896 11676 7903 11793
rect 7936 11767 7943 11843
rect 7956 11687 7963 11873
rect 8136 11863 8143 11893
rect 8236 11887 8243 11913
rect 8116 11856 8143 11863
rect 8096 11827 8103 11843
rect 7676 11183 7683 11393
rect 7716 11387 7723 11663
rect 7836 11467 7843 11676
rect 8056 11676 8063 11693
rect 8096 11676 8103 11753
rect 8136 11707 8143 11773
rect 8296 11707 8303 11903
rect 8836 11896 8843 11913
rect 8676 11863 8683 11873
rect 8136 11676 8143 11693
rect 8076 11627 8083 11663
rect 7836 11427 7843 11453
rect 8116 11447 8123 11663
rect 7836 11387 7843 11413
rect 7676 11176 7703 11183
rect 7696 11167 7703 11176
rect 7656 11156 7683 11163
rect 7516 10907 7523 11033
rect 7636 10943 7643 11033
rect 7616 10936 7643 10943
rect 7556 10916 7563 10933
rect 7576 10876 7603 10883
rect 7576 10463 7583 10773
rect 7596 10707 7603 10876
rect 7636 10727 7643 10936
rect 7656 10907 7663 10923
rect 7676 10867 7683 11156
rect 7716 11067 7723 11373
rect 7776 11287 7783 11383
rect 7916 11307 7923 11393
rect 7736 11087 7743 11183
rect 7776 11087 7783 11273
rect 7896 11196 7903 11233
rect 7936 11196 7943 11353
rect 7976 11196 7983 11313
rect 8036 11267 8043 11413
rect 8216 11383 8223 11693
rect 8236 11627 8243 11693
rect 8316 11676 8323 11773
rect 8256 11647 8263 11663
rect 8236 11427 8243 11613
rect 8196 11376 8223 11383
rect 8196 11327 8203 11376
rect 8196 11307 8203 11313
rect 7916 11167 7923 11183
rect 7956 11163 7963 11183
rect 7956 11156 7983 11163
rect 7676 10736 7703 10743
rect 7676 10727 7683 10736
rect 7676 10667 7683 10713
rect 7736 10703 7743 10773
rect 7716 10696 7743 10703
rect 7556 10456 7583 10463
rect 7536 10427 7543 10443
rect 7476 10256 7503 10263
rect 7496 10236 7503 10256
rect 7316 9923 7323 10213
rect 7476 10203 7483 10223
rect 7516 10216 7523 10253
rect 7476 10196 7503 10203
rect 7456 10127 7463 10193
rect 7336 9947 7343 9953
rect 7336 9927 7343 9933
rect 7296 9916 7323 9923
rect 7076 8496 7103 8503
rect 6936 8007 6943 8193
rect 6996 8007 7003 8023
rect 7016 7947 7023 8233
rect 6956 7836 6983 7843
rect 6876 7567 6883 7713
rect 6856 7487 6863 7543
rect 6876 7347 6883 7453
rect 6896 7407 6903 7793
rect 6976 7787 6983 7836
rect 6996 7807 7003 7853
rect 6956 7356 6963 7453
rect 6976 7367 6983 7673
rect 6996 7387 7003 7753
rect 7016 7607 7023 7893
rect 7036 7667 7043 8293
rect 7056 7567 7063 8273
rect 7076 7687 7083 8496
rect 7116 8467 7123 8503
rect 7136 8336 7143 8353
rect 7096 8183 7103 8313
rect 7116 8287 7123 8303
rect 7116 8227 7123 8273
rect 7096 8176 7123 8183
rect 7116 7856 7123 8176
rect 7136 8007 7143 8193
rect 7156 8087 7163 9233
rect 7196 9227 7203 9243
rect 7256 9067 7263 9853
rect 7276 9527 7283 9793
rect 7276 9167 7283 9393
rect 7176 8227 7183 9033
rect 7196 8847 7203 8983
rect 7196 8816 7243 8823
rect 7196 8807 7203 8816
rect 7256 8796 7263 9033
rect 7296 9027 7303 9916
rect 7316 9776 7323 9793
rect 7336 9567 7343 9743
rect 7336 9476 7343 9513
rect 7396 9483 7403 9713
rect 7416 9587 7423 9953
rect 7456 9943 7463 10113
rect 7436 9936 7463 9943
rect 7376 9476 7403 9483
rect 7316 9207 7323 9463
rect 7276 8807 7283 8833
rect 7316 8643 7323 9053
rect 7336 8847 7343 9433
rect 7376 9276 7383 9373
rect 7396 9067 7403 9263
rect 7436 9207 7443 9913
rect 7456 9147 7463 9936
rect 7476 9743 7483 9933
rect 7496 9887 7503 10196
rect 7516 9756 7523 9793
rect 7576 9787 7583 10393
rect 7596 10387 7603 10453
rect 7556 9763 7563 9773
rect 7556 9756 7583 9763
rect 7496 9743 7503 9753
rect 7576 9747 7583 9756
rect 7476 9736 7503 9743
rect 7476 9507 7483 9736
rect 7536 9707 7543 9743
rect 7496 9647 7503 9673
rect 7476 9347 7483 9473
rect 7476 9123 7483 9313
rect 7496 9267 7503 9633
rect 7516 9307 7523 9633
rect 7556 9447 7563 9493
rect 7596 9487 7603 9973
rect 7616 9467 7623 10633
rect 7676 10436 7683 10493
rect 7636 10236 7643 10413
rect 7676 10236 7683 10393
rect 7696 10387 7703 10403
rect 7656 9987 7663 10223
rect 7696 10216 7703 10253
rect 7636 9807 7643 9963
rect 7656 9907 7663 9943
rect 7656 9783 7663 9873
rect 7716 9783 7723 10013
rect 7636 9776 7663 9783
rect 7696 9776 7723 9783
rect 7596 9327 7603 9443
rect 7636 9367 7643 9776
rect 7696 9756 7703 9776
rect 7676 9723 7683 9743
rect 7716 9736 7723 9753
rect 7656 9716 7683 9723
rect 7576 9276 7583 9293
rect 7556 9256 7563 9273
rect 7476 9116 7503 9123
rect 7456 9007 7463 9113
rect 7376 8907 7383 9003
rect 7376 8803 7383 8873
rect 7436 8867 7443 8983
rect 7456 8807 7463 8993
rect 7356 8796 7383 8803
rect 7396 8796 7423 8803
rect 7316 8636 7343 8643
rect 7196 8507 7203 8633
rect 7196 8127 7203 8493
rect 7156 7967 7163 8043
rect 7196 8036 7203 8093
rect 7176 7927 7183 8023
rect 7096 7807 7103 7823
rect 7036 7523 7043 7543
rect 7036 7516 7063 7523
rect 6816 7216 6843 7223
rect 6836 7096 6843 7216
rect 6776 6596 6783 6693
rect 6696 6267 6703 6393
rect 6716 6387 6723 6583
rect 6736 6407 6743 6533
rect 6756 6527 6763 6583
rect 6816 6567 6823 7053
rect 6836 7027 6843 7053
rect 6856 6887 6863 7083
rect 6896 6903 6903 7353
rect 6976 7336 7003 7343
rect 6916 7047 6923 7093
rect 6876 6896 6903 6903
rect 6876 6876 6883 6896
rect 6916 6876 6923 6913
rect 6776 6396 6783 6533
rect 6816 6427 6823 6493
rect 6756 6307 6763 6383
rect 6796 6376 6803 6393
rect 6816 6347 6823 6373
rect 6836 6307 6843 6873
rect 6856 6447 6863 6853
rect 6896 6827 6903 6863
rect 6936 6856 6943 7313
rect 6996 6943 7003 7336
rect 7036 7127 7043 7193
rect 6976 6936 7003 6943
rect 6896 6727 6903 6813
rect 6956 6687 6963 6713
rect 6976 6647 6983 6936
rect 6936 6607 6943 6633
rect 6896 6596 6923 6603
rect 6856 6347 6863 6413
rect 6876 6367 6883 6413
rect 6656 6156 6683 6163
rect 6636 6107 6643 6123
rect 6576 6087 6583 6103
rect 6536 5916 6543 5973
rect 6496 5827 6503 5913
rect 6516 5883 6523 5913
rect 6516 5876 6543 5883
rect 6516 5636 6523 5853
rect 6496 5547 6503 5623
rect 6496 5427 6503 5533
rect 6376 5176 6403 5183
rect 6276 4543 6283 4813
rect 6336 4696 6343 4713
rect 6316 4567 6323 4683
rect 6276 4536 6303 4543
rect 6196 4443 6203 4533
rect 6236 4456 6243 4493
rect 6196 4436 6223 4443
rect 6176 4267 6183 4273
rect 6136 4216 6143 4253
rect 6056 3996 6063 4033
rect 6096 3996 6103 4013
rect 6116 3976 6123 4173
rect 5996 3496 6023 3503
rect 6056 3487 6063 3513
rect 6076 3507 6083 3573
rect 6096 3567 6103 3913
rect 6156 3687 6163 3703
rect 5956 2987 5963 3023
rect 5916 2687 5923 2753
rect 5936 2707 5943 2763
rect 5976 2756 5983 2793
rect 6036 2747 6043 2813
rect 5896 2263 5903 2513
rect 5936 2276 5943 2653
rect 5956 2556 5963 2613
rect 6036 2556 6043 2633
rect 5976 2327 5983 2543
rect 6056 2343 6063 3253
rect 6096 3223 6103 3553
rect 6136 3536 6143 3573
rect 6156 3523 6163 3533
rect 6176 3523 6183 3693
rect 6156 3516 6183 3523
rect 6096 3216 6123 3223
rect 6036 2336 6063 2343
rect 5896 2256 5913 2263
rect 5956 2127 5963 2263
rect 5856 2076 5883 2083
rect 5896 2076 5923 2083
rect 5796 1796 5823 1803
rect 5756 1776 5783 1783
rect 5696 1596 5703 1613
rect 5736 1596 5743 1653
rect 5436 1436 5463 1443
rect 5376 1107 5383 1133
rect 5396 1127 5403 1293
rect 5436 1116 5443 1133
rect 5436 856 5443 1033
rect 5456 947 5463 1436
rect 5496 1296 5503 1333
rect 5676 1147 5683 1593
rect 5756 1576 5783 1583
rect 5716 1207 5723 1573
rect 5556 1087 5563 1123
rect 5676 1116 5683 1133
rect 5396 636 5403 673
rect 5456 643 5463 843
rect 5556 827 5563 1073
rect 5716 827 5723 873
rect 5756 827 5763 1113
rect 5776 867 5783 1576
rect 5796 1567 5803 1593
rect 5816 1407 5823 1763
rect 5836 1316 5843 1453
rect 5856 1367 5863 2076
rect 5916 2047 5923 2076
rect 5876 1387 5883 2043
rect 5816 1287 5823 1303
rect 5896 1247 5903 2033
rect 5936 1403 5943 2053
rect 5956 1707 5963 2093
rect 6036 1823 6043 2336
rect 6056 2083 6063 2313
rect 6076 2107 6083 3213
rect 6116 2867 6123 3023
rect 6196 2847 6203 4093
rect 6216 3987 6223 4413
rect 6236 3667 6243 4233
rect 6156 2687 6163 2743
rect 6176 2536 6183 2613
rect 6196 2607 6203 2743
rect 6236 2667 6243 3593
rect 6256 3167 6263 4373
rect 6296 4023 6303 4536
rect 6356 4487 6363 4973
rect 6376 4307 6383 5176
rect 6396 4647 6403 4943
rect 6416 4907 6423 5413
rect 6456 5407 6463 5423
rect 6536 5407 6543 5876
rect 6556 5727 6563 5903
rect 6596 5896 6603 5933
rect 6436 5156 6443 5173
rect 6476 5156 6483 5393
rect 6396 4496 6403 4513
rect 6416 4447 6423 4463
rect 6336 4196 6343 4213
rect 6376 4163 6383 4293
rect 6396 4207 6403 4393
rect 6436 4227 6443 5013
rect 6456 5007 6463 5123
rect 6496 5047 6503 5143
rect 6516 4887 6523 5173
rect 6556 5007 6563 5553
rect 6576 5267 6583 5833
rect 6616 5707 6623 6073
rect 6636 5587 6643 6033
rect 6656 5847 6663 6113
rect 6676 6047 6683 6156
rect 6676 5643 6683 5993
rect 6696 5927 6703 6093
rect 6736 6087 6743 6253
rect 6816 6116 6823 6253
rect 6856 6116 6863 6153
rect 6787 6096 6803 6103
rect 6716 5927 6723 6033
rect 6736 5967 6743 6033
rect 6756 5936 6763 5953
rect 6796 5916 6803 5933
rect 6656 5636 6683 5643
rect 6696 5627 6703 5893
rect 6676 5596 6703 5603
rect 6656 5436 6663 5493
rect 6596 5187 6603 5423
rect 6636 5387 6643 5423
rect 6676 5367 6683 5573
rect 6696 5407 6703 5596
rect 6716 5267 6723 5893
rect 6816 5867 6823 5933
rect 6836 5847 6843 6073
rect 6856 5787 6863 6013
rect 6676 5156 6683 5253
rect 6716 5156 6723 5193
rect 6636 5107 6643 5153
rect 6756 5143 6763 5653
rect 6796 5456 6803 5693
rect 6876 5663 6883 6313
rect 6896 6087 6903 6596
rect 6956 6596 6963 6613
rect 6916 6407 6923 6433
rect 6956 6416 6963 6433
rect 6936 6396 6943 6413
rect 6856 5656 6883 5663
rect 6856 5636 6863 5656
rect 6816 5487 6823 5613
rect 6836 5603 6843 5623
rect 6896 5607 6903 5993
rect 6916 5923 6923 6233
rect 6936 6107 6943 6133
rect 6956 6127 6963 6333
rect 6996 6267 7003 6913
rect 7016 6147 7023 6953
rect 7036 6927 7043 6973
rect 7036 6227 7043 6673
rect 7056 6667 7063 7516
rect 7076 7467 7083 7533
rect 7076 7207 7083 7353
rect 7096 7327 7103 7733
rect 7136 7667 7143 7823
rect 7116 7107 7123 7493
rect 7176 7427 7183 7813
rect 7196 7647 7203 7993
rect 7216 7747 7223 7833
rect 7236 7647 7243 8573
rect 7296 8496 7313 8503
rect 7256 8407 7263 8453
rect 7256 7723 7263 8393
rect 7276 8387 7283 8483
rect 7276 8316 7303 8323
rect 7276 7747 7283 8273
rect 7296 8147 7303 8316
rect 7256 7716 7283 7723
rect 7196 7467 7203 7543
rect 7236 7536 7263 7543
rect 7136 7356 7143 7393
rect 7176 7376 7183 7393
rect 7176 7336 7203 7343
rect 7076 7076 7103 7083
rect 7096 7047 7103 7076
rect 7136 6947 7143 7293
rect 7176 7143 7183 7336
rect 7236 7267 7243 7393
rect 7256 7227 7263 7536
rect 7276 7307 7283 7716
rect 7296 7527 7303 8133
rect 7336 7927 7343 8636
rect 7356 8327 7363 8796
rect 7376 8367 7383 8693
rect 7396 8607 7403 8796
rect 7396 8527 7403 8593
rect 7476 8547 7483 9053
rect 7496 8987 7503 9116
rect 7396 8507 7403 8513
rect 7376 8267 7383 8273
rect 7376 8036 7383 8253
rect 7396 8147 7403 8373
rect 7416 8347 7423 8533
rect 7496 8467 7503 8833
rect 7516 8487 7523 8893
rect 7536 8867 7543 9233
rect 7636 9127 7643 9353
rect 7556 8887 7563 9053
rect 7616 8996 7623 9013
rect 7596 8847 7603 8953
rect 7656 8907 7663 9716
rect 7676 9267 7683 9653
rect 7736 9643 7743 10393
rect 7756 10267 7763 10393
rect 7756 10207 7763 10253
rect 7756 9667 7763 9953
rect 7736 9636 7763 9643
rect 7736 9476 7743 9493
rect 7756 9487 7763 9636
rect 7596 8816 7603 8833
rect 7616 8796 7623 8853
rect 7416 8036 7423 8233
rect 7356 8007 7363 8023
rect 7436 7847 7443 8453
rect 7476 8307 7483 8313
rect 7456 8267 7463 8283
rect 7456 8007 7463 8253
rect 7496 8247 7503 8283
rect 7556 8036 7563 8573
rect 7636 8563 7643 8853
rect 7656 8807 7663 8833
rect 7676 8787 7683 9253
rect 7696 8667 7703 9433
rect 7716 9307 7723 9473
rect 7776 9307 7783 10853
rect 7856 10703 7863 10793
rect 7916 10743 7923 10913
rect 7896 10736 7923 10743
rect 7856 10696 7883 10703
rect 7736 9227 7743 9263
rect 7756 9127 7763 9293
rect 7616 8556 7643 8563
rect 7616 8527 7623 8556
rect 7656 8516 7663 8653
rect 7576 8503 7583 8513
rect 7696 8503 7703 8593
rect 7576 8496 7603 8503
rect 7576 8267 7583 8413
rect 7596 8027 7603 8043
rect 7536 8007 7543 8023
rect 7576 7967 7583 8023
rect 7496 7887 7503 7953
rect 7516 7843 7523 7893
rect 7536 7856 7543 7873
rect 7496 7836 7523 7843
rect 7496 7827 7503 7836
rect 7596 7827 7603 7873
rect 7296 7467 7303 7513
rect 7316 7347 7323 7633
rect 7356 7336 7363 7593
rect 7376 7563 7383 7793
rect 7456 7576 7483 7583
rect 7376 7556 7403 7563
rect 7436 7447 7443 7553
rect 7476 7427 7483 7576
rect 7376 7347 7383 7373
rect 7396 7336 7423 7343
rect 7376 7316 7383 7333
rect 7416 7307 7423 7336
rect 7176 7136 7203 7143
rect 7196 7007 7203 7136
rect 7096 6876 7123 6883
rect 7136 6876 7143 6933
rect 7056 6247 7063 6553
rect 7036 6127 7043 6153
rect 7076 6127 7083 6853
rect 7116 6827 7123 6876
rect 7116 6607 7123 6713
rect 7156 6596 7163 6653
rect 7196 6587 7203 6993
rect 7216 6907 7223 6953
rect 7136 6427 7143 6583
rect 7216 6427 7223 6793
rect 7236 6707 7243 6893
rect 7256 6876 7263 6933
rect 7296 6876 7303 6973
rect 7316 6856 7323 6873
rect 7276 6847 7283 6853
rect 7276 6747 7283 6793
rect 7336 6767 7343 7013
rect 7116 6396 7143 6403
rect 7116 6387 7123 6396
rect 7216 6396 7223 6413
rect 7116 6143 7123 6373
rect 7156 6327 7163 6383
rect 7096 6136 7123 6143
rect 6936 5987 6943 6093
rect 6956 5947 6963 6113
rect 7016 6067 7023 6103
rect 6916 5916 6943 5923
rect 6976 5916 6983 6013
rect 7016 5916 7023 6033
rect 7056 5907 7063 6073
rect 7076 6007 7083 6093
rect 7096 6007 7103 6136
rect 6956 5867 6963 5903
rect 6996 5847 7003 5893
rect 7076 5867 7083 5893
rect 6916 5627 6923 5653
rect 6836 5596 6863 5603
rect 6836 5423 6843 5453
rect 6856 5427 6863 5596
rect 6936 5587 6943 5833
rect 6996 5747 7003 5833
rect 6996 5627 7003 5693
rect 6816 5416 6843 5423
rect 6796 5167 6803 5273
rect 6696 5107 6703 5143
rect 6736 5136 6763 5143
rect 6636 4963 6643 5013
rect 6616 4956 6643 4963
rect 6536 4903 6543 4953
rect 6596 4927 6603 4943
rect 6536 4896 6563 4903
rect 6536 4663 6543 4713
rect 6556 4707 6563 4896
rect 6596 4667 6603 4913
rect 6636 4727 6643 4956
rect 6516 4656 6543 4663
rect 6496 4547 6503 4643
rect 6556 4496 6563 4613
rect 6356 4156 6383 4163
rect 6396 4047 6403 4193
rect 6436 4147 6443 4213
rect 6456 4187 6463 4233
rect 6536 4216 6543 4233
rect 6596 4207 6603 4413
rect 6296 4016 6323 4023
rect 6316 3967 6323 4016
rect 6396 3983 6403 4033
rect 6436 3996 6443 4133
rect 6496 3996 6503 4033
rect 6396 3976 6423 3983
rect 6396 3727 6403 3853
rect 6396 3703 6403 3713
rect 6376 3696 6403 3703
rect 6276 3516 6303 3523
rect 6336 3516 6343 3653
rect 6276 3407 6283 3516
rect 6316 3267 6323 3503
rect 6476 3447 6483 3983
rect 6536 3716 6543 3753
rect 6556 3703 6563 3973
rect 6596 3716 6603 4153
rect 6516 3567 6523 3703
rect 6556 3696 6583 3703
rect 6576 3536 6583 3553
rect 6616 3543 6623 4433
rect 6656 4407 6663 4683
rect 6696 4447 6703 5033
rect 6756 4987 6763 5136
rect 6756 4956 6763 4973
rect 6776 4867 6783 4943
rect 6716 4456 6723 4833
rect 6816 4743 6823 5273
rect 6796 4736 6823 4743
rect 6736 4436 6743 4553
rect 6776 4427 6783 4443
rect 6716 4223 6723 4393
rect 6716 4216 6743 4223
rect 6736 4187 6743 4216
rect 6656 4176 6703 4183
rect 6636 4027 6643 4053
rect 6656 3996 6663 4176
rect 6756 4127 6763 4183
rect 6676 4016 6683 4033
rect 6696 3996 6703 4053
rect 6796 4003 6803 4736
rect 6836 4723 6843 5253
rect 6856 5067 6863 5393
rect 6896 5156 6903 5353
rect 6936 5167 6943 5513
rect 7016 5507 7023 5643
rect 7076 5607 7083 5623
rect 6956 5416 6983 5423
rect 6856 4947 6863 5053
rect 6816 4716 6843 4723
rect 6816 4696 6823 4716
rect 6876 4367 6883 5133
rect 6916 5127 6923 5143
rect 6916 4976 6923 4993
rect 6896 4387 6903 4893
rect 6916 4547 6923 4693
rect 6916 4496 6923 4533
rect 6876 4067 6883 4163
rect 6896 4127 6903 4183
rect 6956 4087 6963 4713
rect 6976 4587 6983 5416
rect 6996 5127 7003 5153
rect 6996 4687 7003 4953
rect 7036 4927 7043 5573
rect 7056 5027 7063 5573
rect 7096 5247 7103 5953
rect 7116 5627 7123 6113
rect 7136 6107 7143 6273
rect 7156 6083 7163 6253
rect 7196 6247 7203 6383
rect 7136 6076 7163 6083
rect 7136 5887 7143 6076
rect 7176 6007 7183 6233
rect 7196 6147 7203 6233
rect 7216 6116 7223 6193
rect 7236 6167 7243 6693
rect 7276 6616 7283 6733
rect 7356 6647 7363 7293
rect 7376 6747 7383 6953
rect 7396 6847 7403 6993
rect 7416 6783 7423 6953
rect 7396 6776 7423 6783
rect 7316 6616 7343 6623
rect 7256 6287 7263 6533
rect 7276 6207 7283 6393
rect 7196 6047 7203 6103
rect 7256 6083 7263 6093
rect 7236 6076 7263 6083
rect 7156 5916 7163 5993
rect 7196 5916 7223 5923
rect 7136 5603 7143 5633
rect 7116 5596 7143 5603
rect 7116 5347 7123 5596
rect 7156 5343 7163 5873
rect 7216 5767 7223 5916
rect 7216 5607 7223 5623
rect 7236 5567 7243 6076
rect 7256 5887 7263 6033
rect 7276 5647 7283 6133
rect 7296 5727 7303 6603
rect 7336 6423 7343 6616
rect 7336 6416 7363 6423
rect 7376 6396 7383 6713
rect 7236 5436 7243 5513
rect 7256 5507 7263 5623
rect 7176 5416 7183 5433
rect 7216 5347 7223 5423
rect 7156 5336 7183 5343
rect 7076 5156 7083 5233
rect 7156 5143 7163 5173
rect 7136 5136 7163 5143
rect 7076 4683 7083 4913
rect 7096 4867 7103 5123
rect 7136 4976 7143 5013
rect 7076 4676 7103 4683
rect 7076 4663 7083 4676
rect 6976 4327 6983 4573
rect 7016 4507 7023 4663
rect 7056 4656 7083 4663
rect 6796 3996 6813 4003
rect 6856 3996 6863 4013
rect 6896 3996 6903 4013
rect 6996 3987 7003 4173
rect 7016 4167 7023 4493
rect 7036 4467 7043 4643
rect 7116 4527 7123 4933
rect 7156 4783 7163 4993
rect 7176 4947 7183 5336
rect 7136 4776 7163 4783
rect 7136 4667 7143 4776
rect 7136 4476 7143 4593
rect 7076 4447 7083 4463
rect 7096 4196 7103 4213
rect 7116 4167 7123 4183
rect 6636 3716 6643 3953
rect 6736 3747 6743 3973
rect 6596 3536 6623 3543
rect 6287 3236 6303 3243
rect 6296 3147 6303 3236
rect 6496 3223 6503 3453
rect 6476 3216 6503 3223
rect 6256 3036 6263 3093
rect 6236 2556 6263 2563
rect 6216 2527 6223 2543
rect 6156 2267 6163 2303
rect 6176 2267 6183 2283
rect 6156 2227 6163 2233
rect 6056 2076 6083 2083
rect 6116 2076 6123 2093
rect 6096 2047 6103 2063
rect 6036 1816 6063 1823
rect 5956 1596 5963 1693
rect 5976 1427 5983 1803
rect 6036 1767 6043 1783
rect 5916 1396 5943 1403
rect 5856 823 5863 1193
rect 5896 1096 5903 1193
rect 5916 1127 5923 1396
rect 5956 1187 5963 1253
rect 5956 1116 5963 1173
rect 5976 1107 5983 1353
rect 5836 816 5863 823
rect 5436 636 5463 643
rect 5456 343 5463 513
rect 5476 387 5483 653
rect 5636 647 5643 803
rect 5756 707 5763 813
rect 5436 336 5463 343
rect 5456 227 5463 336
rect 5196 156 5223 163
rect 5216 -17 5223 156
rect 5516 116 5523 393
rect 5536 363 5543 633
rect 5676 607 5683 643
rect 5756 636 5763 693
rect 5616 376 5643 383
rect 5536 356 5563 363
rect 5636 347 5643 376
rect 5536 136 5543 153
rect 5576 123 5583 173
rect 5636 147 5643 333
rect 5736 323 5743 413
rect 5816 367 5823 613
rect 5856 587 5863 816
rect 5996 727 6003 1593
rect 6056 1447 6063 1816
rect 6096 1523 6103 1563
rect 6136 1556 6143 1673
rect 6156 1583 6163 2213
rect 6236 1887 6243 2153
rect 6256 2107 6263 2556
rect 6276 2167 6283 3133
rect 6476 3067 6483 3216
rect 6496 3036 6503 3153
rect 6336 2787 6343 3033
rect 6336 2763 6343 2773
rect 6336 2756 6363 2763
rect 6336 2747 6343 2756
rect 6416 2736 6433 2743
rect 6356 2556 6363 2573
rect 6416 2567 6423 2613
rect 6376 2507 6383 2543
rect 6416 2536 6423 2553
rect 6436 2507 6443 2733
rect 6456 2687 6463 2753
rect 6476 2567 6483 3033
rect 6536 2727 6543 3533
rect 6596 3247 6603 3536
rect 6716 3527 6723 3723
rect 6736 3627 6743 3733
rect 6916 3683 6923 3753
rect 7056 3736 7063 3773
rect 6896 3676 6923 3683
rect 6876 3536 6883 3613
rect 6716 3503 6723 3513
rect 7016 3503 7023 3723
rect 6696 3496 6723 3503
rect 6996 3496 7023 3503
rect 6676 3236 6683 3313
rect 6656 3187 6663 3223
rect 6696 3207 6703 3223
rect 6716 3127 6723 3496
rect 6656 3036 6663 3053
rect 6696 3036 6703 3073
rect 6636 3016 6643 3033
rect 6716 3003 6723 3053
rect 6796 3027 6803 3393
rect 7016 3363 7023 3496
rect 7076 3487 7083 3773
rect 7007 3356 7023 3363
rect 6816 3207 6823 3243
rect 6836 3227 6843 3263
rect 6856 3207 6863 3243
rect 6816 3023 6823 3173
rect 6896 3036 6923 3043
rect 6816 3016 6843 3023
rect 6696 2996 6723 3003
rect 6596 2776 6623 2783
rect 6576 2727 6583 2763
rect 6616 2747 6623 2776
rect 6516 2307 6523 2393
rect 6536 2307 6543 2713
rect 6576 2556 6583 2693
rect 6296 2227 6303 2253
rect 6376 2247 6383 2283
rect 6516 2167 6523 2263
rect 6576 2263 6583 2373
rect 6556 2256 6583 2263
rect 6516 2107 6523 2153
rect 6276 2056 6283 2073
rect 6316 2056 6323 2093
rect 6196 1796 6203 1813
rect 6236 1796 6243 1853
rect 6196 1727 6203 1753
rect 6156 1576 6183 1583
rect 6096 1516 6123 1523
rect 6016 643 6023 1433
rect 6116 1347 6123 1516
rect 6176 1507 6183 1576
rect 6056 883 6063 1323
rect 6096 1287 6103 1313
rect 6076 1136 6123 1143
rect 6076 1083 6083 1136
rect 6136 1116 6143 1173
rect 6076 1076 6103 1083
rect 6036 876 6063 883
rect 6036 827 6043 876
rect 6056 807 6063 843
rect 6096 836 6103 1076
rect 6116 787 6123 823
rect 5996 636 6023 643
rect 5936 356 5943 373
rect 5996 347 6003 636
rect 6036 616 6043 633
rect 6156 627 6163 1313
rect 6176 1167 6183 1373
rect 6196 1303 6203 1713
rect 6216 1647 6223 1763
rect 6276 1327 6283 1873
rect 6396 1807 6403 2093
rect 6436 1796 6443 2073
rect 6476 1987 6483 2033
rect 6356 1596 6363 1613
rect 6296 1576 6303 1593
rect 6376 1587 6383 1783
rect 6416 1747 6423 1763
rect 6456 1547 6463 1753
rect 6476 1547 6483 1973
rect 6496 1607 6503 2053
rect 6516 1747 6523 1873
rect 6536 1623 6543 2253
rect 6556 2127 6563 2256
rect 6596 2107 6603 2513
rect 6636 2487 6643 2543
rect 6556 2087 6563 2093
rect 6596 2067 6603 2093
rect 6616 1787 6623 1873
rect 6596 1747 6603 1783
rect 6536 1616 6563 1623
rect 6536 1547 6543 1563
rect 6376 1307 6383 1393
rect 6196 1296 6223 1303
rect 6016 407 6023 603
rect 5736 316 5763 323
rect 5916 267 5923 343
rect 6016 327 6023 373
rect 6136 356 6143 553
rect 6176 327 6183 1093
rect 6216 616 6223 1233
rect 6236 1127 6243 1283
rect 6256 1247 6263 1303
rect 6276 1096 6283 1133
rect 6336 1116 6343 1193
rect 6356 1107 6363 1213
rect 6256 807 6263 823
rect 6256 767 6263 793
rect 6276 403 6283 693
rect 6376 667 6383 1253
rect 6396 627 6403 1533
rect 6416 847 6423 1313
rect 6496 1303 6503 1533
rect 6476 1296 6503 1303
rect 6456 1136 6463 1153
rect 6496 1116 6503 1273
rect 6476 863 6483 1103
rect 6476 856 6503 863
rect 6416 823 6423 833
rect 6416 816 6443 823
rect 6456 667 6463 673
rect 6456 636 6463 653
rect 6436 587 6443 623
rect 6476 547 6483 823
rect 6496 807 6503 856
rect 6516 827 6523 1373
rect 6536 1307 6543 1413
rect 6536 647 6543 1153
rect 6256 396 6283 403
rect 6256 347 6263 396
rect 6276 356 6303 363
rect 5696 156 5703 213
rect 5756 136 5783 143
rect 5776 127 5783 136
rect 5876 127 5883 193
rect 5956 156 5963 313
rect 6116 187 6123 323
rect 6136 176 6163 183
rect 5936 127 5943 143
rect 6116 127 6123 143
rect 5556 116 5583 123
rect 6156 27 6163 176
rect 6256 156 6263 333
rect 6276 307 6283 356
rect 6336 336 6363 343
rect 6336 323 6343 336
rect 6316 316 6343 323
rect 6296 156 6303 193
rect 6496 156 6503 573
rect 6536 347 6543 413
rect 6556 347 6563 1616
rect 6576 1567 6583 1593
rect 6596 1447 6603 1573
rect 6636 1387 6643 2293
rect 6656 2107 6663 2913
rect 6696 2487 6703 2996
rect 6716 2767 6723 2793
rect 6816 2787 6823 3016
rect 6716 2527 6723 2753
rect 6736 2687 6743 2743
rect 6676 2247 6683 2473
rect 6736 2427 6743 2673
rect 6776 2627 6783 2723
rect 6756 2507 6763 2523
rect 6756 2327 6763 2493
rect 6696 2187 6703 2283
rect 6696 2076 6703 2133
rect 6716 2043 6723 2113
rect 6696 2036 6723 2043
rect 6696 1767 6703 2036
rect 6736 1967 6743 2233
rect 6756 2167 6763 2263
rect 6756 2127 6763 2153
rect 6776 2047 6783 2473
rect 6796 2027 6803 2523
rect 6816 2507 6823 2573
rect 6816 2267 6823 2313
rect 6816 2076 6823 2253
rect 6836 2107 6843 2973
rect 6876 2847 6883 3023
rect 6916 2987 6923 3036
rect 6876 2727 6883 2793
rect 6936 2756 6943 3273
rect 7096 3243 7103 3613
rect 7076 3236 7103 3243
rect 6956 2727 6963 2743
rect 6856 2367 6863 2713
rect 6856 2076 6863 2273
rect 6876 2187 6883 2713
rect 6916 2547 6923 2653
rect 6936 2303 6943 2573
rect 6956 2556 6963 2633
rect 6996 2587 7003 2733
rect 7016 2707 7023 3223
rect 7056 3207 7063 3223
rect 7036 3036 7043 3073
rect 7116 3023 7123 3033
rect 7096 3016 7123 3023
rect 7096 2567 7103 2993
rect 7116 2967 7123 3016
rect 7116 2767 7123 2833
rect 7136 2807 7143 4013
rect 7156 3787 7163 4693
rect 7176 4647 7183 4683
rect 7196 4507 7203 4973
rect 7256 4907 7263 5373
rect 7276 5147 7283 5473
rect 7316 5387 7323 6333
rect 7356 5967 7363 6213
rect 7396 6143 7403 6776
rect 7416 6227 7423 6633
rect 7436 6467 7443 7413
rect 7456 7007 7463 7053
rect 7476 6967 7483 7293
rect 7496 7127 7503 7613
rect 7516 7243 7523 7793
rect 7616 7647 7623 8473
rect 7636 8167 7643 8503
rect 7676 8496 7703 8503
rect 7656 8316 7663 8373
rect 7636 7887 7643 8133
rect 7576 7543 7583 7633
rect 7656 7607 7663 8153
rect 7616 7556 7623 7593
rect 7676 7567 7683 8473
rect 7716 8387 7723 8893
rect 7756 8796 7763 9013
rect 7796 8823 7803 10693
rect 7816 10427 7823 10693
rect 7816 9723 7823 10253
rect 7836 10047 7843 10493
rect 7916 10487 7923 10736
rect 7936 10507 7943 11053
rect 7956 10867 7963 10923
rect 7956 10827 7963 10853
rect 7976 10603 7983 11156
rect 8096 11127 8103 11183
rect 8056 10716 8063 10733
rect 8036 10687 8043 10703
rect 7976 10596 8003 10603
rect 7896 10436 7903 10453
rect 7956 10427 7963 10513
rect 7876 10407 7883 10423
rect 7936 10407 7943 10413
rect 7976 10407 7983 10453
rect 7876 10256 7883 10273
rect 7836 9947 7843 9963
rect 7876 9956 7883 10053
rect 7916 9943 7923 10273
rect 7836 9927 7843 9933
rect 7836 9747 7843 9913
rect 7856 9847 7863 9943
rect 7896 9936 7923 9943
rect 7916 9787 7923 9936
rect 7936 9847 7943 10233
rect 7956 9983 7963 10313
rect 7996 10287 8003 10596
rect 8136 10507 8143 11183
rect 8196 10916 8203 11133
rect 8216 10823 8223 10903
rect 8236 10847 8243 10923
rect 8256 10907 8263 11273
rect 8196 10816 8223 10823
rect 8196 10707 8203 10816
rect 8276 10716 8283 11653
rect 8296 11487 8303 11663
rect 8356 11416 8363 11733
rect 8476 11703 8483 11843
rect 8596 11827 8603 11863
rect 8656 11856 8683 11863
rect 8456 11696 8483 11703
rect 8496 11696 8503 11733
rect 8696 11727 8703 11893
rect 8816 11807 8823 11863
rect 8016 10387 8023 10473
rect 8036 10427 8043 10433
rect 8056 10247 8063 10493
rect 8156 10443 8163 10533
rect 8136 10436 8163 10443
rect 8076 10327 8083 10423
rect 8136 10367 8143 10436
rect 7976 10007 7983 10213
rect 8016 10187 8023 10193
rect 8056 10167 8063 10203
rect 7956 9976 7983 9983
rect 7816 9716 7843 9723
rect 7816 9107 7823 9153
rect 7816 8907 7823 8983
rect 7836 8967 7843 9716
rect 7856 9607 7863 9773
rect 7936 9756 7943 9833
rect 7976 9783 7983 9976
rect 8016 9976 8023 10013
rect 7996 9907 8003 9973
rect 8036 9947 8043 9963
rect 8076 9907 8083 9993
rect 8096 9807 8103 10033
rect 8116 9847 8123 10033
rect 7976 9776 8003 9783
rect 8096 9776 8103 9793
rect 7916 9707 7923 9743
rect 7856 9467 7863 9593
rect 7956 9463 7963 9773
rect 7936 9456 7963 9463
rect 7896 9276 7913 9283
rect 7856 8987 7863 9233
rect 7876 9227 7883 9263
rect 7876 8927 7883 9133
rect 7776 8816 7803 8823
rect 7736 8467 7743 8773
rect 7756 8467 7763 8533
rect 7776 8487 7783 8816
rect 7796 8527 7803 8783
rect 7796 8496 7823 8503
rect 7736 8327 7743 8433
rect 7696 8316 7723 8323
rect 7716 8247 7723 8316
rect 7716 8147 7723 8233
rect 7736 8187 7743 8293
rect 7716 8027 7723 8133
rect 7756 8107 7763 8433
rect 7756 8087 7763 8093
rect 7736 8036 7743 8053
rect 7696 7987 7703 8013
rect 7696 7836 7703 7973
rect 7756 7947 7763 8023
rect 7716 7867 7723 7913
rect 7576 7536 7603 7543
rect 7556 7356 7563 7453
rect 7596 7356 7603 7373
rect 7576 7307 7583 7333
rect 7516 7236 7543 7243
rect 7496 7096 7503 7113
rect 7516 7087 7523 7213
rect 7536 6947 7543 7236
rect 7496 6896 7503 6913
rect 7456 6847 7463 6873
rect 7536 6867 7543 6893
rect 7556 6887 7563 7093
rect 7576 7027 7583 7073
rect 7476 6856 7503 6863
rect 7496 6847 7503 6856
rect 7556 6847 7563 6853
rect 7456 6596 7463 6633
rect 7496 6596 7503 6613
rect 7536 6583 7543 6693
rect 7516 6576 7543 6583
rect 7476 6547 7483 6563
rect 7556 6547 7563 6813
rect 7576 6687 7583 6973
rect 7596 6827 7603 7313
rect 7616 6823 7623 7413
rect 7636 7327 7643 7543
rect 7656 7467 7663 7563
rect 7716 7427 7723 7813
rect 7756 7803 7763 7933
rect 7776 7847 7783 8373
rect 7796 8287 7803 8496
rect 7876 8487 7883 8893
rect 7816 8367 7823 8453
rect 7876 8447 7883 8473
rect 7896 8467 7903 9193
rect 7916 8987 7923 9193
rect 7936 9067 7943 9413
rect 7956 9247 7963 9433
rect 7976 9047 7983 9733
rect 7996 9447 8003 9776
rect 8056 9756 8073 9763
rect 8056 9687 8063 9756
rect 8116 9756 8123 9833
rect 7996 9107 8003 9293
rect 8016 9047 8023 9573
rect 8136 9527 8143 10233
rect 8036 9367 8043 9473
rect 7936 8983 7943 8993
rect 7996 8987 8003 9023
rect 8036 9007 8043 9313
rect 8056 9307 8063 9433
rect 8096 9407 8103 9463
rect 8096 9296 8103 9313
rect 8076 9287 8083 9293
rect 8136 9283 8143 9493
rect 8116 9276 8143 9283
rect 7936 8976 7963 8983
rect 7936 8803 7943 8913
rect 7916 8796 7943 8803
rect 7916 8687 7923 8796
rect 7896 8407 7903 8433
rect 7816 8303 7823 8313
rect 7816 8296 7843 8303
rect 7736 7796 7763 7803
rect 7656 7087 7663 7373
rect 7676 7147 7683 7393
rect 7736 7387 7743 7796
rect 7796 7787 7803 8173
rect 7816 7807 7823 8296
rect 7856 8276 7863 8353
rect 7916 8083 7923 8593
rect 7936 8107 7943 8513
rect 7956 8407 7963 8976
rect 7996 8763 8003 8873
rect 7976 8756 8003 8763
rect 7976 8507 7983 8756
rect 8016 8687 8023 9003
rect 8016 8547 8023 8673
rect 8016 8516 8043 8523
rect 8036 8487 8043 8516
rect 7987 8476 8003 8483
rect 7916 8076 7943 8083
rect 7836 7987 7843 8073
rect 7776 7367 7783 7653
rect 7836 7587 7843 7913
rect 7856 7547 7863 8053
rect 7936 8023 7943 8076
rect 7956 8047 7963 8333
rect 7916 8016 7943 8023
rect 7876 7947 7883 8013
rect 7936 8007 7943 8016
rect 7896 7987 7903 8003
rect 7936 7836 7943 7973
rect 7956 7827 7963 7933
rect 7796 7527 7803 7543
rect 7816 7516 7843 7523
rect 7696 7356 7723 7363
rect 7696 7347 7703 7356
rect 7736 7207 7743 7343
rect 7696 7076 7703 7093
rect 7636 7007 7643 7063
rect 7676 6867 7683 7063
rect 7696 6947 7703 6993
rect 7696 6856 7703 6933
rect 7716 6887 7723 7063
rect 7616 6816 7643 6823
rect 7456 6443 7463 6473
rect 7436 6436 7463 6443
rect 7416 6147 7423 6193
rect 7436 6187 7443 6436
rect 7456 6267 7463 6393
rect 7476 6347 7483 6453
rect 7576 6447 7583 6593
rect 7376 6136 7403 6143
rect 7336 5887 7343 5903
rect 7356 5443 7363 5693
rect 7376 5667 7383 6136
rect 7416 6123 7423 6133
rect 7396 6116 7423 6123
rect 7396 5707 7403 5953
rect 7476 5943 7483 6133
rect 7496 5987 7503 6173
rect 7516 6107 7523 6133
rect 7516 5943 7523 5993
rect 7456 5936 7483 5943
rect 7496 5936 7523 5943
rect 7436 5907 7443 5933
rect 7456 5887 7463 5936
rect 7536 5916 7543 6153
rect 7476 5887 7483 5903
rect 7436 5636 7443 5713
rect 7356 5436 7383 5443
rect 7336 5247 7343 5433
rect 7376 5416 7383 5436
rect 7396 5387 7403 5403
rect 7376 5227 7383 5353
rect 7336 5176 7343 5213
rect 7316 4983 7323 5163
rect 7376 5156 7383 5213
rect 7296 4976 7323 4983
rect 7356 4607 7363 4643
rect 7256 4476 7263 4533
rect 7216 4187 7223 4473
rect 7316 4467 7323 4533
rect 7376 4467 7383 4953
rect 7416 4927 7423 5623
rect 7436 5027 7443 5553
rect 7456 5147 7463 5163
rect 7456 4987 7463 5133
rect 7476 5007 7483 5713
rect 7496 5367 7503 5853
rect 7516 5567 7523 5873
rect 7576 5867 7583 6433
rect 7596 6367 7603 6633
rect 7616 6627 7623 6673
rect 7616 6387 7623 6593
rect 7636 6387 7643 6816
rect 7696 6616 7703 6813
rect 7716 6767 7723 6853
rect 7736 6583 7743 6853
rect 7756 6707 7763 7313
rect 7656 6443 7663 6583
rect 7716 6576 7743 6583
rect 7656 6436 7683 6443
rect 7556 5587 7563 5653
rect 7516 5387 7523 5433
rect 7536 5416 7543 5493
rect 7596 5447 7603 5623
rect 7636 5287 7643 5973
rect 7656 5903 7663 6413
rect 7676 6167 7683 6436
rect 7696 6396 7703 6433
rect 7716 6416 7723 6433
rect 7736 6396 7743 6413
rect 7676 5936 7683 6113
rect 7716 6107 7723 6373
rect 7656 5896 7683 5903
rect 7636 5107 7643 5123
rect 7496 4956 7503 5073
rect 7516 4947 7523 4993
rect 7427 4816 7433 4823
rect 7456 4683 7463 4813
rect 7536 4767 7543 4943
rect 7456 4676 7483 4683
rect 7276 4447 7283 4463
rect 7436 4463 7443 4573
rect 7476 4496 7483 4653
rect 7436 4456 7463 4463
rect 7216 4087 7223 4153
rect 7216 3996 7223 4073
rect 7236 4016 7243 4113
rect 7256 4007 7263 4163
rect 7396 4003 7403 4373
rect 7456 4167 7463 4353
rect 7436 4007 7443 4153
rect 7476 4087 7483 4183
rect 7516 4163 7523 4213
rect 7496 4156 7523 4163
rect 7376 3996 7403 4003
rect 7156 3227 7163 3413
rect 7176 2887 7183 3953
rect 7216 3523 7223 3873
rect 7376 3727 7383 3996
rect 7196 3516 7223 3523
rect 7236 3516 7263 3523
rect 7196 3007 7203 3516
rect 7236 3267 7243 3516
rect 7276 3467 7283 3703
rect 7476 3703 7483 3933
rect 7556 3747 7563 5053
rect 7656 5047 7663 5553
rect 7676 5387 7683 5896
rect 7696 5647 7703 5903
rect 7716 5263 7723 5933
rect 7736 5567 7743 6353
rect 7756 5547 7763 6653
rect 7776 6167 7783 7173
rect 7796 7027 7803 7473
rect 7836 7407 7843 7516
rect 7856 7427 7863 7533
rect 7796 6407 7803 6873
rect 7816 6487 7823 7033
rect 7836 6987 7843 7353
rect 7856 6967 7863 7353
rect 7876 7267 7883 7633
rect 7896 7327 7903 7373
rect 7916 7356 7923 7793
rect 7976 7787 7983 8453
rect 7956 7487 7963 7773
rect 7996 7687 8003 8453
rect 8016 7587 8023 8213
rect 7976 7527 7983 7543
rect 8036 7523 8043 8453
rect 8056 8323 8063 9033
rect 8076 8347 8083 9013
rect 8096 8343 8103 8993
rect 8136 8967 8143 9276
rect 8156 9027 8163 10373
rect 8176 10227 8183 10473
rect 8196 10267 8203 10433
rect 8216 10427 8223 10703
rect 8296 10647 8303 11393
rect 8336 11347 8343 11403
rect 8436 11327 8443 11693
rect 8456 11507 8463 11696
rect 8536 11527 8543 11713
rect 8516 11396 8523 11513
rect 8576 11447 8583 11673
rect 8596 11647 8603 11693
rect 8696 11676 8703 11713
rect 8636 11607 8643 11663
rect 8576 11383 8583 11433
rect 8496 11287 8503 11383
rect 8536 11376 8583 11383
rect 8316 11196 8323 11273
rect 8356 11196 8363 11233
rect 8556 11227 8563 11253
rect 8396 11196 8403 11213
rect 8376 11123 8383 11183
rect 8356 11116 8383 11123
rect 8176 9267 8183 10213
rect 8216 9967 8223 10193
rect 8256 9947 8263 10493
rect 8276 10436 8283 10453
rect 8296 10407 8303 10423
rect 8196 9587 8203 9943
rect 8216 9887 8223 9923
rect 8276 9887 8283 9993
rect 8296 9867 8303 10073
rect 8176 8996 8183 9233
rect 8156 8907 8163 8983
rect 8136 8767 8143 8783
rect 8136 8747 8143 8753
rect 8156 8567 8163 8773
rect 8176 8647 8183 8953
rect 8196 8607 8203 9513
rect 8216 9467 8223 9713
rect 8256 9447 8263 9723
rect 8296 9707 8303 9723
rect 8316 9527 8323 10713
rect 8336 10436 8343 10573
rect 8356 10487 8363 11116
rect 8376 10527 8383 11093
rect 8396 10787 8403 10903
rect 8436 10803 8443 10903
rect 8456 10827 8463 11213
rect 8496 11107 8503 11193
rect 8536 11156 8543 11193
rect 8556 11176 8563 11213
rect 8596 11163 8603 11253
rect 8576 11156 8603 11163
rect 8596 10903 8603 10933
rect 8576 10896 8603 10903
rect 8436 10796 8463 10803
rect 8396 10736 8423 10743
rect 8336 9507 8343 10393
rect 8356 9847 8363 10423
rect 8376 10407 8383 10453
rect 8376 10216 8383 10393
rect 8396 10307 8403 10736
rect 8436 10687 8443 10703
rect 8456 10547 8463 10796
rect 8436 10236 8463 10243
rect 8416 10147 8423 10223
rect 8456 10207 8463 10236
rect 8456 10047 8463 10193
rect 8236 9263 8243 9273
rect 8236 9256 8263 9263
rect 8296 9067 8303 9453
rect 8316 9447 8323 9463
rect 8316 9427 8323 9433
rect 8216 8767 8223 8983
rect 8236 8787 8243 8813
rect 8136 8507 8143 8553
rect 8196 8487 8203 8523
rect 8236 8467 8243 8653
rect 8096 8336 8123 8343
rect 8056 8316 8083 8323
rect 8116 8316 8123 8336
rect 8096 8067 8103 8293
rect 8056 7836 8063 7933
rect 8096 7927 8103 8023
rect 8136 8007 8143 8023
rect 8076 7807 8083 7823
rect 8076 7747 8083 7773
rect 8056 7547 8063 7733
rect 7996 7503 8003 7523
rect 7976 7496 8003 7503
rect 8016 7516 8043 7523
rect 7876 7027 7883 7083
rect 7856 6856 7863 6933
rect 7896 6887 7903 6893
rect 7896 6856 7903 6873
rect 7876 6836 7883 6853
rect 7876 6616 7883 6713
rect 7936 6667 7943 7013
rect 7896 6587 7903 6603
rect 7916 6487 7923 6623
rect 7956 6587 7963 7313
rect 7796 6116 7803 6393
rect 7836 6347 7843 6473
rect 7856 6363 7863 6433
rect 7896 6376 7903 6393
rect 7936 6363 7943 6413
rect 7856 6356 7883 6363
rect 7916 6356 7943 6363
rect 7836 6116 7843 6333
rect 7976 6247 7983 7496
rect 7996 7167 8003 7453
rect 7996 6987 8003 7153
rect 7996 6607 8003 6953
rect 8016 6847 8023 7516
rect 8096 7407 8103 7593
rect 8116 7467 8123 7753
rect 8136 7707 8143 7833
rect 8156 7603 8163 8093
rect 8176 7627 8183 8333
rect 8196 8027 8203 8453
rect 8256 8363 8263 8893
rect 8276 8487 8283 8813
rect 8296 8796 8303 8953
rect 8316 8907 8323 9393
rect 8336 8967 8343 9413
rect 8356 9407 8363 9833
rect 8376 9747 8383 9963
rect 8436 9736 8443 9753
rect 8416 9667 8423 9723
rect 8376 9227 8383 9513
rect 8396 9256 8403 9553
rect 8436 9483 8443 9593
rect 8456 9507 8463 9723
rect 8436 9476 8463 9483
rect 8416 9407 8423 9473
rect 8436 9327 8443 9443
rect 8476 9427 8483 10133
rect 8496 9987 8503 10793
rect 8616 10787 8623 10903
rect 8596 10696 8603 10733
rect 8576 10547 8583 10683
rect 8616 10663 8623 10683
rect 8596 10656 8623 10663
rect 8516 10427 8523 10443
rect 8536 10367 8543 10423
rect 8576 10407 8583 10423
rect 8596 10387 8603 10656
rect 8656 10483 8663 11633
rect 8676 10527 8683 11663
rect 8716 11607 8723 11733
rect 8836 11656 8843 11833
rect 8916 11643 8923 11813
rect 8896 11636 8923 11643
rect 8716 11267 8723 11383
rect 8736 11327 8743 11363
rect 8756 11327 8763 11383
rect 8816 11267 8823 11633
rect 8936 11587 8943 11853
rect 8996 11647 9003 11833
rect 9016 11687 9023 11863
rect 9176 11807 9183 11883
rect 9196 11847 9203 11903
rect 9496 11896 9503 12013
rect 8856 11416 8883 11423
rect 8856 11307 8863 11416
rect 8716 11196 8723 11213
rect 8696 10747 8703 11153
rect 8716 10747 8723 10913
rect 8736 10887 8743 10903
rect 8796 10747 8803 10923
rect 8716 10687 8723 10733
rect 8816 10716 8823 11253
rect 8636 10476 8663 10483
rect 8636 10307 8643 10476
rect 8676 10456 8703 10463
rect 8736 10456 8743 10653
rect 8756 10507 8763 10703
rect 8516 9467 8523 10293
rect 8656 10267 8663 10453
rect 8676 10407 8683 10456
rect 8716 10427 8723 10443
rect 8596 10236 8603 10253
rect 8676 10247 8683 10393
rect 8556 9707 8563 10233
rect 8616 10087 8623 10223
rect 8556 9463 8563 9693
rect 8536 9456 8563 9463
rect 8416 9236 8423 9253
rect 8456 9207 8463 9243
rect 8376 8867 8383 8983
rect 8396 8807 8403 9153
rect 8436 9087 8443 9153
rect 8456 8963 8463 9073
rect 8476 8987 8483 9353
rect 8436 8956 8463 8963
rect 8336 8796 8363 8803
rect 8356 8607 8363 8796
rect 8236 8356 8263 8363
rect 8236 8316 8243 8356
rect 8276 8316 8303 8323
rect 8296 8287 8303 8316
rect 8216 8007 8223 8093
rect 8196 7807 8203 7993
rect 8236 7607 8243 8253
rect 8316 8087 8323 8593
rect 8276 7863 8283 8013
rect 8296 7947 8303 8003
rect 8316 7887 8323 8023
rect 8276 7856 8303 7863
rect 8136 7596 8163 7603
rect 8056 7376 8083 7383
rect 8056 7347 8063 7376
rect 8116 7343 8123 7433
rect 8096 7336 8123 7343
rect 8036 7067 8043 7313
rect 8136 7147 8143 7596
rect 8156 7227 8163 7573
rect 8196 7267 8203 7543
rect 8156 7096 8163 7113
rect 8176 7087 8183 7173
rect 8076 6876 8083 6913
rect 8116 6876 8143 6883
rect 8136 6847 8143 6876
rect 8047 6716 8053 6723
rect 7776 5487 7783 6093
rect 7856 6047 7863 6103
rect 7876 5947 7883 6153
rect 7896 6087 7903 6153
rect 7976 6107 7983 6133
rect 7836 5916 7843 5933
rect 7916 5916 7943 5923
rect 7816 5467 7823 5603
rect 7836 5587 7843 5623
rect 7776 5436 7783 5453
rect 7796 5407 7803 5453
rect 7816 5427 7823 5453
rect 7716 5256 7743 5263
rect 7736 5087 7743 5256
rect 7576 4676 7583 5013
rect 7616 4943 7623 4973
rect 7616 4936 7643 4943
rect 7636 4647 7643 4936
rect 7816 4787 7823 5373
rect 7836 5067 7843 5533
rect 7856 5267 7863 5853
rect 7856 5156 7863 5253
rect 7876 5067 7883 5873
rect 7896 5847 7903 5903
rect 7936 5527 7943 5916
rect 7996 5887 8003 6573
rect 8036 6423 8043 6593
rect 8076 6427 8083 6563
rect 8036 6416 8063 6423
rect 8076 6396 8103 6403
rect 8096 6367 8103 6396
rect 8076 6116 8083 6173
rect 8096 6087 8103 6153
rect 8116 5987 8123 6613
rect 8176 6607 8183 7053
rect 8196 6727 8203 7083
rect 8096 5936 8123 5943
rect 8056 5727 8063 5913
rect 8116 5903 8123 5936
rect 7976 5656 7983 5693
rect 8076 5667 8083 5903
rect 8116 5896 8143 5903
rect 8156 5767 8163 6573
rect 8196 6187 8203 6593
rect 8216 6467 8223 7433
rect 8256 7367 8263 7593
rect 8276 7447 8283 7553
rect 8236 7287 8243 7323
rect 8276 7307 8283 7323
rect 8256 6876 8263 6933
rect 8296 6847 8303 7813
rect 8336 7787 8343 8353
rect 8356 7847 8363 8533
rect 8376 8516 8383 8633
rect 8376 7827 8383 8333
rect 8396 8327 8403 8473
rect 8416 8447 8423 8953
rect 8436 8423 8443 8956
rect 8496 8923 8503 9413
rect 8516 8947 8523 9453
rect 8536 9007 8543 9456
rect 8576 9247 8583 10053
rect 8656 9927 8663 9943
rect 8596 9756 8603 9853
rect 8696 9807 8703 10313
rect 8616 9776 8623 9793
rect 8656 9447 8663 9753
rect 8676 9467 8683 9773
rect 8596 9436 8623 9443
rect 8596 9276 8603 9436
rect 8636 9347 8643 9433
rect 8556 9016 8563 9133
rect 8576 8987 8583 9003
rect 8496 8916 8523 8923
rect 8476 8816 8493 8823
rect 8456 8796 8463 8813
rect 8476 8507 8483 8533
rect 8416 8416 8443 8423
rect 8416 8267 8423 8416
rect 8476 8276 8483 8393
rect 8496 8323 8503 8653
rect 8516 8567 8523 8916
rect 8536 8667 8543 8813
rect 8556 8567 8563 8813
rect 8596 8727 8603 9023
rect 8636 9003 8643 9243
rect 8616 8996 8643 9003
rect 8636 8807 8643 8996
rect 8656 8887 8663 9073
rect 8676 8987 8683 9293
rect 8696 9087 8703 9733
rect 8716 9183 8723 10373
rect 8756 10307 8763 10493
rect 8736 10236 8763 10243
rect 8736 10127 8743 10236
rect 8776 10187 8783 10413
rect 8796 10267 8803 10703
rect 8816 10347 8823 10473
rect 8836 10283 8843 11153
rect 8856 10947 8863 11293
rect 8896 11176 8923 11183
rect 8956 11176 8963 11193
rect 8896 11107 8903 11176
rect 8996 11163 9003 11293
rect 8976 11156 9003 11163
rect 8936 11007 8943 11113
rect 8936 10927 8943 10993
rect 9016 10987 9023 11413
rect 8956 10936 8963 10953
rect 8996 10907 9003 10943
rect 9036 10927 9043 11733
rect 9216 11707 9223 11883
rect 9436 11876 9443 11893
rect 10036 11883 10043 12013
rect 10556 11896 10563 11913
rect 9076 11416 9083 11473
rect 9156 11447 9163 11633
rect 8856 10567 8863 10733
rect 8876 10487 8883 10773
rect 8896 10707 8903 10773
rect 8896 10463 8903 10693
rect 8916 10483 8923 10753
rect 8936 10723 8943 10813
rect 9016 10767 9023 10923
rect 8936 10716 8963 10723
rect 8936 10683 8943 10716
rect 9016 10696 9023 10733
rect 8936 10676 8963 10683
rect 8916 10476 8943 10483
rect 8896 10456 8923 10463
rect 8816 10276 8843 10283
rect 8736 9947 8743 10113
rect 8816 10007 8823 10276
rect 8776 9927 8783 9943
rect 8736 9627 8743 9913
rect 8796 9776 8803 9793
rect 8816 9787 8823 9943
rect 8836 9927 8843 10253
rect 8716 9176 8743 9183
rect 8656 8827 8663 8873
rect 8516 8507 8523 8553
rect 8576 8527 8583 8543
rect 8596 8467 8603 8523
rect 8496 8316 8523 8323
rect 8416 8187 8423 8193
rect 8396 7947 8403 8073
rect 8416 8027 8423 8173
rect 8456 8056 8463 8073
rect 8496 8056 8503 8073
rect 8436 7807 8443 8033
rect 8476 8023 8483 8043
rect 8476 8016 8503 8023
rect 8476 7827 8483 7873
rect 8496 7836 8503 8016
rect 8516 7887 8523 8316
rect 8536 8307 8543 8453
rect 8336 7523 8343 7613
rect 8376 7567 8383 7573
rect 8416 7523 8423 7563
rect 8336 7516 8423 7523
rect 8316 7307 8323 7373
rect 8436 7356 8443 7693
rect 8456 7447 8463 7823
rect 8536 7723 8543 8053
rect 8556 7907 8563 8353
rect 8576 8087 8583 8453
rect 8616 8367 8623 8753
rect 8636 8667 8643 8763
rect 8676 8647 8683 8763
rect 8696 8503 8703 9053
rect 8716 8907 8723 9073
rect 8736 8767 8743 9176
rect 8756 9027 8763 9773
rect 8776 9476 8783 9693
rect 8816 9507 8823 9513
rect 8776 8996 8783 9433
rect 8796 9427 8803 9463
rect 8816 9283 8823 9493
rect 8836 9476 8843 9853
rect 8856 9747 8863 10253
rect 8876 10187 8883 10403
rect 8916 10263 8923 10456
rect 8936 10436 8943 10476
rect 8956 10427 8963 10676
rect 8896 10256 8923 10263
rect 8856 9507 8863 9653
rect 8876 9607 8883 9713
rect 8816 9276 8843 9283
rect 8836 9256 8843 9276
rect 8796 9236 8823 9243
rect 8856 9236 8863 9433
rect 8736 8516 8743 8553
rect 8756 8547 8763 8973
rect 8796 8967 8803 9236
rect 8836 8996 8843 9213
rect 8856 8827 8863 9013
rect 8876 8967 8883 9193
rect 8896 9043 8903 10256
rect 8956 10236 8963 10253
rect 8916 10223 8923 10233
rect 8916 10216 8943 10223
rect 8976 9807 8983 10533
rect 9016 10236 9023 10273
rect 9036 10167 9043 10913
rect 9056 10587 9063 11413
rect 9096 11387 9103 11403
rect 9116 11287 9123 11423
rect 9156 11403 9163 11413
rect 9136 11396 9163 11403
rect 9136 11196 9143 11373
rect 9176 10967 9183 11673
rect 9236 11643 9243 11853
rect 9416 11847 9423 11863
rect 9316 11656 9323 11773
rect 9336 11647 9343 11753
rect 9236 11636 9263 11643
rect 9316 11487 9323 11613
rect 9256 11416 9283 11423
rect 9256 11387 9263 11416
rect 9196 11227 9203 11353
rect 9196 11196 9203 11213
rect 9116 10903 9123 10933
rect 9116 10896 9143 10903
rect 9136 10683 9143 10713
rect 9176 10696 9183 10713
rect 9136 10676 9163 10683
rect 8996 9887 9003 9943
rect 8996 9787 9003 9873
rect 9036 9807 9043 10153
rect 9056 10127 9063 10513
rect 9096 10423 9103 10473
rect 9076 10416 9103 10423
rect 9116 10407 9123 10423
rect 9136 10367 9143 10393
rect 8916 9227 8923 9613
rect 8936 9427 8943 9453
rect 8936 9187 8943 9413
rect 8956 9267 8963 9773
rect 9036 9756 9043 9773
rect 9016 9727 9023 9743
rect 9076 9667 9083 9973
rect 9116 9707 9123 10273
rect 9176 10263 9183 10493
rect 9196 10387 9203 10683
rect 9196 10327 9203 10373
rect 9176 10256 9203 10263
rect 9136 10236 9163 10243
rect 9196 10236 9203 10256
rect 9216 10247 9223 10313
rect 9136 10207 9143 10236
rect 9136 10087 9143 10193
rect 9176 10147 9183 10223
rect 9216 10216 9223 10233
rect 9236 10067 9243 10813
rect 9316 10456 9323 10693
rect 9336 10467 9343 11613
rect 9376 11387 9383 11413
rect 9396 11047 9403 11753
rect 9356 10787 9363 10883
rect 9396 10743 9403 10953
rect 9416 10867 9423 11773
rect 9536 11767 9543 11873
rect 9836 11787 9843 11883
rect 9916 11876 9943 11883
rect 10016 11876 10043 11883
rect 9636 11696 9643 11753
rect 9816 11696 9863 11703
rect 9596 11676 9623 11683
rect 9656 11676 9683 11683
rect 9436 11567 9443 11653
rect 9496 11627 9503 11643
rect 9436 11207 9443 11383
rect 9596 11367 9603 11676
rect 9676 11667 9683 11676
rect 9696 11607 9703 11653
rect 9856 11627 9863 11696
rect 9876 11687 9883 11813
rect 9656 11416 9683 11423
rect 9376 10736 9403 10743
rect 9256 10227 9263 10433
rect 9276 10427 9283 10453
rect 9336 10447 9343 10453
rect 9296 10407 9303 10443
rect 9436 10347 9443 10673
rect 9456 10527 9463 11313
rect 9596 11307 9603 11353
rect 9556 11187 9563 11213
rect 9496 11176 9523 11183
rect 9356 10236 9383 10243
rect 9436 10236 9443 10333
rect 9356 10183 9363 10236
rect 9416 10203 9423 10213
rect 9456 10207 9463 10253
rect 9396 10196 9423 10203
rect 9356 10176 9383 10183
rect 9196 9976 9203 10013
rect 9176 9907 9183 9963
rect 8996 9496 9003 9613
rect 9036 9496 9063 9503
rect 9056 9387 9063 9496
rect 9076 9447 9083 9653
rect 9116 9527 9123 9573
rect 8976 9207 8983 9273
rect 9016 9267 9023 9293
rect 9076 9276 9103 9283
rect 8896 9036 8923 9043
rect 8896 8947 8903 9013
rect 8776 8507 8783 8523
rect 8696 8496 8723 8503
rect 8696 8347 8703 8496
rect 8576 7987 8583 8053
rect 8596 8023 8603 8333
rect 8696 8316 8703 8333
rect 8616 8296 8643 8303
rect 8616 8287 8623 8296
rect 8616 8247 8623 8273
rect 8676 8023 8683 8303
rect 8596 8016 8623 8023
rect 8656 8016 8683 8023
rect 8636 7907 8643 8003
rect 8676 7927 8683 8016
rect 8696 7887 8703 8093
rect 8716 7887 8723 8073
rect 8516 7716 8543 7723
rect 8516 7567 8523 7716
rect 8616 7667 8623 7853
rect 8576 7567 8583 7583
rect 8616 7576 8623 7593
rect 8596 7547 8603 7563
rect 8636 7547 8643 7873
rect 8476 7356 8483 7373
rect 8496 7307 8503 7533
rect 8656 7527 8663 7853
rect 8676 7567 8683 7613
rect 8316 6967 8323 7043
rect 8476 7027 8483 7253
rect 8516 7083 8523 7493
rect 8496 7076 8523 7083
rect 8316 6887 8323 6933
rect 8256 6616 8263 6773
rect 8296 6616 8303 6833
rect 8336 6807 8343 6873
rect 8256 6376 8263 6413
rect 8316 6383 8323 6593
rect 8296 6376 8323 6383
rect 8216 6147 8223 6373
rect 8276 6356 8283 6373
rect 8216 6116 8223 6133
rect 8176 5747 8183 5933
rect 8196 5867 8203 6083
rect 8236 5903 8243 6113
rect 8216 5896 8243 5903
rect 8016 5656 8043 5663
rect 8036 5607 8043 5656
rect 8076 5627 8083 5653
rect 8176 5636 8183 5653
rect 8196 5607 8203 5623
rect 8116 5456 8123 5493
rect 7936 5436 7943 5453
rect 8087 5436 8103 5443
rect 7916 5416 7923 5433
rect 8076 5387 8083 5433
rect 7896 5223 7903 5293
rect 8196 5287 8203 5593
rect 8216 5407 8223 5833
rect 8236 5803 8243 5896
rect 8256 5847 8263 6133
rect 8276 6116 8283 6153
rect 8336 6007 8343 6533
rect 8376 6487 8383 6973
rect 8436 6883 8443 6913
rect 8416 6876 8443 6883
rect 8416 6787 8423 6876
rect 8456 6587 8463 6993
rect 8536 6927 8543 7433
rect 8376 6167 8383 6473
rect 8396 6463 8403 6533
rect 8416 6487 8423 6563
rect 8396 6456 8423 6463
rect 8416 6396 8423 6456
rect 8456 6407 8463 6553
rect 8516 6227 8523 6853
rect 8536 6127 8543 6413
rect 8556 6327 8563 7513
rect 8616 7367 8623 7473
rect 8676 7407 8683 7433
rect 8636 7207 8643 7343
rect 8596 6627 8603 7113
rect 8676 7047 8683 7353
rect 8696 7327 8703 7693
rect 8716 7507 8723 7593
rect 8736 7527 8743 8353
rect 8756 7767 8763 8503
rect 8776 8167 8783 8333
rect 8776 8107 8783 8153
rect 8776 8047 8783 8073
rect 8796 7607 8803 8713
rect 8816 8523 8823 8813
rect 8896 8796 8903 8933
rect 8876 8767 8883 8783
rect 8876 8527 8883 8753
rect 8816 8516 8843 8523
rect 8816 8087 8823 8493
rect 8836 8347 8843 8516
rect 8896 8367 8903 8533
rect 8896 8347 8903 8353
rect 8916 8347 8923 9036
rect 8936 8883 8943 9033
rect 9036 8987 9043 9213
rect 8936 8876 8963 8883
rect 8936 8847 8943 8853
rect 8936 8567 8943 8833
rect 8956 8807 8963 8876
rect 8976 8787 8983 8973
rect 9036 8823 9043 8913
rect 9056 8847 9063 9263
rect 9076 8987 9083 9013
rect 9096 8927 9103 9276
rect 9116 9247 9123 9433
rect 9016 8816 9043 8823
rect 9016 8796 9023 8816
rect 8996 8723 9003 8773
rect 9036 8747 9043 8783
rect 8996 8716 9023 8723
rect 9016 8587 9023 8716
rect 8876 8316 8903 8323
rect 8856 8067 8863 8213
rect 8896 8107 8903 8316
rect 8856 8036 8863 8053
rect 8896 8047 8903 8093
rect 8816 7927 8823 7953
rect 8816 7827 8823 7913
rect 8836 7767 8843 7833
rect 8776 7576 8783 7593
rect 8756 7547 8763 7573
rect 8816 7527 8823 7583
rect 8856 7563 8863 7913
rect 8876 7816 8883 7933
rect 8896 7867 8903 7973
rect 8916 7947 8923 8293
rect 8936 8267 8943 8513
rect 9016 8503 9023 8573
rect 8996 8496 9023 8503
rect 9016 8487 9023 8496
rect 8936 8007 8943 8013
rect 8936 7847 8943 7993
rect 8836 7556 8863 7563
rect 8716 7303 8723 7373
rect 8776 7356 8783 7493
rect 8816 7356 8823 7453
rect 8876 7407 8883 7753
rect 8896 7327 8903 7773
rect 8916 7547 8923 7653
rect 8696 7296 8723 7303
rect 8696 7067 8703 7296
rect 8756 7076 8763 7313
rect 8916 7127 8923 7533
rect 8936 7387 8943 7673
rect 8956 7507 8963 8313
rect 8996 8307 9003 8333
rect 9036 8327 9043 8553
rect 9056 8527 9063 8573
rect 9056 8363 9063 8513
rect 9076 8387 9083 8593
rect 9056 8356 9083 8363
rect 8976 7587 8983 7873
rect 8996 7667 9003 8253
rect 9016 8207 9023 8283
rect 9076 8207 9083 8356
rect 9056 8036 9063 8053
rect 8996 7576 9003 7653
rect 9016 7627 9023 8033
rect 9076 8007 9083 8023
rect 9036 7827 9043 7893
rect 9096 7867 9103 8833
rect 9116 8807 9123 9233
rect 9116 8543 9123 8633
rect 9136 8567 9143 9793
rect 9176 9736 9183 9773
rect 9196 9756 9203 9793
rect 9156 9527 9163 9733
rect 9216 9687 9223 9743
rect 9176 9496 9183 9533
rect 9196 9467 9203 9483
rect 9236 9447 9243 9483
rect 9196 9276 9203 9293
rect 9256 9283 9263 10153
rect 9336 10047 9343 10073
rect 9236 9276 9263 9283
rect 9216 9023 9223 9263
rect 9216 9016 9243 9023
rect 9156 8947 9163 9003
rect 9196 8996 9203 9013
rect 9176 8687 9183 8983
rect 9236 8823 9243 9016
rect 9256 8907 9263 9173
rect 9276 9147 9283 9953
rect 9296 9747 9303 10013
rect 9336 9943 9343 10033
rect 9376 9967 9383 10176
rect 9456 9987 9463 10113
rect 9316 9907 9323 9943
rect 9336 9936 9363 9943
rect 9296 9007 9303 9713
rect 9316 9367 9323 9893
rect 9356 9756 9363 9913
rect 9396 9756 9403 9773
rect 9416 9747 9423 9753
rect 9336 9467 9343 9733
rect 9376 9687 9383 9743
rect 9347 9456 9363 9463
rect 9416 9387 9423 9463
rect 9356 9227 9363 9373
rect 9436 9267 9443 9853
rect 9456 9367 9463 9693
rect 9376 9256 9403 9263
rect 9376 9067 9383 9256
rect 9456 9167 9463 9243
rect 9316 9016 9343 9023
rect 9216 8816 9243 8823
rect 9116 8536 9143 8543
rect 9136 8516 9143 8536
rect 9176 8507 9183 8523
rect 9116 8487 9123 8503
rect 9156 8467 9163 8503
rect 9216 8467 9223 8816
rect 9256 8796 9283 8803
rect 9256 8687 9263 8796
rect 9236 8443 9243 8473
rect 9216 8436 9243 8443
rect 9116 7907 9123 8373
rect 9176 8316 9203 8323
rect 9136 7867 9143 8193
rect 9176 8147 9183 8316
rect 9216 8283 9223 8436
rect 9256 8323 9263 8673
rect 9296 8403 9303 8973
rect 9316 8947 9323 9016
rect 9356 8907 9363 8993
rect 9316 8667 9323 8793
rect 9316 8536 9323 8653
rect 9356 8647 9363 8873
rect 9396 8796 9403 8933
rect 9376 8607 9383 8773
rect 9416 8767 9423 8783
rect 9376 8587 9383 8593
rect 9356 8536 9383 8543
rect 9296 8396 9323 8403
rect 9296 8367 9303 8373
rect 9236 8316 9263 8323
rect 9196 8276 9223 8283
rect 9176 8027 9183 8133
rect 9196 8007 9203 8276
rect 9256 8247 9263 8273
rect 9216 8027 9223 8043
rect 9256 8036 9263 8093
rect 9056 7836 9063 7853
rect 9096 7836 9143 7843
rect 9136 7707 9143 7836
rect 8896 7096 8923 7103
rect 8956 7096 8963 7343
rect 8676 6876 8683 6953
rect 8716 6876 8723 6993
rect 8736 6843 8743 7033
rect 8836 6896 8843 7073
rect 8876 6987 8883 7093
rect 8896 7087 8903 7096
rect 8856 6847 8863 6853
rect 8716 6836 8743 6843
rect 8716 6747 8723 6836
rect 8596 6416 8603 6493
rect 8616 6427 8623 6583
rect 8656 6547 8663 6583
rect 8676 6487 8683 6593
rect 8236 5796 8263 5803
rect 8236 5627 8243 5733
rect 7896 5216 7923 5223
rect 7916 5167 7923 5216
rect 7916 4936 7923 5153
rect 7936 5147 7943 5163
rect 7936 5007 7943 5133
rect 7976 4923 7983 5173
rect 8116 5087 8123 5123
rect 7956 4916 7983 4923
rect 7956 4727 7963 4916
rect 7656 4647 7663 4683
rect 7696 4567 7703 4573
rect 7836 4567 7843 4643
rect 7656 4476 7663 4493
rect 7696 4476 7703 4553
rect 7576 4003 7583 4473
rect 7616 4087 7623 4473
rect 7796 4467 7803 4553
rect 7856 4527 7863 4673
rect 7836 4476 7843 4513
rect 7656 4196 7663 4293
rect 7736 4196 7763 4203
rect 7736 4187 7743 4196
rect 7576 3996 7603 4003
rect 7576 3723 7583 3996
rect 7576 3716 7603 3723
rect 7456 3696 7483 3703
rect 7216 3187 7223 3233
rect 7116 2743 7123 2753
rect 7216 2747 7223 3073
rect 7256 3056 7263 3093
rect 7276 3083 7283 3223
rect 7296 3107 7303 3233
rect 7336 3167 7343 3693
rect 7416 3687 7423 3693
rect 7456 3647 7463 3696
rect 7616 3687 7623 3983
rect 7636 3967 7643 4183
rect 7656 3996 7663 4153
rect 7816 4007 7823 4463
rect 7836 4187 7843 4203
rect 7756 3787 7763 3973
rect 7796 3947 7803 3963
rect 7276 3076 7303 3083
rect 7276 3047 7283 3053
rect 7116 2736 7143 2743
rect 7016 2447 7023 2543
rect 7096 2387 7103 2553
rect 7156 2347 7163 2723
rect 7176 2556 7203 2563
rect 7176 2507 7183 2513
rect 6936 2296 6963 2303
rect 6956 2263 6963 2296
rect 6996 2267 7003 2293
rect 6936 2256 6963 2263
rect 6876 2056 6903 2063
rect 6736 1803 6743 1953
rect 6736 1796 6763 1803
rect 6836 1783 6843 2013
rect 6816 1776 6843 1783
rect 6676 1583 6683 1713
rect 6656 1576 6683 1583
rect 6656 1487 6663 1576
rect 6716 1567 6723 1583
rect 6596 1107 6603 1353
rect 6636 1316 6643 1333
rect 6636 1116 6643 1253
rect 6656 1247 6663 1283
rect 6696 1267 6703 1333
rect 6696 1163 6703 1253
rect 6676 1156 6703 1163
rect 6676 1116 6683 1156
rect 6696 1096 6703 1133
rect 6596 747 6603 823
rect 6616 616 6623 693
rect 6656 627 6663 753
rect 6736 647 6743 1493
rect 6756 1387 6763 1753
rect 6776 1347 6783 1593
rect 6816 1367 6823 1776
rect 6836 1567 6843 1613
rect 6756 1287 6763 1313
rect 6776 1296 6803 1303
rect 6776 1287 6783 1296
rect 6807 1276 6823 1283
rect 6576 187 6583 613
rect 6736 467 6743 613
rect 6696 356 6723 363
rect 6716 307 6723 356
rect 6516 156 6543 163
rect 6696 156 6723 163
rect 6736 156 6743 453
rect 6756 387 6763 1193
rect 6776 827 6783 1273
rect 6856 1207 6863 2033
rect 6896 1787 6903 2056
rect 6916 2047 6923 2073
rect 6936 1827 6943 2173
rect 6956 2147 6963 2256
rect 6956 1807 6963 2093
rect 6996 1867 7003 2113
rect 6936 1767 6943 1783
rect 6896 1616 6903 1633
rect 6876 1596 6883 1613
rect 6936 1603 6943 1753
rect 6976 1747 6983 1783
rect 6996 1727 7003 1803
rect 7016 1667 7023 2333
rect 7036 2247 7043 2313
rect 7096 2276 7103 2293
rect 7136 2276 7143 2313
rect 7156 2147 7163 2263
rect 7036 2056 7043 2113
rect 7096 2076 7123 2083
rect 7076 2047 7083 2063
rect 6927 1596 6943 1603
rect 6816 1087 6823 1153
rect 6876 1116 6883 1153
rect 6856 1087 6863 1103
rect 6896 1096 6903 1113
rect 6796 827 6803 843
rect 6836 836 6843 933
rect 6816 807 6823 823
rect 6856 807 6863 823
rect 6916 747 6923 1373
rect 6956 1307 6963 1653
rect 6996 1316 7003 1633
rect 7036 1596 7043 1813
rect 7076 1767 7083 2013
rect 7096 1807 7103 1853
rect 7116 1783 7123 2076
rect 7136 2027 7143 2073
rect 7176 2047 7183 2493
rect 7196 2247 7203 2556
rect 7236 2467 7243 2693
rect 7256 2547 7263 2713
rect 7276 2547 7283 2993
rect 7296 2567 7303 3076
rect 7336 2887 7343 3153
rect 7356 2767 7363 3293
rect 7376 3227 7383 3633
rect 7576 3536 7583 3673
rect 7676 3547 7683 3713
rect 7396 3496 7403 3513
rect 7696 3496 7723 3503
rect 7716 3367 7723 3496
rect 7396 3047 7403 3213
rect 7416 3187 7423 3223
rect 7396 3016 7403 3033
rect 7416 3007 7423 3053
rect 7436 3016 7443 3073
rect 7316 2747 7323 2763
rect 7336 2727 7343 2743
rect 7376 2727 7383 2743
rect 7216 2067 7223 2373
rect 7276 2347 7283 2533
rect 7376 2527 7383 2633
rect 7396 2536 7403 2753
rect 7416 2727 7423 2853
rect 7436 2727 7443 2893
rect 7516 2827 7523 2993
rect 7556 2947 7563 3253
rect 7516 2756 7523 2813
rect 7496 2727 7503 2743
rect 7536 2727 7543 2743
rect 7436 2527 7443 2613
rect 7556 2587 7563 2763
rect 7576 2747 7583 3193
rect 7596 3036 7603 3213
rect 7616 3187 7623 3243
rect 7656 3147 7663 3243
rect 7616 3007 7623 3023
rect 7656 3016 7663 3033
rect 7296 2307 7303 2493
rect 7336 2387 7343 2523
rect 7376 2307 7383 2313
rect 7316 2276 7323 2293
rect 7256 2096 7263 2253
rect 7336 2167 7343 2263
rect 7376 2167 7383 2293
rect 7236 2087 7243 2093
rect 7276 2076 7303 2083
rect 7196 1816 7203 1973
rect 7156 1787 7163 1813
rect 7116 1776 7143 1783
rect 7116 1596 7123 1753
rect 7036 1287 7043 1323
rect 7016 847 7023 1193
rect 7036 1107 7043 1273
rect 7136 1147 7143 1776
rect 7176 1667 7183 1803
rect 7216 1787 7223 1833
rect 7236 1627 7243 2033
rect 7296 1767 7303 2076
rect 7196 1567 7203 1613
rect 7216 1587 7223 1613
rect 7236 1596 7263 1603
rect 7236 1547 7243 1596
rect 7116 1087 7123 1103
rect 6996 787 7003 823
rect 6776 367 6783 633
rect 6836 596 6843 653
rect 6856 616 6863 713
rect 6876 607 6883 633
rect 6876 327 6883 363
rect 6916 287 6923 713
rect 7016 636 7023 653
rect 7056 636 7063 753
rect 6916 163 6923 273
rect 6976 227 6983 613
rect 7036 607 7043 623
rect 7056 376 7063 393
rect 6856 156 6883 163
rect 6896 156 6923 163
rect 7016 156 7023 293
rect 7076 187 7083 273
rect 7096 267 7103 383
rect 7116 347 7123 353
rect 4996 -24 5023 -17
rect 5156 -24 5183 -17
rect 5196 -24 5223 -17
rect 6116 -24 6123 13
rect 6516 -24 6523 156
rect 6716 -17 6723 156
rect 6876 -17 6883 156
rect 7076 136 7083 173
rect 7136 147 7143 173
rect 7156 147 7163 1473
rect 7236 1427 7243 1533
rect 7196 1327 7203 1343
rect 7176 1307 7183 1323
rect 7176 1027 7183 1293
rect 7216 1167 7223 1323
rect 7256 1307 7263 1473
rect 7236 1167 7243 1253
rect 7276 1247 7283 1493
rect 7236 1116 7243 1153
rect 7176 747 7183 823
rect 7196 616 7203 833
rect 7216 643 7223 823
rect 7256 767 7263 1103
rect 7296 1096 7303 1553
rect 7316 847 7323 1833
rect 7336 1823 7343 2133
rect 7396 2007 7403 2433
rect 7436 2183 7443 2433
rect 7456 2207 7463 2533
rect 7516 2467 7523 2513
rect 7576 2487 7583 2733
rect 7596 2727 7603 2753
rect 7536 2276 7543 2473
rect 7476 2247 7483 2263
rect 7576 2263 7583 2413
rect 7556 2256 7583 2263
rect 7416 2176 7443 2183
rect 7416 2087 7423 2176
rect 7476 2107 7483 2233
rect 7496 2076 7503 2133
rect 7436 1927 7443 2063
rect 7476 2027 7483 2063
rect 7336 1816 7363 1823
rect 7336 1267 7343 1573
rect 7356 1547 7363 1816
rect 7396 1607 7403 1873
rect 7436 1827 7443 1913
rect 7436 1767 7443 1813
rect 7396 1407 7403 1573
rect 7416 1563 7423 1673
rect 7496 1607 7503 1993
rect 7516 1583 7523 2153
rect 7596 2143 7603 2333
rect 7576 2136 7603 2143
rect 7576 2047 7583 2136
rect 7616 2123 7623 2993
rect 7636 2587 7643 2773
rect 7656 2127 7663 2893
rect 7676 2647 7683 3213
rect 7736 2847 7743 3033
rect 7756 3007 7763 3773
rect 7796 3767 7803 3933
rect 7836 3867 7843 3963
rect 7856 3843 7863 4493
rect 7896 4476 7903 4513
rect 8016 4247 8023 4693
rect 8036 4507 8043 5033
rect 8056 4627 8063 5053
rect 8056 4323 8063 4463
rect 8076 4407 8083 5053
rect 8136 4956 8143 4973
rect 8176 4956 8203 4963
rect 8116 4936 8123 4953
rect 8096 4687 8103 4793
rect 8036 4316 8063 4323
rect 7876 3947 7883 4193
rect 8036 4167 8043 4316
rect 8016 4147 8023 4163
rect 8116 3987 8123 4773
rect 8136 4696 8143 4753
rect 8196 4727 8203 4956
rect 8216 4947 8223 5253
rect 8236 4787 8243 5163
rect 8256 5007 8263 5796
rect 8356 5656 8363 5773
rect 8336 5607 8343 5623
rect 8176 4696 8183 4713
rect 8256 4687 8263 4953
rect 8196 4496 8203 4573
rect 8236 4463 8243 4473
rect 8216 4456 8243 4463
rect 8216 4447 8223 4456
rect 8176 4216 8183 4233
rect 8216 4207 8223 4313
rect 8276 4287 8283 5113
rect 8296 5027 8303 5273
rect 8316 5127 8323 5373
rect 8376 5127 8383 5753
rect 8396 5147 8403 5393
rect 8296 4956 8303 5013
rect 8336 4956 8343 5073
rect 8396 5003 8403 5133
rect 8376 4996 8403 5003
rect 8376 4967 8383 4996
rect 8416 4983 8423 5993
rect 8556 5923 8563 6213
rect 8636 6043 8643 6393
rect 8676 6136 8703 6143
rect 8616 6036 8643 6043
rect 8556 5916 8583 5923
rect 8496 5896 8523 5903
rect 8496 5767 8503 5896
rect 8476 5416 8483 5453
rect 8496 5443 8503 5653
rect 8496 5436 8523 5443
rect 8496 5207 8503 5403
rect 8496 5143 8503 5193
rect 8476 5136 8503 5143
rect 8447 5116 8463 5123
rect 8396 4976 8423 4983
rect 8356 4936 8383 4943
rect 8376 4927 8383 4936
rect 8396 4707 8403 4976
rect 8436 4867 8443 5073
rect 8356 4696 8383 4703
rect 8376 4687 8383 4696
rect 8316 4183 8323 4513
rect 8336 4467 8343 4683
rect 8356 4227 8363 4493
rect 8416 4487 8423 4853
rect 8436 4627 8443 4713
rect 8436 4463 8443 4613
rect 8456 4527 8463 4993
rect 8476 4967 8483 5136
rect 8496 4936 8503 4993
rect 8516 4787 8523 5436
rect 8536 5187 8543 5873
rect 8556 5656 8563 5813
rect 8576 5667 8583 5916
rect 8596 5647 8603 6033
rect 8616 5627 8623 6036
rect 8536 4927 8543 5173
rect 8556 5087 8563 5613
rect 8576 5467 8583 5623
rect 8636 5587 8643 5993
rect 8656 5416 8663 5893
rect 8676 5887 8683 6136
rect 8736 6007 8743 6773
rect 8756 6367 8763 6793
rect 8976 6787 8983 7373
rect 8996 6807 9003 7333
rect 9016 6927 9023 7573
rect 9056 7543 9063 7593
rect 9156 7587 9163 7713
rect 9176 7627 9183 7933
rect 9196 7887 9203 7933
rect 9196 7607 9203 7853
rect 9156 7556 9163 7573
rect 9036 7536 9063 7543
rect 9116 7347 9123 7493
rect 9136 7356 9143 7453
rect 9176 7356 9183 7373
rect 9036 6856 9043 7113
rect 9076 7087 9083 7313
rect 9136 7096 9143 7113
rect 9196 6967 9203 7073
rect 9216 7007 9223 7553
rect 9236 7547 9243 8023
rect 9276 8007 9283 8023
rect 9276 7827 9283 7973
rect 9296 7867 9303 8353
rect 9316 7887 9323 8396
rect 9376 8387 9383 8536
rect 9456 8447 9463 8613
rect 9476 8407 9483 10653
rect 9496 10567 9503 11176
rect 9536 11156 9543 11173
rect 9596 11163 9603 11213
rect 9576 11156 9603 11163
rect 9556 10936 9563 10953
rect 9516 10716 9523 10793
rect 9496 10167 9503 10273
rect 9536 10087 9543 10553
rect 9576 10267 9583 10973
rect 9596 10236 9603 10253
rect 9516 9583 9523 9983
rect 9576 9756 9583 10073
rect 9616 9927 9623 10253
rect 9636 10067 9643 11333
rect 9656 11127 9663 11416
rect 9716 11196 9723 11433
rect 9796 11403 9803 11513
rect 9936 11507 9943 11876
rect 10316 11847 10323 11883
rect 10396 11876 10423 11883
rect 10136 11723 10143 11843
rect 10316 11787 10323 11833
rect 10116 11716 10143 11723
rect 10116 11647 10123 11716
rect 10156 11647 10163 11663
rect 10276 11647 10283 11673
rect 10296 11587 10303 11673
rect 10376 11656 10383 11773
rect 10356 11636 10363 11653
rect 9796 11396 9823 11403
rect 9836 11307 9843 11423
rect 9876 11416 9903 11423
rect 9856 11387 9863 11403
rect 9736 11216 9743 11293
rect 9756 11196 9783 11203
rect 9776 10943 9783 11196
rect 9876 10963 9883 11373
rect 9896 11047 9903 11416
rect 9916 11207 9923 11233
rect 9936 11216 9943 11473
rect 9967 11216 9973 11223
rect 9956 11196 9983 11203
rect 9676 10923 9683 10933
rect 9676 10916 9703 10923
rect 9716 10747 9723 10943
rect 9756 10936 9783 10943
rect 9856 10956 9883 10963
rect 9856 10927 9863 10956
rect 9876 10936 9903 10943
rect 9936 10936 9943 11013
rect 9736 10907 9743 10923
rect 9876 10747 9883 10936
rect 9976 10927 9983 11196
rect 9936 10716 9943 10733
rect 9716 10696 9723 10713
rect 9656 10387 9663 10443
rect 9676 10287 9683 10463
rect 9716 10456 9723 10513
rect 9696 10427 9703 10433
rect 9676 10247 9683 10253
rect 9656 10087 9663 10233
rect 9736 10216 9743 10273
rect 9756 10236 9763 10713
rect 9996 10527 10003 11493
rect 10016 11363 10023 11413
rect 10256 11396 10263 11433
rect 10076 11367 10083 11383
rect 10016 11356 10063 11363
rect 9856 10407 9863 10443
rect 9876 10387 9883 10463
rect 9916 10456 9943 10463
rect 9936 10387 9943 10456
rect 9796 10236 9823 10243
rect 9596 9736 9623 9743
rect 9496 9576 9523 9583
rect 9496 9487 9503 9576
rect 9516 9547 9523 9553
rect 9516 9247 9523 9533
rect 9496 8976 9523 8983
rect 9496 8627 9503 8976
rect 9536 8843 9543 9093
rect 9556 9087 9563 9553
rect 9576 9476 9583 9513
rect 9616 9447 9623 9736
rect 9636 9647 9643 9743
rect 9656 9467 9663 9733
rect 9576 9227 9583 9253
rect 9656 9243 9663 9293
rect 9596 9207 9603 9243
rect 9636 9236 9663 9243
rect 9556 8947 9563 8983
rect 9516 8836 9543 8843
rect 9516 8543 9523 8836
rect 9556 8563 9563 8873
rect 9576 8767 9583 8853
rect 9596 8787 9603 9133
rect 9616 8947 9623 9013
rect 9616 8756 9623 8893
rect 9676 8887 9683 10053
rect 9696 9107 9703 10173
rect 9756 9927 9763 9943
rect 9736 9867 9743 9923
rect 9776 9867 9783 10223
rect 9816 10147 9823 10236
rect 9816 9887 9823 10133
rect 9836 10067 9843 10253
rect 9836 9947 9843 10053
rect 9856 9927 9863 10353
rect 9876 10227 9883 10373
rect 9956 10216 9963 10393
rect 9996 10203 10003 10273
rect 9876 9943 9883 10033
rect 9936 10007 9943 10203
rect 9976 10196 10003 10203
rect 10016 10183 10023 11293
rect 10087 11216 10133 11223
rect 10056 11167 10063 11213
rect 10196 11207 10203 11363
rect 10296 11216 10303 11573
rect 10396 11427 10403 11653
rect 10416 11587 10423 11876
rect 10576 11807 10583 11883
rect 10536 11656 10543 11793
rect 10416 11396 10423 11553
rect 10456 11487 10463 11633
rect 10456 11363 10463 11413
rect 10436 11356 10463 11363
rect 10536 11323 10543 11573
rect 10556 11367 10563 11643
rect 10616 11627 10623 11913
rect 10936 11896 10963 11903
rect 10656 11607 10663 11873
rect 10716 11827 10723 11863
rect 10696 11643 10703 11753
rect 10696 11636 10723 11643
rect 10656 11447 10663 11453
rect 10656 11407 10663 11433
rect 10536 11316 10563 11323
rect 10276 11196 10283 11213
rect 10416 11176 10443 11183
rect 10076 10943 10083 11163
rect 10136 11127 10143 11173
rect 10076 10936 10103 10943
rect 10056 10687 10063 10703
rect 10076 10547 10083 10903
rect 10096 10467 10103 10936
rect 10316 10936 10323 10973
rect 10176 10887 10183 10933
rect 10116 10427 10123 10493
rect 10056 10407 10063 10423
rect 10096 10383 10103 10423
rect 10067 10376 10103 10383
rect 10156 10327 10163 10713
rect 10087 10236 10103 10243
rect 10136 10236 10143 10253
rect 9996 10176 10023 10183
rect 9876 9936 9903 9943
rect 9776 9776 9783 9813
rect 9736 9756 9763 9763
rect 9736 9547 9743 9756
rect 9756 9327 9763 9463
rect 9716 9007 9723 9253
rect 9696 8976 9723 8983
rect 9636 8776 9643 8793
rect 9676 8763 9683 8813
rect 9656 8756 9683 8763
rect 9496 8536 9523 8543
rect 9536 8556 9563 8563
rect 9296 7836 9303 7853
rect 9256 7347 9263 7573
rect 9316 7543 9323 7833
rect 9336 7827 9343 8293
rect 9356 7727 9363 8313
rect 9416 8207 9423 8303
rect 9496 8263 9503 8536
rect 9516 8307 9523 8493
rect 9496 8256 9523 8263
rect 9416 8027 9423 8043
rect 9456 8036 9463 8193
rect 9496 8107 9503 8233
rect 9496 8023 9503 8093
rect 9516 8047 9523 8256
rect 9436 7987 9443 8023
rect 9476 8016 9503 8023
rect 9416 7856 9423 7873
rect 9456 7836 9483 7843
rect 9436 7767 9443 7823
rect 9356 7556 9363 7613
rect 9316 7536 9343 7543
rect 9376 7536 9403 7543
rect 9316 7387 9323 7536
rect 9276 7356 9303 7363
rect 9236 7063 9243 7213
rect 9276 7207 9283 7356
rect 9316 7327 9323 7343
rect 9376 7303 9383 7513
rect 9356 7296 9383 7303
rect 9336 7087 9343 7293
rect 9316 7067 9323 7083
rect 9236 7056 9263 7063
rect 9196 6876 9203 6953
rect 9236 6876 9243 6913
rect 9056 6787 9063 6843
rect 8796 6616 8823 6623
rect 8796 6587 8803 6616
rect 8856 6607 8863 6623
rect 8856 6527 8863 6593
rect 8876 6467 8883 6603
rect 9036 6596 9043 6633
rect 9116 6583 9123 6873
rect 9276 6616 9283 6753
rect 9296 6727 9303 7063
rect 8836 6396 8843 6433
rect 8816 6367 8823 6383
rect 8756 6127 8763 6233
rect 8736 5916 8743 5953
rect 8776 5916 8783 5933
rect 8696 5656 8723 5663
rect 8756 5656 8783 5663
rect 8696 5607 8703 5656
rect 8736 5627 8743 5643
rect 8636 5307 8643 5403
rect 8596 5176 8603 5193
rect 8696 4967 8703 5573
rect 8736 5067 8743 5573
rect 8756 5427 8763 5593
rect 8776 5443 8783 5656
rect 8796 5587 8803 6353
rect 8836 5807 8843 6333
rect 8856 6136 8863 6393
rect 8876 6347 8883 6453
rect 8896 6167 8903 6393
rect 8896 6136 8903 6153
rect 8916 6127 8923 6493
rect 8996 6396 9003 6493
rect 9056 6403 9063 6583
rect 9096 6576 9123 6583
rect 9036 6396 9063 6403
rect 8876 5947 8883 6123
rect 8936 5943 8943 6133
rect 9016 6027 9023 6143
rect 9036 6047 9043 6123
rect 8916 5936 8943 5943
rect 8916 5916 8923 5936
rect 9016 5907 9023 6013
rect 8936 5883 8943 5903
rect 8916 5876 8943 5883
rect 8916 5647 8923 5876
rect 8956 5636 8963 5773
rect 8776 5436 8803 5443
rect 8776 5307 8783 5436
rect 8856 5416 8863 5473
rect 8936 5427 8943 5623
rect 8996 5463 9003 5653
rect 8976 5456 9003 5463
rect 8976 5407 8983 5456
rect 9056 5416 9063 5893
rect 8876 5143 8883 5173
rect 8816 4987 8823 5143
rect 8856 5136 8883 5143
rect 8796 4936 8823 4943
rect 8816 4807 8823 4936
rect 8856 4867 8863 4913
rect 8496 4696 8503 4713
rect 8476 4547 8483 4693
rect 8736 4676 8743 4773
rect 8436 4456 8463 4463
rect 8396 4183 8403 4253
rect 8456 4196 8463 4273
rect 8316 4176 8343 4183
rect 8376 4176 8403 4183
rect 8376 4107 8383 4176
rect 8156 3996 8163 4013
rect 8036 3947 8043 3963
rect 7836 3836 7863 3843
rect 7796 3716 7803 3733
rect 7776 3667 7783 3683
rect 7816 3667 7823 3693
rect 7776 3467 7783 3573
rect 7836 3507 7843 3836
rect 7876 3567 7883 3933
rect 7856 3516 7863 3533
rect 7896 3527 7903 3713
rect 7776 3183 7783 3453
rect 7876 3243 7883 3513
rect 7776 3176 7803 3183
rect 7776 2807 7783 3176
rect 7796 3036 7803 3176
rect 7816 3063 7823 3243
rect 7856 3236 7883 3243
rect 7816 3056 7843 3063
rect 7836 3036 7843 3056
rect 7876 3036 7883 3093
rect 7896 3067 7903 3453
rect 7716 2716 7743 2723
rect 7736 2547 7743 2716
rect 7776 2707 7783 2753
rect 7796 2747 7803 2813
rect 7696 2487 7703 2543
rect 7716 2296 7723 2393
rect 7596 2116 7623 2123
rect 7556 2007 7563 2033
rect 7596 2027 7603 2116
rect 7616 2076 7623 2093
rect 7696 2076 7703 2153
rect 7536 1787 7543 1803
rect 7576 1796 7583 1893
rect 7556 1767 7563 1783
rect 7496 1576 7523 1583
rect 7416 1556 7443 1563
rect 7476 1556 7483 1573
rect 7516 1487 7523 1576
rect 7456 1387 7463 1453
rect 7476 1447 7483 1453
rect 7376 1207 7383 1323
rect 7416 1316 7423 1333
rect 7336 827 7343 1113
rect 7356 807 7363 1053
rect 7376 887 7383 1193
rect 7396 1187 7403 1303
rect 7436 1287 7443 1293
rect 7396 836 7403 1093
rect 7416 967 7423 1253
rect 7456 1187 7463 1353
rect 7476 1096 7483 1433
rect 7496 1287 7503 1393
rect 7576 1363 7583 1733
rect 7596 1687 7603 1783
rect 7616 1747 7623 2033
rect 7676 2007 7683 2063
rect 7556 1356 7583 1363
rect 7456 1067 7463 1083
rect 7496 1076 7503 1113
rect 7516 1107 7523 1293
rect 7536 987 7543 1333
rect 7416 803 7423 823
rect 7416 796 7443 803
rect 7256 727 7263 753
rect 7416 656 7423 753
rect 7436 667 7443 796
rect 7216 636 7243 643
rect 7236 627 7243 636
rect 7456 623 7463 713
rect 7436 616 7463 623
rect 7396 587 7403 613
rect 7416 607 7423 613
rect 7236 376 7263 383
rect 7236 327 7243 376
rect 7236 116 7243 153
rect 7256 136 7263 233
rect 7276 163 7283 363
rect 7316 307 7323 363
rect 7276 156 7303 163
rect 7296 123 7303 156
rect 7416 143 7423 453
rect 7456 343 7463 593
rect 7476 407 7483 873
rect 7496 827 7503 973
rect 7516 767 7523 853
rect 7536 667 7543 953
rect 7556 807 7563 1356
rect 7596 1343 7603 1593
rect 7616 1583 7623 1653
rect 7676 1647 7683 1933
rect 7716 1887 7723 2113
rect 7736 2047 7743 2283
rect 7756 2267 7763 2303
rect 7796 2283 7803 2573
rect 7816 2527 7823 2733
rect 7856 2556 7863 3023
rect 7916 2907 7923 3473
rect 7936 2807 7943 3853
rect 8016 3716 8023 3893
rect 7956 3627 7963 3703
rect 7996 3627 8003 3683
rect 8076 3496 8083 3733
rect 8136 3727 8143 3993
rect 8476 3987 8483 4533
rect 8216 3976 8243 3983
rect 8196 3647 8203 3743
rect 8216 3707 8223 3723
rect 8216 3587 8223 3693
rect 8236 3627 8243 3976
rect 8056 3427 8063 3483
rect 8096 3476 8103 3553
rect 8296 3527 8303 3753
rect 8336 3547 8343 3703
rect 8236 3516 8263 3523
rect 8116 3496 8123 3513
rect 8136 3427 8143 3513
rect 7956 3223 7963 3293
rect 7996 3247 8003 3373
rect 8236 3287 8243 3516
rect 7956 3216 7983 3223
rect 8036 3056 8043 3193
rect 8096 3087 8103 3233
rect 8016 2927 8023 3013
rect 7896 2576 7903 2793
rect 7776 2276 7803 2283
rect 7776 2007 7783 2113
rect 7796 2067 7803 2253
rect 7836 2103 7843 2553
rect 7936 2547 7943 2763
rect 7956 2707 7963 2783
rect 7996 2763 8003 2793
rect 8016 2787 8023 2853
rect 7976 2756 8003 2763
rect 7996 2747 8003 2756
rect 8056 2763 8063 3023
rect 8096 2947 8103 3073
rect 8096 2847 8103 2853
rect 8056 2756 8083 2763
rect 7956 2547 7963 2693
rect 7876 2523 7883 2533
rect 7856 2516 7883 2523
rect 7856 2407 7863 2516
rect 7856 2107 7863 2393
rect 7876 2227 7883 2293
rect 7896 2247 7903 2533
rect 7916 2527 7923 2543
rect 7976 2367 7983 2493
rect 7936 2276 7943 2313
rect 7976 2276 7983 2353
rect 7816 2096 7843 2103
rect 7736 1887 7743 1973
rect 7716 1823 7723 1873
rect 7716 1816 7743 1823
rect 7736 1796 7743 1816
rect 7796 1803 7803 1973
rect 7816 1827 7823 2096
rect 7876 2076 7883 2113
rect 7776 1796 7803 1803
rect 7716 1767 7723 1773
rect 7616 1576 7643 1583
rect 7676 1487 7683 1583
rect 7596 1336 7623 1343
rect 7616 1327 7623 1336
rect 7576 1307 7583 1323
rect 7596 1287 7603 1303
rect 7636 1207 7643 1303
rect 7696 1287 7703 1373
rect 7636 1103 7643 1193
rect 7716 1147 7723 1753
rect 7736 1567 7743 1593
rect 7756 1527 7763 1733
rect 7736 1507 7743 1513
rect 7776 1467 7783 1573
rect 7796 1407 7803 1773
rect 7836 1747 7843 1993
rect 7856 1727 7863 2013
rect 7936 2007 7943 2233
rect 7956 2227 7963 2243
rect 7876 1787 7883 1853
rect 7896 1747 7903 1993
rect 7936 1796 7943 1853
rect 7956 1847 7963 2213
rect 7976 2067 7983 2093
rect 7996 2007 8003 2513
rect 8036 2187 8043 2753
rect 8076 2707 8083 2756
rect 8096 2743 8103 2833
rect 8156 2783 8163 3273
rect 8216 3043 8223 3113
rect 8216 3036 8243 3043
rect 8256 3036 8263 3053
rect 8236 2807 8243 3036
rect 8336 3027 8343 3333
rect 8376 3267 8383 3703
rect 8396 3627 8403 3723
rect 8456 3516 8463 3633
rect 8436 3487 8443 3503
rect 8476 3496 8483 3533
rect 8156 2776 8183 2783
rect 8096 2736 8123 2743
rect 8056 2556 8063 2693
rect 8076 2587 8083 2693
rect 8076 2556 8103 2563
rect 7856 1596 7863 1653
rect 7896 1607 7903 1713
rect 7916 1687 7923 1783
rect 7816 1343 7823 1513
rect 7856 1467 7863 1553
rect 7816 1336 7863 1343
rect 7776 1316 7783 1333
rect 7816 1316 7823 1336
rect 7856 1307 7863 1336
rect 7796 1287 7803 1303
rect 7836 1287 7843 1303
rect 7736 1123 7743 1173
rect 7716 1116 7743 1123
rect 7636 1096 7663 1103
rect 7556 656 7563 673
rect 7576 647 7583 823
rect 7596 727 7603 803
rect 7616 787 7623 823
rect 7616 687 7623 773
rect 7636 727 7643 873
rect 7476 376 7483 393
rect 7436 336 7463 343
rect 7456 156 7463 253
rect 7496 156 7523 163
rect 7416 136 7443 143
rect 7276 116 7303 123
rect 7516 107 7523 156
rect 7536 147 7543 333
rect 7616 327 7623 393
rect 7636 356 7643 653
rect 7656 627 7663 793
rect 7696 647 7703 1093
rect 7736 1047 7743 1116
rect 7716 667 7723 913
rect 7756 823 7763 1133
rect 7776 1107 7783 1133
rect 7796 847 7803 1233
rect 7836 907 7843 1173
rect 7856 1096 7863 1273
rect 7876 1247 7883 1553
rect 7896 1367 7903 1513
rect 7916 1447 7923 1673
rect 7936 1527 7943 1733
rect 7996 1687 8003 1893
rect 7896 1267 7903 1333
rect 7916 1307 7923 1333
rect 7916 1187 7923 1273
rect 7916 1116 7923 1133
rect 7896 1007 7903 1103
rect 7836 836 7843 893
rect 7756 816 7783 823
rect 7776 687 7783 816
rect 7656 507 7663 613
rect 7736 567 7743 673
rect 7816 636 7823 653
rect 7836 607 7843 713
rect 7856 647 7863 823
rect 7896 807 7903 833
rect 7936 647 7943 1433
rect 7956 1307 7963 1593
rect 8016 1567 8023 2133
rect 8076 2127 8083 2556
rect 8176 2327 8183 2776
rect 8356 2763 8363 3053
rect 8336 2756 8363 2763
rect 8196 2467 8203 2613
rect 8256 2607 8263 2753
rect 8276 2727 8283 2743
rect 8256 2583 8263 2593
rect 8256 2576 8283 2583
rect 8276 2556 8283 2576
rect 8216 2536 8243 2543
rect 8096 2276 8123 2283
rect 8096 2207 8103 2276
rect 8196 2267 8203 2453
rect 8047 2096 8083 2103
rect 8076 2076 8083 2096
rect 8056 2027 8063 2063
rect 8096 2056 8103 2093
rect 8116 1867 8123 2253
rect 8136 2247 8143 2263
rect 8136 2067 8143 2093
rect 8136 1907 8143 2033
rect 8156 1947 8163 2113
rect 8176 2047 8183 2113
rect 8076 1747 8083 1813
rect 8036 1547 8043 1563
rect 8076 1527 8083 1563
rect 7976 1316 7983 1393
rect 8016 1347 8023 1373
rect 8016 1316 8023 1333
rect 7856 607 7863 633
rect 7656 387 7663 433
rect 7676 407 7683 453
rect 7676 356 7683 393
rect 7716 343 7723 353
rect 7696 336 7723 343
rect 7736 327 7743 533
rect 7616 147 7623 173
rect 7636 136 7643 293
rect 7696 156 7703 173
rect 7796 127 7803 553
rect 7816 347 7823 473
rect 7836 356 7843 373
rect 7876 163 7883 633
rect 7956 627 7963 1273
rect 7996 1127 8003 1283
rect 8036 1267 8043 1303
rect 8056 1247 8063 1453
rect 8096 1287 8103 1813
rect 8116 1347 8123 1853
rect 8156 1796 8163 1873
rect 8176 1827 8183 2033
rect 8196 1847 8203 2233
rect 8216 2087 8223 2473
rect 8236 2387 8243 2536
rect 8236 2147 8243 2373
rect 8256 2127 8263 2313
rect 8276 2127 8283 2333
rect 8316 2287 8323 2493
rect 8356 2387 8363 2756
rect 8376 2527 8383 3193
rect 8396 2927 8403 3233
rect 8416 3187 8423 3223
rect 8456 3087 8463 3223
rect 8496 3207 8503 4613
rect 8516 4203 8523 4513
rect 8536 4456 8543 4513
rect 8716 4496 8723 4663
rect 8756 4647 8763 4663
rect 8776 4647 8783 4693
rect 8736 4447 8743 4473
rect 8516 4196 8543 4203
rect 8516 4187 8523 4196
rect 8516 3976 8523 4173
rect 8816 4047 8823 4473
rect 8836 4456 8843 4793
rect 8856 4443 8863 4853
rect 8876 4727 8883 5136
rect 8896 5127 8903 5153
rect 8936 4927 8943 5213
rect 8976 5207 8983 5393
rect 8976 5176 8983 5193
rect 9016 5176 9023 5233
rect 8956 5027 8963 5053
rect 8956 4923 8963 5013
rect 8956 4916 8983 4923
rect 8876 4663 8883 4713
rect 8876 4656 8903 4663
rect 8856 4436 8883 4443
rect 8876 4227 8883 4436
rect 8976 4247 8983 4916
rect 9016 4907 9023 4923
rect 9076 4627 9083 6413
rect 9096 5883 9103 6333
rect 9116 6087 9123 6576
rect 9256 6407 9263 6453
rect 9276 6387 9283 6453
rect 9176 6376 9203 6383
rect 9176 6167 9183 6376
rect 9116 5927 9123 6073
rect 9176 5947 9183 6153
rect 9216 6116 9223 6353
rect 9236 6027 9243 6083
rect 9296 6047 9303 6613
rect 9336 6347 9343 6893
rect 9276 5887 9283 5913
rect 9316 5896 9323 6093
rect 9096 5876 9123 5883
rect 9096 5667 9103 5876
rect 9116 5636 9123 5813
rect 9156 5687 9163 5873
rect 9356 5747 9363 7296
rect 9396 6907 9403 7536
rect 9416 7067 9423 7733
rect 9476 7567 9483 7836
rect 9516 7447 9523 7673
rect 9536 7527 9543 8556
rect 9576 8503 9583 8613
rect 9696 8547 9703 8773
rect 9556 8496 9583 8503
rect 9576 8336 9583 8433
rect 9556 8316 9563 8333
rect 9596 8316 9603 8333
rect 9616 8056 9623 8333
rect 9656 8227 9663 8493
rect 9696 8463 9703 8503
rect 9676 8456 9703 8463
rect 9676 8187 9683 8456
rect 9716 8367 9723 8976
rect 9736 8927 9743 8983
rect 9736 8887 9743 8913
rect 9736 8516 9743 8833
rect 9756 8603 9763 9313
rect 9776 9276 9803 9283
rect 9836 9276 9863 9283
rect 9776 9247 9783 9276
rect 9856 9087 9863 9276
rect 9876 9047 9883 9853
rect 9896 9796 9943 9803
rect 9896 9787 9903 9796
rect 9936 9783 9943 9796
rect 9936 9776 9963 9783
rect 9916 9756 9923 9773
rect 9956 9756 9963 9776
rect 9976 9747 9983 10173
rect 9936 9607 9943 9743
rect 9896 9487 9903 9593
rect 9916 9496 9923 9573
rect 9956 9527 9963 9653
rect 9956 9496 9963 9513
rect 9856 8996 9883 9003
rect 9916 8996 9923 9353
rect 9936 9027 9943 9473
rect 9996 9467 10003 10176
rect 10076 10007 10083 10233
rect 10116 10127 10123 10223
rect 10156 10216 10163 10313
rect 10036 9976 10063 9983
rect 10096 9976 10103 10013
rect 10036 9667 10043 9976
rect 10076 9947 10083 9963
rect 10116 9783 10123 9973
rect 10156 9927 10163 9993
rect 10096 9776 10123 9783
rect 9807 8836 9843 8843
rect 9796 8796 9803 8813
rect 9836 8796 9843 8836
rect 9756 8596 9783 8603
rect 9716 8327 9723 8333
rect 9696 8187 9703 8313
rect 9576 7827 9583 8053
rect 9596 7836 9603 7853
rect 9616 7667 9623 8013
rect 9636 7927 9643 8033
rect 9636 7836 9643 7853
rect 9556 7576 9563 7593
rect 9616 7583 9623 7653
rect 9596 7576 9623 7583
rect 9576 7507 9583 7563
rect 9536 7407 9543 7433
rect 9456 6947 9463 7373
rect 9556 7356 9563 7453
rect 9476 6967 9483 7063
rect 9476 6867 9483 6953
rect 9576 6863 9583 6873
rect 9556 6856 9583 6863
rect 9616 6616 9623 6873
rect 9416 6596 9443 6603
rect 9376 6447 9383 6573
rect 9396 6527 9403 6563
rect 9376 6396 9383 6433
rect 9396 6416 9403 6453
rect 9436 6403 9443 6596
rect 9416 6396 9443 6403
rect 9436 6167 9443 6293
rect 9536 6287 9543 6613
rect 9596 6567 9603 6603
rect 9556 6363 9563 6393
rect 9596 6376 9603 6433
rect 9636 6427 9643 7773
rect 9656 7507 9663 8063
rect 9716 7527 9723 7853
rect 9736 7787 9743 8253
rect 9756 8247 9763 8283
rect 9756 7587 9763 8213
rect 9776 8087 9783 8596
rect 9796 8107 9803 8453
rect 9816 8227 9823 8733
rect 9836 8267 9843 8573
rect 9856 8267 9863 8996
rect 9876 8587 9883 8953
rect 9896 8947 9903 8963
rect 9896 8907 9903 8933
rect 9876 8536 9883 8553
rect 9916 8536 9923 8793
rect 9936 8567 9943 8983
rect 9956 8967 9963 9453
rect 9996 9256 10003 9293
rect 10016 9236 10023 9533
rect 10036 9507 10043 9653
rect 10096 9476 10103 9776
rect 10116 9756 10143 9763
rect 10156 9756 10163 9913
rect 10176 9807 10183 10753
rect 10196 10727 10203 10933
rect 10236 10716 10243 10733
rect 10116 9407 10123 9433
rect 9976 8943 9983 9213
rect 10036 9067 10043 9133
rect 9956 8936 9983 8943
rect 9776 8067 9783 8073
rect 9816 8056 9823 8133
rect 9776 7823 9783 8033
rect 9796 8027 9803 8053
rect 9856 7836 9863 7853
rect 9776 7816 9803 7823
rect 9876 7667 9883 7833
rect 9767 7576 9783 7583
rect 9736 7547 9743 7563
rect 9776 7556 9783 7576
rect 9896 7547 9903 8523
rect 9936 8296 9943 8513
rect 9956 8403 9963 8936
rect 9996 8776 10003 8813
rect 9976 8527 9983 8763
rect 10016 8756 10023 8793
rect 10036 8776 10043 9053
rect 10056 8543 10063 9013
rect 10036 8536 10063 8543
rect 10036 8507 10043 8536
rect 10076 8527 10083 9353
rect 10136 9347 10143 9756
rect 10196 9367 10203 10453
rect 10136 9207 10143 9333
rect 10196 9296 10203 9313
rect 10216 9303 10223 10703
rect 10256 10696 10263 10913
rect 10416 10696 10423 11176
rect 10456 11156 10463 11313
rect 10516 11167 10523 11193
rect 10536 10903 10543 11193
rect 10516 10896 10543 10903
rect 10396 10627 10403 10683
rect 10256 10267 10263 10443
rect 10276 10347 10283 10423
rect 10316 10347 10323 10423
rect 10316 10327 10323 10333
rect 10316 10216 10323 10253
rect 10336 10236 10343 10313
rect 10396 10267 10403 10613
rect 10376 10236 10383 10253
rect 10396 10187 10403 10253
rect 10256 9927 10263 9943
rect 10276 9496 10283 9513
rect 10256 9447 10263 9483
rect 10296 9327 10303 9893
rect 10316 9736 10323 10093
rect 10396 10007 10403 10153
rect 10416 10047 10423 10513
rect 10436 10467 10443 10683
rect 10536 10467 10543 10896
rect 10556 10607 10563 11316
rect 10636 11223 10643 11403
rect 10616 11216 10643 11223
rect 10656 11216 10663 11273
rect 10436 10407 10443 10433
rect 10456 10427 10463 10443
rect 10416 9907 10423 9943
rect 10436 9927 10443 10393
rect 10476 10387 10483 10423
rect 10496 10327 10503 10373
rect 10516 10347 10523 10423
rect 10536 10367 10543 10433
rect 10576 10327 10583 11173
rect 10616 10883 10623 11216
rect 10676 11196 10703 11203
rect 10696 10887 10703 11196
rect 10616 10876 10643 10883
rect 10616 10767 10623 10876
rect 10596 10667 10603 10683
rect 10636 10667 10643 10683
rect 10596 10527 10603 10633
rect 10376 9756 10383 9773
rect 10216 9296 10243 9303
rect 10156 9276 10183 9283
rect 10156 9227 10163 9276
rect 10096 8767 10103 8973
rect 10116 8803 10123 8983
rect 10156 8887 10163 8933
rect 10116 8796 10143 8803
rect 10156 8796 10163 8873
rect 10176 8823 10183 8993
rect 10196 8967 10203 9253
rect 10236 9167 10243 9296
rect 10176 8816 10203 8823
rect 10196 8796 10203 8816
rect 10216 8807 10223 8853
rect 10047 8496 10063 8503
rect 10096 8467 10103 8503
rect 10116 8487 10123 8513
rect 9956 8396 9983 8403
rect 9916 8147 9923 8283
rect 9956 8267 9963 8283
rect 9976 8243 9983 8396
rect 10076 8347 10083 8373
rect 9956 8236 9983 8243
rect 9916 8027 9923 8133
rect 9936 7827 9943 7973
rect 9956 7867 9963 8236
rect 9976 8023 9983 8093
rect 10056 8023 10063 8233
rect 9976 8016 10003 8023
rect 10036 8016 10063 8023
rect 9736 7383 9743 7533
rect 9756 7487 9763 7543
rect 9796 7527 9803 7543
rect 9796 7507 9803 7513
rect 9716 7376 9743 7383
rect 9836 7356 9843 7433
rect 9876 7356 9883 7533
rect 9696 7087 9703 7343
rect 9896 7307 9903 7373
rect 9676 6847 9683 7063
rect 9716 6907 9723 7053
rect 9876 6887 9883 7063
rect 9896 7027 9903 7083
rect 9736 6876 9763 6883
rect 9656 6567 9663 6613
rect 9676 6587 9683 6833
rect 9736 6807 9743 6876
rect 9776 6847 9783 6863
rect 9756 6596 9763 6793
rect 9556 6356 9583 6363
rect 9616 6347 9623 6363
rect 9436 6116 9443 6153
rect 9676 6147 9683 6573
rect 9716 6416 9743 6423
rect 9716 6287 9723 6416
rect 9776 6367 9783 6583
rect 9796 6567 9803 6603
rect 9796 6387 9803 6553
rect 9816 6147 9823 6713
rect 9896 6587 9903 6633
rect 9916 6627 9923 6843
rect 9956 6767 9963 6843
rect 9976 6687 9983 8016
rect 10016 7996 10043 8003
rect 9996 7887 10003 7913
rect 10016 7816 10023 7873
rect 9996 7783 10003 7803
rect 10036 7796 10043 7996
rect 10056 7816 10063 7993
rect 10096 7967 10103 8303
rect 10116 8287 10123 8333
rect 10096 7827 10103 7953
rect 9996 7776 10023 7783
rect 9996 7367 10003 7653
rect 10016 7547 10023 7776
rect 10076 7576 10103 7583
rect 10136 7576 10143 8796
rect 10216 8776 10223 8793
rect 10196 8503 10203 8753
rect 10236 8727 10243 9153
rect 10256 8983 10263 9313
rect 10276 9267 10283 9313
rect 10316 9287 10323 9493
rect 10356 9387 10363 9743
rect 10396 9427 10403 9513
rect 10416 9447 10423 9853
rect 10456 9807 10463 9943
rect 10496 9907 10503 10233
rect 10556 10147 10563 10203
rect 10496 9723 10503 9813
rect 10536 9736 10543 10113
rect 10496 9716 10523 9723
rect 10436 9496 10443 9573
rect 10476 9496 10483 9713
rect 10396 9296 10403 9413
rect 10356 9276 10363 9293
rect 10256 8976 10283 8983
rect 10276 8887 10283 8976
rect 10296 8927 10303 9273
rect 10436 9263 10443 9273
rect 10416 9256 10443 9263
rect 10456 9247 10463 9483
rect 10216 8567 10223 8593
rect 10196 8496 10223 8503
rect 10156 8047 10163 8473
rect 10236 8447 10243 8483
rect 10196 8063 10203 8393
rect 10236 8347 10243 8353
rect 10236 8316 10243 8333
rect 10276 8323 10283 8833
rect 10296 8367 10303 8913
rect 10316 8467 10323 8973
rect 10336 8747 10343 8973
rect 10356 8787 10363 9213
rect 10496 9207 10503 9693
rect 10516 9267 10523 9716
rect 10576 9707 10583 10233
rect 10596 9987 10603 10513
rect 10616 10267 10623 10453
rect 10636 10347 10643 10653
rect 10676 10467 10683 10673
rect 10716 10587 10723 11613
rect 10656 10387 10663 10443
rect 10736 10387 10743 11573
rect 10756 11007 10763 11863
rect 10776 11416 10783 11433
rect 10796 11387 10803 11403
rect 10836 11367 10843 11793
rect 10856 11287 10863 11833
rect 10896 11656 10903 11853
rect 10916 11847 10923 11883
rect 10936 11687 10943 11713
rect 10936 11643 10943 11673
rect 10876 11627 10883 11643
rect 10916 11636 10943 11643
rect 10796 11196 10823 11203
rect 10596 9747 10603 9943
rect 10656 9927 10663 9963
rect 10576 9283 10583 9513
rect 10596 9347 10603 9483
rect 10616 9447 10623 9503
rect 10656 9496 10663 9553
rect 10676 9507 10683 10333
rect 10696 10247 10703 10373
rect 10756 10267 10763 10753
rect 10796 10747 10803 11196
rect 10816 10767 10823 10903
rect 10856 10723 10863 10893
rect 10876 10727 10883 11613
rect 10896 11147 10903 11413
rect 10956 11407 10963 11896
rect 11236 11896 11263 11903
rect 11296 11896 11303 11913
rect 11056 11747 11063 11873
rect 10836 10716 10863 10723
rect 10816 10683 10823 10703
rect 10796 10676 10823 10683
rect 10776 10367 10783 10433
rect 10796 10307 10803 10676
rect 10856 10667 10863 10716
rect 10716 10236 10723 10253
rect 10756 10236 10783 10243
rect 10696 10027 10703 10173
rect 10736 10127 10743 10223
rect 10756 9927 10763 10193
rect 10776 10147 10783 10236
rect 10776 9987 10783 10133
rect 10696 9727 10703 9743
rect 10716 9527 10723 9693
rect 10576 9276 10603 9283
rect 10376 8987 10383 9053
rect 10396 8783 10403 8873
rect 10376 8776 10403 8783
rect 10436 8727 10443 9193
rect 10376 8536 10403 8543
rect 10436 8536 10443 8653
rect 10276 8316 10303 8323
rect 10216 8287 10223 8313
rect 10236 8107 10243 8253
rect 10196 8056 10223 8063
rect 10216 8047 10223 8056
rect 10236 8036 10243 8093
rect 10176 8007 10183 8023
rect 10216 7856 10223 7873
rect 10076 7527 10083 7576
rect 10116 7527 10123 7563
rect 10016 7107 10023 7373
rect 10036 7356 10043 7473
rect 10076 7356 10083 7373
rect 10036 7096 10063 7103
rect 10036 6987 10043 7096
rect 10076 7067 10083 7083
rect 10156 7027 10163 7853
rect 10176 7836 10203 7843
rect 10236 7836 10243 7993
rect 10176 7427 10183 7836
rect 10296 7583 10303 8316
rect 10316 8007 10323 8333
rect 10336 7907 10343 8453
rect 10376 8107 10383 8536
rect 10456 8527 10463 8953
rect 10456 8296 10463 8513
rect 10476 8287 10483 8453
rect 10516 8267 10523 8773
rect 10396 8056 10403 8173
rect 10536 8127 10543 9233
rect 10556 9187 10563 9243
rect 10596 9236 10603 9276
rect 10556 9027 10563 9073
rect 10556 8987 10563 9013
rect 10576 9007 10583 9093
rect 10576 8776 10583 8993
rect 10596 8987 10603 9093
rect 10556 8747 10563 8763
rect 10556 8207 10563 8733
rect 10616 8647 10623 9193
rect 10596 8516 10603 8633
rect 10616 8423 10623 8483
rect 10636 8467 10643 9433
rect 10656 9267 10663 9453
rect 10656 9187 10663 9253
rect 10716 9107 10723 9493
rect 10716 9007 10723 9033
rect 10676 8867 10683 8963
rect 10676 8427 10683 8813
rect 10696 8796 10723 8803
rect 10696 8687 10703 8796
rect 10696 8467 10703 8673
rect 10616 8416 10643 8423
rect 10636 8307 10643 8416
rect 10676 8283 10683 8313
rect 10616 8267 10623 8283
rect 10656 8276 10683 8283
rect 10336 7883 10343 7893
rect 10336 7876 10363 7883
rect 10336 7667 10343 7853
rect 10356 7836 10363 7876
rect 10416 7867 10423 8073
rect 10596 8036 10603 8113
rect 10616 8067 10623 8253
rect 10576 7967 10583 8023
rect 10636 7987 10643 8053
rect 10416 7816 10423 7853
rect 10276 7576 10303 7583
rect 10276 7556 10283 7576
rect 10336 7563 10343 7653
rect 10456 7627 10463 7813
rect 10316 7556 10343 7563
rect 10456 7576 10483 7583
rect 10256 7507 10263 7543
rect 10296 7387 10303 7543
rect 10176 7376 10223 7383
rect 10176 7347 10183 7376
rect 10416 7376 10423 7413
rect 10436 7387 10443 7493
rect 10236 7356 10243 7373
rect 10376 7356 10403 7363
rect 10436 7356 10443 7373
rect 10456 7367 10463 7576
rect 10496 7387 10503 7553
rect 10516 7507 10523 7583
rect 10556 7563 10563 7853
rect 10616 7836 10623 7893
rect 10596 7767 10603 7793
rect 10536 7556 10563 7563
rect 10636 7547 10643 7953
rect 10696 7747 10703 8433
rect 10716 8027 10723 8433
rect 10716 7843 10723 8013
rect 10736 7867 10743 9893
rect 10756 9627 10763 9773
rect 10776 9547 10783 9953
rect 10796 9527 10803 10253
rect 10816 10167 10823 10573
rect 10896 10487 10903 10713
rect 10876 10387 10883 10423
rect 10876 10287 10883 10373
rect 10896 10243 10903 10313
rect 10916 10267 10923 11393
rect 10996 11363 11003 11413
rect 11016 11387 11023 11433
rect 10956 11356 11003 11363
rect 10936 10347 10943 11353
rect 11036 11307 11043 11693
rect 11096 11627 11103 11643
rect 11016 11216 11043 11223
rect 11036 11087 11043 11216
rect 10996 10936 11023 10943
rect 10996 10907 11003 10936
rect 10976 10787 10983 10903
rect 10976 10743 10983 10773
rect 10976 10736 11003 10743
rect 10956 10716 10983 10723
rect 10956 10627 10963 10716
rect 10956 10427 10963 10613
rect 10896 10236 10923 10243
rect 10916 10216 10923 10236
rect 10876 9943 10883 10053
rect 10856 9936 10883 9943
rect 10856 9736 10863 9873
rect 10896 9767 10903 9993
rect 10916 9887 10923 10113
rect 10936 10027 10943 10203
rect 10956 10003 10963 10253
rect 10976 10007 10983 10493
rect 10936 9996 10963 10003
rect 10836 9607 10843 9723
rect 10756 9487 10763 9513
rect 10776 9496 10803 9503
rect 10776 9467 10783 9496
rect 10776 9347 10783 9433
rect 10776 9256 10783 9333
rect 10816 9243 10823 9313
rect 10756 9207 10763 9243
rect 10796 9236 10823 9243
rect 10756 8827 10763 9193
rect 10776 9027 10783 9173
rect 10776 8803 10783 9013
rect 10756 8796 10783 8803
rect 10776 8767 10783 8796
rect 10796 8767 10803 9093
rect 10816 8987 10823 9236
rect 10836 8967 10843 9453
rect 10856 9307 10863 9533
rect 10876 9507 10883 9723
rect 10876 9427 10883 9493
rect 10896 9467 10903 9753
rect 10916 9447 10923 9733
rect 10936 9347 10943 9996
rect 10996 9976 11003 10736
rect 11016 10727 11023 10873
rect 11036 10463 11043 10713
rect 11056 10507 11063 11183
rect 11076 10967 11083 11493
rect 11096 11447 11103 11613
rect 11116 11167 11123 11363
rect 11136 11227 11143 11273
rect 11136 11176 11143 11213
rect 11136 10627 11143 11073
rect 11156 11067 11163 11893
rect 11176 11167 11183 11593
rect 11196 11347 11203 11793
rect 11236 11527 11243 11896
rect 11936 11896 11963 11903
rect 11276 11747 11283 11883
rect 11296 11656 11303 11673
rect 11336 11643 11343 11713
rect 11316 11636 11343 11643
rect 11296 11407 11303 11423
rect 11276 11307 11283 11403
rect 11356 11383 11363 11773
rect 11376 11607 11383 11833
rect 11396 11587 11403 11873
rect 11416 11627 11423 11863
rect 11596 11847 11603 11863
rect 11636 11847 11643 11863
rect 11476 11696 11483 11753
rect 11436 11676 11463 11683
rect 11336 11376 11363 11383
rect 11316 11216 11323 11373
rect 11336 11207 11343 11376
rect 11156 10723 11163 10933
rect 11216 10916 11223 10933
rect 11196 10727 11203 10883
rect 11236 10847 11243 10903
rect 11156 10716 11183 10723
rect 11176 10696 11183 10716
rect 11016 10456 11043 10463
rect 11016 10067 11023 10456
rect 11116 10443 11123 10553
rect 11096 10436 11123 10443
rect 11036 10287 11043 10423
rect 11136 10307 11143 10573
rect 11156 10387 11163 10683
rect 11036 10127 11043 10273
rect 11056 10256 11063 10293
rect 11096 10223 11103 10253
rect 11076 10216 11103 10223
rect 10976 9947 10983 9963
rect 11016 9767 11023 9973
rect 10956 9327 10963 9753
rect 11036 9716 11043 9873
rect 11056 9847 11063 10213
rect 11076 9947 11083 10013
rect 10996 9647 11003 9673
rect 10996 9487 11003 9633
rect 11016 9456 11043 9463
rect 10896 9276 10913 9283
rect 10896 9243 10903 9276
rect 10956 9276 10963 9293
rect 10896 9236 10923 9243
rect 10836 8787 10843 8953
rect 10856 8887 10863 8983
rect 10916 8963 10923 9236
rect 10936 9227 10943 9263
rect 10876 8927 10883 8963
rect 10896 8956 10923 8963
rect 10896 8867 10903 8956
rect 10916 8887 10923 8913
rect 10796 8503 10803 8713
rect 10836 8547 10843 8773
rect 10836 8507 10843 8533
rect 10776 8496 10803 8503
rect 10796 8316 10803 8496
rect 10816 8487 10823 8503
rect 10816 8327 10823 8413
rect 10836 8107 10843 8213
rect 10756 7887 10763 8043
rect 10796 8036 10803 8053
rect 10836 8023 10843 8093
rect 10816 8016 10843 8023
rect 10716 7836 10743 7843
rect 10776 7836 10783 7893
rect 10856 7867 10863 8273
rect 10796 7816 10803 7853
rect 10856 7847 10863 7853
rect 10876 7827 10883 8633
rect 10896 8327 10903 8853
rect 10916 8796 10923 8873
rect 10956 8707 10963 9233
rect 10916 8287 10923 8553
rect 10916 8187 10923 8273
rect 10936 7963 10943 8693
rect 10976 8647 10983 9113
rect 10996 8567 11003 9333
rect 11016 9267 11023 9433
rect 11016 9067 11023 9253
rect 11036 9107 11043 9456
rect 11096 9303 11103 10053
rect 11116 9987 11123 10253
rect 11156 9967 11163 10113
rect 11196 10007 11203 10613
rect 11216 10427 11223 10693
rect 11256 10547 11263 11053
rect 11296 10507 11303 10993
rect 11316 10847 11323 11173
rect 11336 11047 11343 11173
rect 11356 10923 11363 11073
rect 11416 11067 11423 11593
rect 11436 11507 11443 11676
rect 11516 11643 11523 11833
rect 11496 11636 11523 11643
rect 11456 11247 11463 11573
rect 11476 11267 11483 11383
rect 11467 11156 11483 11163
rect 11456 11107 11463 11153
rect 11436 10936 11443 10953
rect 11356 10916 11383 10923
rect 11336 10696 11343 10733
rect 11356 10667 11363 10683
rect 11316 10443 11323 10553
rect 11296 10436 11323 10443
rect 11216 10247 11223 10393
rect 11236 10267 11243 10423
rect 11227 10236 11243 10243
rect 11236 10216 11243 10236
rect 11216 10187 11223 10203
rect 11116 9407 11123 9953
rect 11136 9927 11143 9943
rect 11156 9447 11163 9733
rect 11176 9447 11183 9873
rect 11196 9867 11203 9963
rect 11216 9807 11223 9953
rect 11236 9907 11243 10173
rect 11276 10047 11283 10373
rect 11256 9947 11263 10033
rect 11196 9547 11203 9773
rect 11216 9756 11223 9793
rect 11236 9776 11243 9833
rect 11276 9787 11283 9993
rect 11256 9756 11283 9763
rect 11196 9487 11203 9513
rect 11136 9367 11143 9433
rect 11156 9307 11163 9393
rect 11076 9296 11103 9303
rect 11076 8987 11083 9296
rect 11156 9256 11163 9293
rect 11176 9247 11183 9393
rect 11016 8967 11023 8983
rect 10956 8447 10963 8503
rect 10976 8467 10983 8483
rect 10976 8387 10983 8453
rect 11016 8347 11023 8793
rect 11036 8627 11043 8963
rect 11036 8507 11043 8613
rect 11056 8347 11063 8953
rect 11076 8807 11083 8953
rect 11116 8947 11123 9233
rect 11116 8796 11123 8933
rect 11136 8763 11143 9173
rect 11196 9047 11203 9433
rect 11216 9427 11223 9443
rect 11216 9187 11223 9353
rect 11236 9327 11243 9533
rect 11256 9047 11263 9593
rect 11276 9527 11283 9756
rect 11296 9503 11303 10413
rect 11276 9496 11303 9503
rect 11156 8887 11163 9033
rect 11116 8756 11143 8763
rect 10996 8067 11003 8293
rect 11016 8047 11023 8253
rect 10916 7956 10943 7963
rect 10716 7543 10723 7713
rect 10696 7536 10723 7543
rect 10376 7307 10383 7356
rect 10276 7096 10283 7293
rect 10296 7047 10303 7093
rect 10316 7047 10323 7063
rect 10036 6827 10043 6853
rect 10056 6767 10063 6893
rect 10076 6827 10083 6843
rect 10016 6596 10023 6613
rect 10056 6583 10063 6753
rect 10196 6607 10203 6873
rect 10236 6836 10263 6843
rect 10236 6583 10243 6836
rect 10316 6607 10323 6853
rect 9616 6136 9643 6143
rect 9136 5187 9143 5623
rect 9176 5607 9183 5623
rect 9216 5416 9223 5593
rect 9256 5407 9263 5453
rect 9196 5327 9203 5403
rect 9236 5396 9253 5403
rect 9216 5156 9223 5173
rect 9276 5143 9283 5453
rect 9176 4936 9183 5133
rect 9196 5027 9203 5143
rect 9236 5136 9283 5143
rect 9236 4943 9243 4953
rect 9236 4936 9263 4943
rect 9096 4647 9103 4663
rect 9096 4476 9103 4633
rect 9116 4467 9123 4513
rect 8696 4016 8703 4033
rect 8836 3983 8843 4203
rect 8816 3976 8843 3983
rect 8836 3847 8843 3976
rect 8556 3716 8563 3773
rect 8616 3647 8623 3703
rect 8656 3516 8663 3713
rect 8776 3676 8803 3683
rect 8516 3307 8523 3513
rect 8676 3496 8703 3503
rect 8536 3227 8543 3293
rect 8616 3236 8623 3313
rect 8696 3287 8703 3496
rect 8676 3236 8683 3253
rect 8476 3036 8483 3053
rect 8416 3016 8423 3033
rect 8456 2987 8463 3023
rect 8416 2607 8423 2873
rect 8456 2743 8463 2813
rect 8456 2736 8483 2743
rect 8416 2556 8423 2593
rect 8376 2283 8383 2313
rect 8436 2287 8443 2573
rect 8456 2563 8463 2693
rect 8556 2567 8563 2743
rect 8456 2556 8483 2563
rect 8356 2276 8383 2283
rect 8296 2207 8303 2253
rect 8336 2243 8343 2263
rect 8316 2236 8343 2243
rect 8276 2076 8283 2093
rect 8216 2027 8223 2053
rect 8256 2047 8263 2063
rect 8296 2056 8303 2133
rect 8316 2023 8323 2236
rect 8296 2016 8323 2023
rect 8216 1823 8223 1893
rect 8196 1816 8223 1823
rect 8196 1796 8203 1816
rect 8136 1763 8143 1783
rect 8136 1756 8163 1763
rect 8136 1567 8143 1573
rect 8136 1287 8143 1553
rect 8156 1307 8163 1756
rect 8176 1587 8183 1763
rect 8196 1596 8223 1603
rect 8196 1427 8203 1596
rect 8216 1427 8223 1533
rect 8056 1136 8063 1233
rect 8076 1027 8083 1093
rect 8016 887 8023 953
rect 8016 856 8023 873
rect 7976 567 7983 603
rect 7896 356 7903 413
rect 7996 387 8003 833
rect 8076 787 8083 1013
rect 8096 867 8103 1013
rect 8136 847 8143 1113
rect 8176 887 8183 1273
rect 8196 1047 8203 1273
rect 8216 1087 8223 1413
rect 8236 1343 8243 1993
rect 8256 1947 8263 2013
rect 8256 1596 8263 1933
rect 8296 1907 8303 2016
rect 8336 2003 8343 2193
rect 8316 1996 8343 2003
rect 8316 1823 8323 1996
rect 8356 1947 8363 2213
rect 8376 1987 8383 2253
rect 8476 2227 8483 2556
rect 8576 2543 8583 2993
rect 8596 2747 8603 3223
rect 8716 3167 8723 3253
rect 8616 3036 8623 3073
rect 8656 2647 8663 2753
rect 8676 2743 8683 2833
rect 8696 2763 8703 3033
rect 8776 3007 8783 3676
rect 8876 3523 8883 3793
rect 8856 3516 8883 3523
rect 8856 3447 8863 3516
rect 8796 3227 8803 3253
rect 8836 3236 8843 3373
rect 8836 3036 8843 3193
rect 8856 3087 8863 3203
rect 8876 3036 8883 3193
rect 8796 3007 8803 3033
rect 8816 3016 8823 3033
rect 8856 2987 8863 3023
rect 8696 2756 8723 2763
rect 8676 2736 8703 2743
rect 8676 2556 8683 2573
rect 8556 2536 8583 2543
rect 8596 2536 8623 2543
rect 8536 2307 8543 2373
rect 8556 2367 8563 2536
rect 8596 2407 8603 2536
rect 8656 2447 8663 2543
rect 8576 2327 8583 2373
rect 8536 2276 8543 2293
rect 8576 2276 8583 2313
rect 8596 2243 8603 2333
rect 8556 2207 8563 2243
rect 8576 2236 8603 2243
rect 8296 1816 8323 1823
rect 8276 1787 8283 1813
rect 8276 1647 8283 1653
rect 8296 1447 8303 1816
rect 8336 1796 8343 1813
rect 8396 1803 8403 2093
rect 8416 2067 8423 2133
rect 8476 2076 8483 2153
rect 8527 2076 8543 2083
rect 8436 2056 8463 2063
rect 8436 1927 8443 2056
rect 8536 2043 8543 2076
rect 8556 2067 8563 2093
rect 8516 2036 8543 2043
rect 8376 1796 8403 1803
rect 8316 1767 8323 1783
rect 8316 1667 8323 1713
rect 8336 1667 8343 1713
rect 8416 1596 8423 1733
rect 8336 1527 8343 1573
rect 8396 1567 8403 1583
rect 8436 1576 8443 1733
rect 8456 1543 8463 1973
rect 8476 1807 8483 1813
rect 8476 1627 8483 1793
rect 8436 1536 8463 1543
rect 8236 1336 8263 1343
rect 8236 847 8243 1313
rect 8256 1127 8263 1336
rect 8276 1096 8283 1193
rect 8316 1147 8323 1513
rect 8316 1096 8323 1133
rect 8396 1107 8403 1323
rect 8436 1136 8443 1536
rect 8456 1307 8463 1333
rect 8476 1187 8483 1533
rect 8156 803 8163 833
rect 8156 796 8203 803
rect 8196 636 8203 673
rect 8216 647 8223 823
rect 8116 616 8143 623
rect 8116 587 8123 616
rect 8216 587 8223 633
rect 8036 343 8043 453
rect 8116 356 8123 393
rect 8036 336 8063 343
rect 8136 307 8143 343
rect 7876 156 7903 163
rect 7816 123 7823 153
rect 7916 147 7923 173
rect 8016 156 8043 163
rect 7816 116 7843 123
rect 7836 103 7843 116
rect 7876 103 7883 113
rect 8016 107 8023 156
rect 8116 143 8123 253
rect 8236 187 8243 573
rect 8256 363 8263 1083
rect 8296 667 8303 913
rect 8316 667 8323 893
rect 8416 836 8423 1093
rect 8476 947 8483 1173
rect 8336 663 8343 833
rect 8356 767 8363 823
rect 8336 656 8363 663
rect 8316 636 8323 653
rect 8356 636 8363 656
rect 8376 616 8383 633
rect 8276 547 8283 613
rect 8336 376 8343 433
rect 8396 427 8403 753
rect 8416 387 8423 653
rect 8476 607 8483 933
rect 8496 807 8503 2033
rect 8516 1767 8523 2036
rect 8576 1987 8583 2236
rect 8536 1787 8543 1803
rect 8576 1796 8583 1873
rect 8596 1867 8603 2213
rect 8616 1783 8623 2393
rect 8636 2307 8643 2313
rect 8636 2067 8643 2293
rect 8676 2267 8683 2353
rect 8696 2107 8703 2736
rect 8716 2547 8723 2756
rect 8736 2727 8743 2743
rect 8736 2347 8743 2713
rect 8796 2707 8803 2753
rect 8856 2727 8863 2813
rect 8776 2556 8803 2563
rect 8836 2556 8843 2653
rect 8776 2547 8783 2556
rect 8776 2467 8783 2533
rect 8756 2323 8763 2333
rect 8736 2316 8763 2323
rect 8736 2307 8743 2316
rect 8756 2276 8763 2293
rect 8856 2267 8863 2593
rect 8776 2256 8803 2263
rect 8716 1967 8723 2063
rect 8736 1967 8743 2113
rect 8596 1776 8623 1783
rect 8516 847 8523 1153
rect 8536 1087 8543 1673
rect 8556 1527 8563 1753
rect 8576 1596 8583 1613
rect 8636 1603 8643 1873
rect 8716 1867 8723 1953
rect 8696 1767 8703 1853
rect 8756 1796 8763 2173
rect 8776 1743 8783 1783
rect 8796 1767 8803 2256
rect 8876 2127 8883 2973
rect 8896 2747 8903 4053
rect 8916 3967 8923 4213
rect 8956 3716 8963 3973
rect 8976 3947 8983 4233
rect 9016 4216 9023 4273
rect 9056 3963 9063 4013
rect 9036 3956 9063 3963
rect 9156 3963 9163 4873
rect 9196 4727 9203 4923
rect 9196 4647 9203 4713
rect 9256 4707 9263 4936
rect 9296 4887 9303 5733
rect 9416 5703 9423 6103
rect 9456 6087 9463 6103
rect 9456 5936 9523 5943
rect 9396 5696 9423 5703
rect 9396 5663 9403 5696
rect 9376 5656 9403 5663
rect 9316 5636 9343 5643
rect 9376 5636 9383 5656
rect 9316 5167 9323 5636
rect 9356 5587 9363 5623
rect 9396 5616 9413 5623
rect 9436 5487 9443 5933
rect 9456 5627 9463 5936
rect 9516 5916 9523 5936
rect 9536 5896 9543 5933
rect 9496 5887 9503 5893
rect 9596 5867 9603 6113
rect 9636 6087 9643 6136
rect 9756 6116 9763 6133
rect 9896 6127 9903 6573
rect 9996 6427 10003 6583
rect 10036 6576 10063 6583
rect 10216 6576 10243 6583
rect 9976 6363 9983 6393
rect 9956 6356 9983 6363
rect 9956 6136 9963 6153
rect 9656 5887 9663 6073
rect 9676 5916 9683 6053
rect 9816 6047 9823 6093
rect 9716 5916 9723 5933
rect 9756 5916 9783 5923
rect 9776 5907 9783 5916
rect 9696 5887 9703 5903
rect 9536 5636 9543 5713
rect 9576 5647 9583 5853
rect 9656 5627 9663 5873
rect 9736 5867 9743 5903
rect 9776 5656 9783 5713
rect 9816 5627 9823 6033
rect 9936 5927 9943 6103
rect 9896 5707 9903 5883
rect 9936 5656 9943 5693
rect 9976 5656 9983 6333
rect 9416 5436 9423 5453
rect 9336 5327 9343 5413
rect 9356 5367 9363 5433
rect 9396 5407 9403 5423
rect 9436 5416 9443 5473
rect 9556 5467 9563 5623
rect 9596 5416 9603 5623
rect 9796 5507 9803 5623
rect 9716 5427 9723 5493
rect 9736 5436 9763 5443
rect 9716 5407 9723 5413
rect 9576 5387 9583 5403
rect 9736 5387 9743 5436
rect 9816 5416 9823 5473
rect 9956 5467 9963 5643
rect 10036 5627 10043 6553
rect 10076 6396 10083 6413
rect 10116 6396 10123 6413
rect 10136 6376 10143 6433
rect 10136 6136 10163 6143
rect 10136 6067 10143 6136
rect 10156 5927 10163 5933
rect 10056 5916 10083 5923
rect 10056 5707 10063 5916
rect 10136 5896 10143 5913
rect 10176 5907 10183 6103
rect 10196 5927 10203 6393
rect 10256 6347 10263 6593
rect 10276 6347 10283 6383
rect 10336 6163 10343 7133
rect 10496 7087 10503 7373
rect 10536 7067 10543 7373
rect 10556 7336 10563 7473
rect 10596 7336 10603 7373
rect 10636 7347 10643 7513
rect 10676 7487 10683 7523
rect 10576 7316 10583 7333
rect 10616 7207 10623 7323
rect 10636 7076 10643 7293
rect 10736 7287 10743 7733
rect 10896 7543 10903 7793
rect 10876 7536 10903 7543
rect 10856 7507 10863 7523
rect 10916 7467 10923 7956
rect 10936 7856 10943 7933
rect 10816 7356 10843 7363
rect 10836 7167 10843 7356
rect 10916 7327 10923 7393
rect 10936 7303 10943 7813
rect 10956 7787 10963 7823
rect 10976 7763 10983 8003
rect 10996 7987 11003 8023
rect 10956 7756 10983 7763
rect 10956 7367 10963 7756
rect 11016 7576 11023 8033
rect 11056 7727 11063 8313
rect 11076 7567 11083 8753
rect 11116 8467 11123 8756
rect 11196 8563 11203 8993
rect 11236 8983 11243 9033
rect 11216 8976 11243 8983
rect 11216 8787 11223 8976
rect 11256 8867 11263 9013
rect 11276 8927 11283 9496
rect 11236 8796 11243 8853
rect 11256 8816 11263 8853
rect 11276 8827 11283 8833
rect 11276 8796 11283 8813
rect 11296 8807 11303 9473
rect 11316 9287 11323 10413
rect 11336 10127 11343 10613
rect 11336 9787 11343 9933
rect 11356 9547 11363 10453
rect 11376 10427 11383 10873
rect 11416 10827 11423 10923
rect 11456 10887 11463 11053
rect 11476 10807 11483 10973
rect 11496 10783 11503 11636
rect 11516 11416 11523 11433
rect 11536 11427 11543 11673
rect 11556 11607 11563 11643
rect 11536 11327 11543 11383
rect 11516 10987 11523 11233
rect 11536 11127 11543 11193
rect 11476 10776 11503 10783
rect 11396 10427 11403 10553
rect 11376 10227 11383 10393
rect 11396 10207 11403 10293
rect 11416 10267 11423 10753
rect 11436 10667 11443 10713
rect 11456 10467 11463 10773
rect 11476 10627 11483 10776
rect 11516 10767 11523 10953
rect 11536 10887 11543 11033
rect 11556 10967 11563 11493
rect 11576 11447 11583 11833
rect 11616 11787 11623 11843
rect 11596 11656 11623 11663
rect 11576 10943 11583 11413
rect 11556 10936 11583 10943
rect 11496 10716 11503 10733
rect 11556 10727 11563 10936
rect 11516 10527 11523 10703
rect 11496 10427 11503 10443
rect 11436 10227 11443 10233
rect 11407 10196 11423 10203
rect 11376 9976 11383 10013
rect 11396 9907 11403 9943
rect 11416 9927 11423 10173
rect 11376 9647 11383 9853
rect 11416 9827 11423 9893
rect 11436 9887 11443 10113
rect 11456 9947 11463 10193
rect 11396 9756 11403 9793
rect 11416 9776 11423 9813
rect 11356 9476 11363 9513
rect 11396 9467 11403 9483
rect 11336 9407 11343 9463
rect 11376 9447 11383 9463
rect 11336 9276 11343 9313
rect 11396 9307 11403 9453
rect 11376 9276 11383 9293
rect 11316 9007 11323 9133
rect 11356 9047 11363 9263
rect 11396 9027 11403 9273
rect 11336 9016 11363 9023
rect 11336 8927 11343 9016
rect 11196 8556 11223 8563
rect 11176 8536 11203 8543
rect 11096 8087 11103 8333
rect 11116 8327 11123 8433
rect 11116 8127 11123 8293
rect 11136 8107 11143 8393
rect 11196 8383 11203 8536
rect 11216 8407 11223 8556
rect 11176 8376 11203 8383
rect 11156 8267 11163 8333
rect 11176 8243 11183 8376
rect 11236 8323 11243 8533
rect 11256 8487 11263 8773
rect 11296 8483 11303 8793
rect 11316 8547 11323 8913
rect 11276 8476 11303 8483
rect 11236 8316 11263 8323
rect 11196 8267 11203 8273
rect 11176 8236 11193 8243
rect 11096 7687 11103 8053
rect 11156 8036 11163 8053
rect 11196 8007 11203 8233
rect 11236 8227 11243 8283
rect 11216 7967 11223 8113
rect 11136 7816 11143 7853
rect 11176 7816 11183 7953
rect 11236 7607 11243 8093
rect 11256 7827 11263 8316
rect 11276 8047 11283 8476
rect 11276 7987 11283 8033
rect 11296 7887 11303 8453
rect 11316 8207 11323 8493
rect 11336 8347 11343 8913
rect 11356 8487 11363 8493
rect 11376 8367 11383 8853
rect 11416 8803 11423 9513
rect 11436 8947 11443 9533
rect 11396 8796 11423 8803
rect 11436 8796 11443 8873
rect 11456 8827 11463 9913
rect 11476 9527 11483 10253
rect 11496 9767 11503 10213
rect 11496 9747 11503 9753
rect 11476 8823 11483 9493
rect 11496 9323 11503 9573
rect 11516 9507 11523 10493
rect 11536 9847 11543 10533
rect 11576 10483 11583 10793
rect 11556 10476 11583 10483
rect 11556 10227 11563 10476
rect 11596 10407 11603 11613
rect 11616 11527 11623 11656
rect 11696 11567 11703 11893
rect 11756 11863 11763 11873
rect 11756 11856 11783 11863
rect 11816 11767 11823 11863
rect 11716 11696 11723 11713
rect 11616 11223 11623 11293
rect 11636 11247 11643 11433
rect 11656 11383 11663 11553
rect 11656 11376 11683 11383
rect 11616 11216 11643 11223
rect 11656 11196 11663 11333
rect 11676 11163 11683 11376
rect 11656 11156 11683 11163
rect 11616 10947 11623 10993
rect 11616 10747 11623 10903
rect 11636 10767 11643 11133
rect 11616 10687 11623 10733
rect 11616 10567 11623 10673
rect 11636 10527 11643 10713
rect 11656 10707 11663 11156
rect 11676 10936 11683 11093
rect 11696 10787 11703 11233
rect 11716 11107 11723 11163
rect 11676 10716 11703 10723
rect 11616 10256 11623 10493
rect 11676 10487 11683 10716
rect 11716 10567 11723 10923
rect 11736 10747 11743 11553
rect 11756 11176 11763 11513
rect 11776 11047 11783 11453
rect 11796 11387 11803 11413
rect 11816 11407 11823 11533
rect 11836 11347 11843 11413
rect 11856 11027 11863 11473
rect 11916 11467 11923 11853
rect 11936 11587 11943 11896
rect 11976 11867 11983 11883
rect 11976 11567 11983 11663
rect 11996 11487 12003 11753
rect 11916 11367 11923 11423
rect 11936 11387 11943 11403
rect 11876 11216 11883 11353
rect 12016 11147 12023 11733
rect 11736 10667 11743 10683
rect 11656 10436 11663 10453
rect 11636 10287 11643 10423
rect 11636 10267 11643 10273
rect 11576 10236 11603 10243
rect 11636 10236 11643 10253
rect 11556 9976 11563 10193
rect 11576 10007 11583 10236
rect 11596 9976 11623 9983
rect 11556 9507 11563 9933
rect 11576 9867 11583 9953
rect 11616 9927 11623 9976
rect 11596 9547 11603 9733
rect 11576 9447 11583 9483
rect 11596 9467 11603 9493
rect 11616 9487 11623 9893
rect 11636 9887 11643 10153
rect 11656 10087 11663 10353
rect 11676 10167 11683 10393
rect 11696 10143 11703 10413
rect 11716 10367 11723 10453
rect 11716 10207 11723 10293
rect 11676 10136 11703 10143
rect 11496 9316 11523 9323
rect 11516 9296 11523 9316
rect 11536 9276 11563 9283
rect 11556 9267 11563 9276
rect 11496 9007 11503 9153
rect 11476 8816 11503 8823
rect 11396 8567 11403 8796
rect 11456 8747 11463 8783
rect 11416 8347 11423 8513
rect 11336 8227 11343 8333
rect 11376 8316 11383 8333
rect 11276 7623 11283 7853
rect 11316 7807 11323 8153
rect 11336 8056 11343 8073
rect 11356 8027 11363 8043
rect 11376 8007 11383 8063
rect 11396 7867 11403 8043
rect 11356 7767 11363 7803
rect 11276 7616 11303 7623
rect 11196 7576 11223 7583
rect 11036 7547 11043 7563
rect 11176 7447 11183 7573
rect 11196 7487 11203 7576
rect 11236 7543 11243 7563
rect 11236 7536 11253 7543
rect 11296 7527 11303 7616
rect 11176 7376 11183 7433
rect 11316 7383 11323 7753
rect 11356 7547 11363 7553
rect 11376 7547 11383 7793
rect 11396 7787 11403 7813
rect 11436 7603 11443 8553
rect 11496 8543 11503 8816
rect 11516 8607 11523 9233
rect 11536 9016 11543 9033
rect 11616 8987 11623 9373
rect 11636 9247 11643 9833
rect 11656 8967 11663 10073
rect 11676 9907 11683 10136
rect 11736 9987 11743 10513
rect 11756 10447 11763 10673
rect 11776 10427 11783 10733
rect 11796 10427 11803 10693
rect 11756 10027 11763 10413
rect 11776 10247 11783 10313
rect 11796 10216 11803 10353
rect 11816 10243 11823 11013
rect 11836 10367 11843 10833
rect 11916 10696 11923 10753
rect 11936 10667 11943 10683
rect 11936 10507 11943 10653
rect 11816 10236 11843 10243
rect 11696 9907 11703 9943
rect 11536 8587 11543 8813
rect 11556 8747 11563 8913
rect 11576 8807 11583 8853
rect 11476 8536 11503 8543
rect 11456 8027 11463 8353
rect 11456 7787 11463 7853
rect 11416 7596 11443 7603
rect 11387 7536 11403 7543
rect 11296 7376 11323 7383
rect 10976 7336 10983 7373
rect 10936 7296 10963 7303
rect 10816 7083 10823 7133
rect 10436 7007 10443 7063
rect 10607 7056 10623 7063
rect 10676 7027 10683 7083
rect 10816 7076 10843 7083
rect 10856 6947 10863 7063
rect 10896 6947 10903 7063
rect 10456 6807 10463 6863
rect 10576 6827 10583 6893
rect 10636 6876 10643 6933
rect 10416 6616 10443 6623
rect 10356 6447 10363 6603
rect 10436 6567 10443 6616
rect 10456 6383 10463 6753
rect 10676 6607 10683 6893
rect 10856 6876 10863 6913
rect 10776 6856 10803 6863
rect 10776 6787 10783 6856
rect 10776 6627 10783 6773
rect 10616 6596 10643 6603
rect 10556 6547 10563 6583
rect 10476 6396 10483 6473
rect 10636 6447 10643 6596
rect 10816 6596 10823 6833
rect 10876 6787 10883 6873
rect 10916 6867 10923 7053
rect 10676 6416 10683 6593
rect 10756 6567 10763 6583
rect 10796 6467 10803 6583
rect 10516 6396 10543 6403
rect 10536 6387 10543 6396
rect 10436 6376 10463 6383
rect 10316 6156 10343 6163
rect 10316 6136 10323 6156
rect 10356 6136 10363 6333
rect 10096 5887 10103 5893
rect 10196 5623 10203 5913
rect 10236 5647 10243 5913
rect 10256 5907 10263 5933
rect 10276 5916 10283 5933
rect 10336 5896 10343 6123
rect 10356 5647 10363 5913
rect 10176 5616 10203 5623
rect 10156 5507 10163 5603
rect 10176 5487 10183 5616
rect 9936 5427 9943 5453
rect 10016 5416 10023 5453
rect 9356 5176 9363 5193
rect 9396 5176 9403 5313
rect 9576 5247 9583 5373
rect 9556 5147 9563 5163
rect 9956 5156 9963 5193
rect 9576 5107 9583 5143
rect 9636 5107 9643 5153
rect 9776 5127 9783 5143
rect 9816 5127 9823 5143
rect 10036 5127 10043 5413
rect 10056 5407 10063 5433
rect 10076 5167 10083 5433
rect 10136 5227 10143 5453
rect 10196 5436 10203 5453
rect 10236 5447 10243 5633
rect 10216 5416 10223 5433
rect 10116 5156 10123 5173
rect 10156 5156 10163 5193
rect 10076 5143 10083 5153
rect 10076 5136 10103 5143
rect 9976 5007 9983 5123
rect 9276 4647 9283 4663
rect 9316 4487 9323 4993
rect 9336 4936 9343 4993
rect 9536 4807 9543 4933
rect 9616 4843 9623 4973
rect 9656 4907 9663 4933
rect 9816 4923 9823 4953
rect 9996 4936 10003 4953
rect 9896 4923 9903 4933
rect 9596 4836 9623 4843
rect 9456 4696 9463 4713
rect 9596 4667 9603 4836
rect 9656 4767 9663 4893
rect 9676 4867 9683 4923
rect 9816 4916 9843 4923
rect 9876 4916 9903 4923
rect 10036 4923 10043 4953
rect 10056 4927 10063 4973
rect 10016 4916 10043 4923
rect 9236 4227 9243 4443
rect 9256 4196 9263 4273
rect 9296 4207 9303 4213
rect 9296 4183 9303 4193
rect 9356 4187 9363 4653
rect 9696 4627 9703 4673
rect 9716 4667 9723 4713
rect 9796 4696 9803 4733
rect 9836 4696 9843 4713
rect 9436 4476 9443 4493
rect 9476 4476 9503 4483
rect 9496 4207 9503 4476
rect 9516 4447 9523 4463
rect 9596 4456 9603 4473
rect 9876 4456 9903 4463
rect 9876 4327 9883 4456
rect 9916 4443 9923 4853
rect 9996 4676 10003 4713
rect 10136 4687 10143 5143
rect 10176 5047 10183 5143
rect 10196 4987 10203 5213
rect 10216 4947 10223 4973
rect 10176 4927 10183 4943
rect 10236 4676 10243 4893
rect 10276 4807 10283 5493
rect 10316 5163 10323 5613
rect 10336 5447 10343 5623
rect 10376 5467 10383 5623
rect 10416 5483 10423 5633
rect 10436 5627 10443 6376
rect 10816 6376 10823 6433
rect 10836 6427 10843 6583
rect 10876 6407 10883 6413
rect 10936 6387 10943 6413
rect 10656 6347 10663 6373
rect 10956 6367 10963 7296
rect 10996 7287 11003 7323
rect 11156 7307 11163 7343
rect 11016 7076 11023 7093
rect 11156 7063 11163 7153
rect 11156 7056 11183 7063
rect 10976 6876 10983 6933
rect 11036 6887 11043 7053
rect 10996 6807 11003 6863
rect 10976 6407 10983 6603
rect 10996 6447 11003 6583
rect 11036 6547 11043 6583
rect 11056 6427 11063 6593
rect 10996 6416 11043 6423
rect 10996 6387 11003 6416
rect 11056 6396 11063 6413
rect 10496 6067 10503 6103
rect 10456 5903 10463 6053
rect 10496 5936 10503 5993
rect 10536 5947 10543 6103
rect 10556 6087 10563 6123
rect 10576 6007 10583 6113
rect 10456 5896 10483 5903
rect 10476 5607 10483 5713
rect 10556 5663 10563 5913
rect 10576 5907 10583 5933
rect 10536 5656 10563 5663
rect 10496 5636 10503 5653
rect 10536 5636 10543 5656
rect 10556 5483 10563 5623
rect 10396 5476 10443 5483
rect 10396 5427 10403 5476
rect 10436 5456 10443 5476
rect 10536 5476 10563 5483
rect 10416 5436 10423 5453
rect 10376 5187 10383 5423
rect 10316 5156 10343 5163
rect 10336 5067 10343 5156
rect 10416 5143 10423 5173
rect 10516 5163 10523 5433
rect 10536 5427 10543 5476
rect 10556 5436 10563 5453
rect 10516 5156 10543 5163
rect 10576 5156 10583 5413
rect 10396 5136 10423 5143
rect 10316 4936 10323 4993
rect 10336 4927 10343 5033
rect 10396 4923 10403 4973
rect 10376 4916 10403 4923
rect 10296 4707 10303 4913
rect 10016 4507 10023 4663
rect 10216 4567 10223 4663
rect 10036 4456 10063 4463
rect 10336 4456 10343 4473
rect 10376 4467 10383 4733
rect 10436 4727 10443 5153
rect 10536 5007 10543 5156
rect 10636 5147 10643 5393
rect 10536 4936 10543 4993
rect 10556 4987 10563 5143
rect 10596 4987 10603 4993
rect 10596 4956 10603 4973
rect 10436 4696 10463 4703
rect 10456 4687 10463 4696
rect 10416 4667 10423 4683
rect 9916 4436 9933 4443
rect 10056 4327 10063 4456
rect 10476 4287 10483 4733
rect 10496 4587 10503 4933
rect 10576 4907 10583 4943
rect 10536 4647 10543 4793
rect 10556 4696 10583 4703
rect 10616 4696 10623 4793
rect 10556 4567 10563 4696
rect 10556 4496 10563 4553
rect 10576 4476 10583 4633
rect 10596 4487 10603 4683
rect 10656 4387 10663 6313
rect 10776 6103 10783 6133
rect 10716 6007 10723 6103
rect 10756 6096 10783 6103
rect 10876 6087 10883 6153
rect 10956 6116 10983 6123
rect 10736 6007 10743 6073
rect 10716 5947 10723 5993
rect 10676 5916 10683 5933
rect 10736 5907 10743 5993
rect 10696 5727 10703 5903
rect 10756 5647 10763 5913
rect 10716 5587 10723 5643
rect 10696 5187 10703 5433
rect 10736 5427 10743 5623
rect 10776 5467 10783 5613
rect 10836 5607 10843 5813
rect 10876 5803 10883 5933
rect 10896 5927 10903 6103
rect 10976 6087 10983 6116
rect 10956 5916 10963 6073
rect 10876 5796 10903 5803
rect 10896 5667 10903 5796
rect 10896 5636 10903 5653
rect 10916 5643 10923 5873
rect 10936 5827 10943 5903
rect 10916 5636 10943 5643
rect 10796 5447 10803 5453
rect 10836 5447 10843 5573
rect 10856 5427 10863 5633
rect 10956 5487 10963 5623
rect 10736 5187 10743 5413
rect 10976 5407 10983 5423
rect 10696 5143 10703 5173
rect 10916 5143 10923 5173
rect 10696 5136 10723 5143
rect 10756 4983 10763 5143
rect 10916 5136 10943 5143
rect 10996 5127 11003 5613
rect 11016 5147 11023 5393
rect 10956 5107 10963 5123
rect 10736 4976 10763 4983
rect 10736 4967 10743 4976
rect 10816 4956 10823 5013
rect 10756 4696 10763 4913
rect 10776 4527 10783 4683
rect 10796 4476 10803 4613
rect 10856 4467 10863 4753
rect 10936 4707 10943 4973
rect 10936 4676 10943 4693
rect 10956 4627 10963 4643
rect 10976 4547 10983 4993
rect 10996 4956 11003 5113
rect 10976 4496 10983 4533
rect 10496 4247 10503 4253
rect 9756 4196 9763 4233
rect 9236 4167 9243 4183
rect 9276 4176 9303 4183
rect 9576 4183 9583 4193
rect 9196 4003 9203 4093
rect 9176 3996 9203 4003
rect 9156 3956 9183 3963
rect 8916 3207 8923 3473
rect 8916 3027 8923 3113
rect 8936 2987 8943 3133
rect 8896 2687 8903 2733
rect 8896 2287 8903 2673
rect 8916 2327 8923 2763
rect 8956 2756 8963 3513
rect 8976 3407 8983 3703
rect 8996 3627 9003 3953
rect 9056 3927 9063 3956
rect 9016 3687 9023 3713
rect 8996 3507 9003 3613
rect 9016 3516 9023 3533
rect 9116 3527 9123 3683
rect 9176 3547 9183 3956
rect 9196 3887 9203 3996
rect 9316 3967 9323 3993
rect 9376 3987 9383 4013
rect 9396 3996 9403 4053
rect 9416 4027 9423 4183
rect 9436 4003 9443 4153
rect 9456 4147 9463 4183
rect 9576 4176 9603 4183
rect 9436 3996 9463 4003
rect 9316 3947 9323 3953
rect 9256 3687 9263 3753
rect 9316 3716 9323 3933
rect 9076 3487 9083 3503
rect 8976 3227 8983 3253
rect 9016 3236 9023 3293
rect 8996 3147 9003 3223
rect 9096 3223 9103 3433
rect 9076 3216 9103 3223
rect 9116 3207 9123 3353
rect 9176 3307 9183 3533
rect 9276 3516 9283 3613
rect 9196 3496 9223 3503
rect 9176 3267 9183 3273
rect 8976 2867 8983 3013
rect 8996 2787 9003 3053
rect 9076 3003 9083 3053
rect 9056 2996 9083 3003
rect 9016 2907 9023 2993
rect 8936 2607 8943 2743
rect 8956 2543 8963 2713
rect 8976 2627 8983 2743
rect 8996 2576 9003 2773
rect 9016 2707 9023 2893
rect 9036 2727 9043 2873
rect 9056 2547 9063 2693
rect 8956 2536 8983 2543
rect 8956 2307 8963 2536
rect 8976 2276 8983 2293
rect 8816 2076 8843 2083
rect 8816 2067 8823 2076
rect 8776 1736 8803 1743
rect 8616 1596 8643 1603
rect 8776 1596 8783 1693
rect 8596 1547 8603 1583
rect 8556 1407 8563 1513
rect 8696 1467 8703 1573
rect 8796 1547 8803 1736
rect 8816 1596 8823 1733
rect 8856 1727 8863 2063
rect 8896 2056 8903 2253
rect 8916 2207 8923 2263
rect 8596 1327 8603 1433
rect 8576 1067 8583 1303
rect 8596 1083 8603 1193
rect 8676 1083 8683 1313
rect 8696 1123 8703 1453
rect 8716 1307 8723 1313
rect 8796 1303 8803 1393
rect 8727 1296 8743 1303
rect 8776 1296 8803 1303
rect 8696 1116 8723 1123
rect 8596 1076 8623 1083
rect 8656 1076 8683 1083
rect 8676 1027 8683 1076
rect 8536 947 8543 973
rect 8596 847 8603 873
rect 8496 636 8523 643
rect 8556 636 8563 693
rect 8256 356 8283 363
rect 8476 347 8483 593
rect 8496 547 8503 636
rect 8496 407 8503 533
rect 8536 527 8543 623
rect 8576 616 8583 793
rect 8056 127 8063 143
rect 8096 136 8123 143
rect 8236 136 8243 173
rect 8256 156 8263 213
rect 8276 127 8283 143
rect 8396 127 8403 173
rect 8416 156 8423 273
rect 8476 163 8483 333
rect 8536 323 8543 393
rect 8596 367 8603 773
rect 8616 707 8623 823
rect 8636 747 8643 973
rect 8696 907 8703 1093
rect 8616 687 8623 693
rect 8616 447 8623 653
rect 8656 647 8663 833
rect 8676 527 8683 633
rect 8696 627 8703 893
rect 8716 747 8723 1116
rect 8716 567 8723 673
rect 8736 667 8743 1253
rect 8756 1207 8763 1283
rect 8876 1143 8883 1953
rect 8896 1247 8903 1733
rect 8916 1707 8923 2093
rect 8936 1907 8943 2073
rect 8956 1807 8963 2263
rect 8976 1987 8983 2113
rect 8996 2047 9003 2153
rect 8996 1783 9003 1793
rect 8976 1776 9003 1783
rect 8936 1387 8943 1733
rect 8956 1627 8963 1763
rect 9016 1687 9023 2473
rect 9036 1867 9043 2513
rect 9076 2507 9083 2773
rect 9056 2076 9063 2413
rect 9076 2267 9083 2313
rect 9096 2107 9103 2993
rect 9116 2827 9123 3173
rect 9136 3007 9143 3033
rect 9136 2756 9143 2913
rect 9156 2787 9163 3193
rect 9176 3067 9183 3253
rect 9196 2907 9203 3496
rect 9236 3287 9243 3413
rect 9236 3236 9243 3273
rect 9256 3267 9263 3503
rect 9296 3467 9303 3673
rect 9316 3267 9323 3293
rect 9276 3236 9303 3243
rect 9256 3187 9263 3203
rect 9216 3036 9223 3153
rect 9176 2756 9183 2813
rect 9116 2647 9123 2743
rect 9136 2507 9143 2533
rect 9156 2307 9163 2653
rect 9236 2587 9243 2893
rect 9196 2507 9203 2523
rect 9136 2076 9143 2113
rect 9156 2067 9163 2273
rect 9176 2247 9183 2353
rect 9076 2007 9083 2063
rect 8976 1583 8983 1613
rect 8996 1596 9003 1653
rect 9036 1603 9043 1753
rect 9036 1596 9063 1603
rect 8956 1576 8983 1583
rect 8956 1407 8963 1576
rect 9016 1547 9023 1583
rect 9056 1567 9063 1596
rect 8936 1316 8943 1333
rect 8976 1316 8983 1533
rect 8996 1487 9003 1513
rect 9016 1303 9023 1333
rect 8876 1136 8903 1143
rect 8856 1116 8883 1123
rect 8776 1096 8803 1103
rect 8776 1007 8783 1096
rect 8836 1087 8843 1103
rect 8756 687 8763 823
rect 8796 787 8803 823
rect 8747 636 8763 643
rect 8816 627 8823 733
rect 8516 316 8543 323
rect 8456 156 8483 163
rect 8616 156 8623 433
rect 8656 356 8663 373
rect 8696 347 8703 363
rect 8716 347 8723 553
rect 8736 347 8743 373
rect 8676 267 8683 343
rect 8756 156 8763 333
rect 8816 163 8823 493
rect 8796 156 8823 163
rect 8836 147 8843 833
rect 8856 487 8863 1073
rect 8876 1067 8883 1116
rect 8896 847 8903 1136
rect 8916 887 8923 1303
rect 8956 1087 8963 1303
rect 8996 1296 9023 1303
rect 8976 1116 8983 1153
rect 9036 1096 9043 1473
rect 9056 1327 9063 1353
rect 9076 1267 9083 1993
rect 9116 1947 9123 2053
rect 9116 1867 9123 1933
rect 9096 1796 9103 1853
rect 9156 1763 9163 1783
rect 9136 1756 9163 1763
rect 9096 1667 9103 1673
rect 8896 816 8923 823
rect 8876 567 8883 633
rect 8896 627 8903 816
rect 8956 807 8963 823
rect 8916 636 8923 733
rect 8936 663 8943 793
rect 8996 767 9003 823
rect 9016 807 9023 833
rect 9076 827 9083 1233
rect 9096 1127 9103 1653
rect 9116 1307 9123 1713
rect 9136 1487 9143 1756
rect 9176 1727 9183 2073
rect 9196 1767 9203 2493
rect 9216 2007 9223 2093
rect 9236 1887 9243 2523
rect 9256 2307 9263 3133
rect 9276 2487 9283 3173
rect 9296 3147 9303 3236
rect 9296 2887 9303 3033
rect 9316 2907 9323 3253
rect 9336 3027 9343 3073
rect 9316 2887 9323 2893
rect 9296 2763 9303 2853
rect 9356 2847 9363 3873
rect 9416 3867 9423 3953
rect 9376 3407 9383 3613
rect 9376 3207 9383 3393
rect 9396 3347 9403 3533
rect 9416 3516 9423 3853
rect 9456 3527 9463 3996
rect 9476 3987 9483 4053
rect 9396 3236 9403 3253
rect 9436 3236 9443 3253
rect 9376 3036 9383 3053
rect 9416 3036 9423 3093
rect 9396 2807 9403 2853
rect 9296 2756 9323 2763
rect 9336 2727 9343 2743
rect 9316 2347 9323 2553
rect 9336 2547 9343 2633
rect 9336 2283 9343 2453
rect 9316 2276 9343 2283
rect 9216 1767 9223 1793
rect 9236 1596 9243 1873
rect 9256 1827 9263 2253
rect 9276 2076 9283 2133
rect 9296 2127 9303 2263
rect 9356 2167 9363 2633
rect 9376 2587 9383 2743
rect 9356 2063 9363 2113
rect 9336 2056 9363 2063
rect 9296 1796 9303 1973
rect 9156 1576 9183 1583
rect 9156 1547 9163 1576
rect 9196 1307 9203 1343
rect 9216 1247 9223 1323
rect 9236 1247 9243 1533
rect 9256 1447 9263 1553
rect 9216 1167 9223 1233
rect 9256 1183 9263 1333
rect 9276 1287 9283 1573
rect 9276 1267 9283 1273
rect 9256 1176 9283 1183
rect 8936 656 8963 663
rect 8956 636 8963 656
rect 8896 587 8903 613
rect 8936 567 8943 623
rect 8856 287 8863 363
rect 8896 356 8903 413
rect 8876 307 8883 343
rect 8936 156 8943 173
rect 8976 156 8983 233
rect 8996 136 9003 673
rect 9036 387 9043 693
rect 9076 547 9083 813
rect 9116 687 9123 1153
rect 9256 1096 9263 1153
rect 9196 1063 9203 1083
rect 9196 1056 9223 1063
rect 9216 843 9223 1056
rect 9196 836 9223 843
rect 9176 816 9203 823
rect 9116 616 9123 673
rect 9176 636 9183 673
rect 9156 607 9163 623
rect 9196 527 9203 816
rect 9096 356 9103 513
rect 9016 147 9023 253
rect 9156 156 9163 353
rect 9216 327 9223 653
rect 9236 376 9243 573
rect 9256 507 9263 853
rect 9276 667 9283 1176
rect 9276 376 9283 633
rect 9216 187 9223 313
rect 9216 163 9223 173
rect 9196 156 9223 163
rect 9296 127 9303 1653
rect 9316 1607 9323 1763
rect 9316 1327 9323 1393
rect 9336 1347 9343 2033
rect 9356 1827 9363 2056
rect 9356 1627 9363 1773
rect 9376 1747 9383 2413
rect 9396 2407 9403 2753
rect 9436 2563 9443 3093
rect 9456 3067 9463 3223
rect 9416 2556 9443 2563
rect 9436 2447 9443 2473
rect 9456 2467 9463 2753
rect 9476 2607 9483 3703
rect 9496 3387 9503 4013
rect 9536 3996 9563 4003
rect 9596 3996 9603 4013
rect 9536 3947 9543 3996
rect 9616 3976 9643 3983
rect 9636 3747 9643 3976
rect 9536 3703 9543 3733
rect 9516 3696 9543 3703
rect 9656 3627 9663 4113
rect 9696 3987 9703 4033
rect 9716 3987 9723 4153
rect 9976 4127 9983 4183
rect 9996 4167 10003 4193
rect 10176 4187 10183 4203
rect 9756 3996 9763 4053
rect 9676 3647 9683 3703
rect 9656 3516 9663 3613
rect 9556 3167 9563 3233
rect 9556 3056 9563 3073
rect 9516 3036 9543 3043
rect 9576 3036 9583 3373
rect 9596 3047 9603 3503
rect 9636 3367 9643 3503
rect 9616 3183 9623 3243
rect 9656 3236 9663 3293
rect 9636 3203 9643 3223
rect 9636 3196 9663 3203
rect 9616 3176 9643 3183
rect 9516 3007 9523 3036
rect 9576 2743 9583 2793
rect 9556 2736 9583 2743
rect 9516 2687 9523 2723
rect 9456 2447 9463 2453
rect 9476 2347 9483 2593
rect 9496 2547 9503 2573
rect 9396 1963 9403 2333
rect 9416 2247 9423 2333
rect 9416 2067 9423 2133
rect 9436 2047 9443 2333
rect 9516 2323 9523 2613
rect 9596 2587 9603 2753
rect 9616 2707 9623 2733
rect 9636 2727 9643 3176
rect 9656 3167 9663 3196
rect 9576 2527 9583 2543
rect 9516 2316 9543 2323
rect 9456 2267 9463 2283
rect 9476 2103 9483 2303
rect 9496 2127 9503 2283
rect 9476 2096 9503 2103
rect 9496 2076 9503 2096
rect 9536 2087 9543 2316
rect 9476 2047 9483 2063
rect 9396 1956 9423 1963
rect 9396 1787 9403 1933
rect 9376 1616 9383 1653
rect 9356 1596 9363 1613
rect 9416 1587 9423 1956
rect 9476 1867 9483 2033
rect 9356 1316 9363 1333
rect 9316 687 9323 1213
rect 9336 967 9343 1303
rect 9376 967 9383 1303
rect 9396 1116 9403 1253
rect 9416 1187 9423 1533
rect 9436 1187 9443 1853
rect 9496 1816 9503 1993
rect 9556 1987 9563 2273
rect 9576 2267 9583 2513
rect 9616 2287 9623 2693
rect 9416 1136 9423 1173
rect 9456 1167 9463 1733
rect 9516 1347 9523 1853
rect 9536 1367 9543 1873
rect 9556 1627 9563 1853
rect 9576 1687 9583 2053
rect 9596 1787 9603 2253
rect 9636 2243 9643 2553
rect 9656 2427 9663 2913
rect 9676 2667 9683 3223
rect 9696 3207 9703 3293
rect 9716 3187 9723 3973
rect 9736 3927 9743 3993
rect 9816 3976 9823 4073
rect 9996 4007 10003 4153
rect 10116 4087 10123 4183
rect 10156 4047 10163 4183
rect 9736 3187 9743 3703
rect 9756 3447 9763 3493
rect 9776 3483 9783 3933
rect 9776 3476 9803 3483
rect 9836 3287 9843 3433
rect 9776 3236 9803 3243
rect 9836 3236 9843 3273
rect 9856 3263 9863 3993
rect 9996 3976 10003 3993
rect 10036 3963 10043 3993
rect 10196 3976 10203 4213
rect 10316 4107 10323 4183
rect 10356 4007 10363 4183
rect 10496 4183 10503 4233
rect 10476 4176 10503 4183
rect 10236 3976 10243 3993
rect 10336 3976 10363 3983
rect 10396 3976 10403 4013
rect 10016 3956 10043 3963
rect 9876 3707 9883 3723
rect 9936 3687 9943 3703
rect 9956 3687 9963 3933
rect 10036 3747 10043 3933
rect 9896 3487 9903 3653
rect 9976 3547 9983 3713
rect 9856 3256 9883 3263
rect 9696 3027 9703 3073
rect 9776 3036 9783 3236
rect 9816 3167 9823 3203
rect 9716 2927 9723 3023
rect 9716 2767 9723 2913
rect 9696 2727 9703 2743
rect 9676 2407 9683 2593
rect 9696 2527 9703 2713
rect 9716 2707 9723 2723
rect 9756 2707 9763 2753
rect 9676 2276 9683 2393
rect 9716 2347 9723 2573
rect 9736 2556 9743 2613
rect 9776 2556 9783 2773
rect 9796 2707 9803 2973
rect 9836 2807 9843 3153
rect 9756 2527 9763 2543
rect 9796 2536 9823 2543
rect 9636 2236 9663 2243
rect 9616 1867 9623 2113
rect 9636 1967 9643 2073
rect 9656 2007 9663 2236
rect 9696 2167 9703 2263
rect 9696 2076 9703 2113
rect 9736 2076 9743 2393
rect 9716 1987 9723 2063
rect 9636 1807 9643 1823
rect 9616 1747 9623 1803
rect 9596 1596 9603 1653
rect 9616 1567 9623 1583
rect 9656 1447 9663 1773
rect 9516 1267 9523 1313
rect 9556 1247 9563 1323
rect 9596 1316 9603 1353
rect 9576 1283 9583 1303
rect 9576 1276 9603 1283
rect 9596 1127 9603 1276
rect 9676 1127 9683 1753
rect 9696 1727 9703 1953
rect 9696 1167 9703 1613
rect 9716 1547 9723 1973
rect 9736 1587 9743 1993
rect 9756 1967 9763 2513
rect 9816 2487 9823 2536
rect 9776 2087 9783 2333
rect 9816 2327 9823 2473
rect 9796 2087 9803 2153
rect 9776 2047 9783 2073
rect 9756 1807 9763 1893
rect 9756 1627 9763 1773
rect 9776 1767 9783 1993
rect 9796 1947 9803 2053
rect 9816 1967 9823 2253
rect 9836 2047 9843 2533
rect 9856 2287 9863 3173
rect 9876 2547 9883 3256
rect 9896 3227 9903 3273
rect 9896 2807 9903 3013
rect 9916 2787 9923 3533
rect 9956 3516 9983 3523
rect 10016 3516 10023 3553
rect 9956 3167 9963 3516
rect 10036 3496 10043 3733
rect 10056 3687 10063 3703
rect 10056 3487 10063 3673
rect 10096 3667 10103 3703
rect 10116 3547 10123 3723
rect 9996 3247 10003 3333
rect 10036 3236 10043 3413
rect 9996 3047 10003 3233
rect 10016 3147 10023 3223
rect 9996 3016 10003 3033
rect 9936 2987 9943 3003
rect 9976 2996 9983 3013
rect 9927 2776 9943 2783
rect 9896 2723 9903 2763
rect 9936 2756 9943 2776
rect 9976 2767 9983 2793
rect 9896 2716 9923 2723
rect 9916 2707 9923 2716
rect 9896 2307 9903 2693
rect 9916 2447 9923 2673
rect 9936 2547 9943 2713
rect 9956 2556 9963 2693
rect 9996 2576 10003 2733
rect 10016 2647 10023 3053
rect 9896 2276 9903 2293
rect 9976 2247 9983 2333
rect 9916 2167 9923 2243
rect 9876 2096 9883 2113
rect 9856 2047 9863 2063
rect 9936 2047 9943 2113
rect 9796 1616 9803 1893
rect 9896 1803 9903 2033
rect 9936 1907 9943 2033
rect 9956 2007 9963 2073
rect 9976 2067 9983 2213
rect 9996 2187 10003 2233
rect 9876 1796 9903 1803
rect 9816 1767 9823 1783
rect 9756 1583 9763 1593
rect 9756 1576 9783 1583
rect 9756 1527 9763 1576
rect 9716 1307 9723 1433
rect 9727 1296 9743 1303
rect 9756 1227 9763 1283
rect 9776 1247 9783 1303
rect 9436 1116 9463 1123
rect 9456 1067 9463 1116
rect 9596 1096 9623 1103
rect 9356 667 9363 843
rect 9396 836 9403 853
rect 9416 647 9423 823
rect 9436 707 9443 953
rect 9456 747 9463 1053
rect 9476 907 9483 953
rect 9476 667 9483 893
rect 9536 843 9543 1073
rect 9516 836 9543 843
rect 9576 1036 9593 1043
rect 9516 667 9523 836
rect 9576 807 9583 1036
rect 9616 967 9623 1096
rect 9636 823 9643 1113
rect 9676 1087 9683 1113
rect 9696 1087 9703 1133
rect 9616 816 9643 823
rect 9416 607 9423 633
rect 9476 623 9483 653
rect 9476 616 9503 623
rect 9536 603 9543 623
rect 9536 596 9563 603
rect 9556 587 9563 596
rect 9436 376 9443 453
rect 9476 227 9483 383
rect 9516 363 9523 533
rect 9496 356 9523 363
rect 9556 227 9563 573
rect 9576 367 9583 653
rect 9596 627 9603 653
rect 9356 156 9363 213
rect 9516 156 9523 173
rect 9556 156 9563 213
rect 9576 147 9583 353
rect 9596 343 9603 593
rect 9636 356 9643 793
rect 9656 587 9663 833
rect 9676 403 9683 1013
rect 9736 807 9743 1173
rect 9776 1096 9783 1153
rect 9756 1067 9763 1083
rect 9796 1076 9803 1113
rect 9816 1096 9823 1113
rect 9836 907 9843 1613
rect 9856 1147 9863 1713
rect 9756 636 9763 893
rect 9796 847 9803 853
rect 9876 823 9883 1653
rect 9916 1596 9923 1693
rect 9956 1596 9963 1893
rect 9976 1567 9983 1853
rect 9996 1803 10003 2173
rect 10016 2007 10023 2543
rect 10036 2167 10043 2973
rect 10056 2367 10063 2993
rect 10096 2867 10103 3133
rect 10116 3067 10123 3513
rect 10136 3167 10143 3673
rect 10156 3667 10163 3953
rect 10176 3907 10183 3963
rect 10216 3956 10223 3973
rect 10336 3947 10343 3976
rect 10336 3927 10343 3933
rect 10356 3907 10363 3933
rect 10196 3516 10203 3733
rect 10316 3727 10323 3743
rect 10296 3707 10303 3723
rect 10336 3667 10343 3723
rect 10236 3516 10243 3593
rect 10276 3516 10283 3553
rect 10176 3367 10183 3473
rect 10156 3327 10163 3353
rect 10176 3003 10183 3353
rect 10216 3287 10223 3503
rect 10256 3447 10263 3503
rect 10116 2983 10123 3003
rect 10156 2996 10183 3003
rect 10196 3256 10223 3263
rect 10256 3256 10263 3393
rect 10116 2976 10143 2983
rect 10136 2907 10143 2976
rect 10096 2743 10103 2853
rect 10136 2743 10143 2893
rect 10156 2747 10163 2996
rect 10076 2736 10103 2743
rect 10116 2736 10143 2743
rect 10076 2407 10083 2736
rect 10116 2727 10123 2736
rect 10056 2327 10063 2353
rect 10016 1847 10023 1993
rect 10056 1987 10063 2293
rect 10116 2287 10123 2573
rect 10176 2556 10183 2953
rect 10196 2627 10203 3256
rect 10216 2587 10223 3153
rect 10256 2767 10263 3053
rect 10276 2907 10283 3273
rect 10296 3267 10303 3633
rect 10336 3347 10343 3653
rect 10296 3167 10303 3253
rect 10336 3207 10343 3253
rect 10296 3036 10303 3073
rect 10356 3067 10363 3893
rect 10456 3743 10463 4173
rect 10656 4127 10663 4183
rect 10696 4167 10703 4183
rect 10436 3736 10463 3743
rect 10436 3703 10443 3736
rect 10536 3727 10543 4033
rect 10576 4007 10583 4093
rect 10656 4047 10663 4073
rect 10696 4067 10703 4153
rect 10596 3996 10603 4033
rect 10636 3996 10643 4013
rect 10576 3976 10583 3993
rect 10436 3696 10463 3703
rect 10476 3647 10483 3683
rect 10456 3547 10463 3613
rect 10496 3503 10503 3533
rect 10436 3347 10443 3503
rect 10476 3496 10503 3503
rect 10376 3256 10383 3273
rect 10416 3256 10443 3263
rect 10396 3207 10403 3243
rect 10436 3207 10443 3256
rect 10316 3007 10323 3023
rect 10296 2743 10303 2773
rect 10276 2736 10303 2743
rect 10276 2607 10283 2736
rect 10216 2556 10243 2563
rect 10156 2523 10163 2543
rect 10156 2516 10183 2523
rect 10136 2276 10143 2353
rect 10116 2227 10123 2243
rect 10076 2076 10103 2083
rect 10116 2076 10143 2083
rect 10096 1947 10103 2076
rect 10136 2027 10143 2076
rect 9996 1796 10023 1803
rect 10056 1787 10063 1803
rect 9916 1307 9923 1493
rect 9936 1207 9943 1323
rect 10016 1303 10023 1593
rect 10076 1343 10083 1713
rect 10096 1607 10103 1933
rect 10116 1727 10123 1973
rect 10116 1576 10123 1653
rect 10136 1543 10143 1553
rect 10116 1536 10143 1543
rect 10076 1336 10103 1343
rect 9996 1296 10023 1303
rect 10076 1287 10083 1313
rect 9696 607 9703 623
rect 9676 396 9703 403
rect 9596 336 9623 343
rect 9696 247 9703 396
rect 9696 156 9703 233
rect 9736 156 9743 373
rect 9776 367 9783 633
rect 9816 587 9823 823
rect 9856 816 9883 823
rect 9856 567 9863 713
rect 9876 407 9883 613
rect 9876 356 9883 393
rect 9896 387 9903 1193
rect 10036 1167 10043 1233
rect 10007 1136 10013 1143
rect 9936 1107 9943 1113
rect 9956 1096 9963 1133
rect 9976 1116 9983 1133
rect 10036 1123 10043 1153
rect 10016 1116 10043 1123
rect 9916 787 9923 893
rect 9936 727 9943 873
rect 9976 836 9983 1053
rect 9996 847 10003 1103
rect 10036 1067 10043 1093
rect 10016 836 10023 853
rect 9936 636 9943 653
rect 9976 636 9983 733
rect 9916 616 9923 633
rect 9996 627 10003 673
rect 10016 356 10023 513
rect 10056 367 10063 653
rect 10076 647 10083 1173
rect 10096 667 10103 1336
rect 10116 1227 10123 1536
rect 10156 1387 10163 2273
rect 10176 1567 10183 2516
rect 10196 2047 10203 2293
rect 10216 2267 10223 2313
rect 10216 2127 10223 2233
rect 10236 2167 10243 2556
rect 10256 2507 10263 2553
rect 10276 2387 10283 2573
rect 10296 2467 10303 2553
rect 10316 2467 10323 2753
rect 10336 2547 10343 2853
rect 10356 2847 10363 3023
rect 10396 2647 10403 3153
rect 10436 2927 10443 3033
rect 10456 3003 10463 3333
rect 10516 3267 10523 3513
rect 10536 3507 10543 3593
rect 10556 3507 10563 3913
rect 10656 3843 10663 4033
rect 10696 3887 10703 3993
rect 10636 3836 10663 3843
rect 10636 3723 10643 3836
rect 10636 3716 10663 3723
rect 10696 3716 10703 3753
rect 10636 3707 10643 3716
rect 10676 3683 10683 3703
rect 10676 3676 10703 3683
rect 10576 3516 10603 3523
rect 10636 3516 10643 3553
rect 10576 3267 10583 3516
rect 10476 3027 10483 3173
rect 10536 3036 10543 3253
rect 10616 3236 10623 3453
rect 10696 3423 10703 3676
rect 10716 3567 10723 3703
rect 10696 3416 10723 3423
rect 10556 3087 10563 3223
rect 10596 3207 10603 3223
rect 10636 3207 10643 3223
rect 10596 3067 10603 3193
rect 10456 2996 10483 3003
rect 10416 2736 10443 2743
rect 10376 2536 10383 2573
rect 10336 2523 10343 2533
rect 10416 2523 10423 2593
rect 10336 2516 10363 2523
rect 10396 2516 10423 2523
rect 10436 2503 10443 2736
rect 10416 2496 10443 2503
rect 10276 2276 10283 2373
rect 10296 2327 10303 2453
rect 10316 2247 10323 2283
rect 10196 1783 10203 1953
rect 10216 1907 10223 2113
rect 10236 1887 10243 2153
rect 10256 2056 10263 2213
rect 10276 2076 10283 2133
rect 10296 2047 10303 2063
rect 10236 1796 10243 1813
rect 10336 1787 10343 2393
rect 10196 1776 10223 1783
rect 10256 1647 10263 1783
rect 10296 1727 10303 1783
rect 10356 1627 10363 2273
rect 10376 1847 10383 2413
rect 10256 1616 10283 1623
rect 10196 1447 10203 1553
rect 10256 1467 10263 1616
rect 10196 1303 10203 1433
rect 10216 1307 10223 1433
rect 10176 1296 10203 1303
rect 10116 667 10123 1213
rect 10136 1116 10183 1123
rect 10216 1116 10243 1123
rect 10136 1107 10143 1116
rect 10196 867 10203 1103
rect 10236 1027 10243 1116
rect 10276 1047 10283 1513
rect 10296 1287 10303 1303
rect 10356 1247 10363 1313
rect 10196 836 10203 853
rect 10236 803 10243 993
rect 10216 796 10243 803
rect 10256 767 10263 833
rect 10156 616 10163 653
rect 10176 567 10183 633
rect 10116 367 10123 393
rect 9856 287 9863 343
rect 9896 307 9903 343
rect 9876 176 9883 253
rect 9376 127 9383 143
rect 9916 143 9923 193
rect 9996 147 10003 353
rect 10016 303 10023 313
rect 10016 296 10043 303
rect 10036 156 10043 296
rect 10076 287 10083 343
rect 10076 156 10083 173
rect 10136 147 10143 273
rect 10216 267 10223 633
rect 10236 376 10243 693
rect 10256 687 10263 753
rect 10256 627 10263 673
rect 10276 403 10283 1033
rect 10296 827 10303 1233
rect 10396 1187 10403 2493
rect 10416 2027 10423 2496
rect 10456 2447 10463 2653
rect 10476 2507 10483 2996
rect 10436 2147 10443 2313
rect 10456 2103 10463 2433
rect 10496 2307 10503 2573
rect 10516 2287 10523 2993
rect 10556 2587 10563 3023
rect 10596 3007 10603 3033
rect 10636 2907 10643 3193
rect 10596 2747 10603 2813
rect 10656 2776 10663 2813
rect 10636 2687 10643 2763
rect 10576 2576 10583 2673
rect 10596 2527 10603 2543
rect 10556 2407 10563 2513
rect 10536 2276 10543 2313
rect 10436 2096 10463 2103
rect 10476 2087 10483 2263
rect 10496 1823 10503 2133
rect 10476 1816 10503 1823
rect 10456 1767 10463 1783
rect 10456 1616 10463 1633
rect 10416 1596 10443 1603
rect 10476 1596 10483 1816
rect 10496 1767 10503 1773
rect 10416 1307 10423 1596
rect 10496 1587 10503 1633
rect 10436 1147 10443 1373
rect 10456 1327 10463 1393
rect 10516 1387 10523 1833
rect 10536 1507 10543 2073
rect 10556 2067 10563 2393
rect 10596 2083 10603 2293
rect 10616 2107 10623 2633
rect 10636 2527 10643 2553
rect 10656 2267 10663 2333
rect 10676 2327 10683 3053
rect 10696 2547 10703 3073
rect 10716 3016 10723 3416
rect 10736 3167 10743 4233
rect 10756 3996 10763 4033
rect 10756 3187 10763 3953
rect 10796 3507 10803 3853
rect 10816 3527 10823 4093
rect 10836 3667 10843 4193
rect 10856 3987 10863 4183
rect 10996 4016 11003 4093
rect 10936 3996 10963 4003
rect 10936 3867 10943 3996
rect 10976 3927 10983 3983
rect 11036 3807 11043 6353
rect 11096 6327 11103 7033
rect 11116 6567 11123 6813
rect 11136 6596 11143 6913
rect 11176 6596 11183 6893
rect 11296 6767 11303 7093
rect 11376 7067 11383 7083
rect 11336 6876 11343 6913
rect 11376 6876 11383 6893
rect 11316 6607 11323 6873
rect 11396 6867 11403 6873
rect 11356 6827 11363 6863
rect 11416 6647 11423 7596
rect 11456 7527 11463 7543
rect 11196 6427 11203 6583
rect 11156 6396 11183 6403
rect 11156 6347 11163 6396
rect 11236 6376 11243 6433
rect 11356 6407 11363 6593
rect 11416 6547 11423 6553
rect 11096 6116 11103 6153
rect 11076 6087 11083 6103
rect 11096 5947 11103 5993
rect 11136 5947 11143 6113
rect 11156 6107 11163 6133
rect 11356 6127 11363 6393
rect 11296 6087 11303 6103
rect 11096 5896 11103 5933
rect 11156 5916 11163 6073
rect 11176 5907 11183 6013
rect 11136 5636 11163 5643
rect 11076 5603 11083 5633
rect 11076 5596 11103 5603
rect 11096 5167 11103 5473
rect 11136 5467 11143 5636
rect 11196 5627 11203 5933
rect 11256 5903 11263 6073
rect 11356 6047 11363 6113
rect 11296 5936 11303 6013
rect 11256 5896 11283 5903
rect 11376 5663 11383 6433
rect 11416 6427 11423 6533
rect 11436 6423 11443 7353
rect 11456 7336 11463 7373
rect 11476 7367 11483 8536
rect 11576 8523 11583 8793
rect 11556 8516 11583 8523
rect 11536 8483 11543 8503
rect 11516 8476 11543 8483
rect 11496 8327 11503 8433
rect 11516 7987 11523 8476
rect 11596 8403 11603 8933
rect 11616 8796 11623 8833
rect 11596 8396 11623 8403
rect 11556 8316 11583 8323
rect 11596 8316 11603 8373
rect 11576 8067 11583 8316
rect 11556 7996 11583 8003
rect 11516 7836 11523 7853
rect 11556 7843 11563 7973
rect 11576 7907 11583 7996
rect 11556 7836 11583 7843
rect 11496 7807 11503 7833
rect 11536 7327 11543 7773
rect 11556 7567 11563 7836
rect 11576 7563 11583 7793
rect 11616 7627 11623 8396
rect 11636 8027 11643 8593
rect 11656 8047 11663 8633
rect 11676 8407 11683 9873
rect 11696 9727 11703 9753
rect 11716 9667 11723 9913
rect 11736 9767 11743 9933
rect 11756 9807 11763 10013
rect 11736 9627 11743 9733
rect 11816 9703 11823 10173
rect 11796 9696 11823 9703
rect 11696 9307 11703 9493
rect 11756 9447 11763 9513
rect 11696 9287 11703 9293
rect 11776 9267 11783 9473
rect 11796 9467 11803 9696
rect 11816 9287 11823 9613
rect 11776 9027 11783 9253
rect 11796 9207 11803 9263
rect 11716 8947 11723 8983
rect 11716 8867 11723 8933
rect 11736 8907 11743 8963
rect 11756 8907 11763 8973
rect 11796 8887 11803 9193
rect 11816 8967 11823 9273
rect 11716 8667 11723 8813
rect 11736 8547 11743 8873
rect 11756 8807 11763 8853
rect 11776 8796 11783 8833
rect 11796 8816 11803 8853
rect 11756 8483 11763 8793
rect 11776 8507 11783 8613
rect 11716 8427 11723 8483
rect 11736 8476 11763 8483
rect 11676 8107 11683 8333
rect 11716 8147 11723 8333
rect 11736 8316 11743 8476
rect 11776 8327 11783 8493
rect 11736 8056 11743 8253
rect 11716 7823 11723 8033
rect 11696 7816 11723 7823
rect 11736 7816 11743 7893
rect 11576 7556 11603 7563
rect 11616 7547 11623 7583
rect 11656 7576 11663 7633
rect 11616 7327 11623 7533
rect 11676 7383 11683 7613
rect 11736 7547 11743 7773
rect 11656 7376 11683 7383
rect 11516 7067 11523 7323
rect 11536 7096 11543 7273
rect 11576 7096 11603 7103
rect 11596 7047 11603 7096
rect 11536 6896 11543 6913
rect 11576 6863 11583 6933
rect 11556 6856 11583 6863
rect 11456 6527 11463 6593
rect 11436 6416 11463 6423
rect 11356 5656 11383 5663
rect 11156 5436 11163 5453
rect 11176 5407 11183 5423
rect 11216 5187 11223 5433
rect 11096 4987 11103 5153
rect 11116 5027 11123 5163
rect 11136 5047 11143 5143
rect 11176 5127 11183 5143
rect 11096 4947 11103 4973
rect 11136 4956 11143 5013
rect 11196 4943 11203 5033
rect 11196 4936 11223 4943
rect 11056 4696 11083 4703
rect 11116 4696 11143 4703
rect 11056 4687 11063 4696
rect 11056 4467 11063 4673
rect 11096 4587 11103 4683
rect 11136 4667 11143 4696
rect 11216 4687 11223 4936
rect 11236 4663 11243 4953
rect 11256 4703 11263 5453
rect 11336 5436 11343 5643
rect 11376 5467 11383 5656
rect 11396 5416 11403 5433
rect 11276 5267 11283 5413
rect 11276 5167 11283 5253
rect 11336 5176 11363 5183
rect 11356 5147 11363 5176
rect 11376 4976 11383 5173
rect 11356 4767 11363 4943
rect 11276 4703 11283 4713
rect 11256 4696 11283 4703
rect 11276 4676 11283 4696
rect 11236 4656 11263 4663
rect 11236 4627 11243 4656
rect 11136 4467 11143 4553
rect 11316 4487 11323 4673
rect 11216 4447 11223 4453
rect 11336 4443 11343 4573
rect 11356 4567 11363 4753
rect 11396 4647 11403 4973
rect 11336 4436 11363 4443
rect 11096 4207 11103 4223
rect 10896 3716 10903 3733
rect 10856 3647 10863 3713
rect 10876 3627 10883 3703
rect 10856 3516 10883 3523
rect 10876 3507 10883 3516
rect 10736 3036 10743 3113
rect 10776 3087 10783 3273
rect 10876 3227 10883 3493
rect 10896 3367 10903 3653
rect 10916 3407 10923 3513
rect 10776 3036 10783 3073
rect 10796 3047 10803 3223
rect 10836 3147 10843 3223
rect 10756 3007 10763 3023
rect 10736 2647 10743 2773
rect 10756 2667 10763 2973
rect 10796 2807 10803 3033
rect 10776 2796 10793 2803
rect 10776 2763 10783 2796
rect 10836 2767 10843 3113
rect 10916 3087 10923 3393
rect 10936 3127 10943 3573
rect 11016 3567 11023 3733
rect 11016 3536 11023 3553
rect 10996 3327 11003 3503
rect 11036 3367 11043 3503
rect 11076 3387 11083 4193
rect 11116 4167 11123 4203
rect 11116 3707 11123 4153
rect 11156 3983 11163 4213
rect 11256 4047 11263 4193
rect 11276 4187 11283 4223
rect 11276 4127 11283 4173
rect 11256 4007 11263 4033
rect 11136 3976 11163 3983
rect 11136 3967 11143 3976
rect 11096 3667 11103 3703
rect 11256 3703 11263 3993
rect 11236 3696 11263 3703
rect 11276 3687 11283 3703
rect 10956 3256 10963 3293
rect 10996 3256 11023 3263
rect 10976 3047 10983 3243
rect 10936 3016 10943 3033
rect 10876 2827 10883 2893
rect 10776 2756 10803 2763
rect 10876 2743 10883 2813
rect 10996 2783 11003 3153
rect 11016 3047 11023 3256
rect 11016 2867 11023 3033
rect 11036 2803 11043 3273
rect 11096 3127 11103 3653
rect 11276 3516 11283 3573
rect 11196 3467 11203 3513
rect 11176 3236 11183 3273
rect 10976 2776 11003 2783
rect 11016 2796 11043 2803
rect 10776 2587 10783 2593
rect 10736 2536 10743 2553
rect 10776 2536 10783 2573
rect 10676 2187 10683 2283
rect 10596 2076 10623 2083
rect 10656 2076 10663 2153
rect 10576 2056 10603 2063
rect 10556 1427 10563 2053
rect 10336 1116 10363 1123
rect 10396 1116 10403 1133
rect 10336 1107 10343 1116
rect 10316 823 10323 973
rect 10316 816 10343 823
rect 10296 636 10303 733
rect 10356 647 10363 933
rect 10356 616 10363 633
rect 10376 427 10383 813
rect 10476 627 10483 1373
rect 10536 1336 10563 1343
rect 10556 1307 10563 1336
rect 10576 1227 10583 2056
rect 10576 1207 10583 1213
rect 10536 1116 10543 1153
rect 10576 1116 10583 1133
rect 10516 823 10523 1093
rect 10596 827 10603 2013
rect 10636 1623 10643 1783
rect 10676 1723 10683 1993
rect 10696 1827 10703 2093
rect 10756 2023 10763 2353
rect 10736 2016 10763 2023
rect 10716 1796 10723 1833
rect 10696 1747 10703 1783
rect 10676 1716 10703 1723
rect 10636 1616 10663 1623
rect 10616 1596 10623 1613
rect 10656 1596 10663 1616
rect 10676 1576 10683 1613
rect 10516 816 10543 823
rect 10576 816 10593 823
rect 10536 727 10543 816
rect 10516 636 10523 713
rect 10556 656 10563 693
rect 10616 627 10623 1493
rect 10636 1147 10643 1373
rect 10636 947 10643 1133
rect 10656 807 10663 1453
rect 10696 1316 10703 1716
rect 10736 1527 10743 2016
rect 10736 1307 10743 1323
rect 10676 1287 10683 1303
rect 10676 667 10683 1273
rect 10716 1127 10723 1233
rect 10716 1096 10723 1113
rect 10696 1067 10703 1083
rect 10696 1007 10703 1053
rect 10736 1047 10743 1083
rect 10696 687 10703 913
rect 10736 836 10743 1013
rect 10776 927 10783 2493
rect 10816 2307 10823 2743
rect 10856 2736 10883 2743
rect 10836 2527 10843 2693
rect 10896 2563 10903 2753
rect 10876 2556 10903 2563
rect 10856 2487 10863 2533
rect 10876 2523 10883 2556
rect 10956 2523 10963 2573
rect 10876 2516 10903 2523
rect 10936 2516 10963 2523
rect 10856 2327 10863 2473
rect 10896 2307 10903 2516
rect 10916 2276 10923 2473
rect 10836 2187 10843 2273
rect 10936 2243 10943 2273
rect 10896 2227 10903 2243
rect 10916 2236 10943 2243
rect 10896 2107 10903 2213
rect 10916 2127 10923 2236
rect 10796 1807 10803 2063
rect 10816 1596 10823 2053
rect 10836 1347 10843 2053
rect 10856 1816 10863 1913
rect 10916 1847 10923 2113
rect 10896 1807 10903 1823
rect 10876 1623 10883 1793
rect 10916 1667 10923 1803
rect 10876 1616 10903 1623
rect 10856 1596 10883 1603
rect 10876 1567 10883 1596
rect 10896 1316 10903 1616
rect 10936 1387 10943 2113
rect 10956 2067 10963 2133
rect 10976 2107 10983 2776
rect 11016 2756 11023 2796
rect 11056 2767 11063 3013
rect 11076 2967 11083 3073
rect 11096 3023 11103 3053
rect 11096 3016 11123 3023
rect 11076 2867 11083 2933
rect 10996 2687 11003 2743
rect 11076 2727 11083 2853
rect 10996 2107 11003 2633
rect 11016 2207 11023 2253
rect 11016 2076 11023 2193
rect 11036 2067 11043 2673
rect 11076 2556 11083 2633
rect 11096 2587 11103 2813
rect 11116 2587 11123 2753
rect 11136 2607 11143 3113
rect 11156 3036 11163 3073
rect 11196 2987 11203 3223
rect 11156 2743 11163 2953
rect 11216 2787 11223 3373
rect 11156 2736 11183 2743
rect 11216 2627 11223 2733
rect 11156 2556 11163 2613
rect 11096 2527 11103 2543
rect 11096 2367 11103 2513
rect 11136 2447 11143 2543
rect 11116 2276 11123 2293
rect 11096 2207 11103 2243
rect 11096 2167 11103 2193
rect 11156 2103 11163 2213
rect 11176 2127 11183 2593
rect 11156 2096 11183 2103
rect 11096 2067 11103 2093
rect 11116 2076 11143 2083
rect 11176 2076 11183 2096
rect 11196 2087 11203 2573
rect 11216 2447 11223 2573
rect 11236 2527 11243 3473
rect 11316 3467 11323 4013
rect 11336 3996 11343 4013
rect 11396 4007 11403 4193
rect 11396 3976 11403 3993
rect 11356 3567 11363 3973
rect 11416 3743 11423 6153
rect 11456 6143 11463 6416
rect 11476 6167 11483 6633
rect 11516 6596 11543 6603
rect 11576 6596 11583 6613
rect 11516 6587 11523 6596
rect 11516 6407 11523 6573
rect 11556 6527 11563 6563
rect 11516 6147 11523 6393
rect 11536 6367 11543 6453
rect 11436 6136 11463 6143
rect 11436 4227 11443 6136
rect 11476 6123 11483 6133
rect 11456 6116 11483 6123
rect 11476 6067 11483 6083
rect 11456 5407 11463 5973
rect 11476 5787 11483 6053
rect 11516 5987 11523 6103
rect 11496 5896 11503 5953
rect 11556 5947 11563 6413
rect 11616 6403 11623 6813
rect 11596 6396 11623 6403
rect 11596 6107 11603 6396
rect 11656 6147 11663 7376
rect 11736 7356 11743 7393
rect 11676 6347 11683 7213
rect 11756 7187 11763 7803
rect 11776 7227 11783 7873
rect 11796 7867 11803 8533
rect 11816 7787 11823 8753
rect 11836 7587 11843 10236
rect 11856 9287 11863 10333
rect 11876 10207 11883 10403
rect 11876 9976 11883 10193
rect 11896 10187 11903 10353
rect 11916 10147 11923 10373
rect 11936 10327 11943 10433
rect 11956 10387 11963 10813
rect 11936 10236 11943 10273
rect 11956 10256 11963 10293
rect 11976 10287 11983 10973
rect 11996 10347 12003 11033
rect 12016 10647 12023 10893
rect 12036 10727 12043 11373
rect 12056 11327 12063 11383
rect 12056 11227 12063 11253
rect 12056 11176 12063 11213
rect 12056 10827 12063 11133
rect 12076 10907 12083 11913
rect 12096 11676 12103 11793
rect 12116 11507 12123 11663
rect 12156 11656 12163 11693
rect 12116 11367 12123 11383
rect 12136 11223 12143 11413
rect 12116 11216 12143 11223
rect 12116 11007 12123 11216
rect 12056 10716 12083 10723
rect 12116 10716 12123 10993
rect 12136 10987 12143 11183
rect 12036 10467 12043 10693
rect 12056 10687 12063 10716
rect 12056 10487 12063 10673
rect 12096 10667 12103 10703
rect 12096 10443 12103 10473
rect 12076 10436 12103 10443
rect 11916 9976 11943 9983
rect 11896 9943 11903 9963
rect 11876 9936 11903 9943
rect 11876 9687 11883 9936
rect 11936 9927 11943 9976
rect 11896 9523 11903 9773
rect 11976 9747 11983 10153
rect 11996 9907 12003 10273
rect 12016 10267 12023 10423
rect 12116 10343 12123 10633
rect 12096 10336 12123 10343
rect 11996 9787 12003 9893
rect 11996 9767 12003 9773
rect 11876 9516 11903 9523
rect 11876 9507 11883 9516
rect 11916 9507 11923 9513
rect 11856 8547 11863 9273
rect 11876 8767 11883 9453
rect 11896 9447 11903 9483
rect 11896 9016 11903 9293
rect 11936 9227 11943 9673
rect 11976 9343 11983 9733
rect 11956 9336 11983 9343
rect 11896 8627 11903 8973
rect 11916 8847 11923 9003
rect 11956 8947 11963 9336
rect 11996 9296 12003 9413
rect 12016 9287 12023 10133
rect 12036 9947 12043 10253
rect 12096 10143 12103 10336
rect 12136 10267 12143 10593
rect 12156 10247 12163 11513
rect 12176 11267 12183 11653
rect 12176 10967 12183 11253
rect 12176 10587 12183 10913
rect 12156 10227 12163 10233
rect 12096 10136 12123 10143
rect 12116 9943 12123 10136
rect 12047 9936 12063 9943
rect 12096 9936 12123 9943
rect 12036 9463 12043 9933
rect 12056 9507 12063 9793
rect 12076 9707 12083 9913
rect 12096 9743 12103 9936
rect 12096 9736 12123 9743
rect 12096 9496 12103 9533
rect 12036 9456 12063 9463
rect 11936 8803 11943 8893
rect 11956 8816 11963 8913
rect 11916 8796 11943 8803
rect 11916 8567 11923 8796
rect 11996 8787 12003 9253
rect 11936 8503 11943 8533
rect 11956 8507 11963 8773
rect 11916 8496 11943 8503
rect 11876 8476 11903 8483
rect 11856 8267 11863 8473
rect 11876 8247 11883 8476
rect 11916 8347 11923 8393
rect 11956 8363 11963 8493
rect 11936 8356 11963 8363
rect 11936 8327 11943 8356
rect 11976 8347 11983 8553
rect 12016 8447 12023 9013
rect 12036 8987 12043 9433
rect 12056 9247 12063 9456
rect 12076 9387 12083 9483
rect 12116 9463 12123 9736
rect 12156 9727 12163 10213
rect 12096 9456 12123 9463
rect 12076 9083 12083 9273
rect 12096 9227 12103 9456
rect 12176 9287 12183 10573
rect 12056 9076 12083 9083
rect 12036 8527 12043 8953
rect 12056 8807 12063 9076
rect 12116 9027 12123 9273
rect 12176 9227 12183 9243
rect 12076 8967 12083 8983
rect 12096 8787 12103 8963
rect 12116 8847 12123 8983
rect 12116 8796 12123 8833
rect 12036 8503 12043 8513
rect 12116 8503 12123 8533
rect 12036 8496 12063 8503
rect 12096 8496 12123 8503
rect 11956 8307 11963 8333
rect 12056 8316 12063 8333
rect 11856 7807 11863 8093
rect 11876 8056 11883 8093
rect 11916 8056 11923 8293
rect 11896 8007 11903 8043
rect 11776 7063 11783 7193
rect 11756 7056 11783 7063
rect 11696 6876 11703 6913
rect 11796 6647 11803 7573
rect 11856 7556 11863 7793
rect 11896 7543 11903 7573
rect 11956 7567 11963 8293
rect 11976 7807 11983 7853
rect 11976 7567 11983 7653
rect 11996 7587 12003 7853
rect 12016 7807 12023 8053
rect 12036 8023 12043 8193
rect 12036 8016 12063 8023
rect 12056 7583 12063 7893
rect 12096 7867 12103 8013
rect 12116 7907 12123 8333
rect 12136 7927 12143 8773
rect 12096 7816 12103 7833
rect 12136 7803 12143 7913
rect 12116 7796 12143 7803
rect 12036 7576 12063 7583
rect 11876 7536 11903 7543
rect 11736 6567 11743 6583
rect 11796 6487 11803 6603
rect 11716 6363 11723 6373
rect 11796 6363 11803 6413
rect 11716 6356 11743 6363
rect 11776 6356 11803 6363
rect 11816 6347 11823 7533
rect 11876 7336 11883 7473
rect 11896 7356 11903 7393
rect 11936 7387 11943 7553
rect 11936 7356 11943 7373
rect 11876 7063 11883 7233
rect 11956 7063 11963 7453
rect 12016 7327 12023 7373
rect 12036 7323 12043 7473
rect 12056 7447 12063 7576
rect 12076 7487 12083 7793
rect 12056 7367 12063 7433
rect 12076 7336 12083 7453
rect 12036 7316 12063 7323
rect 11876 7056 11903 7063
rect 11936 7056 11963 7063
rect 11916 6903 11923 7043
rect 11896 6896 11923 6903
rect 11616 6087 11623 6133
rect 11636 6067 11643 6113
rect 11656 6087 11663 6103
rect 11716 6047 11723 6123
rect 11556 5916 11563 5933
rect 11516 5627 11523 5643
rect 11576 5627 11583 5713
rect 11596 5667 11603 5973
rect 11676 5916 11683 5953
rect 11716 5916 11723 5933
rect 11656 5587 11663 5913
rect 11736 5896 11743 5913
rect 11676 5656 11683 5693
rect 11716 5656 11723 5673
rect 11716 5456 11723 5573
rect 11456 4947 11463 5393
rect 11476 5187 11483 5453
rect 11596 5436 11623 5443
rect 11576 5407 11583 5423
rect 11496 5156 11503 5393
rect 11616 5367 11623 5436
rect 11556 5163 11563 5353
rect 11536 5156 11563 5163
rect 11476 5127 11483 5143
rect 11516 5007 11523 5143
rect 11536 4987 11543 5156
rect 11496 4956 11503 4973
rect 11556 4936 11563 4993
rect 11516 4703 11523 4933
rect 11616 4747 11623 5193
rect 11636 4947 11643 5413
rect 11656 5207 11663 5453
rect 11656 5176 11683 5183
rect 11716 5176 11723 5233
rect 11656 4967 11663 5176
rect 11496 4696 11523 4703
rect 11496 4663 11503 4696
rect 11476 4656 11503 4663
rect 11516 4456 11523 4473
rect 11536 4436 11543 4533
rect 11556 4456 11563 4513
rect 11616 4427 11623 4713
rect 11656 4676 11663 4933
rect 11676 4923 11683 4993
rect 11676 4916 11703 4923
rect 11736 4663 11743 4673
rect 11716 4656 11743 4663
rect 11676 4443 11683 4513
rect 11716 4456 11723 4493
rect 11676 4436 11703 4443
rect 11436 3987 11443 4183
rect 11476 4167 11483 4183
rect 11476 4147 11483 4153
rect 11396 3736 11423 3743
rect 11356 3507 11363 3553
rect 11256 3207 11263 3293
rect 11256 2507 11263 3133
rect 11276 2867 11283 3253
rect 11296 3047 11303 3153
rect 11316 3127 11323 3453
rect 11376 3347 11383 3513
rect 11396 3363 11403 3736
rect 11416 3587 11423 3703
rect 11456 3667 11463 3703
rect 11476 3667 11483 3993
rect 11476 3516 11483 3653
rect 11396 3356 11423 3363
rect 11396 3307 11403 3333
rect 11396 3223 11403 3293
rect 11376 3216 11403 3223
rect 11356 3187 11363 3203
rect 11336 3036 11343 3053
rect 11316 3007 11323 3023
rect 11356 3016 11363 3033
rect 11376 3027 11383 3113
rect 11276 2587 11283 2773
rect 11296 2587 11303 2993
rect 11316 2607 11323 2993
rect 11376 2907 11383 3013
rect 11396 2787 11403 3173
rect 11416 3047 11423 3356
rect 11416 2887 11423 3033
rect 11436 2987 11443 3473
rect 11456 3467 11463 3503
rect 11376 2707 11383 2763
rect 11416 2756 11423 2813
rect 11336 2556 11353 2563
rect 11276 2523 11283 2553
rect 11276 2516 11303 2523
rect 11116 2047 11123 2076
rect 10936 1316 10943 1333
rect 10916 1207 10923 1303
rect 10956 1223 10963 1303
rect 10976 1267 10983 1813
rect 10996 1543 11003 2033
rect 11076 1816 11083 1893
rect 11216 1867 11223 2413
rect 11236 2027 11243 2263
rect 11136 1707 11143 1833
rect 11256 1823 11263 2313
rect 11296 2267 11303 2516
rect 11316 2507 11323 2543
rect 11316 2287 11323 2493
rect 11276 2247 11283 2263
rect 11316 2247 11323 2273
rect 11236 1816 11263 1823
rect 11236 1796 11243 1816
rect 11036 1596 11043 1613
rect 11076 1596 11083 1673
rect 11016 1576 11023 1593
rect 10996 1536 11023 1543
rect 10936 1216 10963 1223
rect 10936 1123 10943 1216
rect 10856 1116 10883 1123
rect 10916 1116 10943 1123
rect 10856 867 10863 1116
rect 10896 1027 10903 1103
rect 10956 1007 10963 1193
rect 10776 836 10783 853
rect 10696 636 10703 673
rect 10736 636 10743 733
rect 10276 396 10303 403
rect 10296 183 10303 396
rect 10376 387 10383 413
rect 10456 356 10463 573
rect 10536 387 10543 613
rect 10536 347 10543 373
rect 10396 187 10403 343
rect 10476 327 10483 333
rect 10276 176 10303 183
rect 10276 156 10283 176
rect 10476 176 10483 213
rect 10436 156 10443 173
rect 9896 136 9923 143
rect 10296 127 10303 143
rect 10516 143 10523 173
rect 10536 147 10543 333
rect 10556 147 10563 433
rect 10576 367 10583 613
rect 10676 356 10683 393
rect 10616 207 10623 313
rect 10616 156 10623 193
rect 10656 156 10663 173
rect 10716 163 10723 433
rect 10796 347 10803 823
rect 10916 807 10923 993
rect 10956 836 10963 873
rect 10816 607 10823 713
rect 10876 636 10883 713
rect 10916 636 10923 693
rect 10936 667 10943 823
rect 10936 616 10943 633
rect 10956 607 10963 793
rect 10976 787 10983 823
rect 10816 347 10823 593
rect 10856 356 10863 373
rect 10896 356 10903 593
rect 10696 156 10723 163
rect 10816 147 10823 173
rect 10496 136 10523 143
rect 10836 143 10843 343
rect 10876 227 10883 323
rect 10976 287 10983 713
rect 10996 607 11003 833
rect 11016 727 11023 1536
rect 11036 647 11043 1313
rect 11056 847 11063 1273
rect 11076 1147 11083 1413
rect 11096 1303 11103 1593
rect 11136 1316 11143 1693
rect 11196 1596 11203 1773
rect 11256 1687 11263 1783
rect 11256 1576 11263 1593
rect 11296 1587 11303 2073
rect 11316 1787 11323 2233
rect 11336 2067 11343 2233
rect 11356 2227 11363 2453
rect 11356 2076 11363 2193
rect 11336 1607 11343 2053
rect 11356 1727 11363 2033
rect 11376 1827 11383 2693
rect 11416 2547 11423 2573
rect 11396 2167 11403 2533
rect 11436 2527 11443 2593
rect 11416 2463 11423 2513
rect 11416 2456 11443 2463
rect 11396 2076 11403 2113
rect 11396 1787 11403 1853
rect 11416 1847 11423 2433
rect 11436 2427 11443 2456
rect 11456 2307 11463 3033
rect 11476 2563 11483 3273
rect 11496 3047 11503 4213
rect 11516 3507 11523 4173
rect 11536 3487 11543 4393
rect 11556 3996 11563 4013
rect 11556 3507 11563 3693
rect 11576 3323 11583 3793
rect 11636 3716 11643 3953
rect 11656 3807 11663 4173
rect 11756 4163 11763 6333
rect 11776 4407 11783 6333
rect 11756 4156 11783 4163
rect 11676 3907 11683 3973
rect 11696 3956 11723 3963
rect 11656 3667 11663 3703
rect 11696 3667 11703 3956
rect 11596 3516 11603 3533
rect 11636 3516 11643 3593
rect 11676 3516 11683 3613
rect 11576 3316 11603 3323
rect 11516 3147 11523 3223
rect 11516 2996 11523 3073
rect 11576 3003 11583 3173
rect 11556 2996 11583 3003
rect 11496 2687 11503 2973
rect 11596 2927 11603 3316
rect 11516 2667 11523 2913
rect 11556 2787 11563 2833
rect 11636 2823 11643 3473
rect 11656 3187 11663 3503
rect 11716 3487 11723 3933
rect 11736 3467 11743 3573
rect 11756 3487 11763 3953
rect 11776 3947 11783 4156
rect 11796 3727 11803 6133
rect 11816 5707 11823 5933
rect 11816 4927 11823 5233
rect 11816 4907 11823 4913
rect 11816 4647 11823 4693
rect 11816 3967 11823 4173
rect 11796 3627 11803 3683
rect 11816 3567 11823 3703
rect 11756 3347 11763 3473
rect 11656 2843 11663 3153
rect 11676 3047 11683 3313
rect 11716 3256 11743 3263
rect 11716 3227 11723 3256
rect 11696 3207 11703 3223
rect 11736 3216 11763 3223
rect 11716 3187 11723 3213
rect 11736 3167 11743 3216
rect 11776 3207 11783 3533
rect 11836 3527 11843 6633
rect 11896 6447 11903 6896
rect 11936 6427 11943 6863
rect 11996 6627 12003 6863
rect 12076 6827 12083 7063
rect 12116 6927 12123 7063
rect 12096 6896 12123 6903
rect 11956 6587 11963 6603
rect 12036 6583 12043 6613
rect 12096 6607 12103 6896
rect 11856 6367 11863 6393
rect 11876 6143 11883 6373
rect 11856 6136 11883 6143
rect 11916 6136 11923 6333
rect 11856 6107 11863 6136
rect 11956 6127 11963 6573
rect 11976 6367 11983 6583
rect 12016 6576 12043 6583
rect 12016 6487 12023 6576
rect 11896 5987 11903 6123
rect 11916 5896 11923 6093
rect 11956 5896 11963 6113
rect 11896 5727 11903 5883
rect 11976 5707 11983 6133
rect 11876 5656 11883 5693
rect 12016 5687 12023 6393
rect 12096 6376 12103 6573
rect 12156 6396 12163 6563
rect 12176 6487 12183 6583
rect 12056 5947 12063 6143
rect 12076 6107 12083 6123
rect 12196 5963 12203 11813
rect 12176 5956 12203 5963
rect 12096 5887 12103 5903
rect 11856 4787 11863 5653
rect 11896 5467 11903 5643
rect 11936 5456 11943 5653
rect 12016 5487 12023 5673
rect 12036 5667 12043 5873
rect 12076 5656 12083 5673
rect 11876 5436 11903 5443
rect 11876 5247 11883 5436
rect 12016 5427 12023 5473
rect 12076 5436 12083 5473
rect 11916 5187 11923 5413
rect 12056 5203 12063 5433
rect 12096 5403 12103 5653
rect 12096 5396 12123 5403
rect 12056 5196 12083 5203
rect 11876 5047 11883 5163
rect 11956 5147 11963 5173
rect 12076 5167 12083 5196
rect 11936 5136 11953 5143
rect 11896 4927 11903 4943
rect 11916 4927 11923 5033
rect 11856 4707 11863 4773
rect 11876 4683 11883 4733
rect 11856 4676 11883 4683
rect 11896 4676 11903 4753
rect 12016 4707 12023 4933
rect 12076 4907 12083 4923
rect 12096 4696 12103 5143
rect 12116 4987 12123 5163
rect 11856 4443 11863 4613
rect 12056 4476 12083 4483
rect 11856 4436 11883 4443
rect 11916 4427 11923 4443
rect 11676 2867 11683 3033
rect 11716 3016 11723 3033
rect 11696 2987 11703 3003
rect 11756 2987 11763 3193
rect 11776 3067 11783 3093
rect 11656 2836 11683 2843
rect 11636 2816 11663 2823
rect 11536 2707 11543 2773
rect 11556 2743 11563 2773
rect 11636 2743 11643 2793
rect 11556 2736 11583 2743
rect 11616 2736 11643 2743
rect 11507 2576 11513 2583
rect 11476 2556 11503 2563
rect 11536 2556 11543 2573
rect 11556 2536 11563 2713
rect 11476 2487 11483 2533
rect 11496 2276 11503 2313
rect 11516 2247 11523 2263
rect 11536 2227 11543 2293
rect 11436 1867 11443 2153
rect 11456 1927 11463 2213
rect 11476 1867 11483 2193
rect 11416 1787 11423 1803
rect 11216 1363 11223 1573
rect 11196 1356 11223 1363
rect 11096 1296 11123 1303
rect 11196 1247 11203 1356
rect 11116 1147 11123 1173
rect 11076 1096 11083 1113
rect 11116 1096 11123 1133
rect 11136 1027 11143 1083
rect 11156 867 11163 1073
rect 11036 447 11043 633
rect 11056 627 11063 673
rect 11076 616 11083 653
rect 11096 627 11103 853
rect 11156 667 11163 823
rect 11116 636 11163 643
rect 11116 616 11123 636
rect 11096 596 11103 613
rect 10996 327 11003 353
rect 11096 347 11103 393
rect 11116 367 11123 413
rect 11156 407 11163 636
rect 11216 367 11223 1333
rect 11276 1307 11283 1353
rect 11256 1127 11263 1273
rect 11256 1083 11263 1113
rect 11296 1096 11303 1453
rect 11336 1316 11343 1593
rect 11356 1347 11363 1713
rect 11396 1576 11403 1713
rect 11376 1316 11383 1413
rect 11416 1287 11423 1553
rect 11436 1243 11443 1813
rect 11456 1787 11463 1803
rect 11416 1236 11443 1243
rect 11336 1083 11343 1233
rect 11416 1087 11423 1236
rect 11456 1227 11463 1773
rect 11496 1567 11503 2093
rect 11516 2076 11523 2213
rect 11536 2107 11543 2213
rect 11556 2207 11563 2313
rect 11556 2076 11563 2153
rect 11576 2127 11583 2653
rect 11596 2247 11603 2673
rect 11596 2076 11603 2093
rect 11536 2047 11543 2063
rect 11436 1116 11443 1133
rect 11476 1116 11483 1373
rect 11516 1347 11523 1833
rect 11536 1387 11543 1853
rect 11556 1447 11563 1913
rect 11596 1767 11603 1783
rect 11596 1576 11603 1633
rect 11616 1603 11623 2633
rect 11636 2287 11643 2713
rect 11656 2507 11663 2816
rect 11676 2667 11683 2836
rect 11676 2303 11683 2573
rect 11696 2327 11703 2853
rect 11716 2647 11723 2853
rect 11776 2827 11783 3053
rect 11736 2583 11743 2813
rect 11776 2756 11783 2793
rect 11796 2767 11803 3513
rect 11856 3467 11863 3483
rect 11816 2867 11823 3293
rect 11876 3207 11883 4153
rect 11896 3983 11903 3993
rect 11976 3983 11983 3993
rect 11896 3976 11923 3983
rect 11956 3976 11983 3983
rect 11896 3507 11903 3553
rect 11896 3267 11903 3493
rect 11896 3187 11903 3223
rect 11836 3007 11843 3173
rect 11876 3036 11883 3173
rect 11916 3067 11923 3976
rect 11996 3743 12003 4473
rect 12076 4247 12083 4476
rect 12016 4167 12023 4183
rect 12136 3996 12143 4233
rect 11976 3736 12003 3743
rect 11936 3267 11943 3713
rect 11956 3147 11963 3703
rect 11816 2756 11823 2773
rect 11756 2727 11763 2743
rect 11796 2707 11803 2723
rect 11736 2576 11763 2583
rect 11756 2556 11763 2576
rect 11676 2296 11703 2303
rect 11696 2276 11703 2296
rect 11636 2067 11643 2193
rect 11656 2027 11663 2253
rect 11716 2123 11723 2253
rect 11696 2116 11723 2123
rect 11696 1907 11703 2116
rect 11736 2103 11743 2553
rect 11756 2207 11763 2313
rect 11796 2267 11803 2693
rect 11816 2547 11823 2653
rect 11816 2267 11823 2333
rect 11716 2096 11743 2103
rect 11756 2096 11763 2153
rect 11656 1647 11663 1793
rect 11616 1596 11643 1603
rect 11556 1316 11563 1433
rect 11576 1327 11583 1563
rect 11496 1283 11503 1303
rect 11596 1287 11603 1313
rect 11496 1276 11523 1283
rect 11256 1076 11283 1083
rect 11316 1076 11343 1083
rect 11456 1047 11463 1103
rect 11496 1096 11503 1193
rect 11516 1107 11523 1276
rect 11536 1267 11543 1283
rect 11616 1247 11623 1553
rect 11636 1267 11643 1596
rect 11656 1567 11663 1613
rect 11676 1347 11683 1633
rect 11696 1607 11703 1773
rect 11696 1587 11703 1593
rect 11716 1343 11723 2096
rect 11796 2076 11803 2173
rect 11736 1787 11743 2063
rect 11776 1823 11783 2063
rect 11836 1847 11843 2753
rect 11856 2747 11863 2973
rect 11896 2847 11903 3023
rect 11936 3016 11943 3053
rect 11876 2727 11883 2773
rect 11896 2647 11903 2833
rect 11856 2567 11863 2633
rect 11896 2563 11903 2573
rect 11916 2563 11923 2873
rect 11976 2783 11983 3736
rect 11996 3667 12003 3703
rect 11996 3516 12003 3653
rect 12036 3527 12043 3873
rect 12056 3547 12063 3993
rect 12016 3487 12023 3503
rect 12056 3496 12063 3533
rect 12076 3307 12083 3513
rect 12096 3287 12103 3693
rect 12176 3687 12183 5956
rect 12196 3687 12203 3703
rect 11976 2776 12003 2783
rect 11896 2556 11923 2563
rect 11916 2536 11943 2543
rect 11936 2507 11943 2536
rect 11976 2507 11983 2743
rect 11916 2247 11923 2263
rect 11756 1816 11783 1823
rect 11756 1767 11763 1816
rect 11816 1767 11823 1783
rect 11836 1707 11843 1803
rect 11756 1616 11763 1633
rect 11736 1567 11743 1583
rect 11716 1336 11743 1343
rect 11336 836 11343 933
rect 11456 847 11463 1033
rect 11356 836 11383 843
rect 11356 747 11363 836
rect 11256 387 11263 653
rect 11296 587 11303 603
rect 11256 356 11263 373
rect 11296 356 11303 393
rect 10916 156 10923 213
rect 10836 136 10863 143
rect 11056 136 11063 273
rect 11116 156 11123 353
rect 11136 127 11143 353
rect 11236 307 11243 343
rect 11216 147 11223 193
rect 11336 187 11343 593
rect 11356 587 11363 653
rect 11376 607 11383 633
rect 11376 327 11383 573
rect 11396 343 11403 733
rect 11456 587 11463 833
rect 11476 823 11483 933
rect 11476 816 11503 823
rect 11536 727 11543 823
rect 11476 616 11483 713
rect 11496 636 11503 673
rect 11536 636 11543 653
rect 11516 587 11523 623
rect 11436 356 11443 373
rect 11576 347 11583 1193
rect 11636 1096 11643 1113
rect 11656 1107 11663 1313
rect 11676 1127 11683 1293
rect 11716 1267 11723 1303
rect 11736 1123 11743 1336
rect 11716 1116 11743 1123
rect 11616 627 11623 1093
rect 11716 883 11723 1116
rect 11736 1047 11743 1093
rect 11756 1087 11763 1333
rect 11776 887 11783 1213
rect 11796 1087 11803 1373
rect 11716 876 11743 883
rect 11736 863 11743 876
rect 11776 867 11783 873
rect 11676 856 11703 863
rect 11736 856 11763 863
rect 11676 827 11683 856
rect 11616 607 11623 613
rect 11636 587 11643 613
rect 11656 383 11663 713
rect 11696 627 11703 813
rect 11756 667 11763 856
rect 11736 616 11743 633
rect 11756 607 11763 653
rect 11656 376 11683 383
rect 11676 367 11683 376
rect 11396 336 11423 343
rect 11456 323 11463 343
rect 11716 343 11723 373
rect 11796 347 11803 1053
rect 11696 336 11723 343
rect 11436 316 11463 323
rect 11276 156 11283 173
rect 11336 167 11343 173
rect 11436 156 11443 316
rect 11476 156 11483 193
rect 11496 147 11503 193
rect 11636 176 11643 333
rect 11796 207 11803 333
rect 11816 247 11823 1573
rect 11876 1427 11883 2093
rect 11896 1407 11903 2113
rect 11936 2076 11943 2133
rect 11956 2107 11963 2293
rect 11976 2076 11983 2093
rect 11996 2087 12003 2776
rect 12016 2127 12023 3253
rect 12056 3227 12063 3253
rect 12096 3223 12103 3273
rect 12076 3216 12103 3223
rect 12036 2563 12043 3193
rect 12076 3067 12083 3216
rect 12056 3036 12083 3043
rect 12116 3036 12143 3043
rect 12056 2807 12063 3036
rect 12136 3007 12143 3036
rect 12036 2556 12063 2563
rect 12036 2307 12043 2556
rect 12056 2276 12063 2393
rect 12076 2307 12083 2793
rect 12036 2227 12043 2263
rect 11916 1367 11923 2073
rect 11956 2047 11963 2063
rect 11936 1627 11943 1833
rect 12016 1796 12023 2093
rect 12056 1796 12063 2013
rect 12096 1783 12103 2053
rect 11936 1596 11943 1613
rect 11976 1596 11983 1613
rect 11996 1607 12003 1783
rect 12036 1747 12043 1783
rect 12076 1776 12103 1783
rect 12076 1707 12083 1776
rect 12116 1727 12123 2743
rect 12216 2047 12223 11673
rect 11996 1576 12023 1583
rect 11836 387 11843 1233
rect 11876 1227 11883 1343
rect 11896 1287 11903 1323
rect 11876 1096 11883 1173
rect 11856 727 11863 1073
rect 11936 907 11943 1213
rect 11956 1087 11963 1353
rect 11976 1227 11983 1413
rect 12016 1287 12023 1576
rect 12036 1567 12043 1613
rect 11976 1127 11983 1133
rect 11936 887 11943 893
rect 11896 827 11903 843
rect 11916 727 11923 863
rect 11956 843 11963 1073
rect 11936 836 11963 843
rect 11856 636 11863 693
rect 11956 607 11963 836
rect 11976 647 11983 1113
rect 11996 1107 12003 1233
rect 12036 1143 12043 1393
rect 12056 1316 12063 1373
rect 12116 1287 12123 1303
rect 12076 1247 12083 1283
rect 12036 1136 12063 1143
rect 12056 1116 12063 1136
rect 12076 1096 12103 1103
rect 12096 1063 12103 1096
rect 12076 1056 12103 1063
rect 12036 823 12043 873
rect 12036 816 12063 823
rect 12076 767 12083 1056
rect 12056 616 12063 753
rect 12096 603 12103 813
rect 12076 596 12103 603
rect 11876 376 11883 593
rect 11856 347 11863 363
rect 11956 347 11963 593
rect 12016 376 12023 393
rect 12076 347 12083 363
rect 11836 176 11843 233
rect 11816 156 11823 173
rect 12036 167 12043 333
rect 11996 156 12023 163
rect 11256 127 11263 143
rect 7836 96 7883 103
rect 12016 -17 12023 156
rect 6696 -24 6723 -17
rect 6856 -24 6883 -17
rect 11996 -24 12023 -17
<< m3contact >>
rect 493 12013 507 12027
rect 1213 12013 1227 12027
rect 193 11913 207 11927
rect 153 11873 167 11887
rect 293 11893 307 11907
rect 253 11873 267 11887
rect 93 11853 107 11867
rect 133 11853 147 11867
rect 253 11833 267 11847
rect 173 11813 187 11827
rect 353 11853 367 11867
rect 333 11833 347 11847
rect 353 11813 367 11827
rect 133 11673 147 11687
rect 213 11673 227 11687
rect 313 11673 327 11687
rect 153 11653 167 11667
rect 93 11373 107 11387
rect 213 11413 227 11427
rect 373 11653 387 11667
rect 733 11913 747 11927
rect 873 11913 887 11927
rect 513 11893 527 11907
rect 553 11893 567 11907
rect 533 11873 547 11887
rect 693 11873 707 11887
rect 793 11893 807 11907
rect 753 11833 767 11847
rect 793 11833 807 11847
rect 773 11813 787 11827
rect 713 11713 727 11727
rect 633 11693 647 11707
rect 673 11673 687 11687
rect 793 11673 807 11687
rect 633 11413 647 11427
rect 753 11413 767 11427
rect 393 11393 407 11407
rect 433 11393 447 11407
rect 373 11373 387 11387
rect 833 11393 847 11407
rect 813 11373 827 11387
rect 353 11353 367 11367
rect 413 11353 427 11367
rect 573 11353 587 11367
rect 593 11353 607 11367
rect 773 11353 787 11367
rect 153 11213 167 11227
rect 373 11213 387 11227
rect 133 11193 147 11207
rect 233 11193 247 11207
rect 353 11193 367 11207
rect 213 11173 227 11187
rect 193 11073 207 11087
rect 373 10973 387 10987
rect 333 10933 347 10947
rect 753 11193 767 11207
rect 573 11173 587 11187
rect 733 11173 747 11187
rect 553 11153 567 11167
rect 413 10933 427 10947
rect 553 10933 567 10947
rect 353 10913 367 10927
rect 233 10893 247 10907
rect 373 10893 387 10907
rect 173 10873 187 10887
rect 53 10473 67 10487
rect 513 10913 527 10927
rect 773 11073 787 11087
rect 733 10933 747 10947
rect 593 10913 607 10927
rect 693 10913 707 10927
rect 413 10873 427 10887
rect 373 10713 387 10727
rect 113 10533 127 10547
rect 173 10533 187 10547
rect 113 10453 127 10467
rect 133 10433 147 10447
rect 273 10453 287 10467
rect 313 10433 327 10447
rect 353 10433 367 10447
rect 393 10433 407 10447
rect 173 10393 187 10407
rect 373 10393 387 10407
rect 193 10333 207 10347
rect 333 10333 347 10347
rect 373 10213 387 10227
rect 393 10213 407 10227
rect 73 9953 87 9967
rect 753 10893 767 10907
rect 573 10873 587 10887
rect 713 10873 727 10887
rect 533 10853 547 10867
rect 573 10853 587 10867
rect 493 10713 507 10727
rect 613 10713 627 10727
rect 693 10713 707 10727
rect 433 10513 447 10527
rect 433 10473 447 10487
rect 453 10453 467 10467
rect 473 10433 487 10447
rect 433 10393 447 10407
rect 413 10193 427 10207
rect 713 10693 727 10707
rect 813 10913 827 10927
rect 773 10493 787 10507
rect 1053 11893 1067 11907
rect 1073 11873 1087 11887
rect 893 11853 907 11867
rect 953 11853 967 11867
rect 933 11813 947 11827
rect 913 11693 927 11707
rect 1153 11873 1167 11887
rect 1113 11813 1127 11827
rect 1093 11673 1107 11687
rect 1133 11673 1147 11687
rect 893 11653 907 11667
rect 933 11653 947 11667
rect 973 11653 987 11667
rect 1073 11653 1087 11667
rect 1113 11653 1127 11667
rect 993 11433 1007 11447
rect 933 11393 947 11407
rect 913 11373 927 11387
rect 953 11373 967 11387
rect 993 11373 1007 11387
rect 973 11353 987 11367
rect 873 10733 887 10747
rect 853 10693 867 10707
rect 833 10473 847 10487
rect 873 10473 887 10487
rect 793 10453 807 10467
rect 833 10433 847 10447
rect 853 10433 867 10447
rect 433 9993 447 10007
rect 493 10213 507 10227
rect 573 10033 587 10047
rect 53 9933 67 9947
rect 373 9933 387 9947
rect 153 9773 167 9787
rect 73 9753 87 9767
rect 73 9633 87 9647
rect 13 6413 27 6427
rect 53 5853 67 5867
rect 33 5113 47 5127
rect 333 9773 347 9787
rect 353 9773 367 9787
rect 193 9753 207 9767
rect 213 9593 227 9607
rect 113 9453 127 9467
rect 173 9453 187 9467
rect 153 9293 167 9307
rect 153 9253 167 9267
rect 393 9753 407 9767
rect 473 9913 487 9927
rect 793 10313 807 10327
rect 673 10233 687 10247
rect 833 10233 847 10247
rect 633 10213 647 10227
rect 773 10213 787 10227
rect 613 10053 627 10067
rect 653 10053 667 10067
rect 613 9993 627 10007
rect 593 9973 607 9987
rect 633 9913 647 9927
rect 633 9833 647 9847
rect 573 9773 587 9787
rect 593 9753 607 9767
rect 513 9593 527 9607
rect 433 9573 447 9587
rect 733 9953 747 9967
rect 693 9813 707 9827
rect 693 9753 707 9767
rect 733 9753 747 9767
rect 793 9933 807 9947
rect 613 9733 627 9747
rect 653 9733 667 9747
rect 753 9733 767 9747
rect 813 9733 827 9747
rect 793 9713 807 9727
rect 553 9473 567 9487
rect 593 9473 607 9487
rect 793 9473 807 9487
rect 653 9373 667 9387
rect 713 9313 727 9327
rect 393 9293 407 9307
rect 553 9293 567 9307
rect 373 9273 387 9287
rect 333 9253 347 9267
rect 313 9233 327 9247
rect 353 9233 367 9247
rect 393 9233 407 9247
rect 393 9053 407 9067
rect 173 9013 187 9027
rect 253 9013 267 9027
rect 113 8973 127 8987
rect 173 8993 187 9007
rect 233 8993 247 9007
rect 153 8973 167 8987
rect 193 8973 207 8987
rect 233 8913 247 8927
rect 153 8813 167 8827
rect 133 8733 147 8747
rect 333 8993 347 9007
rect 353 8933 367 8947
rect 273 8813 287 8827
rect 253 8753 267 8767
rect 113 8553 127 8567
rect 233 8553 247 8567
rect 153 8533 167 8547
rect 133 8513 147 8527
rect 153 8453 167 8467
rect 313 8773 327 8787
rect 293 8753 307 8767
rect 333 8753 347 8767
rect 313 8513 327 8527
rect 273 8493 287 8507
rect 333 8473 347 8487
rect 213 8453 227 8467
rect 173 8413 187 8427
rect 193 8313 207 8327
rect 153 8273 167 8287
rect 133 8073 147 8087
rect 173 8053 187 8067
rect 233 8413 247 8427
rect 313 8333 327 8347
rect 313 8313 327 8327
rect 353 8313 367 8327
rect 373 8273 387 8287
rect 253 8073 267 8087
rect 333 8073 347 8087
rect 233 8053 247 8067
rect 193 8033 207 8047
rect 213 8033 227 8047
rect 113 7833 127 7847
rect 153 7833 167 7847
rect 153 7813 167 7827
rect 133 7793 147 7807
rect 233 7793 247 7807
rect 173 7693 187 7707
rect 213 7693 227 7707
rect 153 7613 167 7627
rect 193 7553 207 7567
rect 133 7533 147 7547
rect 173 7513 187 7527
rect 173 7353 187 7367
rect 233 7513 247 7527
rect 113 7313 127 7327
rect 213 7333 227 7347
rect 413 8353 427 8367
rect 393 8053 407 8067
rect 333 8033 347 8047
rect 353 7993 367 8007
rect 393 7993 407 8007
rect 413 7993 427 8007
rect 393 7873 407 7887
rect 353 7813 367 7827
rect 413 7813 427 7827
rect 513 9273 527 9287
rect 813 9453 827 9467
rect 873 9353 887 9367
rect 933 11233 947 11247
rect 953 11153 967 11167
rect 1013 11133 1027 11147
rect 953 10973 967 10987
rect 993 10913 1007 10927
rect 913 10893 927 10907
rect 933 10893 947 10907
rect 1153 11393 1167 11407
rect 1193 11373 1207 11387
rect 1113 11353 1127 11367
rect 1113 11193 1127 11207
rect 1153 11173 1167 11187
rect 1093 11153 1107 11167
rect 1133 11153 1147 11167
rect 1073 10993 1087 11007
rect 1033 10933 1047 10947
rect 1173 11133 1187 11147
rect 1133 11053 1147 11067
rect 5993 12013 6007 12027
rect 6213 12013 6227 12027
rect 1513 11933 1527 11947
rect 1673 11933 1687 11947
rect 5793 11933 5807 11947
rect 1253 11873 1267 11887
rect 1393 11873 1407 11887
rect 1233 11833 1247 11847
rect 1273 11833 1287 11847
rect 1253 11773 1267 11787
rect 1233 11193 1247 11207
rect 1173 11013 1187 11027
rect 1213 11013 1227 11027
rect 1153 10953 1167 10967
rect 1013 10893 1027 10907
rect 1033 10793 1047 10807
rect 973 10693 987 10707
rect 1013 10453 1027 10467
rect 973 10433 987 10447
rect 993 10433 1007 10447
rect 1033 10433 1047 10447
rect 933 10213 947 10227
rect 993 10213 1007 10227
rect 913 9953 927 9967
rect 973 10193 987 10207
rect 1013 10193 1027 10207
rect 993 9953 1007 9967
rect 1113 10913 1127 10927
rect 1153 10913 1167 10927
rect 1213 10993 1227 11007
rect 1173 10473 1187 10487
rect 1173 10453 1187 10467
rect 1093 10433 1107 10447
rect 1073 10253 1087 10267
rect 1053 10213 1067 10227
rect 1013 9933 1027 9947
rect 1033 9933 1047 9947
rect 1133 10293 1147 10307
rect 1193 10273 1207 10287
rect 1173 10253 1187 10267
rect 1133 10233 1147 10247
rect 1193 10213 1207 10227
rect 1153 10193 1167 10207
rect 1133 9933 1147 9947
rect 1093 9913 1107 9927
rect 973 9873 987 9887
rect 1113 9873 1127 9887
rect 993 9793 1007 9807
rect 913 9773 927 9787
rect 993 9773 1007 9787
rect 953 9753 967 9767
rect 1153 9813 1167 9827
rect 1333 11693 1347 11707
rect 1273 11673 1287 11687
rect 1273 11633 1287 11647
rect 1313 11633 1327 11647
rect 1353 11633 1367 11647
rect 1313 11373 1327 11387
rect 1333 11373 1347 11387
rect 1353 11333 1367 11347
rect 1313 11213 1327 11227
rect 1353 11213 1367 11227
rect 1293 11193 1307 11207
rect 1333 11193 1347 11207
rect 1253 11173 1267 11187
rect 1273 11173 1287 11187
rect 1313 11173 1327 11187
rect 1273 11133 1287 11147
rect 1313 10933 1327 10947
rect 1293 10913 1307 10927
rect 1233 10753 1247 10767
rect 1313 10733 1327 10747
rect 1293 10693 1307 10707
rect 1373 10333 1387 10347
rect 1333 10293 1347 10307
rect 1353 10213 1367 10227
rect 1293 9993 1307 10007
rect 1273 9953 1287 9967
rect 1413 11853 1427 11867
rect 1473 11813 1487 11827
rect 1613 11853 1627 11867
rect 2253 11913 2267 11927
rect 2613 11913 2627 11927
rect 2933 11913 2947 11927
rect 3813 11913 3827 11927
rect 4753 11913 4767 11927
rect 5133 11913 5147 11927
rect 5773 11913 5787 11927
rect 2033 11893 2047 11907
rect 1813 11873 1827 11887
rect 1593 11713 1607 11727
rect 1493 11653 1507 11667
rect 1533 11653 1547 11667
rect 1473 11433 1487 11447
rect 1453 11413 1467 11427
rect 1513 11413 1527 11427
rect 1593 11653 1607 11667
rect 1573 11353 1587 11367
rect 1633 11833 1647 11847
rect 1693 11713 1707 11727
rect 1673 11633 1687 11647
rect 1713 11633 1727 11647
rect 1653 11373 1667 11387
rect 1533 11333 1547 11347
rect 1593 11333 1607 11347
rect 1613 11333 1627 11347
rect 1553 11313 1567 11327
rect 1513 11273 1527 11287
rect 1473 11193 1487 11207
rect 1533 11213 1547 11227
rect 1473 11073 1487 11087
rect 1473 11013 1487 11027
rect 1573 10973 1587 10987
rect 1553 10933 1567 10947
rect 1493 10873 1507 10887
rect 1513 10753 1527 10767
rect 1433 10733 1447 10747
rect 1473 10713 1487 10727
rect 1453 10693 1467 10707
rect 1493 10693 1507 10707
rect 1493 10433 1507 10447
rect 1533 10513 1547 10527
rect 1513 10313 1527 10327
rect 1533 10313 1547 10327
rect 1433 10193 1447 10207
rect 1553 10193 1567 10207
rect 1213 9873 1227 9887
rect 1173 9753 1187 9767
rect 1233 9753 1247 9767
rect 1013 9733 1027 9747
rect 973 9713 987 9727
rect 973 9573 987 9587
rect 993 9453 1007 9467
rect 953 9433 967 9447
rect 893 9333 907 9347
rect 733 9293 747 9307
rect 773 9293 787 9307
rect 833 9293 847 9307
rect 913 9293 927 9307
rect 493 9253 507 9267
rect 533 9233 547 9247
rect 593 9233 607 9247
rect 533 9033 547 9047
rect 473 8973 487 8987
rect 493 8953 507 8967
rect 533 8953 547 8967
rect 553 8813 567 8827
rect 493 8773 507 8787
rect 513 8773 527 8787
rect 573 8773 587 8787
rect 513 8513 527 8527
rect 493 8493 507 8507
rect 533 8493 547 8507
rect 873 9273 887 9287
rect 733 9253 747 9267
rect 693 9033 707 9047
rect 933 9253 947 9267
rect 653 9013 667 9027
rect 833 9013 847 9027
rect 893 9013 907 9027
rect 673 8953 687 8967
rect 653 8933 667 8947
rect 693 8913 707 8927
rect 793 8833 807 8847
rect 753 8813 767 8827
rect 773 8813 787 8827
rect 613 8793 627 8807
rect 633 8793 647 8807
rect 593 8493 607 8507
rect 573 8473 587 8487
rect 473 8453 487 8467
rect 673 8533 687 8547
rect 653 8513 667 8527
rect 693 8513 707 8527
rect 633 8353 647 8367
rect 573 8313 587 8327
rect 473 7853 487 7867
rect 453 7833 467 7847
rect 473 7813 487 7827
rect 473 7793 487 7807
rect 413 7613 427 7627
rect 373 7553 387 7567
rect 333 7533 347 7547
rect 393 7533 407 7547
rect 393 7513 407 7527
rect 353 7453 367 7467
rect 313 7353 327 7367
rect 353 7353 367 7367
rect 273 7333 287 7347
rect 333 7333 347 7347
rect 373 7333 387 7347
rect 253 7293 267 7307
rect 153 7093 167 7107
rect 133 7073 147 7087
rect 193 7073 207 7087
rect 173 7053 187 7067
rect 153 7033 167 7047
rect 93 6913 107 6927
rect 173 6893 187 6907
rect 133 6853 147 6867
rect 333 7293 347 7307
rect 293 7073 307 7087
rect 333 7073 347 7087
rect 273 7053 287 7067
rect 153 6833 167 6847
rect 193 6833 207 6847
rect 153 6613 167 6627
rect 173 6573 187 6587
rect 133 6433 147 6447
rect 173 6413 187 6427
rect 133 6393 147 6407
rect 353 7033 367 7047
rect 333 6873 347 6887
rect 333 6853 347 6867
rect 353 6833 367 6847
rect 393 6633 407 6647
rect 393 6613 407 6627
rect 453 7573 467 7587
rect 433 6613 447 6627
rect 353 6593 367 6607
rect 333 6573 347 6587
rect 413 6553 427 6567
rect 373 6493 387 6507
rect 313 6413 327 6427
rect 313 6393 327 6407
rect 353 6393 367 6407
rect 333 6353 347 6367
rect 313 5933 327 5947
rect 293 5913 307 5927
rect 333 5913 347 5927
rect 373 5913 387 5927
rect 153 5893 167 5907
rect 313 5893 327 5907
rect 353 5893 367 5907
rect 133 5873 147 5887
rect 173 5853 187 5867
rect 593 8293 607 8307
rect 693 8493 707 8507
rect 653 8253 667 8267
rect 733 8413 747 8427
rect 813 8793 827 8807
rect 893 8993 907 9007
rect 933 8993 947 9007
rect 873 8953 887 8967
rect 993 8973 1007 8987
rect 933 8913 947 8927
rect 913 8873 927 8887
rect 853 8833 867 8847
rect 873 8793 887 8807
rect 973 8793 987 8807
rect 913 8773 927 8787
rect 953 8773 967 8787
rect 873 8753 887 8767
rect 853 8493 867 8507
rect 893 8493 907 8507
rect 833 8473 847 8487
rect 873 8473 887 8487
rect 773 8433 787 8447
rect 753 8293 767 8307
rect 793 8413 807 8427
rect 1273 9713 1287 9727
rect 1353 9953 1367 9967
rect 1393 9953 1407 9967
rect 1413 9953 1427 9967
rect 1333 9913 1347 9927
rect 1293 9693 1307 9707
rect 1373 9853 1387 9867
rect 1493 9953 1507 9967
rect 1533 9953 1547 9967
rect 1473 9933 1487 9947
rect 1513 9893 1527 9907
rect 1433 9813 1447 9827
rect 1413 9753 1427 9767
rect 1393 9733 1407 9747
rect 1413 9713 1427 9727
rect 1373 9693 1387 9707
rect 1053 9593 1067 9607
rect 1333 9593 1347 9607
rect 1193 9573 1207 9587
rect 1033 9333 1047 9347
rect 1093 9433 1107 9447
rect 1113 9373 1127 9387
rect 1133 9353 1147 9367
rect 1093 9233 1107 9247
rect 1073 9053 1087 9067
rect 1073 9033 1087 9047
rect 1093 8973 1107 8987
rect 1053 8953 1067 8967
rect 1053 8813 1067 8827
rect 1033 8613 1047 8627
rect 1073 8793 1087 8807
rect 1113 8773 1127 8787
rect 1053 8533 1067 8547
rect 1093 8533 1107 8547
rect 1033 8513 1047 8527
rect 1073 8513 1087 8527
rect 1013 8333 1027 8347
rect 773 8273 787 8287
rect 813 8273 827 8287
rect 993 8293 1007 8307
rect 973 8273 987 8287
rect 873 8233 887 8247
rect 1013 8233 1027 8247
rect 693 8133 707 8147
rect 853 8133 867 8147
rect 693 8053 707 8067
rect 553 7993 567 8007
rect 573 7873 587 7887
rect 613 7873 627 7887
rect 673 7853 687 7867
rect 613 7833 627 7847
rect 633 7833 647 7847
rect 593 7813 607 7827
rect 533 7793 547 7807
rect 573 7793 587 7807
rect 653 7793 667 7807
rect 773 7973 787 7987
rect 733 7913 747 7927
rect 833 7893 847 7907
rect 773 7853 787 7867
rect 493 7573 507 7587
rect 593 7573 607 7587
rect 493 7553 507 7567
rect 533 7553 547 7567
rect 713 7633 727 7647
rect 793 7633 807 7647
rect 693 7573 707 7587
rect 733 7573 747 7587
rect 713 7553 727 7567
rect 673 7513 687 7527
rect 653 7393 667 7407
rect 573 7373 587 7387
rect 533 7353 547 7367
rect 713 7393 727 7407
rect 613 7353 627 7367
rect 673 7353 687 7367
rect 553 7313 567 7327
rect 633 7333 647 7347
rect 653 7313 667 7327
rect 593 7113 607 7127
rect 493 7053 507 7067
rect 533 7033 547 7047
rect 533 7013 547 7027
rect 473 6873 487 6887
rect 693 7333 707 7347
rect 693 7073 707 7087
rect 673 6973 687 6987
rect 693 6913 707 6927
rect 553 6893 567 6907
rect 653 6893 667 6907
rect 573 6853 587 6867
rect 533 6813 547 6827
rect 513 6653 527 6667
rect 493 6573 507 6587
rect 513 6573 527 6587
rect 553 6573 567 6587
rect 593 6573 607 6587
rect 533 6533 547 6547
rect 573 6533 587 6547
rect 493 6433 507 6447
rect 573 6513 587 6527
rect 533 6353 547 6367
rect 453 6153 467 6167
rect 453 6133 467 6147
rect 513 6133 527 6147
rect 553 6113 567 6127
rect 533 5953 547 5967
rect 433 5913 447 5927
rect 433 5873 447 5887
rect 513 5893 527 5907
rect 473 5853 487 5867
rect 313 5773 327 5787
rect 413 5773 427 5787
rect 133 5653 147 5667
rect 113 5633 127 5647
rect 973 8033 987 8047
rect 1033 8033 1047 8047
rect 953 7993 967 8007
rect 873 7853 887 7867
rect 873 7813 887 7827
rect 1113 8333 1127 8347
rect 1093 8033 1107 8047
rect 1053 8013 1067 8027
rect 1093 7993 1107 8007
rect 1053 7913 1067 7927
rect 933 7713 947 7727
rect 1033 7713 1047 7727
rect 893 7553 907 7567
rect 1093 7813 1107 7827
rect 973 7653 987 7667
rect 953 7513 967 7527
rect 873 7493 887 7507
rect 913 7493 927 7507
rect 853 7433 867 7447
rect 813 7373 827 7387
rect 793 7313 807 7327
rect 873 7213 887 7227
rect 753 7093 767 7107
rect 733 7053 747 7067
rect 733 6973 747 6987
rect 793 6853 807 6867
rect 713 6833 727 6847
rect 693 6633 707 6647
rect 753 6573 767 6587
rect 713 6553 727 6567
rect 733 6553 747 6567
rect 693 6533 707 6547
rect 713 6373 727 6387
rect 733 6353 747 6367
rect 833 6253 847 6267
rect 653 6153 667 6167
rect 653 5913 667 5927
rect 573 5893 587 5907
rect 653 5853 667 5867
rect 333 5733 347 5747
rect 473 5733 487 5747
rect 533 5733 547 5747
rect 273 5633 287 5647
rect 313 5633 327 5647
rect 373 5633 387 5647
rect 393 5613 407 5627
rect 253 5193 267 5207
rect 313 5193 327 5207
rect 293 5173 307 5187
rect 133 5153 147 5167
rect 253 5153 267 5167
rect 333 5153 347 5167
rect 273 5133 287 5147
rect 313 5133 327 5147
rect 113 5113 127 5127
rect 173 5053 187 5067
rect 133 4953 147 4967
rect 113 4933 127 4947
rect 313 4933 327 4947
rect 293 4913 307 4927
rect 173 4893 187 4907
rect 73 4633 87 4647
rect 193 4653 207 4667
rect 333 4893 347 4907
rect 353 4653 367 4667
rect 173 4633 187 4647
rect 153 4613 167 4627
rect 33 4433 47 4447
rect 53 4433 67 4447
rect 193 4613 207 4627
rect 333 4413 347 4427
rect 333 4353 347 4367
rect 93 4293 107 4307
rect 173 4293 187 4307
rect 293 4293 307 4307
rect 53 3953 67 3967
rect 33 3253 47 3267
rect 13 2973 27 2987
rect 73 2913 87 2927
rect 133 4173 147 4187
rect 193 4113 207 4127
rect 633 5653 647 5667
rect 493 5573 507 5587
rect 613 5433 627 5447
rect 693 5953 707 5967
rect 713 5913 727 5927
rect 673 5613 687 5627
rect 513 5173 527 5187
rect 573 5173 587 5187
rect 593 5173 607 5187
rect 493 5153 507 5167
rect 453 5133 467 5147
rect 433 5053 447 5067
rect 373 4413 387 4427
rect 373 4353 387 4367
rect 393 4293 407 4307
rect 353 4273 367 4287
rect 393 4273 407 4287
rect 373 4193 387 4207
rect 353 4153 367 4167
rect 393 4153 407 4167
rect 313 4113 327 4127
rect 293 4073 307 4087
rect 173 3893 187 3907
rect 373 4073 387 4087
rect 373 3993 387 4007
rect 353 3833 367 3847
rect 393 3833 407 3847
rect 353 3713 367 3727
rect 133 3693 147 3707
rect 133 3153 147 3167
rect 113 3053 127 3067
rect 313 3693 327 3707
rect 413 3713 427 3727
rect 413 3653 427 3667
rect 193 3613 207 3627
rect 333 3613 347 3627
rect 473 5113 487 5127
rect 513 4953 527 4967
rect 553 4953 567 4967
rect 453 4913 467 4927
rect 473 4913 487 4927
rect 453 4853 467 4867
rect 453 4453 467 4467
rect 453 4173 467 4187
rect 533 4913 547 4927
rect 513 4673 527 4687
rect 533 4633 547 4647
rect 493 4493 507 4507
rect 573 4553 587 4567
rect 593 4513 607 4527
rect 573 4473 587 4487
rect 533 4453 547 4467
rect 573 4433 587 4447
rect 533 4233 547 4247
rect 513 4193 527 4207
rect 473 3993 487 4007
rect 453 3973 467 3987
rect 373 3493 387 3507
rect 393 3493 407 3507
rect 393 3233 407 3247
rect 193 3153 207 3167
rect 193 3133 207 3147
rect 173 3073 187 3087
rect 333 3113 347 3127
rect 253 3093 267 3107
rect 113 3013 127 3027
rect 153 3013 167 3027
rect 193 3013 207 3027
rect 33 2833 47 2847
rect 93 2833 107 2847
rect 133 2733 147 2747
rect 173 2553 187 2567
rect 133 2533 147 2547
rect 33 2333 47 2347
rect 13 2233 27 2247
rect 313 3073 327 3087
rect 273 2913 287 2927
rect 353 3053 367 3067
rect 333 3033 347 3047
rect 373 3033 387 3047
rect 393 2873 407 2887
rect 293 2573 307 2587
rect 433 3513 447 3527
rect 493 3973 507 3987
rect 513 3953 527 3967
rect 513 3793 527 3807
rect 653 5213 667 5227
rect 693 5433 707 5447
rect 733 5873 747 5887
rect 633 5153 647 5167
rect 633 5113 647 5127
rect 633 4473 647 4487
rect 713 5173 727 5187
rect 713 5133 727 5147
rect 693 5113 707 5127
rect 673 5093 687 5107
rect 673 5033 687 5047
rect 713 4973 727 4987
rect 673 4953 687 4967
rect 693 4893 707 4907
rect 713 4693 727 4707
rect 693 4653 707 4667
rect 653 4293 667 4307
rect 713 4293 727 4307
rect 613 4233 627 4247
rect 553 4173 567 4187
rect 613 4173 627 4187
rect 853 5893 867 5907
rect 853 5653 867 5667
rect 853 5633 867 5647
rect 833 5613 847 5627
rect 773 5593 787 5607
rect 813 5453 827 5467
rect 833 5453 847 5467
rect 773 5433 787 5447
rect 773 5393 787 5407
rect 753 5293 767 5307
rect 813 5413 827 5427
rect 933 7093 947 7107
rect 953 7033 967 7047
rect 933 6953 947 6967
rect 893 6853 907 6867
rect 933 6853 947 6867
rect 993 7633 1007 7647
rect 993 7493 1007 7507
rect 1153 9293 1167 9307
rect 1173 9273 1187 9287
rect 1153 9253 1167 9267
rect 1393 9473 1407 9487
rect 1433 9473 1447 9487
rect 1373 9453 1387 9467
rect 1313 9373 1327 9387
rect 1213 9273 1227 9287
rect 1253 9253 1267 9267
rect 1293 9253 1307 9267
rect 1193 9233 1207 9247
rect 1233 9233 1247 9247
rect 1273 9073 1287 9087
rect 1173 8953 1187 8967
rect 1253 8953 1267 8967
rect 1273 8953 1287 8967
rect 1233 8833 1247 8847
rect 1173 8813 1187 8827
rect 1213 8793 1227 8807
rect 1153 8773 1167 8787
rect 1193 8773 1207 8787
rect 1233 8773 1247 8787
rect 1233 8553 1247 8567
rect 1173 8533 1187 8547
rect 1193 8513 1207 8527
rect 1433 9433 1447 9447
rect 1513 9873 1527 9887
rect 1473 9473 1487 9487
rect 1453 9333 1467 9347
rect 1433 9313 1447 9327
rect 1493 9293 1507 9307
rect 1453 9273 1467 9287
rect 1473 9253 1487 9267
rect 1653 11173 1667 11187
rect 1693 11333 1707 11347
rect 1693 11213 1707 11227
rect 1693 11193 1707 11207
rect 1753 11193 1767 11207
rect 1773 11193 1787 11207
rect 1613 11093 1627 11107
rect 1713 11173 1727 11187
rect 1733 11153 1747 11167
rect 1773 11153 1787 11167
rect 1753 11033 1767 11047
rect 1653 11013 1667 11027
rect 1693 10993 1707 11007
rect 1833 11833 1847 11847
rect 1973 11813 1987 11827
rect 1953 11693 1967 11707
rect 1913 11673 1927 11687
rect 1853 11593 1867 11607
rect 1913 11573 1927 11587
rect 1873 11433 1887 11447
rect 1873 11413 1887 11427
rect 1833 11353 1847 11367
rect 1833 11313 1847 11327
rect 1893 11253 1907 11267
rect 1913 11173 1927 11187
rect 1933 11153 1947 11167
rect 1853 11133 1867 11147
rect 1833 11053 1847 11067
rect 1753 10973 1767 10987
rect 1793 10973 1807 10987
rect 1613 10873 1627 10887
rect 1653 10873 1667 10887
rect 1693 10853 1707 10867
rect 1633 10753 1647 10767
rect 1673 10673 1687 10687
rect 1633 10433 1647 10447
rect 1593 10293 1607 10307
rect 1613 10293 1627 10307
rect 1593 10253 1607 10267
rect 1593 10193 1607 10207
rect 1593 9953 1607 9967
rect 1713 10333 1727 10347
rect 1673 10253 1687 10267
rect 1653 10233 1667 10247
rect 1673 10233 1687 10247
rect 1733 10293 1747 10307
rect 2013 11853 2027 11867
rect 2053 11773 2067 11787
rect 2133 11713 2147 11727
rect 2013 11653 2027 11667
rect 2073 11633 2087 11647
rect 1993 11473 2007 11487
rect 1973 11413 1987 11427
rect 2113 11453 2127 11467
rect 2073 11433 2087 11447
rect 2033 11413 2047 11427
rect 2053 11393 2067 11407
rect 2093 11293 2107 11307
rect 2073 11173 2087 11187
rect 2213 11873 2227 11887
rect 2433 11893 2447 11907
rect 2553 11893 2567 11907
rect 2913 11893 2927 11907
rect 2973 11893 2987 11907
rect 2413 11873 2427 11887
rect 2193 11813 2207 11827
rect 2373 11813 2387 11827
rect 2333 11793 2347 11807
rect 2173 11693 2187 11707
rect 2153 11633 2167 11647
rect 2273 11673 2287 11687
rect 2273 11653 2287 11667
rect 2313 11653 2327 11667
rect 2173 11613 2187 11627
rect 2253 11613 2267 11627
rect 2193 11593 2207 11607
rect 2133 11373 2147 11387
rect 2113 11273 2127 11287
rect 2153 11233 2167 11247
rect 2113 11193 2127 11207
rect 2153 11173 2167 11187
rect 2133 11153 2147 11167
rect 2093 11113 2107 11127
rect 1993 11053 2007 11067
rect 2013 10973 2027 10987
rect 1833 10893 1847 10907
rect 1793 10873 1807 10887
rect 1813 10733 1827 10747
rect 1893 10733 1907 10747
rect 1873 10693 1887 10707
rect 1893 10693 1907 10707
rect 1813 10673 1827 10687
rect 1793 10413 1807 10427
rect 1633 9913 1647 9927
rect 1633 9833 1647 9847
rect 1633 9813 1647 9827
rect 1593 9773 1607 9787
rect 1573 9733 1587 9747
rect 1613 9713 1627 9727
rect 1553 9693 1567 9707
rect 1573 9593 1587 9607
rect 1533 9353 1547 9367
rect 1553 9293 1567 9307
rect 1533 9253 1547 9267
rect 1373 8973 1387 8987
rect 1413 8953 1427 8967
rect 1393 8913 1407 8927
rect 1433 8873 1447 8887
rect 1353 8813 1367 8827
rect 1433 8813 1447 8827
rect 1393 8793 1407 8807
rect 1333 8773 1347 8787
rect 1313 8633 1327 8647
rect 1353 8533 1367 8547
rect 1213 8453 1227 8467
rect 1293 8473 1307 8487
rect 1253 8433 1267 8447
rect 1213 8393 1227 8407
rect 1193 8333 1207 8347
rect 1233 8333 1247 8347
rect 1273 8333 1287 8347
rect 1173 8293 1187 8307
rect 1253 8273 1267 8287
rect 1213 8253 1227 8267
rect 1133 8153 1147 8167
rect 1173 8053 1187 8067
rect 1133 8033 1147 8047
rect 1193 8013 1207 8027
rect 1153 7953 1167 7967
rect 1133 7813 1147 7827
rect 1253 7853 1267 7867
rect 1413 8593 1427 8607
rect 1393 8273 1407 8287
rect 1353 8253 1367 8267
rect 1393 8073 1407 8087
rect 1333 8033 1347 8047
rect 1353 7993 1367 8007
rect 1353 7953 1367 7967
rect 1293 7873 1307 7887
rect 1353 7873 1367 7887
rect 1273 7813 1287 7827
rect 1313 7793 1327 7807
rect 1053 7493 1067 7507
rect 1093 7393 1107 7407
rect 1213 7653 1227 7667
rect 1293 7513 1307 7527
rect 1233 7453 1247 7467
rect 1193 7433 1207 7447
rect 1153 7353 1167 7367
rect 1093 7073 1107 7087
rect 1053 7033 1067 7047
rect 1053 6993 1067 7007
rect 1113 7053 1127 7067
rect 1133 7033 1147 7047
rect 1013 6873 1027 6887
rect 1133 6973 1147 6987
rect 1073 6853 1087 6867
rect 1153 6753 1167 6767
rect 1153 6633 1167 6647
rect 913 6573 927 6587
rect 933 6553 947 6567
rect 973 6573 987 6587
rect 1093 6553 1107 6567
rect 1113 6533 1127 6547
rect 953 6513 967 6527
rect 893 6493 907 6507
rect 1173 6413 1187 6427
rect 1053 6253 1067 6267
rect 893 6213 907 6227
rect 1033 6133 1047 6147
rect 1173 6133 1187 6147
rect 893 5893 907 5907
rect 893 5653 907 5667
rect 873 5613 887 5627
rect 793 5193 807 5207
rect 793 5153 807 5167
rect 813 5113 827 5127
rect 773 5073 787 5087
rect 873 5073 887 5087
rect 913 5633 927 5647
rect 973 6113 987 6127
rect 973 5973 987 5987
rect 1093 6093 1107 6107
rect 1133 6033 1147 6047
rect 1093 5973 1107 5987
rect 1033 5953 1047 5967
rect 993 5893 1007 5907
rect 1033 5673 1047 5687
rect 913 5453 927 5467
rect 973 5413 987 5427
rect 1073 5633 1087 5647
rect 1053 5613 1067 5627
rect 1113 5613 1127 5627
rect 1093 5553 1107 5567
rect 993 5373 1007 5387
rect 1033 5293 1047 5307
rect 1093 5413 1107 5427
rect 913 5153 927 5167
rect 933 5053 947 5067
rect 913 4993 927 5007
rect 893 4973 907 4987
rect 893 4933 907 4947
rect 1093 5153 1107 5167
rect 1133 5593 1147 5607
rect 1133 5493 1147 5507
rect 1253 7353 1267 7367
rect 1333 7493 1347 7507
rect 1513 8973 1527 8987
rect 1493 8573 1507 8587
rect 1693 10213 1707 10227
rect 1733 10213 1747 10227
rect 1793 10073 1807 10087
rect 1673 9953 1687 9967
rect 1713 9953 1727 9967
rect 1753 9953 1767 9967
rect 1833 10473 1847 10487
rect 1813 9933 1827 9947
rect 1693 9913 1707 9927
rect 1673 9893 1687 9907
rect 1733 9733 1747 9747
rect 1653 9573 1667 9587
rect 1653 9533 1667 9547
rect 1613 9473 1627 9487
rect 1593 9453 1607 9467
rect 1633 9433 1647 9447
rect 1573 9113 1587 9127
rect 1553 9093 1567 9107
rect 1633 9253 1647 9267
rect 1593 9013 1607 9027
rect 1553 8973 1567 8987
rect 1573 8933 1587 8947
rect 1553 8913 1567 8927
rect 1533 8833 1547 8847
rect 1593 8793 1607 8807
rect 1553 8773 1567 8787
rect 1433 8493 1447 8507
rect 1493 8513 1507 8527
rect 1473 8493 1487 8507
rect 1573 8573 1587 8587
rect 1553 8513 1567 8527
rect 1453 8473 1467 8487
rect 1453 8433 1467 8447
rect 1633 8633 1647 8647
rect 1713 9473 1727 9487
rect 1673 9433 1687 9447
rect 1693 9333 1707 9347
rect 1673 8993 1687 9007
rect 1713 9293 1727 9307
rect 1733 9173 1747 9187
rect 1793 9853 1807 9867
rect 1773 9713 1787 9727
rect 1853 10413 1867 10427
rect 1853 10213 1867 10227
rect 1853 9973 1867 9987
rect 1853 9893 1867 9907
rect 1853 9793 1867 9807
rect 1833 9533 1847 9547
rect 1913 10673 1927 10687
rect 1913 10413 1927 10427
rect 1993 10913 2007 10927
rect 1953 10873 1967 10887
rect 1953 10733 1967 10747
rect 1993 10733 2007 10747
rect 2073 10733 2087 10747
rect 2053 10693 2067 10707
rect 1973 10513 1987 10527
rect 1953 10313 1967 10327
rect 1933 10293 1947 10307
rect 1953 10233 1967 10247
rect 2013 10493 2027 10507
rect 1993 10193 2007 10207
rect 1933 10053 1947 10067
rect 1893 9913 1907 9927
rect 1953 9933 1967 9947
rect 1933 9913 1947 9927
rect 1913 9893 1927 9907
rect 1933 9833 1947 9847
rect 1873 9673 1887 9687
rect 1953 9793 1967 9807
rect 1993 9633 2007 9647
rect 1973 9573 1987 9587
rect 1893 9553 1907 9567
rect 1893 9493 1907 9507
rect 1873 9453 1887 9467
rect 1853 9433 1867 9447
rect 1913 9433 1927 9447
rect 1833 9273 1847 9287
rect 1793 9253 1807 9267
rect 1873 9213 1887 9227
rect 1753 9153 1767 9167
rect 1993 9493 2007 9507
rect 1993 9433 2007 9447
rect 2053 10453 2067 10467
rect 2133 11053 2147 11067
rect 2293 11533 2307 11547
rect 2253 11373 2267 11387
rect 2313 11373 2327 11387
rect 2213 11313 2227 11327
rect 2233 11313 2247 11327
rect 2273 11313 2287 11327
rect 2233 11273 2247 11287
rect 2193 10933 2207 10947
rect 2193 10913 2207 10927
rect 2253 11193 2267 11207
rect 2253 11113 2267 11127
rect 2553 11753 2567 11767
rect 2453 11673 2467 11687
rect 2393 11593 2407 11607
rect 2393 11453 2407 11467
rect 2753 11833 2767 11847
rect 2613 11753 2627 11767
rect 2873 11753 2887 11767
rect 2793 11733 2807 11747
rect 2693 11693 2707 11707
rect 2773 11693 2787 11707
rect 2833 11693 2847 11707
rect 2653 11673 2667 11687
rect 2713 11673 2727 11687
rect 2633 11653 2647 11667
rect 2593 11633 2607 11647
rect 2693 11633 2707 11647
rect 2673 11613 2687 11627
rect 2653 11593 2667 11607
rect 2493 11493 2507 11507
rect 2433 11433 2447 11447
rect 2433 11413 2447 11427
rect 2413 11393 2427 11407
rect 2413 11373 2427 11387
rect 2393 11353 2407 11367
rect 2373 11253 2387 11267
rect 2393 11253 2407 11267
rect 2333 11213 2347 11227
rect 2293 11193 2307 11207
rect 2313 11153 2327 11167
rect 2353 11153 2367 11167
rect 2433 11173 2447 11187
rect 2313 11113 2327 11127
rect 2413 11113 2427 11127
rect 2313 11093 2327 11107
rect 2133 10453 2147 10467
rect 2073 10413 2087 10427
rect 2113 10353 2127 10367
rect 2273 10753 2287 10767
rect 2233 10713 2247 10727
rect 2473 11413 2487 11427
rect 2513 11453 2527 11467
rect 2573 11433 2587 11447
rect 2633 11433 2647 11447
rect 2573 11393 2587 11407
rect 2613 11393 2627 11407
rect 2553 11373 2567 11387
rect 2593 11373 2607 11387
rect 2513 11233 2527 11247
rect 2553 11233 2567 11247
rect 2453 10993 2467 11007
rect 2513 11193 2527 11207
rect 2573 11213 2587 11227
rect 2493 11173 2507 11187
rect 2533 11173 2547 11187
rect 2573 11173 2587 11187
rect 2693 11393 2707 11407
rect 2673 11353 2687 11367
rect 2653 11313 2667 11327
rect 2673 11293 2687 11307
rect 2673 11273 2687 11287
rect 2853 11653 2867 11667
rect 2753 11473 2767 11487
rect 2733 11373 2747 11387
rect 2833 11413 2847 11427
rect 2793 11393 2807 11407
rect 2793 11333 2807 11347
rect 2713 11293 2727 11307
rect 2793 11233 2807 11247
rect 2713 11133 2727 11147
rect 2633 10973 2647 10987
rect 2353 10933 2367 10947
rect 2473 10933 2487 10947
rect 2373 10873 2387 10887
rect 2553 10913 2567 10927
rect 2453 10873 2467 10887
rect 2473 10873 2487 10887
rect 2533 10873 2547 10887
rect 2593 10873 2607 10887
rect 2393 10833 2407 10847
rect 2593 10793 2607 10807
rect 2493 10773 2507 10787
rect 2213 10693 2227 10707
rect 2253 10693 2267 10707
rect 2293 10693 2307 10707
rect 2353 10633 2367 10647
rect 2273 10593 2287 10607
rect 2513 10713 2527 10727
rect 2653 10933 2667 10947
rect 2733 11053 2747 11067
rect 2773 11013 2787 11027
rect 2713 10913 2727 10927
rect 2433 10673 2447 10687
rect 2393 10593 2407 10607
rect 2353 10453 2367 10467
rect 2313 10433 2327 10447
rect 2473 10433 2487 10447
rect 2173 10393 2187 10407
rect 2293 10393 2307 10407
rect 2053 10253 2067 10267
rect 2153 10333 2167 10347
rect 2373 10413 2387 10427
rect 2433 10393 2447 10407
rect 2393 10353 2407 10367
rect 2333 10333 2347 10347
rect 2313 10313 2327 10327
rect 2293 10153 2307 10167
rect 2253 10113 2267 10127
rect 2213 9993 2227 10007
rect 2093 9953 2107 9967
rect 2133 9953 2147 9967
rect 2073 9933 2087 9947
rect 2033 9753 2047 9767
rect 2113 9873 2127 9887
rect 2133 9813 2147 9827
rect 2113 9753 2127 9767
rect 2033 9473 2047 9487
rect 2093 9453 2107 9467
rect 2073 9433 2087 9447
rect 2013 9313 2027 9327
rect 2013 9293 2027 9307
rect 1973 9273 1987 9287
rect 2033 9273 2047 9287
rect 1993 9213 2007 9227
rect 2153 9733 2167 9747
rect 2293 10053 2307 10067
rect 2333 10273 2347 10287
rect 2373 10053 2387 10067
rect 2293 9753 2307 9767
rect 2253 9733 2267 9747
rect 2273 9693 2287 9707
rect 2233 9673 2247 9687
rect 2193 9633 2207 9647
rect 2353 9633 2367 9647
rect 2273 9493 2287 9507
rect 2313 9493 2327 9507
rect 2173 9413 2187 9427
rect 2153 9393 2167 9407
rect 2133 9133 2147 9147
rect 1793 9093 1807 9107
rect 1953 9093 1967 9107
rect 1773 9073 1787 9087
rect 1733 9053 1747 9067
rect 1733 9013 1747 9027
rect 1753 8853 1767 8867
rect 1853 9073 1867 9087
rect 1833 9033 1847 9047
rect 1813 8853 1827 8867
rect 1793 8813 1807 8827
rect 1733 8793 1747 8807
rect 1773 8793 1787 8807
rect 1693 8733 1707 8747
rect 1653 8593 1667 8607
rect 1633 8573 1647 8587
rect 1593 8553 1607 8567
rect 1613 8553 1627 8567
rect 1593 8493 1607 8507
rect 1573 8373 1587 8387
rect 1433 8313 1447 8327
rect 1453 8313 1467 8327
rect 1413 8033 1427 8047
rect 1393 7913 1407 7927
rect 1593 8333 1607 8347
rect 1693 8513 1707 8527
rect 1673 8493 1687 8507
rect 1693 8473 1707 8487
rect 1673 8413 1687 8427
rect 1653 8373 1667 8387
rect 1553 8313 1567 8327
rect 1613 8293 1627 8307
rect 1573 8273 1587 8287
rect 1533 8173 1547 8187
rect 1493 8053 1507 8067
rect 1533 8033 1547 8047
rect 1473 8013 1487 8027
rect 1513 8013 1527 8027
rect 1573 8013 1587 8027
rect 1493 7873 1507 7887
rect 1453 7833 1467 7847
rect 1533 7853 1547 7867
rect 1513 7793 1527 7807
rect 1553 7653 1567 7667
rect 1413 7553 1427 7567
rect 1533 7553 1547 7567
rect 1553 7553 1567 7567
rect 1593 7513 1607 7527
rect 1273 7333 1287 7347
rect 1333 7313 1347 7327
rect 1333 7153 1347 7167
rect 1333 7093 1347 7107
rect 1393 7153 1407 7167
rect 1293 7053 1307 7067
rect 1313 7053 1327 7067
rect 1313 7033 1327 7047
rect 1353 7033 1367 7047
rect 1233 6873 1247 6887
rect 1213 6853 1227 6867
rect 1213 6573 1227 6587
rect 1213 6113 1227 6127
rect 1273 6853 1287 6867
rect 1353 6973 1367 6987
rect 1253 6833 1267 6847
rect 1313 6833 1327 6847
rect 1253 6813 1267 6827
rect 1273 6593 1287 6607
rect 1313 6593 1327 6607
rect 1253 6573 1267 6587
rect 1333 6413 1347 6427
rect 1313 6373 1327 6387
rect 1373 6373 1387 6387
rect 1653 8073 1667 8087
rect 1633 7293 1647 7307
rect 1553 7233 1567 7247
rect 1453 7053 1467 7067
rect 1513 7073 1527 7087
rect 1533 7053 1547 7067
rect 1493 7013 1507 7027
rect 1473 6993 1487 7007
rect 1433 6853 1447 6867
rect 1413 6833 1427 6847
rect 1453 6793 1467 6807
rect 1473 6613 1487 6627
rect 1453 6553 1467 6567
rect 1493 6553 1507 6567
rect 1533 6413 1547 6427
rect 1473 6373 1487 6387
rect 1393 6353 1407 6367
rect 1373 6213 1387 6227
rect 1393 5973 1407 5987
rect 1513 5973 1527 5987
rect 1513 5913 1527 5927
rect 1393 5893 1407 5907
rect 1473 5893 1487 5907
rect 1433 5733 1447 5747
rect 1373 5673 1387 5687
rect 1313 5653 1327 5667
rect 1393 5633 1407 5647
rect 1293 5573 1307 5587
rect 1273 5553 1287 5567
rect 1373 5553 1387 5567
rect 1333 5513 1347 5527
rect 1373 5513 1387 5527
rect 1193 5473 1207 5487
rect 1213 5413 1227 5427
rect 1233 5293 1247 5307
rect 1213 5133 1227 5147
rect 1533 5813 1547 5827
rect 1753 8753 1767 8767
rect 1753 8513 1767 8527
rect 1733 8413 1747 8427
rect 1713 8353 1727 8367
rect 1833 8533 1847 8547
rect 1933 8873 1947 8887
rect 1893 8773 1907 8787
rect 1853 8513 1867 8527
rect 1813 8473 1827 8487
rect 1853 8453 1867 8467
rect 1773 8353 1787 8367
rect 1753 8333 1767 8347
rect 1733 8313 1747 8327
rect 1693 8293 1707 8307
rect 1813 8313 1827 8327
rect 1753 8293 1767 8307
rect 1793 8293 1807 8307
rect 1733 8273 1747 8287
rect 1753 8153 1767 8167
rect 1693 8133 1707 8147
rect 1733 8093 1747 8107
rect 1693 7893 1707 7907
rect 1813 8273 1827 8287
rect 1793 8053 1807 8067
rect 1773 7993 1787 8007
rect 1693 7873 1707 7887
rect 1713 7813 1727 7827
rect 1753 7893 1767 7907
rect 1733 7773 1747 7787
rect 1833 8133 1847 8147
rect 1833 7993 1847 8007
rect 1813 7973 1827 7987
rect 1833 7953 1847 7967
rect 1813 7933 1827 7947
rect 1793 7873 1807 7887
rect 1773 7633 1787 7647
rect 1773 7573 1787 7587
rect 1813 7813 1827 7827
rect 1733 7553 1747 7567
rect 1753 7533 1767 7547
rect 1673 7493 1687 7507
rect 1673 7413 1687 7427
rect 1653 7213 1667 7227
rect 1713 7093 1727 7107
rect 1653 7053 1667 7067
rect 1693 7053 1707 7067
rect 1713 7053 1727 7067
rect 1573 7033 1587 7047
rect 1653 7033 1667 7047
rect 1673 6953 1687 6967
rect 1653 6893 1667 6907
rect 1613 6873 1627 6887
rect 1633 6853 1647 6867
rect 1593 6733 1607 6747
rect 1573 6413 1587 6427
rect 1693 6613 1707 6627
rect 1613 6593 1627 6607
rect 1653 6593 1667 6607
rect 1633 6573 1647 6587
rect 1673 6493 1687 6507
rect 1613 6473 1627 6487
rect 1613 6373 1627 6387
rect 1593 6253 1607 6267
rect 1633 6253 1647 6267
rect 1693 6333 1707 6347
rect 1673 6133 1687 6147
rect 1633 5933 1647 5947
rect 1613 5893 1627 5907
rect 1553 5733 1567 5747
rect 1513 5633 1527 5647
rect 1473 5353 1487 5367
rect 1393 5213 1407 5227
rect 1433 5213 1447 5227
rect 1293 5193 1307 5207
rect 1333 5193 1347 5207
rect 1373 5193 1387 5207
rect 1233 5013 1247 5027
rect 1373 5153 1387 5167
rect 1353 5133 1367 5147
rect 1313 5113 1327 5127
rect 1373 5113 1387 5127
rect 1253 4993 1267 5007
rect 1293 4993 1307 5007
rect 1233 4973 1247 4987
rect 1013 4953 1027 4967
rect 1053 4953 1067 4967
rect 1093 4953 1107 4967
rect 1113 4953 1127 4967
rect 1133 4953 1147 4967
rect 1193 4953 1207 4967
rect 993 4873 1007 4887
rect 833 4713 847 4727
rect 893 4713 907 4727
rect 773 4693 787 4707
rect 833 4633 847 4647
rect 813 4613 827 4627
rect 793 4433 807 4447
rect 953 4553 967 4567
rect 873 4453 887 4467
rect 893 4453 907 4467
rect 853 4413 867 4427
rect 733 4193 747 4207
rect 733 4153 747 4167
rect 653 4073 667 4087
rect 713 4073 727 4087
rect 553 3913 567 3927
rect 493 3733 507 3747
rect 533 3733 547 3747
rect 473 3493 487 3507
rect 453 3473 467 3487
rect 533 3693 547 3707
rect 673 4013 687 4027
rect 853 3993 867 4007
rect 713 3773 727 3787
rect 653 3633 667 3647
rect 653 3613 667 3627
rect 573 3573 587 3587
rect 613 3533 627 3547
rect 573 3513 587 3527
rect 773 3713 787 3727
rect 973 4433 987 4447
rect 1113 4893 1127 4907
rect 1133 4893 1147 4907
rect 1073 4733 1087 4747
rect 1033 4693 1047 4707
rect 1353 4973 1367 4987
rect 1273 4933 1287 4947
rect 1353 4933 1367 4947
rect 1313 4913 1327 4927
rect 1233 4693 1247 4707
rect 1013 4613 1027 4627
rect 1013 4533 1027 4547
rect 1013 4493 1027 4507
rect 1053 4433 1067 4447
rect 1053 4413 1067 4427
rect 953 4233 967 4247
rect 993 4233 1007 4247
rect 933 4133 947 4147
rect 913 3993 927 4007
rect 933 3973 947 3987
rect 993 4213 1007 4227
rect 973 4193 987 4207
rect 993 4133 1007 4147
rect 1033 3993 1047 4007
rect 993 3933 1007 3947
rect 973 3813 987 3827
rect 953 3773 967 3787
rect 913 3733 927 3747
rect 953 3733 967 3747
rect 893 3713 907 3727
rect 933 3713 947 3727
rect 873 3693 887 3707
rect 873 3653 887 3667
rect 753 3553 767 3567
rect 733 3533 747 3547
rect 813 3533 827 3547
rect 593 3493 607 3507
rect 833 3513 847 3527
rect 953 3633 967 3647
rect 513 3473 527 3487
rect 633 3473 647 3487
rect 913 3513 927 3527
rect 893 3433 907 3447
rect 853 3413 867 3427
rect 573 3373 587 3387
rect 773 3373 787 3387
rect 513 3253 527 3267
rect 853 3233 867 3247
rect 673 3193 687 3207
rect 553 3173 567 3187
rect 493 3093 507 3107
rect 433 3033 447 3047
rect 453 3033 467 3047
rect 513 3033 527 3047
rect 913 3193 927 3207
rect 893 3133 907 3147
rect 753 3053 767 3067
rect 893 3033 907 3047
rect 493 3013 507 3027
rect 633 3013 647 3027
rect 933 3013 947 3027
rect 453 2993 467 3007
rect 1013 3873 1027 3887
rect 1013 3793 1027 3807
rect 1113 4573 1127 4587
rect 1273 4653 1287 4667
rect 1253 4573 1267 4587
rect 1313 4553 1327 4567
rect 1113 4493 1127 4507
rect 1073 4253 1087 4267
rect 1213 4493 1227 4507
rect 1613 5493 1627 5507
rect 1653 5433 1667 5447
rect 1713 5633 1727 5647
rect 1593 5393 1607 5407
rect 1633 5393 1647 5407
rect 1533 5193 1547 5207
rect 1473 5173 1487 5187
rect 1513 5173 1527 5187
rect 1533 5153 1547 5167
rect 1433 5133 1447 5147
rect 1693 5393 1707 5407
rect 1673 5333 1687 5347
rect 1713 5213 1727 5227
rect 1653 5193 1667 5207
rect 1573 5113 1587 5127
rect 1593 5113 1607 5127
rect 1553 5093 1567 5107
rect 1533 5013 1547 5027
rect 1453 4973 1467 4987
rect 1433 4953 1447 4967
rect 1493 4913 1507 4927
rect 1433 4893 1447 4907
rect 1433 4713 1447 4727
rect 1573 5013 1587 5027
rect 1613 4993 1627 5007
rect 1793 7513 1807 7527
rect 1773 7373 1787 7387
rect 1793 7333 1807 7347
rect 1753 7093 1767 7107
rect 1953 8793 1967 8807
rect 2253 9293 2267 9307
rect 2173 9273 2187 9287
rect 2213 9273 2227 9287
rect 2193 9253 2207 9267
rect 2233 9253 2247 9267
rect 2213 9233 2227 9247
rect 2193 9093 2207 9107
rect 2173 8993 2187 9007
rect 2033 8813 2047 8827
rect 1933 8753 1947 8767
rect 1953 8733 1967 8747
rect 1913 8513 1927 8527
rect 1933 8493 1947 8507
rect 2013 8773 2027 8787
rect 1973 8533 1987 8547
rect 1993 8513 2007 8527
rect 2033 8513 2047 8527
rect 1973 8493 1987 8507
rect 1933 8313 1947 8327
rect 1893 8273 1907 8287
rect 1913 8273 1927 8287
rect 1933 8113 1947 8127
rect 1913 8053 1927 8067
rect 1953 8053 1967 8067
rect 1873 8013 1887 8027
rect 1853 7873 1867 7887
rect 1933 8013 1947 8027
rect 1893 7853 1907 7867
rect 1913 7853 1927 7867
rect 1953 7853 1967 7867
rect 1873 7833 1887 7847
rect 1993 8473 2007 8487
rect 2033 8493 2047 8507
rect 2013 8453 2027 8467
rect 2013 8253 2027 8267
rect 1993 8113 2007 8127
rect 2013 8113 2027 8127
rect 2013 8093 2027 8107
rect 1993 8013 2007 8027
rect 1993 7913 2007 7927
rect 1853 7813 1867 7827
rect 1873 7793 1887 7807
rect 1853 7333 1867 7347
rect 1833 7233 1847 7247
rect 1873 7233 1887 7247
rect 1813 7213 1827 7227
rect 1933 7813 1947 7827
rect 1973 7813 1987 7827
rect 1993 7553 2007 7567
rect 1933 7533 1947 7547
rect 1973 7533 1987 7547
rect 1953 7513 1967 7527
rect 2053 8233 2067 8247
rect 2073 8133 2087 8147
rect 2093 8113 2107 8127
rect 2113 8113 2127 8127
rect 2153 8813 2167 8827
rect 2193 8513 2207 8527
rect 2233 9113 2247 9127
rect 2253 8993 2267 9007
rect 2293 8993 2307 9007
rect 2273 8913 2287 8927
rect 2253 8833 2267 8847
rect 2213 8493 2227 8507
rect 2233 8493 2247 8507
rect 2173 8473 2187 8487
rect 2233 8373 2247 8387
rect 2173 8353 2187 8367
rect 2193 8333 2207 8347
rect 2173 8313 2187 8327
rect 2233 8273 2247 8287
rect 2113 8033 2127 8047
rect 2133 8033 2147 8047
rect 2093 7993 2107 8007
rect 2033 7953 2047 7967
rect 2053 7953 2067 7967
rect 2033 7853 2047 7867
rect 1953 7493 1967 7507
rect 2013 7493 2027 7507
rect 1933 7453 1947 7467
rect 1933 7373 1947 7387
rect 1893 7173 1907 7187
rect 1893 7153 1907 7167
rect 1833 7053 1847 7067
rect 1933 7293 1947 7307
rect 1913 7053 1927 7067
rect 1853 7033 1867 7047
rect 1793 6953 1807 6967
rect 1813 6933 1827 6947
rect 1893 6913 1907 6927
rect 1833 6893 1847 6907
rect 1873 6833 1887 6847
rect 1793 6613 1807 6627
rect 1833 6613 1847 6627
rect 1753 6413 1767 6427
rect 1773 6313 1787 6327
rect 1873 6593 1887 6607
rect 1853 6573 1867 6587
rect 1813 6473 1827 6487
rect 1833 6353 1847 6367
rect 1813 6313 1827 6327
rect 1813 6273 1827 6287
rect 1753 6173 1767 6187
rect 1793 6173 1807 6187
rect 1813 6173 1827 6187
rect 1833 6173 1847 6187
rect 1793 6133 1807 6147
rect 1813 6093 1827 6107
rect 1813 5973 1827 5987
rect 1833 5873 1847 5887
rect 1753 5633 1767 5647
rect 1793 5633 1807 5647
rect 1733 5173 1747 5187
rect 1833 5613 1847 5627
rect 1793 5453 1807 5467
rect 1753 5153 1767 5167
rect 1833 5413 1847 5427
rect 1913 6873 1927 6887
rect 1913 6793 1927 6807
rect 1973 7313 1987 7327
rect 2073 7913 2087 7927
rect 2113 7913 2127 7927
rect 2133 7833 2147 7847
rect 2113 7793 2127 7807
rect 2133 7773 2147 7787
rect 2053 7713 2067 7727
rect 2333 9313 2347 9327
rect 2313 8933 2327 8947
rect 2333 8873 2347 8887
rect 2473 10373 2487 10387
rect 2473 10193 2487 10207
rect 2473 9993 2487 10007
rect 2433 9953 2447 9967
rect 2513 10433 2527 10447
rect 2633 10413 2647 10427
rect 2533 10393 2547 10407
rect 2733 10813 2747 10827
rect 2953 11833 2967 11847
rect 3153 11853 3167 11867
rect 3113 11793 3127 11807
rect 2993 11733 3007 11747
rect 2933 11653 2947 11667
rect 2953 11653 2967 11667
rect 2913 11533 2927 11547
rect 3073 11713 3087 11727
rect 3033 11653 3047 11667
rect 3053 11633 3067 11647
rect 3033 11533 3047 11547
rect 3013 11473 3027 11487
rect 2953 11413 2967 11427
rect 3053 11473 3067 11487
rect 2933 11393 2947 11407
rect 2973 11393 2987 11407
rect 3293 11853 3307 11867
rect 3253 11733 3267 11747
rect 3193 11713 3207 11727
rect 3233 11653 3247 11667
rect 3253 11633 3267 11647
rect 3253 11573 3267 11587
rect 3453 11753 3467 11767
rect 3413 11693 3427 11707
rect 3453 11693 3467 11707
rect 3313 11673 3327 11687
rect 3313 11653 3327 11667
rect 3153 11433 3167 11447
rect 3053 11393 3067 11407
rect 2913 11333 2927 11347
rect 2873 11213 2887 11227
rect 2833 11193 2847 11207
rect 2913 11193 2927 11207
rect 2893 11173 2907 11187
rect 2993 11373 3007 11387
rect 3113 11353 3127 11367
rect 2993 11293 3007 11307
rect 2973 10973 2987 10987
rect 2793 10773 2807 10787
rect 2913 10933 2927 10947
rect 2913 10913 2927 10927
rect 2873 10893 2887 10907
rect 2933 10893 2947 10907
rect 2893 10873 2907 10887
rect 2973 10893 2987 10907
rect 2953 10853 2967 10867
rect 2873 10773 2887 10787
rect 2873 10733 2887 10747
rect 2813 10713 2827 10727
rect 2853 10713 2867 10727
rect 2693 10693 2707 10707
rect 2753 10693 2767 10707
rect 2693 10453 2707 10467
rect 2893 10713 2907 10727
rect 2973 10713 2987 10727
rect 2833 10653 2847 10667
rect 2773 10453 2787 10467
rect 2893 10673 2907 10687
rect 3053 11213 3067 11227
rect 3013 11053 3027 11067
rect 3013 10693 3027 10707
rect 3033 10673 3047 10687
rect 2993 10613 3007 10627
rect 2933 10453 2947 10467
rect 2893 10433 2907 10447
rect 2913 10413 2927 10427
rect 2673 10373 2687 10387
rect 2653 10313 2667 10327
rect 2793 10273 2807 10287
rect 2813 10273 2827 10287
rect 2913 10253 2927 10267
rect 2953 10213 2967 10227
rect 2573 10053 2587 10067
rect 2533 9953 2547 9967
rect 2673 9993 2687 10007
rect 2493 9933 2507 9947
rect 2633 9953 2647 9967
rect 2713 9953 2727 9967
rect 2453 9913 2467 9927
rect 2613 9933 2627 9947
rect 2693 9913 2707 9927
rect 2593 9893 2607 9907
rect 2633 9873 2647 9887
rect 2553 9773 2567 9787
rect 2393 9733 2407 9747
rect 2373 9493 2387 9507
rect 2453 9493 2467 9507
rect 2533 9473 2547 9487
rect 2453 9433 2467 9447
rect 2433 9373 2447 9387
rect 2373 9353 2387 9367
rect 2473 9333 2487 9347
rect 2533 9333 2547 9347
rect 2453 9273 2467 9287
rect 2413 9253 2427 9267
rect 2513 9253 2527 9267
rect 2493 9213 2507 9227
rect 2493 9073 2507 9087
rect 2413 8993 2427 9007
rect 2473 8993 2487 9007
rect 2433 8973 2447 8987
rect 2393 8953 2407 8967
rect 2493 8973 2507 8987
rect 2533 8973 2547 8987
rect 2573 9733 2587 9747
rect 2773 9873 2787 9887
rect 2613 9473 2627 9487
rect 2653 9453 2667 9467
rect 2593 9433 2607 9447
rect 2773 9733 2787 9747
rect 3213 11393 3227 11407
rect 3153 11373 3167 11387
rect 3153 11333 3167 11347
rect 3133 11293 3147 11307
rect 3133 11273 3147 11287
rect 3153 11233 3167 11247
rect 3073 11133 3087 11147
rect 3213 11373 3227 11387
rect 3193 11153 3207 11167
rect 3133 11113 3147 11127
rect 3193 11113 3207 11127
rect 3173 11093 3187 11107
rect 3073 11053 3087 11067
rect 3113 10913 3127 10927
rect 3153 10913 3167 10927
rect 3133 10893 3147 10907
rect 3093 10873 3107 10887
rect 3113 10873 3127 10887
rect 3073 10653 3087 10667
rect 3073 10453 3087 10467
rect 3133 10733 3147 10747
rect 3133 10613 3147 10627
rect 3093 10433 3107 10447
rect 3053 10293 3067 10307
rect 3033 10253 3047 10267
rect 3113 10393 3127 10407
rect 3053 10213 3067 10227
rect 3073 10213 3087 10227
rect 3093 10213 3107 10227
rect 3013 9933 3027 9947
rect 2833 9913 2847 9927
rect 2993 9913 3007 9927
rect 2973 9893 2987 9907
rect 3013 9873 3027 9887
rect 2913 9533 2927 9547
rect 2773 9373 2787 9387
rect 2713 9353 2727 9367
rect 3013 9433 3027 9447
rect 2973 9293 2987 9307
rect 2593 9273 2607 9287
rect 2793 9273 2807 9287
rect 2633 9133 2647 9147
rect 2413 8933 2427 8947
rect 2473 8933 2487 8947
rect 2353 8813 2367 8827
rect 2333 8793 2347 8807
rect 2293 8333 2307 8347
rect 2373 8533 2387 8547
rect 2453 8773 2467 8787
rect 2593 8933 2607 8947
rect 2513 8793 2527 8807
rect 2533 8773 2547 8787
rect 2413 8513 2427 8527
rect 2333 8473 2347 8487
rect 2313 8293 2327 8307
rect 2353 8433 2367 8447
rect 2393 8373 2407 8387
rect 2373 8333 2387 8347
rect 2353 8293 2367 8307
rect 2233 7993 2247 8007
rect 2253 7993 2267 8007
rect 2213 7913 2227 7927
rect 2173 7693 2187 7707
rect 2153 7613 2167 7627
rect 2213 7593 2227 7607
rect 2173 7553 2187 7567
rect 2113 7513 2127 7527
rect 2193 7493 2207 7507
rect 2353 8233 2367 8247
rect 2293 8013 2307 8027
rect 2433 8253 2447 8267
rect 2573 8733 2587 8747
rect 2493 8513 2507 8527
rect 2453 8213 2467 8227
rect 2413 8173 2427 8187
rect 2453 8173 2467 8187
rect 2393 8133 2407 8147
rect 2273 7873 2287 7887
rect 2313 7873 2327 7887
rect 2273 7833 2287 7847
rect 2333 7853 2347 7867
rect 2513 8493 2527 8507
rect 2533 8493 2547 8507
rect 2613 8773 2627 8787
rect 2553 8473 2567 8487
rect 2593 8433 2607 8447
rect 2613 8373 2627 8387
rect 2593 8333 2607 8347
rect 2553 8313 2567 8327
rect 2613 8293 2627 8307
rect 2573 8273 2587 8287
rect 2553 8213 2567 8227
rect 2513 8193 2527 8207
rect 2493 8153 2507 8167
rect 2453 8093 2467 8107
rect 2513 8093 2527 8107
rect 2473 8053 2487 8067
rect 2413 8033 2427 8047
rect 2493 8033 2507 8047
rect 2513 7973 2527 7987
rect 2473 7833 2487 7847
rect 2553 7833 2567 7847
rect 2413 7813 2427 7827
rect 2393 7773 2407 7787
rect 2453 7793 2467 7807
rect 2493 7793 2507 7807
rect 2293 7613 2307 7627
rect 2373 7573 2387 7587
rect 2353 7533 2367 7547
rect 2393 7533 2407 7547
rect 2293 7493 2307 7507
rect 2233 7433 2247 7447
rect 2333 7473 2347 7487
rect 2293 7413 2307 7427
rect 2133 7333 2147 7347
rect 2073 7153 2087 7167
rect 2033 7133 2047 7147
rect 2033 7073 2047 7087
rect 2113 7113 2127 7127
rect 2053 6993 2067 7007
rect 1953 6973 1967 6987
rect 2033 6933 2047 6947
rect 1933 6553 1947 6567
rect 1993 6873 2007 6887
rect 1973 6833 1987 6847
rect 2013 6833 2027 6847
rect 2033 6833 2047 6847
rect 1993 6793 2007 6807
rect 2093 6773 2107 6787
rect 2033 6613 2047 6627
rect 1993 6593 2007 6607
rect 2033 6593 2047 6607
rect 2013 6533 2027 6547
rect 2053 6493 2067 6507
rect 2233 7133 2247 7147
rect 2273 7093 2287 7107
rect 2253 7033 2267 7047
rect 2233 6913 2247 6927
rect 2193 6893 2207 6907
rect 2273 6873 2287 6887
rect 2233 6853 2247 6867
rect 2213 6833 2227 6847
rect 2173 6813 2187 6827
rect 2273 6733 2287 6747
rect 2193 6633 2207 6647
rect 2233 6633 2247 6647
rect 2293 6613 2307 6627
rect 2193 6573 2207 6587
rect 2253 6573 2267 6587
rect 2213 6553 2227 6567
rect 2153 6533 2167 6547
rect 2133 6453 2147 6467
rect 1993 6433 2007 6447
rect 2173 6373 2187 6387
rect 2173 6313 2187 6327
rect 1973 6253 1987 6267
rect 2013 6253 2027 6267
rect 1993 6113 2007 6127
rect 1933 6093 1947 6107
rect 1973 6093 1987 6107
rect 1953 6073 1967 6087
rect 1993 5973 2007 5987
rect 1973 5613 1987 5627
rect 1893 5593 1907 5607
rect 1933 5593 1947 5607
rect 2133 6113 2147 6127
rect 2273 6533 2287 6547
rect 2233 6453 2247 6467
rect 2213 6213 2227 6227
rect 2113 6073 2127 6087
rect 2033 6013 2047 6027
rect 2153 6013 2167 6027
rect 2213 5993 2227 6007
rect 2213 5913 2227 5927
rect 2193 5873 2207 5887
rect 2273 6413 2287 6427
rect 2313 6473 2327 6487
rect 2293 6373 2307 6387
rect 2273 6133 2287 6147
rect 2233 5773 2247 5787
rect 2293 6113 2307 6127
rect 2353 7033 2367 7047
rect 2393 7333 2407 7347
rect 2533 7773 2547 7787
rect 2493 7673 2507 7687
rect 2553 7653 2567 7667
rect 2493 7613 2507 7627
rect 2553 7613 2567 7627
rect 2473 7573 2487 7587
rect 2453 7533 2467 7547
rect 2533 7553 2547 7567
rect 2593 8213 2607 8227
rect 2613 8153 2627 8167
rect 2593 8053 2607 8067
rect 2593 7553 2607 7567
rect 2493 7433 2507 7447
rect 2433 7153 2447 7167
rect 2473 7153 2487 7167
rect 2413 7133 2427 7147
rect 2373 6973 2387 6987
rect 2393 6893 2407 6907
rect 2373 6793 2387 6807
rect 2413 6773 2427 6787
rect 2393 6753 2407 6767
rect 2393 6673 2407 6687
rect 2373 6653 2387 6667
rect 2373 6573 2387 6587
rect 2433 6633 2447 6647
rect 2453 6573 2467 6587
rect 2433 6433 2447 6447
rect 2473 6393 2487 6407
rect 2333 6333 2347 6347
rect 2333 6253 2347 6267
rect 2453 6253 2467 6267
rect 2333 6133 2347 6147
rect 2373 6133 2387 6147
rect 2573 7513 2587 7527
rect 2573 7433 2587 7447
rect 2573 7393 2587 7407
rect 2533 7373 2547 7387
rect 2513 7333 2527 7347
rect 2933 9233 2947 9247
rect 2953 9093 2967 9107
rect 2993 9233 3007 9247
rect 2993 9113 3007 9127
rect 2773 9073 2787 9087
rect 2953 9073 2967 9087
rect 2973 9073 2987 9087
rect 2993 9013 3007 9027
rect 2813 8993 2827 9007
rect 2753 8973 2767 8987
rect 2653 8953 2667 8967
rect 2753 8773 2767 8787
rect 2693 8753 2707 8767
rect 2733 8753 2747 8767
rect 2713 8733 2727 8747
rect 2693 8613 2707 8627
rect 2693 8493 2707 8507
rect 2673 8453 2687 8467
rect 2653 8413 2667 8427
rect 2653 8313 2667 8327
rect 2653 8253 2667 8267
rect 2653 8153 2667 8167
rect 2653 8113 2667 8127
rect 2693 8293 2707 8307
rect 2673 8073 2687 8087
rect 2693 8073 2707 8087
rect 2673 8053 2687 8067
rect 2773 8493 2787 8507
rect 2753 8353 2767 8367
rect 2733 8333 2747 8347
rect 2733 8213 2747 8227
rect 2733 8113 2747 8127
rect 2653 8033 2667 8047
rect 2733 8033 2747 8047
rect 2653 8013 2667 8027
rect 2693 7873 2707 7887
rect 2633 7853 2647 7867
rect 2733 7833 2747 7847
rect 2673 7813 2687 7827
rect 2633 7733 2647 7747
rect 2633 7713 2647 7727
rect 2633 7693 2647 7707
rect 2553 7313 2567 7327
rect 2613 7313 2627 7327
rect 2533 7113 2547 7127
rect 2533 6573 2547 6587
rect 2513 6473 2527 6487
rect 2413 6173 2427 6187
rect 2433 6133 2447 6147
rect 2353 6113 2367 6127
rect 2393 6113 2407 6127
rect 2453 6113 2467 6127
rect 2353 5933 2367 5947
rect 2393 5913 2407 5927
rect 2393 5853 2407 5867
rect 2593 7273 2607 7287
rect 2573 7153 2587 7167
rect 2613 7133 2627 7147
rect 2593 7093 2607 7107
rect 2653 7553 2667 7567
rect 2693 7553 2707 7567
rect 2733 7553 2747 7567
rect 2713 7533 2727 7547
rect 3093 9953 3107 9967
rect 3093 9733 3107 9747
rect 3073 9533 3087 9547
rect 3093 9473 3107 9487
rect 3193 10913 3207 10927
rect 3173 10893 3187 10907
rect 3233 11333 3247 11347
rect 3213 10853 3227 10867
rect 3193 10793 3207 10807
rect 3433 11673 3447 11687
rect 3433 11633 3447 11647
rect 3433 11613 3447 11627
rect 3373 11493 3387 11507
rect 3693 11893 3707 11907
rect 3773 11893 3787 11907
rect 3813 11893 3827 11907
rect 3613 11813 3627 11827
rect 3493 11773 3507 11787
rect 3473 11613 3487 11627
rect 3453 11513 3467 11527
rect 3333 11413 3347 11427
rect 3313 11393 3327 11407
rect 3353 11353 3367 11367
rect 3373 11353 3387 11367
rect 3313 11193 3327 11207
rect 3273 11133 3287 11147
rect 3253 10893 3267 10907
rect 3233 10753 3247 10767
rect 3273 10753 3287 10767
rect 3393 11293 3407 11307
rect 3433 11293 3447 11307
rect 3433 11253 3447 11267
rect 3433 11193 3447 11207
rect 3573 11753 3587 11767
rect 3633 11653 3647 11667
rect 3533 11533 3547 11547
rect 3533 11473 3547 11487
rect 3593 11573 3607 11587
rect 3613 11553 3627 11567
rect 3593 11533 3607 11547
rect 3553 11453 3567 11467
rect 3553 11413 3567 11427
rect 3493 11373 3507 11387
rect 3393 11133 3407 11147
rect 3313 10953 3327 10967
rect 3373 10953 3387 10967
rect 3333 10913 3347 10927
rect 3313 10893 3327 10907
rect 3233 10733 3247 10747
rect 3293 10733 3307 10747
rect 3273 10713 3287 10727
rect 3293 10713 3307 10727
rect 3213 10693 3227 10707
rect 3293 10673 3307 10687
rect 3373 10873 3387 10887
rect 3513 11193 3527 11207
rect 3573 11153 3587 11167
rect 3553 11053 3567 11067
rect 3513 10933 3527 10947
rect 3653 11473 3667 11487
rect 3633 11253 3647 11267
rect 3793 11853 3807 11867
rect 3753 11753 3767 11767
rect 3733 11653 3747 11667
rect 3773 11653 3787 11667
rect 3993 11773 4007 11787
rect 3973 11673 3987 11687
rect 3913 11653 3927 11667
rect 3953 11653 3967 11667
rect 3873 11633 3887 11647
rect 3813 11553 3827 11567
rect 4133 11893 4147 11907
rect 4153 11873 4167 11887
rect 4493 11873 4507 11887
rect 4533 11873 4547 11887
rect 4573 11873 4587 11887
rect 4313 11853 4327 11867
rect 4193 11833 4207 11847
rect 4333 11833 4347 11847
rect 4133 11773 4147 11787
rect 4293 11713 4307 11727
rect 4293 11693 4307 11707
rect 4013 11673 4027 11687
rect 4073 11673 4087 11687
rect 4113 11673 4127 11687
rect 3913 11533 3927 11547
rect 3933 11533 3947 11547
rect 3953 11533 3967 11547
rect 3773 11473 3787 11487
rect 3713 11373 3727 11387
rect 3753 11373 3767 11387
rect 3733 11353 3747 11367
rect 3733 11273 3747 11287
rect 3733 11233 3747 11247
rect 3713 11213 3727 11227
rect 3633 11193 3647 11207
rect 3693 11193 3707 11207
rect 3613 11093 3627 11107
rect 3693 11173 3707 11187
rect 3673 11153 3687 11167
rect 3753 11213 3767 11227
rect 3673 11113 3687 11127
rect 3653 11093 3667 11107
rect 3633 10973 3647 10987
rect 3333 10833 3347 10847
rect 3453 10833 3467 10847
rect 3373 10733 3387 10747
rect 3433 10733 3447 10747
rect 3253 10633 3267 10647
rect 3173 10473 3187 10487
rect 3153 10233 3167 10247
rect 3253 10453 3267 10467
rect 3253 10293 3267 10307
rect 3233 10193 3247 10207
rect 3233 10053 3247 10067
rect 3173 9993 3187 10007
rect 3213 9953 3227 9967
rect 3313 10233 3327 10247
rect 3393 10713 3407 10727
rect 3453 10713 3467 10727
rect 3473 10713 3487 10727
rect 3413 10673 3427 10687
rect 3473 10453 3487 10467
rect 3393 10313 3407 10327
rect 3633 10773 3647 10787
rect 3533 10733 3547 10747
rect 3513 10413 3527 10427
rect 3453 10253 3467 10267
rect 3433 10233 3447 10247
rect 3473 10233 3487 10247
rect 3413 10213 3427 10227
rect 3453 10193 3467 10207
rect 3613 10713 3627 10727
rect 3573 10693 3587 10707
rect 3553 10353 3567 10367
rect 3533 10293 3547 10307
rect 3373 10173 3387 10187
rect 3313 10013 3327 10027
rect 3453 10013 3467 10027
rect 3313 9913 3327 9927
rect 3553 10033 3567 10047
rect 3493 9933 3507 9947
rect 3533 9933 3547 9947
rect 3473 9913 3487 9927
rect 3533 9873 3547 9887
rect 3293 9853 3307 9867
rect 3333 9853 3347 9867
rect 3353 9853 3367 9867
rect 3453 9853 3467 9867
rect 3213 9773 3227 9787
rect 3253 9773 3267 9787
rect 3213 9733 3227 9747
rect 3233 9733 3247 9747
rect 3133 9573 3147 9587
rect 3233 9473 3247 9487
rect 3053 9453 3067 9467
rect 3013 8953 3027 8967
rect 2973 8913 2987 8927
rect 2873 8813 2887 8827
rect 2833 8793 2847 8807
rect 2853 8793 2867 8807
rect 2833 8753 2847 8767
rect 2853 8633 2867 8647
rect 2813 8553 2827 8567
rect 2793 8353 2807 8367
rect 2853 8493 2867 8507
rect 2833 8373 2847 8387
rect 2813 8313 2827 8327
rect 2793 8293 2807 8307
rect 2773 8213 2787 8227
rect 2893 8793 2907 8807
rect 2953 8793 2967 8807
rect 2993 8793 3007 8807
rect 2913 8753 2927 8767
rect 3113 9433 3127 9447
rect 3073 9413 3087 9427
rect 3233 9373 3247 9387
rect 3313 9493 3327 9507
rect 3273 9473 3287 9487
rect 3373 9573 3387 9587
rect 3373 9513 3387 9527
rect 3353 9473 3367 9487
rect 3133 9353 3147 9367
rect 3253 9353 3267 9367
rect 3113 9113 3127 9127
rect 3093 9013 3107 9027
rect 3093 8973 3107 8987
rect 3073 8813 3087 8827
rect 3333 9453 3347 9467
rect 3153 9333 3167 9347
rect 3293 9333 3307 9347
rect 3313 9333 3327 9347
rect 3233 9173 3247 9187
rect 3173 9113 3187 9127
rect 3193 8973 3207 8987
rect 3153 8953 3167 8967
rect 3093 8733 3107 8747
rect 3053 8653 3067 8667
rect 2993 8613 3007 8627
rect 2913 8553 2927 8567
rect 2913 8533 2927 8547
rect 2953 8533 2967 8547
rect 2933 8513 2947 8527
rect 2993 8513 3007 8527
rect 3033 8513 3047 8527
rect 2973 8473 2987 8487
rect 3013 8473 3027 8487
rect 2933 8433 2947 8447
rect 2993 8433 3007 8447
rect 2853 8213 2867 8227
rect 2873 8213 2887 8227
rect 2973 8333 2987 8347
rect 2953 8313 2967 8327
rect 2993 8213 3007 8227
rect 2973 8193 2987 8207
rect 2793 8053 2807 8067
rect 2773 7773 2787 7787
rect 2753 7473 2767 7487
rect 2753 7393 2767 7407
rect 2713 7373 2727 7387
rect 2773 7373 2787 7387
rect 2733 7333 2747 7347
rect 2773 7333 2787 7347
rect 2693 7313 2707 7327
rect 2673 7293 2687 7307
rect 2913 8073 2927 8087
rect 2833 8053 2847 8067
rect 2853 7953 2867 7967
rect 2833 7893 2847 7907
rect 2813 7813 2827 7827
rect 2813 7333 2827 7347
rect 2813 7313 2827 7327
rect 2713 7153 2727 7167
rect 2793 7153 2807 7167
rect 2653 7073 2667 7087
rect 2633 7013 2647 7027
rect 2613 6913 2627 6927
rect 2633 6913 2647 6927
rect 2593 6893 2607 6907
rect 2573 6873 2587 6887
rect 2593 6853 2607 6867
rect 2573 6713 2587 6727
rect 2693 6853 2707 6867
rect 2653 6633 2667 6647
rect 2593 6593 2607 6607
rect 2633 6593 2647 6607
rect 2613 6573 2627 6587
rect 2673 6573 2687 6587
rect 2653 6553 2667 6567
rect 2593 6433 2607 6447
rect 2593 6413 2607 6427
rect 2613 6373 2627 6387
rect 2753 7073 2767 7087
rect 2733 7053 2747 7067
rect 2853 7873 2867 7887
rect 2893 8033 2907 8047
rect 2893 7993 2907 8007
rect 2873 7853 2887 7867
rect 2913 7873 2927 7887
rect 2933 7833 2947 7847
rect 2873 7813 2887 7827
rect 2873 7773 2887 7787
rect 2913 7773 2927 7787
rect 2933 7773 2947 7787
rect 2953 7773 2967 7787
rect 2853 7653 2867 7667
rect 2833 7053 2847 7067
rect 2773 7033 2787 7047
rect 2793 7033 2807 7047
rect 2713 6513 2727 6527
rect 2733 6413 2747 6427
rect 2673 6353 2687 6367
rect 2773 6893 2787 6907
rect 2793 6853 2807 6867
rect 2793 6753 2807 6767
rect 2833 6633 2847 6647
rect 2893 7553 2907 7567
rect 2913 7513 2927 7527
rect 3193 8793 3207 8807
rect 3333 9273 3347 9287
rect 3513 9493 3527 9507
rect 3473 9473 3487 9487
rect 3433 9453 3447 9467
rect 3373 9233 3387 9247
rect 3373 9173 3387 9187
rect 3353 8933 3367 8947
rect 3413 8933 3427 8947
rect 3413 8873 3427 8887
rect 3313 8813 3327 8827
rect 3273 8793 3287 8807
rect 3193 8773 3207 8787
rect 3233 8773 3247 8787
rect 3153 8573 3167 8587
rect 3153 8513 3167 8527
rect 3113 8493 3127 8507
rect 3333 8673 3347 8687
rect 3193 8473 3207 8487
rect 3173 8433 3187 8447
rect 3173 8373 3187 8387
rect 3033 8313 3047 8327
rect 3153 8293 3167 8307
rect 3293 8333 3307 8347
rect 3293 8273 3307 8287
rect 3153 8213 3167 8227
rect 3333 8393 3347 8407
rect 3493 9313 3507 9327
rect 3513 9253 3527 9267
rect 3673 10973 3687 10987
rect 3693 10873 3707 10887
rect 3713 10833 3727 10847
rect 3733 10833 3747 10847
rect 3653 10733 3667 10747
rect 3613 10433 3627 10447
rect 3633 10413 3647 10427
rect 3673 10393 3687 10407
rect 3693 10293 3707 10307
rect 3633 10253 3647 10267
rect 3673 10253 3687 10267
rect 3693 10233 3707 10247
rect 3573 9973 3587 9987
rect 3653 10213 3667 10227
rect 3633 10173 3647 10187
rect 3593 9913 3607 9927
rect 3573 9513 3587 9527
rect 3613 9853 3627 9867
rect 3613 9713 3627 9727
rect 3613 9693 3627 9707
rect 3613 9513 3627 9527
rect 3673 9973 3687 9987
rect 3653 9953 3667 9967
rect 3733 10753 3747 10767
rect 3833 11413 3847 11427
rect 3873 11393 3887 11407
rect 3893 11373 3907 11387
rect 3993 11493 4007 11507
rect 3953 11353 3967 11367
rect 3873 11333 3887 11347
rect 3913 11333 3927 11347
rect 3933 11333 3947 11347
rect 3933 11313 3947 11327
rect 3913 11193 3927 11207
rect 3873 11173 3887 11187
rect 3893 11133 3907 11147
rect 3893 11113 3907 11127
rect 3913 11073 3927 11087
rect 3833 10933 3847 10947
rect 3773 10893 3787 10907
rect 3753 10513 3767 10527
rect 3753 10473 3767 10487
rect 3873 10913 3887 10927
rect 3853 10873 3867 10887
rect 3833 10853 3847 10867
rect 3873 10853 3887 10867
rect 3793 10793 3807 10807
rect 3873 10833 3887 10847
rect 4333 11673 4347 11687
rect 4393 11853 4407 11867
rect 4553 11853 4567 11867
rect 4373 11673 4387 11687
rect 4293 11653 4307 11667
rect 4253 11593 4267 11607
rect 4173 11553 4187 11567
rect 4093 11453 4107 11467
rect 4113 11433 4127 11447
rect 4073 11273 4087 11287
rect 4073 11213 4087 11227
rect 4273 11533 4287 11547
rect 4253 11493 4267 11507
rect 4233 11413 4247 11427
rect 4353 11653 4367 11667
rect 4353 11633 4367 11647
rect 4373 11633 4387 11647
rect 4313 11573 4327 11587
rect 4293 11513 4307 11527
rect 4353 11493 4367 11507
rect 4353 11473 4367 11487
rect 4333 11453 4347 11467
rect 4233 11373 4247 11387
rect 4173 11353 4187 11367
rect 4173 11293 4187 11307
rect 4133 11273 4147 11287
rect 4153 11273 4167 11287
rect 4153 11213 4167 11227
rect 4133 11173 4147 11187
rect 4073 11073 4087 11087
rect 4053 11013 4067 11027
rect 4113 10913 4127 10927
rect 4133 10913 4147 10927
rect 4033 10853 4047 10867
rect 4313 11413 4327 11427
rect 4273 11373 4287 11387
rect 4293 11293 4307 11307
rect 4313 11253 4327 11267
rect 4173 11173 4187 11187
rect 4293 11193 4307 11207
rect 4693 11853 4707 11867
rect 4733 11853 4747 11867
rect 4513 11793 4527 11807
rect 4553 11793 4567 11807
rect 4573 11793 4587 11807
rect 4493 11773 4507 11787
rect 4433 11693 4447 11707
rect 4413 11553 4427 11567
rect 4353 11193 4367 11207
rect 4373 11193 4387 11207
rect 4393 11193 4407 11207
rect 4233 11173 4247 11187
rect 4273 11173 4287 11187
rect 4333 11173 4347 11187
rect 4193 11033 4207 11047
rect 4353 11013 4367 11027
rect 4293 10973 4307 10987
rect 4213 10913 4227 10927
rect 4193 10893 4207 10907
rect 4153 10873 4167 10887
rect 4233 10853 4247 10867
rect 4113 10773 4127 10787
rect 3993 10753 4007 10767
rect 4033 10713 4047 10727
rect 4173 10713 4187 10727
rect 4253 10713 4267 10727
rect 4013 10693 4027 10707
rect 4113 10693 4127 10707
rect 4213 10693 4227 10707
rect 4233 10673 4247 10687
rect 3913 10653 3927 10667
rect 3973 10653 3987 10667
rect 3813 10633 3827 10647
rect 3793 10433 3807 10447
rect 3813 10413 3827 10427
rect 3913 10393 3927 10407
rect 3773 10313 3787 10327
rect 3973 10293 3987 10307
rect 3933 10253 3947 10267
rect 3813 10233 3827 10247
rect 3873 10233 3887 10247
rect 3933 10233 3947 10247
rect 4153 10293 4167 10307
rect 4213 10293 4227 10307
rect 4093 10273 4107 10287
rect 3993 10253 4007 10267
rect 4153 10253 4167 10267
rect 4173 10253 4187 10267
rect 3793 10213 3807 10227
rect 3733 9933 3747 9947
rect 3713 9793 3727 9807
rect 3713 9773 3727 9787
rect 3793 9933 3807 9947
rect 3773 9813 3787 9827
rect 3773 9793 3787 9807
rect 3793 9773 3807 9787
rect 3813 9773 3827 9787
rect 3713 9633 3727 9647
rect 3693 9613 3707 9627
rect 3673 9573 3687 9587
rect 3773 9753 3787 9767
rect 3753 9733 3767 9747
rect 3853 9953 3867 9967
rect 3953 10213 3967 10227
rect 4133 10233 4147 10247
rect 4153 10213 4167 10227
rect 4193 10213 4207 10227
rect 4153 9993 4167 10007
rect 3873 9913 3887 9927
rect 3973 9913 3987 9927
rect 4153 9873 4167 9887
rect 4193 9873 4207 9887
rect 3913 9773 3927 9787
rect 4013 9773 4027 9787
rect 3993 9753 4007 9767
rect 3893 9733 3907 9747
rect 3913 9733 3927 9747
rect 3833 9693 3847 9707
rect 3853 9693 3867 9707
rect 3933 9633 3947 9647
rect 3593 9433 3607 9447
rect 3553 9333 3567 9347
rect 3633 9473 3647 9487
rect 3733 9473 3747 9487
rect 3873 9473 3887 9487
rect 3733 9433 3747 9447
rect 3853 9353 3867 9367
rect 3633 9313 3647 9327
rect 3813 9273 3827 9287
rect 3613 9253 3627 9267
rect 3473 9233 3487 9247
rect 3533 9233 3547 9247
rect 3473 9213 3487 9227
rect 3513 9053 3527 9067
rect 3573 8993 3587 9007
rect 3713 8993 3727 9007
rect 3733 8993 3747 9007
rect 3813 8993 3827 9007
rect 3433 8833 3447 8847
rect 3473 8793 3487 8807
rect 3493 8773 3507 8787
rect 3533 8773 3547 8787
rect 3533 8733 3547 8747
rect 3453 8713 3467 8727
rect 3473 8553 3487 8567
rect 3553 8533 3567 8547
rect 3453 8493 3467 8507
rect 3593 8953 3607 8967
rect 3593 8793 3607 8807
rect 3373 8333 3387 8347
rect 3413 8333 3427 8347
rect 3153 8153 3167 8167
rect 3313 8153 3327 8167
rect 3133 8133 3147 8147
rect 3153 8133 3167 8147
rect 3033 8053 3047 8067
rect 3013 8033 3027 8047
rect 2953 7553 2967 7567
rect 2953 7513 2967 7527
rect 3073 7873 3087 7887
rect 3193 8073 3207 8087
rect 3113 7853 3127 7867
rect 3153 7853 3167 7867
rect 3093 7833 3107 7847
rect 3153 7833 3167 7847
rect 3133 7813 3147 7827
rect 3073 7773 3087 7787
rect 3033 7593 3047 7607
rect 3073 7553 3087 7567
rect 2993 7413 3007 7427
rect 2993 7393 3007 7407
rect 2933 7373 2947 7387
rect 2893 7353 2907 7367
rect 2913 7333 2927 7347
rect 2953 7333 2967 7347
rect 2893 7213 2907 7227
rect 2993 7333 3007 7347
rect 2973 7113 2987 7127
rect 2933 7093 2947 7107
rect 2973 7093 2987 7107
rect 3093 7513 3107 7527
rect 3053 7353 3067 7367
rect 2933 7013 2947 7027
rect 2993 7013 3007 7027
rect 2973 6893 2987 6907
rect 2993 6873 3007 6887
rect 2913 6853 2927 6867
rect 2893 6813 2907 6827
rect 2813 6533 2827 6547
rect 2833 6513 2847 6527
rect 2793 6473 2807 6487
rect 2973 6733 2987 6747
rect 2953 6573 2967 6587
rect 2953 6553 2967 6567
rect 2933 6533 2947 6547
rect 2873 6473 2887 6487
rect 2793 6353 2807 6367
rect 2773 6313 2787 6327
rect 2773 6233 2787 6247
rect 2573 6073 2587 6087
rect 2733 6073 2747 6087
rect 2533 5993 2547 6007
rect 2433 5933 2447 5947
rect 2473 5933 2487 5947
rect 2473 5913 2487 5927
rect 2493 5913 2507 5927
rect 2413 5833 2427 5847
rect 2393 5733 2407 5747
rect 2353 5693 2367 5707
rect 2273 5653 2287 5667
rect 2113 5633 2127 5647
rect 2313 5633 2327 5647
rect 2093 5613 2107 5627
rect 2253 5613 2267 5627
rect 2073 5533 2087 5547
rect 2013 5493 2027 5507
rect 2033 5453 2047 5467
rect 1853 5373 1867 5387
rect 1873 5373 1887 5387
rect 1813 5353 1827 5367
rect 1833 5153 1847 5167
rect 1693 5133 1707 5147
rect 1733 5133 1747 5147
rect 1793 5133 1807 5147
rect 1773 5033 1787 5047
rect 1673 4953 1687 4967
rect 1593 4933 1607 4947
rect 1633 4933 1647 4947
rect 2013 5413 2027 5427
rect 1993 5373 2007 5387
rect 1973 5333 1987 5347
rect 1973 5133 1987 5147
rect 1933 5113 1947 5127
rect 1853 5093 1867 5107
rect 1853 4953 1867 4967
rect 1553 4733 1567 4747
rect 1453 4653 1467 4667
rect 1413 4613 1427 4627
rect 1393 4533 1407 4547
rect 1433 4533 1447 4547
rect 1393 4473 1407 4487
rect 1413 4453 1427 4467
rect 1373 4253 1387 4267
rect 1393 4253 1407 4267
rect 1113 4233 1127 4247
rect 1153 4233 1167 4247
rect 1193 4233 1207 4247
rect 1073 4173 1087 4187
rect 1053 3753 1067 3767
rect 1033 3713 1047 3727
rect 1053 3693 1067 3707
rect 1093 4013 1107 4027
rect 1333 4213 1347 4227
rect 1193 4193 1207 4207
rect 1353 4193 1367 4207
rect 1133 4173 1147 4187
rect 1173 4153 1187 4167
rect 1213 4013 1227 4027
rect 1293 4013 1307 4027
rect 1373 4013 1387 4027
rect 1273 3993 1287 4007
rect 1113 3973 1127 3987
rect 1213 3973 1227 3987
rect 1153 3933 1167 3947
rect 1333 3933 1347 3947
rect 1353 3713 1367 3727
rect 1333 3673 1347 3687
rect 1173 3653 1187 3667
rect 1073 3573 1087 3587
rect 1033 3533 1047 3547
rect 1053 3373 1067 3387
rect 1073 3273 1087 3287
rect 1053 3233 1067 3247
rect 993 3113 1007 3127
rect 973 3013 987 3027
rect 1013 3013 1027 3027
rect 593 2773 607 2787
rect 613 2773 627 2787
rect 553 2753 567 2767
rect 753 2753 767 2767
rect 513 2733 527 2747
rect 653 2733 667 2747
rect 573 2693 587 2707
rect 633 2633 647 2647
rect 433 2573 447 2587
rect 393 2553 407 2567
rect 413 2553 427 2567
rect 1253 3593 1267 3607
rect 1213 3553 1227 3567
rect 1153 3473 1167 3487
rect 1193 3473 1207 3487
rect 1373 3653 1387 3667
rect 1513 4433 1527 4447
rect 1873 4793 1887 4807
rect 1873 4673 1887 4687
rect 1913 4653 1927 4667
rect 1693 4633 1707 4647
rect 1913 4613 1927 4627
rect 1653 4593 1667 4607
rect 1633 4573 1647 4587
rect 1953 5093 1967 5107
rect 1953 4993 1967 5007
rect 1973 4953 1987 4967
rect 2133 5573 2147 5587
rect 2293 5513 2307 5527
rect 2173 5473 2187 5487
rect 2093 5213 2107 5227
rect 2033 5173 2047 5187
rect 2133 5173 2147 5187
rect 2213 5433 2227 5447
rect 2193 5173 2207 5187
rect 2033 5133 2047 5147
rect 2093 5113 2107 5127
rect 2173 5133 2187 5147
rect 2153 5033 2167 5047
rect 1993 4893 2007 4907
rect 1973 4853 1987 4867
rect 2073 4933 2087 4947
rect 2133 4933 2147 4947
rect 2053 4913 2067 4927
rect 2013 4793 2027 4807
rect 1953 4733 1967 4747
rect 1933 4573 1947 4587
rect 2153 4913 2167 4927
rect 2093 4893 2107 4907
rect 2153 4693 2167 4707
rect 2213 4693 2227 4707
rect 2073 4673 2087 4687
rect 1793 4553 1807 4567
rect 2053 4553 2067 4567
rect 1653 4453 1667 4467
rect 1693 4453 1707 4467
rect 1773 4453 1787 4467
rect 1633 4433 1647 4447
rect 1593 4373 1607 4387
rect 1573 4313 1587 4327
rect 1553 4253 1567 4267
rect 1453 4233 1467 4247
rect 1513 4213 1527 4227
rect 1533 4193 1547 4207
rect 1453 4093 1467 4107
rect 1513 4033 1527 4047
rect 1493 4013 1507 4027
rect 1433 3973 1447 3987
rect 1473 3853 1487 3867
rect 1673 4313 1687 4327
rect 1733 4333 1747 4347
rect 1753 4313 1767 4327
rect 1653 4193 1667 4207
rect 1713 4213 1727 4227
rect 1693 4193 1707 4207
rect 1673 4173 1687 4187
rect 1693 4013 1707 4027
rect 1733 4013 1747 4027
rect 1653 3993 1667 4007
rect 2133 4633 2147 4647
rect 2113 4613 2127 4627
rect 2073 4533 2087 4547
rect 2133 4533 2147 4547
rect 1893 4513 1907 4527
rect 2073 4473 2087 4487
rect 1813 4333 1827 4347
rect 1733 3993 1747 4007
rect 1793 3993 1807 4007
rect 1673 3973 1687 3987
rect 1713 3973 1727 3987
rect 1673 3953 1687 3967
rect 1593 3833 1607 3847
rect 1433 3773 1447 3787
rect 1413 3713 1427 3727
rect 1693 3813 1707 3827
rect 1473 3673 1487 3687
rect 1573 3653 1587 3667
rect 1633 3693 1647 3707
rect 1653 3653 1667 3667
rect 1393 3593 1407 3607
rect 1453 3593 1467 3607
rect 1613 3593 1627 3607
rect 1093 3253 1107 3267
rect 1173 3453 1187 3467
rect 1293 3453 1307 3467
rect 1253 3333 1267 3347
rect 1173 3273 1187 3287
rect 1113 3213 1127 3227
rect 1233 3253 1247 3267
rect 1533 3253 1547 3267
rect 1213 3233 1227 3247
rect 1173 3213 1187 3227
rect 1153 3013 1167 3027
rect 1513 3213 1527 3227
rect 1193 3053 1207 3067
rect 1233 3053 1247 3067
rect 1453 3133 1467 3147
rect 1433 3053 1447 3067
rect 1333 3033 1347 3047
rect 1213 3013 1227 3027
rect 1513 3093 1527 3107
rect 1373 3013 1387 3027
rect 1413 3013 1427 3027
rect 1453 3013 1467 3027
rect 1233 2993 1247 3007
rect 1353 2993 1367 3007
rect 1073 2773 1087 2787
rect 1053 2673 1067 2687
rect 953 2653 967 2667
rect 933 2613 947 2627
rect 673 2573 687 2587
rect 893 2573 907 2587
rect 293 2533 307 2547
rect 273 2333 287 2347
rect 133 2313 147 2327
rect 193 2313 207 2327
rect 173 2293 187 2307
rect 113 2053 127 2067
rect 193 2233 207 2247
rect 153 1793 167 1807
rect 133 1773 147 1787
rect 413 2313 427 2327
rect 393 2293 407 2307
rect 293 2233 307 2247
rect 393 2093 407 2107
rect 273 2053 287 2067
rect 633 2553 647 2567
rect 513 2293 527 2307
rect 673 2293 687 2307
rect 513 2253 527 2267
rect 633 2253 647 2267
rect 693 2253 707 2267
rect 953 2573 967 2587
rect 1593 3233 1607 3247
rect 1613 3213 1627 3227
rect 1773 3953 1787 3967
rect 1773 3793 1787 3807
rect 1713 3773 1727 3787
rect 1733 3553 1747 3567
rect 1813 3913 1827 3927
rect 1793 3773 1807 3787
rect 2173 4473 2187 4487
rect 2153 4453 2167 4467
rect 2253 5413 2267 5427
rect 2313 5413 2327 5427
rect 2273 5393 2287 5407
rect 2273 5373 2287 5387
rect 2313 5193 2327 5207
rect 2353 5153 2367 5167
rect 2293 5133 2307 5147
rect 2333 5073 2347 5087
rect 2253 4973 2267 4987
rect 2293 4733 2307 4747
rect 2353 4713 2367 4727
rect 2313 4673 2327 4687
rect 2373 4653 2387 4667
rect 2333 4613 2347 4627
rect 2233 4593 2247 4607
rect 2333 4513 2347 4527
rect 2353 4513 2367 4527
rect 2293 4473 2307 4487
rect 2453 5713 2467 5727
rect 2433 5653 2447 5667
rect 2493 5653 2507 5667
rect 2473 5633 2487 5647
rect 2433 5613 2447 5627
rect 2433 5513 2447 5527
rect 2433 5413 2447 5427
rect 2753 5993 2767 6007
rect 2753 5933 2767 5947
rect 2613 5893 2627 5907
rect 2653 5893 2667 5907
rect 2633 5873 2647 5887
rect 2633 5673 2647 5687
rect 2753 5793 2767 5807
rect 2633 5653 2647 5667
rect 2673 5653 2687 5667
rect 2733 5653 2747 5667
rect 2613 5633 2627 5647
rect 2593 5513 2607 5527
rect 2573 5373 2587 5387
rect 2513 5153 2527 5167
rect 2533 5113 2547 5127
rect 2433 4793 2447 4807
rect 2413 4633 2427 4647
rect 2413 4613 2427 4627
rect 2313 4373 2327 4387
rect 2213 4233 2227 4247
rect 2313 4213 2327 4227
rect 2233 4193 2247 4207
rect 1853 4173 1867 4187
rect 1973 4153 1987 4167
rect 1953 4133 1967 4147
rect 1913 4033 1927 4047
rect 1873 3993 1887 4007
rect 2153 4033 2167 4047
rect 1953 3993 1967 4007
rect 1833 3873 1847 3887
rect 1813 3693 1827 3707
rect 1893 3973 1907 3987
rect 2033 3973 2047 3987
rect 2133 3973 2147 3987
rect 1933 3913 1947 3927
rect 1993 3873 2007 3887
rect 2193 3873 2207 3887
rect 2253 3833 2267 3847
rect 1933 3813 1947 3827
rect 2193 3813 2207 3827
rect 1933 3773 1947 3787
rect 2153 3773 2167 3787
rect 2033 3733 2047 3747
rect 2013 3713 2027 3727
rect 1973 3693 1987 3707
rect 1933 3633 1947 3647
rect 1933 3613 1947 3627
rect 1853 3573 1867 3587
rect 1793 3553 1807 3567
rect 1893 3533 1907 3547
rect 1773 3513 1787 3527
rect 1793 3513 1807 3527
rect 1773 3493 1787 3507
rect 1693 3393 1707 3407
rect 1653 3133 1667 3147
rect 1613 3053 1627 3067
rect 1573 3013 1587 3027
rect 1513 2853 1527 2867
rect 1553 2853 1567 2867
rect 1393 2733 1407 2747
rect 1393 2693 1407 2707
rect 1673 2753 1687 2767
rect 2073 3693 2087 3707
rect 1873 3493 1887 3507
rect 1913 3493 1927 3507
rect 2053 3493 2067 3507
rect 2113 3533 2127 3547
rect 1973 3473 1987 3487
rect 2093 3473 2107 3487
rect 2233 3713 2247 3727
rect 2213 3653 2227 3667
rect 2173 3573 2187 3587
rect 2213 3533 2227 3547
rect 2173 3513 2187 3527
rect 1833 3233 1847 3247
rect 1793 3213 1807 3227
rect 1753 3113 1767 3127
rect 1793 3133 1807 3147
rect 1773 3053 1787 3067
rect 1833 3113 1847 3127
rect 1753 3033 1767 3047
rect 1773 3013 1787 3027
rect 1953 3333 1967 3347
rect 1913 3253 1927 3267
rect 2113 3453 2127 3467
rect 2113 3413 2127 3427
rect 1993 3273 2007 3287
rect 1993 3253 2007 3267
rect 1933 3233 1947 3247
rect 1973 3233 1987 3247
rect 2013 3153 2027 3167
rect 2133 3153 2147 3167
rect 2093 3133 2107 3147
rect 2193 3093 2207 3107
rect 1853 2993 1867 3007
rect 1993 2993 2007 3007
rect 2173 2993 2187 3007
rect 1973 2893 1987 2907
rect 1873 2753 1887 2767
rect 1913 2753 1927 2767
rect 2093 2753 2107 2767
rect 2113 2753 2127 2767
rect 1693 2713 1707 2727
rect 1893 2733 1907 2747
rect 1973 2733 1987 2747
rect 1933 2713 1947 2727
rect 2053 2713 2067 2727
rect 1733 2693 1747 2707
rect 2053 2693 2067 2707
rect 1713 2673 1727 2687
rect 1933 2673 1947 2687
rect 1433 2653 1447 2667
rect 1553 2653 1567 2667
rect 1653 2653 1667 2667
rect 2073 2653 2087 2667
rect 1173 2593 1187 2607
rect 1133 2573 1147 2587
rect 1373 2573 1387 2587
rect 1193 2533 1207 2547
rect 1253 2533 1267 2547
rect 1073 2513 1087 2527
rect 1213 2513 1227 2527
rect 1553 2493 1567 2507
rect 1433 2333 1447 2347
rect 1073 2293 1087 2307
rect 1313 2293 1327 2307
rect 813 2253 827 2267
rect 853 2253 867 2267
rect 893 2253 907 2267
rect 1033 2253 1047 2267
rect 473 2053 487 2067
rect 413 2033 427 2047
rect 153 1653 167 1667
rect 33 1573 47 1587
rect 113 1573 127 1587
rect 313 1813 327 1827
rect 333 1793 347 1807
rect 353 1753 367 1767
rect 593 2093 607 2107
rect 573 2073 587 2087
rect 713 2233 727 2247
rect 753 2233 767 2247
rect 833 2233 847 2247
rect 693 2093 707 2107
rect 493 1793 507 1807
rect 513 1773 527 1787
rect 633 2033 647 2047
rect 593 1813 607 1827
rect 1013 2093 1027 2107
rect 853 2073 867 2087
rect 813 2053 827 2067
rect 833 2033 847 2047
rect 993 2033 1007 2047
rect 453 1733 467 1747
rect 533 1713 547 1727
rect 373 1653 387 1667
rect 273 1573 287 1587
rect 93 1533 107 1547
rect 153 1533 167 1547
rect 213 1533 227 1547
rect 33 1433 47 1447
rect 173 1313 187 1327
rect 133 1153 147 1167
rect 373 1573 387 1587
rect 553 1573 567 1587
rect 733 1813 747 1827
rect 793 1813 807 1827
rect 1253 2253 1267 2267
rect 1193 2233 1207 2247
rect 1293 2233 1307 2247
rect 1133 2093 1147 2107
rect 1173 2093 1187 2107
rect 1233 2093 1247 2107
rect 1253 2093 1267 2107
rect 1153 2073 1167 2087
rect 1193 2073 1207 2087
rect 1233 2033 1247 2047
rect 1133 2013 1147 2027
rect 1513 2113 1527 2127
rect 1353 2053 1367 2067
rect 1373 2033 1387 2047
rect 1473 2073 1487 2087
rect 1573 2293 1587 2307
rect 1393 2013 1407 2027
rect 1413 2013 1427 2027
rect 673 1773 687 1787
rect 713 1773 727 1787
rect 853 1793 867 1807
rect 873 1773 887 1787
rect 853 1753 867 1767
rect 893 1753 907 1767
rect 893 1733 907 1747
rect 1013 1753 1027 1767
rect 913 1693 927 1707
rect 793 1633 807 1647
rect 653 1613 667 1627
rect 773 1613 787 1627
rect 613 1573 627 1587
rect 933 1613 947 1627
rect 1033 1613 1047 1627
rect 953 1593 967 1607
rect 793 1573 807 1587
rect 593 1553 607 1567
rect 473 1433 487 1447
rect 953 1553 967 1567
rect 893 1533 907 1547
rect 353 1293 367 1307
rect 193 1153 207 1167
rect 173 1133 187 1147
rect 233 1133 247 1147
rect 93 1093 107 1107
rect 153 1093 167 1107
rect 193 1093 207 1107
rect 153 833 167 847
rect 93 633 107 647
rect 173 793 187 807
rect 153 653 167 667
rect 193 633 207 647
rect 333 1093 347 1107
rect 373 1093 387 1107
rect 613 1313 627 1327
rect 653 1313 667 1327
rect 693 1313 707 1327
rect 713 1313 727 1327
rect 473 1093 487 1107
rect 513 1093 527 1107
rect 633 1293 647 1307
rect 673 1273 687 1287
rect 693 1113 707 1127
rect 893 1353 907 1367
rect 793 1293 807 1307
rect 933 1293 947 1307
rect 793 1113 807 1127
rect 733 1093 747 1107
rect 753 1093 767 1107
rect 493 1053 507 1067
rect 533 1053 547 1067
rect 593 1053 607 1067
rect 253 853 267 867
rect 233 793 247 807
rect 393 833 407 847
rect 333 793 347 807
rect 353 793 367 807
rect 313 713 327 727
rect 273 673 287 687
rect 253 653 267 667
rect 173 573 187 587
rect 213 573 227 587
rect 173 553 187 567
rect 153 373 167 387
rect 93 353 107 367
rect 133 353 147 367
rect 133 153 147 167
rect 393 793 407 807
rect 473 773 487 787
rect 373 673 387 687
rect 733 1073 747 1087
rect 533 1033 547 1047
rect 693 1033 707 1047
rect 753 853 767 867
rect 573 833 587 847
rect 873 1273 887 1287
rect 913 1273 927 1287
rect 893 1133 907 1147
rect 913 1113 927 1127
rect 1213 1793 1227 1807
rect 1293 1753 1307 1767
rect 1073 1713 1087 1727
rect 1313 1653 1327 1667
rect 1453 1653 1467 1667
rect 1073 1593 1087 1607
rect 1273 1593 1287 1607
rect 1113 1573 1127 1587
rect 1493 1573 1507 1587
rect 1133 1553 1147 1567
rect 1293 1553 1307 1567
rect 1333 1473 1347 1487
rect 1053 1373 1067 1387
rect 1433 1353 1447 1367
rect 1033 1333 1047 1347
rect 1033 1133 1047 1147
rect 1333 1153 1347 1167
rect 993 1113 1007 1127
rect 1233 1133 1247 1147
rect 1113 1113 1127 1127
rect 1213 1113 1227 1127
rect 853 1093 867 1107
rect 953 1093 967 1107
rect 853 1053 867 1067
rect 513 793 527 807
rect 553 753 567 767
rect 733 813 747 827
rect 933 953 947 967
rect 973 853 987 867
rect 1053 1073 1067 1087
rect 1093 1073 1107 1087
rect 1013 1053 1027 1067
rect 953 833 967 847
rect 993 833 1007 847
rect 1113 1033 1127 1047
rect 1073 953 1087 967
rect 1033 853 1047 867
rect 773 793 787 807
rect 853 793 867 807
rect 893 773 907 787
rect 653 753 667 767
rect 853 753 867 767
rect 593 713 607 727
rect 493 673 507 687
rect 373 553 387 567
rect 393 553 407 567
rect 813 593 827 607
rect 793 573 807 587
rect 513 393 527 407
rect 273 373 287 387
rect 253 353 267 367
rect 493 233 507 247
rect 233 113 247 127
rect 373 173 387 187
rect 473 173 487 187
rect 433 153 447 167
rect 293 133 307 147
rect 453 133 467 147
rect 633 373 647 387
rect 553 353 567 367
rect 873 673 887 687
rect 853 373 867 387
rect 1013 673 1027 687
rect 993 653 1007 667
rect 1293 1113 1307 1127
rect 1333 1113 1347 1127
rect 1313 1093 1327 1107
rect 1253 1053 1267 1067
rect 1493 1313 1507 1327
rect 1453 1213 1467 1227
rect 1453 1153 1467 1167
rect 1833 2533 1847 2547
rect 1873 2313 1887 2327
rect 1733 2273 1747 2287
rect 1813 2273 1827 2287
rect 1993 2293 2007 2307
rect 2013 2293 2027 2307
rect 1933 2273 1947 2287
rect 1713 2233 1727 2247
rect 1893 2253 1907 2267
rect 1953 2253 1967 2267
rect 1813 2053 1827 2067
rect 1993 2053 2007 2067
rect 2033 2053 2047 2067
rect 1653 1953 1667 1967
rect 1673 1953 1687 1967
rect 1813 1853 1827 1867
rect 1813 1813 1827 1827
rect 1573 1793 1587 1807
rect 1713 1793 1727 1807
rect 1553 1473 1567 1487
rect 1533 1233 1547 1247
rect 1513 1133 1527 1147
rect 1613 1753 1627 1767
rect 1613 1633 1627 1647
rect 1593 1613 1607 1627
rect 2073 1913 2087 1927
rect 2233 3493 2247 3507
rect 2233 3013 2247 3027
rect 2233 2933 2247 2947
rect 2213 2733 2227 2747
rect 2173 2713 2187 2727
rect 2213 2593 2227 2607
rect 2133 2573 2147 2587
rect 2113 2273 2127 2287
rect 2153 2273 2167 2287
rect 2113 2053 2127 2067
rect 2093 1833 2107 1847
rect 2093 1793 2107 1807
rect 2033 1773 2047 1787
rect 1853 1693 1867 1707
rect 1633 1593 1647 1607
rect 1613 1553 1627 1567
rect 1813 1613 1827 1627
rect 1693 1593 1707 1607
rect 1673 1553 1687 1567
rect 2033 1653 2047 1667
rect 2013 1633 2027 1647
rect 1953 1593 1967 1607
rect 1653 1533 1667 1547
rect 1873 1533 1887 1547
rect 2133 1913 2147 1927
rect 2273 3573 2287 3587
rect 2373 4273 2387 4287
rect 2413 4213 2427 4227
rect 2513 4853 2527 4867
rect 2473 4713 2487 4727
rect 2493 4673 2507 4687
rect 2473 4653 2487 4667
rect 2473 4633 2487 4647
rect 2453 4533 2467 4547
rect 2373 4193 2387 4207
rect 2393 4193 2407 4207
rect 2433 4193 2447 4207
rect 2413 4173 2427 4187
rect 2353 4133 2367 4147
rect 2453 4133 2467 4147
rect 2433 4013 2447 4027
rect 2333 3973 2347 3987
rect 2553 4693 2567 4707
rect 2533 4593 2547 4607
rect 2513 4573 2527 4587
rect 2533 4513 2547 4527
rect 2493 4353 2507 4367
rect 2473 3833 2487 3847
rect 2393 3793 2407 3807
rect 2433 3713 2447 3727
rect 2353 3673 2367 3687
rect 2313 3533 2327 3547
rect 2353 3533 2367 3547
rect 2313 3513 2327 3527
rect 2333 3493 2347 3507
rect 2293 3453 2307 3467
rect 2353 3453 2367 3467
rect 2293 3373 2307 3387
rect 2413 3693 2427 3707
rect 2433 3673 2447 3687
rect 2413 3613 2427 3627
rect 2393 3253 2407 3267
rect 2313 3113 2327 3127
rect 2273 3013 2287 3027
rect 2313 3013 2327 3027
rect 2453 3633 2467 3647
rect 2553 4453 2567 4467
rect 2553 4413 2567 4427
rect 2533 4253 2547 4267
rect 2513 4193 2527 4207
rect 2513 3873 2527 3887
rect 2493 3613 2507 3627
rect 2453 3453 2467 3467
rect 2413 3173 2427 3187
rect 2333 2953 2347 2967
rect 2253 2873 2267 2887
rect 2273 2753 2287 2767
rect 2313 2753 2327 2767
rect 2373 2753 2387 2767
rect 2293 2733 2307 2747
rect 2333 2673 2347 2687
rect 2253 2573 2267 2587
rect 2293 2553 2307 2567
rect 2353 2453 2367 2467
rect 2353 2313 2367 2327
rect 2293 2273 2307 2287
rect 2233 2233 2247 2247
rect 2153 1813 2167 1827
rect 2333 2253 2347 2267
rect 2353 2073 2367 2087
rect 2353 2033 2367 2047
rect 2193 1793 2207 1807
rect 2113 1633 2127 1647
rect 2133 1613 2147 1627
rect 2053 1593 2067 1607
rect 1593 1293 1607 1307
rect 1793 1333 1807 1347
rect 1953 1333 1967 1347
rect 1733 1273 1747 1287
rect 2013 1313 2027 1327
rect 1973 1293 1987 1307
rect 1813 1253 1827 1267
rect 1773 1193 1787 1207
rect 2093 1333 2107 1347
rect 2133 1313 2147 1327
rect 2133 1273 2147 1287
rect 2173 1253 2187 1267
rect 1573 1173 1587 1187
rect 1973 1173 1987 1187
rect 2073 1173 2087 1187
rect 1533 1113 1547 1127
rect 1473 1073 1487 1087
rect 1233 1033 1247 1047
rect 1433 1033 1447 1047
rect 1533 1033 1547 1047
rect 1213 953 1227 967
rect 1293 853 1307 867
rect 1093 773 1107 787
rect 1173 733 1187 747
rect 1033 653 1047 667
rect 1073 653 1087 667
rect 1393 833 1407 847
rect 1293 733 1307 747
rect 1373 673 1387 687
rect 1313 653 1327 667
rect 1033 613 1047 627
rect 1133 613 1147 627
rect 1053 593 1067 607
rect 1273 633 1287 647
rect 1633 853 1647 867
rect 1453 833 1467 847
rect 1473 833 1487 847
rect 1553 833 1567 847
rect 1333 633 1347 647
rect 1373 633 1387 647
rect 953 573 967 587
rect 893 353 907 367
rect 773 333 787 347
rect 713 293 727 307
rect 593 253 607 267
rect 673 253 687 267
rect 513 133 527 147
rect 873 333 887 347
rect 813 233 827 247
rect 993 353 1007 367
rect 953 273 967 287
rect 993 313 1007 327
rect 893 133 907 147
rect 553 113 567 127
rect 1033 113 1047 127
rect 1433 633 1447 647
rect 1393 593 1407 607
rect 1353 573 1367 587
rect 1393 573 1407 587
rect 1153 393 1167 407
rect 1133 333 1147 347
rect 1193 333 1207 347
rect 1393 353 1407 367
rect 1573 813 1587 827
rect 1853 1133 1867 1147
rect 1873 1133 1887 1147
rect 1793 993 1807 1007
rect 1753 933 1767 947
rect 1733 853 1747 867
rect 1613 813 1627 827
rect 1593 773 1607 787
rect 1673 813 1687 827
rect 1653 713 1667 727
rect 1713 713 1727 727
rect 1713 553 1727 567
rect 1553 413 1567 427
rect 1553 353 1567 367
rect 1373 333 1387 347
rect 1413 333 1427 347
rect 1433 333 1447 347
rect 1533 333 1547 347
rect 1573 333 1587 347
rect 1353 313 1367 327
rect 1533 313 1547 327
rect 1173 293 1187 307
rect 1073 273 1087 287
rect 1353 273 1367 287
rect 1713 353 1727 367
rect 1613 333 1627 347
rect 1593 233 1607 247
rect 1193 173 1207 187
rect 1373 133 1387 147
rect 1453 133 1467 147
rect 1593 133 1607 147
rect 1953 1093 1967 1107
rect 1853 933 1867 947
rect 1793 833 1807 847
rect 1773 793 1787 807
rect 1813 773 1827 787
rect 1853 773 1867 787
rect 1773 633 1787 647
rect 1753 613 1767 627
rect 1953 633 1967 647
rect 2153 1133 2167 1147
rect 2053 1113 2067 1127
rect 2033 853 2047 867
rect 2053 853 2067 867
rect 1993 833 2007 847
rect 2013 813 2027 827
rect 2053 813 2067 827
rect 2133 1113 2147 1127
rect 2153 1093 2167 1107
rect 2113 993 2127 1007
rect 2233 1773 2247 1787
rect 2273 1733 2287 1747
rect 2213 1633 2227 1647
rect 2213 1613 2227 1627
rect 2233 1613 2247 1627
rect 2273 1533 2287 1547
rect 2273 1353 2287 1367
rect 2613 5453 2627 5467
rect 2613 5433 2627 5447
rect 2613 5213 2627 5227
rect 2613 4413 2627 4427
rect 2653 5633 2667 5647
rect 2693 5633 2707 5647
rect 2673 5573 2687 5587
rect 2653 5553 2667 5567
rect 2713 5253 2727 5267
rect 2673 5133 2687 5147
rect 2813 6153 2827 6167
rect 2793 5713 2807 5727
rect 2773 5473 2787 5487
rect 2693 5113 2707 5127
rect 2753 5033 2767 5047
rect 2653 5013 2667 5027
rect 2733 5013 2747 5027
rect 2753 5013 2767 5027
rect 2693 4973 2707 4987
rect 2713 4933 2727 4947
rect 2733 4913 2747 4927
rect 2673 4893 2687 4907
rect 2693 4673 2707 4687
rect 2713 4673 2727 4687
rect 2713 4553 2727 4567
rect 2673 4473 2687 4487
rect 2853 6093 2867 6107
rect 2933 6373 2947 6387
rect 2893 6313 2907 6327
rect 2873 6073 2887 6087
rect 2953 6293 2967 6307
rect 2913 6133 2927 6147
rect 2833 5893 2847 5907
rect 2853 5893 2867 5907
rect 2853 5793 2867 5807
rect 2913 5893 2927 5907
rect 2873 5633 2887 5647
rect 2853 5613 2867 5627
rect 2813 5513 2827 5527
rect 2813 5493 2827 5507
rect 2853 5433 2867 5447
rect 2793 5413 2807 5427
rect 2833 5413 2847 5427
rect 2873 5413 2887 5427
rect 2933 5433 2947 5447
rect 2913 5393 2927 5407
rect 2913 5373 2927 5387
rect 2933 5373 2947 5387
rect 2893 5273 2907 5287
rect 2793 5193 2807 5207
rect 2893 5193 2907 5207
rect 2873 5133 2887 5147
rect 2813 4973 2827 4987
rect 2873 4933 2887 4947
rect 2933 5113 2947 5127
rect 2933 4993 2947 5007
rect 2813 4893 2827 4907
rect 2833 4893 2847 4907
rect 2773 4613 2787 4627
rect 2633 4393 2647 4407
rect 2633 4373 2647 4387
rect 2593 4253 2607 4267
rect 2793 4473 2807 4487
rect 2733 4453 2747 4467
rect 2713 4433 2727 4447
rect 2893 4913 2907 4927
rect 2913 4913 2927 4927
rect 2853 4853 2867 4867
rect 2853 4693 2867 4707
rect 2853 4573 2867 4587
rect 2693 4333 2707 4347
rect 2693 4233 2707 4247
rect 2593 4193 2607 4207
rect 2633 4193 2647 4207
rect 2673 4193 2687 4207
rect 2593 4153 2607 4167
rect 2613 4153 2627 4167
rect 2653 4153 2667 4167
rect 2573 4033 2587 4047
rect 2653 4033 2667 4047
rect 2593 3973 2607 3987
rect 2653 3973 2667 3987
rect 2633 3933 2647 3947
rect 2673 3673 2687 3687
rect 2613 3653 2627 3667
rect 2633 3653 2647 3667
rect 2553 3633 2567 3647
rect 2553 3573 2567 3587
rect 2753 4333 2767 4347
rect 2733 4193 2747 4207
rect 2833 4433 2847 4447
rect 2833 4273 2847 4287
rect 2793 4193 2807 4207
rect 2853 4213 2867 4227
rect 2753 4173 2767 4187
rect 2853 4173 2867 4187
rect 2813 4113 2827 4127
rect 2793 4093 2807 4107
rect 2773 4033 2787 4047
rect 2753 4013 2767 4027
rect 2793 3993 2807 4007
rect 2833 3993 2847 4007
rect 2773 3973 2787 3987
rect 2773 3953 2787 3967
rect 2733 3793 2747 3807
rect 2713 3713 2727 3727
rect 2713 3673 2727 3687
rect 2853 3953 2867 3967
rect 2833 3933 2847 3947
rect 2893 4853 2907 4867
rect 2993 6593 3007 6607
rect 2993 6573 3007 6587
rect 2973 6133 2987 6147
rect 3113 7393 3127 7407
rect 3093 7373 3107 7387
rect 3393 8193 3407 8207
rect 3373 8153 3387 8167
rect 3213 8033 3227 8047
rect 3353 8033 3367 8047
rect 3353 7993 3367 8007
rect 3513 8433 3527 8447
rect 3493 8313 3507 8327
rect 3533 8353 3547 8367
rect 3553 8313 3567 8327
rect 3573 8313 3587 8327
rect 3533 8293 3547 8307
rect 3493 8273 3507 8287
rect 3453 8173 3467 8187
rect 3533 8173 3547 8187
rect 3413 8133 3427 8147
rect 3373 7913 3387 7927
rect 3433 7913 3447 7927
rect 3233 7893 3247 7907
rect 3393 7893 3407 7907
rect 3253 7853 3267 7867
rect 3233 7833 3247 7847
rect 3293 7833 3307 7847
rect 3333 7833 3347 7847
rect 3353 7833 3367 7847
rect 3253 7793 3267 7807
rect 3313 7793 3327 7807
rect 3233 7773 3247 7787
rect 3213 7693 3227 7707
rect 3193 7593 3207 7607
rect 3193 7573 3207 7587
rect 3173 7493 3187 7507
rect 3133 7373 3147 7387
rect 3093 7353 3107 7367
rect 3153 7313 3167 7327
rect 3073 7213 3087 7227
rect 3133 7173 3147 7187
rect 3113 7153 3127 7167
rect 3073 7013 3087 7027
rect 3073 6993 3087 7007
rect 3053 6853 3067 6867
rect 3073 6773 3087 6787
rect 3313 7693 3327 7707
rect 3293 7593 3307 7607
rect 3253 7573 3267 7587
rect 3253 7533 3267 7547
rect 3233 7513 3247 7527
rect 3213 7293 3227 7307
rect 3193 7153 3207 7167
rect 3153 7093 3167 7107
rect 3193 7093 3207 7107
rect 3213 7073 3227 7087
rect 3173 7053 3187 7067
rect 3153 6873 3167 6887
rect 3213 6873 3227 6887
rect 3133 6833 3147 6847
rect 3113 6733 3127 6747
rect 3173 6733 3187 6747
rect 3273 7473 3287 7487
rect 3313 7553 3327 7567
rect 3373 7753 3387 7767
rect 3353 7693 3367 7707
rect 3353 7613 3367 7627
rect 3373 7613 3387 7627
rect 3353 7593 3367 7607
rect 3333 7513 3347 7527
rect 3253 7113 3267 7127
rect 3253 7073 3267 7087
rect 3193 6693 3207 6707
rect 3233 6693 3247 6707
rect 3013 6553 3027 6567
rect 3033 6513 3047 6527
rect 3053 6433 3067 6447
rect 3153 6433 3167 6447
rect 3033 6393 3047 6407
rect 3113 6413 3127 6427
rect 3073 6393 3087 6407
rect 3133 6393 3147 6407
rect 3053 6373 3067 6387
rect 3093 6333 3107 6347
rect 3013 6313 3027 6327
rect 3093 6253 3107 6267
rect 2993 6113 3007 6127
rect 3053 6113 3067 6127
rect 3013 6093 3027 6107
rect 3033 6093 3047 6107
rect 2973 6073 2987 6087
rect 3033 6053 3047 6067
rect 3013 6033 3027 6047
rect 3013 5993 3027 6007
rect 3173 6253 3187 6267
rect 3333 7413 3347 7427
rect 3293 7353 3307 7367
rect 3313 7333 3327 7347
rect 3353 7173 3367 7187
rect 3293 7133 3307 7147
rect 3413 7813 3427 7827
rect 3413 7773 3427 7787
rect 3513 8153 3527 8167
rect 3533 8153 3547 8167
rect 3653 8773 3667 8787
rect 3693 8773 3707 8787
rect 3633 8753 3647 8767
rect 3653 8693 3667 8707
rect 3753 8933 3767 8947
rect 3753 8853 3767 8867
rect 3913 9273 3927 9287
rect 3893 9253 3907 9267
rect 3873 9033 3887 9047
rect 3993 9593 4007 9607
rect 3953 9573 3967 9587
rect 3973 9553 3987 9567
rect 3953 9133 3967 9147
rect 3933 9013 3947 9027
rect 3893 8993 3907 9007
rect 3953 8993 3967 9007
rect 3813 8833 3827 8847
rect 3753 8813 3767 8827
rect 3713 8733 3727 8747
rect 3693 8693 3707 8707
rect 3673 8593 3687 8607
rect 3693 8533 3707 8547
rect 3733 8533 3747 8547
rect 3773 8793 3787 8807
rect 3873 8813 3887 8827
rect 3953 8813 3967 8827
rect 3853 8793 3867 8807
rect 3873 8793 3887 8807
rect 3873 8773 3887 8787
rect 3833 8713 3847 8727
rect 3773 8593 3787 8607
rect 3853 8533 3867 8547
rect 3793 8493 3807 8507
rect 3753 8473 3767 8487
rect 3753 8333 3767 8347
rect 3713 8273 3727 8287
rect 3773 8273 3787 8287
rect 3753 8193 3767 8207
rect 3733 8173 3747 8187
rect 3753 8173 3767 8187
rect 3733 8153 3747 8167
rect 3533 8133 3547 8147
rect 3593 8133 3607 8147
rect 3713 8133 3727 8147
rect 3493 7973 3507 7987
rect 3473 7913 3487 7927
rect 3513 7953 3527 7967
rect 3493 7833 3507 7847
rect 3453 7753 3467 7767
rect 3433 7593 3447 7607
rect 3453 7573 3467 7587
rect 3433 7553 3447 7567
rect 3393 7533 3407 7547
rect 3433 7533 3447 7547
rect 3413 7353 3427 7367
rect 3393 7113 3407 7127
rect 3313 7073 3327 7087
rect 3373 7073 3387 7087
rect 3413 7073 3427 7087
rect 3293 7053 3307 7067
rect 3293 6633 3307 6647
rect 3353 7053 3367 7067
rect 3513 7793 3527 7807
rect 3633 8053 3647 8067
rect 3673 7993 3687 8007
rect 3673 7973 3687 7987
rect 3653 7953 3667 7967
rect 3753 7973 3767 7987
rect 3733 7893 3747 7907
rect 3913 8493 3927 8507
rect 3833 8433 3847 8447
rect 3813 8333 3827 8347
rect 3813 8213 3827 8227
rect 3773 7853 3787 7867
rect 3533 7773 3547 7787
rect 3933 8393 3947 8407
rect 3873 8313 3887 8327
rect 4153 9493 4167 9507
rect 4193 9473 4207 9487
rect 4253 10233 4267 10247
rect 4233 10213 4247 10227
rect 4233 10173 4247 10187
rect 4253 9933 4267 9947
rect 4253 9813 4267 9827
rect 4253 9653 4267 9667
rect 4173 9433 4187 9447
rect 4213 9433 4227 9447
rect 4133 9393 4147 9407
rect 4013 9353 4027 9367
rect 4013 9253 4027 9267
rect 4053 9233 4067 9247
rect 4113 9213 4127 9227
rect 4013 9033 4027 9047
rect 4053 9013 4067 9027
rect 4093 9013 4107 9027
rect 4073 8993 4087 9007
rect 3973 8753 3987 8767
rect 4053 8793 4067 8807
rect 4273 9513 4287 9527
rect 4313 10653 4327 10667
rect 4393 11173 4407 11187
rect 4393 11073 4407 11087
rect 4533 11673 4547 11687
rect 4513 11633 4527 11647
rect 4473 11553 4487 11567
rect 4533 11553 4547 11567
rect 4493 11393 4507 11407
rect 4433 11373 4447 11387
rect 4893 11893 4907 11907
rect 4973 11893 4987 11907
rect 4933 11873 4947 11887
rect 4753 11813 4767 11827
rect 4593 11753 4607 11767
rect 4713 11753 4727 11767
rect 4673 11673 4687 11687
rect 4733 11673 4747 11687
rect 4613 11653 4627 11667
rect 4573 11593 4587 11607
rect 4593 11593 4607 11607
rect 4573 11493 4587 11507
rect 4553 11453 4567 11467
rect 4473 11353 4487 11367
rect 4493 11233 4507 11247
rect 4453 11173 4467 11187
rect 4713 11553 4727 11567
rect 4733 11433 4747 11447
rect 4653 11233 4667 11247
rect 4913 11853 4927 11867
rect 4873 11793 4887 11807
rect 4873 11753 4887 11767
rect 4893 11693 4907 11707
rect 5453 11893 5467 11907
rect 5113 11873 5127 11887
rect 5233 11873 5247 11887
rect 5073 11833 5087 11847
rect 4973 11773 4987 11787
rect 5113 11813 5127 11827
rect 5313 11873 5327 11887
rect 5333 11853 5347 11867
rect 5473 11853 5487 11867
rect 5293 11833 5307 11847
rect 5313 11833 5327 11847
rect 5453 11833 5467 11847
rect 5253 11813 5267 11827
rect 5233 11793 5247 11807
rect 5073 11753 5087 11767
rect 4973 11713 4987 11727
rect 4913 11673 4927 11687
rect 4953 11673 4967 11687
rect 5113 11673 5127 11687
rect 5273 11653 5287 11667
rect 4933 11613 4947 11627
rect 4973 11613 4987 11627
rect 5093 11613 5107 11627
rect 4813 11413 4827 11427
rect 4873 11373 4887 11387
rect 4693 11353 4707 11367
rect 4753 11353 4767 11367
rect 4793 11333 4807 11347
rect 4953 11333 4967 11347
rect 4853 11293 4867 11307
rect 4813 11213 4827 11227
rect 4833 11193 4847 11207
rect 4933 11193 4947 11207
rect 4433 11133 4447 11147
rect 4673 11133 4687 11147
rect 4433 11073 4447 11087
rect 4473 11073 4487 11087
rect 4533 11073 4547 11087
rect 4453 11033 4467 11047
rect 4413 11013 4427 11027
rect 4373 10933 4387 10947
rect 4373 10913 4387 10927
rect 4433 10893 4447 10907
rect 4473 10993 4487 11007
rect 4413 10833 4427 10847
rect 4393 10733 4407 10747
rect 4513 10953 4527 10967
rect 4513 10853 4527 10867
rect 4373 10713 4387 10727
rect 4413 10713 4427 10727
rect 4473 10713 4487 10727
rect 4353 10453 4367 10467
rect 4653 11053 4667 11067
rect 4593 10873 4607 10887
rect 4613 10873 4627 10887
rect 4633 10853 4647 10867
rect 4573 10693 4587 10707
rect 4633 10633 4647 10647
rect 4313 10233 4327 10247
rect 4413 10373 4427 10387
rect 4353 10253 4367 10267
rect 4333 10213 4347 10227
rect 4373 10233 4387 10247
rect 4393 10213 4407 10227
rect 4373 9993 4387 10007
rect 4413 9953 4427 9967
rect 4353 9933 4367 9947
rect 4413 9933 4427 9947
rect 4313 9913 4327 9927
rect 4393 9913 4407 9927
rect 4453 9773 4467 9787
rect 4373 9753 4387 9767
rect 4413 9753 4427 9767
rect 4633 10413 4647 10427
rect 4513 10373 4527 10387
rect 4533 10333 4547 10347
rect 4573 10253 4587 10267
rect 4593 10233 4607 10247
rect 4553 10213 4567 10227
rect 4813 10893 4827 10907
rect 5053 11373 5067 11387
rect 5133 11393 5147 11407
rect 5033 11353 5047 11367
rect 5093 11353 5107 11367
rect 5013 11313 5027 11327
rect 5013 11253 5027 11267
rect 4993 11213 5007 11227
rect 4993 11173 5007 11187
rect 5033 11193 5047 11207
rect 5053 11193 5067 11207
rect 4973 11053 4987 11067
rect 5073 11173 5087 11187
rect 5193 11373 5207 11387
rect 5293 11493 5307 11507
rect 5233 11333 5247 11347
rect 5253 11333 5267 11347
rect 5213 11213 5227 11227
rect 5193 11193 5207 11207
rect 5213 11153 5227 11167
rect 5133 11113 5147 11127
rect 5173 11113 5187 11127
rect 5173 11093 5187 11107
rect 5133 11053 5147 11067
rect 5073 10933 5087 10947
rect 5013 10913 5027 10927
rect 5053 10913 5067 10927
rect 4993 10893 5007 10907
rect 4753 10793 4767 10807
rect 4733 10733 4747 10747
rect 4693 10713 4707 10727
rect 4793 10873 4807 10887
rect 5433 11733 5447 11747
rect 5413 11693 5427 11707
rect 5433 11693 5447 11707
rect 5513 11773 5527 11787
rect 5713 11773 5727 11787
rect 5693 11733 5707 11747
rect 5653 11673 5667 11687
rect 5333 11653 5347 11667
rect 5333 11573 5347 11587
rect 5493 11653 5507 11667
rect 5553 11653 5567 11667
rect 5593 11653 5607 11667
rect 5553 11613 5567 11627
rect 5593 11573 5607 11587
rect 5433 11493 5447 11507
rect 5453 11493 5467 11507
rect 5373 11333 5387 11347
rect 5413 11353 5427 11367
rect 5393 11313 5407 11327
rect 5333 11213 5347 11227
rect 5353 11153 5367 11167
rect 5313 11033 5327 11047
rect 5153 10893 5167 10907
rect 5693 11653 5707 11667
rect 5673 11633 5687 11647
rect 5713 11593 5727 11607
rect 5713 11493 5727 11507
rect 5633 11453 5647 11467
rect 5493 11413 5507 11427
rect 5573 11413 5587 11427
rect 5633 11413 5647 11427
rect 5573 11373 5587 11387
rect 5493 11233 5507 11247
rect 5433 11213 5447 11227
rect 5473 11193 5487 11207
rect 4753 10693 4767 10707
rect 4653 10393 4667 10407
rect 4713 10413 4727 10427
rect 4713 10393 4727 10407
rect 4673 10353 4687 10367
rect 4593 10153 4607 10167
rect 4513 9953 4527 9967
rect 4553 9953 4567 9967
rect 4753 10333 4767 10347
rect 4833 10833 4847 10847
rect 5333 10833 5347 10847
rect 5193 10773 5207 10787
rect 4853 10513 4867 10527
rect 4893 10453 4907 10467
rect 4873 10433 4887 10447
rect 4813 10413 4827 10427
rect 5253 10733 5267 10747
rect 5373 10733 5387 10747
rect 5153 10653 5167 10667
rect 4973 10533 4987 10547
rect 4953 10393 4967 10407
rect 4813 10253 4827 10267
rect 4793 10153 4807 10167
rect 4713 9953 4727 9967
rect 4473 9753 4487 9767
rect 4753 9933 4767 9947
rect 4573 9913 4587 9927
rect 4613 9913 4627 9927
rect 4693 9913 4707 9927
rect 4933 9953 4947 9967
rect 5033 10473 5047 10487
rect 5113 10453 5127 10467
rect 5073 10433 5087 10447
rect 5033 10413 5047 10427
rect 4993 10273 5007 10287
rect 5093 10393 5107 10407
rect 5053 10373 5067 10387
rect 5053 10353 5067 10367
rect 5353 10693 5367 10707
rect 5333 10673 5347 10687
rect 5513 11193 5527 11207
rect 5533 11193 5547 11207
rect 5733 11413 5747 11427
rect 6093 11913 6107 11927
rect 6013 11893 6027 11907
rect 6053 11833 6067 11847
rect 6833 11913 6847 11927
rect 7573 11913 7587 11927
rect 8233 11913 8247 11927
rect 8833 11913 8847 11927
rect 6793 11893 6807 11907
rect 6353 11873 6367 11887
rect 6093 11833 6107 11847
rect 6533 11833 6547 11847
rect 6513 11813 6527 11827
rect 6753 11873 6767 11887
rect 6673 11813 6687 11827
rect 6713 11813 6727 11827
rect 5893 11793 5907 11807
rect 5973 11793 5987 11807
rect 6073 11793 6087 11807
rect 6553 11793 6567 11807
rect 5853 11773 5867 11787
rect 5873 11773 5887 11787
rect 5933 11673 5947 11687
rect 5873 11653 5887 11667
rect 5933 11633 5947 11647
rect 5893 11613 5907 11627
rect 5933 11613 5947 11627
rect 5853 11573 5867 11587
rect 5893 11573 5907 11587
rect 5793 11413 5807 11427
rect 5913 11413 5927 11427
rect 6313 11753 6327 11767
rect 6033 11673 6047 11687
rect 6073 11673 6087 11687
rect 6213 11673 6227 11687
rect 6233 11673 6247 11687
rect 6053 11473 6067 11487
rect 5893 11393 5907 11407
rect 5933 11393 5947 11407
rect 5973 11393 5987 11407
rect 6233 11653 6247 11667
rect 6273 11653 6287 11667
rect 6293 11633 6307 11647
rect 6293 11593 6307 11607
rect 6113 11433 6127 11447
rect 6073 11413 6087 11427
rect 6733 11713 6747 11727
rect 6393 11693 6407 11707
rect 6433 11693 6447 11707
rect 6613 11693 6627 11707
rect 5633 11373 5647 11387
rect 5713 11373 5727 11387
rect 5753 11373 5767 11387
rect 6053 11373 6067 11387
rect 5593 11353 5607 11367
rect 5753 11353 5767 11367
rect 6193 11393 6207 11407
rect 5733 11333 5747 11347
rect 6133 11333 6147 11347
rect 6093 11273 6107 11287
rect 6173 11273 6187 11287
rect 5733 11253 5747 11267
rect 5693 11213 5707 11227
rect 5713 11213 5727 11227
rect 5753 11213 5767 11227
rect 5493 11173 5507 11187
rect 5553 11173 5567 11187
rect 5533 11113 5547 11127
rect 5513 10913 5527 10927
rect 5893 11193 5907 11207
rect 5933 11193 5947 11207
rect 5913 11173 5927 11187
rect 5913 11153 5927 11167
rect 5953 11153 5967 11167
rect 5753 11113 5767 11127
rect 5593 10973 5607 10987
rect 5873 10973 5887 10987
rect 5793 10953 5807 10967
rect 5853 10933 5867 10947
rect 5793 10913 5807 10927
rect 5493 10873 5507 10887
rect 5533 10873 5547 10887
rect 5693 10873 5707 10887
rect 5933 10933 5947 10947
rect 5953 10933 5967 10947
rect 5593 10833 5607 10847
rect 5653 10833 5667 10847
rect 5953 10833 5967 10847
rect 5553 10693 5567 10707
rect 5473 10673 5487 10687
rect 5533 10673 5547 10687
rect 6013 11193 6027 11207
rect 6153 11253 6167 11267
rect 6133 11193 6147 11207
rect 6113 11173 6127 11187
rect 6013 11093 6027 11107
rect 6173 11073 6187 11087
rect 6033 10913 6047 10927
rect 6073 10913 6087 10927
rect 6093 10913 6107 10927
rect 6053 10833 6067 10847
rect 6133 10833 6147 10847
rect 6093 10813 6107 10827
rect 5993 10773 6007 10787
rect 6133 10753 6147 10767
rect 5753 10733 5767 10747
rect 5993 10733 6007 10747
rect 5733 10693 5747 10707
rect 5653 10673 5667 10687
rect 5773 10673 5787 10687
rect 5393 10653 5407 10667
rect 5853 10693 5867 10707
rect 5813 10653 5827 10667
rect 5653 10533 5667 10547
rect 5393 10473 5407 10487
rect 5333 10453 5347 10467
rect 5293 10433 5307 10447
rect 5353 10413 5367 10427
rect 5313 10393 5327 10407
rect 5273 10333 5287 10347
rect 5273 10313 5287 10327
rect 5553 10393 5567 10407
rect 5813 10433 5827 10447
rect 5733 10373 5747 10387
rect 5653 10333 5667 10347
rect 5233 10293 5247 10307
rect 5273 10293 5287 10307
rect 5393 10293 5407 10307
rect 5433 10293 5447 10307
rect 5173 10273 5187 10287
rect 5133 10253 5147 10267
rect 5173 10253 5187 10267
rect 5073 10213 5087 10227
rect 5033 10193 5047 10207
rect 5053 10173 5067 10187
rect 4913 9913 4927 9927
rect 4993 9933 5007 9947
rect 4953 9893 4967 9907
rect 4793 9873 4807 9887
rect 4873 9753 4887 9767
rect 4433 9733 4447 9747
rect 4293 9493 4307 9507
rect 4273 9453 4287 9467
rect 4293 9413 4307 9427
rect 4373 9493 4387 9507
rect 4513 9733 4527 9747
rect 4533 9693 4547 9707
rect 4573 9673 4587 9687
rect 4513 9513 4527 9527
rect 4553 9493 4567 9507
rect 4353 9473 4367 9487
rect 4493 9473 4507 9487
rect 4533 9473 4547 9487
rect 4313 9353 4327 9367
rect 4453 9273 4467 9287
rect 4273 9233 4287 9247
rect 4253 9173 4267 9187
rect 4273 9173 4287 9187
rect 4173 8933 4187 8947
rect 4153 8793 4167 8807
rect 4113 8753 4127 8767
rect 4033 8673 4047 8687
rect 4093 8653 4107 8667
rect 4033 8573 4047 8587
rect 4053 8573 4067 8587
rect 4033 8493 4047 8507
rect 4053 8493 4067 8507
rect 4033 8473 4047 8487
rect 3953 8353 3967 8367
rect 4013 8333 4027 8347
rect 3853 8253 3867 8267
rect 3873 8253 3887 8267
rect 3953 8213 3967 8227
rect 3913 8193 3927 8207
rect 3953 8133 3967 8147
rect 3893 8053 3907 8067
rect 3873 8013 3887 8027
rect 3953 7993 3967 8007
rect 3833 7973 3847 7987
rect 3893 7973 3907 7987
rect 3873 7913 3887 7927
rect 3853 7893 3867 7907
rect 3573 7653 3587 7667
rect 3533 7593 3547 7607
rect 3473 7493 3487 7507
rect 3473 7453 3487 7467
rect 3453 7413 3467 7427
rect 3553 7553 3567 7567
rect 3533 7413 3547 7427
rect 3513 7353 3527 7367
rect 3533 7333 3547 7347
rect 3553 7333 3567 7347
rect 3453 7313 3467 7327
rect 3493 7313 3507 7327
rect 3453 7293 3467 7307
rect 3373 7033 3387 7047
rect 3393 7033 3407 7047
rect 3353 7013 3367 7027
rect 3353 6913 3367 6927
rect 3373 6873 3387 6887
rect 3293 6593 3307 6607
rect 3393 6853 3407 6867
rect 3393 6813 3407 6827
rect 3373 6593 3387 6607
rect 3273 6433 3287 6447
rect 3293 6393 3307 6407
rect 3273 6333 3287 6347
rect 3273 6173 3287 6187
rect 3193 6153 3207 6167
rect 3173 6113 3187 6127
rect 3153 6053 3167 6067
rect 3053 6033 3067 6047
rect 3233 6113 3247 6127
rect 3193 6013 3207 6027
rect 3053 5973 3067 5987
rect 3213 5993 3227 6007
rect 3233 5933 3247 5947
rect 2973 5793 2987 5807
rect 3033 5793 3047 5807
rect 3053 5793 3067 5807
rect 3013 5653 3027 5667
rect 3113 5653 3127 5667
rect 3053 5453 3067 5467
rect 3033 5413 3047 5427
rect 3073 5413 3087 5427
rect 3013 5353 3027 5367
rect 3053 5353 3067 5367
rect 2973 5333 2987 5347
rect 3013 5333 3027 5347
rect 2953 4893 2967 4907
rect 2913 4673 2927 4687
rect 3093 5213 3107 5227
rect 3073 5173 3087 5187
rect 3073 5133 3087 5147
rect 3153 5633 3167 5647
rect 3133 5133 3147 5147
rect 3133 5073 3147 5087
rect 3073 4973 3087 4987
rect 3113 4973 3127 4987
rect 3093 4913 3107 4927
rect 3133 4753 3147 4767
rect 3073 4693 3087 4707
rect 3053 4673 3067 4687
rect 3013 4653 3027 4667
rect 3093 4653 3107 4667
rect 3273 6033 3287 6047
rect 3253 5573 3267 5587
rect 3253 5513 3267 5527
rect 3253 5473 3267 5487
rect 3213 5453 3227 5467
rect 3313 6313 3327 6327
rect 3333 6213 3347 6227
rect 3313 5893 3327 5907
rect 3433 6913 3447 6927
rect 3473 7273 3487 7287
rect 3473 7213 3487 7227
rect 3513 7213 3527 7227
rect 3473 7113 3487 7127
rect 3473 6893 3487 6907
rect 3433 6793 3447 6807
rect 3453 6793 3467 6807
rect 3473 6793 3487 6807
rect 3453 6633 3467 6647
rect 3453 6593 3467 6607
rect 3533 7073 3547 7087
rect 3593 7573 3607 7587
rect 3633 7553 3647 7567
rect 3653 7513 3667 7527
rect 3613 7473 3627 7487
rect 3633 7473 3647 7487
rect 3613 7353 3627 7367
rect 3633 7253 3647 7267
rect 3633 7173 3647 7187
rect 3613 7153 3627 7167
rect 3553 7053 3567 7067
rect 3593 7053 3607 7067
rect 3573 7033 3587 7047
rect 3533 6873 3547 6887
rect 3593 6893 3607 6907
rect 3513 6653 3527 6667
rect 3833 7613 3847 7627
rect 3873 7613 3887 7627
rect 3813 7533 3827 7547
rect 3933 7893 3947 7907
rect 3933 7833 3947 7847
rect 4073 8453 4087 8467
rect 4073 8353 4087 8367
rect 4193 8853 4207 8867
rect 4233 8793 4247 8807
rect 4253 8773 4267 8787
rect 4213 8713 4227 8727
rect 4173 8633 4187 8647
rect 4333 8793 4347 8807
rect 4313 8753 4327 8767
rect 4313 8533 4327 8547
rect 4213 8453 4227 8467
rect 4153 8333 4167 8347
rect 4213 8333 4227 8347
rect 4253 8333 4267 8347
rect 4073 8293 4087 8307
rect 4053 8213 4067 8227
rect 4133 8293 4147 8307
rect 4193 8313 4207 8327
rect 4233 8313 4247 8327
rect 4213 8293 4227 8307
rect 4213 8253 4227 8267
rect 4173 8213 4187 8227
rect 4133 8193 4147 8207
rect 4093 8073 4107 8087
rect 4073 8033 4087 8047
rect 4013 8013 4027 8027
rect 4033 8013 4047 8027
rect 4013 7973 4027 7987
rect 4053 7913 4067 7927
rect 4093 8013 4107 8027
rect 4113 7953 4127 7967
rect 4073 7873 4087 7887
rect 4033 7813 4047 7827
rect 3973 7793 3987 7807
rect 3993 7793 4007 7807
rect 3913 7753 3927 7767
rect 3953 7753 3967 7767
rect 3693 7413 3707 7427
rect 3733 7393 3747 7407
rect 3673 7373 3687 7387
rect 3733 7373 3747 7387
rect 3693 7353 3707 7367
rect 3793 7353 3807 7367
rect 3713 7333 3727 7347
rect 3713 7213 3727 7227
rect 3713 7193 3727 7207
rect 3653 7153 3667 7167
rect 3673 7153 3687 7167
rect 3693 7133 3707 7147
rect 3653 7053 3667 7067
rect 3693 7053 3707 7067
rect 3633 6873 3647 6887
rect 3553 6593 3567 6607
rect 3393 6213 3407 6227
rect 3533 6573 3547 6587
rect 3473 6473 3487 6487
rect 3493 6473 3507 6487
rect 3513 6433 3527 6447
rect 3473 6413 3487 6427
rect 3433 6353 3447 6367
rect 3473 6353 3487 6367
rect 3413 6153 3427 6167
rect 3433 6153 3447 6167
rect 3353 5873 3367 5887
rect 3413 6053 3427 6067
rect 3393 5953 3407 5967
rect 3553 6473 3567 6487
rect 3573 6433 3587 6447
rect 3553 6413 3567 6427
rect 3533 6353 3547 6367
rect 3553 6333 3567 6347
rect 3493 5973 3507 5987
rect 3513 5973 3527 5987
rect 3453 5933 3467 5947
rect 3393 5913 3407 5927
rect 3533 5913 3547 5927
rect 3573 6053 3587 6067
rect 3573 5993 3587 6007
rect 3393 5893 3407 5907
rect 3293 5573 3307 5587
rect 3193 5413 3207 5427
rect 3233 5413 3247 5427
rect 3273 5413 3287 5427
rect 3193 5373 3207 5387
rect 3173 4873 3187 4887
rect 3173 4713 3187 4727
rect 3213 5353 3227 5367
rect 3293 5393 3307 5407
rect 3233 5253 3247 5267
rect 3373 5753 3387 5767
rect 3333 5733 3347 5747
rect 3353 5633 3367 5647
rect 3513 5893 3527 5907
rect 3553 5893 3567 5907
rect 3513 5873 3527 5887
rect 3513 5813 3527 5827
rect 3553 5813 3567 5827
rect 3613 6433 3627 6447
rect 3653 6813 3667 6827
rect 3653 6773 3667 6787
rect 3653 6713 3667 6727
rect 3673 6713 3687 6727
rect 3693 6653 3707 6667
rect 3793 7193 3807 7207
rect 3793 7153 3807 7167
rect 3753 7093 3767 7107
rect 3753 7073 3767 7087
rect 3873 7413 3887 7427
rect 3833 7113 3847 7127
rect 3733 7053 3747 7067
rect 3773 7033 3787 7047
rect 3833 7073 3847 7087
rect 3833 6893 3847 6907
rect 3773 6853 3787 6867
rect 3773 6813 3787 6827
rect 3733 6733 3747 6747
rect 3753 6613 3767 6627
rect 3713 6593 3727 6607
rect 3693 6573 3707 6587
rect 3753 6573 3767 6587
rect 3653 6533 3667 6547
rect 3653 6493 3667 6507
rect 3713 6493 3727 6507
rect 3693 6473 3707 6487
rect 3653 6453 3667 6467
rect 3633 6393 3647 6407
rect 3613 6373 3627 6387
rect 3653 6373 3667 6387
rect 3673 6333 3687 6347
rect 3633 6293 3647 6307
rect 3673 6293 3687 6307
rect 3693 6253 3707 6267
rect 3693 6193 3707 6207
rect 3613 6133 3627 6147
rect 3633 6093 3647 6107
rect 3613 5973 3627 5987
rect 3593 5853 3607 5867
rect 3653 5953 3667 5967
rect 3673 5893 3687 5907
rect 3753 6453 3767 6467
rect 3733 6393 3747 6407
rect 3573 5793 3587 5807
rect 3613 5793 3627 5807
rect 3453 5633 3467 5647
rect 3533 5633 3547 5647
rect 3593 5573 3607 5587
rect 3393 5493 3407 5507
rect 3453 5453 3467 5467
rect 3433 5433 3447 5447
rect 3313 5333 3327 5347
rect 3593 5373 3607 5387
rect 3433 5313 3447 5327
rect 3533 5313 3547 5327
rect 3553 5313 3567 5327
rect 3433 5293 3447 5307
rect 3293 5173 3307 5187
rect 3353 5173 3367 5187
rect 3313 5153 3327 5167
rect 3293 5133 3307 5147
rect 3333 5133 3347 5147
rect 3273 5093 3287 5107
rect 3473 5173 3487 5187
rect 3473 5153 3487 5167
rect 3513 5153 3527 5167
rect 3433 5133 3447 5147
rect 3493 5113 3507 5127
rect 3413 5093 3427 5107
rect 3213 5033 3227 5047
rect 3233 4973 3247 4987
rect 3273 4953 3287 4967
rect 3213 4933 3227 4947
rect 3253 4933 3267 4947
rect 3313 4773 3327 4787
rect 3453 4933 3467 4947
rect 3513 4853 3527 4867
rect 3413 4833 3427 4847
rect 3333 4713 3347 4727
rect 3193 4693 3207 4707
rect 3493 4693 3507 4707
rect 3213 4673 3227 4687
rect 3233 4653 3247 4667
rect 3053 4593 3067 4607
rect 3133 4593 3147 4607
rect 3153 4593 3167 4607
rect 2953 4573 2967 4587
rect 2933 4533 2947 4547
rect 2953 4513 2967 4527
rect 2993 4513 3007 4527
rect 2973 4473 2987 4487
rect 2993 4433 3007 4447
rect 2973 4393 2987 4407
rect 3113 4533 3127 4547
rect 3153 4513 3167 4527
rect 3093 4453 3107 4467
rect 3213 4453 3227 4467
rect 3133 4433 3147 4447
rect 3053 4253 3067 4267
rect 3273 4593 3287 4607
rect 3013 4233 3027 4247
rect 3153 4233 3167 4247
rect 3213 4233 3227 4247
rect 2993 4173 3007 4187
rect 3053 4173 3067 4187
rect 2933 4093 2947 4107
rect 2873 3913 2887 3927
rect 2733 3613 2747 3627
rect 2753 3593 2767 3607
rect 2733 3573 2747 3587
rect 2713 3553 2727 3567
rect 2733 3513 2747 3527
rect 2693 3473 2707 3487
rect 2533 3353 2547 3367
rect 2673 3353 2687 3367
rect 2493 3333 2507 3347
rect 2633 3113 2647 3127
rect 2473 3093 2487 3107
rect 2593 3073 2607 3087
rect 2653 3073 2667 3087
rect 2653 3013 2667 3027
rect 2613 2953 2627 2967
rect 2733 3073 2747 3087
rect 2673 2793 2687 2807
rect 2453 2693 2467 2707
rect 2493 2713 2507 2727
rect 2493 2693 2507 2707
rect 2473 2613 2487 2627
rect 2433 2553 2447 2567
rect 2693 2773 2707 2787
rect 2673 2733 2687 2747
rect 2633 2713 2647 2727
rect 2533 2633 2547 2647
rect 2633 2633 2647 2647
rect 2573 2553 2587 2567
rect 2453 2533 2467 2547
rect 2513 2453 2527 2467
rect 2413 2253 2427 2267
rect 2513 2233 2527 2247
rect 2493 2213 2507 2227
rect 2533 2213 2547 2227
rect 2413 2093 2427 2107
rect 2393 2073 2407 2087
rect 2473 2053 2487 2067
rect 2453 1993 2467 2007
rect 2373 1973 2387 1987
rect 2413 1973 2427 1987
rect 2393 1953 2407 1967
rect 2373 1793 2387 1807
rect 2433 1793 2447 1807
rect 2413 1653 2427 1667
rect 2413 1633 2427 1647
rect 2393 1613 2407 1627
rect 2433 1613 2447 1627
rect 2653 2533 2667 2547
rect 2713 2753 2727 2767
rect 2713 2573 2727 2587
rect 2693 2513 2707 2527
rect 2673 2273 2687 2287
rect 2573 2233 2587 2247
rect 2553 2173 2567 2187
rect 2553 2113 2567 2127
rect 2593 2073 2607 2087
rect 2693 2013 2707 2027
rect 2553 1753 2567 1767
rect 2533 1673 2547 1687
rect 2613 1673 2627 1687
rect 2473 1653 2487 1667
rect 2393 1573 2407 1587
rect 2413 1373 2427 1387
rect 2433 1373 2447 1387
rect 2353 1313 2367 1327
rect 2273 1293 2287 1307
rect 2333 1293 2347 1307
rect 2373 1293 2387 1307
rect 2353 1273 2367 1287
rect 2333 1253 2347 1267
rect 2293 1133 2307 1147
rect 2273 853 2287 867
rect 2333 853 2347 867
rect 2193 833 2207 847
rect 2313 833 2327 847
rect 2373 833 2387 847
rect 2393 813 2407 827
rect 2073 793 2087 807
rect 2173 793 2187 807
rect 2353 773 2367 787
rect 2213 693 2227 707
rect 2253 693 2267 707
rect 2213 673 2227 687
rect 2013 633 2027 647
rect 1813 593 1827 607
rect 1753 553 1767 567
rect 1813 373 1827 387
rect 1873 373 1887 387
rect 1853 353 1867 367
rect 1733 213 1747 227
rect 1633 173 1647 187
rect 1673 153 1687 167
rect 1653 133 1667 147
rect 1733 133 1747 147
rect 253 13 267 27
rect 293 13 307 27
rect 953 13 967 27
rect 993 13 1007 27
rect 1793 173 1807 187
rect 1833 173 1847 187
rect 1813 133 1827 147
rect 2133 613 2147 627
rect 2133 393 2147 407
rect 2153 293 2167 307
rect 2073 213 2087 227
rect 1973 193 1987 207
rect 1873 113 1887 127
rect 1953 173 1967 187
rect 1993 173 2007 187
rect 1953 133 1967 147
rect 2133 193 2147 207
rect 2093 153 2107 167
rect 2073 133 2087 147
rect 2113 133 2127 147
rect 2113 13 2127 27
rect 2233 353 2247 367
rect 2373 653 2387 667
rect 2353 613 2367 627
rect 2453 1333 2467 1347
rect 2433 833 2447 847
rect 2593 1593 2607 1607
rect 2573 1373 2587 1387
rect 2493 1313 2507 1327
rect 2533 1313 2547 1327
rect 2473 1293 2487 1307
rect 2493 1253 2507 1267
rect 2553 1293 2567 1307
rect 2593 1293 2607 1307
rect 2733 2493 2747 2507
rect 2973 3653 2987 3667
rect 3253 4193 3267 4207
rect 3233 4173 3247 4187
rect 3333 4533 3347 4547
rect 3473 4513 3487 4527
rect 3293 4213 3307 4227
rect 3213 4153 3227 4167
rect 3173 4133 3187 4147
rect 3193 4133 3207 4147
rect 3153 3933 3167 3947
rect 3193 3973 3207 3987
rect 3193 3933 3207 3947
rect 3213 3933 3227 3947
rect 3073 3833 3087 3847
rect 3053 3633 3067 3647
rect 2873 3613 2887 3627
rect 2933 3613 2947 3627
rect 2993 3613 3007 3627
rect 2833 3573 2847 3587
rect 2793 3333 2807 3347
rect 2853 3333 2867 3347
rect 2813 3253 2827 3267
rect 2813 3093 2827 3107
rect 2813 3073 2827 3087
rect 2833 3033 2847 3047
rect 2773 2793 2787 2807
rect 2753 2053 2767 2067
rect 2733 1773 2747 1787
rect 2793 2753 2807 2767
rect 2853 2893 2867 2907
rect 2893 3293 2907 3307
rect 2893 3113 2907 3127
rect 2873 2773 2887 2787
rect 2853 2713 2867 2727
rect 2873 2673 2887 2687
rect 2833 2553 2847 2567
rect 2793 2533 2807 2547
rect 2813 2513 2827 2527
rect 2793 2493 2807 2507
rect 2913 2453 2927 2467
rect 2913 2313 2927 2327
rect 2833 2253 2847 2267
rect 2893 2253 2907 2267
rect 2953 3553 2967 3567
rect 3033 3553 3047 3567
rect 2993 3513 3007 3527
rect 3013 3493 3027 3507
rect 2973 3473 2987 3487
rect 3033 3293 3047 3307
rect 3053 3273 3067 3287
rect 3013 3233 3027 3247
rect 2993 3173 3007 3187
rect 2973 3113 2987 3127
rect 2973 3073 2987 3087
rect 2953 2913 2967 2927
rect 2953 2733 2967 2747
rect 2953 2313 2967 2327
rect 2933 2213 2947 2227
rect 2873 2153 2887 2167
rect 2793 2073 2807 2087
rect 2813 1793 2827 1807
rect 2633 1613 2647 1627
rect 2713 1613 2727 1627
rect 2753 1613 2767 1627
rect 2773 1613 2787 1627
rect 2833 1613 2847 1627
rect 2673 1593 2687 1607
rect 2633 1353 2647 1367
rect 2613 1253 2627 1267
rect 2633 1253 2647 1267
rect 2473 1133 2487 1147
rect 2513 1133 2527 1147
rect 2513 1093 2527 1107
rect 2533 1073 2547 1087
rect 2573 993 2587 1007
rect 2473 853 2487 867
rect 2473 833 2487 847
rect 2533 833 2547 847
rect 2453 813 2467 827
rect 2433 613 2447 627
rect 2593 813 2607 827
rect 2553 753 2567 767
rect 2653 1153 2667 1167
rect 2633 673 2647 687
rect 2533 653 2547 667
rect 2573 633 2587 647
rect 2553 613 2567 627
rect 2553 593 2567 607
rect 2473 573 2487 587
rect 2513 573 2527 587
rect 2433 413 2447 427
rect 2413 373 2427 387
rect 2373 353 2387 367
rect 2393 353 2407 367
rect 2513 333 2527 347
rect 2453 313 2467 327
rect 2413 293 2427 307
rect 2333 213 2347 227
rect 2493 173 2507 187
rect 2453 153 2467 167
rect 2313 133 2327 147
rect 2333 133 2347 147
rect 2473 133 2487 147
rect 2593 413 2607 427
rect 2653 393 2667 407
rect 2613 333 2627 347
rect 2573 313 2587 327
rect 2633 313 2647 327
rect 2553 253 2567 267
rect 2613 253 2627 267
rect 2593 213 2607 227
rect 2573 113 2587 127
rect 2253 13 2267 27
rect 2273 13 2287 27
rect 2313 13 2327 27
rect 2693 1413 2707 1427
rect 2693 1293 2707 1307
rect 2753 1253 2767 1267
rect 2713 1153 2727 1167
rect 2713 1093 2727 1107
rect 2693 1073 2707 1087
rect 2733 1073 2747 1087
rect 2773 1073 2787 1087
rect 2713 1053 2727 1067
rect 2673 213 2687 227
rect 2773 853 2787 867
rect 2753 833 2767 847
rect 2733 793 2747 807
rect 2773 653 2787 667
rect 2833 653 2847 667
rect 2733 633 2747 647
rect 2753 613 2767 627
rect 2793 593 2807 607
rect 2833 553 2847 567
rect 2753 373 2767 387
rect 2793 373 2807 387
rect 2813 353 2827 367
rect 2793 253 2807 267
rect 2873 2053 2887 2067
rect 2893 1953 2907 1967
rect 2893 1853 2907 1867
rect 2873 1773 2887 1787
rect 2913 1793 2927 1807
rect 2993 3013 3007 3027
rect 3093 3713 3107 3727
rect 3113 3673 3127 3687
rect 3173 3713 3187 3727
rect 3233 3813 3247 3827
rect 3233 3733 3247 3747
rect 3273 3973 3287 3987
rect 3373 4253 3387 4267
rect 3353 4193 3367 4207
rect 3313 3993 3327 4007
rect 3413 4213 3427 4227
rect 3393 4193 3407 4207
rect 3473 4193 3487 4207
rect 3373 4173 3387 4187
rect 3433 4173 3447 4187
rect 3353 3973 3367 3987
rect 3353 3913 3367 3927
rect 3293 3813 3307 3827
rect 3293 3733 3307 3747
rect 3333 3733 3347 3747
rect 3253 3653 3267 3667
rect 3313 3713 3327 3727
rect 3273 3573 3287 3587
rect 3193 3533 3207 3547
rect 3233 3533 3247 3547
rect 3193 3513 3207 3527
rect 3173 3493 3187 3507
rect 3213 3493 3227 3507
rect 3173 3373 3187 3387
rect 3173 3293 3187 3307
rect 3113 3253 3127 3267
rect 3133 3253 3147 3267
rect 3113 3233 3127 3247
rect 3213 3233 3227 3247
rect 3273 3493 3287 3507
rect 3193 3213 3207 3227
rect 3233 3213 3247 3227
rect 3113 3193 3127 3207
rect 3133 3113 3147 3127
rect 3073 3013 3087 3027
rect 3413 4153 3427 4167
rect 3393 4133 3407 4147
rect 3373 3753 3387 3767
rect 3593 5213 3607 5227
rect 3553 5153 3567 5167
rect 3593 5133 3607 5147
rect 3653 5633 3667 5647
rect 3633 5433 3647 5447
rect 3653 5393 3667 5407
rect 3633 5373 3647 5387
rect 3713 5873 3727 5887
rect 3793 6713 3807 6727
rect 3833 6853 3847 6867
rect 4033 7773 4047 7787
rect 3993 7613 4007 7627
rect 3973 7593 3987 7607
rect 4073 7753 4087 7767
rect 4073 7613 4087 7627
rect 4093 7553 4107 7567
rect 3973 7453 3987 7467
rect 3973 7393 3987 7407
rect 3953 7373 3967 7387
rect 3993 7373 4007 7387
rect 3953 7353 3967 7367
rect 3893 7333 3907 7347
rect 3893 7253 3907 7267
rect 3873 7033 3887 7047
rect 4053 7513 4067 7527
rect 4093 7473 4107 7487
rect 4053 7433 4067 7447
rect 4113 7433 4127 7447
rect 4033 7373 4047 7387
rect 4013 7313 4027 7327
rect 3933 7193 3947 7207
rect 3993 7173 4007 7187
rect 3953 7073 3967 7087
rect 3913 7053 3927 7067
rect 3933 7013 3947 7027
rect 3953 6893 3967 6907
rect 4193 8033 4207 8047
rect 4193 7993 4207 8007
rect 4153 7953 4167 7967
rect 4153 7913 4167 7927
rect 4313 8313 4327 8327
rect 4293 8293 4307 8307
rect 4273 8113 4287 8127
rect 4233 8073 4247 8087
rect 4173 7833 4187 7847
rect 4213 7833 4227 7847
rect 4213 7813 4227 7827
rect 4193 7793 4207 7807
rect 4313 8073 4327 8087
rect 4293 7853 4307 7867
rect 4253 7773 4267 7787
rect 4233 7753 4247 7767
rect 4233 7573 4247 7587
rect 4273 7553 4287 7567
rect 4173 7513 4187 7527
rect 4213 7533 4227 7547
rect 4253 7533 4267 7547
rect 4253 7513 4267 7527
rect 4293 7513 4307 7527
rect 4193 7473 4207 7487
rect 4173 7433 4187 7447
rect 4113 7373 4127 7387
rect 4133 7373 4147 7387
rect 4093 7353 4107 7367
rect 4213 7353 4227 7367
rect 4293 7473 4307 7487
rect 4413 9013 4427 9027
rect 4533 9013 4547 9027
rect 4373 8993 4387 9007
rect 4473 8993 4487 9007
rect 4433 8853 4447 8867
rect 4953 9733 4967 9747
rect 4713 9593 4727 9607
rect 4633 9513 4647 9527
rect 4673 9513 4687 9527
rect 4613 9353 4627 9367
rect 4673 9493 4687 9507
rect 4933 9513 4947 9527
rect 4833 9493 4847 9507
rect 4893 9493 4907 9507
rect 4753 9473 4767 9487
rect 4733 9453 4747 9467
rect 4633 9313 4647 9327
rect 4673 9293 4687 9307
rect 4653 9273 4667 9287
rect 4633 9233 4647 9247
rect 4573 8953 4587 8967
rect 4493 8873 4507 8887
rect 4413 8633 4427 8647
rect 4373 8553 4387 8567
rect 4593 8613 4607 8627
rect 4553 8593 4567 8607
rect 4453 8513 4467 8527
rect 4433 8473 4447 8487
rect 4453 8473 4467 8487
rect 4513 8373 4527 8387
rect 4353 8293 4367 8307
rect 4493 8293 4507 8307
rect 4333 7793 4347 7807
rect 4333 7773 4347 7787
rect 4393 8273 4407 8287
rect 4473 8273 4487 8287
rect 4533 8293 4547 8307
rect 4573 8313 4587 8327
rect 4413 8113 4427 8127
rect 4553 8093 4567 8107
rect 4513 8053 4527 8067
rect 4613 8553 4627 8567
rect 4713 9253 4727 9267
rect 4733 9233 4747 9247
rect 4913 9473 4927 9487
rect 5073 9913 5087 9927
rect 5113 9853 5127 9867
rect 5253 10233 5267 10247
rect 5193 10173 5207 10187
rect 5353 10273 5367 10287
rect 5273 10133 5287 10147
rect 5433 10253 5447 10267
rect 5473 10233 5487 10247
rect 5413 10213 5427 10227
rect 5673 10293 5687 10307
rect 5513 10193 5527 10207
rect 5453 10093 5467 10107
rect 5653 10193 5667 10207
rect 5193 9893 5207 9907
rect 5613 9953 5627 9967
rect 5473 9913 5487 9927
rect 5493 9913 5507 9927
rect 5593 9913 5607 9927
rect 5293 9853 5307 9867
rect 5353 9853 5367 9867
rect 5173 9813 5187 9827
rect 5313 9813 5327 9827
rect 5133 9733 5147 9747
rect 5073 9713 5087 9727
rect 5113 9613 5127 9627
rect 5113 9513 5127 9527
rect 5073 9473 5087 9487
rect 5053 9453 5067 9467
rect 4933 9413 4947 9427
rect 4873 9313 4887 9327
rect 4853 9293 4867 9307
rect 4913 9233 4927 9247
rect 4893 9053 4907 9067
rect 4833 9013 4847 9027
rect 4853 9013 4867 9027
rect 4873 8993 4887 9007
rect 4693 8973 4707 8987
rect 4633 8513 4647 8527
rect 4853 8773 4867 8787
rect 4893 8773 4907 8787
rect 4773 8753 4787 8767
rect 4773 8733 4787 8747
rect 4733 8693 4747 8707
rect 4713 8593 4727 8607
rect 4713 8493 4727 8507
rect 5033 9253 5047 9267
rect 5073 9253 5087 9267
rect 5113 9253 5127 9267
rect 5093 9233 5107 9247
rect 5113 9213 5127 9227
rect 5113 9013 5127 9027
rect 5033 8993 5047 9007
rect 5073 8993 5087 9007
rect 5053 8973 5067 8987
rect 5293 9753 5307 9767
rect 5213 9493 5227 9507
rect 5213 9473 5227 9487
rect 5253 9453 5267 9467
rect 5293 9453 5307 9467
rect 5253 9313 5267 9327
rect 5273 9293 5287 9307
rect 5293 9273 5307 9287
rect 5173 9033 5187 9047
rect 5153 9013 5167 9027
rect 5273 9253 5287 9267
rect 5293 9053 5307 9067
rect 5133 8953 5147 8967
rect 5033 8893 5047 8907
rect 5133 8893 5147 8907
rect 5013 8853 5027 8867
rect 4953 8793 4967 8807
rect 4953 8733 4967 8747
rect 4873 8613 4887 8627
rect 4973 8553 4987 8567
rect 5053 8733 5067 8747
rect 5053 8613 5067 8627
rect 4753 8493 4767 8507
rect 4813 8493 4827 8507
rect 4893 8493 4907 8507
rect 4913 8493 4927 8507
rect 4813 8473 4827 8487
rect 4873 8473 4887 8487
rect 4733 8453 4747 8467
rect 4793 8453 4807 8467
rect 4673 8313 4687 8327
rect 4693 8293 4707 8307
rect 4733 8293 4747 8307
rect 4913 8453 4927 8467
rect 4873 8433 4887 8447
rect 4893 8433 4907 8447
rect 4893 8413 4907 8427
rect 4593 8273 4607 8287
rect 4593 8093 4607 8107
rect 4513 7953 4527 7967
rect 4533 7813 4547 7827
rect 5033 8493 5047 8507
rect 5073 8553 5087 8567
rect 4993 8453 5007 8467
rect 5053 8453 5067 8467
rect 4953 8413 4967 8427
rect 5053 8293 5067 8307
rect 4973 8193 4987 8207
rect 4893 8133 4907 8147
rect 4753 8053 4767 8067
rect 4893 8053 4907 8067
rect 4733 7993 4747 8007
rect 4673 7933 4687 7947
rect 4713 7933 4727 7947
rect 4633 7853 4647 7867
rect 4393 7793 4407 7807
rect 4453 7793 4467 7807
rect 4513 7793 4527 7807
rect 4553 7793 4567 7807
rect 4593 7793 4607 7807
rect 4373 7773 4387 7787
rect 4373 7613 4387 7627
rect 4353 7553 4367 7567
rect 4413 7693 4427 7707
rect 4393 7573 4407 7587
rect 4373 7513 4387 7527
rect 4333 7473 4347 7487
rect 4313 7373 4327 7387
rect 4353 7373 4367 7387
rect 4333 7353 4347 7367
rect 4173 7333 4187 7347
rect 4113 7213 4127 7227
rect 4033 7193 4047 7207
rect 4193 7133 4207 7147
rect 4053 7093 4067 7107
rect 4033 7033 4047 7047
rect 3853 6813 3867 6827
rect 3973 6873 3987 6887
rect 4013 6873 4027 6887
rect 3973 6813 3987 6827
rect 4013 6813 4027 6827
rect 3913 6713 3927 6727
rect 3813 6693 3827 6707
rect 3933 6693 3947 6707
rect 3873 6633 3887 6647
rect 3833 6593 3847 6607
rect 3913 6613 3927 6627
rect 3853 6573 3867 6587
rect 3893 6573 3907 6587
rect 3913 6553 3927 6567
rect 3913 6533 3927 6547
rect 3853 6473 3867 6487
rect 3813 6433 3827 6447
rect 3873 6373 3887 6387
rect 3833 6293 3847 6307
rect 3773 6253 3787 6267
rect 3873 6213 3887 6227
rect 3793 6113 3807 6127
rect 3833 6113 3847 6127
rect 3753 6073 3767 6087
rect 3793 6073 3807 6087
rect 3773 6053 3787 6067
rect 3753 5973 3767 5987
rect 3853 6093 3867 6107
rect 3813 6053 3827 6067
rect 3773 5833 3787 5847
rect 3853 5933 3867 5947
rect 3813 5893 3827 5907
rect 3793 5713 3807 5727
rect 3733 5653 3747 5667
rect 3773 5653 3787 5667
rect 3693 5633 3707 5647
rect 3673 5313 3687 5327
rect 3713 5493 3727 5507
rect 3753 5553 3767 5567
rect 3733 5433 3747 5447
rect 3713 5413 3727 5427
rect 3753 5413 3767 5427
rect 3753 5393 3767 5407
rect 3693 5173 3707 5187
rect 3653 5153 3667 5167
rect 3693 5153 3707 5167
rect 3733 5153 3747 5167
rect 3633 5113 3647 5127
rect 3673 5133 3687 5147
rect 3673 5113 3687 5127
rect 3713 5113 3727 5127
rect 3633 5033 3647 5047
rect 3653 5033 3667 5047
rect 3653 4953 3667 4967
rect 3653 4713 3667 4727
rect 3613 4633 3627 4647
rect 3613 4573 3627 4587
rect 3653 4493 3667 4507
rect 3553 4213 3567 4227
rect 3613 4213 3627 4227
rect 3653 4213 3667 4227
rect 3493 4133 3507 4147
rect 3493 4013 3507 4027
rect 3453 3973 3467 3987
rect 3433 3913 3447 3927
rect 3413 3893 3427 3907
rect 3453 3873 3467 3887
rect 3373 3453 3387 3467
rect 3413 3413 3427 3427
rect 3353 3253 3367 3267
rect 3393 3233 3407 3247
rect 3353 3133 3367 3147
rect 3333 3093 3347 3107
rect 3353 3053 3367 3067
rect 3293 3013 3307 3027
rect 3333 3013 3347 3027
rect 3053 2993 3067 3007
rect 3113 2993 3127 3007
rect 2993 2833 3007 2847
rect 3313 2993 3327 3007
rect 3293 2973 3307 2987
rect 3173 2913 3187 2927
rect 3153 2793 3167 2807
rect 3133 2773 3147 2787
rect 3233 2793 3247 2807
rect 3013 2753 3027 2767
rect 3053 2713 3067 2727
rect 3213 2733 3227 2747
rect 3033 2593 3047 2607
rect 3093 2593 3107 2607
rect 2993 2573 3007 2587
rect 3013 2293 3027 2307
rect 2973 2253 2987 2267
rect 3193 2573 3207 2587
rect 3133 2493 3147 2507
rect 3053 2293 3067 2307
rect 3033 2273 3047 2287
rect 3033 2253 3047 2267
rect 3013 2233 3027 2247
rect 3073 2233 3087 2247
rect 3113 2253 3127 2267
rect 3213 2553 3227 2567
rect 3633 4173 3647 4187
rect 3633 4033 3647 4047
rect 3753 5093 3767 5107
rect 3733 4973 3747 4987
rect 3713 4913 3727 4927
rect 3693 4213 3707 4227
rect 3793 5253 3807 5267
rect 3833 5813 3847 5827
rect 3893 6153 3907 6167
rect 3873 5873 3887 5887
rect 3953 6593 3967 6607
rect 4053 6873 4067 6887
rect 4173 7093 4187 7107
rect 4153 7073 4167 7087
rect 4133 7033 4147 7047
rect 4173 6893 4187 6907
rect 4033 6733 4047 6747
rect 4073 6693 4087 6707
rect 4013 6653 4027 6667
rect 3973 6533 3987 6547
rect 4153 6853 4167 6867
rect 4133 6833 4147 6847
rect 4213 7033 4227 7047
rect 4213 6853 4227 6867
rect 4113 6813 4127 6827
rect 4153 6813 4167 6827
rect 4133 6733 4147 6747
rect 4093 6653 4107 6667
rect 4113 6653 4127 6667
rect 4053 6593 4067 6607
rect 4113 6573 4127 6587
rect 4013 6473 4027 6487
rect 4013 6413 4027 6427
rect 4033 6333 4047 6347
rect 4033 6293 4047 6307
rect 3953 6253 3967 6267
rect 3933 6213 3947 6227
rect 3913 5893 3927 5907
rect 3933 5833 3947 5847
rect 3933 5673 3947 5687
rect 3893 5633 3907 5647
rect 3933 5633 3947 5647
rect 3913 5613 3927 5627
rect 3993 6253 4007 6267
rect 3993 6153 4007 6167
rect 3993 6113 4007 6127
rect 4073 6553 4087 6567
rect 4073 6473 4087 6487
rect 4053 6173 4067 6187
rect 3973 6053 3987 6067
rect 3993 6053 4007 6067
rect 4053 5993 4067 6007
rect 4033 5933 4047 5947
rect 3993 5893 4007 5907
rect 3973 5873 3987 5887
rect 3973 5853 3987 5867
rect 3913 5493 3927 5507
rect 3953 5493 3967 5507
rect 3873 5453 3887 5467
rect 3913 5453 3927 5467
rect 3893 5413 3907 5427
rect 3933 5413 3947 5427
rect 3853 5293 3867 5307
rect 3913 5293 3927 5307
rect 3833 5193 3847 5207
rect 3873 5193 3887 5207
rect 3933 5173 3947 5187
rect 3913 5153 3927 5167
rect 3793 5113 3807 5127
rect 3813 5113 3827 5127
rect 3873 5113 3887 5127
rect 3793 5093 3807 5107
rect 3773 4953 3787 4967
rect 3853 4953 3867 4967
rect 3833 4933 3847 4947
rect 3813 4913 3827 4927
rect 3733 4793 3747 4807
rect 3753 4713 3767 4727
rect 3733 4633 3747 4647
rect 3733 4593 3747 4607
rect 3693 4013 3707 4027
rect 3713 4013 3727 4027
rect 3653 3973 3667 3987
rect 3673 3973 3687 3987
rect 3613 3933 3627 3947
rect 3573 3913 3587 3927
rect 3613 3913 3627 3927
rect 3533 3753 3547 3767
rect 3473 3713 3487 3727
rect 3513 3693 3527 3707
rect 3553 3673 3567 3687
rect 3553 3573 3567 3587
rect 3533 3473 3547 3487
rect 3573 3473 3587 3487
rect 3553 3453 3567 3467
rect 3593 3453 3607 3467
rect 3493 3413 3507 3427
rect 3533 3193 3547 3207
rect 3573 3193 3587 3207
rect 3573 3153 3587 3167
rect 3533 3053 3547 3067
rect 3513 3013 3527 3027
rect 3473 2993 3487 3007
rect 3513 2993 3527 3007
rect 3493 2953 3507 2967
rect 3453 2933 3467 2947
rect 3393 2873 3407 2887
rect 3473 2793 3487 2807
rect 3313 2773 3327 2787
rect 3353 2593 3367 2607
rect 3513 2793 3527 2807
rect 3513 2693 3527 2707
rect 3573 2973 3587 2987
rect 3553 2773 3567 2787
rect 3533 2613 3547 2627
rect 3513 2573 3527 2587
rect 3553 2573 3567 2587
rect 3493 2553 3507 2567
rect 3373 2533 3387 2547
rect 3473 2533 3487 2547
rect 3333 2513 3347 2527
rect 3193 2373 3207 2387
rect 3233 2373 3247 2387
rect 3173 2273 3187 2287
rect 3153 2213 3167 2227
rect 3093 2193 3107 2207
rect 3053 2173 3067 2187
rect 3053 2153 3067 2167
rect 3433 2313 3447 2327
rect 3473 2273 3487 2287
rect 3413 2073 3427 2087
rect 3233 2053 3247 2067
rect 3293 2053 3307 2067
rect 3313 2013 3327 2027
rect 3033 1953 3047 1967
rect 3093 1953 3107 1967
rect 2953 1813 2967 1827
rect 3053 1813 3067 1827
rect 3113 1833 3127 1847
rect 2933 1773 2947 1787
rect 2913 1613 2927 1627
rect 3013 1753 3027 1767
rect 3013 1613 3027 1627
rect 2933 1573 2947 1587
rect 2973 1573 2987 1587
rect 2893 1113 2907 1127
rect 2913 1093 2927 1107
rect 2993 1253 3007 1267
rect 2993 1173 3007 1187
rect 2933 1073 2947 1087
rect 2913 853 2927 867
rect 2893 833 2907 847
rect 2933 833 2947 847
rect 2973 833 2987 847
rect 3073 1713 3087 1727
rect 3133 1773 3147 1787
rect 3033 1533 3047 1547
rect 3053 1453 3067 1467
rect 3033 1093 3047 1107
rect 3033 893 3047 907
rect 3033 853 3047 867
rect 3133 1453 3147 1467
rect 3093 1373 3107 1387
rect 3113 1353 3127 1367
rect 3193 1373 3207 1387
rect 3153 1333 3167 1347
rect 3173 1333 3187 1347
rect 3393 1853 3407 1867
rect 3333 1613 3347 1627
rect 3253 1553 3267 1567
rect 3313 1533 3327 1547
rect 3233 1353 3247 1367
rect 3253 1353 3267 1367
rect 3233 1333 3247 1347
rect 3113 1293 3127 1307
rect 3173 1293 3187 1307
rect 3213 1293 3227 1307
rect 3133 1273 3147 1287
rect 3173 1273 3187 1287
rect 3113 1093 3127 1107
rect 3133 1093 3147 1107
rect 3133 1073 3147 1087
rect 3193 1073 3207 1087
rect 3113 1053 3127 1067
rect 3173 1053 3187 1067
rect 3273 1313 3287 1327
rect 3353 1313 3367 1327
rect 3253 1293 3267 1307
rect 3453 2053 3467 2067
rect 3433 2013 3447 2027
rect 3433 1853 3447 1867
rect 3453 1793 3467 1807
rect 3413 1613 3427 1627
rect 3533 2533 3547 2547
rect 3553 2293 3567 2307
rect 3513 2233 3527 2247
rect 3553 2233 3567 2247
rect 3513 1993 3527 2007
rect 3513 1793 3527 1807
rect 3493 1733 3507 1747
rect 3493 1693 3507 1707
rect 3393 1273 3407 1287
rect 3373 1253 3387 1267
rect 3473 1573 3487 1587
rect 3473 1273 3487 1287
rect 3353 1153 3367 1167
rect 3233 1053 3247 1067
rect 3193 1013 3207 1027
rect 3313 1093 3327 1107
rect 3293 1073 3307 1087
rect 3313 1053 3327 1067
rect 3253 993 3267 1007
rect 3133 833 3147 847
rect 3053 813 3067 827
rect 3333 833 3347 847
rect 3173 813 3187 827
rect 3253 813 3267 827
rect 3133 793 3147 807
rect 3153 793 3167 807
rect 3033 773 3047 787
rect 3013 713 3027 727
rect 3013 673 3027 687
rect 2993 653 3007 667
rect 2933 633 2947 647
rect 2873 613 2887 627
rect 2973 613 2987 627
rect 2993 593 3007 607
rect 2953 573 2967 587
rect 2953 413 2967 427
rect 2913 393 2927 407
rect 2933 393 2947 407
rect 2833 233 2847 247
rect 2853 233 2867 247
rect 2893 233 2907 247
rect 2733 173 2747 187
rect 2713 133 2727 147
rect 2933 353 2947 367
rect 2993 373 3007 387
rect 3233 793 3247 807
rect 3173 673 3187 687
rect 3193 493 3207 507
rect 3013 313 3027 327
rect 2973 273 2987 287
rect 3153 413 3167 427
rect 3193 373 3207 387
rect 3233 353 3247 367
rect 3173 313 3187 327
rect 3213 313 3227 327
rect 3133 193 3147 207
rect 3173 193 3187 207
rect 2813 13 2827 27
rect 2893 13 2907 27
rect 3153 113 3167 127
rect 3373 813 3387 827
rect 3373 793 3387 807
rect 3433 1253 3447 1267
rect 3473 1173 3487 1187
rect 3493 1093 3507 1107
rect 3413 1073 3427 1087
rect 3353 573 3367 587
rect 3393 373 3407 387
rect 3373 353 3387 367
rect 3493 893 3507 907
rect 3453 873 3467 887
rect 3433 593 3447 607
rect 3433 353 3447 367
rect 3413 333 3427 347
rect 3313 153 3327 167
rect 3433 173 3447 187
rect 3313 133 3327 147
rect 3353 133 3367 147
rect 3293 113 3307 127
rect 3353 113 3367 127
rect 3333 93 3347 107
rect 3553 1173 3567 1187
rect 3593 2773 3607 2787
rect 3593 2693 3607 2707
rect 3593 2273 3607 2287
rect 3593 2073 3607 2087
rect 3753 4473 3767 4487
rect 3773 4473 3787 4487
rect 3733 3733 3747 3747
rect 3653 3713 3667 3727
rect 3633 3253 3647 3267
rect 3833 4893 3847 4907
rect 3853 4653 3867 4667
rect 3833 4593 3847 4607
rect 3813 4493 3827 4507
rect 3833 4473 3847 4487
rect 3793 4433 3807 4447
rect 3773 4193 3787 4207
rect 3893 4953 3907 4967
rect 3953 5153 3967 5167
rect 4013 5813 4027 5827
rect 3993 5773 4007 5787
rect 4013 5733 4027 5747
rect 4013 5593 4027 5607
rect 3993 5173 4007 5187
rect 3973 4953 3987 4967
rect 3993 4933 4007 4947
rect 3933 4893 3947 4907
rect 4013 4893 4027 4907
rect 3893 4693 3907 4707
rect 3913 4673 3927 4687
rect 3953 4673 3967 4687
rect 4053 5853 4067 5867
rect 4053 5673 4067 5687
rect 4133 6533 4147 6547
rect 4113 6453 4127 6467
rect 4093 6433 4107 6447
rect 4093 6313 4107 6327
rect 4093 6133 4107 6147
rect 4093 6053 4107 6067
rect 4093 5673 4107 5687
rect 4233 6813 4247 6827
rect 4313 7293 4327 7307
rect 4273 7273 4287 7287
rect 4253 6753 4267 6767
rect 4233 6733 4247 6747
rect 4233 6593 4247 6607
rect 4373 7333 4387 7347
rect 4353 7233 4367 7247
rect 4353 7193 4367 7207
rect 4313 7173 4327 7187
rect 4293 7113 4307 7127
rect 4353 7093 4367 7107
rect 4333 7073 4347 7087
rect 4293 7033 4307 7047
rect 4333 6913 4347 6927
rect 4333 6833 4347 6847
rect 4353 6833 4367 6847
rect 4313 6813 4327 6827
rect 4293 6713 4307 6727
rect 4313 6593 4327 6607
rect 4233 6573 4247 6587
rect 4213 6553 4227 6567
rect 4193 6373 4207 6387
rect 4153 6193 4167 6207
rect 4213 6353 4227 6367
rect 4213 6213 4227 6227
rect 4173 6173 4187 6187
rect 4173 6113 4187 6127
rect 4193 6073 4207 6087
rect 4293 6573 4307 6587
rect 4293 6553 4307 6567
rect 4253 6473 4267 6487
rect 4253 6353 4267 6367
rect 4253 6113 4267 6127
rect 4153 6053 4167 6067
rect 4233 6053 4247 6067
rect 4313 6373 4327 6387
rect 4313 6313 4327 6327
rect 4313 6133 4327 6147
rect 4293 6113 4307 6127
rect 4173 5953 4187 5967
rect 4253 5953 4267 5967
rect 4153 5913 4167 5927
rect 4133 5653 4147 5667
rect 4073 5633 4087 5647
rect 4113 5633 4127 5647
rect 4053 5573 4067 5587
rect 4233 5913 4247 5927
rect 4213 5793 4227 5807
rect 4273 5873 4287 5887
rect 4233 5753 4247 5767
rect 4193 5673 4207 5687
rect 4153 5553 4167 5567
rect 4073 5453 4087 5467
rect 4133 5393 4147 5407
rect 4093 5273 4107 5287
rect 4113 5273 4127 5287
rect 4073 5173 4087 5187
rect 4053 5093 4067 5107
rect 4053 4993 4067 5007
rect 4033 4613 4047 4627
rect 3933 4493 3947 4507
rect 3993 4493 4007 4507
rect 3933 4453 3947 4467
rect 3973 4433 3987 4447
rect 3873 4373 3887 4387
rect 3793 4173 3807 4187
rect 4033 4313 4047 4327
rect 3993 4193 4007 4207
rect 4253 5593 4267 5607
rect 4313 6093 4327 6107
rect 4573 7673 4587 7687
rect 4493 7593 4507 7607
rect 4453 7553 4467 7567
rect 4533 7573 4547 7587
rect 4413 7513 4427 7527
rect 4433 7513 4447 7527
rect 4473 7513 4487 7527
rect 4393 7293 4407 7307
rect 4493 7413 4507 7427
rect 4453 7353 4467 7367
rect 4593 7573 4607 7587
rect 4633 7513 4647 7527
rect 4633 7453 4647 7467
rect 4653 7453 4667 7467
rect 4733 7913 4747 7927
rect 4953 8073 4967 8087
rect 4833 8033 4847 8047
rect 4853 8033 4867 8047
rect 4933 8033 4947 8047
rect 4753 7853 4767 7867
rect 4753 7693 4767 7707
rect 4813 7833 4827 7847
rect 4793 7773 4807 7787
rect 4813 7773 4827 7787
rect 4773 7613 4787 7627
rect 4753 7533 4767 7547
rect 4873 7913 4887 7927
rect 4853 7893 4867 7907
rect 4833 7673 4847 7687
rect 4813 7573 4827 7587
rect 4953 7853 4967 7867
rect 4913 7833 4927 7847
rect 4893 7793 4907 7807
rect 4913 7793 4927 7807
rect 4893 7773 4907 7787
rect 4633 7353 4647 7367
rect 4433 7253 4447 7267
rect 4413 7153 4427 7167
rect 4433 6973 4447 6987
rect 4413 6913 4427 6927
rect 4413 6893 4427 6907
rect 4393 6833 4407 6847
rect 4373 6713 4387 6727
rect 4353 6553 4367 6567
rect 4353 6453 4367 6467
rect 4513 7333 4527 7347
rect 4573 7333 4587 7347
rect 4533 7313 4547 7327
rect 4513 7213 4527 7227
rect 4513 7133 4527 7147
rect 4573 7253 4587 7267
rect 4613 7193 4627 7207
rect 4593 7153 4607 7167
rect 4493 6893 4507 6907
rect 4473 6853 4487 6867
rect 4533 6993 4547 7007
rect 4473 6593 4487 6607
rect 4473 6553 4487 6567
rect 4413 6373 4427 6387
rect 4433 6373 4447 6387
rect 4413 6353 4427 6367
rect 4453 6353 4467 6367
rect 4453 6313 4467 6327
rect 4373 6293 4387 6307
rect 4353 6253 4367 6267
rect 4433 6173 4447 6187
rect 4353 6153 4367 6167
rect 4393 6153 4407 6167
rect 4313 6073 4327 6087
rect 4333 6073 4347 6087
rect 4413 6073 4427 6087
rect 4333 6053 4347 6067
rect 4373 6053 4387 6067
rect 4313 5813 4327 5827
rect 4253 5533 4267 5547
rect 4293 5473 4307 5487
rect 4233 5393 4247 5407
rect 4193 5293 4207 5307
rect 4213 5153 4227 5167
rect 4313 5413 4327 5427
rect 4293 5153 4307 5167
rect 4133 5133 4147 5147
rect 4193 5133 4207 5147
rect 4193 5113 4207 5127
rect 4173 4993 4187 5007
rect 4133 4973 4147 4987
rect 4153 4933 4167 4947
rect 4213 4953 4227 4967
rect 4133 4913 4147 4927
rect 4113 4893 4127 4907
rect 4133 4813 4147 4827
rect 4093 4733 4107 4747
rect 4213 4913 4227 4927
rect 4273 4993 4287 5007
rect 4253 4953 4267 4967
rect 4173 4893 4187 4907
rect 4233 4893 4247 4907
rect 4093 4673 4107 4687
rect 4133 4673 4147 4687
rect 4153 4673 4167 4687
rect 4073 4653 4087 4667
rect 4073 4633 4087 4647
rect 4133 4653 4147 4667
rect 4093 4613 4107 4627
rect 4113 4613 4127 4627
rect 4233 4853 4247 4867
rect 4213 4713 4227 4727
rect 4193 4693 4207 4707
rect 4193 4653 4207 4667
rect 4173 4633 4187 4647
rect 4173 4533 4187 4547
rect 4153 4493 4167 4507
rect 4133 4453 4147 4467
rect 4273 4933 4287 4947
rect 4293 4853 4307 4867
rect 4293 4673 4307 4687
rect 4233 4493 4247 4507
rect 4233 4473 4247 4487
rect 4193 4453 4207 4467
rect 4213 4433 4227 4447
rect 4093 4413 4107 4427
rect 4073 4353 4087 4367
rect 4153 4193 4167 4207
rect 4193 4193 4207 4207
rect 4133 4173 4147 4187
rect 3813 4113 3827 4127
rect 3833 4113 3847 4127
rect 3773 3993 3787 4007
rect 3753 3693 3767 3707
rect 3973 4033 3987 4047
rect 3973 3973 3987 3987
rect 3833 3913 3847 3927
rect 3953 3733 3967 3747
rect 3873 3713 3887 3727
rect 3893 3613 3907 3627
rect 3773 3593 3787 3607
rect 3933 3593 3947 3607
rect 3693 3573 3707 3587
rect 3753 3533 3767 3547
rect 3773 3293 3787 3307
rect 3753 3273 3767 3287
rect 3713 3253 3727 3267
rect 3853 3273 3867 3287
rect 3733 3233 3747 3247
rect 3773 3233 3787 3247
rect 3873 3233 3887 3247
rect 3893 3093 3907 3107
rect 3653 3073 3667 3087
rect 3853 3053 3867 3067
rect 3873 3053 3887 3067
rect 3693 3033 3707 3047
rect 3833 3033 3847 3047
rect 3653 3013 3667 3027
rect 3673 2993 3687 3007
rect 3713 2973 3727 2987
rect 3693 2553 3707 2567
rect 3793 2773 3807 2787
rect 3773 2753 3787 2767
rect 3813 2753 3827 2767
rect 3753 2553 3767 2567
rect 3733 2533 3747 2547
rect 3773 2533 3787 2547
rect 3713 2513 3727 2527
rect 3813 2333 3827 2347
rect 3733 2313 3747 2327
rect 3773 2313 3787 2327
rect 3633 2213 3647 2227
rect 3633 2193 3647 2207
rect 3633 2093 3647 2107
rect 3653 1813 3667 1827
rect 3713 1813 3727 1827
rect 3613 1613 3627 1627
rect 3673 1773 3687 1787
rect 3713 1773 3727 1787
rect 3693 1633 3707 1647
rect 3633 1593 3647 1607
rect 3653 1553 3667 1567
rect 3693 1593 3707 1607
rect 3753 2253 3767 2267
rect 3793 2213 3807 2227
rect 3753 2033 3767 2047
rect 3753 1773 3767 1787
rect 3753 1653 3767 1667
rect 3733 1373 3747 1387
rect 3593 1313 3607 1327
rect 3513 873 3527 887
rect 3573 873 3587 887
rect 3513 853 3527 867
rect 3553 853 3567 867
rect 3493 833 3507 847
rect 3533 833 3547 847
rect 3573 833 3587 847
rect 3693 1313 3707 1327
rect 3773 1313 3787 1327
rect 3713 1293 3727 1307
rect 3873 2893 3887 2907
rect 3873 2773 3887 2787
rect 3933 3233 3947 3247
rect 3933 3193 3947 3207
rect 3973 3213 3987 3227
rect 3953 3173 3967 3187
rect 4053 4153 4067 4167
rect 4133 3953 4147 3967
rect 4173 4013 4187 4027
rect 4153 3873 4167 3887
rect 4113 3733 4127 3747
rect 4013 3413 4027 3427
rect 4073 3713 4087 3727
rect 4053 3653 4067 3667
rect 4093 3513 4107 3527
rect 4033 3293 4047 3307
rect 4093 3273 4107 3287
rect 4013 3213 4027 3227
rect 4053 3213 4067 3227
rect 4093 3213 4107 3227
rect 3993 3133 4007 3147
rect 3973 2993 3987 3007
rect 4033 3053 4047 3067
rect 4093 3033 4107 3047
rect 4073 3013 4087 3027
rect 4093 2993 4107 3007
rect 4013 2953 4027 2967
rect 4033 2753 4047 2767
rect 3993 2733 4007 2747
rect 3933 2673 3947 2687
rect 4193 3953 4207 3967
rect 4253 4433 4267 4447
rect 4253 4413 4267 4427
rect 4233 4333 4247 4347
rect 4433 6013 4447 6027
rect 4373 5893 4387 5907
rect 4413 5893 4427 5907
rect 4453 5893 4467 5907
rect 4353 5833 4367 5847
rect 4353 5753 4367 5767
rect 4473 5713 4487 5727
rect 4433 5673 4447 5687
rect 4473 5653 4487 5667
rect 4453 5633 4467 5647
rect 4373 5593 4387 5607
rect 4413 5453 4427 5467
rect 4453 5433 4467 5447
rect 4513 6553 4527 6567
rect 4593 6853 4607 6867
rect 4673 7353 4687 7367
rect 4713 7353 4727 7367
rect 4793 7473 4807 7487
rect 4773 7353 4787 7367
rect 4733 7333 4747 7347
rect 4693 7313 4707 7327
rect 4713 7273 4727 7287
rect 4673 7093 4687 7107
rect 4653 7053 4667 7067
rect 4633 6873 4647 6887
rect 4633 6853 4647 6867
rect 4613 6833 4627 6847
rect 4553 6753 4567 6767
rect 4573 6733 4587 6747
rect 4553 6633 4567 6647
rect 4613 6593 4627 6607
rect 4573 6473 4587 6487
rect 4593 6473 4607 6487
rect 4533 6413 4547 6427
rect 4573 6413 4587 6427
rect 4593 6413 4607 6427
rect 4773 7153 4787 7167
rect 4793 7113 4807 7127
rect 4793 7093 4807 7107
rect 4773 7073 4787 7087
rect 4693 7053 4707 7067
rect 4753 7053 4767 7067
rect 4733 7033 4747 7047
rect 4713 7013 4727 7027
rect 4693 6873 4707 6887
rect 4753 6993 4767 7007
rect 4873 7513 4887 7527
rect 4833 7033 4847 7047
rect 4813 7013 4827 7027
rect 4793 6913 4807 6927
rect 4813 6913 4827 6927
rect 4753 6893 4767 6907
rect 4773 6893 4787 6907
rect 4733 6873 4747 6887
rect 4773 6873 4787 6887
rect 4933 7673 4947 7687
rect 4993 8093 5007 8107
rect 4973 7793 4987 7807
rect 4953 7593 4967 7607
rect 5113 8533 5127 8547
rect 5093 8513 5107 8527
rect 5093 8313 5107 8327
rect 5113 8233 5127 8247
rect 5093 8213 5107 8227
rect 5073 8073 5087 8087
rect 5233 8993 5247 9007
rect 5213 8913 5227 8927
rect 5233 8873 5247 8887
rect 5273 8913 5287 8927
rect 5253 8793 5267 8807
rect 5173 8693 5187 8707
rect 5253 8553 5267 8567
rect 5153 8533 5167 8547
rect 5193 8513 5207 8527
rect 5233 8513 5247 8527
rect 5213 8493 5227 8507
rect 5173 8433 5187 8447
rect 5153 8413 5167 8427
rect 5133 8193 5147 8207
rect 5173 8393 5187 8407
rect 5153 8093 5167 8107
rect 5053 8013 5067 8027
rect 5013 7913 5027 7927
rect 5073 7853 5087 7867
rect 5153 7853 5167 7867
rect 5013 7833 5027 7847
rect 5033 7833 5047 7847
rect 5013 7793 5027 7807
rect 4993 7553 5007 7567
rect 5013 7513 5027 7527
rect 4933 7473 4947 7487
rect 4993 7433 5007 7447
rect 4913 7393 4927 7407
rect 4953 7353 4967 7367
rect 5113 7833 5127 7847
rect 5133 7813 5147 7827
rect 5073 7773 5087 7787
rect 5053 7593 5067 7607
rect 5033 7373 5047 7387
rect 4893 7333 4907 7347
rect 4973 7333 4987 7347
rect 4873 6913 4887 6927
rect 4753 6853 4767 6867
rect 4793 6853 4807 6867
rect 4853 6873 4867 6887
rect 4713 6833 4727 6847
rect 4753 6833 4767 6847
rect 4793 6833 4807 6847
rect 4833 6833 4847 6847
rect 4673 6813 4687 6827
rect 4673 6733 4687 6747
rect 4673 6653 4687 6667
rect 4713 6613 4727 6627
rect 4673 6593 4687 6607
rect 4693 6573 4707 6587
rect 4733 6553 4747 6567
rect 4653 6533 4667 6547
rect 4553 6393 4567 6407
rect 4733 6513 4747 6527
rect 4673 6473 4687 6487
rect 4733 6473 4747 6487
rect 4653 6393 4667 6407
rect 4533 6373 4547 6387
rect 4613 6373 4627 6387
rect 4653 6373 4667 6387
rect 4573 6213 4587 6227
rect 4533 6193 4547 6207
rect 4533 6153 4547 6167
rect 4613 6113 4627 6127
rect 4533 6093 4547 6107
rect 4553 6073 4567 6087
rect 4513 6013 4527 6027
rect 4553 6013 4567 6027
rect 4573 6013 4587 6027
rect 4533 5953 4547 5967
rect 4513 5833 4527 5847
rect 4433 5413 4447 5427
rect 4493 5413 4507 5427
rect 4493 5393 4507 5407
rect 4453 5153 4467 5167
rect 4433 5133 4447 5147
rect 4513 5173 4527 5187
rect 4493 5133 4507 5147
rect 4413 5073 4427 5087
rect 4453 5073 4467 5087
rect 4393 5033 4407 5047
rect 4573 5933 4587 5947
rect 4613 5913 4627 5927
rect 4593 5873 4607 5887
rect 4713 6393 4727 6407
rect 4733 6393 4747 6407
rect 4773 6713 4787 6727
rect 4813 6793 4827 6807
rect 4813 6613 4827 6627
rect 4793 6593 4807 6607
rect 4773 6573 4787 6587
rect 4793 6553 4807 6567
rect 4793 6413 4807 6427
rect 4773 6393 4787 6407
rect 4933 7313 4947 7327
rect 4953 7213 4967 7227
rect 4933 7173 4947 7187
rect 5053 7213 5067 7227
rect 4973 7173 4987 7187
rect 4933 7073 4947 7087
rect 4953 7073 4967 7087
rect 4913 7053 4927 7067
rect 4953 7013 4967 7027
rect 4993 6913 5007 6927
rect 5033 6913 5047 6927
rect 4973 6873 4987 6887
rect 5013 6873 5027 6887
rect 4953 6853 4967 6867
rect 4893 6793 4907 6807
rect 4873 6693 4887 6707
rect 4933 6773 4947 6787
rect 4953 6773 4967 6787
rect 4893 6633 4907 6647
rect 4933 6573 4947 6587
rect 4833 6513 4847 6527
rect 4753 6373 4767 6387
rect 4733 6313 4747 6327
rect 4713 6293 4727 6307
rect 4673 6213 4687 6227
rect 4693 6213 4707 6227
rect 4653 5753 4667 5767
rect 4713 6153 4727 6167
rect 4773 6153 4787 6167
rect 4813 6153 4827 6167
rect 4813 6113 4827 6127
rect 4733 6093 4747 6107
rect 4753 6093 4767 6107
rect 4773 5993 4787 6007
rect 4913 6553 4927 6567
rect 4893 6533 4907 6547
rect 4993 6693 5007 6707
rect 4973 6633 4987 6647
rect 4973 6593 4987 6607
rect 4993 6593 5007 6607
rect 4993 6533 5007 6547
rect 4993 6473 5007 6487
rect 4933 6413 4947 6427
rect 4973 6413 4987 6427
rect 4893 6373 4907 6387
rect 4873 6193 4887 6207
rect 4873 6113 4887 6127
rect 4793 5933 4807 5947
rect 4853 5953 4867 5967
rect 4833 5933 4847 5947
rect 4813 5913 4827 5927
rect 4753 5893 4767 5907
rect 4793 5893 4807 5907
rect 4713 5793 4727 5807
rect 4693 5673 4707 5687
rect 4613 5633 4627 5647
rect 4593 5613 4607 5627
rect 4673 5593 4687 5607
rect 4633 5553 4647 5567
rect 4693 5513 4707 5527
rect 4613 5493 4627 5507
rect 4553 5453 4567 5467
rect 4653 5433 4667 5447
rect 4633 5413 4647 5427
rect 4673 5413 4687 5427
rect 4693 5313 4707 5327
rect 4673 5253 4687 5267
rect 4613 5173 4627 5187
rect 4573 5153 4587 5167
rect 4653 5153 4667 5167
rect 4533 5113 4547 5127
rect 4533 5053 4547 5067
rect 4553 5053 4567 5067
rect 4533 5033 4547 5047
rect 4513 4993 4527 5007
rect 4413 4973 4427 4987
rect 4553 5013 4567 5027
rect 4593 5133 4607 5147
rect 4693 5133 4707 5147
rect 4713 5133 4727 5147
rect 4673 5073 4687 5087
rect 4693 5013 4707 5027
rect 4573 4993 4587 5007
rect 4573 4973 4587 4987
rect 4373 4953 4387 4967
rect 4393 4933 4407 4947
rect 4553 4933 4567 4947
rect 4333 4893 4347 4907
rect 4393 4893 4407 4907
rect 4333 4733 4347 4747
rect 4333 4573 4347 4587
rect 4293 4473 4307 4487
rect 4313 4473 4327 4487
rect 4353 4193 4367 4207
rect 4433 4753 4447 4767
rect 4473 4693 4487 4707
rect 4453 4673 4467 4687
rect 4413 4613 4427 4627
rect 4413 4453 4427 4467
rect 4333 4153 4347 4167
rect 4393 4153 4407 4167
rect 4273 4133 4287 4147
rect 4333 4133 4347 4147
rect 4253 3733 4267 3747
rect 4233 3713 4247 3727
rect 4493 4373 4507 4387
rect 4553 4253 4567 4267
rect 4633 4853 4647 4867
rect 4773 5653 4787 5667
rect 4753 5633 4767 5647
rect 4753 5413 4767 5427
rect 4753 5393 4767 5407
rect 4813 5653 4827 5667
rect 4793 5633 4807 5647
rect 4953 6393 4967 6407
rect 4993 6393 5007 6407
rect 4973 6313 4987 6327
rect 5053 6873 5067 6887
rect 5073 6873 5087 6887
rect 5053 6833 5067 6847
rect 5153 7673 5167 7687
rect 5133 7593 5147 7607
rect 5233 8293 5247 8307
rect 5193 8113 5207 8127
rect 5273 8093 5287 8107
rect 5233 8053 5247 8067
rect 5273 8033 5287 8047
rect 5253 7993 5267 8007
rect 5273 7913 5287 7927
rect 5473 9773 5487 9787
rect 5393 9473 5407 9487
rect 5473 9473 5487 9487
rect 5353 9313 5367 9327
rect 5333 9273 5347 9287
rect 5333 9193 5347 9207
rect 5333 9153 5347 9167
rect 5313 8773 5327 8787
rect 5313 8313 5327 8327
rect 6173 10693 6187 10707
rect 6013 10473 6027 10487
rect 5913 10433 5927 10447
rect 5933 10433 5947 10447
rect 5973 10433 5987 10447
rect 5933 10413 5947 10427
rect 5913 10393 5927 10407
rect 5853 10373 5867 10387
rect 5953 10393 5967 10407
rect 5853 10273 5867 10287
rect 5833 10193 5847 10207
rect 5753 10133 5767 10147
rect 5733 9953 5747 9967
rect 5673 9873 5687 9887
rect 5633 9533 5647 9547
rect 5433 9453 5447 9467
rect 5493 9453 5507 9467
rect 5613 9453 5627 9467
rect 5413 9433 5427 9447
rect 5473 9293 5487 9307
rect 5433 9273 5447 9287
rect 5513 9273 5527 9287
rect 5533 9273 5547 9287
rect 5453 9253 5467 9267
rect 5493 9253 5507 9267
rect 5453 9233 5467 9247
rect 5513 9193 5527 9207
rect 5433 9173 5447 9187
rect 5453 9173 5467 9187
rect 5453 9133 5467 9147
rect 5433 9033 5447 9047
rect 5453 9013 5467 9027
rect 5613 9173 5627 9187
rect 5573 9013 5587 9027
rect 5373 8973 5387 8987
rect 5413 8973 5427 8987
rect 5353 8893 5367 8907
rect 5533 8893 5547 8907
rect 5353 8793 5367 8807
rect 5393 8793 5407 8807
rect 5473 8793 5487 8807
rect 5373 8773 5387 8787
rect 5413 8773 5427 8787
rect 5513 8773 5527 8787
rect 5393 8533 5407 8547
rect 5413 8513 5427 8527
rect 5473 8533 5487 8547
rect 5513 8513 5527 8527
rect 5453 8433 5467 8447
rect 5493 8413 5507 8427
rect 5593 8953 5607 8967
rect 5573 8873 5587 8887
rect 5573 8773 5587 8787
rect 5553 8553 5567 8567
rect 5573 8513 5587 8527
rect 5533 8373 5547 8387
rect 5513 8293 5527 8307
rect 5353 8193 5367 8207
rect 5333 8113 5347 8127
rect 5313 7953 5327 7967
rect 5293 7893 5307 7907
rect 5573 8193 5587 8207
rect 5513 8133 5527 8147
rect 5393 8093 5407 8107
rect 5413 8093 5427 8107
rect 5373 8053 5387 8067
rect 5373 7973 5387 7987
rect 5353 7913 5367 7927
rect 5373 7893 5387 7907
rect 5373 7833 5387 7847
rect 5293 7813 5307 7827
rect 5273 7793 5287 7807
rect 5213 7753 5227 7767
rect 5173 7593 5187 7607
rect 5153 7573 5167 7587
rect 5193 7573 5207 7587
rect 5153 7533 5167 7547
rect 5173 7533 5187 7547
rect 5133 7513 5147 7527
rect 5113 7473 5127 7487
rect 5153 7473 5167 7487
rect 5233 7713 5247 7727
rect 5153 7453 5167 7467
rect 5213 7453 5227 7467
rect 5133 7353 5147 7367
rect 5193 7353 5207 7367
rect 5213 7353 5227 7367
rect 5113 7333 5127 7347
rect 5153 7233 5167 7247
rect 5193 7133 5207 7147
rect 5133 7053 5147 7067
rect 5113 7033 5127 7047
rect 5193 7013 5207 7027
rect 5173 6913 5187 6927
rect 5213 6913 5227 6927
rect 5133 6893 5147 6907
rect 5173 6893 5187 6907
rect 5433 8053 5447 8067
rect 5453 8013 5467 8027
rect 5493 8033 5507 8047
rect 5473 7953 5487 7967
rect 5573 8073 5587 8087
rect 5613 8293 5627 8307
rect 5613 8233 5627 8247
rect 5613 8073 5627 8087
rect 5713 9493 5727 9507
rect 5673 9453 5687 9467
rect 5653 9393 5667 9407
rect 5673 9253 5687 9267
rect 5693 9213 5707 9227
rect 5653 9173 5667 9187
rect 5853 9913 5867 9927
rect 5813 9813 5827 9827
rect 5813 9793 5827 9807
rect 5933 10213 5947 10227
rect 5993 10193 6007 10207
rect 5933 10173 5947 10187
rect 5933 10093 5947 10107
rect 6293 11393 6307 11407
rect 6293 11373 6307 11387
rect 6413 11673 6427 11687
rect 6493 11653 6507 11667
rect 6713 11673 6727 11687
rect 6653 11653 6667 11667
rect 6453 11633 6467 11647
rect 6553 11633 6567 11647
rect 6633 11633 6647 11647
rect 6693 11633 6707 11647
rect 6573 11613 6587 11627
rect 6673 11613 6687 11627
rect 6553 11533 6567 11547
rect 6453 11373 6467 11387
rect 6433 11233 6447 11247
rect 6333 11193 6347 11207
rect 6313 11173 6327 11187
rect 6353 11173 6367 11187
rect 6473 11333 6487 11347
rect 6353 11133 6367 11147
rect 6413 11133 6427 11147
rect 6253 11013 6267 11027
rect 6233 10913 6247 10927
rect 6213 10893 6227 10907
rect 6253 10833 6267 10847
rect 6293 10913 6307 10927
rect 6373 10913 6387 10927
rect 6353 10813 6367 10827
rect 6273 10733 6287 10747
rect 6133 10433 6147 10447
rect 6113 10313 6127 10327
rect 6193 10433 6207 10447
rect 6393 10733 6407 10747
rect 6373 10673 6387 10687
rect 6413 10653 6427 10667
rect 6373 10453 6387 10467
rect 6333 10433 6347 10447
rect 6293 10413 6307 10427
rect 6173 10393 6187 10407
rect 6313 10353 6327 10367
rect 6153 10293 6167 10307
rect 6313 10293 6327 10307
rect 6133 10273 6147 10287
rect 6153 10253 6167 10267
rect 5913 9893 5927 9907
rect 5973 9913 5987 9927
rect 5973 9893 5987 9907
rect 5953 9853 5967 9867
rect 5953 9813 5967 9827
rect 5873 9793 5887 9807
rect 5773 9593 5787 9607
rect 5733 9273 5747 9287
rect 5793 9493 5807 9507
rect 5833 9493 5847 9507
rect 5813 9473 5827 9487
rect 5813 9273 5827 9287
rect 5893 9773 5907 9787
rect 5913 9733 5927 9747
rect 5893 9553 5907 9567
rect 5873 9493 5887 9507
rect 5893 9473 5907 9487
rect 5913 9473 5927 9487
rect 5873 9333 5887 9347
rect 5773 9213 5787 9227
rect 5773 8993 5787 9007
rect 5793 8973 5807 8987
rect 5753 8953 5767 8967
rect 5713 8913 5727 8927
rect 5773 8913 5787 8927
rect 5753 8793 5767 8807
rect 5733 8773 5747 8787
rect 5813 8813 5827 8827
rect 5813 8793 5827 8807
rect 5713 8713 5727 8727
rect 5473 7893 5487 7907
rect 5513 7893 5527 7907
rect 5413 7793 5427 7807
rect 5433 7793 5447 7807
rect 5393 7573 5407 7587
rect 5253 7533 5267 7547
rect 5333 7533 5347 7547
rect 5353 7373 5367 7387
rect 5393 7373 5407 7387
rect 5273 7353 5287 7367
rect 5273 7293 5287 7307
rect 5273 7133 5287 7147
rect 5273 7093 5287 7107
rect 5253 7053 5267 7067
rect 5393 7353 5407 7367
rect 5373 7333 5387 7347
rect 5413 7333 5427 7347
rect 5333 7313 5347 7327
rect 5353 7273 5367 7287
rect 5413 7213 5427 7227
rect 5393 7173 5407 7187
rect 5313 7053 5327 7067
rect 5333 7053 5347 7067
rect 5373 7053 5387 7067
rect 5293 7033 5307 7047
rect 5333 7033 5347 7047
rect 5393 7033 5407 7047
rect 5253 6893 5267 6907
rect 5273 6893 5287 6907
rect 5313 6893 5327 6907
rect 5113 6853 5127 6867
rect 5073 6813 5087 6827
rect 5093 6813 5107 6827
rect 5133 6833 5147 6847
rect 5193 6853 5207 6867
rect 5113 6773 5127 6787
rect 5053 6713 5067 6727
rect 5113 6693 5127 6707
rect 5213 6813 5227 6827
rect 5173 6793 5187 6807
rect 5193 6713 5207 6727
rect 5173 6633 5187 6647
rect 5153 6613 5167 6627
rect 5093 6553 5107 6567
rect 5113 6553 5127 6567
rect 5033 6473 5047 6487
rect 5093 6473 5107 6487
rect 5073 6353 5087 6367
rect 4933 6253 4947 6267
rect 4933 6113 4947 6127
rect 5013 6253 5027 6267
rect 5033 6253 5047 6267
rect 5013 6113 5027 6127
rect 4893 6093 4907 6107
rect 4993 6093 5007 6107
rect 4953 6013 4967 6027
rect 4913 5973 4927 5987
rect 4913 5953 4927 5967
rect 4893 5913 4907 5927
rect 4873 5893 4887 5907
rect 4833 5633 4847 5647
rect 4793 5593 4807 5607
rect 4793 5533 4807 5547
rect 4793 5453 4807 5467
rect 4873 5453 4887 5467
rect 4773 5373 4787 5387
rect 4753 5193 4767 5207
rect 4733 5013 4747 5027
rect 4853 5433 4867 5447
rect 4793 5153 4807 5167
rect 4773 5133 4787 5147
rect 4813 5133 4827 5147
rect 4793 5113 4807 5127
rect 4693 4833 4707 4847
rect 4673 4753 4687 4767
rect 4653 4633 4667 4647
rect 4633 4493 4647 4507
rect 4633 4233 4647 4247
rect 4573 4173 4587 4187
rect 4613 4193 4627 4207
rect 4633 4193 4647 4207
rect 4533 4113 4547 4127
rect 4413 4093 4427 4107
rect 4573 4093 4587 4107
rect 4353 4013 4367 4027
rect 4353 3973 4367 3987
rect 4533 3973 4547 3987
rect 4393 3813 4407 3827
rect 4333 3613 4347 3627
rect 4373 3593 4387 3607
rect 4553 3653 4567 3667
rect 4513 3613 4527 3627
rect 4413 3593 4427 3607
rect 4153 3513 4167 3527
rect 4173 3493 4187 3507
rect 4373 3493 4387 3507
rect 4233 3253 4247 3267
rect 4613 3813 4627 3827
rect 4573 3533 4587 3547
rect 4553 3253 4567 3267
rect 4133 3233 4147 3247
rect 4213 3233 4227 3247
rect 4413 3233 4427 3247
rect 4393 3173 4407 3187
rect 4373 3133 4387 3147
rect 4173 3053 4187 3067
rect 4233 3053 4247 3067
rect 4293 2953 4307 2967
rect 4253 2893 4267 2907
rect 4173 2793 4187 2807
rect 4253 2773 4267 2787
rect 4293 2773 4307 2787
rect 4233 2753 4247 2767
rect 4273 2753 4287 2767
rect 4173 2733 4187 2747
rect 4193 2733 4207 2747
rect 4133 2713 4147 2727
rect 3933 2653 3947 2667
rect 4113 2653 4127 2667
rect 3913 2593 3927 2607
rect 3853 2573 3867 2587
rect 3893 2573 3907 2587
rect 3913 2533 3927 2547
rect 3913 2293 3927 2307
rect 3893 2273 3907 2287
rect 3853 2253 3867 2267
rect 3873 2233 3887 2247
rect 3913 2233 3927 2247
rect 3873 2173 3887 2187
rect 3873 2113 3887 2127
rect 3833 2093 3847 2107
rect 3833 2073 3847 2087
rect 3813 2053 3827 2067
rect 3893 1773 3907 1787
rect 3893 1633 3907 1647
rect 3873 1613 3887 1627
rect 3853 1573 3867 1587
rect 3833 1413 3847 1427
rect 3793 1293 3807 1307
rect 3873 1253 3887 1267
rect 3673 1153 3687 1167
rect 3653 1133 3667 1147
rect 3713 1133 3727 1147
rect 3633 1093 3647 1107
rect 3673 1093 3687 1107
rect 3613 1073 3627 1087
rect 3653 1073 3667 1087
rect 3613 1013 3627 1027
rect 3613 853 3627 867
rect 3593 773 3607 787
rect 3493 653 3507 667
rect 3513 633 3527 647
rect 3473 573 3487 587
rect 3553 513 3567 527
rect 3753 1113 3767 1127
rect 3673 433 3687 447
rect 3533 373 3547 387
rect 3473 293 3487 307
rect 3573 353 3587 367
rect 3473 173 3487 187
rect 3533 173 3547 187
rect 3493 133 3507 147
rect 3593 133 3607 147
rect 3533 113 3547 127
rect 3453 13 3467 27
rect 3493 13 3507 27
rect 3653 133 3667 147
rect 3813 1093 3827 1107
rect 3953 2593 3967 2607
rect 4313 2693 4327 2707
rect 4393 3053 4407 3067
rect 4433 3033 4447 3047
rect 4493 3033 4507 3047
rect 4413 2973 4427 2987
rect 4493 2993 4507 3007
rect 4473 2953 4487 2967
rect 4433 2753 4447 2767
rect 4553 3053 4567 3067
rect 4513 2753 4527 2767
rect 4413 2733 4427 2747
rect 4493 2733 4507 2747
rect 4453 2713 4467 2727
rect 4413 2693 4427 2707
rect 4373 2573 4387 2587
rect 4313 2553 4327 2567
rect 3973 2493 3987 2507
rect 4393 2533 4407 2547
rect 4033 2493 4047 2507
rect 3953 2273 3967 2287
rect 3953 2193 3967 2207
rect 3933 1613 3947 1627
rect 3913 1133 3927 1147
rect 3913 1113 3927 1127
rect 3813 893 3827 907
rect 3893 1073 3907 1087
rect 3953 1133 3967 1147
rect 3933 1033 3947 1047
rect 3873 873 3887 887
rect 3773 813 3787 827
rect 3853 813 3867 827
rect 3713 653 3727 667
rect 3733 653 3747 667
rect 3893 853 3907 867
rect 3873 673 3887 687
rect 3753 633 3767 647
rect 3913 813 3927 827
rect 3893 653 3907 667
rect 4093 2293 4107 2307
rect 4253 2273 4267 2287
rect 4073 2253 4087 2267
rect 4113 2253 4127 2267
rect 4233 2253 4247 2267
rect 4553 2733 4567 2747
rect 4513 2533 4527 2547
rect 4493 2513 4507 2527
rect 4453 2273 4467 2287
rect 4293 2233 4307 2247
rect 4473 2233 4487 2247
rect 4273 2213 4287 2227
rect 4353 2213 4367 2227
rect 4393 2093 4407 2107
rect 4553 2513 4567 2527
rect 4533 2273 4547 2287
rect 4513 2133 4527 2147
rect 4533 2113 4547 2127
rect 4393 2073 4407 2087
rect 4473 2073 4487 2087
rect 4493 2073 4507 2087
rect 4093 2053 4107 2067
rect 4233 2053 4247 2067
rect 4293 2053 4307 2067
rect 4053 2033 4067 2047
rect 4173 1793 4187 1807
rect 4233 1773 4247 1787
rect 4333 1993 4347 2007
rect 4313 1773 4327 1787
rect 4193 1753 4207 1767
rect 3993 1713 4007 1727
rect 3993 1693 4007 1707
rect 4173 1653 4187 1667
rect 4153 1613 4167 1627
rect 4373 1933 4387 1947
rect 4553 1773 4567 1787
rect 4453 1753 4467 1767
rect 4373 1613 4387 1627
rect 4393 1613 4407 1627
rect 4553 1653 4567 1667
rect 4553 1633 4567 1647
rect 4313 1553 4327 1567
rect 4453 1553 4467 1567
rect 4193 1333 4207 1347
rect 4073 1313 4087 1327
rect 4153 1313 4167 1327
rect 4093 1273 4107 1287
rect 4113 1273 4127 1287
rect 4053 1213 4067 1227
rect 3973 873 3987 887
rect 4013 1093 4027 1107
rect 4273 1333 4287 1347
rect 4253 1313 4267 1327
rect 4453 1393 4467 1407
rect 4453 1373 4467 1387
rect 4533 1353 4547 1367
rect 4213 1153 4227 1167
rect 4273 1153 4287 1167
rect 4193 1133 4207 1147
rect 4153 1113 4167 1127
rect 4013 873 4027 887
rect 3993 853 4007 867
rect 3993 833 4007 847
rect 3973 713 3987 727
rect 3973 653 3987 667
rect 3873 533 3887 547
rect 3953 533 3967 547
rect 3853 453 3867 467
rect 3753 333 3767 347
rect 3833 353 3847 367
rect 3853 333 3867 347
rect 3833 313 3847 327
rect 3793 213 3807 227
rect 3833 213 3847 227
rect 3713 173 3727 187
rect 3773 13 3787 27
rect 3813 13 3827 27
rect 3953 493 3967 507
rect 3913 353 3927 367
rect 3993 393 4007 407
rect 3973 373 3987 387
rect 4033 853 4047 867
rect 4153 853 4167 867
rect 4013 353 4027 367
rect 3893 333 3907 347
rect 3933 333 3947 347
rect 3993 333 4007 347
rect 3973 313 3987 327
rect 3993 293 4007 307
rect 3953 173 3967 187
rect 4013 113 4027 127
rect 4053 793 4067 807
rect 4253 1093 4267 1107
rect 4213 1053 4227 1067
rect 4213 1033 4227 1047
rect 4113 653 4127 667
rect 4093 633 4107 647
rect 4173 633 4187 647
rect 4133 613 4147 627
rect 4073 493 4087 507
rect 4113 453 4127 467
rect 4093 433 4107 447
rect 4193 493 4207 507
rect 4173 393 4187 407
rect 4093 353 4107 367
rect 4133 353 4147 367
rect 4253 873 4267 887
rect 4253 853 4267 867
rect 4253 813 4267 827
rect 4233 713 4247 727
rect 4293 853 4307 867
rect 4333 853 4347 867
rect 4273 653 4287 667
rect 4293 653 4307 667
rect 4253 633 4267 647
rect 4313 633 4327 647
rect 4433 1273 4447 1287
rect 4473 1273 4487 1287
rect 4433 1133 4447 1147
rect 4533 1133 4547 1147
rect 4413 1093 4427 1107
rect 4553 1113 4567 1127
rect 4533 1033 4547 1047
rect 4473 873 4487 887
rect 4513 853 4527 867
rect 4453 673 4467 687
rect 4433 613 4447 627
rect 4433 593 4447 607
rect 4413 413 4427 427
rect 4253 393 4267 407
rect 4273 373 4287 387
rect 4253 353 4267 367
rect 4213 273 4227 287
rect 4333 353 4347 367
rect 4313 313 4327 327
rect 4393 373 4407 387
rect 4393 333 4407 347
rect 4673 4433 4687 4447
rect 4873 5373 4887 5387
rect 4833 4933 4847 4947
rect 4813 4713 4827 4727
rect 4833 4693 4847 4707
rect 4793 4673 4807 4687
rect 4833 4673 4847 4687
rect 4773 4653 4787 4667
rect 4853 4653 4867 4667
rect 4733 4633 4747 4647
rect 4813 4633 4827 4647
rect 4813 4493 4827 4507
rect 4733 4433 4747 4447
rect 4713 4253 4727 4267
rect 4693 4193 4707 4207
rect 4933 5933 4947 5947
rect 4973 5913 4987 5927
rect 5033 6093 5047 6107
rect 5053 6093 5067 6107
rect 5013 6053 5027 6067
rect 5033 6053 5047 6067
rect 5013 6013 5027 6027
rect 4953 5873 4967 5887
rect 5033 5893 5047 5907
rect 4933 5753 4947 5767
rect 5013 5753 5027 5767
rect 4913 5413 4927 5427
rect 4893 5093 4907 5107
rect 4953 5653 4967 5667
rect 5013 5613 5027 5627
rect 5053 5833 5067 5847
rect 5053 5733 5067 5747
rect 5053 5593 5067 5607
rect 5173 6473 5187 6487
rect 5273 6873 5287 6887
rect 5293 6873 5307 6887
rect 5273 6773 5287 6787
rect 5253 6713 5267 6727
rect 5313 6853 5327 6867
rect 5293 6613 5307 6627
rect 5233 6593 5247 6607
rect 5213 6553 5227 6567
rect 5273 6573 5287 6587
rect 5313 6573 5327 6587
rect 5253 6553 5267 6567
rect 5273 6553 5287 6567
rect 5373 6873 5387 6887
rect 5353 6853 5367 6867
rect 5393 6733 5407 6747
rect 5353 6613 5367 6627
rect 5333 6493 5347 6507
rect 5373 6593 5387 6607
rect 5353 6473 5367 6487
rect 5193 6393 5207 6407
rect 5233 6393 5247 6407
rect 5153 6373 5167 6387
rect 5233 6353 5247 6367
rect 5133 6253 5147 6267
rect 5113 6173 5127 6187
rect 5113 6073 5127 6087
rect 5233 6153 5247 6167
rect 5173 6113 5187 6127
rect 5153 6093 5167 6107
rect 5133 6033 5147 6047
rect 5193 6033 5207 6047
rect 5113 6013 5127 6027
rect 5213 6013 5227 6027
rect 5093 5973 5107 5987
rect 5133 5933 5147 5947
rect 5193 5933 5207 5947
rect 5113 5913 5127 5927
rect 5173 5913 5187 5927
rect 5093 5693 5107 5707
rect 5073 5553 5087 5567
rect 5033 5473 5047 5487
rect 5033 5453 5047 5467
rect 5073 5453 5087 5467
rect 4973 5433 4987 5447
rect 5013 5433 5027 5447
rect 5053 5433 5067 5447
rect 4953 5413 4967 5427
rect 4973 5373 4987 5387
rect 4933 5273 4947 5287
rect 4953 5173 4967 5187
rect 4933 5113 4947 5127
rect 4893 4933 4907 4947
rect 4973 4793 4987 4807
rect 4953 4773 4967 4787
rect 4913 4673 4927 4687
rect 4893 4633 4907 4647
rect 4873 4193 4887 4207
rect 4953 4653 4967 4667
rect 5033 5413 5047 5427
rect 5033 5193 5047 5207
rect 5153 5893 5167 5907
rect 5113 5673 5127 5687
rect 5213 5693 5227 5707
rect 5213 5633 5227 5647
rect 5313 6393 5327 6407
rect 5293 6373 5307 6387
rect 5273 6353 5287 6367
rect 5333 6353 5347 6367
rect 5333 6333 5347 6347
rect 5313 6153 5327 6167
rect 5293 6133 5307 6147
rect 5273 6033 5287 6047
rect 5273 5773 5287 5787
rect 5253 5633 5267 5647
rect 5233 5593 5247 5607
rect 5173 5573 5187 5587
rect 5193 5573 5207 5587
rect 5153 5513 5167 5527
rect 5133 5413 5147 5427
rect 5233 5473 5247 5487
rect 5393 6473 5407 6487
rect 5393 6293 5407 6307
rect 5393 6193 5407 6207
rect 5373 6133 5387 6147
rect 5353 6113 5367 6127
rect 5453 7533 5467 7547
rect 5453 7173 5467 7187
rect 5453 7153 5467 7167
rect 5453 7073 5467 7087
rect 5553 7873 5567 7887
rect 5513 7813 5527 7827
rect 5493 7793 5507 7807
rect 5533 7773 5547 7787
rect 5653 8053 5667 8067
rect 5613 8033 5627 8047
rect 5593 8013 5607 8027
rect 5593 7993 5607 8007
rect 5613 7993 5627 8007
rect 5633 7973 5647 7987
rect 5633 7953 5647 7967
rect 5613 7913 5627 7927
rect 5593 7893 5607 7907
rect 5593 7813 5607 7827
rect 5593 7773 5607 7787
rect 5573 7753 5587 7767
rect 5553 7673 5567 7687
rect 5593 7673 5607 7687
rect 5533 7593 5547 7607
rect 5513 7573 5527 7587
rect 5693 7853 5707 7867
rect 5673 7793 5687 7807
rect 5673 7753 5687 7767
rect 5653 7613 5667 7627
rect 5573 7353 5587 7367
rect 5513 7293 5527 7307
rect 5653 7533 5667 7547
rect 5653 7513 5667 7527
rect 5633 7453 5647 7467
rect 5653 7453 5667 7467
rect 5613 7353 5627 7367
rect 5553 7233 5567 7247
rect 5533 7213 5547 7227
rect 5613 7213 5627 7227
rect 5593 7113 5607 7127
rect 5573 7073 5587 7087
rect 5473 7053 5487 7067
rect 5493 7053 5507 7067
rect 5453 6913 5467 6927
rect 5473 6913 5487 6927
rect 5453 6713 5467 6727
rect 5453 6613 5467 6627
rect 5473 6593 5487 6607
rect 5453 6533 5467 6547
rect 5473 6533 5487 6547
rect 5453 6493 5467 6507
rect 5433 6413 5447 6427
rect 5433 6373 5447 6387
rect 5433 6233 5447 6247
rect 5413 6173 5427 6187
rect 5373 6093 5387 6107
rect 5333 6033 5347 6047
rect 5313 6013 5327 6027
rect 5353 6013 5367 6027
rect 5333 5993 5347 6007
rect 5413 5993 5427 6007
rect 5353 5933 5367 5947
rect 5373 5933 5387 5947
rect 5393 5913 5407 5927
rect 5393 5833 5407 5847
rect 5393 5773 5407 5787
rect 5313 5633 5327 5647
rect 5353 5633 5367 5647
rect 5333 5613 5347 5627
rect 5373 5593 5387 5607
rect 5293 5473 5307 5487
rect 5253 5453 5267 5467
rect 5293 5453 5307 5467
rect 5213 5413 5227 5427
rect 5253 5413 5267 5427
rect 5153 5253 5167 5267
rect 5153 5193 5167 5207
rect 5113 5153 5127 5167
rect 5313 5413 5327 5427
rect 5553 7013 5567 7027
rect 5553 6873 5567 6887
rect 5553 6853 5567 6867
rect 5513 6773 5527 6787
rect 5613 7013 5627 7027
rect 5593 6853 5607 6867
rect 5613 6833 5627 6847
rect 5553 6813 5567 6827
rect 5533 6753 5547 6767
rect 5653 7333 5667 7347
rect 5673 7333 5687 7347
rect 5653 7213 5667 7227
rect 5933 9393 5947 9407
rect 5913 9293 5927 9307
rect 6293 9893 6307 9907
rect 6333 10273 6347 10287
rect 6353 10253 6367 10267
rect 6413 10293 6427 10307
rect 6433 10253 6447 10267
rect 6453 10193 6467 10207
rect 6393 10093 6407 10107
rect 6453 9973 6467 9987
rect 6413 9953 6427 9967
rect 6213 9853 6227 9867
rect 6073 9793 6087 9807
rect 6053 9773 6067 9787
rect 6013 9753 6027 9767
rect 5993 9733 6007 9747
rect 6013 9713 6027 9727
rect 6013 9513 6027 9527
rect 6213 9753 6227 9767
rect 6153 9653 6167 9667
rect 6153 9533 6167 9547
rect 6173 9473 6187 9487
rect 6213 9473 6227 9487
rect 6153 9453 6167 9467
rect 6033 9413 6047 9427
rect 6013 9373 6027 9387
rect 6073 9313 6087 9327
rect 6093 9293 6107 9307
rect 6133 9173 6147 9187
rect 6113 9133 6127 9147
rect 6013 9053 6027 9067
rect 5993 9013 6007 9027
rect 5973 8993 5987 9007
rect 5933 8933 5947 8947
rect 5953 8933 5967 8947
rect 5993 8953 6007 8967
rect 5973 8913 5987 8927
rect 5893 8793 5907 8807
rect 5953 8793 5967 8807
rect 6073 8973 6087 8987
rect 6053 8873 6067 8887
rect 6033 8833 6047 8847
rect 6033 8813 6047 8827
rect 5833 8733 5847 8747
rect 5793 8693 5807 8707
rect 5813 8693 5827 8707
rect 5773 8493 5787 8507
rect 5733 8453 5747 8467
rect 5753 8433 5767 8447
rect 5733 7813 5747 7827
rect 5933 8773 5947 8787
rect 5913 8733 5927 8747
rect 5953 8733 5967 8747
rect 5973 8733 5987 8747
rect 5873 8573 5887 8587
rect 5833 8433 5847 8447
rect 5833 8353 5847 8367
rect 5853 8313 5867 8327
rect 5773 8273 5787 8287
rect 5793 8273 5807 8287
rect 5773 8133 5787 8147
rect 5953 8553 5967 8567
rect 5893 8493 5907 8507
rect 5933 8413 5947 8427
rect 5973 8393 5987 8407
rect 5953 8373 5967 8387
rect 5913 8333 5927 8347
rect 5853 8053 5867 8067
rect 5793 8033 5807 8047
rect 5833 8033 5847 8047
rect 5773 8013 5787 8027
rect 5753 7673 5767 7687
rect 5933 8073 5947 8087
rect 5913 7953 5927 7967
rect 5793 7933 5807 7947
rect 5873 7933 5887 7947
rect 5973 8353 5987 8367
rect 5993 8333 6007 8347
rect 6093 8773 6107 8787
rect 6073 8593 6087 8607
rect 6053 8513 6067 8527
rect 6213 9433 6227 9447
rect 6193 9413 6207 9427
rect 6173 9293 6187 9307
rect 6153 9133 6167 9147
rect 6273 9293 6287 9307
rect 6253 9273 6267 9287
rect 6213 9213 6227 9227
rect 6213 9073 6227 9087
rect 6173 9013 6187 9027
rect 6173 8933 6187 8947
rect 6193 8813 6207 8827
rect 6153 8793 6167 8807
rect 6193 8793 6207 8807
rect 6133 8773 6147 8787
rect 6173 8773 6187 8787
rect 6113 8733 6127 8747
rect 6173 8513 6187 8527
rect 6113 8493 6127 8507
rect 6153 8493 6167 8507
rect 6073 8273 6087 8287
rect 6033 8213 6047 8227
rect 6113 8093 6127 8107
rect 6093 8053 6107 8067
rect 6053 8033 6067 8047
rect 6073 8013 6087 8027
rect 6033 7993 6047 8007
rect 6073 7993 6087 8007
rect 5953 7973 5967 7987
rect 5973 7973 5987 7987
rect 6013 7973 6027 7987
rect 5933 7913 5947 7927
rect 5993 7853 6007 7867
rect 5853 7833 5867 7847
rect 5793 7533 5807 7547
rect 5753 7433 5767 7447
rect 5773 7373 5787 7387
rect 5753 7353 5767 7367
rect 5993 7813 6007 7827
rect 5853 7793 5867 7807
rect 5973 7713 5987 7727
rect 5913 7693 5927 7707
rect 5893 7573 5907 7587
rect 5893 7533 5907 7547
rect 5853 7513 5867 7527
rect 5833 7493 5847 7507
rect 5833 7353 5847 7367
rect 5753 7113 5767 7127
rect 5693 7093 5707 7107
rect 5653 7073 5667 7087
rect 5713 7073 5727 7087
rect 5713 7053 5727 7067
rect 5833 7133 5847 7147
rect 5953 7673 5967 7687
rect 5973 7673 5987 7687
rect 5933 7573 5947 7587
rect 5973 7573 5987 7587
rect 5953 7553 5967 7567
rect 5973 7333 5987 7347
rect 5933 7233 5947 7247
rect 5873 7173 5887 7187
rect 5933 7153 5947 7167
rect 5833 7093 5847 7107
rect 5853 7093 5867 7107
rect 5893 7093 5907 7107
rect 5653 7033 5667 7047
rect 5613 6793 5627 6807
rect 5633 6793 5647 6807
rect 5553 6613 5567 6627
rect 5533 6593 5547 6607
rect 5613 6593 5627 6607
rect 5653 6593 5667 6607
rect 5533 6533 5547 6547
rect 5533 6433 5547 6447
rect 5513 6413 5527 6427
rect 5553 6373 5567 6387
rect 5453 5893 5467 5907
rect 5433 5753 5447 5767
rect 5573 6353 5587 6367
rect 5533 6213 5547 6227
rect 5513 6173 5527 6187
rect 5573 6313 5587 6327
rect 5553 6133 5567 6147
rect 5553 6093 5567 6107
rect 5513 6073 5527 6087
rect 5533 5933 5547 5947
rect 5513 5913 5527 5927
rect 5653 6573 5667 6587
rect 5633 6333 5647 6347
rect 5633 6273 5647 6287
rect 5613 6193 5627 6207
rect 5613 6093 5627 6107
rect 5593 5953 5607 5967
rect 5593 5913 5607 5927
rect 5573 5893 5587 5907
rect 5573 5753 5587 5767
rect 5493 5733 5507 5747
rect 5473 5713 5487 5727
rect 5473 5633 5487 5647
rect 5513 5633 5527 5647
rect 5553 5633 5567 5647
rect 5493 5613 5507 5627
rect 5453 5533 5467 5547
rect 5413 5513 5427 5527
rect 5473 5473 5487 5487
rect 5393 5453 5407 5467
rect 5453 5453 5467 5467
rect 5433 5433 5447 5447
rect 5533 5593 5547 5607
rect 5513 5553 5527 5567
rect 5453 5413 5467 5427
rect 5493 5413 5507 5427
rect 5293 5353 5307 5367
rect 5313 5353 5327 5367
rect 5293 5213 5307 5227
rect 5073 4973 5087 4987
rect 5033 4953 5047 4967
rect 5073 4953 5087 4967
rect 5173 5133 5187 5147
rect 5193 5133 5207 5147
rect 5353 5333 5367 5347
rect 5353 5233 5367 5247
rect 5313 5173 5327 5187
rect 5373 5173 5387 5187
rect 5333 5153 5347 5167
rect 5233 5093 5247 5107
rect 5153 4973 5167 4987
rect 5053 4933 5067 4947
rect 5133 4933 5147 4947
rect 5093 4913 5107 4927
rect 5033 4853 5047 4867
rect 5093 4853 5107 4867
rect 5073 4773 5087 4787
rect 4993 4713 5007 4727
rect 5033 4673 5047 4687
rect 5013 4653 5027 4667
rect 4913 4613 4927 4627
rect 4733 4133 4747 4147
rect 4693 3973 4707 3987
rect 4713 3973 4727 3987
rect 4673 3753 4687 3767
rect 4713 3733 4727 3747
rect 4673 3713 4687 3727
rect 4693 3533 4707 3547
rect 5053 4633 5067 4647
rect 4993 4613 5007 4627
rect 5033 4573 5047 4587
rect 4993 4193 5007 4207
rect 4993 4173 5007 4187
rect 4973 4113 4987 4127
rect 4973 4073 4987 4087
rect 4933 3993 4947 4007
rect 4773 3973 4787 3987
rect 4813 3973 4827 3987
rect 4913 3833 4927 3847
rect 4813 3773 4827 3787
rect 4833 3733 4847 3747
rect 4753 3713 4767 3727
rect 4673 3493 4687 3507
rect 4653 3133 4667 3147
rect 4633 3053 4647 3067
rect 4653 3033 4667 3047
rect 4593 2773 4607 2787
rect 4633 2753 4647 2767
rect 4633 2573 4647 2587
rect 4613 2533 4627 2547
rect 4653 2533 4667 2547
rect 4713 3373 4727 3387
rect 4833 3253 4847 3267
rect 4993 3953 5007 3967
rect 5033 4173 5047 4187
rect 5053 3853 5067 3867
rect 5213 4953 5227 4967
rect 5213 4813 5227 4827
rect 5213 4693 5227 4707
rect 5193 4653 5207 4667
rect 5153 4593 5167 4607
rect 5213 4493 5227 4507
rect 5193 4473 5207 4487
rect 5133 4453 5147 4467
rect 5173 4453 5187 4467
rect 5173 4433 5187 4447
rect 5133 4413 5147 4427
rect 5153 4193 5167 4207
rect 5353 5073 5367 5087
rect 5293 5013 5307 5027
rect 5253 4953 5267 4967
rect 5273 4933 5287 4947
rect 5413 5393 5427 5407
rect 5453 5393 5467 5407
rect 5413 5333 5427 5347
rect 5413 5293 5427 5307
rect 5313 4833 5327 4847
rect 5393 4833 5407 4847
rect 5453 5153 5467 5167
rect 5433 4953 5447 4967
rect 5413 4753 5427 4767
rect 5333 4713 5347 4727
rect 5293 4693 5307 4707
rect 5293 4653 5307 4667
rect 5253 4613 5267 4627
rect 5093 4173 5107 4187
rect 5113 4153 5127 4167
rect 5213 4133 5227 4147
rect 5253 4113 5267 4127
rect 5253 4033 5267 4047
rect 5373 4653 5387 4667
rect 5393 4633 5407 4647
rect 5413 4613 5427 4627
rect 5513 5293 5527 5307
rect 5533 5173 5547 5187
rect 5513 5153 5527 5167
rect 5533 5113 5547 5127
rect 5533 4993 5547 5007
rect 5493 4973 5507 4987
rect 5473 4953 5487 4967
rect 5513 4953 5527 4967
rect 5493 4933 5507 4947
rect 5493 4913 5507 4927
rect 5353 4533 5367 4547
rect 5373 4413 5387 4427
rect 5373 4333 5387 4347
rect 5573 5613 5587 5627
rect 5613 5513 5627 5527
rect 5693 7013 5707 7027
rect 5693 6893 5707 6907
rect 5773 7033 5787 7047
rect 5753 6993 5767 7007
rect 5733 6913 5747 6927
rect 5713 6853 5727 6867
rect 5733 6853 5747 6867
rect 5693 6813 5707 6827
rect 5693 6793 5707 6807
rect 5733 6793 5747 6807
rect 5713 6613 5727 6627
rect 5693 6573 5707 6587
rect 5713 6513 5727 6527
rect 5753 6593 5767 6607
rect 5793 6993 5807 7007
rect 5813 6913 5827 6927
rect 5873 7073 5887 7087
rect 5773 6473 5787 6487
rect 5693 6293 5707 6307
rect 5753 6353 5767 6367
rect 5733 6333 5747 6347
rect 5713 6133 5727 6147
rect 5753 6153 5767 6167
rect 5833 6593 5847 6607
rect 5813 6373 5827 6387
rect 5813 6253 5827 6267
rect 5793 6153 5807 6167
rect 5793 6133 5807 6147
rect 5653 6093 5667 6107
rect 5653 6073 5667 6087
rect 5753 6113 5767 6127
rect 5773 6113 5787 6127
rect 5693 6093 5707 6107
rect 5673 5853 5687 5867
rect 5673 5753 5687 5767
rect 5673 5553 5687 5567
rect 5753 6073 5767 6087
rect 5793 6053 5807 6067
rect 5733 5913 5747 5927
rect 5733 5873 5747 5887
rect 5753 5873 5767 5887
rect 5813 5873 5827 5887
rect 5773 5813 5787 5827
rect 5753 5773 5767 5787
rect 5753 5633 5767 5647
rect 5813 5733 5827 5747
rect 5713 5613 5727 5627
rect 5813 5613 5827 5627
rect 5753 5593 5767 5607
rect 5753 5553 5767 5567
rect 5693 5533 5707 5547
rect 5773 5533 5787 5547
rect 5753 5513 5767 5527
rect 5693 5473 5707 5487
rect 5673 5453 5687 5467
rect 5733 5453 5747 5467
rect 5653 5433 5667 5447
rect 5633 5413 5647 5427
rect 5713 5433 5727 5447
rect 5693 5413 5707 5427
rect 5693 5353 5707 5367
rect 5613 5293 5627 5307
rect 5713 5293 5727 5307
rect 5593 5153 5607 5167
rect 5653 5253 5667 5267
rect 5693 5193 5707 5207
rect 5693 5173 5707 5187
rect 5673 5133 5687 5147
rect 5713 5133 5727 5147
rect 5633 5093 5647 5107
rect 5613 5033 5627 5047
rect 5593 4933 5607 4947
rect 5653 4993 5667 5007
rect 5673 4933 5687 4947
rect 5613 4853 5627 4867
rect 5573 4813 5587 4827
rect 5573 4693 5587 4707
rect 5653 4813 5667 4827
rect 5453 4513 5467 4527
rect 5533 4513 5547 4527
rect 5393 4153 5407 4167
rect 5213 4013 5227 4027
rect 5333 4013 5347 4027
rect 5013 3733 5027 3747
rect 4893 3673 4907 3687
rect 4933 3673 4947 3687
rect 4893 3653 4907 3667
rect 4973 3513 4987 3527
rect 4853 3113 4867 3127
rect 4753 3093 4767 3107
rect 4813 3073 4827 3087
rect 4693 3053 4707 3067
rect 4713 3033 4727 3047
rect 4793 3013 4807 3027
rect 4833 3013 4847 3027
rect 4753 2973 4767 2987
rect 4893 3233 4907 3247
rect 5113 3953 5127 3967
rect 5093 3753 5107 3767
rect 5073 3693 5087 3707
rect 5193 3653 5207 3667
rect 5173 3613 5187 3627
rect 5193 3533 5207 3547
rect 5013 3493 5027 3507
rect 5053 3493 5067 3507
rect 5133 3473 5147 3487
rect 5313 3993 5327 4007
rect 5393 3993 5407 4007
rect 5333 3953 5347 3967
rect 5533 4493 5547 4507
rect 5553 4493 5567 4507
rect 5473 4473 5487 4487
rect 5513 4473 5527 4487
rect 5453 4153 5467 4167
rect 5593 4653 5607 4667
rect 5513 4153 5527 4167
rect 5633 4193 5647 4207
rect 5593 4173 5607 4187
rect 5573 4153 5587 4167
rect 5553 4013 5567 4027
rect 5473 3993 5487 4007
rect 5633 4013 5647 4027
rect 5493 3973 5507 3987
rect 5533 3973 5547 3987
rect 5573 3973 5587 3987
rect 5433 3913 5447 3927
rect 5533 3773 5547 3787
rect 5533 3733 5547 3747
rect 5313 3613 5327 3627
rect 5253 3553 5267 3567
rect 5213 3333 5227 3347
rect 5173 3233 5187 3247
rect 5353 3533 5367 3547
rect 5373 3493 5387 3507
rect 5633 3633 5647 3647
rect 5593 3533 5607 3547
rect 5553 3513 5567 3527
rect 5573 3493 5587 3507
rect 5733 4893 5747 4907
rect 5793 5513 5807 5527
rect 5773 5273 5787 5287
rect 5773 5253 5787 5267
rect 5753 4813 5767 4827
rect 5733 4753 5747 4767
rect 5953 7053 5967 7067
rect 5893 7013 5907 7027
rect 5873 6853 5887 6867
rect 5973 6913 5987 6927
rect 5913 6893 5927 6907
rect 5933 6873 5947 6887
rect 5913 6853 5927 6867
rect 5953 6853 5967 6867
rect 5953 6833 5967 6847
rect 5933 6813 5947 6827
rect 5893 6733 5907 6747
rect 5913 6533 5927 6547
rect 5873 6433 5887 6447
rect 5853 5853 5867 5867
rect 5853 5833 5867 5847
rect 6073 7893 6087 7907
rect 6093 7893 6107 7907
rect 6233 8453 6247 8467
rect 6193 8333 6207 8347
rect 6173 8313 6187 8327
rect 6393 9753 6407 9767
rect 6453 9753 6467 9767
rect 6373 9733 6387 9747
rect 6333 9713 6347 9727
rect 6313 9493 6327 9507
rect 6313 9213 6327 9227
rect 6453 9693 6467 9707
rect 6753 11693 6767 11707
rect 6713 11613 6727 11627
rect 6733 11613 6747 11627
rect 6693 11573 6707 11587
rect 6613 11393 6627 11407
rect 6653 11393 6667 11407
rect 6633 11373 6647 11387
rect 6733 11373 6747 11387
rect 6653 11273 6667 11287
rect 6573 11213 6587 11227
rect 6553 11133 6567 11147
rect 6773 11553 6787 11567
rect 6773 11373 6787 11387
rect 6913 11893 6927 11907
rect 7133 11893 7147 11907
rect 6873 11873 6887 11887
rect 7013 11873 7027 11887
rect 7093 11873 7107 11887
rect 7313 11873 7327 11887
rect 7353 11873 7367 11887
rect 7453 11873 7467 11887
rect 6933 11833 6947 11847
rect 6893 11753 6907 11767
rect 6813 11673 6827 11687
rect 6853 11673 6867 11687
rect 6893 11673 6907 11687
rect 6833 11613 6847 11627
rect 6893 11593 6907 11607
rect 6813 11373 6827 11387
rect 6833 11353 6847 11367
rect 6793 11333 6807 11347
rect 6733 11013 6747 11027
rect 6753 10913 6767 10927
rect 6793 11153 6807 11167
rect 6833 11153 6847 11167
rect 6673 10893 6687 10907
rect 6773 10893 6787 10907
rect 6493 10833 6507 10847
rect 6593 10813 6607 10827
rect 6773 10813 6787 10827
rect 6613 10753 6627 10767
rect 6553 10713 6567 10727
rect 6593 10713 6607 10727
rect 6493 10433 6507 10447
rect 6533 10433 6547 10447
rect 6553 10393 6567 10407
rect 6513 10373 6527 10387
rect 6553 10253 6567 10267
rect 6513 10233 6527 10247
rect 6493 10173 6507 10187
rect 6593 10213 6607 10227
rect 6573 10093 6587 10107
rect 6493 10073 6507 10087
rect 6473 9673 6487 9687
rect 6433 9633 6447 9647
rect 6413 9573 6427 9587
rect 6353 9493 6367 9507
rect 6373 9473 6387 9487
rect 6413 9453 6427 9467
rect 6453 9353 6467 9367
rect 6433 9333 6447 9347
rect 6413 9313 6427 9327
rect 6373 9273 6387 9287
rect 6353 8973 6367 8987
rect 6553 9953 6567 9967
rect 6513 9893 6527 9907
rect 6533 9773 6547 9787
rect 6633 10453 6647 10467
rect 6733 10433 6747 10447
rect 6753 10413 6767 10427
rect 6713 10373 6727 10387
rect 6733 10233 6747 10247
rect 6773 10213 6787 10227
rect 6653 10193 6667 10207
rect 6713 10193 6727 10207
rect 6813 11093 6827 11107
rect 6913 11353 6927 11367
rect 7073 11853 7087 11867
rect 7113 11853 7127 11867
rect 7153 11833 7167 11847
rect 7053 11813 7067 11827
rect 7373 11833 7387 11847
rect 7333 11813 7347 11827
rect 7293 11773 7307 11787
rect 7373 11773 7387 11787
rect 7113 11653 7127 11667
rect 7173 11653 7187 11667
rect 7033 11633 7047 11647
rect 6993 11613 7007 11627
rect 6953 11393 6967 11407
rect 6973 11373 6987 11387
rect 7073 11473 7087 11487
rect 7073 11413 7087 11427
rect 6953 11353 6967 11367
rect 6933 11033 6947 11047
rect 6893 10993 6907 11007
rect 6853 10953 6867 10967
rect 7013 11213 7027 11227
rect 6993 11193 7007 11207
rect 7053 11193 7067 11207
rect 7213 11413 7227 11427
rect 7093 11393 7107 11407
rect 7133 11393 7147 11407
rect 7033 11173 7047 11187
rect 7073 11173 7087 11187
rect 7053 11033 7067 11047
rect 7033 10973 7047 10987
rect 6973 10933 6987 10947
rect 7013 10933 7027 10947
rect 7033 10893 7047 10907
rect 6853 10853 6867 10867
rect 6953 10693 6967 10707
rect 7013 10873 7027 10887
rect 6993 10813 7007 10827
rect 6913 10433 6927 10447
rect 6973 10413 6987 10427
rect 6993 10413 7007 10427
rect 6953 10393 6967 10407
rect 7033 10813 7047 10827
rect 7013 10393 7027 10407
rect 6973 10373 6987 10387
rect 6913 10293 6927 10307
rect 6893 10253 6907 10267
rect 6893 10233 6907 10247
rect 7033 10273 7047 10287
rect 6953 10233 6967 10247
rect 6933 10213 6947 10227
rect 6793 10053 6807 10067
rect 6853 10053 6867 10067
rect 6713 9973 6727 9987
rect 6753 9953 6767 9967
rect 6673 9933 6687 9947
rect 6633 9913 6647 9927
rect 6773 9773 6787 9787
rect 6613 9753 6627 9767
rect 6653 9753 6667 9767
rect 6813 9753 6827 9767
rect 6573 9713 6587 9727
rect 6833 9733 6847 9747
rect 6793 9713 6807 9727
rect 6633 9693 6647 9707
rect 6593 9653 6607 9667
rect 6513 9433 6527 9447
rect 6733 9473 6747 9487
rect 6593 9453 6607 9467
rect 6713 9453 6727 9467
rect 6753 9433 6767 9447
rect 6833 9473 6847 9487
rect 6833 9433 6847 9447
rect 6553 9413 6567 9427
rect 6773 9413 6787 9427
rect 6613 9333 6627 9347
rect 6593 9293 6607 9307
rect 6573 9273 6587 9287
rect 6753 9313 6767 9327
rect 6793 9293 6807 9307
rect 6833 9293 6847 9307
rect 6433 9253 6447 9267
rect 6493 9253 6507 9267
rect 6733 9253 6747 9267
rect 6573 9193 6587 9207
rect 6433 9013 6447 9027
rect 6453 8993 6467 9007
rect 6373 8953 6387 8967
rect 6353 8933 6367 8947
rect 6533 8893 6547 8907
rect 6353 8853 6367 8867
rect 6353 8813 6367 8827
rect 6393 8793 6407 8807
rect 6373 8773 6387 8787
rect 6373 8633 6387 8647
rect 6473 8793 6487 8807
rect 6533 8793 6547 8807
rect 6413 8593 6427 8607
rect 6313 8573 6327 8587
rect 6273 8553 6287 8567
rect 6333 8553 6347 8567
rect 6313 8513 6327 8527
rect 6253 8353 6267 8367
rect 6213 8293 6227 8307
rect 6253 8293 6267 8307
rect 6153 8073 6167 8087
rect 6153 8013 6167 8027
rect 6273 8133 6287 8147
rect 6193 8053 6207 8067
rect 6173 7813 6187 7827
rect 6033 7653 6047 7667
rect 6013 7533 6027 7547
rect 6053 7473 6067 7487
rect 6033 7373 6047 7387
rect 6013 7113 6027 7127
rect 6013 6893 6027 6907
rect 6013 6853 6027 6867
rect 6013 6833 6027 6847
rect 5973 6753 5987 6767
rect 5993 6753 6007 6767
rect 6013 6633 6027 6647
rect 6013 6593 6027 6607
rect 6153 7613 6167 7627
rect 6113 7553 6127 7567
rect 6153 7553 6167 7567
rect 6113 7473 6127 7487
rect 6073 7453 6087 7467
rect 6093 7453 6107 7467
rect 6173 7533 6187 7547
rect 6213 7993 6227 8007
rect 6213 7573 6227 7587
rect 6193 7473 6207 7487
rect 6133 7433 6147 7447
rect 6253 7973 6267 7987
rect 6513 8733 6527 8747
rect 6553 8733 6567 8747
rect 6353 8413 6367 8427
rect 6353 8373 6367 8387
rect 6393 8313 6407 8327
rect 6373 8293 6387 8307
rect 6413 8273 6427 8287
rect 6513 8493 6527 8507
rect 6513 8433 6527 8447
rect 6493 8393 6507 8407
rect 6493 8313 6507 8327
rect 6473 8173 6487 8187
rect 6373 8133 6387 8147
rect 6413 8133 6427 8147
rect 6453 8133 6467 8147
rect 6333 8053 6347 8067
rect 6453 8073 6467 8087
rect 6413 8053 6427 8067
rect 6493 8053 6507 8067
rect 6373 8033 6387 8047
rect 6433 8033 6447 8047
rect 6293 7913 6307 7927
rect 6293 7873 6307 7887
rect 6333 7853 6347 7867
rect 6293 7833 6307 7847
rect 6373 7833 6387 7847
rect 6353 7813 6367 7827
rect 6313 7793 6327 7807
rect 6413 8013 6427 8027
rect 6453 8013 6467 8027
rect 6433 7993 6447 8007
rect 6413 7873 6427 7887
rect 6533 8333 6547 8347
rect 6813 9253 6827 9267
rect 6873 9953 6887 9967
rect 7073 10913 7087 10927
rect 7153 11373 7167 11387
rect 7313 11433 7327 11447
rect 7273 11373 7287 11387
rect 7393 11413 7407 11427
rect 7373 11393 7387 11407
rect 7333 11313 7347 11327
rect 7353 11253 7367 11267
rect 7313 11193 7327 11207
rect 7193 11173 7207 11187
rect 7153 11153 7167 11167
rect 7353 11173 7367 11187
rect 7373 11113 7387 11127
rect 7393 11073 7407 11087
rect 7133 11053 7147 11067
rect 7173 10953 7187 10967
rect 7393 10953 7407 10967
rect 7213 10933 7227 10947
rect 7113 10893 7127 10907
rect 7233 10913 7247 10927
rect 7353 10913 7367 10927
rect 7073 10733 7087 10747
rect 7333 10893 7347 10907
rect 7373 10873 7387 10887
rect 7233 10793 7247 10807
rect 7413 10793 7427 10807
rect 7153 10753 7167 10767
rect 7293 10753 7307 10767
rect 7153 10733 7167 10747
rect 7113 10713 7127 10727
rect 7093 10693 7107 10707
rect 7073 10653 7087 10667
rect 7073 10473 7087 10487
rect 7073 10373 7087 10387
rect 7053 10253 7067 10267
rect 7133 10333 7147 10347
rect 7093 10273 7107 10287
rect 7173 10693 7187 10707
rect 7273 10693 7287 10707
rect 7293 10433 7307 10447
rect 7173 10273 7187 10287
rect 7073 10233 7087 10247
rect 7153 10213 7167 10227
rect 7113 9973 7127 9987
rect 7153 9973 7167 9987
rect 6873 9913 6887 9927
rect 6953 9853 6967 9867
rect 6873 9733 6887 9747
rect 6993 9793 7007 9807
rect 6973 9773 6987 9787
rect 7033 9713 7047 9727
rect 6953 9673 6967 9687
rect 6973 9633 6987 9647
rect 7033 9633 7047 9647
rect 7013 9493 7027 9507
rect 6873 9473 6887 9487
rect 6933 9473 6947 9487
rect 6973 9473 6987 9487
rect 6953 9453 6967 9467
rect 6973 9393 6987 9407
rect 6873 9353 6887 9367
rect 6853 9253 6867 9267
rect 6773 9153 6787 9167
rect 6633 9093 6647 9107
rect 6733 9093 6747 9107
rect 6993 9293 7007 9307
rect 6933 9233 6947 9247
rect 6933 9213 6947 9227
rect 6873 9173 6887 9187
rect 6933 9133 6947 9147
rect 6833 9113 6847 9127
rect 6653 8993 6667 9007
rect 6773 9013 6787 9027
rect 6813 9013 6827 9027
rect 6873 9013 6887 9027
rect 6693 8993 6707 9007
rect 6893 8993 6907 9007
rect 6673 8973 6687 8987
rect 6853 8973 6867 8987
rect 6673 8953 6687 8967
rect 6773 8853 6787 8867
rect 6753 8833 6767 8847
rect 6693 8813 6707 8827
rect 6713 8793 6727 8807
rect 6673 8633 6687 8647
rect 6633 8593 6647 8607
rect 6573 8553 6587 8567
rect 6713 8513 6727 8527
rect 6693 8493 6707 8507
rect 6733 8493 6747 8507
rect 6613 8373 6627 8387
rect 6553 8313 6567 8327
rect 6613 8313 6627 8327
rect 6753 8433 6767 8447
rect 6753 8333 6767 8347
rect 6793 8813 6807 8827
rect 6773 8313 6787 8327
rect 6533 8293 6547 8307
rect 6573 8293 6587 8307
rect 6593 8233 6607 8247
rect 6573 8173 6587 8187
rect 6533 8013 6547 8027
rect 6513 7853 6527 7867
rect 6393 7793 6407 7807
rect 6513 7793 6527 7807
rect 6553 7793 6567 7807
rect 6373 7773 6387 7787
rect 6233 7413 6247 7427
rect 6133 7373 6147 7387
rect 6173 7373 6187 7387
rect 6053 7333 6067 7347
rect 6073 7153 6087 7167
rect 6053 7053 6067 7067
rect 5953 6453 5967 6467
rect 5893 6353 5907 6367
rect 5933 6353 5947 6367
rect 5933 6253 5947 6267
rect 5933 6173 5947 6187
rect 5913 6053 5927 6067
rect 5933 5933 5947 5947
rect 5993 6533 6007 6547
rect 5993 6393 6007 6407
rect 5973 6373 5987 6387
rect 5973 6353 5987 6367
rect 5953 5913 5967 5927
rect 5913 5893 5927 5907
rect 5993 6293 6007 6307
rect 5993 6013 6007 6027
rect 5893 5873 5907 5887
rect 5913 5873 5927 5887
rect 5893 5833 5907 5847
rect 5873 5793 5887 5807
rect 5853 5773 5867 5787
rect 5893 5733 5907 5747
rect 5893 5653 5907 5667
rect 5993 5853 6007 5867
rect 5973 5653 5987 5667
rect 5913 5633 5927 5647
rect 5953 5633 5967 5647
rect 5893 5613 5907 5627
rect 5893 5593 5907 5607
rect 5833 5453 5847 5467
rect 5853 5433 5867 5447
rect 5913 5433 5927 5447
rect 5833 5413 5847 5427
rect 5933 5413 5947 5427
rect 5873 5393 5887 5407
rect 5913 5393 5927 5407
rect 5833 5353 5847 5367
rect 5853 5273 5867 5287
rect 5833 5173 5847 5187
rect 5833 5153 5847 5167
rect 5813 5093 5827 5107
rect 5793 4953 5807 4967
rect 5753 4673 5767 4687
rect 5793 4633 5807 4647
rect 5833 4953 5847 4967
rect 5873 5213 5887 5227
rect 5893 5113 5907 5127
rect 5913 5073 5927 5087
rect 5913 5033 5927 5047
rect 5933 4973 5947 4987
rect 5873 4953 5887 4967
rect 5833 4853 5847 4867
rect 5893 4853 5907 4867
rect 5673 4193 5687 4207
rect 5753 4573 5767 4587
rect 5813 4573 5827 4587
rect 5713 4533 5727 4547
rect 5713 4513 5727 4527
rect 5733 4493 5747 4507
rect 5793 4493 5807 4507
rect 5773 4453 5787 4467
rect 5753 4213 5767 4227
rect 5713 4193 5727 4207
rect 5693 4133 5707 4147
rect 5793 4213 5807 4227
rect 5833 4213 5847 4227
rect 5773 4193 5787 4207
rect 5813 4193 5827 4207
rect 5753 4153 5767 4167
rect 5733 3973 5747 3987
rect 6073 7013 6087 7027
rect 6073 6793 6087 6807
rect 6113 7313 6127 7327
rect 6153 7233 6167 7247
rect 6113 7073 6127 7087
rect 6193 7313 6207 7327
rect 6173 7173 6187 7187
rect 6213 7293 6227 7307
rect 6213 7233 6227 7247
rect 6193 7113 6207 7127
rect 6233 7073 6247 7087
rect 6133 7053 6147 7067
rect 6173 7013 6187 7027
rect 6173 6993 6187 7007
rect 6133 6853 6147 6867
rect 6113 6773 6127 6787
rect 6113 6593 6127 6607
rect 6113 6533 6127 6547
rect 6193 6853 6207 6867
rect 6193 6813 6207 6827
rect 6273 7493 6287 7507
rect 6293 7493 6307 7507
rect 6453 7453 6467 7467
rect 6293 7413 6307 7427
rect 6253 6993 6267 7007
rect 6253 6933 6267 6947
rect 6893 8813 6907 8827
rect 6873 8773 6887 8787
rect 6873 8753 6887 8767
rect 6813 8613 6827 8627
rect 6853 8613 6867 8627
rect 6833 8593 6847 8607
rect 6813 8553 6827 8567
rect 6813 8513 6827 8527
rect 6873 8513 6887 8527
rect 6893 8493 6907 8507
rect 6913 8453 6927 8467
rect 6873 8433 6887 8447
rect 6853 8333 6867 8347
rect 6813 8273 6827 8287
rect 6793 8173 6807 8187
rect 6633 8113 6647 8127
rect 6813 8113 6827 8127
rect 6593 8053 6607 8067
rect 6753 8093 6767 8107
rect 6613 8013 6627 8027
rect 6593 7833 6607 7847
rect 6593 7793 6607 7807
rect 6613 7613 6627 7627
rect 6633 7613 6647 7627
rect 6473 7433 6487 7447
rect 6493 7233 6507 7247
rect 6433 7153 6447 7167
rect 6453 7153 6467 7167
rect 6373 7093 6387 7107
rect 6433 7093 6447 7107
rect 6633 7413 6647 7427
rect 6633 7373 6647 7387
rect 6693 8053 6707 8067
rect 6673 7933 6687 7947
rect 6753 8013 6767 8027
rect 6733 7833 6747 7847
rect 6713 7793 6727 7807
rect 6733 7673 6747 7687
rect 6693 7593 6707 7607
rect 6553 7173 6567 7187
rect 6593 7173 6607 7187
rect 6533 7113 6547 7127
rect 6553 7093 6567 7107
rect 6333 6993 6347 7007
rect 6313 6893 6327 6907
rect 6353 6913 6367 6927
rect 6313 6853 6327 6867
rect 6433 6853 6447 6867
rect 6273 6833 6287 6847
rect 6253 6753 6267 6767
rect 6173 6633 6187 6647
rect 6153 6553 6167 6567
rect 6153 6473 6167 6487
rect 6213 6573 6227 6587
rect 6193 6533 6207 6547
rect 6193 6513 6207 6527
rect 6173 6413 6187 6427
rect 6393 6733 6407 6747
rect 6293 6713 6307 6727
rect 6233 6413 6247 6427
rect 6273 6413 6287 6427
rect 6193 6393 6207 6407
rect 6133 6293 6147 6307
rect 6193 6273 6207 6287
rect 6173 6253 6187 6267
rect 6113 6173 6127 6187
rect 6093 6133 6107 6147
rect 6033 5933 6047 5947
rect 6053 5913 6067 5927
rect 6033 5633 6047 5647
rect 6033 5613 6047 5627
rect 6033 5573 6047 5587
rect 5993 5553 6007 5567
rect 6013 5553 6027 5567
rect 6133 6013 6147 6027
rect 6153 6013 6167 6027
rect 6133 5973 6147 5987
rect 6133 5933 6147 5947
rect 6173 5973 6187 5987
rect 6273 6373 6287 6387
rect 6233 6353 6247 6367
rect 6213 6193 6227 6207
rect 6213 6133 6227 6147
rect 6213 6093 6227 6107
rect 6093 5873 6107 5887
rect 6073 5753 6087 5767
rect 6093 5753 6107 5767
rect 6053 5513 6067 5527
rect 6033 5453 6047 5467
rect 6073 5433 6087 5447
rect 5973 5273 5987 5287
rect 6053 5413 6067 5427
rect 5973 5233 5987 5247
rect 5993 5233 6007 5247
rect 5953 4913 5967 4927
rect 6073 5253 6087 5267
rect 6153 5873 6167 5887
rect 6173 5833 6187 5847
rect 6153 5813 6167 5827
rect 6173 5813 6187 5827
rect 6113 5733 6127 5747
rect 6133 5733 6147 5747
rect 6153 5653 6167 5667
rect 6133 5633 6147 5647
rect 6153 5553 6167 5567
rect 6133 5493 6147 5507
rect 6113 5373 6127 5387
rect 6113 5293 6127 5307
rect 6113 5193 6127 5207
rect 6053 5133 6067 5147
rect 6033 5113 6047 5127
rect 6013 5013 6027 5027
rect 6093 5113 6107 5127
rect 6053 5073 6067 5087
rect 6093 5033 6107 5047
rect 6053 4973 6067 4987
rect 6093 4973 6107 4987
rect 6033 4933 6047 4947
rect 6073 4933 6087 4947
rect 6033 4913 6047 4927
rect 5973 4853 5987 4867
rect 5933 4693 5947 4707
rect 5933 4673 5947 4687
rect 5913 4653 5927 4667
rect 5953 4653 5967 4667
rect 5973 4653 5987 4667
rect 5933 4633 5947 4647
rect 5893 4613 5907 4627
rect 5953 4573 5967 4587
rect 5933 4533 5947 4547
rect 5973 4493 5987 4507
rect 5873 4453 5887 4467
rect 5953 4453 5967 4467
rect 5913 4433 5927 4447
rect 5873 4213 5887 4227
rect 5993 4233 6007 4247
rect 6013 4213 6027 4227
rect 5873 4173 5887 4187
rect 5993 4173 6007 4187
rect 6013 4133 6027 4147
rect 5933 4013 5947 4027
rect 5853 3973 5867 3987
rect 5773 3953 5787 3967
rect 5913 3933 5927 3947
rect 5673 3633 5687 3647
rect 5693 3573 5707 3587
rect 5653 3553 5667 3567
rect 5693 3493 5707 3507
rect 5853 3673 5867 3687
rect 5753 3573 5767 3587
rect 5733 3553 5747 3567
rect 5773 3533 5787 3547
rect 5833 3513 5847 3527
rect 5733 3473 5747 3487
rect 5693 3413 5707 3427
rect 5493 3353 5507 3367
rect 5313 3253 5327 3267
rect 5333 3173 5347 3187
rect 4913 3093 4927 3107
rect 4893 3053 4907 3067
rect 4893 2953 4907 2967
rect 4753 2773 4767 2787
rect 4733 2753 4747 2767
rect 4813 2753 4827 2767
rect 4713 2713 4727 2727
rect 4693 2553 4707 2567
rect 4693 2473 4707 2487
rect 4673 2333 4687 2347
rect 4613 2253 4627 2267
rect 4633 2253 4647 2267
rect 4773 2713 4787 2727
rect 4813 2693 4827 2707
rect 4733 2673 4747 2687
rect 5153 3073 5167 3087
rect 4973 3053 4987 3067
rect 5253 2993 5267 3007
rect 5133 2913 5147 2927
rect 4933 2773 4947 2787
rect 4973 2753 4987 2767
rect 5013 2753 5027 2767
rect 4953 2673 4967 2687
rect 4873 2573 4887 2587
rect 4733 2473 4747 2487
rect 5053 2553 5067 2567
rect 5033 2493 5047 2507
rect 4673 2253 4687 2267
rect 4653 2193 4667 2207
rect 4613 2073 4627 2087
rect 4593 1773 4607 1787
rect 4593 1593 4607 1607
rect 4693 1593 4707 1607
rect 4713 1553 4727 1567
rect 4673 1373 4687 1387
rect 4713 1373 4727 1387
rect 4593 1313 4607 1327
rect 4653 1313 4667 1327
rect 4613 1233 4627 1247
rect 4693 1253 4707 1267
rect 4613 1133 4627 1147
rect 4673 1133 4687 1147
rect 4593 1053 4607 1067
rect 4613 853 4627 867
rect 4653 853 4667 867
rect 4713 853 4727 867
rect 4593 813 4607 827
rect 4533 333 4547 347
rect 4513 313 4527 327
rect 4513 273 4527 287
rect 4413 193 4427 207
rect 4373 173 4387 187
rect 4153 133 4167 147
rect 4133 113 4147 127
rect 4093 13 4107 27
rect 4133 13 4147 27
rect 4433 153 4447 167
rect 4473 153 4487 167
rect 4613 633 4627 647
rect 4593 613 4607 627
rect 4593 593 4607 607
rect 4633 333 4647 347
rect 4673 813 4687 827
rect 4713 813 4727 827
rect 4693 693 4707 707
rect 4893 2253 4907 2267
rect 4853 2233 4867 2247
rect 4833 2133 4847 2147
rect 4873 2033 4887 2047
rect 4753 1593 4767 1607
rect 5153 2793 5167 2807
rect 5173 2733 5187 2747
rect 5173 2593 5187 2607
rect 5213 2593 5227 2607
rect 5193 2553 5207 2567
rect 5233 2553 5247 2567
rect 5273 2833 5287 2847
rect 5273 2573 5287 2587
rect 5273 2553 5287 2567
rect 5293 2553 5307 2567
rect 5253 2493 5267 2507
rect 5173 2313 5187 2327
rect 5233 2313 5247 2327
rect 5213 2293 5227 2307
rect 5173 2273 5187 2287
rect 5133 2253 5147 2267
rect 5153 2253 5167 2267
rect 5053 2233 5067 2247
rect 4993 2113 5007 2127
rect 4953 2093 4967 2107
rect 4813 1773 4827 1787
rect 4853 1773 4867 1787
rect 4913 1773 4927 1787
rect 5013 1773 5027 1787
rect 4973 1733 4987 1747
rect 5033 1653 5047 1667
rect 4873 1613 4887 1627
rect 4933 1613 4947 1627
rect 5133 1913 5147 1927
rect 5053 1613 5067 1627
rect 4893 1573 4907 1587
rect 4873 1353 4887 1367
rect 4953 1553 4967 1567
rect 5093 1553 5107 1567
rect 5053 1353 5067 1367
rect 4953 1333 4967 1347
rect 5013 1333 5027 1347
rect 5073 1333 5087 1347
rect 4893 1313 4907 1327
rect 4993 1313 5007 1327
rect 4793 1133 4807 1147
rect 4753 1113 4767 1127
rect 5073 1293 5087 1307
rect 5033 1253 5047 1267
rect 4833 1193 4847 1207
rect 4953 1173 4967 1187
rect 4833 1133 4847 1147
rect 4853 1133 4867 1147
rect 4813 1053 4827 1067
rect 4853 1053 4867 1067
rect 4853 893 4867 907
rect 4893 853 4907 867
rect 4833 833 4847 847
rect 4813 813 4827 827
rect 4873 793 4887 807
rect 4813 693 4827 707
rect 4793 633 4807 647
rect 4773 613 4787 627
rect 4833 593 4847 607
rect 4913 833 4927 847
rect 4933 773 4947 787
rect 4913 653 4927 667
rect 4913 413 4927 427
rect 4893 393 4907 407
rect 4693 333 4707 347
rect 4733 333 4747 347
rect 4713 313 4727 327
rect 4693 173 4707 187
rect 4613 153 4627 167
rect 4653 153 4667 167
rect 4653 133 4667 147
rect 4633 113 4647 127
rect 4853 373 4867 387
rect 4853 353 4867 367
rect 4913 333 4927 347
rect 5073 1133 5087 1147
rect 4973 1073 4987 1087
rect 5033 1093 5047 1107
rect 5033 1073 5047 1087
rect 4993 1053 5007 1067
rect 5053 853 5067 867
rect 5093 853 5107 867
rect 5033 813 5047 827
rect 5053 813 5067 827
rect 4993 793 5007 807
rect 4973 653 4987 667
rect 4993 653 5007 667
rect 5073 773 5087 787
rect 5033 593 5047 607
rect 5013 393 5027 407
rect 5033 353 5047 367
rect 4953 333 4967 347
rect 5033 333 5047 347
rect 4933 313 4947 327
rect 4873 193 4887 207
rect 5073 313 5087 327
rect 5173 2233 5187 2247
rect 5213 2093 5227 2107
rect 5293 2273 5307 2287
rect 5253 2253 5267 2267
rect 5273 2253 5287 2267
rect 5173 1773 5187 1787
rect 5173 1633 5187 1647
rect 5233 1633 5247 1647
rect 5273 1653 5287 1667
rect 5273 1593 5287 1607
rect 5273 1393 5287 1407
rect 5193 1353 5207 1367
rect 5253 1353 5267 1367
rect 5233 1313 5247 1327
rect 5653 3233 5667 3247
rect 5473 3193 5487 3207
rect 5653 3113 5667 3127
rect 5373 2993 5387 3007
rect 5433 2853 5447 2867
rect 5353 2833 5367 2847
rect 5393 2833 5407 2847
rect 5373 2773 5387 2787
rect 5353 2733 5367 2747
rect 5373 2553 5387 2567
rect 5373 2253 5387 2267
rect 5753 3353 5767 3367
rect 5833 3193 5847 3207
rect 5713 3113 5727 3127
rect 5813 3053 5827 3067
rect 5693 2933 5707 2947
rect 5513 2753 5527 2767
rect 5533 2733 5547 2747
rect 5413 2713 5427 2727
rect 5513 2693 5527 2707
rect 5473 2093 5487 2107
rect 5453 2053 5467 2067
rect 5593 2753 5607 2767
rect 5573 2733 5587 2747
rect 5593 2613 5607 2627
rect 5613 2613 5627 2627
rect 5673 2553 5687 2567
rect 5573 2533 5587 2547
rect 5573 2493 5587 2507
rect 5593 2253 5607 2267
rect 5673 2473 5687 2487
rect 5693 2273 5707 2287
rect 5673 2093 5687 2107
rect 5413 1973 5427 1987
rect 5453 1973 5467 1987
rect 5333 1813 5347 1827
rect 5373 1793 5387 1807
rect 5393 1753 5407 1767
rect 5373 1613 5387 1627
rect 5353 1393 5367 1407
rect 5333 1353 5347 1367
rect 5213 1273 5227 1287
rect 5293 1293 5307 1307
rect 5293 1273 5307 1287
rect 5313 1273 5327 1287
rect 5233 1253 5247 1267
rect 5253 1253 5267 1267
rect 5193 1173 5207 1187
rect 5153 913 5167 927
rect 5153 693 5167 707
rect 5213 1113 5227 1127
rect 5273 1053 5287 1067
rect 5213 893 5227 907
rect 5273 873 5287 887
rect 5233 833 5247 847
rect 5333 1253 5347 1267
rect 5313 1033 5327 1047
rect 5213 353 5227 367
rect 5293 653 5307 667
rect 5273 333 5287 347
rect 5133 173 5147 187
rect 5153 173 5167 187
rect 4833 113 4847 127
rect 4673 13 4687 27
rect 4753 13 4767 27
rect 4793 13 4807 27
rect 4833 13 4847 27
rect 5393 1593 5407 1607
rect 5533 2033 5547 2047
rect 5673 2073 5687 2087
rect 5593 1833 5607 1847
rect 5653 2053 5667 2067
rect 5693 2013 5707 2027
rect 5633 1833 5647 1847
rect 5593 1813 5607 1827
rect 5613 1813 5627 1827
rect 5553 1793 5567 1807
rect 5673 1813 5687 1827
rect 5473 1773 5487 1787
rect 5493 1773 5507 1787
rect 5533 1773 5547 1787
rect 5573 1773 5587 1787
rect 5453 1753 5467 1767
rect 5573 1673 5587 1687
rect 5533 1633 5547 1647
rect 5533 1593 5547 1607
rect 5633 1773 5647 1787
rect 5613 1653 5627 1667
rect 5693 1793 5707 1807
rect 5693 1753 5707 1767
rect 5733 2713 5747 2727
rect 5733 2593 5747 2607
rect 5773 2593 5787 2607
rect 5773 2553 5787 2567
rect 5753 2533 5767 2547
rect 5793 2533 5807 2547
rect 5773 2473 5787 2487
rect 5733 2453 5747 2467
rect 5733 2313 5747 2327
rect 5733 2273 5747 2287
rect 5813 2313 5827 2327
rect 5733 2253 5747 2267
rect 5753 2233 5767 2247
rect 5733 1833 5747 1847
rect 5713 1733 5727 1747
rect 5753 1813 5767 1827
rect 5793 1813 5807 1827
rect 5833 2293 5847 2307
rect 5893 3613 5907 3627
rect 5873 3233 5887 3247
rect 5893 3193 5907 3207
rect 5873 2873 5887 2887
rect 5853 2253 5867 2267
rect 5833 2213 5847 2227
rect 5833 2193 5847 2207
rect 5833 2073 5847 2087
rect 6013 3693 6027 3707
rect 5973 3533 5987 3547
rect 5933 3513 5947 3527
rect 5953 3493 5967 3507
rect 6113 4893 6127 4907
rect 6153 5073 6167 5087
rect 6113 4833 6127 4847
rect 6133 4833 6147 4847
rect 6093 4733 6107 4747
rect 6093 4693 6107 4707
rect 6133 4693 6147 4707
rect 6053 4633 6067 4647
rect 6073 4513 6087 4527
rect 6113 4513 6127 4527
rect 6093 4473 6107 4487
rect 6133 4473 6147 4487
rect 6113 4433 6127 4447
rect 6133 4433 6147 4447
rect 6153 4413 6167 4427
rect 6273 6273 6287 6287
rect 6253 6133 6267 6147
rect 6273 6093 6287 6107
rect 6253 6073 6267 6087
rect 6233 5753 6247 5767
rect 6233 5653 6247 5667
rect 6273 6053 6287 6067
rect 6413 6713 6427 6727
rect 6393 6693 6407 6707
rect 6333 6633 6347 6647
rect 6393 6573 6407 6587
rect 6373 6553 6387 6567
rect 6353 6533 6367 6547
rect 6513 7073 6527 7087
rect 6573 7033 6587 7047
rect 6553 6993 6567 7007
rect 6513 6933 6527 6947
rect 6533 6933 6547 6947
rect 6453 6813 6467 6827
rect 6453 6693 6467 6707
rect 6433 6553 6447 6567
rect 6413 6533 6427 6547
rect 6393 6493 6407 6507
rect 6433 6493 6447 6507
rect 6433 6393 6447 6407
rect 6373 6373 6387 6387
rect 6353 6353 6367 6367
rect 6333 6073 6347 6087
rect 6313 6053 6327 6067
rect 6293 5973 6307 5987
rect 6533 6913 6547 6927
rect 6553 6913 6567 6927
rect 6513 6813 6527 6827
rect 6573 6873 6587 6887
rect 6573 6833 6587 6847
rect 6553 6793 6567 6807
rect 6533 6693 6547 6707
rect 6513 6573 6527 6587
rect 6553 6573 6567 6587
rect 6513 6553 6527 6567
rect 6473 6433 6487 6447
rect 6493 6393 6507 6407
rect 6453 6353 6467 6367
rect 6393 6293 6407 6307
rect 6433 6293 6447 6307
rect 6413 6193 6427 6207
rect 6433 6173 6447 6187
rect 6393 6153 6407 6167
rect 6413 6153 6427 6167
rect 6473 6153 6487 6167
rect 6433 6113 6447 6127
rect 6473 6113 6487 6127
rect 6433 6093 6447 6107
rect 6413 5993 6427 6007
rect 6373 5933 6387 5947
rect 6313 5913 6327 5927
rect 6353 5913 6367 5927
rect 6293 5893 6307 5907
rect 6333 5833 6347 5847
rect 6413 5873 6427 5887
rect 6373 5733 6387 5747
rect 6333 5653 6347 5667
rect 6293 5633 6307 5647
rect 6233 5593 6247 5607
rect 6253 5593 6267 5607
rect 6273 5593 6287 5607
rect 6213 5433 6227 5447
rect 6333 5593 6347 5607
rect 6313 5513 6327 5527
rect 6273 5473 6287 5487
rect 6313 5413 6327 5427
rect 6253 5393 6267 5407
rect 6273 5153 6287 5167
rect 6253 5133 6267 5147
rect 6233 4933 6247 4947
rect 6393 5593 6407 5607
rect 6353 5533 6367 5547
rect 6353 5513 6367 5527
rect 6373 5433 6387 5447
rect 6373 5393 6387 5407
rect 6353 5213 6367 5227
rect 6473 6033 6487 6047
rect 6453 5993 6467 6007
rect 6453 5873 6467 5887
rect 6613 7073 6627 7087
rect 6713 7373 6727 7387
rect 6713 7213 6727 7227
rect 6693 7173 6707 7187
rect 6673 7073 6687 7087
rect 6693 7033 6707 7047
rect 6653 6973 6667 6987
rect 6713 6973 6727 6987
rect 6713 6893 6727 6907
rect 6693 6873 6707 6887
rect 6813 8033 6827 8047
rect 6793 8013 6807 8027
rect 6833 7973 6847 7987
rect 6853 7793 6867 7807
rect 6813 7753 6827 7767
rect 6793 7433 6807 7447
rect 6753 7373 6767 7387
rect 6633 6753 6647 6767
rect 6633 6693 6647 6707
rect 6633 6673 6647 6687
rect 6613 6553 6627 6567
rect 6593 6533 6607 6547
rect 6553 6513 6567 6527
rect 6613 6413 6627 6427
rect 6553 6333 6567 6347
rect 6593 6333 6607 6347
rect 6693 6773 6707 6787
rect 6673 6753 6687 6767
rect 6653 6613 6667 6627
rect 6673 6593 6687 6607
rect 6653 6573 6667 6587
rect 6653 6433 6667 6447
rect 6593 6273 6607 6287
rect 6613 6273 6627 6287
rect 6553 6173 6567 6187
rect 6593 6173 6607 6187
rect 6513 6093 6527 6107
rect 6533 6033 6547 6047
rect 6713 6693 6727 6707
rect 6773 7273 6787 7287
rect 6773 7213 6787 7227
rect 6773 6913 6787 6927
rect 6773 6893 6787 6907
rect 6953 8433 6967 8447
rect 6953 8393 6967 8407
rect 6913 8333 6927 8347
rect 6933 8333 6947 8347
rect 7033 9473 7047 9487
rect 7033 9373 7047 9387
rect 7073 9273 7087 9287
rect 7093 9273 7107 9287
rect 7073 9073 7087 9087
rect 6993 9013 7007 9027
rect 7033 8993 7047 9007
rect 7073 8953 7087 8967
rect 7053 8913 7067 8927
rect 7033 8813 7047 8827
rect 6993 8753 7007 8767
rect 7013 8693 7027 8707
rect 7153 9913 7167 9927
rect 7233 10273 7247 10287
rect 7193 10253 7207 10267
rect 7213 10233 7227 10247
rect 7193 9813 7207 9827
rect 7173 9793 7187 9807
rect 7173 9713 7187 9727
rect 7173 9653 7187 9667
rect 7213 9653 7227 9667
rect 7213 9593 7227 9607
rect 7153 9473 7167 9487
rect 7193 9473 7207 9487
rect 7133 9433 7147 9447
rect 7133 9373 7147 9387
rect 7173 9373 7187 9387
rect 7173 9253 7187 9267
rect 7273 10253 7287 10267
rect 7353 10413 7367 10427
rect 7493 11853 7507 11867
rect 7653 11893 7667 11907
rect 7513 11753 7527 11767
rect 7473 11693 7487 11707
rect 7573 11693 7587 11707
rect 7513 11533 7527 11547
rect 7493 11433 7507 11447
rect 7473 10813 7487 10827
rect 7473 10553 7487 10567
rect 7453 10393 7467 10407
rect 7353 10353 7367 10367
rect 7313 10333 7327 10347
rect 7333 10313 7347 10327
rect 7453 10313 7467 10327
rect 7573 11413 7587 11427
rect 7533 11393 7547 11407
rect 7573 11393 7587 11407
rect 7553 11373 7567 11387
rect 7593 11373 7607 11387
rect 7553 11213 7567 11227
rect 7533 11193 7547 11207
rect 7693 11853 7707 11867
rect 8133 11893 8147 11907
rect 7913 11873 7927 11887
rect 7953 11873 7967 11887
rect 7713 11833 7727 11847
rect 7713 11813 7727 11827
rect 7893 11793 7907 11807
rect 7753 11713 7767 11727
rect 7693 11693 7707 11707
rect 7873 11693 7887 11707
rect 7933 11753 7947 11767
rect 8073 11853 8087 11867
rect 8253 11893 8267 11907
rect 8233 11873 8247 11887
rect 8273 11873 8287 11887
rect 8093 11813 8107 11827
rect 8133 11773 8147 11787
rect 8093 11753 8107 11767
rect 8053 11693 8067 11707
rect 7673 11393 7687 11407
rect 7953 11673 7967 11687
rect 8633 11893 8647 11907
rect 8693 11893 8707 11907
rect 8313 11873 8327 11887
rect 8453 11873 8467 11887
rect 8673 11873 8687 11887
rect 8313 11773 8327 11787
rect 8133 11693 8147 11707
rect 8213 11693 8227 11707
rect 8233 11693 8247 11707
rect 8273 11693 8287 11707
rect 8293 11693 8307 11707
rect 8073 11613 8087 11627
rect 7833 11453 7847 11467
rect 8113 11433 8127 11447
rect 7833 11413 7847 11427
rect 7913 11413 7927 11427
rect 7953 11413 7967 11427
rect 8033 11413 8047 11427
rect 7893 11393 7907 11407
rect 7913 11393 7927 11407
rect 7933 11393 7947 11407
rect 7713 11373 7727 11387
rect 7733 11373 7747 11387
rect 7593 11073 7607 11087
rect 7633 11033 7647 11047
rect 7553 10933 7567 10947
rect 7513 10893 7527 10907
rect 7573 10773 7587 10787
rect 7553 10693 7567 10707
rect 7513 10453 7527 10467
rect 7653 10893 7667 10907
rect 7693 11153 7707 11167
rect 7753 11353 7767 11367
rect 7833 11373 7847 11387
rect 7933 11353 7947 11367
rect 7913 11293 7927 11307
rect 7773 11273 7787 11287
rect 7893 11233 7907 11247
rect 7973 11313 7987 11327
rect 8133 11393 8147 11407
rect 8173 11393 8187 11407
rect 8113 11373 8127 11387
rect 8153 11373 8167 11387
rect 8353 11733 8367 11747
rect 8273 11653 8287 11667
rect 8253 11633 8267 11647
rect 8233 11613 8247 11627
rect 8233 11413 8247 11427
rect 8193 11313 8207 11327
rect 8193 11293 8207 11307
rect 8253 11273 8267 11287
rect 8033 11253 8047 11267
rect 8113 11213 8127 11227
rect 8153 11193 8167 11207
rect 7913 11153 7927 11167
rect 7733 11073 7747 11087
rect 7773 11073 7787 11087
rect 7713 11053 7727 11067
rect 7933 11053 7947 11067
rect 7913 10913 7927 10927
rect 7773 10873 7787 10887
rect 7673 10853 7687 10867
rect 7773 10853 7787 10867
rect 7733 10773 7747 10787
rect 7633 10713 7647 10727
rect 7673 10713 7687 10727
rect 7593 10693 7607 10707
rect 7673 10653 7687 10667
rect 7613 10633 7627 10647
rect 7593 10453 7607 10467
rect 7533 10413 7547 10427
rect 7573 10393 7587 10407
rect 7493 10273 7507 10287
rect 7513 10253 7527 10267
rect 7313 10213 7327 10227
rect 7293 9953 7307 9967
rect 7273 9913 7287 9927
rect 7453 10193 7467 10207
rect 7453 10113 7467 10127
rect 7333 9953 7347 9967
rect 7413 9953 7427 9967
rect 7333 9933 7347 9947
rect 7253 9853 7267 9867
rect 7153 9233 7167 9247
rect 7133 8893 7147 8907
rect 7113 8533 7127 8547
rect 7033 8293 7047 8307
rect 6973 8233 6987 8247
rect 7013 8233 7027 8247
rect 6933 8193 6947 8207
rect 6953 8013 6967 8027
rect 6933 7993 6947 8007
rect 6973 7993 6987 8007
rect 6993 7993 7007 8007
rect 7013 7933 7027 7947
rect 7013 7893 7027 7907
rect 6913 7853 6927 7867
rect 6993 7853 7007 7867
rect 6893 7813 6907 7827
rect 6933 7813 6947 7827
rect 6893 7793 6907 7807
rect 6873 7713 6887 7727
rect 6833 7553 6847 7567
rect 6873 7553 6887 7567
rect 6853 7473 6867 7487
rect 6873 7453 6887 7467
rect 6993 7793 7007 7807
rect 6973 7773 6987 7787
rect 6993 7753 7007 7767
rect 6973 7673 6987 7687
rect 6953 7453 6967 7467
rect 6893 7353 6907 7367
rect 6913 7353 6927 7367
rect 7053 8273 7067 8287
rect 7033 7653 7047 7667
rect 7013 7593 7027 7607
rect 7113 8453 7127 8467
rect 7133 8353 7147 8367
rect 7093 8313 7107 8327
rect 7113 8273 7127 8287
rect 7113 8213 7127 8227
rect 7133 8193 7147 8207
rect 7233 9233 7247 9247
rect 7193 9213 7207 9227
rect 7273 9793 7287 9807
rect 7273 9513 7287 9527
rect 7273 9393 7287 9407
rect 7273 9153 7287 9167
rect 7253 9053 7267 9067
rect 7173 9033 7187 9047
rect 7253 9033 7267 9047
rect 7233 8973 7247 8987
rect 7213 8953 7227 8967
rect 7193 8833 7207 8847
rect 7193 8793 7207 8807
rect 7213 8793 7227 8807
rect 7333 9913 7347 9927
rect 7313 9793 7327 9807
rect 7393 9713 7407 9727
rect 7333 9553 7347 9567
rect 7333 9513 7347 9527
rect 7433 9913 7447 9927
rect 7413 9573 7427 9587
rect 7353 9453 7367 9467
rect 7333 9433 7347 9447
rect 7313 9193 7327 9207
rect 7313 9053 7327 9067
rect 7293 9013 7307 9027
rect 7273 8833 7287 8847
rect 7273 8793 7287 8807
rect 7193 8633 7207 8647
rect 7373 9373 7387 9387
rect 7413 9273 7427 9287
rect 7353 9253 7367 9267
rect 7433 9193 7447 9207
rect 7473 9933 7487 9947
rect 7493 9873 7507 9887
rect 7513 9793 7527 9807
rect 7493 9753 7507 9767
rect 7593 10373 7607 10387
rect 7593 9973 7607 9987
rect 7553 9773 7567 9787
rect 7573 9773 7587 9787
rect 7573 9733 7587 9747
rect 7533 9693 7547 9707
rect 7493 9673 7507 9687
rect 7493 9633 7507 9647
rect 7513 9633 7527 9647
rect 7473 9493 7487 9507
rect 7473 9473 7487 9487
rect 7473 9333 7487 9347
rect 7473 9313 7487 9327
rect 7453 9133 7467 9147
rect 7453 9113 7467 9127
rect 7553 9493 7567 9507
rect 7533 9473 7547 9487
rect 7593 9473 7607 9487
rect 7673 10493 7687 10507
rect 7713 10433 7727 10447
rect 7633 10413 7647 10427
rect 7733 10413 7747 10427
rect 7673 10393 7687 10407
rect 7733 10393 7747 10407
rect 7693 10373 7707 10387
rect 7693 10253 7707 10267
rect 7713 10013 7727 10027
rect 7653 9973 7667 9987
rect 7673 9953 7687 9967
rect 7693 9933 7707 9947
rect 7653 9893 7667 9907
rect 7653 9873 7667 9887
rect 7633 9793 7647 9807
rect 7573 9453 7587 9467
rect 7613 9453 7627 9467
rect 7553 9433 7567 9447
rect 7653 9753 7667 9767
rect 7713 9753 7727 9767
rect 7633 9353 7647 9367
rect 7593 9313 7607 9327
rect 7513 9293 7527 9307
rect 7573 9293 7587 9307
rect 7553 9273 7567 9287
rect 7613 9273 7627 9287
rect 7493 9253 7507 9267
rect 7593 9253 7607 9267
rect 7533 9233 7547 9247
rect 7393 9053 7407 9067
rect 7473 9053 7487 9067
rect 7413 8993 7427 9007
rect 7453 8993 7467 9007
rect 7393 8973 7407 8987
rect 7373 8893 7387 8907
rect 7373 8873 7387 8887
rect 7333 8833 7347 8847
rect 7433 8853 7447 8867
rect 7233 8573 7247 8587
rect 7193 8493 7207 8507
rect 7173 8213 7187 8227
rect 7193 8113 7207 8127
rect 7193 8093 7207 8107
rect 7153 8073 7167 8087
rect 7133 7993 7147 8007
rect 7153 7953 7167 7967
rect 7213 8013 7227 8027
rect 7193 7993 7207 8007
rect 7173 7913 7187 7927
rect 7153 7833 7167 7847
rect 7093 7793 7107 7807
rect 7093 7733 7107 7747
rect 7073 7673 7087 7687
rect 7013 7553 7027 7567
rect 7053 7553 7067 7567
rect 7073 7533 7087 7547
rect 6993 7373 7007 7387
rect 6973 7353 6987 7367
rect 6873 7333 6887 7347
rect 6873 7093 6887 7107
rect 6813 7053 6827 7067
rect 6833 7053 6847 7067
rect 6773 6793 6787 6807
rect 6773 6693 6787 6707
rect 6753 6613 6767 6627
rect 6733 6593 6747 6607
rect 6673 6413 6687 6427
rect 6693 6393 6707 6407
rect 6733 6533 6747 6547
rect 6793 6573 6807 6587
rect 6833 7013 6847 7027
rect 6933 7333 6947 7347
rect 6933 7313 6947 7327
rect 6913 7093 6927 7107
rect 6913 7033 6927 7047
rect 6913 6913 6927 6927
rect 6833 6873 6847 6887
rect 6853 6873 6867 6887
rect 6813 6553 6827 6567
rect 6773 6533 6787 6547
rect 6753 6513 6767 6527
rect 6733 6393 6747 6407
rect 6813 6493 6827 6507
rect 6793 6393 6807 6407
rect 6713 6373 6727 6387
rect 6813 6373 6827 6387
rect 6813 6333 6827 6347
rect 7033 7193 7047 7207
rect 7033 7113 7047 7127
rect 7013 7073 7027 7087
rect 7033 7033 7047 7047
rect 7033 6973 7047 6987
rect 7013 6953 7027 6967
rect 6893 6813 6907 6827
rect 6893 6713 6907 6727
rect 6953 6713 6967 6727
rect 6953 6673 6967 6687
rect 6993 6913 7007 6927
rect 6933 6633 6947 6647
rect 6973 6633 6987 6647
rect 6953 6613 6967 6627
rect 6853 6433 6867 6447
rect 6853 6413 6867 6427
rect 6873 6413 6887 6427
rect 6873 6353 6887 6367
rect 6853 6333 6867 6347
rect 6873 6313 6887 6327
rect 6753 6293 6767 6307
rect 6833 6293 6847 6307
rect 6693 6253 6707 6267
rect 6733 6253 6747 6267
rect 6813 6253 6827 6267
rect 6653 6113 6667 6127
rect 6613 6093 6627 6107
rect 6573 6073 6587 6087
rect 6613 6073 6627 6087
rect 6493 5993 6507 6007
rect 6553 5993 6567 6007
rect 6533 5973 6547 5987
rect 6493 5913 6507 5927
rect 6513 5913 6527 5927
rect 6593 5933 6607 5947
rect 6573 5913 6587 5927
rect 6513 5853 6527 5867
rect 6493 5813 6507 5827
rect 6473 5633 6487 5647
rect 6453 5553 6467 5567
rect 6493 5533 6507 5547
rect 6433 5493 6447 5507
rect 6433 5453 6447 5467
rect 6473 5433 6487 5447
rect 6413 5413 6427 5427
rect 6353 5133 6367 5147
rect 6353 4973 6367 4987
rect 6333 4913 6347 4927
rect 6293 4853 6307 4867
rect 6273 4813 6287 4827
rect 6253 4773 6267 4787
rect 6213 4693 6227 4707
rect 6193 4533 6207 4547
rect 6333 4713 6347 4727
rect 6293 4693 6307 4707
rect 6313 4553 6327 4567
rect 6233 4493 6247 4507
rect 6253 4433 6267 4447
rect 6213 4413 6227 4427
rect 6173 4273 6187 4287
rect 6133 4253 6147 4267
rect 6173 4253 6187 4267
rect 6113 4213 6127 4227
rect 6173 4213 6187 4227
rect 6153 4193 6167 4207
rect 6113 4173 6127 4187
rect 6053 4033 6067 4047
rect 6093 4013 6107 4027
rect 6073 3973 6087 3987
rect 6193 4093 6207 4107
rect 6093 3913 6107 3927
rect 6073 3573 6087 3587
rect 6033 3513 6047 3527
rect 6053 3513 6067 3527
rect 6113 3693 6127 3707
rect 6173 3693 6187 3707
rect 6153 3673 6167 3687
rect 6133 3573 6147 3587
rect 6093 3553 6107 3567
rect 6073 3493 6087 3507
rect 6053 3473 6067 3487
rect 6053 3253 6067 3267
rect 5933 3053 5947 3067
rect 5953 2973 5967 2987
rect 5913 2913 5927 2927
rect 6033 2813 6047 2827
rect 5973 2793 5987 2807
rect 5913 2753 5927 2767
rect 5953 2733 5967 2747
rect 5993 2733 6007 2747
rect 6033 2733 6047 2747
rect 5933 2693 5947 2707
rect 5913 2673 5927 2687
rect 5933 2653 5947 2667
rect 5893 2513 5907 2527
rect 6033 2633 6047 2647
rect 5953 2613 5967 2627
rect 5993 2553 6007 2567
rect 6013 2533 6027 2547
rect 6073 3213 6087 3227
rect 6153 3533 6167 3547
rect 6113 3513 6127 3527
rect 5973 2313 5987 2327
rect 5973 2273 5987 2287
rect 5913 2253 5927 2267
rect 5953 2113 5967 2127
rect 5953 2093 5967 2107
rect 5833 1793 5847 1807
rect 5733 1673 5747 1687
rect 5733 1653 5747 1667
rect 5693 1613 5707 1627
rect 5673 1593 5687 1607
rect 5793 1593 5807 1607
rect 5473 1573 5487 1587
rect 5433 1313 5447 1327
rect 5393 1293 5407 1307
rect 5373 1133 5387 1147
rect 5413 1273 5427 1287
rect 5433 1133 5447 1147
rect 5393 1113 5407 1127
rect 5373 1093 5387 1107
rect 5433 1033 5447 1047
rect 5493 1333 5507 1347
rect 5573 1293 5587 1307
rect 5613 1293 5627 1307
rect 5713 1573 5727 1587
rect 5713 1193 5727 1207
rect 5673 1133 5687 1147
rect 5633 1113 5647 1127
rect 5753 1113 5767 1127
rect 5553 1073 5567 1087
rect 5453 933 5467 947
rect 5473 853 5487 867
rect 5393 673 5407 687
rect 5413 653 5427 667
rect 5713 873 5727 887
rect 5793 1553 5807 1567
rect 5833 1453 5847 1467
rect 5813 1393 5827 1407
rect 5933 2053 5947 2067
rect 5893 2033 5907 2047
rect 5913 2033 5927 2047
rect 5873 1373 5887 1387
rect 5853 1353 5867 1367
rect 5873 1313 5887 1327
rect 5853 1293 5867 1307
rect 5813 1273 5827 1287
rect 5913 1593 5927 1607
rect 6053 2313 6067 2327
rect 6133 3053 6147 3067
rect 6113 2853 6127 2867
rect 6253 4373 6267 4387
rect 6233 4233 6247 4247
rect 6213 3973 6227 3987
rect 6233 3653 6247 3667
rect 6233 3593 6247 3607
rect 6193 2833 6207 2847
rect 6133 2753 6147 2767
rect 6173 2753 6187 2767
rect 6113 2733 6127 2747
rect 6153 2673 6167 2687
rect 6173 2613 6187 2627
rect 6353 4473 6367 4487
rect 6493 5413 6507 5427
rect 6573 5833 6587 5847
rect 6553 5713 6567 5727
rect 6553 5553 6567 5567
rect 6473 5393 6487 5407
rect 6533 5393 6547 5407
rect 6433 5173 6447 5187
rect 6513 5173 6527 5187
rect 6433 5013 6447 5027
rect 6413 4893 6427 4907
rect 6393 4633 6407 4647
rect 6393 4513 6407 4527
rect 6413 4433 6427 4447
rect 6393 4393 6407 4407
rect 6373 4293 6387 4307
rect 6333 4213 6347 4227
rect 6493 5033 6507 5047
rect 6453 4993 6467 5007
rect 6633 6033 6647 6047
rect 6613 5693 6627 5707
rect 6693 6093 6707 6107
rect 6673 6033 6687 6047
rect 6673 5993 6687 6007
rect 6653 5833 6667 5847
rect 6853 6153 6867 6167
rect 6733 6073 6747 6087
rect 6833 6073 6847 6087
rect 6713 6033 6727 6047
rect 6733 6033 6747 6047
rect 6733 5953 6747 5967
rect 6753 5953 6767 5967
rect 6793 5933 6807 5947
rect 6813 5933 6827 5947
rect 6693 5913 6707 5927
rect 6713 5893 6727 5907
rect 6733 5893 6747 5907
rect 6773 5893 6787 5907
rect 6693 5613 6707 5627
rect 6633 5573 6647 5587
rect 6673 5573 6687 5587
rect 6653 5493 6667 5507
rect 6613 5453 6627 5467
rect 6573 5253 6587 5267
rect 6633 5373 6647 5387
rect 6693 5393 6707 5407
rect 6673 5353 6687 5367
rect 6813 5853 6827 5867
rect 6853 6013 6867 6027
rect 6833 5833 6847 5847
rect 6853 5773 6867 5787
rect 6793 5693 6807 5707
rect 6753 5653 6767 5667
rect 6673 5253 6687 5267
rect 6713 5253 6727 5267
rect 6593 5173 6607 5187
rect 6633 5153 6647 5167
rect 6713 5193 6727 5207
rect 6653 5133 6667 5147
rect 6933 6593 6947 6607
rect 6973 6573 6987 6587
rect 6933 6553 6947 6567
rect 6913 6433 6927 6447
rect 6953 6433 6967 6447
rect 6913 6393 6927 6407
rect 6973 6393 6987 6407
rect 6953 6333 6967 6347
rect 6913 6233 6927 6247
rect 6893 6073 6907 6087
rect 6893 5993 6907 6007
rect 6813 5633 6827 5647
rect 6813 5613 6827 5627
rect 6873 5613 6887 5627
rect 6933 6133 6947 6147
rect 6993 6253 7007 6267
rect 7033 6913 7047 6927
rect 7033 6673 7047 6687
rect 7073 7453 7087 7467
rect 7073 7353 7087 7367
rect 7173 7813 7187 7827
rect 7133 7653 7147 7667
rect 7113 7493 7127 7507
rect 7093 7313 7107 7327
rect 7073 7193 7087 7207
rect 7213 7833 7227 7847
rect 7213 7733 7227 7747
rect 7253 8493 7267 8507
rect 7253 8453 7267 8467
rect 7253 8393 7267 8407
rect 7273 8373 7287 8387
rect 7273 8273 7287 8287
rect 7313 8313 7327 8327
rect 7293 8133 7307 8147
rect 7273 7733 7287 7747
rect 7193 7633 7207 7647
rect 7233 7633 7247 7647
rect 7213 7553 7227 7567
rect 7253 7553 7267 7567
rect 7193 7453 7207 7467
rect 7173 7413 7187 7427
rect 7133 7393 7147 7407
rect 7173 7393 7187 7407
rect 7233 7393 7247 7407
rect 7153 7333 7167 7347
rect 7133 7293 7147 7307
rect 7113 7093 7127 7107
rect 7093 7033 7107 7047
rect 7233 7253 7247 7267
rect 7373 8693 7387 8707
rect 7453 8793 7467 8807
rect 7393 8593 7407 8607
rect 7493 8973 7507 8987
rect 7513 8893 7527 8907
rect 7493 8833 7507 8847
rect 7413 8533 7427 8547
rect 7473 8533 7487 8547
rect 7393 8513 7407 8527
rect 7393 8373 7407 8387
rect 7373 8353 7387 8367
rect 7353 8313 7367 8327
rect 7373 8273 7387 8287
rect 7373 8253 7387 8267
rect 7433 8493 7447 8507
rect 7473 8493 7487 8507
rect 7453 8473 7467 8487
rect 7633 9113 7647 9127
rect 7553 9053 7567 9067
rect 7613 9013 7627 9027
rect 7573 8993 7587 9007
rect 7593 8973 7607 8987
rect 7633 8973 7647 8987
rect 7593 8953 7607 8967
rect 7553 8873 7567 8887
rect 7533 8853 7547 8867
rect 7673 9653 7687 9667
rect 7753 10253 7767 10267
rect 7753 10193 7767 10207
rect 7753 9953 7767 9967
rect 7753 9653 7767 9667
rect 7733 9493 7747 9507
rect 7713 9473 7727 9487
rect 7753 9473 7767 9487
rect 7693 9433 7707 9447
rect 7673 9253 7687 9267
rect 7653 8893 7667 8907
rect 7613 8853 7627 8867
rect 7633 8853 7647 8867
rect 7593 8833 7607 8847
rect 7573 8793 7587 8807
rect 7553 8573 7567 8587
rect 7513 8473 7527 8487
rect 7433 8453 7447 8467
rect 7493 8453 7507 8467
rect 7413 8333 7427 8347
rect 7413 8233 7427 8247
rect 7393 8133 7407 8147
rect 7353 7993 7367 8007
rect 7393 7993 7407 8007
rect 7333 7913 7347 7927
rect 7473 8313 7487 8327
rect 7473 8293 7487 8307
rect 7453 8253 7467 8267
rect 7493 8233 7507 8247
rect 7653 8833 7667 8847
rect 7653 8793 7667 8807
rect 7673 8773 7687 8787
rect 7753 9433 7767 9447
rect 7853 10793 7867 10807
rect 7793 10693 7807 10707
rect 7813 10693 7827 10707
rect 7713 9293 7727 9307
rect 7753 9293 7767 9307
rect 7773 9293 7787 9307
rect 7733 9213 7747 9227
rect 7753 9113 7767 9127
rect 7753 9013 7767 9027
rect 7713 8893 7727 8907
rect 7653 8653 7667 8667
rect 7693 8653 7707 8667
rect 7573 8513 7587 8527
rect 7613 8513 7627 8527
rect 7693 8593 7707 8607
rect 7613 8473 7627 8487
rect 7573 8413 7587 8427
rect 7573 8253 7587 8267
rect 7453 7993 7467 8007
rect 7533 7993 7547 8007
rect 7493 7953 7507 7967
rect 7573 7953 7587 7967
rect 7513 7893 7527 7907
rect 7493 7873 7507 7887
rect 7333 7833 7347 7847
rect 7373 7833 7387 7847
rect 7433 7833 7447 7847
rect 7533 7873 7547 7887
rect 7593 7873 7607 7887
rect 7553 7833 7567 7847
rect 7313 7813 7327 7827
rect 7353 7813 7367 7827
rect 7493 7813 7507 7827
rect 7593 7813 7607 7827
rect 7373 7793 7387 7807
rect 7513 7793 7527 7807
rect 7313 7633 7327 7647
rect 7293 7513 7307 7527
rect 7293 7453 7307 7467
rect 7353 7593 7367 7607
rect 7313 7333 7327 7347
rect 7493 7613 7507 7627
rect 7413 7573 7427 7587
rect 7433 7553 7447 7567
rect 7433 7433 7447 7447
rect 7433 7413 7447 7427
rect 7473 7413 7487 7427
rect 7373 7373 7387 7387
rect 7373 7333 7387 7347
rect 7333 7313 7347 7327
rect 7273 7293 7287 7307
rect 7353 7293 7367 7307
rect 7413 7293 7427 7307
rect 7253 7213 7267 7227
rect 7153 7073 7167 7087
rect 7333 7033 7347 7047
rect 7333 7013 7347 7027
rect 7193 6993 7207 7007
rect 7133 6933 7147 6947
rect 7073 6853 7087 6867
rect 7053 6653 7067 6667
rect 7053 6553 7067 6567
rect 7053 6233 7067 6247
rect 7033 6213 7047 6227
rect 7033 6153 7047 6167
rect 7013 6133 7027 6147
rect 7113 6813 7127 6827
rect 7113 6713 7127 6727
rect 7153 6653 7167 6667
rect 7113 6593 7127 6607
rect 7293 6973 7307 6987
rect 7213 6953 7227 6967
rect 7253 6933 7267 6947
rect 7213 6893 7227 6907
rect 7233 6893 7247 6907
rect 7213 6793 7227 6807
rect 7193 6573 7207 6587
rect 7313 6873 7327 6887
rect 7273 6853 7287 6867
rect 7273 6833 7287 6847
rect 7273 6793 7287 6807
rect 7333 6753 7347 6767
rect 7273 6733 7287 6747
rect 7233 6693 7247 6707
rect 7133 6413 7147 6427
rect 7213 6413 7227 6427
rect 7173 6393 7187 6407
rect 7113 6373 7127 6387
rect 7153 6313 7167 6327
rect 7133 6273 7147 6287
rect 6953 6113 6967 6127
rect 6993 6113 7007 6127
rect 7033 6113 7047 6127
rect 7073 6113 7087 6127
rect 6933 6093 6947 6107
rect 6933 5973 6947 5987
rect 6973 6093 6987 6107
rect 7053 6093 7067 6107
rect 7073 6093 7087 6107
rect 7053 6073 7067 6087
rect 7013 6053 7027 6067
rect 7013 6033 7027 6047
rect 6973 6013 6987 6027
rect 6953 5933 6967 5947
rect 7113 6113 7127 6127
rect 7073 5993 7087 6007
rect 7093 5993 7107 6007
rect 7093 5953 7107 5967
rect 6993 5893 7007 5907
rect 7053 5893 7067 5907
rect 7073 5893 7087 5907
rect 6953 5853 6967 5867
rect 7073 5853 7087 5867
rect 6933 5833 6947 5847
rect 6993 5833 7007 5847
rect 6913 5653 6927 5667
rect 6913 5613 6927 5627
rect 6813 5473 6827 5487
rect 6833 5453 6847 5467
rect 6893 5593 6907 5607
rect 6993 5733 7007 5747
rect 6993 5693 7007 5707
rect 6993 5613 7007 5627
rect 6933 5573 6947 5587
rect 6933 5513 6947 5527
rect 6853 5413 6867 5427
rect 6853 5393 6867 5407
rect 6793 5273 6807 5287
rect 6813 5273 6827 5287
rect 6793 5153 6807 5167
rect 6633 5093 6647 5107
rect 6693 5093 6707 5107
rect 6693 5033 6707 5047
rect 6633 5013 6647 5027
rect 6553 4993 6567 5007
rect 6533 4953 6547 4967
rect 6573 4953 6587 4967
rect 6553 4933 6567 4947
rect 6593 4913 6607 4927
rect 6513 4873 6527 4887
rect 6533 4713 6547 4727
rect 6473 4653 6487 4667
rect 6553 4693 6567 4707
rect 6633 4713 6647 4727
rect 6633 4693 6647 4707
rect 6673 4693 6687 4707
rect 6593 4653 6607 4667
rect 6553 4613 6567 4627
rect 6493 4533 6507 4547
rect 6573 4453 6587 4467
rect 6613 4433 6627 4447
rect 6593 4413 6607 4427
rect 6453 4233 6467 4247
rect 6533 4233 6547 4247
rect 6433 4213 6447 4227
rect 6393 4193 6407 4207
rect 6493 4213 6507 4227
rect 6473 4193 6487 4207
rect 6513 4193 6527 4207
rect 6593 4193 6607 4207
rect 6453 4173 6467 4187
rect 6593 4153 6607 4167
rect 6433 4133 6447 4147
rect 6393 4033 6407 4047
rect 6273 3973 6287 3987
rect 6493 4033 6507 4047
rect 6313 3953 6327 3967
rect 6393 3853 6407 3867
rect 6393 3713 6407 3727
rect 6333 3693 6347 3707
rect 6333 3653 6347 3667
rect 6273 3393 6287 3407
rect 6353 3493 6367 3507
rect 6553 3973 6567 3987
rect 6533 3753 6547 3767
rect 6513 3553 6527 3567
rect 6573 3553 6587 3567
rect 6533 3533 6547 3547
rect 6753 4973 6767 4987
rect 6773 4853 6787 4867
rect 6713 4833 6727 4847
rect 6833 5253 6847 5267
rect 6733 4553 6747 4567
rect 6693 4433 6707 4447
rect 6753 4453 6767 4467
rect 6773 4413 6787 4427
rect 6633 4053 6647 4067
rect 6633 4013 6647 4027
rect 6733 4173 6747 4187
rect 6753 4113 6767 4127
rect 6693 4053 6707 4067
rect 6673 4033 6687 4047
rect 6893 5353 6907 5367
rect 7053 5633 7067 5647
rect 7033 5613 7047 5627
rect 7073 5593 7087 5607
rect 7033 5573 7047 5587
rect 7053 5573 7067 5587
rect 7013 5493 7027 5507
rect 6973 5453 6987 5467
rect 7013 5433 7027 5447
rect 6933 5153 6947 5167
rect 6873 5133 6887 5147
rect 6853 5053 6867 5067
rect 6853 4933 6867 4947
rect 6853 4693 6867 4707
rect 6833 4673 6847 4687
rect 6953 5133 6967 5147
rect 6913 5113 6927 5127
rect 6913 4993 6927 5007
rect 6953 4953 6967 4967
rect 6893 4933 6907 4947
rect 6933 4933 6947 4947
rect 6893 4893 6907 4907
rect 6953 4713 6967 4727
rect 6913 4693 6927 4707
rect 6913 4533 6927 4547
rect 6933 4453 6947 4467
rect 6893 4373 6907 4387
rect 6873 4353 6887 4367
rect 6853 4173 6867 4187
rect 6893 4113 6907 4127
rect 6993 5413 7007 5427
rect 6993 5153 7007 5167
rect 6993 5113 7007 5127
rect 6993 4953 7007 4967
rect 7153 6253 7167 6267
rect 7133 6093 7147 6107
rect 7173 6233 7187 6247
rect 7193 6233 7207 6247
rect 7213 6193 7227 6207
rect 7193 6133 7207 6147
rect 7393 6993 7407 7007
rect 7373 6953 7387 6967
rect 7413 6953 7427 6967
rect 7393 6833 7407 6847
rect 7373 6733 7387 6747
rect 7373 6713 7387 6727
rect 7353 6633 7367 6647
rect 7253 6533 7267 6547
rect 7273 6393 7287 6407
rect 7253 6273 7267 6287
rect 7273 6193 7287 6207
rect 7233 6153 7247 6167
rect 7273 6133 7287 6147
rect 7253 6113 7267 6127
rect 7233 6093 7247 6107
rect 7193 6033 7207 6047
rect 7153 5993 7167 6007
rect 7173 5993 7187 6007
rect 7173 5933 7187 5947
rect 7133 5873 7147 5887
rect 7153 5873 7167 5887
rect 7133 5633 7147 5647
rect 7113 5613 7127 5627
rect 7113 5333 7127 5347
rect 7213 5753 7227 5767
rect 7213 5593 7227 5607
rect 7253 6033 7267 6047
rect 7253 5873 7267 5887
rect 7333 6393 7347 6407
rect 7313 6333 7327 6347
rect 7293 5713 7307 5727
rect 7273 5633 7287 5647
rect 7233 5553 7247 5567
rect 7233 5513 7247 5527
rect 7173 5433 7187 5447
rect 7193 5433 7207 5447
rect 7253 5493 7267 5507
rect 7273 5473 7287 5487
rect 7253 5373 7267 5387
rect 7073 5233 7087 5247
rect 7093 5233 7107 5247
rect 7153 5173 7167 5187
rect 7113 5153 7127 5167
rect 7053 5013 7067 5027
rect 7033 4913 7047 4927
rect 7073 4913 7087 4927
rect 6993 4673 7007 4687
rect 7133 5013 7147 5027
rect 7153 4993 7167 5007
rect 7113 4933 7127 4947
rect 7093 4853 7107 4867
rect 6973 4573 6987 4587
rect 7013 4493 7027 4507
rect 6973 4313 6987 4327
rect 6993 4173 7007 4187
rect 6953 4073 6967 4087
rect 6873 4053 6887 4067
rect 6853 4013 6867 4027
rect 6893 4013 6907 4027
rect 6813 3993 6827 4007
rect 7213 5333 7227 5347
rect 7193 4973 7207 4987
rect 7173 4933 7187 4947
rect 7153 4693 7167 4707
rect 7133 4653 7147 4667
rect 7133 4593 7147 4607
rect 7113 4513 7127 4527
rect 7093 4493 7107 4507
rect 7033 4453 7047 4467
rect 7113 4453 7127 4467
rect 7073 4433 7087 4447
rect 7093 4213 7107 4227
rect 7053 4193 7067 4207
rect 7073 4173 7087 4187
rect 7013 4153 7027 4167
rect 7053 4013 7067 4027
rect 7133 4013 7147 4027
rect 7033 3993 7047 4007
rect 7073 3993 7087 4007
rect 6733 3973 6747 3987
rect 6833 3973 6847 3987
rect 6873 3973 6887 3987
rect 6993 3973 7007 3987
rect 6633 3953 6647 3967
rect 7053 3773 7067 3787
rect 7073 3773 7087 3787
rect 6913 3753 6927 3767
rect 6733 3733 6747 3747
rect 6513 3493 6527 3507
rect 6493 3453 6507 3467
rect 6473 3433 6487 3447
rect 6313 3253 6327 3267
rect 6273 3233 6287 3247
rect 6253 3153 6267 3167
rect 6313 3233 6327 3247
rect 6433 3213 6447 3227
rect 6273 3133 6287 3147
rect 6293 3133 6307 3147
rect 6253 3093 6267 3107
rect 6233 2653 6247 2667
rect 6193 2593 6207 2607
rect 6193 2553 6207 2567
rect 6213 2513 6227 2527
rect 6113 2293 6127 2307
rect 6133 2273 6147 2287
rect 6173 2253 6187 2267
rect 6153 2233 6167 2247
rect 6153 2213 6167 2227
rect 6073 2093 6087 2107
rect 6113 2093 6127 2107
rect 6053 2053 6067 2067
rect 6093 2033 6107 2047
rect 5953 1693 5967 1707
rect 6013 1793 6027 1807
rect 5993 1773 6007 1787
rect 6033 1753 6047 1767
rect 5993 1593 6007 1607
rect 5973 1413 5987 1427
rect 5893 1233 5907 1247
rect 5853 1193 5867 1207
rect 5893 1193 5907 1207
rect 5773 853 5787 867
rect 5553 813 5567 827
rect 5613 813 5627 827
rect 5653 813 5667 827
rect 5713 813 5727 827
rect 5753 813 5767 827
rect 5793 813 5807 827
rect 5973 1353 5987 1367
rect 5953 1253 5967 1267
rect 5953 1173 5967 1187
rect 5913 1113 5927 1127
rect 5933 1093 5947 1107
rect 5973 1093 5987 1107
rect 5473 653 5487 667
rect 5353 593 5367 607
rect 5453 513 5467 527
rect 5373 353 5387 367
rect 5413 353 5427 367
rect 5393 333 5407 347
rect 5753 693 5767 707
rect 5533 633 5547 647
rect 5633 633 5647 647
rect 5513 393 5527 407
rect 5473 373 5487 387
rect 5453 213 5467 227
rect 5333 173 5347 187
rect 5293 153 5307 167
rect 5353 133 5367 147
rect 5493 133 5507 147
rect 5613 613 5627 627
rect 5793 633 5807 647
rect 5813 613 5827 627
rect 5593 593 5607 607
rect 5633 593 5647 607
rect 5673 593 5687 607
rect 5733 413 5747 427
rect 5573 373 5587 387
rect 5593 353 5607 367
rect 5633 333 5647 347
rect 5573 173 5587 187
rect 5533 153 5547 167
rect 6133 1673 6147 1687
rect 6113 1573 6127 1587
rect 6233 2153 6247 2167
rect 6493 3153 6507 3167
rect 6473 3053 6487 3067
rect 6293 3033 6307 3047
rect 6333 3033 6347 3047
rect 6453 3033 6467 3047
rect 6473 3033 6487 3047
rect 6333 2773 6347 2787
rect 6393 2753 6407 2767
rect 6453 2753 6467 2767
rect 6333 2733 6347 2747
rect 6373 2733 6387 2747
rect 6433 2733 6447 2747
rect 6413 2613 6427 2627
rect 6353 2573 6367 2587
rect 6393 2553 6407 2567
rect 6413 2553 6427 2567
rect 6453 2673 6467 2687
rect 6553 3513 6567 3527
rect 6733 3613 6747 3627
rect 6873 3613 6887 3627
rect 6713 3513 6727 3527
rect 6613 3493 6627 3507
rect 6673 3313 6687 3327
rect 6593 3233 6607 3247
rect 6633 3233 6647 3247
rect 6693 3193 6707 3207
rect 6653 3173 6667 3187
rect 6793 3393 6807 3407
rect 6713 3113 6727 3127
rect 6693 3073 6707 3087
rect 6653 3053 6667 3067
rect 6633 3033 6647 3047
rect 6713 3053 6727 3067
rect 6673 3013 6687 3027
rect 7093 3613 7107 3627
rect 7033 3473 7047 3487
rect 7073 3473 7087 3487
rect 6933 3273 6947 3287
rect 6873 3253 6887 3267
rect 6833 3213 6847 3227
rect 6813 3193 6827 3207
rect 6853 3193 6867 3207
rect 6813 3173 6827 3187
rect 6793 3013 6807 3027
rect 6853 3033 6867 3047
rect 6653 2913 6667 2927
rect 6553 2773 6567 2787
rect 6613 2733 6627 2747
rect 6533 2713 6547 2727
rect 6573 2713 6587 2727
rect 6473 2553 6487 2567
rect 6373 2493 6387 2507
rect 6433 2493 6447 2507
rect 6513 2393 6527 2407
rect 6573 2693 6587 2707
rect 6613 2573 6627 2587
rect 6593 2533 6607 2547
rect 6573 2373 6587 2387
rect 6313 2293 6327 2307
rect 6353 2293 6367 2307
rect 6513 2293 6527 2307
rect 6533 2293 6547 2307
rect 6333 2273 6347 2287
rect 6373 2233 6387 2247
rect 6293 2213 6307 2227
rect 6533 2253 6547 2267
rect 6273 2153 6287 2167
rect 6513 2153 6527 2167
rect 6253 2093 6267 2107
rect 6313 2093 6327 2107
rect 6393 2093 6407 2107
rect 6513 2093 6527 2107
rect 6273 2073 6287 2087
rect 6253 2033 6267 2047
rect 6293 2033 6307 2047
rect 6233 1873 6247 1887
rect 6273 1873 6287 1887
rect 6233 1853 6247 1867
rect 6193 1813 6207 1827
rect 6173 1773 6187 1787
rect 6193 1753 6207 1767
rect 6193 1713 6207 1727
rect 6013 1433 6027 1447
rect 6053 1433 6067 1447
rect 5993 713 6007 727
rect 6173 1493 6187 1507
rect 6173 1373 6187 1387
rect 6033 1333 6047 1347
rect 6073 1333 6087 1347
rect 6113 1333 6127 1347
rect 6093 1313 6107 1327
rect 6153 1313 6167 1327
rect 6093 1273 6107 1287
rect 6133 1173 6147 1187
rect 6093 1113 6107 1127
rect 6033 813 6047 827
rect 6073 813 6087 827
rect 6053 793 6067 807
rect 6113 773 6127 787
rect 5853 573 5867 587
rect 5933 373 5947 387
rect 5773 353 5787 367
rect 5813 353 5827 367
rect 5973 353 5987 367
rect 6033 633 6047 647
rect 6213 1633 6227 1647
rect 6433 2073 6447 2087
rect 6473 2073 6487 2087
rect 6513 2073 6527 2087
rect 6393 1793 6407 1807
rect 6453 2053 6467 2067
rect 6493 2053 6507 2067
rect 6473 2033 6487 2047
rect 6473 1973 6487 1987
rect 6353 1613 6367 1627
rect 6293 1593 6307 1607
rect 6313 1593 6327 1607
rect 6453 1753 6467 1767
rect 6413 1733 6427 1747
rect 6333 1573 6347 1587
rect 6373 1573 6387 1587
rect 6513 1873 6527 1887
rect 6513 1733 6527 1747
rect 6553 2113 6567 2127
rect 6633 2473 6647 2487
rect 6633 2293 6647 2307
rect 6593 2093 6607 2107
rect 6553 2073 6567 2087
rect 6593 2053 6607 2067
rect 6613 1873 6627 1887
rect 6553 1773 6567 1787
rect 6573 1753 6587 1767
rect 6613 1773 6627 1787
rect 6593 1733 6607 1747
rect 6493 1593 6507 1607
rect 6513 1573 6527 1587
rect 6493 1553 6507 1567
rect 6393 1533 6407 1547
rect 6473 1533 6487 1547
rect 6533 1533 6547 1547
rect 6373 1393 6387 1407
rect 6273 1313 6287 1327
rect 6213 1233 6227 1247
rect 6173 1153 6187 1167
rect 6173 1093 6187 1107
rect 6153 613 6167 627
rect 6053 593 6067 607
rect 6133 553 6147 567
rect 6013 393 6027 407
rect 6013 373 6027 387
rect 5953 333 5967 347
rect 5993 333 6007 347
rect 6373 1293 6387 1307
rect 6373 1253 6387 1267
rect 6253 1233 6267 1247
rect 6353 1213 6367 1227
rect 6333 1193 6347 1207
rect 6273 1133 6287 1147
rect 6233 1113 6247 1127
rect 6293 1113 6307 1127
rect 6313 1093 6327 1107
rect 6353 1093 6367 1107
rect 6293 813 6307 827
rect 6253 793 6267 807
rect 6253 753 6267 767
rect 6273 693 6287 707
rect 6253 613 6267 627
rect 6193 593 6207 607
rect 6233 593 6247 607
rect 6373 653 6387 667
rect 6413 1313 6427 1327
rect 6453 1313 6467 1327
rect 6433 1293 6447 1307
rect 6533 1413 6547 1427
rect 6513 1373 6527 1387
rect 6493 1273 6507 1287
rect 6453 1153 6467 1167
rect 6433 1093 6447 1107
rect 6413 833 6427 847
rect 6453 673 6467 687
rect 6453 653 6467 667
rect 6413 633 6427 647
rect 6393 613 6407 627
rect 6433 573 6447 587
rect 6533 1293 6547 1307
rect 6533 1153 6547 1167
rect 6513 813 6527 827
rect 6493 793 6507 807
rect 6533 633 6547 647
rect 6493 573 6507 587
rect 6473 533 6487 547
rect 6253 333 6267 347
rect 5953 313 5967 327
rect 6013 313 6027 327
rect 5913 253 5927 267
rect 5693 213 5707 227
rect 5873 193 5887 207
rect 5733 153 5747 167
rect 5633 133 5647 147
rect 5713 133 5727 147
rect 5913 173 5927 187
rect 6173 313 6187 327
rect 6113 173 6127 187
rect 5893 133 5907 147
rect 5773 113 5787 127
rect 6113 113 6127 127
rect 6173 153 6187 167
rect 6433 333 6447 347
rect 6473 333 6487 347
rect 6273 293 6287 307
rect 6293 193 6307 207
rect 6533 413 6547 427
rect 6573 1593 6587 1607
rect 6593 1573 6607 1587
rect 6573 1553 6587 1567
rect 6593 1433 6607 1447
rect 6713 2793 6727 2807
rect 6833 2973 6847 2987
rect 6813 2773 6827 2787
rect 6713 2753 6727 2767
rect 6753 2753 6767 2767
rect 6793 2753 6807 2767
rect 6733 2673 6747 2687
rect 6673 2473 6687 2487
rect 6693 2473 6707 2487
rect 6773 2613 6787 2627
rect 6813 2573 6827 2587
rect 6773 2533 6787 2547
rect 6753 2493 6767 2507
rect 6733 2413 6747 2427
rect 6773 2473 6787 2487
rect 6753 2313 6767 2327
rect 6673 2233 6687 2247
rect 6733 2273 6747 2287
rect 6713 2253 6727 2267
rect 6733 2233 6747 2247
rect 6693 2173 6707 2187
rect 6693 2133 6707 2147
rect 6673 2093 6687 2107
rect 6653 2073 6667 2087
rect 6713 2113 6727 2127
rect 6753 2153 6767 2167
rect 6753 2113 6767 2127
rect 6773 2033 6787 2047
rect 6813 2493 6827 2507
rect 6813 2313 6827 2327
rect 6813 2253 6827 2267
rect 6913 2973 6927 2987
rect 6873 2833 6887 2847
rect 6873 2793 6887 2807
rect 7033 3233 7047 3247
rect 6973 2753 6987 2767
rect 6913 2733 6927 2747
rect 6993 2733 7007 2747
rect 6853 2713 6867 2727
rect 6873 2713 6887 2727
rect 6953 2713 6967 2727
rect 6853 2353 6867 2367
rect 6853 2273 6867 2287
rect 6833 2093 6847 2107
rect 6913 2653 6927 2667
rect 6953 2633 6967 2647
rect 6933 2573 6947 2587
rect 6913 2533 6927 2547
rect 7053 3193 7067 3207
rect 7033 3073 7047 3087
rect 7073 3053 7087 3067
rect 7113 3033 7127 3047
rect 7053 3013 7067 3027
rect 7093 2993 7107 3007
rect 7013 2693 7027 2707
rect 6993 2573 7007 2587
rect 7113 2953 7127 2967
rect 7113 2833 7127 2847
rect 7173 4633 7187 4647
rect 7353 6213 7367 6227
rect 7413 6633 7427 6647
rect 7473 7293 7487 7307
rect 7453 7073 7467 7087
rect 7453 7053 7467 7067
rect 7453 6993 7467 7007
rect 7673 8473 7687 8487
rect 7653 8373 7667 8387
rect 7633 8153 7647 8167
rect 7653 8153 7667 8167
rect 7633 8133 7647 8147
rect 7633 7873 7647 7887
rect 7573 7633 7587 7647
rect 7613 7633 7627 7647
rect 7613 7593 7627 7607
rect 7653 7593 7667 7607
rect 7733 8813 7747 8827
rect 7773 8973 7787 8987
rect 7833 10493 7847 10507
rect 7813 10413 7827 10427
rect 7813 10253 7827 10267
rect 7953 10853 7967 10867
rect 7953 10813 7967 10827
rect 8093 11113 8107 11127
rect 8033 10913 8047 10927
rect 8053 10733 8067 10747
rect 8013 10713 8027 10727
rect 8073 10693 8087 10707
rect 8033 10673 8047 10687
rect 7953 10513 7967 10527
rect 7913 10473 7927 10487
rect 7893 10453 7907 10467
rect 7933 10433 7947 10447
rect 7973 10453 7987 10467
rect 7913 10413 7927 10427
rect 7953 10413 7967 10427
rect 7933 10393 7947 10407
rect 7973 10393 7987 10407
rect 7953 10313 7967 10327
rect 7873 10273 7887 10287
rect 7913 10273 7927 10287
rect 7853 10233 7867 10247
rect 7893 10233 7907 10247
rect 7873 10053 7887 10067
rect 7833 10033 7847 10047
rect 7833 9933 7847 9947
rect 7933 10233 7947 10247
rect 7833 9913 7847 9927
rect 7853 9833 7867 9847
rect 8193 11133 8207 11147
rect 8173 10893 8187 10907
rect 8253 10893 8267 10907
rect 8233 10833 8247 10847
rect 8233 10733 8247 10747
rect 8293 11473 8307 11487
rect 8313 11413 8327 11427
rect 8433 11693 8447 11707
rect 8593 11813 8607 11827
rect 8493 11733 8507 11747
rect 8873 11853 8887 11867
rect 8933 11853 8947 11867
rect 8833 11833 8847 11847
rect 8813 11793 8827 11807
rect 8713 11733 8727 11747
rect 8533 11713 8547 11727
rect 8693 11713 8707 11727
rect 8293 11393 8307 11407
rect 8193 10693 8207 10707
rect 8153 10533 8167 10547
rect 8013 10473 8027 10487
rect 8033 10433 8047 10447
rect 8013 10373 8027 10387
rect 7993 10273 8007 10287
rect 8093 10433 8107 10447
rect 8173 10473 8187 10487
rect 8113 10413 8127 10427
rect 8153 10373 8167 10387
rect 8133 10353 8147 10367
rect 8073 10313 8087 10327
rect 8053 10233 8067 10247
rect 8133 10233 8147 10247
rect 7973 10213 7987 10227
rect 8033 10213 8047 10227
rect 8013 10193 8027 10207
rect 8013 10173 8027 10187
rect 8053 10153 8067 10167
rect 8093 10033 8107 10047
rect 8113 10033 8127 10047
rect 8013 10013 8027 10027
rect 7973 9993 7987 10007
rect 7933 9833 7947 9847
rect 7853 9773 7867 9787
rect 7913 9773 7927 9787
rect 7833 9733 7847 9747
rect 7813 9153 7827 9167
rect 7813 9093 7827 9107
rect 7893 9753 7907 9767
rect 7953 9773 7967 9787
rect 7993 9973 8007 9987
rect 8073 9993 8087 10007
rect 8053 9973 8067 9987
rect 8033 9933 8047 9947
rect 7993 9893 8007 9907
rect 8073 9893 8087 9907
rect 8113 9833 8127 9847
rect 8093 9793 8107 9807
rect 7873 9733 7887 9747
rect 7913 9693 7927 9707
rect 7853 9593 7867 9607
rect 7853 9453 7867 9467
rect 7893 9453 7907 9467
rect 7973 9733 7987 9747
rect 7913 9433 7927 9447
rect 7953 9433 7967 9447
rect 7933 9413 7947 9427
rect 7853 9273 7867 9287
rect 7853 9233 7867 9247
rect 7913 9253 7927 9267
rect 7873 9213 7887 9227
rect 7893 9193 7907 9207
rect 7873 9133 7887 9147
rect 7853 8973 7867 8987
rect 7833 8953 7847 8967
rect 7873 8913 7887 8927
rect 7813 8893 7827 8907
rect 7873 8893 7887 8907
rect 7733 8773 7747 8787
rect 7753 8533 7767 8547
rect 7793 8513 7807 8527
rect 7773 8473 7787 8487
rect 7733 8453 7747 8467
rect 7733 8433 7747 8447
rect 7753 8433 7767 8447
rect 7713 8373 7727 8387
rect 7733 8293 7747 8307
rect 7713 8233 7727 8247
rect 7733 8173 7747 8187
rect 7713 8133 7727 8147
rect 7773 8373 7787 8387
rect 7753 8093 7767 8107
rect 7753 8073 7767 8087
rect 7733 8053 7747 8067
rect 7693 8013 7707 8027
rect 7693 7973 7707 7987
rect 7753 7933 7767 7947
rect 7713 7913 7727 7927
rect 7713 7853 7727 7867
rect 7733 7833 7747 7847
rect 7713 7813 7727 7827
rect 7553 7453 7567 7467
rect 7613 7413 7627 7427
rect 7593 7373 7607 7387
rect 7533 7333 7547 7347
rect 7573 7333 7587 7347
rect 7593 7313 7607 7327
rect 7573 7293 7587 7307
rect 7493 7113 7507 7127
rect 7513 7073 7527 7087
rect 7473 6953 7487 6967
rect 7553 7093 7567 7107
rect 7533 6933 7547 6947
rect 7493 6913 7507 6927
rect 7533 6893 7547 6907
rect 7453 6873 7467 6887
rect 7573 7073 7587 7087
rect 7573 7013 7587 7027
rect 7573 6973 7587 6987
rect 7553 6873 7567 6887
rect 7533 6853 7547 6867
rect 7553 6853 7567 6867
rect 7453 6833 7467 6847
rect 7553 6813 7567 6827
rect 7533 6693 7547 6707
rect 7453 6633 7467 6647
rect 7493 6613 7507 6627
rect 7593 6813 7607 6827
rect 7673 7553 7687 7567
rect 7653 7453 7667 7467
rect 7853 8493 7867 8507
rect 7833 8473 7847 8487
rect 7953 9233 7967 9247
rect 7933 9053 7947 9067
rect 8073 9753 8087 9767
rect 8053 9673 8067 9687
rect 8013 9573 8027 9587
rect 7993 9433 8007 9447
rect 7993 9093 8007 9107
rect 8133 9513 8147 9527
rect 8133 9493 8147 9507
rect 8033 9473 8047 9487
rect 8073 9473 8087 9487
rect 8113 9473 8127 9487
rect 8053 9453 8067 9467
rect 8053 9433 8067 9447
rect 8033 9353 8047 9367
rect 8033 9313 8047 9327
rect 7973 9033 7987 9047
rect 8013 9033 8027 9047
rect 7953 9013 7967 9027
rect 7933 8993 7947 9007
rect 7973 8993 7987 9007
rect 7913 8973 7927 8987
rect 8093 9393 8107 9407
rect 8093 9313 8107 9327
rect 8073 9293 8087 9307
rect 8073 9273 8087 9287
rect 8053 9033 8067 9047
rect 7933 8913 7947 8927
rect 7913 8673 7927 8687
rect 7913 8593 7927 8607
rect 7873 8433 7887 8447
rect 7893 8433 7907 8447
rect 7893 8393 7907 8407
rect 7813 8353 7827 8367
rect 7853 8353 7867 8367
rect 7793 8273 7807 8287
rect 7793 8173 7807 8187
rect 7773 7833 7787 7847
rect 7713 7413 7727 7427
rect 7673 7393 7687 7407
rect 7653 7373 7667 7387
rect 7633 7313 7647 7327
rect 7873 8293 7887 8307
rect 7893 8273 7907 8287
rect 7833 8073 7847 8087
rect 7933 8513 7947 8527
rect 7993 8973 8007 8987
rect 7993 8873 8007 8887
rect 7973 8793 7987 8807
rect 8033 8993 8047 9007
rect 8013 8673 8027 8687
rect 8013 8533 8027 8547
rect 7973 8493 7987 8507
rect 8033 8473 8047 8487
rect 7993 8453 8007 8467
rect 8033 8453 8047 8467
rect 7953 8393 7967 8407
rect 7953 8333 7967 8347
rect 7933 8093 7947 8107
rect 7853 8053 7867 8067
rect 7833 7973 7847 7987
rect 7833 7913 7847 7927
rect 7813 7793 7827 7807
rect 7793 7773 7807 7787
rect 7773 7653 7787 7667
rect 7733 7373 7747 7387
rect 7833 7573 7847 7587
rect 7873 8013 7887 8027
rect 7953 8033 7967 8047
rect 7933 7993 7947 8007
rect 7893 7973 7907 7987
rect 7933 7973 7947 7987
rect 7873 7933 7887 7947
rect 7893 7833 7907 7847
rect 7953 7933 7967 7947
rect 7873 7813 7887 7827
rect 7913 7813 7927 7827
rect 7953 7813 7967 7827
rect 7913 7793 7927 7807
rect 7873 7633 7887 7647
rect 7833 7533 7847 7547
rect 7853 7533 7867 7547
rect 7793 7513 7807 7527
rect 7793 7473 7807 7487
rect 7753 7353 7767 7367
rect 7693 7333 7707 7347
rect 7773 7333 7787 7347
rect 7753 7313 7767 7327
rect 7733 7193 7747 7207
rect 7673 7133 7687 7147
rect 7693 7093 7707 7107
rect 7653 7073 7667 7087
rect 7633 6993 7647 7007
rect 7693 6993 7707 7007
rect 7693 6933 7707 6947
rect 7653 6853 7667 6867
rect 7673 6853 7687 6867
rect 7713 6873 7727 6887
rect 7713 6853 7727 6867
rect 7733 6853 7747 6867
rect 7633 6833 7647 6847
rect 7673 6833 7687 6847
rect 7573 6673 7587 6687
rect 7613 6673 7627 6687
rect 7593 6633 7607 6647
rect 7573 6593 7587 6607
rect 7473 6533 7487 6547
rect 7553 6533 7567 6547
rect 7453 6473 7467 6487
rect 7413 6213 7427 6227
rect 7413 6193 7427 6207
rect 7453 6393 7467 6407
rect 7573 6433 7587 6447
rect 7533 6393 7547 6407
rect 7553 6373 7567 6387
rect 7473 6333 7487 6347
rect 7453 6253 7467 6267
rect 7433 6173 7447 6187
rect 7493 6173 7507 6187
rect 7353 5953 7367 5967
rect 7353 5933 7367 5947
rect 7333 5873 7347 5887
rect 7333 5433 7347 5447
rect 7473 6133 7487 6147
rect 7433 6113 7447 6127
rect 7453 6093 7467 6107
rect 7413 6073 7427 6087
rect 7393 5953 7407 5967
rect 7433 5933 7447 5947
rect 7533 6153 7547 6167
rect 7513 6133 7527 6147
rect 7513 6093 7527 6107
rect 7513 5993 7527 6007
rect 7493 5973 7507 5987
rect 7433 5893 7447 5907
rect 7513 5893 7527 5907
rect 7453 5873 7467 5887
rect 7473 5873 7487 5887
rect 7513 5873 7527 5887
rect 7493 5853 7507 5867
rect 7433 5713 7447 5727
rect 7473 5713 7487 5727
rect 7373 5653 7387 5667
rect 7393 5633 7407 5647
rect 7313 5373 7327 5387
rect 7353 5393 7367 5407
rect 7373 5353 7387 5367
rect 7333 5233 7347 5247
rect 7333 5213 7347 5227
rect 7373 5213 7387 5227
rect 7293 5173 7307 5187
rect 7273 5133 7287 5147
rect 7373 4953 7387 4967
rect 7273 4933 7287 4947
rect 7253 4893 7267 4907
rect 7353 4593 7367 4607
rect 7253 4533 7267 4547
rect 7313 4533 7327 4547
rect 7193 4493 7207 4507
rect 7213 4473 7227 4487
rect 7293 4473 7307 4487
rect 7453 5613 7467 5627
rect 7433 5553 7447 5567
rect 7453 5133 7467 5147
rect 7433 5013 7447 5027
rect 7613 6613 7627 6627
rect 7613 6593 7627 6607
rect 7693 6813 7707 6827
rect 7713 6753 7727 6767
rect 7773 7173 7787 7187
rect 7753 6693 7767 6707
rect 7753 6653 7767 6667
rect 7653 6413 7667 6427
rect 7613 6373 7627 6387
rect 7633 6373 7647 6387
rect 7593 6353 7607 6367
rect 7593 6133 7607 6147
rect 7633 6133 7647 6147
rect 7613 6113 7627 6127
rect 7633 5973 7647 5987
rect 7573 5853 7587 5867
rect 7553 5653 7567 5667
rect 7613 5653 7627 5667
rect 7553 5573 7567 5587
rect 7513 5553 7527 5567
rect 7533 5493 7547 5507
rect 7513 5433 7527 5447
rect 7553 5433 7567 5447
rect 7593 5433 7607 5447
rect 7573 5413 7587 5427
rect 7493 5353 7507 5367
rect 7693 6433 7707 6447
rect 7713 6433 7727 6447
rect 7733 6413 7747 6427
rect 7713 6373 7727 6387
rect 7673 6153 7687 6167
rect 7673 6113 7687 6127
rect 7733 6353 7747 6367
rect 7713 6093 7727 6107
rect 7713 5933 7727 5947
rect 7653 5613 7667 5627
rect 7653 5553 7667 5567
rect 7633 5273 7647 5287
rect 7633 5093 7647 5107
rect 7493 5073 7507 5087
rect 7473 4993 7487 5007
rect 7453 4973 7467 4987
rect 7453 4953 7467 4967
rect 7553 5053 7567 5067
rect 7513 4993 7527 5007
rect 7433 4933 7447 4947
rect 7473 4933 7487 4947
rect 7513 4933 7527 4947
rect 7413 4913 7427 4927
rect 7433 4813 7447 4827
rect 7453 4813 7467 4827
rect 7533 4753 7547 4767
rect 7513 4693 7527 4707
rect 7473 4653 7487 4667
rect 7433 4573 7447 4587
rect 7313 4453 7327 4467
rect 7373 4453 7387 4467
rect 7513 4473 7527 4487
rect 7493 4453 7507 4467
rect 7273 4433 7287 4447
rect 7393 4373 7407 4387
rect 7213 4173 7227 4187
rect 7233 4173 7247 4187
rect 7273 4173 7287 4187
rect 7233 4113 7247 4127
rect 7213 4073 7227 4087
rect 7253 3993 7267 4007
rect 7453 4353 7467 4367
rect 7433 4193 7447 4207
rect 7513 4213 7527 4227
rect 7433 4153 7447 4167
rect 7453 4153 7467 4167
rect 7473 4073 7487 4087
rect 7173 3953 7187 3967
rect 7153 3773 7167 3787
rect 7153 3413 7167 3427
rect 7153 3213 7167 3227
rect 7213 3873 7227 3887
rect 7433 3993 7447 4007
rect 7473 3933 7487 3947
rect 7373 3713 7387 3727
rect 7233 3693 7247 3707
rect 7333 3693 7347 3707
rect 7413 3693 7427 3707
rect 7693 5633 7707 5647
rect 7673 5373 7687 5387
rect 7733 5553 7747 5567
rect 7853 7413 7867 7427
rect 7833 7393 7847 7407
rect 7833 7353 7847 7367
rect 7813 7033 7827 7047
rect 7793 7013 7807 7027
rect 7793 6873 7807 6887
rect 7833 6973 7847 6987
rect 7893 7373 7907 7387
rect 7953 7773 7967 7787
rect 7973 7773 7987 7787
rect 8013 8213 8027 8227
rect 7993 7673 8007 7687
rect 8013 7573 8027 7587
rect 8013 7533 8027 7547
rect 7973 7513 7987 7527
rect 8073 9013 8087 9027
rect 8093 8993 8107 9007
rect 8073 8333 8087 8347
rect 8193 10433 8207 10447
rect 8253 10693 8267 10707
rect 8333 11333 8347 11347
rect 8473 11673 8487 11687
rect 8513 11673 8527 11687
rect 8593 11693 8607 11707
rect 8653 11693 8667 11707
rect 8573 11673 8587 11687
rect 8513 11513 8527 11527
rect 8533 11513 8547 11527
rect 8453 11493 8467 11507
rect 8593 11633 8607 11647
rect 8653 11633 8667 11647
rect 8633 11593 8647 11607
rect 8573 11433 8587 11447
rect 8553 11393 8567 11407
rect 8433 11313 8447 11327
rect 8313 11273 8327 11287
rect 8493 11273 8507 11287
rect 8553 11253 8567 11267
rect 8593 11253 8607 11267
rect 8353 11233 8367 11247
rect 8393 11213 8407 11227
rect 8453 11213 8467 11227
rect 8553 11213 8567 11227
rect 8333 11173 8347 11187
rect 8313 10713 8327 10727
rect 8293 10633 8307 10647
rect 8213 10413 8227 10427
rect 8193 10253 8207 10267
rect 8173 10213 8187 10227
rect 8213 10213 8227 10227
rect 8213 10193 8227 10207
rect 8213 9953 8227 9967
rect 8273 10453 8287 10467
rect 8293 10393 8307 10407
rect 8293 10073 8307 10087
rect 8273 9993 8287 10007
rect 8233 9933 8247 9947
rect 8253 9933 8267 9947
rect 8213 9873 8227 9887
rect 8273 9873 8287 9887
rect 8293 9853 8307 9867
rect 8273 9733 8287 9747
rect 8213 9713 8227 9727
rect 8193 9573 8207 9587
rect 8193 9513 8207 9527
rect 8173 9253 8187 9267
rect 8173 9233 8187 9247
rect 8153 9013 8167 9027
rect 8133 8953 8147 8967
rect 8173 8953 8187 8967
rect 8153 8893 8167 8907
rect 8113 8813 8127 8827
rect 8153 8773 8167 8787
rect 8133 8753 8147 8767
rect 8133 8733 8147 8747
rect 8173 8633 8187 8647
rect 8213 9453 8227 9467
rect 8293 9693 8307 9707
rect 8333 10573 8347 10587
rect 8373 11093 8387 11107
rect 8413 10873 8427 10887
rect 8513 11173 8527 11187
rect 8493 11093 8507 11107
rect 8593 10933 8607 10947
rect 8453 10813 8467 10827
rect 8393 10773 8407 10787
rect 8373 10513 8387 10527
rect 8353 10473 8367 10487
rect 8373 10453 8387 10467
rect 8333 10393 8347 10407
rect 8313 9513 8327 9527
rect 8373 10393 8387 10407
rect 8433 10673 8447 10687
rect 8493 10793 8507 10807
rect 8453 10533 8467 10547
rect 8393 10293 8407 10307
rect 8393 10233 8407 10247
rect 8453 10193 8467 10207
rect 8413 10133 8427 10147
rect 8473 10133 8487 10147
rect 8453 10033 8467 10047
rect 8393 9973 8407 9987
rect 8433 9973 8447 9987
rect 8353 9833 8367 9847
rect 8333 9493 8347 9507
rect 8273 9453 8287 9467
rect 8293 9453 8307 9467
rect 8253 9433 8267 9447
rect 8273 9293 8287 9307
rect 8233 9273 8247 9287
rect 8313 9433 8327 9447
rect 8313 9413 8327 9427
rect 8333 9413 8347 9427
rect 8313 9393 8327 9407
rect 8293 9053 8307 9067
rect 8233 8993 8247 9007
rect 8293 8953 8307 8967
rect 8253 8893 8267 8907
rect 8233 8813 8247 8827
rect 8233 8773 8247 8787
rect 8213 8753 8227 8767
rect 8233 8653 8247 8667
rect 8193 8593 8207 8607
rect 8133 8553 8147 8567
rect 8153 8553 8167 8567
rect 8173 8533 8187 8547
rect 8213 8533 8227 8547
rect 8153 8513 8167 8527
rect 8133 8493 8147 8507
rect 8193 8473 8207 8487
rect 8193 8453 8207 8467
rect 8233 8453 8247 8467
rect 8173 8333 8187 8347
rect 8053 8293 8067 8307
rect 8093 8293 8107 8307
rect 8153 8093 8167 8107
rect 8093 8053 8107 8067
rect 8073 8033 8087 8047
rect 8113 8033 8127 8047
rect 8053 7933 8067 7947
rect 8093 7913 8107 7927
rect 8093 7833 8107 7847
rect 8133 7833 8147 7847
rect 8113 7813 8127 7827
rect 8073 7793 8087 7807
rect 8073 7773 8087 7787
rect 8113 7753 8127 7767
rect 8053 7733 8067 7747
rect 8073 7733 8087 7747
rect 8093 7593 8107 7607
rect 8053 7533 8067 7547
rect 7953 7473 7967 7487
rect 7933 7373 7947 7387
rect 7953 7353 7967 7367
rect 7893 7313 7907 7327
rect 7953 7313 7967 7327
rect 7873 7253 7887 7267
rect 7913 7073 7927 7087
rect 7893 7053 7907 7067
rect 7933 7053 7947 7067
rect 7873 7013 7887 7027
rect 7933 7013 7947 7027
rect 7853 6953 7867 6967
rect 7853 6933 7867 6947
rect 7893 6893 7907 6907
rect 7893 6873 7907 6887
rect 7873 6853 7887 6867
rect 7833 6833 7847 6847
rect 7873 6713 7887 6727
rect 7933 6653 7947 6667
rect 7893 6573 7907 6587
rect 7933 6593 7947 6607
rect 7953 6573 7967 6587
rect 7813 6473 7827 6487
rect 7833 6473 7847 6487
rect 7913 6473 7927 6487
rect 7793 6393 7807 6407
rect 7773 6153 7787 6167
rect 7853 6433 7867 6447
rect 7933 6413 7947 6427
rect 7893 6393 7907 6407
rect 7833 6333 7847 6347
rect 7993 7453 8007 7467
rect 7993 7153 8007 7167
rect 7993 6973 8007 6987
rect 7993 6953 8007 6967
rect 8133 7693 8147 7707
rect 8273 8813 8287 8827
rect 8413 9953 8427 9967
rect 8433 9753 8447 9767
rect 8373 9733 8387 9747
rect 8413 9653 8427 9667
rect 8433 9593 8447 9607
rect 8393 9553 8407 9567
rect 8373 9513 8387 9527
rect 8353 9393 8367 9407
rect 8413 9473 8427 9487
rect 8453 9493 8467 9507
rect 8413 9393 8427 9407
rect 8613 10773 8627 10787
rect 8593 10733 8607 10747
rect 8573 10533 8587 10547
rect 8553 10433 8567 10447
rect 8513 10413 8527 10427
rect 8573 10393 8587 10407
rect 8913 11813 8927 11827
rect 8873 11653 8887 11667
rect 8813 11633 8827 11647
rect 8853 11633 8867 11647
rect 8713 11593 8727 11607
rect 8733 11313 8747 11327
rect 8753 11313 8767 11327
rect 8993 11833 9007 11847
rect 9053 11853 9067 11867
rect 9033 11833 9047 11847
rect 9233 11893 9247 11907
rect 9433 11893 9447 11907
rect 9973 11893 9987 11907
rect 9193 11833 9207 11847
rect 9173 11793 9187 11807
rect 9033 11733 9047 11747
rect 9013 11673 9027 11687
rect 8993 11633 9007 11647
rect 8933 11573 8947 11587
rect 8913 11413 8927 11427
rect 9013 11413 9027 11427
rect 8893 11393 8907 11407
rect 8853 11293 8867 11307
rect 8993 11293 9007 11307
rect 8713 11253 8727 11267
rect 8813 11253 8827 11267
rect 8713 11213 8727 11227
rect 8773 11193 8787 11207
rect 8693 11153 8707 11167
rect 8753 11153 8767 11167
rect 8713 10913 8727 10927
rect 8753 10913 8767 10927
rect 8773 10893 8787 10907
rect 8733 10873 8747 10887
rect 8693 10733 8707 10747
rect 8713 10733 8727 10747
rect 8773 10733 8787 10747
rect 8793 10733 8807 10747
rect 8833 11153 8847 11167
rect 8713 10673 8727 10687
rect 8733 10653 8747 10667
rect 8673 10513 8687 10527
rect 8593 10373 8607 10387
rect 8533 10353 8547 10367
rect 8653 10453 8667 10467
rect 8753 10493 8767 10507
rect 8513 10293 8527 10307
rect 8633 10293 8647 10307
rect 8493 9973 8507 9987
rect 8713 10413 8727 10427
rect 8673 10393 8687 10407
rect 8593 10253 8607 10267
rect 8653 10253 8667 10267
rect 8553 10233 8567 10247
rect 8713 10373 8727 10387
rect 8693 10313 8707 10327
rect 8633 10233 8647 10247
rect 8673 10233 8687 10247
rect 8573 10213 8587 10227
rect 8613 10073 8627 10087
rect 8573 10053 8587 10067
rect 8553 9693 8567 9707
rect 8513 9453 8527 9467
rect 8473 9413 8487 9427
rect 8493 9413 8507 9427
rect 8473 9353 8487 9367
rect 8433 9313 8447 9327
rect 8413 9253 8427 9267
rect 8433 9253 8447 9267
rect 8373 9213 8387 9227
rect 8453 9193 8467 9207
rect 8393 9153 8407 9167
rect 8433 9153 8447 9167
rect 8333 8953 8347 8967
rect 8313 8893 8327 8907
rect 8373 8853 8387 8867
rect 8313 8813 8327 8827
rect 8433 9073 8447 9087
rect 8453 9073 8467 9087
rect 8413 8973 8427 8987
rect 8413 8953 8427 8967
rect 8473 8973 8487 8987
rect 8393 8793 8407 8807
rect 8373 8633 8387 8647
rect 8313 8593 8327 8607
rect 8353 8593 8367 8607
rect 8273 8473 8287 8487
rect 8253 8333 8267 8347
rect 8293 8273 8307 8287
rect 8233 8253 8247 8267
rect 8213 8093 8227 8107
rect 8193 8013 8207 8027
rect 8193 7993 8207 8007
rect 8193 7793 8207 7807
rect 8173 7613 8187 7627
rect 8353 8533 8367 8547
rect 8333 8353 8347 8367
rect 8313 8073 8327 8087
rect 8273 8013 8287 8027
rect 8293 7933 8307 7947
rect 8313 7873 8327 7887
rect 8273 7813 8287 7827
rect 8293 7813 8307 7827
rect 8113 7453 8127 7467
rect 8113 7433 8127 7447
rect 8093 7393 8107 7407
rect 8053 7333 8067 7347
rect 8033 7313 8047 7327
rect 8233 7593 8247 7607
rect 8253 7593 8267 7607
rect 8153 7573 8167 7587
rect 8173 7553 8187 7567
rect 8213 7553 8227 7567
rect 8233 7533 8247 7547
rect 8213 7433 8227 7447
rect 8193 7253 8207 7267
rect 8153 7213 8167 7227
rect 8173 7173 8187 7187
rect 8133 7133 8147 7147
rect 8153 7113 8167 7127
rect 8173 7073 8187 7087
rect 8033 7053 8047 7067
rect 8053 7053 8067 7067
rect 8093 7053 8107 7067
rect 8173 7053 8187 7067
rect 8073 7033 8087 7047
rect 8073 6913 8087 6927
rect 8033 6873 8047 6887
rect 8053 6853 8067 6867
rect 8093 6853 8107 6867
rect 8013 6833 8027 6847
rect 8133 6833 8147 6847
rect 8053 6713 8067 6727
rect 8113 6613 8127 6627
rect 7993 6573 8007 6587
rect 7973 6233 7987 6247
rect 7873 6153 7887 6167
rect 7893 6153 7907 6167
rect 7773 6093 7787 6107
rect 7813 6093 7827 6107
rect 7753 5533 7767 5547
rect 7853 6033 7867 6047
rect 7973 6133 7987 6147
rect 7973 6093 7987 6107
rect 7893 6073 7907 6087
rect 7833 5933 7847 5947
rect 7873 5933 7887 5947
rect 7873 5913 7887 5927
rect 7853 5893 7867 5907
rect 7873 5873 7887 5887
rect 7853 5853 7867 5867
rect 7793 5613 7807 5627
rect 7773 5473 7787 5487
rect 7833 5573 7847 5587
rect 7833 5533 7847 5547
rect 7753 5453 7767 5467
rect 7793 5453 7807 5467
rect 7733 5433 7747 5447
rect 7813 5413 7827 5427
rect 7793 5393 7807 5407
rect 7813 5373 7827 5387
rect 7793 5173 7807 5187
rect 7753 5153 7767 5167
rect 7733 5073 7747 5087
rect 7653 5033 7667 5047
rect 7573 5013 7587 5027
rect 7613 4973 7627 4987
rect 7793 4973 7807 4987
rect 7853 5253 7867 5267
rect 7893 5833 7907 5847
rect 8053 6573 8067 6587
rect 8093 6573 8107 6587
rect 8073 6413 8087 6427
rect 8033 6393 8047 6407
rect 8093 6353 8107 6367
rect 8073 6173 8087 6187
rect 8033 6113 8047 6127
rect 8093 6153 8107 6167
rect 8013 6093 8027 6107
rect 8053 6073 8067 6087
rect 8093 6073 8107 6087
rect 8193 6713 8207 6727
rect 8173 6593 8187 6607
rect 8193 6593 8207 6607
rect 8153 6573 8167 6587
rect 8113 5973 8127 5987
rect 8053 5913 8067 5927
rect 7993 5873 8007 5887
rect 8053 5713 8067 5727
rect 7973 5693 7987 5707
rect 8273 7553 8287 7567
rect 8273 7433 8287 7447
rect 8253 7353 8267 7367
rect 8253 7333 8267 7347
rect 8273 7293 8287 7307
rect 8233 7273 8247 7287
rect 8253 6933 8267 6947
rect 8393 8473 8407 8487
rect 8373 8333 8387 8347
rect 8353 7833 8367 7847
rect 8413 8433 8427 8447
rect 8593 9953 8607 9967
rect 8633 9953 8647 9967
rect 8613 9933 8627 9947
rect 8653 9913 8667 9927
rect 8593 9853 8607 9867
rect 8613 9793 8627 9807
rect 8693 9793 8707 9807
rect 8673 9773 8687 9787
rect 8633 9753 8647 9767
rect 8653 9753 8667 9767
rect 8593 9453 8607 9467
rect 8633 9453 8647 9467
rect 8693 9733 8707 9747
rect 8673 9453 8687 9467
rect 8633 9433 8647 9447
rect 8653 9433 8667 9447
rect 8633 9333 8647 9347
rect 8673 9293 8687 9307
rect 8653 9273 8667 9287
rect 8573 9233 8587 9247
rect 8553 9133 8567 9147
rect 8533 8993 8547 9007
rect 8573 8973 8587 8987
rect 8513 8933 8527 8947
rect 8453 8813 8467 8827
rect 8493 8793 8507 8807
rect 8493 8653 8507 8667
rect 8473 8533 8487 8547
rect 8473 8493 8487 8507
rect 8393 8313 8407 8327
rect 8473 8393 8487 8407
rect 8453 8293 8467 8307
rect 8433 8273 8447 8287
rect 8533 8813 8547 8827
rect 8533 8653 8547 8667
rect 8653 9073 8667 9087
rect 8773 10413 8787 10427
rect 8753 10293 8767 10307
rect 8813 10473 8827 10487
rect 8813 10333 8827 10347
rect 8953 11193 8967 11207
rect 8933 11153 8947 11167
rect 8933 11113 8947 11127
rect 8893 11093 8907 11107
rect 8933 10993 8947 11007
rect 8853 10933 8867 10947
rect 9013 10973 9027 10987
rect 8953 10953 8967 10967
rect 8933 10913 8947 10927
rect 8973 10913 8987 10927
rect 9393 11873 9407 11887
rect 9533 11873 9547 11887
rect 10553 11913 10567 11927
rect 10613 11913 10627 11927
rect 11293 11913 11307 11927
rect 12073 11913 12087 11927
rect 10593 11893 10607 11907
rect 9233 11853 9247 11867
rect 9213 11693 9227 11707
rect 9173 11673 9187 11687
rect 9073 11653 9087 11667
rect 9113 11653 9127 11667
rect 9053 11633 9067 11647
rect 9093 11633 9107 11647
rect 9153 11633 9167 11647
rect 9073 11473 9087 11487
rect 9053 11413 9067 11427
rect 8993 10893 9007 10907
rect 8933 10813 8947 10827
rect 8873 10773 8887 10787
rect 8893 10773 8907 10787
rect 8853 10733 8867 10747
rect 8853 10553 8867 10567
rect 8913 10753 8927 10767
rect 8893 10693 8907 10707
rect 8873 10473 8887 10487
rect 9033 10913 9047 10927
rect 9013 10753 9027 10767
rect 9013 10733 9027 10747
rect 8993 10713 9007 10727
rect 8973 10693 8987 10707
rect 8893 10413 8907 10427
rect 8793 10253 8807 10267
rect 8793 10233 8807 10247
rect 8773 10173 8787 10187
rect 8733 10113 8747 10127
rect 8833 10253 8847 10267
rect 8853 10253 8867 10267
rect 8813 9993 8827 10007
rect 8733 9933 8747 9947
rect 8733 9913 8747 9927
rect 8773 9913 8787 9927
rect 8793 9913 8807 9927
rect 8793 9793 8807 9807
rect 8753 9773 8767 9787
rect 8833 9913 8847 9927
rect 8833 9853 8847 9867
rect 8813 9773 8827 9787
rect 8733 9613 8747 9627
rect 8693 9073 8707 9087
rect 8713 9073 8727 9087
rect 8693 9053 8707 9067
rect 8673 8973 8687 8987
rect 8653 8873 8667 8887
rect 8653 8813 8667 8827
rect 8633 8793 8647 8807
rect 8653 8773 8667 8787
rect 8613 8753 8627 8767
rect 8593 8713 8607 8727
rect 8513 8553 8527 8567
rect 8553 8553 8567 8567
rect 8533 8533 8547 8547
rect 8553 8513 8567 8527
rect 8573 8513 8587 8527
rect 8513 8493 8527 8507
rect 8533 8453 8547 8467
rect 8573 8453 8587 8467
rect 8593 8453 8607 8467
rect 8493 8293 8507 8307
rect 8413 8253 8427 8267
rect 8413 8193 8427 8207
rect 8413 8173 8427 8187
rect 8433 8033 8447 8047
rect 8413 8013 8427 8027
rect 8393 7933 8407 7947
rect 8373 7813 8387 7827
rect 8473 7873 8487 7887
rect 8553 8353 8567 8367
rect 8533 8293 8547 8307
rect 8533 8053 8547 8067
rect 8513 7873 8527 7887
rect 8433 7793 8447 7807
rect 8333 7773 8347 7787
rect 8433 7693 8447 7707
rect 8333 7613 8347 7627
rect 8373 7573 8387 7587
rect 8373 7553 8387 7567
rect 8353 7533 8367 7547
rect 8393 7533 8407 7547
rect 8313 7373 8327 7387
rect 8473 7813 8487 7827
rect 8513 7813 8527 7827
rect 8633 8653 8647 8667
rect 8673 8633 8687 8647
rect 8713 8893 8727 8907
rect 8773 9753 8787 9767
rect 8813 9753 8827 9767
rect 8773 9693 8787 9707
rect 8813 9513 8827 9527
rect 8813 9493 8827 9507
rect 8773 9433 8787 9447
rect 8753 9013 8767 9027
rect 8793 9413 8807 9427
rect 8973 10533 8987 10547
rect 8953 10413 8967 10427
rect 8873 10173 8887 10187
rect 8853 9733 8867 9747
rect 8873 9713 8887 9727
rect 8853 9653 8867 9667
rect 8873 9593 8887 9607
rect 8853 9493 8867 9507
rect 8853 9453 8867 9467
rect 8853 9433 8867 9447
rect 8873 9253 8887 9267
rect 8753 8973 8767 8987
rect 8733 8753 8747 8767
rect 8733 8553 8747 8567
rect 8833 9213 8847 9227
rect 8873 9193 8887 9207
rect 8853 9013 8867 9027
rect 8813 8973 8827 8987
rect 8793 8953 8807 8967
rect 8953 10253 8967 10267
rect 8913 10233 8927 10247
rect 8953 9933 8967 9947
rect 9013 10273 9027 10287
rect 8993 10213 9007 10227
rect 9093 11373 9107 11387
rect 9153 11413 9167 11427
rect 9113 11273 9127 11287
rect 9153 11153 9167 11167
rect 9453 11853 9467 11867
rect 9413 11833 9427 11847
rect 9313 11773 9327 11787
rect 9413 11773 9427 11787
rect 9273 11653 9287 11667
rect 9333 11753 9347 11767
rect 9393 11753 9407 11767
rect 9293 11633 9307 11647
rect 9333 11633 9347 11647
rect 9313 11613 9327 11627
rect 9333 11613 9347 11627
rect 9313 11473 9327 11487
rect 9313 11413 9327 11427
rect 9293 11393 9307 11407
rect 9253 11373 9267 11387
rect 9193 11353 9207 11367
rect 9193 11213 9207 11227
rect 9313 11193 9327 11207
rect 9173 10953 9187 10967
rect 9113 10933 9127 10947
rect 9153 10913 9167 10927
rect 9193 10913 9207 10927
rect 9173 10893 9187 10907
rect 9213 10893 9227 10907
rect 9233 10813 9247 10827
rect 9133 10713 9147 10727
rect 9173 10713 9187 10727
rect 9053 10573 9067 10587
rect 9053 10513 9067 10527
rect 9033 10153 9047 10167
rect 8993 9873 9007 9887
rect 8973 9793 8987 9807
rect 9173 10493 9187 10507
rect 9093 10473 9107 10487
rect 9113 10393 9127 10407
rect 9133 10393 9147 10407
rect 9133 10353 9147 10367
rect 9113 10273 9127 10287
rect 9053 10113 9067 10127
rect 9073 9973 9087 9987
rect 9033 9793 9047 9807
rect 8953 9773 8967 9787
rect 8993 9773 9007 9787
rect 9033 9773 9047 9787
rect 8913 9613 8927 9627
rect 8933 9453 8947 9467
rect 8933 9413 8947 9427
rect 8913 9213 8927 9227
rect 8993 9753 9007 9767
rect 8973 9733 8987 9747
rect 9013 9713 9027 9727
rect 9193 10373 9207 10387
rect 9193 10313 9207 10327
rect 9213 10313 9227 10327
rect 9213 10233 9227 10247
rect 9133 10193 9147 10207
rect 9173 10133 9187 10147
rect 9133 10073 9147 10087
rect 9313 10693 9327 10707
rect 9273 10453 9287 10467
rect 9373 11413 9387 11427
rect 9373 11373 9387 11387
rect 9373 11193 9387 11207
rect 9353 11153 9367 11167
rect 9393 11033 9407 11047
rect 9393 10953 9407 10967
rect 9373 10913 9387 10927
rect 9353 10773 9367 10787
rect 9653 11833 9667 11847
rect 9873 11813 9887 11827
rect 9833 11773 9847 11787
rect 9533 11753 9547 11767
rect 9633 11753 9647 11767
rect 9433 11653 9447 11667
rect 9473 11653 9487 11667
rect 9453 11633 9467 11647
rect 9493 11613 9507 11627
rect 9433 11553 9447 11567
rect 9473 11413 9487 11427
rect 9493 11373 9507 11387
rect 9793 11673 9807 11687
rect 9833 11673 9847 11687
rect 9673 11653 9687 11667
rect 9693 11653 9707 11667
rect 9873 11673 9887 11687
rect 9853 11613 9867 11627
rect 9693 11593 9707 11607
rect 9793 11513 9807 11527
rect 9713 11433 9727 11447
rect 9633 11373 9647 11387
rect 9593 11353 9607 11367
rect 9453 11313 9467 11327
rect 9433 11193 9447 11207
rect 9413 10853 9427 10867
rect 9353 10713 9367 10727
rect 9393 10713 9407 10727
rect 9433 10673 9447 10687
rect 9333 10453 9347 10467
rect 9253 10433 9267 10447
rect 9273 10413 9287 10427
rect 9333 10433 9347 10447
rect 9293 10393 9307 10407
rect 9633 11333 9647 11347
rect 9593 11293 9607 11307
rect 9553 11213 9567 11227
rect 9593 11213 9607 11227
rect 9473 10653 9487 10667
rect 9453 10513 9467 10527
rect 9453 10413 9467 10427
rect 9433 10333 9447 10347
rect 9453 10253 9467 10267
rect 9253 10213 9267 10227
rect 9413 10213 9427 10227
rect 9453 10193 9467 10207
rect 9253 10153 9267 10167
rect 9233 10053 9247 10067
rect 9193 10013 9207 10027
rect 9153 9973 9167 9987
rect 9173 9893 9187 9907
rect 9133 9793 9147 9807
rect 9193 9793 9207 9807
rect 9113 9693 9127 9707
rect 9073 9653 9087 9667
rect 8993 9613 9007 9627
rect 9013 9473 9027 9487
rect 9113 9573 9127 9587
rect 9113 9513 9127 9527
rect 9073 9433 9087 9447
rect 9113 9433 9127 9447
rect 9053 9373 9067 9387
rect 9013 9293 9027 9307
rect 8973 9273 8987 9287
rect 8953 9253 8967 9267
rect 9033 9273 9047 9287
rect 9013 9253 9027 9267
rect 9033 9213 9047 9227
rect 8973 9193 8987 9207
rect 8933 9173 8947 9187
rect 8893 9013 8907 9027
rect 8873 8953 8887 8967
rect 8893 8933 8907 8947
rect 8813 8813 8827 8827
rect 8853 8813 8867 8827
rect 8793 8713 8807 8727
rect 8753 8533 8767 8547
rect 8613 8353 8627 8367
rect 8733 8353 8747 8367
rect 8593 8333 8607 8347
rect 8693 8333 8707 8347
rect 8573 8053 8587 8067
rect 8653 8313 8667 8327
rect 8613 8273 8627 8287
rect 8613 8233 8627 8247
rect 8573 7973 8587 7987
rect 8673 7913 8687 7927
rect 8553 7893 8567 7907
rect 8633 7893 8647 7907
rect 8713 8073 8727 8087
rect 8633 7873 8647 7887
rect 8693 7873 8707 7887
rect 8713 7873 8727 7887
rect 8613 7853 8627 7867
rect 8553 7833 8567 7847
rect 8613 7653 8627 7667
rect 8613 7593 8627 7607
rect 8513 7553 8527 7567
rect 8553 7553 8567 7567
rect 8573 7553 8587 7567
rect 8653 7853 8667 7867
rect 8693 7853 8707 7867
rect 8493 7533 8507 7547
rect 8593 7533 8607 7547
rect 8633 7533 8647 7547
rect 8453 7433 8467 7447
rect 8453 7373 8467 7387
rect 8473 7373 8487 7387
rect 8673 7833 8687 7847
rect 8713 7833 8727 7847
rect 8693 7693 8707 7707
rect 8673 7613 8687 7627
rect 8673 7553 8687 7567
rect 8553 7513 8567 7527
rect 8653 7513 8667 7527
rect 8513 7493 8527 7507
rect 8313 7293 8327 7307
rect 8493 7293 8507 7307
rect 8473 7253 8487 7267
rect 8533 7433 8547 7447
rect 8473 7013 8487 7027
rect 8453 6993 8467 7007
rect 8373 6973 8387 6987
rect 8313 6953 8327 6967
rect 8313 6933 8327 6947
rect 8313 6873 8327 6887
rect 8333 6873 8347 6887
rect 8273 6833 8287 6847
rect 8293 6833 8307 6847
rect 8253 6773 8267 6787
rect 8333 6793 8347 6807
rect 8273 6593 8287 6607
rect 8313 6593 8327 6607
rect 8213 6453 8227 6467
rect 8253 6413 8267 6427
rect 8213 6373 8227 6387
rect 8273 6373 8287 6387
rect 8333 6533 8347 6547
rect 8193 6173 8207 6187
rect 8233 6353 8247 6367
rect 8273 6153 8287 6167
rect 8213 6133 8227 6147
rect 8253 6133 8267 6147
rect 8233 6113 8247 6127
rect 8173 5933 8187 5947
rect 8153 5753 8167 5767
rect 8193 5853 8207 5867
rect 8213 5833 8227 5847
rect 8173 5733 8187 5747
rect 7993 5633 8007 5647
rect 8073 5653 8087 5667
rect 8173 5653 8187 5667
rect 8133 5633 8147 5647
rect 8073 5613 8087 5627
rect 8153 5613 8167 5627
rect 8033 5593 8047 5607
rect 8193 5593 8207 5607
rect 7933 5513 7947 5527
rect 8113 5493 8127 5507
rect 7933 5453 7947 5467
rect 7913 5433 7927 5447
rect 7973 5433 7987 5447
rect 8073 5433 8087 5447
rect 8133 5433 8147 5447
rect 7953 5413 7967 5427
rect 8073 5373 8087 5387
rect 8433 6913 8447 6927
rect 8413 6773 8427 6787
rect 8433 6593 8447 6607
rect 8533 6913 8547 6927
rect 8493 6873 8507 6887
rect 8513 6853 8527 6867
rect 8473 6833 8487 6847
rect 8453 6573 8467 6587
rect 8393 6533 8407 6547
rect 8373 6473 8387 6487
rect 8453 6553 8467 6567
rect 8413 6473 8427 6487
rect 8433 6413 8447 6427
rect 8453 6393 8467 6407
rect 8533 6413 8547 6427
rect 8513 6213 8527 6227
rect 8373 6153 8387 6167
rect 8613 7473 8627 7487
rect 8673 7433 8687 7447
rect 8673 7393 8687 7407
rect 8613 7353 8627 7367
rect 8673 7353 8687 7367
rect 8633 7193 8647 7207
rect 8593 7113 8607 7127
rect 8573 7073 8587 7087
rect 8713 7593 8727 7607
rect 8773 8493 8787 8507
rect 8773 8333 8787 8347
rect 8773 8153 8787 8167
rect 8773 8073 8787 8087
rect 8773 8033 8787 8047
rect 8853 8793 8867 8807
rect 8833 8773 8847 8787
rect 8873 8753 8887 8767
rect 8893 8533 8907 8547
rect 8813 8493 8827 8507
rect 8873 8513 8887 8527
rect 8893 8353 8907 8367
rect 8933 9033 8947 9047
rect 8953 9013 8967 9027
rect 8993 9013 9007 9027
rect 8973 8993 8987 9007
rect 8973 8973 8987 8987
rect 9033 8973 9047 8987
rect 8933 8853 8947 8867
rect 8933 8833 8947 8847
rect 8953 8793 8967 8807
rect 9033 8913 9047 8927
rect 9073 9013 9087 9027
rect 9073 8973 9087 8987
rect 9113 9233 9127 9247
rect 9093 8913 9107 8927
rect 9053 8833 9067 8847
rect 9093 8833 9107 8847
rect 9053 8793 9067 8807
rect 8973 8773 8987 8787
rect 8993 8773 9007 8787
rect 9073 8773 9087 8787
rect 9033 8733 9047 8747
rect 9073 8593 9087 8607
rect 9013 8573 9027 8587
rect 9053 8573 9067 8587
rect 8933 8553 8947 8567
rect 8933 8513 8947 8527
rect 8973 8513 8987 8527
rect 8833 8333 8847 8347
rect 8853 8333 8867 8347
rect 8913 8333 8927 8347
rect 8833 8313 8847 8327
rect 8853 8213 8867 8227
rect 8813 8073 8827 8087
rect 8913 8293 8927 8307
rect 8893 8093 8907 8107
rect 8853 8053 8867 8067
rect 8813 8033 8827 8047
rect 8893 8033 8907 8047
rect 8833 8013 8847 8027
rect 8873 8013 8887 8027
rect 8893 7973 8907 7987
rect 8813 7953 8827 7967
rect 8873 7933 8887 7947
rect 8813 7913 8827 7927
rect 8853 7913 8867 7927
rect 8833 7833 8847 7847
rect 8813 7813 8827 7827
rect 8833 7753 8847 7767
rect 8773 7593 8787 7607
rect 8793 7593 8807 7607
rect 8753 7573 8767 7587
rect 8793 7553 8807 7567
rect 8753 7533 8767 7547
rect 8953 8493 8967 8507
rect 9033 8553 9047 8567
rect 9013 8473 9027 8487
rect 8953 8313 8967 8327
rect 8933 8013 8947 8027
rect 8933 7993 8947 8007
rect 8913 7933 8927 7947
rect 8893 7853 8907 7867
rect 8893 7833 8907 7847
rect 8933 7833 8947 7847
rect 8913 7813 8927 7827
rect 8893 7773 8907 7787
rect 8733 7513 8747 7527
rect 8813 7513 8827 7527
rect 8713 7373 8727 7387
rect 8693 7313 8707 7327
rect 8813 7453 8827 7467
rect 8793 7373 8807 7387
rect 8873 7393 8887 7407
rect 8933 7673 8947 7687
rect 8913 7653 8927 7667
rect 8913 7533 8927 7547
rect 8753 7313 8767 7327
rect 8893 7313 8907 7327
rect 8713 7073 8727 7087
rect 9053 8513 9067 8527
rect 9033 8313 9047 8327
rect 8993 8293 9007 8307
rect 9033 8293 9047 8307
rect 8973 7873 8987 7887
rect 9053 8273 9067 8287
rect 9013 8193 9027 8207
rect 9073 8193 9087 8207
rect 9053 8053 9067 8067
rect 9013 8033 9027 8047
rect 8993 7653 9007 7667
rect 8973 7573 8987 7587
rect 9033 8013 9047 8027
rect 9073 7993 9087 8007
rect 9033 7893 9047 7907
rect 9113 8793 9127 8807
rect 9113 8633 9127 8647
rect 9173 9773 9187 9787
rect 9153 9733 9167 9747
rect 9233 9753 9247 9767
rect 9213 9673 9227 9687
rect 9173 9533 9187 9547
rect 9153 9513 9167 9527
rect 9213 9493 9227 9507
rect 9193 9453 9207 9467
rect 9233 9433 9247 9447
rect 9193 9293 9207 9307
rect 9333 10073 9347 10087
rect 9333 10033 9347 10047
rect 9293 10013 9307 10027
rect 9273 9953 9287 9967
rect 9193 9013 9207 9027
rect 9253 9253 9267 9267
rect 9253 9173 9267 9187
rect 9153 8933 9167 8947
rect 9213 8973 9227 8987
rect 9453 10113 9467 10127
rect 9453 9973 9467 9987
rect 9373 9953 9387 9967
rect 9353 9913 9367 9927
rect 9313 9893 9327 9907
rect 9293 9733 9307 9747
rect 9293 9713 9307 9727
rect 9273 9133 9287 9147
rect 9433 9853 9447 9867
rect 9393 9773 9407 9787
rect 9413 9753 9427 9767
rect 9333 9733 9347 9747
rect 9413 9733 9427 9747
rect 9373 9673 9387 9687
rect 9393 9493 9407 9507
rect 9333 9453 9347 9467
rect 9353 9373 9367 9387
rect 9413 9373 9427 9387
rect 9313 9353 9327 9367
rect 9453 9693 9467 9707
rect 9453 9353 9467 9367
rect 9353 9213 9367 9227
rect 9433 9253 9447 9267
rect 9413 9233 9427 9247
rect 9453 9153 9467 9167
rect 9373 9053 9387 9067
rect 9293 8993 9307 9007
rect 9293 8973 9307 8987
rect 9253 8893 9267 8907
rect 9173 8673 9187 8687
rect 9133 8553 9147 8567
rect 9113 8473 9127 8487
rect 9173 8493 9187 8507
rect 9233 8793 9247 8807
rect 9253 8673 9267 8687
rect 9233 8473 9247 8487
rect 9153 8453 9167 8467
rect 9213 8453 9227 8467
rect 9133 8193 9147 8207
rect 9113 7893 9127 7907
rect 9373 9013 9387 9027
rect 9353 8993 9367 9007
rect 9313 8933 9327 8947
rect 9393 8933 9407 8947
rect 9353 8893 9367 8907
rect 9353 8873 9367 8887
rect 9313 8793 9327 8807
rect 9313 8653 9327 8667
rect 9433 8793 9447 8807
rect 9373 8773 9387 8787
rect 9353 8633 9367 8647
rect 9453 8773 9467 8787
rect 9413 8753 9427 8767
rect 9453 8613 9467 8627
rect 9373 8593 9387 8607
rect 9373 8573 9387 8587
rect 9333 8513 9347 8527
rect 9293 8373 9307 8387
rect 9293 8353 9307 8367
rect 9173 8133 9187 8147
rect 9173 8013 9187 8027
rect 9253 8273 9267 8287
rect 9253 8233 9267 8247
rect 9253 8093 9267 8107
rect 9213 8013 9227 8027
rect 9193 7993 9207 8007
rect 9173 7933 9187 7947
rect 9193 7933 9207 7947
rect 9053 7853 9067 7867
rect 9093 7853 9107 7867
rect 9033 7813 9047 7827
rect 9073 7813 9087 7827
rect 9113 7813 9127 7827
rect 9153 7713 9167 7727
rect 9133 7693 9147 7707
rect 9013 7613 9027 7627
rect 9053 7593 9067 7607
rect 9013 7573 9027 7587
rect 8973 7533 8987 7547
rect 8953 7493 8967 7507
rect 8933 7373 8947 7387
rect 8973 7373 8987 7387
rect 8913 7113 8927 7127
rect 8873 7093 8887 7107
rect 8833 7073 8847 7087
rect 8693 7053 8707 7067
rect 8773 7053 8787 7067
rect 8673 7033 8687 7047
rect 8733 7033 8747 7047
rect 8713 6993 8727 7007
rect 8673 6953 8687 6967
rect 8653 6853 8667 6867
rect 8693 6853 8707 6867
rect 8893 7073 8907 7087
rect 8933 7073 8947 7087
rect 8873 6973 8887 6987
rect 8853 6853 8867 6867
rect 8853 6833 8867 6847
rect 8753 6793 8767 6807
rect 8733 6773 8747 6787
rect 8713 6733 8727 6747
rect 8593 6613 8607 6627
rect 8593 6593 8607 6607
rect 8633 6593 8647 6607
rect 8673 6593 8687 6607
rect 8573 6573 8587 6587
rect 8593 6493 8607 6507
rect 8653 6533 8667 6547
rect 8673 6473 8687 6487
rect 8613 6413 8627 6427
rect 8633 6393 8647 6407
rect 8613 6373 8627 6387
rect 8553 6313 8567 6327
rect 8553 6213 8567 6227
rect 8353 6113 8367 6127
rect 8533 6113 8547 6127
rect 8533 6073 8547 6087
rect 8333 5993 8347 6007
rect 8413 5993 8427 6007
rect 8393 5933 8407 5947
rect 8253 5833 8267 5847
rect 8233 5733 8247 5747
rect 8233 5613 8247 5627
rect 8213 5393 8227 5407
rect 8193 5273 8207 5287
rect 8213 5253 8227 5267
rect 7973 5173 7987 5187
rect 7913 5153 7927 5167
rect 7833 5053 7847 5067
rect 7873 5053 7887 5067
rect 7933 5133 7947 5147
rect 7933 4993 7947 5007
rect 8113 5073 8127 5087
rect 8053 5053 8067 5067
rect 8073 5053 8087 5067
rect 8033 5033 8047 5047
rect 7813 4773 7827 4787
rect 7953 4713 7967 4727
rect 7993 4693 8007 4707
rect 8013 4693 8027 4707
rect 7853 4673 7867 4687
rect 7953 4673 7967 4687
rect 7633 4633 7647 4647
rect 7653 4633 7667 4647
rect 7693 4573 7707 4587
rect 7693 4553 7707 4567
rect 7793 4553 7807 4567
rect 7833 4553 7847 4567
rect 7653 4493 7667 4507
rect 7673 4493 7687 4507
rect 7573 4473 7587 4487
rect 7613 4473 7627 4487
rect 7833 4513 7847 4527
rect 7853 4513 7867 4527
rect 7893 4513 7907 4527
rect 7853 4493 7867 4507
rect 7793 4453 7807 4467
rect 7653 4293 7667 4307
rect 7713 4193 7727 4207
rect 7613 4073 7627 4087
rect 7553 3733 7567 3747
rect 7313 3493 7327 3507
rect 7273 3453 7287 3467
rect 7233 3253 7247 3267
rect 7213 3233 7227 3247
rect 7253 3233 7267 3247
rect 7293 3233 7307 3247
rect 7233 3213 7247 3227
rect 7213 3173 7227 3187
rect 7253 3093 7267 3107
rect 7213 3073 7227 3087
rect 7193 2993 7207 3007
rect 7173 2873 7187 2887
rect 7133 2793 7147 2807
rect 7113 2753 7127 2767
rect 7413 3673 7427 3687
rect 7693 4173 7707 4187
rect 7733 4173 7747 4187
rect 7653 4153 7667 4167
rect 7833 4173 7847 4187
rect 7813 3993 7827 4007
rect 7673 3973 7687 3987
rect 7753 3973 7767 3987
rect 7813 3973 7827 3987
rect 7633 3953 7647 3967
rect 7793 3933 7807 3947
rect 7753 3773 7767 3787
rect 7633 3713 7647 3727
rect 7673 3713 7687 3727
rect 7573 3673 7587 3687
rect 7613 3673 7627 3687
rect 7373 3633 7387 3647
rect 7453 3633 7467 3647
rect 7353 3293 7367 3307
rect 7333 3153 7347 3167
rect 7293 3093 7307 3107
rect 7273 3053 7287 3067
rect 7233 3033 7247 3047
rect 7273 3033 7287 3047
rect 7273 2993 7287 3007
rect 7173 2733 7187 2747
rect 7213 2733 7227 2747
rect 7093 2553 7107 2567
rect 7133 2553 7147 2567
rect 6973 2533 6987 2547
rect 7013 2433 7027 2447
rect 7093 2373 7107 2387
rect 7253 2713 7267 2727
rect 7233 2693 7247 2707
rect 7173 2513 7187 2527
rect 7173 2493 7187 2507
rect 7013 2333 7027 2347
rect 7153 2333 7167 2347
rect 6893 2253 6907 2267
rect 6993 2293 7007 2307
rect 6913 2233 6927 2247
rect 6873 2173 6887 2187
rect 6933 2173 6947 2187
rect 6913 2073 6927 2087
rect 6833 2053 6847 2067
rect 6853 2033 6867 2047
rect 6793 2013 6807 2027
rect 6833 2013 6847 2027
rect 6733 1953 6747 1967
rect 6793 1793 6807 1807
rect 6773 1773 6787 1787
rect 6693 1753 6707 1767
rect 6753 1753 6767 1767
rect 6673 1713 6687 1727
rect 6693 1593 6707 1607
rect 6733 1593 6747 1607
rect 6713 1553 6727 1567
rect 6733 1493 6747 1507
rect 6653 1473 6667 1487
rect 6633 1373 6647 1387
rect 6593 1353 6607 1367
rect 6633 1333 6647 1347
rect 6693 1333 6707 1347
rect 6673 1313 6687 1327
rect 6613 1293 6627 1307
rect 6633 1253 6647 1267
rect 6693 1253 6707 1267
rect 6653 1233 6667 1247
rect 6693 1133 6707 1147
rect 6593 1093 6607 1107
rect 6653 1093 6667 1107
rect 6633 813 6647 827
rect 6653 753 6667 767
rect 6593 733 6607 747
rect 6613 693 6627 707
rect 6573 613 6587 627
rect 6773 1593 6787 1607
rect 6753 1373 6767 1387
rect 6833 1553 6847 1567
rect 6813 1353 6827 1367
rect 6773 1333 6787 1347
rect 6753 1313 6767 1327
rect 6833 1293 6847 1307
rect 6773 1273 6787 1287
rect 6753 1193 6767 1207
rect 6653 613 6667 627
rect 6733 613 6747 627
rect 6533 333 6547 347
rect 6553 333 6567 347
rect 6593 593 6607 607
rect 6633 593 6647 607
rect 6733 453 6747 467
rect 6673 313 6687 327
rect 6713 293 6727 307
rect 6573 173 6587 187
rect 6913 2033 6927 2047
rect 6993 2253 7007 2267
rect 6953 2133 6967 2147
rect 6993 2113 7007 2127
rect 6953 2093 6967 2107
rect 6933 1813 6947 1827
rect 6953 1793 6967 1807
rect 6893 1773 6907 1787
rect 6933 1753 6947 1767
rect 6893 1633 6907 1647
rect 6913 1593 6927 1607
rect 6973 1733 6987 1747
rect 6993 1713 7007 1727
rect 7033 2313 7047 2327
rect 7133 2313 7147 2327
rect 7093 2293 7107 2307
rect 7073 2253 7087 2267
rect 7113 2253 7127 2267
rect 7033 2233 7047 2247
rect 7153 2133 7167 2147
rect 7033 2113 7047 2127
rect 7053 2073 7067 2087
rect 7073 2033 7087 2047
rect 7073 2013 7087 2027
rect 7033 1813 7047 1827
rect 6913 1373 6927 1387
rect 6853 1193 6867 1207
rect 6813 1153 6827 1167
rect 6873 1153 6887 1167
rect 6833 1113 6847 1127
rect 6893 1113 6907 1127
rect 6813 1073 6827 1087
rect 6853 1073 6867 1087
rect 6833 933 6847 947
rect 6773 813 6787 827
rect 6793 813 6807 827
rect 6813 793 6827 807
rect 6853 793 6867 807
rect 6993 1633 7007 1647
rect 7093 1793 7107 1807
rect 7133 2073 7147 2087
rect 7333 2873 7347 2887
rect 7673 3533 7687 3547
rect 7393 3513 7407 3527
rect 7733 3473 7747 3487
rect 7553 3253 7567 3267
rect 7593 3253 7607 3267
rect 7633 3253 7647 3267
rect 7373 3213 7387 3227
rect 7393 3213 7407 3227
rect 7453 3213 7467 3227
rect 7433 3193 7447 3207
rect 7413 3173 7427 3187
rect 7433 3073 7447 3087
rect 7413 3053 7427 3067
rect 7393 3033 7407 3047
rect 7413 2993 7427 3007
rect 7453 2993 7467 3007
rect 7513 2993 7527 3007
rect 7433 2893 7447 2907
rect 7413 2853 7427 2867
rect 7353 2753 7367 2767
rect 7393 2753 7407 2767
rect 7313 2733 7327 2747
rect 7333 2713 7347 2727
rect 7373 2633 7387 2647
rect 7293 2553 7307 2567
rect 7253 2533 7267 2547
rect 7273 2533 7287 2547
rect 7353 2533 7367 2547
rect 7233 2453 7247 2467
rect 7213 2373 7227 2387
rect 7193 2233 7207 2247
rect 7593 3213 7607 3227
rect 7573 3193 7587 3207
rect 7553 2933 7567 2947
rect 7513 2813 7527 2827
rect 7533 2713 7547 2727
rect 7433 2613 7447 2627
rect 7613 3173 7627 3187
rect 7673 3213 7687 3227
rect 7653 3133 7667 3147
rect 7633 3033 7647 3047
rect 7653 3033 7667 3047
rect 7613 2993 7627 3007
rect 7593 2753 7607 2767
rect 7573 2733 7587 2747
rect 7553 2573 7567 2587
rect 7453 2533 7467 2547
rect 7533 2533 7547 2547
rect 7293 2493 7307 2507
rect 7273 2333 7287 2347
rect 7373 2513 7387 2527
rect 7433 2513 7447 2527
rect 7393 2433 7407 2447
rect 7433 2433 7447 2447
rect 7333 2373 7347 2387
rect 7373 2313 7387 2327
rect 7293 2293 7307 2307
rect 7313 2293 7327 2307
rect 7373 2293 7387 2307
rect 7273 2273 7287 2287
rect 7253 2253 7267 2267
rect 7233 2093 7247 2107
rect 7293 2233 7307 2247
rect 7333 2153 7347 2167
rect 7373 2153 7387 2167
rect 7333 2133 7347 2147
rect 7233 2073 7247 2087
rect 7213 2053 7227 2067
rect 7173 2033 7187 2047
rect 7233 2033 7247 2047
rect 7133 2013 7147 2027
rect 7193 1973 7207 1987
rect 7153 1813 7167 1827
rect 7213 1833 7227 1847
rect 7133 1793 7147 1807
rect 7073 1593 7087 1607
rect 7053 1573 7067 1587
rect 7093 1573 7107 1587
rect 6953 1293 6967 1307
rect 6973 1293 6987 1307
rect 7013 1293 7027 1307
rect 7033 1273 7047 1287
rect 7013 1193 7027 1207
rect 7153 1773 7167 1787
rect 7213 1773 7227 1787
rect 7173 1653 7187 1667
rect 7313 1833 7327 1847
rect 7293 1753 7307 1767
rect 7213 1613 7227 1627
rect 7273 1613 7287 1627
rect 7213 1573 7227 1587
rect 7193 1553 7207 1567
rect 7293 1593 7307 1607
rect 7293 1553 7307 1567
rect 7233 1533 7247 1547
rect 7153 1473 7167 1487
rect 7093 1133 7107 1147
rect 7133 1133 7147 1147
rect 7053 1113 7067 1127
rect 7033 1093 7047 1107
rect 7073 1093 7087 1107
rect 7113 1073 7127 1087
rect 7013 833 7027 847
rect 7053 833 7067 847
rect 7033 793 7047 807
rect 6993 773 7007 787
rect 7053 753 7067 767
rect 6913 733 6927 747
rect 6853 713 6867 727
rect 6913 713 6927 727
rect 6833 653 6847 667
rect 6753 373 6767 387
rect 6813 613 6827 627
rect 6793 593 6807 607
rect 6873 633 6887 647
rect 6873 593 6887 607
rect 6853 373 6867 387
rect 6893 373 6907 387
rect 6773 353 6787 367
rect 6833 353 6847 367
rect 6873 313 6887 327
rect 7013 653 7027 667
rect 6973 613 6987 627
rect 6993 613 7007 627
rect 6913 273 6927 287
rect 7033 593 7047 607
rect 7053 393 7067 407
rect 7073 353 7087 367
rect 7013 293 7027 307
rect 6973 213 6987 227
rect 7073 273 7087 287
rect 7113 353 7127 367
rect 7113 333 7127 347
rect 7093 253 7107 267
rect 7073 173 7087 187
rect 7133 173 7147 187
rect 6113 13 6127 27
rect 6153 13 6167 27
rect 7053 153 7067 167
rect 7033 133 7047 147
rect 7273 1493 7287 1507
rect 7253 1473 7267 1487
rect 7233 1413 7247 1427
rect 7233 1333 7247 1347
rect 7193 1313 7207 1327
rect 7173 1293 7187 1307
rect 7253 1293 7267 1307
rect 7233 1253 7247 1267
rect 7273 1233 7287 1247
rect 7213 1153 7227 1167
rect 7233 1153 7247 1167
rect 7273 1113 7287 1127
rect 7173 1013 7187 1027
rect 7193 833 7207 847
rect 7173 733 7187 747
rect 7513 2513 7527 2527
rect 7553 2513 7567 2527
rect 7593 2713 7607 2727
rect 7533 2473 7547 2487
rect 7573 2473 7587 2487
rect 7513 2453 7527 2467
rect 7493 2273 7507 2287
rect 7573 2413 7587 2427
rect 7513 2253 7527 2267
rect 7593 2333 7607 2347
rect 7473 2233 7487 2247
rect 7453 2193 7467 2207
rect 7513 2153 7527 2167
rect 7493 2133 7507 2147
rect 7473 2093 7487 2107
rect 7413 2073 7427 2087
rect 7453 2073 7467 2087
rect 7393 1993 7407 2007
rect 7473 2013 7487 2027
rect 7493 1993 7507 2007
rect 7433 1913 7447 1927
rect 7393 1873 7407 1887
rect 7333 1773 7347 1787
rect 7333 1573 7347 1587
rect 7373 1773 7387 1787
rect 7433 1813 7447 1827
rect 7433 1753 7447 1767
rect 7413 1673 7427 1687
rect 7393 1593 7407 1607
rect 7393 1573 7407 1587
rect 7353 1533 7367 1547
rect 7493 1593 7507 1607
rect 7453 1573 7467 1587
rect 7473 1573 7487 1587
rect 7653 2893 7667 2907
rect 7633 2773 7647 2787
rect 7633 2573 7647 2587
rect 7733 3033 7747 3047
rect 7833 3853 7847 3867
rect 7873 4453 7887 4467
rect 8053 4613 8067 4627
rect 8033 4493 8047 4507
rect 8133 4973 8147 4987
rect 8113 4953 8127 4967
rect 8153 4933 8167 4947
rect 8113 4773 8127 4787
rect 8093 4673 8107 4687
rect 8073 4393 8087 4407
rect 8013 4233 8027 4247
rect 7873 4193 7887 4207
rect 8033 4153 8047 4167
rect 8013 4133 8027 4147
rect 8133 4753 8147 4767
rect 8213 4933 8227 4947
rect 8353 5773 8367 5787
rect 8373 5753 8387 5767
rect 8333 5593 8347 5607
rect 8313 5453 8327 5467
rect 8293 5413 8307 5427
rect 8313 5373 8327 5387
rect 8293 5273 8307 5287
rect 8273 5173 8287 5187
rect 8273 5113 8287 5127
rect 8253 4993 8267 5007
rect 8253 4953 8267 4967
rect 8173 4713 8187 4727
rect 8193 4713 8207 4727
rect 8153 4673 8167 4687
rect 8253 4673 8267 4687
rect 8193 4573 8207 4587
rect 8233 4473 8247 4487
rect 8213 4433 8227 4447
rect 8173 4233 8187 4247
rect 8393 5613 8407 5627
rect 8393 5393 8407 5407
rect 8393 5133 8407 5147
rect 8373 5113 8387 5127
rect 8333 5073 8347 5087
rect 8293 5013 8307 5027
rect 8593 6033 8607 6047
rect 8653 6113 8667 6127
rect 8533 5873 8547 5887
rect 8553 5873 8567 5887
rect 8493 5653 8507 5667
rect 8473 5453 8487 5467
rect 8513 5613 8527 5627
rect 8453 5393 8467 5407
rect 8493 5193 8507 5207
rect 8433 5133 8447 5147
rect 8433 5073 8447 5087
rect 8373 4953 8387 4967
rect 8313 4933 8327 4947
rect 8373 4913 8387 4927
rect 8413 4933 8427 4947
rect 8453 4993 8467 5007
rect 8413 4853 8427 4867
rect 8433 4853 8447 4867
rect 8313 4693 8327 4707
rect 8393 4693 8407 4707
rect 8313 4513 8327 4527
rect 8273 4273 8287 4287
rect 8133 4193 8147 4207
rect 8213 4193 8227 4207
rect 8373 4673 8387 4687
rect 8353 4493 8367 4507
rect 8393 4493 8407 4507
rect 8333 4453 8347 4467
rect 8433 4613 8447 4627
rect 8373 4473 8387 4487
rect 8413 4473 8427 4487
rect 8493 4993 8507 5007
rect 8473 4953 8487 4967
rect 8553 5813 8567 5827
rect 8573 5653 8587 5667
rect 8593 5633 8607 5647
rect 8633 5993 8647 6007
rect 8553 5613 8567 5627
rect 8533 5173 8547 5187
rect 8613 5613 8627 5627
rect 8653 5893 8667 5907
rect 8633 5573 8647 5587
rect 8573 5453 8587 5467
rect 8993 7333 9007 7347
rect 9193 7873 9207 7887
rect 9173 7613 9187 7627
rect 9193 7593 9207 7607
rect 9153 7573 9167 7587
rect 9193 7553 9207 7567
rect 9213 7553 9227 7567
rect 9113 7493 9127 7507
rect 9133 7453 9147 7467
rect 9173 7373 9187 7387
rect 9113 7333 9127 7347
rect 9153 7333 9167 7347
rect 9073 7313 9087 7327
rect 9033 7113 9047 7127
rect 9013 6913 9027 6927
rect 9133 7113 9147 7127
rect 9093 7093 9107 7107
rect 9073 7073 9087 7087
rect 9113 7073 9127 7087
rect 9193 7073 9207 7087
rect 9273 7993 9287 8007
rect 9273 7973 9287 7987
rect 9253 7833 9267 7847
rect 9453 8433 9467 8447
rect 9533 11173 9547 11187
rect 9553 11173 9567 11187
rect 9573 10973 9587 10987
rect 9553 10953 9567 10967
rect 9513 10933 9527 10947
rect 9533 10913 9547 10927
rect 9513 10793 9527 10807
rect 9533 10733 9547 10747
rect 9553 10713 9567 10727
rect 9493 10553 9507 10567
rect 9533 10553 9547 10567
rect 9493 10453 9507 10467
rect 9513 10413 9527 10427
rect 9493 10273 9507 10287
rect 9493 10153 9507 10167
rect 9573 10253 9587 10267
rect 9553 10233 9567 10247
rect 9533 10073 9547 10087
rect 9573 10073 9587 10087
rect 9493 9953 9507 9967
rect 9553 9973 9567 9987
rect 9533 9953 9547 9967
rect 9693 11373 9707 11387
rect 10313 11833 10327 11847
rect 10313 11773 10327 11787
rect 10373 11773 10387 11787
rect 10013 11693 10027 11707
rect 9993 11673 10007 11687
rect 10033 11673 10047 11687
rect 10133 11693 10147 11707
rect 10273 11673 10287 11687
rect 10293 11673 10307 11687
rect 10113 11633 10127 11647
rect 10153 11633 10167 11647
rect 10273 11633 10287 11647
rect 10333 11653 10347 11667
rect 10353 11653 10367 11667
rect 10393 11653 10407 11667
rect 10313 11633 10327 11647
rect 10293 11573 10307 11587
rect 9933 11473 9947 11487
rect 9853 11373 9867 11387
rect 9873 11373 9887 11387
rect 9733 11293 9747 11307
rect 9833 11293 9847 11307
rect 9653 11113 9667 11127
rect 9673 10933 9687 10947
rect 9913 11233 9927 11247
rect 9953 11213 9967 11227
rect 9913 11193 9927 11207
rect 9893 11033 9907 11047
rect 9933 11013 9947 11027
rect 9853 10913 9867 10927
rect 9733 10893 9747 10907
rect 9913 10913 9927 10927
rect 9973 10913 9987 10927
rect 9713 10733 9727 10747
rect 9873 10733 9887 10747
rect 9913 10733 9927 10747
rect 9933 10733 9947 10747
rect 9713 10713 9727 10727
rect 9753 10713 9767 10727
rect 9893 10713 9907 10727
rect 9693 10673 9707 10687
rect 9733 10673 9747 10687
rect 9713 10513 9727 10527
rect 9653 10373 9667 10387
rect 9693 10433 9707 10447
rect 9693 10413 9707 10427
rect 9673 10273 9687 10287
rect 9733 10273 9747 10287
rect 9653 10233 9667 10247
rect 9673 10233 9687 10247
rect 10253 11433 10267 11447
rect 10013 11413 10027 11427
rect 10033 11373 10047 11387
rect 10213 11373 10227 11387
rect 10073 11353 10087 11367
rect 10013 11293 10027 11307
rect 9993 10513 10007 10527
rect 9853 10393 9867 10407
rect 9893 10433 9907 10447
rect 9953 10393 9967 10407
rect 9873 10373 9887 10387
rect 9853 10353 9867 10367
rect 9833 10253 9847 10267
rect 9693 10173 9707 10187
rect 9653 10073 9667 10087
rect 9613 9913 9627 9927
rect 9613 9773 9627 9787
rect 9513 9553 9527 9567
rect 9553 9553 9567 9567
rect 9513 9533 9527 9547
rect 9493 9473 9507 9487
rect 9513 9233 9527 9247
rect 9533 9093 9547 9107
rect 9573 9513 9587 9527
rect 9653 9733 9667 9747
rect 9633 9633 9647 9647
rect 9653 9453 9667 9467
rect 9593 9433 9607 9447
rect 9613 9433 9627 9447
rect 9653 9293 9667 9307
rect 9573 9253 9587 9267
rect 9613 9253 9627 9267
rect 9573 9213 9587 9227
rect 9593 9193 9607 9207
rect 9593 9133 9607 9147
rect 9553 9073 9567 9087
rect 9553 8933 9567 8947
rect 9553 8873 9567 8887
rect 9493 8613 9507 8627
rect 9573 8853 9587 8867
rect 9613 9013 9627 9027
rect 9613 8933 9627 8947
rect 9613 8893 9627 8907
rect 9593 8773 9607 8787
rect 9573 8753 9587 8767
rect 9713 9933 9727 9947
rect 9753 9913 9767 9927
rect 9813 10133 9827 10147
rect 9833 10053 9847 10067
rect 9833 9933 9847 9947
rect 9873 10213 9887 10227
rect 9993 10273 10007 10287
rect 9873 10033 9887 10047
rect 9973 10173 9987 10187
rect 10053 11213 10067 11227
rect 10533 11793 10547 11807
rect 10573 11793 10587 11807
rect 10493 11653 10507 11667
rect 10453 11633 10467 11647
rect 10513 11633 10527 11647
rect 10413 11573 10427 11587
rect 10413 11553 10427 11567
rect 10393 11413 10407 11427
rect 10533 11573 10547 11587
rect 10453 11473 10467 11487
rect 10453 11413 10467 11427
rect 10453 11313 10467 11327
rect 10893 11893 10907 11907
rect 10653 11873 10667 11887
rect 10613 11613 10627 11627
rect 10713 11813 10727 11827
rect 10693 11753 10707 11767
rect 10673 11673 10687 11687
rect 10733 11673 10747 11687
rect 10713 11613 10727 11627
rect 10653 11593 10667 11607
rect 10653 11453 10667 11467
rect 10573 11413 10587 11427
rect 10613 11413 10627 11427
rect 10593 11393 10607 11407
rect 10553 11353 10567 11367
rect 10193 11193 10207 11207
rect 10313 11193 10327 11207
rect 10093 11173 10107 11187
rect 10133 11173 10147 11187
rect 10053 11153 10067 11167
rect 10113 11153 10127 11167
rect 10133 11113 10147 11127
rect 10313 10973 10327 10987
rect 10033 10733 10047 10747
rect 10053 10673 10067 10687
rect 10073 10533 10087 10547
rect 10113 10933 10127 10947
rect 10173 10933 10187 10947
rect 10193 10933 10207 10947
rect 10273 10933 10287 10947
rect 10133 10893 10147 10907
rect 10173 10873 10187 10887
rect 10173 10753 10187 10767
rect 10153 10713 10167 10727
rect 10113 10493 10127 10507
rect 10093 10453 10107 10467
rect 10053 10393 10067 10407
rect 10073 10393 10087 10407
rect 10113 10413 10127 10427
rect 10153 10313 10167 10327
rect 10133 10253 10147 10267
rect 10073 10233 10087 10247
rect 9933 9993 9947 10007
rect 9933 9933 9947 9947
rect 9853 9913 9867 9927
rect 9913 9913 9927 9927
rect 9813 9873 9827 9887
rect 9733 9853 9747 9867
rect 9773 9853 9787 9867
rect 9873 9853 9887 9867
rect 9773 9813 9787 9827
rect 9793 9753 9807 9767
rect 9733 9533 9747 9547
rect 9713 9453 9727 9467
rect 9733 9433 9747 9447
rect 9753 9313 9767 9327
rect 9713 9253 9727 9267
rect 9693 9093 9707 9107
rect 9713 8993 9727 9007
rect 9673 8873 9687 8887
rect 9673 8813 9687 8827
rect 9633 8793 9647 8807
rect 9693 8773 9707 8787
rect 9573 8613 9587 8627
rect 9473 8393 9487 8407
rect 9373 8373 9387 8387
rect 9353 8313 9367 8327
rect 9393 8313 9407 8327
rect 9433 8313 9447 8327
rect 9333 8293 9347 8307
rect 9313 7873 9327 7887
rect 9293 7853 9307 7867
rect 9313 7833 9327 7847
rect 9273 7813 9287 7827
rect 9253 7573 9267 7587
rect 9233 7533 9247 7547
rect 9333 7813 9347 7827
rect 9373 8293 9387 8307
rect 9513 8493 9527 8507
rect 9513 8293 9527 8307
rect 9493 8233 9507 8247
rect 9413 8193 9427 8207
rect 9453 8193 9467 8207
rect 9493 8093 9507 8107
rect 9413 8013 9427 8027
rect 9513 8033 9527 8047
rect 9433 7973 9447 7987
rect 9413 7873 9427 7887
rect 9393 7813 9407 7827
rect 9433 7753 9447 7767
rect 9413 7733 9427 7747
rect 9353 7713 9367 7727
rect 9353 7613 9367 7627
rect 9393 7553 9407 7567
rect 9373 7513 9387 7527
rect 9313 7373 9327 7387
rect 9253 7333 9267 7347
rect 9233 7213 9247 7227
rect 9333 7353 9347 7367
rect 9353 7333 9367 7347
rect 9313 7313 9327 7327
rect 9333 7293 9347 7307
rect 9273 7193 9287 7207
rect 9273 7073 9287 7087
rect 9333 7073 9347 7087
rect 9213 6993 9227 7007
rect 9193 6953 9207 6967
rect 9113 6873 9127 6887
rect 9233 6913 9247 6927
rect 9213 6893 9227 6907
rect 9013 6833 9027 6847
rect 8993 6793 9007 6807
rect 8973 6773 8987 6787
rect 9053 6773 9067 6787
rect 9033 6633 9047 6647
rect 8833 6593 8847 6607
rect 8853 6593 8867 6607
rect 8793 6573 8807 6587
rect 8853 6513 8867 6527
rect 9073 6593 9087 6607
rect 9013 6573 9027 6587
rect 9273 6753 9287 6767
rect 9233 6613 9247 6627
rect 9313 7053 9327 7067
rect 9333 6893 9347 6907
rect 9293 6713 9307 6727
rect 9293 6613 9307 6627
rect 9253 6593 9267 6607
rect 8913 6493 8927 6507
rect 8993 6493 9007 6507
rect 8873 6453 8887 6467
rect 8833 6433 8847 6447
rect 8793 6393 8807 6407
rect 8853 6393 8867 6407
rect 8773 6373 8787 6387
rect 8753 6353 8767 6367
rect 8793 6353 8807 6367
rect 8813 6353 8827 6367
rect 8753 6113 8767 6127
rect 8733 5993 8747 6007
rect 8733 5953 8747 5967
rect 8773 5933 8787 5947
rect 8713 5893 8727 5907
rect 8753 5893 8767 5907
rect 8673 5873 8687 5887
rect 8733 5613 8747 5627
rect 8693 5593 8707 5607
rect 8753 5593 8767 5607
rect 8693 5573 8707 5587
rect 8733 5573 8747 5587
rect 8673 5393 8687 5407
rect 8633 5293 8647 5307
rect 8593 5193 8607 5207
rect 8633 5173 8647 5187
rect 8613 5153 8627 5167
rect 8553 5073 8567 5087
rect 8673 4973 8687 4987
rect 8833 6333 8847 6347
rect 8893 6393 8907 6407
rect 8873 6333 8887 6347
rect 8893 6153 8907 6167
rect 8953 6393 8967 6407
rect 9073 6413 9087 6427
rect 8973 6373 8987 6387
rect 9013 6373 9027 6387
rect 8933 6133 8947 6147
rect 8913 6113 8927 6127
rect 8873 5933 8887 5947
rect 8993 6113 9007 6127
rect 9053 6133 9067 6147
rect 9033 6033 9047 6047
rect 9013 6013 9027 6027
rect 8953 5913 8967 5927
rect 8993 5913 9007 5927
rect 8973 5893 8987 5907
rect 9013 5893 9027 5907
rect 9053 5893 9067 5907
rect 8833 5793 8847 5807
rect 8953 5773 8967 5787
rect 8913 5633 8927 5647
rect 8993 5653 9007 5667
rect 8893 5613 8907 5627
rect 8793 5573 8807 5587
rect 8853 5473 8867 5487
rect 8753 5413 8767 5427
rect 8833 5433 8847 5447
rect 8813 5413 8827 5427
rect 8973 5613 8987 5627
rect 8933 5413 8947 5427
rect 8993 5433 9007 5447
rect 9033 5433 9047 5447
rect 9013 5413 9027 5427
rect 8973 5393 8987 5407
rect 8773 5293 8787 5307
rect 8933 5213 8947 5227
rect 8873 5173 8887 5187
rect 8793 5153 8807 5167
rect 8833 5153 8847 5167
rect 8893 5153 8907 5167
rect 8733 5053 8747 5067
rect 8813 4973 8827 4987
rect 8693 4953 8707 4967
rect 8533 4913 8547 4927
rect 8833 4913 8847 4927
rect 8853 4913 8867 4927
rect 8853 4853 8867 4867
rect 8513 4773 8527 4787
rect 8733 4773 8747 4787
rect 8473 4693 8487 4707
rect 8533 4693 8547 4707
rect 8513 4673 8527 4687
rect 8693 4673 8707 4687
rect 8773 4693 8787 4707
rect 8493 4613 8507 4627
rect 8473 4533 8487 4547
rect 8453 4513 8467 4527
rect 8453 4273 8467 4287
rect 8393 4253 8407 4267
rect 8353 4213 8367 4227
rect 8373 4093 8387 4107
rect 8153 4013 8167 4027
rect 8393 4013 8407 4027
rect 8133 3993 8147 4007
rect 8193 3993 8207 4007
rect 8013 3973 8027 3987
rect 8113 3973 8127 3987
rect 7993 3953 8007 3967
rect 7873 3933 7887 3947
rect 8033 3933 8047 3947
rect 7793 3753 7807 3767
rect 7793 3733 7807 3747
rect 7813 3693 7827 3707
rect 7773 3653 7787 3667
rect 7813 3653 7827 3667
rect 7773 3573 7787 3587
rect 8013 3893 8027 3907
rect 7933 3853 7947 3867
rect 7893 3713 7907 3727
rect 7873 3553 7887 3567
rect 7853 3533 7867 3547
rect 7873 3513 7887 3527
rect 7893 3513 7907 3527
rect 7833 3493 7847 3507
rect 7773 3453 7787 3467
rect 7793 3253 7807 3267
rect 7833 3253 7847 3267
rect 7913 3473 7927 3487
rect 7893 3453 7907 3467
rect 7753 2993 7767 3007
rect 7733 2833 7747 2847
rect 7873 3093 7887 3107
rect 7893 3053 7907 3067
rect 7813 3013 7827 3027
rect 7793 2813 7807 2827
rect 7773 2793 7787 2807
rect 7693 2753 7707 2767
rect 7733 2753 7747 2767
rect 7773 2753 7787 2767
rect 7753 2733 7767 2747
rect 7673 2633 7687 2647
rect 7713 2573 7727 2587
rect 7793 2733 7807 2747
rect 7813 2733 7827 2747
rect 7773 2693 7787 2707
rect 7793 2573 7807 2587
rect 7733 2533 7747 2547
rect 7693 2473 7707 2487
rect 7713 2393 7727 2407
rect 7693 2153 7707 2167
rect 7553 2033 7567 2047
rect 7573 2033 7587 2047
rect 7653 2113 7667 2127
rect 7613 2093 7627 2107
rect 7653 2073 7667 2087
rect 7713 2113 7727 2127
rect 7633 2053 7647 2067
rect 7613 2033 7627 2047
rect 7593 2013 7607 2027
rect 7553 1993 7567 2007
rect 7573 1893 7587 1907
rect 7533 1773 7547 1787
rect 7553 1753 7567 1767
rect 7573 1733 7587 1747
rect 7513 1473 7527 1487
rect 7453 1453 7467 1467
rect 7473 1453 7487 1467
rect 7393 1393 7407 1407
rect 7473 1433 7487 1447
rect 7453 1373 7467 1387
rect 7453 1353 7467 1367
rect 7413 1333 7427 1347
rect 7333 1253 7347 1267
rect 7373 1193 7387 1207
rect 7333 1113 7347 1127
rect 7313 833 7327 847
rect 7353 1053 7367 1067
rect 7333 813 7347 827
rect 7433 1293 7447 1307
rect 7433 1273 7447 1287
rect 7413 1253 7427 1267
rect 7393 1173 7407 1187
rect 7393 1093 7407 1107
rect 7373 873 7387 887
rect 7453 1173 7467 1187
rect 7493 1393 7507 1407
rect 7673 1993 7687 2007
rect 7673 1933 7687 1947
rect 7613 1733 7627 1747
rect 7593 1673 7607 1687
rect 7613 1653 7627 1667
rect 7593 1593 7607 1607
rect 7533 1333 7547 1347
rect 7513 1293 7527 1307
rect 7493 1273 7507 1287
rect 7493 1113 7507 1127
rect 7513 1093 7527 1107
rect 7453 1053 7467 1067
rect 7493 973 7507 987
rect 7533 973 7547 987
rect 7413 953 7427 967
rect 7473 873 7487 887
rect 7433 833 7447 847
rect 7373 813 7387 827
rect 7353 793 7367 807
rect 7453 813 7467 827
rect 7253 753 7267 767
rect 7413 753 7427 767
rect 7253 713 7267 727
rect 7453 713 7467 727
rect 7433 653 7447 667
rect 7373 633 7387 647
rect 7233 613 7247 627
rect 7393 613 7407 627
rect 7413 613 7427 627
rect 7173 593 7187 607
rect 7213 593 7227 607
rect 7393 573 7407 587
rect 7413 453 7427 467
rect 7293 373 7307 387
rect 7233 313 7247 327
rect 7253 233 7267 247
rect 7233 153 7247 167
rect 7133 133 7147 147
rect 7153 133 7167 147
rect 7213 133 7227 147
rect 7313 293 7327 307
rect 7533 953 7547 967
rect 7513 853 7527 867
rect 7493 813 7507 827
rect 7513 753 7527 767
rect 7833 2553 7847 2567
rect 7913 2893 7927 2907
rect 7973 3713 7987 3727
rect 8073 3733 8087 3747
rect 7953 3613 7967 3627
rect 7993 3613 8007 3627
rect 8173 3973 8187 3987
rect 8153 3733 8167 3747
rect 8133 3713 8147 3727
rect 8173 3713 8187 3727
rect 8213 3693 8227 3707
rect 8193 3633 8207 3647
rect 8373 3973 8387 3987
rect 8433 3973 8447 3987
rect 8473 3973 8487 3987
rect 8293 3753 8307 3767
rect 8233 3613 8247 3627
rect 8213 3573 8227 3587
rect 8093 3553 8107 3567
rect 8273 3533 8287 3547
rect 8353 3713 8367 3727
rect 8333 3533 8347 3547
rect 8113 3513 8127 3527
rect 8133 3513 8147 3527
rect 8053 3413 8067 3427
rect 8133 3413 8147 3427
rect 7993 3373 8007 3387
rect 7953 3293 7967 3307
rect 8293 3513 8307 3527
rect 8333 3333 8347 3347
rect 8153 3273 8167 3287
rect 8233 3273 8247 3287
rect 7993 3233 8007 3247
rect 8033 3233 8047 3247
rect 8093 3233 8107 3247
rect 8013 3213 8027 3227
rect 8033 3193 8047 3207
rect 8093 3073 8107 3087
rect 8073 3033 8087 3047
rect 8013 3013 8027 3027
rect 8013 2913 8027 2927
rect 8013 2853 8027 2867
rect 7893 2793 7907 2807
rect 7933 2793 7947 2807
rect 7993 2793 8007 2807
rect 7913 2773 7927 2787
rect 7813 2513 7827 2527
rect 7753 2253 7767 2267
rect 7793 2253 7807 2267
rect 7773 2113 7787 2127
rect 7733 2033 7747 2047
rect 8013 2773 8027 2787
rect 8033 2753 8047 2767
rect 8093 2933 8107 2947
rect 8093 2853 8107 2867
rect 8093 2833 8107 2847
rect 7993 2733 8007 2747
rect 7953 2693 7967 2707
rect 7873 2533 7887 2547
rect 7893 2533 7907 2547
rect 7853 2393 7867 2407
rect 7873 2293 7887 2307
rect 7933 2533 7947 2547
rect 7953 2533 7967 2547
rect 7913 2513 7927 2527
rect 7993 2513 8007 2527
rect 7973 2493 7987 2507
rect 7973 2353 7987 2367
rect 7933 2313 7947 2327
rect 7913 2253 7927 2267
rect 7893 2233 7907 2247
rect 7933 2233 7947 2247
rect 7873 2213 7887 2227
rect 7873 2113 7887 2127
rect 7793 2053 7807 2067
rect 7773 1993 7787 2007
rect 7733 1973 7747 1987
rect 7793 1973 7807 1987
rect 7713 1873 7727 1887
rect 7733 1873 7747 1887
rect 7853 2093 7867 2107
rect 7833 2073 7847 2087
rect 7913 2073 7927 2087
rect 7853 2053 7867 2067
rect 7893 2053 7907 2067
rect 7853 2013 7867 2027
rect 7833 1993 7847 2007
rect 7813 1813 7827 1827
rect 7713 1773 7727 1787
rect 7753 1773 7767 1787
rect 7793 1773 7807 1787
rect 7713 1753 7727 1767
rect 7673 1633 7687 1647
rect 7653 1593 7667 1607
rect 7693 1593 7707 1607
rect 7673 1473 7687 1487
rect 7693 1373 7707 1387
rect 7613 1313 7627 1327
rect 7573 1293 7587 1307
rect 7593 1273 7607 1287
rect 7693 1273 7707 1287
rect 7633 1193 7647 1207
rect 7753 1733 7767 1747
rect 7733 1593 7747 1607
rect 7733 1553 7747 1567
rect 7773 1573 7787 1587
rect 7733 1513 7747 1527
rect 7753 1513 7767 1527
rect 7773 1453 7787 1467
rect 7833 1733 7847 1747
rect 7953 2213 7967 2227
rect 7893 1993 7907 2007
rect 7933 1993 7947 2007
rect 7873 1853 7887 1867
rect 7873 1773 7887 1787
rect 7933 1853 7947 1867
rect 7973 2053 7987 2067
rect 8173 3233 8187 3247
rect 8213 3233 8227 3247
rect 8233 3213 8247 3227
rect 8193 3193 8207 3207
rect 8213 3113 8227 3127
rect 8253 3053 8267 3067
rect 8453 3633 8467 3647
rect 8393 3613 8407 3627
rect 8413 3513 8427 3527
rect 8473 3533 8487 3547
rect 8433 3473 8447 3487
rect 8373 3253 8387 3267
rect 8393 3233 8407 3247
rect 8433 3233 8447 3247
rect 8373 3193 8387 3207
rect 8353 3053 8367 3067
rect 8333 3013 8347 3027
rect 8233 2793 8247 2807
rect 8153 2733 8167 2747
rect 8133 2713 8147 2727
rect 8053 2693 8067 2707
rect 8073 2693 8087 2707
rect 8073 2573 8087 2587
rect 8033 2173 8047 2187
rect 8013 2133 8027 2147
rect 7993 1993 8007 2007
rect 7993 1893 8007 1907
rect 7953 1833 7967 1847
rect 7973 1793 7987 1807
rect 7893 1733 7907 1747
rect 7853 1653 7867 1667
rect 7953 1773 7967 1787
rect 7933 1733 7947 1747
rect 7913 1673 7927 1687
rect 7893 1593 7907 1607
rect 7833 1573 7847 1587
rect 7873 1573 7887 1587
rect 7853 1553 7867 1567
rect 7873 1553 7887 1567
rect 7793 1393 7807 1407
rect 7773 1333 7787 1347
rect 7853 1453 7867 1467
rect 7753 1293 7767 1307
rect 7853 1293 7867 1307
rect 7793 1273 7807 1287
rect 7853 1273 7867 1287
rect 7793 1233 7807 1247
rect 7733 1173 7747 1187
rect 7713 1133 7727 1147
rect 7673 1113 7687 1127
rect 7753 1133 7767 1147
rect 7773 1133 7787 1147
rect 7693 1093 7707 1107
rect 7633 873 7647 887
rect 7553 793 7567 807
rect 7553 673 7567 687
rect 7533 653 7547 667
rect 7613 773 7627 787
rect 7593 713 7607 727
rect 7653 793 7667 807
rect 7633 713 7647 727
rect 7613 673 7627 687
rect 7633 653 7647 667
rect 7573 633 7587 647
rect 7613 613 7627 627
rect 7473 393 7487 407
rect 7613 393 7627 407
rect 7493 333 7507 347
rect 7533 333 7547 347
rect 7453 253 7467 267
rect 7473 133 7487 147
rect 7733 1033 7747 1047
rect 7713 913 7727 927
rect 7773 1093 7787 1107
rect 7833 1173 7847 1187
rect 7893 1513 7907 1527
rect 7993 1673 8007 1687
rect 7953 1593 7967 1607
rect 7933 1513 7947 1527
rect 7913 1433 7927 1447
rect 7933 1433 7947 1447
rect 7893 1333 7907 1347
rect 7913 1293 7927 1307
rect 7893 1253 7907 1267
rect 7873 1233 7887 1247
rect 7913 1173 7927 1187
rect 7913 1133 7927 1147
rect 7873 1113 7887 1127
rect 7893 993 7907 1007
rect 7833 893 7847 907
rect 7793 833 7807 847
rect 7893 833 7907 847
rect 7813 813 7827 827
rect 7833 713 7847 727
rect 7733 673 7747 687
rect 7773 673 7787 687
rect 7713 653 7727 667
rect 7693 633 7707 647
rect 7653 613 7667 627
rect 7813 653 7827 667
rect 7773 633 7787 647
rect 7893 793 7907 807
rect 8253 2753 8267 2767
rect 8293 2753 8307 2767
rect 8193 2613 8207 2627
rect 8313 2733 8327 2747
rect 8273 2713 8287 2727
rect 8253 2593 8267 2607
rect 8233 2573 8247 2587
rect 8213 2473 8227 2487
rect 8193 2453 8207 2467
rect 8173 2313 8187 2327
rect 8153 2273 8167 2287
rect 8113 2253 8127 2267
rect 8093 2193 8107 2207
rect 8073 2113 8087 2127
rect 8033 2073 8047 2087
rect 8093 2093 8107 2107
rect 8053 2013 8067 2027
rect 8173 2253 8187 2267
rect 8193 2253 8207 2267
rect 8133 2233 8147 2247
rect 8193 2233 8207 2247
rect 8153 2113 8167 2127
rect 8173 2113 8187 2127
rect 8133 2093 8147 2107
rect 8133 2033 8147 2047
rect 8173 2033 8187 2047
rect 8153 1933 8167 1947
rect 8133 1893 8147 1907
rect 8153 1873 8167 1887
rect 8113 1853 8127 1867
rect 8073 1813 8087 1827
rect 8093 1813 8107 1827
rect 8073 1733 8087 1747
rect 8053 1573 8067 1587
rect 8013 1553 8027 1567
rect 8033 1533 8047 1547
rect 8073 1513 8087 1527
rect 8053 1453 8067 1467
rect 7973 1393 7987 1407
rect 8013 1373 8027 1387
rect 7953 1273 7967 1287
rect 7853 633 7867 647
rect 7873 633 7887 647
rect 7933 633 7947 647
rect 7833 593 7847 607
rect 7853 593 7867 607
rect 7733 553 7747 567
rect 7793 553 7807 567
rect 7733 533 7747 547
rect 7653 493 7667 507
rect 7673 453 7687 467
rect 7653 433 7667 447
rect 7673 393 7687 407
rect 7653 373 7667 387
rect 7713 353 7727 367
rect 7613 313 7627 327
rect 7653 313 7667 327
rect 7733 313 7747 327
rect 7633 293 7647 307
rect 7613 173 7627 187
rect 7533 133 7547 147
rect 7613 133 7627 147
rect 7693 173 7707 187
rect 7653 153 7667 167
rect 7673 133 7687 147
rect 7813 473 7827 487
rect 7833 373 7847 387
rect 7813 333 7827 347
rect 7853 333 7867 347
rect 7813 153 7827 167
rect 7833 153 7847 167
rect 8033 1253 8047 1267
rect 8253 2533 8267 2547
rect 8313 2493 8327 2507
rect 8233 2373 8247 2387
rect 8273 2333 8287 2347
rect 8253 2313 8267 2327
rect 8233 2133 8247 2147
rect 8413 3173 8427 3187
rect 8513 4513 8527 4527
rect 8533 4513 8547 4527
rect 8753 4633 8767 4647
rect 8773 4633 8787 4647
rect 8733 4473 8747 4487
rect 8813 4473 8827 4487
rect 8733 4433 8747 4447
rect 8513 4173 8527 4187
rect 8713 4153 8727 4167
rect 8893 5113 8907 5127
rect 9013 5233 9027 5247
rect 8973 5193 8987 5207
rect 8993 5153 9007 5167
rect 8953 5053 8967 5067
rect 8953 5013 8967 5027
rect 8933 4913 8947 4927
rect 8993 4933 9007 4947
rect 8873 4713 8887 4727
rect 8933 4653 8947 4667
rect 9013 4893 9027 4907
rect 9053 4653 9067 4667
rect 9093 6333 9107 6347
rect 9253 6453 9267 6467
rect 9273 6453 9287 6467
rect 9213 6393 9227 6407
rect 9253 6393 9267 6407
rect 9233 6373 9247 6387
rect 9273 6373 9287 6387
rect 9213 6353 9227 6367
rect 9173 6153 9187 6167
rect 9113 6073 9127 6087
rect 9333 6333 9347 6347
rect 9313 6093 9327 6107
rect 9293 6033 9307 6047
rect 9233 6013 9247 6027
rect 9173 5933 9187 5947
rect 9113 5913 9127 5927
rect 9273 5913 9287 5927
rect 9133 5893 9147 5907
rect 9153 5873 9167 5887
rect 9273 5873 9287 5887
rect 9293 5873 9307 5887
rect 9333 5873 9347 5887
rect 9113 5813 9127 5827
rect 9093 5653 9107 5667
rect 9513 7673 9527 7687
rect 9473 7553 9487 7567
rect 9693 8533 9707 8547
rect 9653 8493 9667 8507
rect 9573 8433 9587 8447
rect 9553 8333 9567 8347
rect 9613 8333 9627 8347
rect 9573 8053 9587 8067
rect 9673 8473 9687 8487
rect 9653 8213 9667 8227
rect 9733 8913 9747 8927
rect 9733 8873 9747 8887
rect 9813 9293 9827 9307
rect 9773 9233 9787 9247
rect 9853 9073 9867 9087
rect 9893 9773 9907 9787
rect 9913 9773 9927 9787
rect 9973 9733 9987 9747
rect 9953 9653 9967 9667
rect 9893 9593 9907 9607
rect 9933 9593 9947 9607
rect 9913 9573 9927 9587
rect 9953 9513 9967 9527
rect 9893 9473 9907 9487
rect 9933 9473 9947 9487
rect 9913 9353 9927 9367
rect 9873 9033 9887 9047
rect 10113 10113 10127 10127
rect 10093 10013 10107 10027
rect 10073 9993 10087 10007
rect 10153 9993 10167 10007
rect 10113 9973 10127 9987
rect 10073 9933 10087 9947
rect 10153 9913 10167 9927
rect 10033 9653 10047 9667
rect 10013 9533 10027 9547
rect 9953 9453 9967 9467
rect 9993 9453 10007 9467
rect 9933 9013 9947 9027
rect 9793 8813 9807 8827
rect 9813 8813 9827 8827
rect 9813 8733 9827 8747
rect 9713 8353 9727 8367
rect 9693 8313 9707 8327
rect 9713 8313 9727 8327
rect 9733 8293 9747 8307
rect 9713 8273 9727 8287
rect 9733 8253 9747 8267
rect 9673 8173 9687 8187
rect 9693 8173 9707 8187
rect 9633 8033 9647 8047
rect 9613 8013 9627 8027
rect 9593 7853 9607 7867
rect 9573 7813 9587 7827
rect 9633 7913 9647 7927
rect 9633 7853 9647 7867
rect 9633 7773 9647 7787
rect 9613 7653 9627 7667
rect 9553 7593 9567 7607
rect 9533 7513 9547 7527
rect 9573 7493 9587 7507
rect 9553 7453 9567 7467
rect 9513 7433 9527 7447
rect 9533 7433 9547 7447
rect 9533 7393 9547 7407
rect 9453 7373 9467 7387
rect 9533 7373 9547 7387
rect 9413 7053 9427 7067
rect 9513 7353 9527 7367
rect 9513 7053 9527 7067
rect 9493 7033 9507 7047
rect 9473 6953 9487 6967
rect 9453 6933 9467 6947
rect 9393 6893 9407 6907
rect 9533 6873 9547 6887
rect 9573 6873 9587 6887
rect 9613 6873 9627 6887
rect 9373 6853 9387 6867
rect 9473 6853 9487 6867
rect 9533 6613 9547 6627
rect 9573 6613 9587 6627
rect 9373 6573 9387 6587
rect 9393 6513 9407 6527
rect 9393 6453 9407 6467
rect 9373 6433 9387 6447
rect 9433 6293 9447 6307
rect 9593 6553 9607 6567
rect 9593 6433 9607 6447
rect 9553 6393 9567 6407
rect 9673 8033 9687 8047
rect 9713 7853 9727 7867
rect 9753 8233 9767 8247
rect 9753 8213 9767 8227
rect 9733 7773 9747 7787
rect 9793 8453 9807 8467
rect 9833 8573 9847 8587
rect 9873 8953 9887 8967
rect 9893 8933 9907 8947
rect 9893 8893 9907 8907
rect 9913 8793 9927 8807
rect 9873 8573 9887 8587
rect 9873 8553 9887 8567
rect 9993 9293 10007 9307
rect 9973 9233 9987 9247
rect 10033 9493 10047 9507
rect 10253 10913 10267 10927
rect 10293 10913 10307 10927
rect 10233 10733 10247 10747
rect 10193 10713 10207 10727
rect 10193 10453 10207 10467
rect 10173 9793 10187 9807
rect 10113 9433 10127 9447
rect 10113 9393 10127 9407
rect 10073 9353 10087 9367
rect 10033 9253 10047 9267
rect 9973 9213 9987 9227
rect 9953 8953 9967 8967
rect 10033 9133 10047 9147
rect 10033 9053 10047 9067
rect 9933 8553 9947 8567
rect 9833 8253 9847 8267
rect 9853 8253 9867 8267
rect 9813 8213 9827 8227
rect 9813 8133 9827 8147
rect 9793 8093 9807 8107
rect 9773 8073 9787 8087
rect 9773 8053 9787 8067
rect 9793 8053 9807 8067
rect 9853 8053 9867 8067
rect 9773 8033 9787 8047
rect 9833 8033 9847 8047
rect 9793 8013 9807 8027
rect 9853 7853 9867 7867
rect 9813 7833 9827 7847
rect 9873 7833 9887 7847
rect 9833 7813 9847 7827
rect 9873 7653 9887 7667
rect 9753 7573 9767 7587
rect 9933 8513 9947 8527
rect 9993 8813 10007 8827
rect 10013 8793 10027 8807
rect 10053 9013 10067 9027
rect 9973 8513 9987 8527
rect 10193 9353 10207 9367
rect 10133 9333 10147 9347
rect 10193 9313 10207 9327
rect 10513 11193 10527 11207
rect 10533 11193 10547 11207
rect 10473 11173 10487 11187
rect 10493 11153 10507 11167
rect 10513 11153 10527 11167
rect 10473 10893 10487 10907
rect 10493 10873 10507 10887
rect 10393 10613 10407 10627
rect 10293 10433 10307 10447
rect 10273 10333 10287 10347
rect 10313 10333 10327 10347
rect 10313 10313 10327 10327
rect 10333 10313 10347 10327
rect 10253 10253 10267 10267
rect 10313 10253 10327 10267
rect 10413 10513 10427 10527
rect 10393 10253 10407 10267
rect 10353 10213 10367 10227
rect 10393 10173 10407 10187
rect 10313 10093 10327 10107
rect 10293 9933 10307 9947
rect 10253 9913 10267 9927
rect 10273 9913 10287 9927
rect 10293 9893 10307 9907
rect 10233 9493 10247 9507
rect 10253 9433 10267 9447
rect 10653 11393 10667 11407
rect 10653 11273 10667 11287
rect 10573 11173 10587 11187
rect 10553 10593 10567 10607
rect 10433 10453 10447 10467
rect 10533 10453 10547 10467
rect 10433 10433 10447 10447
rect 10493 10433 10507 10447
rect 10533 10433 10547 10447
rect 10453 10413 10467 10427
rect 10433 10393 10447 10407
rect 10413 10033 10427 10047
rect 10393 9993 10407 10007
rect 10473 10373 10487 10387
rect 10493 10373 10507 10387
rect 10533 10353 10547 10367
rect 10513 10333 10527 10347
rect 10633 11193 10647 11207
rect 10653 10913 10667 10927
rect 10693 10873 10707 10887
rect 10613 10753 10627 10767
rect 10613 10693 10627 10707
rect 10673 10673 10687 10687
rect 10593 10653 10607 10667
rect 10633 10653 10647 10667
rect 10593 10633 10607 10647
rect 10593 10513 10607 10527
rect 10493 10313 10507 10327
rect 10573 10313 10587 10327
rect 10493 10233 10507 10247
rect 10433 9913 10447 9927
rect 10413 9893 10427 9907
rect 10413 9853 10427 9867
rect 10373 9773 10387 9787
rect 10333 9753 10347 9767
rect 10313 9493 10327 9507
rect 10273 9313 10287 9327
rect 10213 9273 10227 9287
rect 10193 9253 10207 9267
rect 10153 9213 10167 9227
rect 10133 9193 10147 9207
rect 10093 8993 10107 9007
rect 10133 8993 10147 9007
rect 10173 8993 10187 9007
rect 10093 8973 10107 8987
rect 10153 8973 10167 8987
rect 10153 8933 10167 8947
rect 10153 8873 10167 8887
rect 10233 9153 10247 9167
rect 10193 8953 10207 8967
rect 10213 8853 10227 8867
rect 10093 8753 10107 8767
rect 10073 8513 10087 8527
rect 10113 8513 10127 8527
rect 10033 8493 10047 8507
rect 10073 8473 10087 8487
rect 10113 8473 10127 8487
rect 10093 8453 10107 8467
rect 9953 8253 9967 8267
rect 10073 8373 10087 8387
rect 10073 8333 10087 8347
rect 9913 8133 9927 8147
rect 9913 8013 9927 8027
rect 9933 7973 9947 7987
rect 10053 8233 10067 8247
rect 9973 8093 9987 8107
rect 9953 7853 9967 7867
rect 9933 7813 9947 7827
rect 9733 7533 9747 7547
rect 9713 7513 9727 7527
rect 9653 7493 9667 7507
rect 9873 7533 9887 7547
rect 9893 7533 9907 7547
rect 9913 7533 9927 7547
rect 9953 7533 9967 7547
rect 9793 7513 9807 7527
rect 9793 7493 9807 7507
rect 9753 7473 9767 7487
rect 9833 7433 9847 7447
rect 9853 7373 9867 7387
rect 9933 7513 9947 7527
rect 9893 7373 9907 7387
rect 9893 7293 9907 7307
rect 9653 7073 9667 7087
rect 9693 7073 9707 7087
rect 9853 7073 9867 7087
rect 9713 7053 9727 7067
rect 9833 7053 9847 7067
rect 9713 6893 9727 6907
rect 9893 7013 9907 7027
rect 9693 6873 9707 6887
rect 9713 6853 9727 6867
rect 9673 6833 9687 6847
rect 9653 6613 9667 6627
rect 9873 6873 9887 6887
rect 9933 6853 9947 6867
rect 9773 6833 9787 6847
rect 9733 6793 9747 6807
rect 9753 6793 9767 6807
rect 9813 6713 9827 6727
rect 9673 6573 9687 6587
rect 9733 6573 9747 6587
rect 9653 6553 9667 6567
rect 9633 6413 9647 6427
rect 9613 6333 9627 6347
rect 9533 6273 9547 6287
rect 9433 6153 9447 6167
rect 9393 6113 9407 6127
rect 9753 6373 9767 6387
rect 9793 6553 9807 6567
rect 9793 6373 9807 6387
rect 9773 6353 9787 6367
rect 9713 6273 9727 6287
rect 9893 6633 9907 6647
rect 9953 6753 9967 6767
rect 9993 7913 10007 7927
rect 9993 7873 10007 7887
rect 10013 7873 10027 7887
rect 10053 7993 10067 8007
rect 10113 8273 10127 8287
rect 10093 7953 10107 7967
rect 10093 7813 10107 7827
rect 9993 7653 10007 7667
rect 10213 8793 10227 8807
rect 10173 8773 10187 8787
rect 10193 8753 10207 8767
rect 10533 10213 10547 10227
rect 10513 10193 10527 10207
rect 10553 10133 10567 10147
rect 10533 10113 10547 10127
rect 10493 9893 10507 9907
rect 10493 9813 10507 9827
rect 10453 9793 10467 9807
rect 10473 9713 10487 9727
rect 10433 9573 10447 9587
rect 10493 9693 10507 9707
rect 10413 9433 10427 9447
rect 10393 9413 10407 9427
rect 10353 9373 10367 9387
rect 10353 9293 10367 9307
rect 10293 9273 10307 9287
rect 10313 9273 10327 9287
rect 10433 9273 10447 9287
rect 10273 9253 10287 9267
rect 10373 9253 10387 9267
rect 10453 9233 10467 9247
rect 10353 9213 10367 9227
rect 10313 8973 10327 8987
rect 10333 8973 10347 8987
rect 10293 8913 10307 8927
rect 10273 8873 10287 8887
rect 10273 8833 10287 8847
rect 10233 8713 10247 8727
rect 10213 8593 10227 8607
rect 10213 8553 10227 8567
rect 10253 8493 10267 8507
rect 10153 8473 10167 8487
rect 10233 8433 10247 8447
rect 10193 8393 10207 8407
rect 10233 8353 10247 8367
rect 10253 8333 10267 8347
rect 10213 8313 10227 8327
rect 10553 9713 10567 9727
rect 10613 10453 10627 10467
rect 10733 11573 10747 11587
rect 10713 10573 10727 10587
rect 10673 10453 10687 10467
rect 10693 10433 10707 10447
rect 10673 10413 10687 10427
rect 10713 10413 10727 10427
rect 10893 11853 10907 11867
rect 10853 11833 10867 11847
rect 10833 11793 10847 11807
rect 10813 11413 10827 11427
rect 10793 11373 10807 11387
rect 10913 11833 10927 11847
rect 10933 11713 10947 11727
rect 10933 11673 10947 11687
rect 10873 11613 10887 11627
rect 10853 11273 10867 11287
rect 10833 11213 10847 11227
rect 10753 10993 10767 11007
rect 10753 10753 10767 10767
rect 10653 10373 10667 10387
rect 10693 10373 10707 10387
rect 10733 10373 10747 10387
rect 10633 10333 10647 10347
rect 10673 10333 10687 10347
rect 10613 10253 10627 10267
rect 10593 9973 10607 9987
rect 10613 9953 10627 9967
rect 10633 9933 10647 9947
rect 10653 9913 10667 9927
rect 10593 9733 10607 9747
rect 10573 9693 10587 9707
rect 10653 9553 10667 9567
rect 10573 9513 10587 9527
rect 10853 11193 10867 11207
rect 10853 10893 10867 10907
rect 10833 10873 10847 10887
rect 10813 10753 10827 10767
rect 10793 10733 10807 10747
rect 10793 10713 10807 10727
rect 10893 11413 10907 11427
rect 11153 11893 11167 11907
rect 11053 11873 11067 11887
rect 11093 11873 11107 11887
rect 11073 11833 11087 11847
rect 11053 11733 11067 11747
rect 11033 11693 11047 11707
rect 11013 11433 11027 11447
rect 10993 11413 11007 11427
rect 10913 11393 10927 11407
rect 10953 11393 10967 11407
rect 10893 11133 10907 11147
rect 10773 10693 10787 10707
rect 10773 10433 10787 10447
rect 10773 10353 10787 10367
rect 10873 10713 10887 10727
rect 10893 10713 10907 10727
rect 10853 10653 10867 10667
rect 10813 10573 10827 10587
rect 10793 10293 10807 10307
rect 10713 10253 10727 10267
rect 10753 10253 10767 10267
rect 10793 10253 10807 10267
rect 10693 10213 10707 10227
rect 10693 10173 10707 10187
rect 10753 10193 10767 10207
rect 10733 10113 10747 10127
rect 10693 10013 10707 10027
rect 10773 10133 10787 10147
rect 10773 9973 10787 9987
rect 10773 9953 10787 9967
rect 10753 9913 10767 9927
rect 10733 9893 10747 9907
rect 10713 9773 10727 9787
rect 10693 9713 10707 9727
rect 10713 9693 10727 9707
rect 10713 9513 10727 9527
rect 10673 9493 10687 9507
rect 10713 9493 10727 9507
rect 10633 9473 10647 9487
rect 10653 9453 10667 9467
rect 10613 9433 10627 9447
rect 10633 9433 10647 9447
rect 10593 9333 10607 9347
rect 10513 9253 10527 9267
rect 10573 9253 10587 9267
rect 10533 9233 10547 9247
rect 10433 9193 10447 9207
rect 10493 9193 10507 9207
rect 10373 9053 10387 9067
rect 10373 8973 10387 8987
rect 10393 8873 10407 8887
rect 10353 8773 10367 8787
rect 10413 8773 10427 8787
rect 10333 8733 10347 8747
rect 10473 8993 10487 9007
rect 10513 8993 10527 9007
rect 10453 8973 10467 8987
rect 10493 8973 10507 8987
rect 10453 8953 10467 8967
rect 10433 8713 10447 8727
rect 10433 8653 10447 8667
rect 10313 8453 10327 8467
rect 10333 8453 10347 8467
rect 10293 8353 10307 8367
rect 10313 8333 10327 8347
rect 10213 8273 10227 8287
rect 10233 8253 10247 8267
rect 10233 8093 10247 8107
rect 10153 8033 10167 8047
rect 10193 8033 10207 8047
rect 10213 8033 10227 8047
rect 10173 7993 10187 8007
rect 10213 7993 10227 8007
rect 10233 7993 10247 8007
rect 10213 7873 10227 7887
rect 10153 7853 10167 7867
rect 10013 7533 10027 7547
rect 10073 7513 10087 7527
rect 10113 7513 10127 7527
rect 10033 7473 10047 7487
rect 10013 7373 10027 7387
rect 9993 7353 10007 7367
rect 10053 7373 10067 7387
rect 10073 7373 10087 7387
rect 10013 7093 10027 7107
rect 10093 7093 10107 7107
rect 10113 7073 10127 7087
rect 10073 7053 10087 7067
rect 10313 7993 10327 8007
rect 10513 8773 10527 8787
rect 10413 8513 10427 8527
rect 10453 8513 10467 8527
rect 10473 8453 10487 8467
rect 10493 8293 10507 8307
rect 10433 8273 10447 8287
rect 10473 8273 10487 8287
rect 10513 8253 10527 8267
rect 10393 8173 10407 8187
rect 10373 8093 10387 8107
rect 10353 8053 10367 8067
rect 10613 9253 10627 9267
rect 10613 9193 10627 9207
rect 10553 9173 10567 9187
rect 10573 9093 10587 9107
rect 10593 9093 10607 9107
rect 10553 9073 10567 9087
rect 10553 9013 10567 9027
rect 10573 8993 10587 9007
rect 10553 8973 10567 8987
rect 10593 8973 10607 8987
rect 10593 8753 10607 8767
rect 10553 8733 10567 8747
rect 10593 8633 10607 8647
rect 10613 8633 10627 8647
rect 10653 9253 10667 9267
rect 10653 9173 10667 9187
rect 10713 9033 10727 9047
rect 10713 8993 10727 9007
rect 10653 8973 10667 8987
rect 10693 8973 10707 8987
rect 10673 8853 10687 8867
rect 10673 8813 10687 8827
rect 10633 8453 10647 8467
rect 10693 8673 10707 8687
rect 10693 8453 10707 8467
rect 10693 8433 10707 8447
rect 10713 8433 10727 8447
rect 10673 8413 10687 8427
rect 10673 8313 10687 8327
rect 10633 8293 10647 8307
rect 10613 8253 10627 8267
rect 10553 8193 10567 8207
rect 10533 8113 10547 8127
rect 10593 8113 10607 8127
rect 10413 8073 10427 8087
rect 10373 8033 10387 8047
rect 10333 7893 10347 7907
rect 10333 7853 10347 7867
rect 10553 8033 10567 8047
rect 10613 8053 10627 8067
rect 10633 8053 10647 8067
rect 10613 8013 10627 8027
rect 10633 7973 10647 7987
rect 10573 7953 10587 7967
rect 10633 7953 10647 7967
rect 10613 7893 10627 7907
rect 10413 7853 10427 7867
rect 10553 7853 10567 7867
rect 10593 7853 10607 7867
rect 10393 7833 10407 7847
rect 10373 7813 10387 7827
rect 10453 7813 10467 7827
rect 10333 7653 10347 7667
rect 10453 7613 10467 7627
rect 10253 7493 10267 7507
rect 10173 7413 10187 7427
rect 10433 7493 10447 7507
rect 10413 7413 10427 7427
rect 10233 7373 10247 7387
rect 10293 7373 10307 7387
rect 10193 7353 10207 7367
rect 10493 7553 10507 7567
rect 10573 7833 10587 7847
rect 10593 7793 10607 7807
rect 10593 7753 10607 7767
rect 10713 8013 10727 8027
rect 10753 9773 10767 9787
rect 10753 9613 10767 9627
rect 10773 9533 10787 9547
rect 10893 10473 10907 10487
rect 10853 10433 10867 10447
rect 10893 10433 10907 10447
rect 10833 10413 10847 10427
rect 10873 10373 10887 10387
rect 10893 10313 10907 10327
rect 10873 10273 10887 10287
rect 10933 11373 10947 11387
rect 10973 11373 10987 11387
rect 11013 11373 11027 11387
rect 11053 11673 11067 11687
rect 11113 11673 11127 11687
rect 11093 11613 11107 11627
rect 11073 11493 11087 11507
rect 11033 11293 11047 11307
rect 10993 11173 11007 11187
rect 11033 11073 11047 11087
rect 10993 10893 11007 10907
rect 11033 10893 11047 10907
rect 11013 10873 11027 10887
rect 10973 10773 10987 10787
rect 10953 10613 10967 10627
rect 10973 10493 10987 10507
rect 10953 10413 10967 10427
rect 10933 10333 10947 10347
rect 10913 10253 10927 10267
rect 10953 10253 10967 10267
rect 10893 10193 10907 10207
rect 10813 10153 10827 10167
rect 10913 10113 10927 10127
rect 10873 10053 10887 10067
rect 10813 9933 10827 9947
rect 10893 9993 10907 10007
rect 10833 9913 10847 9927
rect 10853 9873 10867 9887
rect 10933 10013 10947 10027
rect 10913 9873 10927 9887
rect 10893 9753 10907 9767
rect 10833 9593 10847 9607
rect 10853 9533 10867 9547
rect 10753 9513 10767 9527
rect 10793 9513 10807 9527
rect 10753 9473 10767 9487
rect 10833 9493 10847 9507
rect 10813 9473 10827 9487
rect 10773 9453 10787 9467
rect 10833 9453 10847 9467
rect 10773 9433 10787 9447
rect 10773 9333 10787 9347
rect 10813 9313 10827 9327
rect 10753 9193 10767 9207
rect 10773 9173 10787 9187
rect 10773 9013 10787 9027
rect 10753 8813 10767 8827
rect 10813 8973 10827 8987
rect 10873 9493 10887 9507
rect 10913 9733 10927 9747
rect 10893 9453 10907 9467
rect 10913 9433 10927 9447
rect 10873 9413 10887 9427
rect 10973 9993 10987 10007
rect 10953 9973 10967 9987
rect 11013 10713 11027 10727
rect 11033 10713 11047 10727
rect 11093 11433 11107 11447
rect 11133 11393 11147 11407
rect 11133 11273 11147 11287
rect 11133 11213 11147 11227
rect 11113 11153 11127 11167
rect 11133 11073 11147 11087
rect 11073 10953 11087 10967
rect 11193 11793 11207 11807
rect 11173 11593 11187 11607
rect 11693 11893 11707 11907
rect 11393 11873 11407 11887
rect 11373 11833 11387 11847
rect 11353 11773 11367 11787
rect 11273 11733 11287 11747
rect 11333 11713 11347 11727
rect 11293 11673 11307 11687
rect 11253 11653 11267 11667
rect 11273 11633 11287 11647
rect 11233 11513 11247 11527
rect 11333 11413 11347 11427
rect 11193 11333 11207 11347
rect 11293 11393 11307 11407
rect 11313 11393 11327 11407
rect 11313 11373 11327 11387
rect 11453 11853 11467 11867
rect 11433 11833 11447 11847
rect 11573 11833 11587 11847
rect 11473 11753 11487 11767
rect 11413 11613 11427 11627
rect 11393 11573 11407 11587
rect 11273 11293 11287 11307
rect 11333 11193 11347 11207
rect 11313 11173 11327 11187
rect 11333 11173 11347 11187
rect 11173 11153 11187 11167
rect 11153 11053 11167 11067
rect 11253 11053 11267 11067
rect 11153 10933 11167 10947
rect 11213 10933 11227 10947
rect 11173 10913 11187 10927
rect 11233 10833 11247 10847
rect 11193 10713 11207 10727
rect 11213 10693 11227 10707
rect 11133 10613 11147 10627
rect 11133 10573 11147 10587
rect 11113 10553 11127 10567
rect 11053 10493 11067 10507
rect 11053 10433 11067 10447
rect 11073 10413 11087 10427
rect 11193 10673 11207 10687
rect 11193 10613 11207 10627
rect 11153 10373 11167 10387
rect 11053 10293 11067 10307
rect 11133 10293 11147 10307
rect 11033 10273 11047 10287
rect 11093 10253 11107 10267
rect 11113 10253 11127 10267
rect 11053 10213 11067 10227
rect 11033 10113 11047 10127
rect 11013 10053 11027 10067
rect 11013 9973 11027 9987
rect 10973 9933 10987 9947
rect 11033 9873 11047 9887
rect 10953 9753 10967 9767
rect 11013 9753 11027 9767
rect 10933 9333 10947 9347
rect 11013 9733 11027 9747
rect 11093 10053 11107 10067
rect 11073 10013 11087 10027
rect 11073 9933 11087 9947
rect 11053 9833 11067 9847
rect 11053 9733 11067 9747
rect 11073 9713 11087 9727
rect 10993 9673 11007 9687
rect 10993 9633 11007 9647
rect 10993 9473 11007 9487
rect 11033 9473 11047 9487
rect 10973 9453 10987 9467
rect 11013 9433 11027 9447
rect 10993 9333 11007 9347
rect 10953 9313 10967 9327
rect 10853 9293 10867 9307
rect 10953 9293 10967 9307
rect 10913 9273 10927 9287
rect 10833 8953 10847 8967
rect 10893 8973 10907 8987
rect 10973 9253 10987 9267
rect 10953 9233 10967 9247
rect 10933 9213 10947 9227
rect 10873 8913 10887 8927
rect 10853 8873 10867 8887
rect 10913 8913 10927 8927
rect 10913 8873 10927 8887
rect 10893 8853 10907 8867
rect 10833 8773 10847 8787
rect 10773 8753 10787 8767
rect 10793 8753 10807 8767
rect 10793 8713 10807 8727
rect 10873 8633 10887 8647
rect 10833 8533 10847 8547
rect 10833 8493 10847 8507
rect 10813 8473 10827 8487
rect 10813 8413 10827 8427
rect 10813 8313 10827 8327
rect 10833 8313 10847 8327
rect 10853 8273 10867 8287
rect 10833 8213 10847 8227
rect 10833 8093 10847 8107
rect 10793 8053 10807 8067
rect 10773 8013 10787 8027
rect 10773 7893 10787 7907
rect 10753 7873 10767 7887
rect 10733 7853 10747 7867
rect 10793 7853 10807 7867
rect 10853 7853 10867 7867
rect 10753 7813 10767 7827
rect 10853 7833 10867 7847
rect 10933 8773 10947 8787
rect 10973 9113 10987 9127
rect 10933 8693 10947 8707
rect 10953 8693 10967 8707
rect 10913 8553 10927 8567
rect 10893 8313 10907 8327
rect 10913 8273 10927 8287
rect 10913 8173 10927 8187
rect 10973 8633 10987 8647
rect 11013 9253 11027 9267
rect 11153 10113 11167 10127
rect 11113 9973 11127 9987
rect 11293 10993 11307 11007
rect 11253 10533 11267 10547
rect 11353 11073 11367 11087
rect 11493 11673 11507 11687
rect 11533 11673 11547 11687
rect 11453 11573 11467 11587
rect 11433 11493 11447 11507
rect 11473 11253 11487 11267
rect 11453 11233 11467 11247
rect 11433 11173 11447 11187
rect 11453 11153 11467 11167
rect 11453 11093 11467 11107
rect 11413 11053 11427 11067
rect 11453 11053 11467 11067
rect 11433 10953 11447 10967
rect 11393 10933 11407 10947
rect 11373 10873 11387 10887
rect 11313 10833 11327 10847
rect 11333 10733 11347 10747
rect 11313 10673 11327 10687
rect 11353 10653 11367 10667
rect 11333 10613 11347 10627
rect 11313 10553 11327 10567
rect 11293 10493 11307 10507
rect 11253 10433 11267 10447
rect 11213 10413 11227 10427
rect 11213 10393 11227 10407
rect 11273 10413 11287 10427
rect 11293 10413 11307 10427
rect 11313 10413 11327 10427
rect 11273 10373 11287 10387
rect 11233 10253 11247 10267
rect 11213 10233 11227 10247
rect 11253 10193 11267 10207
rect 11213 10173 11227 10187
rect 11233 10173 11247 10187
rect 11193 9993 11207 10007
rect 11113 9953 11127 9967
rect 11153 9953 11167 9967
rect 11173 9933 11187 9947
rect 11133 9913 11147 9927
rect 11173 9873 11187 9887
rect 11153 9733 11167 9747
rect 11213 9953 11227 9967
rect 11193 9853 11207 9867
rect 11253 10033 11267 10047
rect 11273 10033 11287 10047
rect 11273 9993 11287 10007
rect 11253 9933 11267 9947
rect 11233 9893 11247 9907
rect 11233 9833 11247 9847
rect 11213 9793 11227 9807
rect 11193 9773 11207 9787
rect 11273 9773 11287 9787
rect 11253 9593 11267 9607
rect 11193 9533 11207 9547
rect 11233 9533 11247 9547
rect 11193 9513 11207 9527
rect 11193 9473 11207 9487
rect 11153 9433 11167 9447
rect 11193 9433 11207 9447
rect 11173 9393 11187 9407
rect 11133 9353 11147 9367
rect 11033 9093 11047 9107
rect 11013 9053 11027 9067
rect 11153 9293 11167 9307
rect 11093 9273 11107 9287
rect 11133 9273 11147 9287
rect 11113 9253 11127 9267
rect 11113 9233 11127 9247
rect 11173 9233 11187 9247
rect 11053 8973 11067 8987
rect 11013 8953 11027 8967
rect 11013 8793 11027 8807
rect 10993 8553 11007 8567
rect 10993 8493 11007 8507
rect 10973 8453 10987 8467
rect 10953 8433 10967 8447
rect 10973 8373 10987 8387
rect 11073 8953 11087 8967
rect 11033 8613 11047 8627
rect 11033 8493 11047 8507
rect 11133 9173 11147 9187
rect 11113 8933 11127 8947
rect 11093 8813 11107 8827
rect 11073 8793 11087 8807
rect 11073 8753 11087 8767
rect 11213 9413 11227 9427
rect 11213 9353 11227 9367
rect 11233 9313 11247 9327
rect 11213 9173 11227 9187
rect 11273 9513 11287 9527
rect 11153 9033 11167 9047
rect 11193 9033 11207 9047
rect 11233 9033 11247 9047
rect 11253 9033 11267 9047
rect 11173 9013 11187 9027
rect 11213 9013 11227 9027
rect 11193 8993 11207 9007
rect 11153 8873 11167 8887
rect 11013 8333 11027 8347
rect 11053 8333 11067 8347
rect 10973 8313 10987 8327
rect 11013 8313 11027 8327
rect 11053 8313 11067 8327
rect 10993 8293 11007 8307
rect 11033 8293 11047 8307
rect 11013 8253 11027 8267
rect 10993 8053 11007 8067
rect 11013 8033 11027 8047
rect 10953 8013 10967 8027
rect 10873 7813 10887 7827
rect 10893 7793 10907 7807
rect 10693 7733 10707 7747
rect 10733 7733 10747 7747
rect 10713 7713 10727 7727
rect 10633 7533 10647 7547
rect 10653 7533 10667 7547
rect 10633 7513 10647 7527
rect 10513 7493 10527 7507
rect 10553 7473 10567 7487
rect 10493 7373 10507 7387
rect 10173 7333 10187 7347
rect 10453 7353 10467 7367
rect 10273 7293 10287 7307
rect 10373 7293 10387 7307
rect 10333 7133 10347 7147
rect 10293 7093 10307 7107
rect 10253 7053 10267 7067
rect 10293 7033 10307 7047
rect 10313 7033 10327 7047
rect 10153 7013 10167 7027
rect 10033 6973 10047 6987
rect 10053 6893 10067 6907
rect 10033 6853 10047 6867
rect 10033 6813 10047 6827
rect 10193 6873 10207 6887
rect 10093 6853 10107 6867
rect 10113 6833 10127 6847
rect 10073 6813 10087 6827
rect 10053 6753 10067 6767
rect 9973 6673 9987 6687
rect 9913 6613 9927 6627
rect 10013 6613 10027 6627
rect 9973 6593 9987 6607
rect 9893 6573 9907 6587
rect 9953 6573 9967 6587
rect 10273 6853 10287 6867
rect 10313 6853 10327 6867
rect 10153 6593 10167 6607
rect 10193 6593 10207 6607
rect 10293 6833 10307 6847
rect 10253 6593 10267 6607
rect 10313 6593 10327 6607
rect 9573 6133 9587 6147
rect 9593 6113 9607 6127
rect 9373 6093 9387 6107
rect 9293 5733 9307 5747
rect 9353 5733 9367 5747
rect 9153 5673 9167 5687
rect 9153 5633 9167 5647
rect 9093 5613 9107 5627
rect 9173 5593 9187 5607
rect 9213 5593 9227 5607
rect 9253 5453 9267 5467
rect 9273 5453 9287 5467
rect 9253 5393 9267 5407
rect 9193 5313 9207 5327
rect 9133 5173 9147 5187
rect 9213 5173 9227 5187
rect 9173 5153 9187 5167
rect 9173 5133 9187 5147
rect 9193 5013 9207 5027
rect 9233 4953 9247 4967
rect 9153 4913 9167 4927
rect 9153 4873 9167 4887
rect 9093 4633 9107 4647
rect 9073 4613 9087 4627
rect 9053 4473 9067 4487
rect 9113 4513 9127 4527
rect 9033 4453 9047 4467
rect 9073 4453 9087 4467
rect 9113 4453 9127 4467
rect 9013 4273 9027 4287
rect 8973 4233 8987 4247
rect 8873 4213 8887 4227
rect 8913 4213 8927 4227
rect 8693 4033 8707 4047
rect 8813 4033 8827 4047
rect 8893 4053 8907 4067
rect 8853 3953 8867 3967
rect 8873 3793 8887 3807
rect 8553 3773 8567 3787
rect 8593 3713 8607 3727
rect 8653 3713 8667 3727
rect 8773 3713 8787 3727
rect 8533 3693 8547 3707
rect 8573 3693 8587 3707
rect 8613 3633 8627 3647
rect 8513 3513 8527 3527
rect 8613 3513 8627 3527
rect 8633 3493 8647 3507
rect 8613 3313 8627 3327
rect 8513 3293 8527 3307
rect 8533 3293 8547 3307
rect 8693 3273 8707 3287
rect 8673 3253 8687 3267
rect 8713 3253 8727 3267
rect 8533 3213 8547 3227
rect 8493 3193 8507 3207
rect 8453 3073 8467 3087
rect 8473 3053 8487 3067
rect 8413 3033 8427 3047
rect 8433 3033 8447 3047
rect 8573 2993 8587 3007
rect 8453 2973 8467 2987
rect 8393 2913 8407 2927
rect 8413 2873 8427 2887
rect 8453 2813 8467 2827
rect 8493 2753 8507 2767
rect 8533 2753 8547 2767
rect 8513 2733 8527 2747
rect 8453 2693 8467 2707
rect 8413 2593 8427 2607
rect 8433 2573 8447 2587
rect 8373 2513 8387 2527
rect 8353 2373 8367 2387
rect 8373 2313 8387 2327
rect 8313 2273 8327 2287
rect 8433 2273 8447 2287
rect 8293 2253 8307 2267
rect 8373 2253 8387 2267
rect 8293 2193 8307 2207
rect 8293 2133 8307 2147
rect 8253 2113 8267 2127
rect 8273 2113 8287 2127
rect 8273 2093 8287 2107
rect 8213 2073 8227 2087
rect 8233 2073 8247 2087
rect 8253 2033 8267 2047
rect 8213 2013 8227 2027
rect 8253 2013 8267 2027
rect 8353 2213 8367 2227
rect 8333 2193 8347 2207
rect 8233 1993 8247 2007
rect 8193 1833 8207 1847
rect 8173 1813 8187 1827
rect 8133 1573 8147 1587
rect 8133 1553 8147 1567
rect 8113 1333 8127 1347
rect 8173 1573 8187 1587
rect 8213 1533 8227 1547
rect 8193 1413 8207 1427
rect 8213 1413 8227 1427
rect 8193 1313 8207 1327
rect 8153 1293 8167 1307
rect 8093 1273 8107 1287
rect 8133 1273 8147 1287
rect 8173 1273 8187 1287
rect 8193 1273 8207 1287
rect 8053 1233 8067 1247
rect 7993 1113 8007 1127
rect 8093 1113 8107 1127
rect 8133 1113 8147 1127
rect 8033 1093 8047 1107
rect 8073 1093 8087 1107
rect 8073 1013 8087 1027
rect 8093 1013 8107 1027
rect 8013 953 8027 967
rect 8013 873 8027 887
rect 7973 853 7987 867
rect 7993 833 8007 847
rect 7953 613 7967 627
rect 7933 593 7947 607
rect 7973 553 7987 567
rect 7893 413 7907 427
rect 8093 853 8107 867
rect 8253 1933 8267 1947
rect 8273 1813 8287 1827
rect 8553 2553 8567 2567
rect 8653 3213 8667 3227
rect 8713 3153 8727 3167
rect 8613 3073 8627 3087
rect 8653 3053 8667 3067
rect 8693 3033 8707 3047
rect 8633 3013 8647 3027
rect 8673 3013 8687 3027
rect 8673 2833 8687 2847
rect 8653 2753 8667 2767
rect 8593 2733 8607 2747
rect 8833 3513 8847 3527
rect 8853 3433 8867 3447
rect 8833 3373 8847 3387
rect 8793 3253 8807 3267
rect 8873 3233 8887 3247
rect 8793 3213 8807 3227
rect 8813 3213 8827 3227
rect 8833 3193 8847 3207
rect 8793 3033 8807 3047
rect 8813 3033 8827 3047
rect 8873 3193 8887 3207
rect 8853 3073 8867 3087
rect 8773 2993 8787 3007
rect 8793 2993 8807 3007
rect 8853 2973 8867 2987
rect 8873 2973 8887 2987
rect 8853 2813 8867 2827
rect 8653 2633 8667 2647
rect 8673 2573 8687 2587
rect 8633 2553 8647 2567
rect 8533 2373 8547 2387
rect 8653 2433 8667 2447
rect 8593 2393 8607 2407
rect 8613 2393 8627 2407
rect 8573 2373 8587 2387
rect 8553 2353 8567 2367
rect 8593 2333 8607 2347
rect 8573 2313 8587 2327
rect 8513 2253 8527 2267
rect 8473 2213 8487 2227
rect 8553 2193 8567 2207
rect 8473 2153 8487 2167
rect 8413 2133 8427 2147
rect 8393 2093 8407 2107
rect 8373 1973 8387 1987
rect 8353 1933 8367 1947
rect 8273 1773 8287 1787
rect 8273 1653 8287 1667
rect 8333 1813 8347 1827
rect 8553 2093 8567 2107
rect 8513 2073 8527 2087
rect 8413 2053 8427 2067
rect 8493 2053 8507 2067
rect 8493 2033 8507 2047
rect 8553 2053 8567 2067
rect 8453 1973 8467 1987
rect 8433 1913 8447 1927
rect 8353 1773 8367 1787
rect 8313 1753 8327 1767
rect 8413 1733 8427 1747
rect 8433 1733 8447 1747
rect 8313 1713 8327 1727
rect 8333 1713 8347 1727
rect 8313 1653 8327 1667
rect 8373 1593 8387 1607
rect 8333 1573 8347 1587
rect 8393 1553 8407 1567
rect 8473 1813 8487 1827
rect 8473 1793 8487 1807
rect 8313 1513 8327 1527
rect 8333 1513 8347 1527
rect 8293 1433 8307 1447
rect 8233 1313 8247 1327
rect 8213 1073 8227 1087
rect 8193 1033 8207 1047
rect 8173 873 8187 887
rect 8273 1193 8287 1207
rect 8253 1113 8267 1127
rect 8353 1313 8367 1327
rect 8333 1293 8347 1307
rect 8373 1293 8387 1307
rect 8313 1133 8327 1147
rect 8473 1533 8487 1547
rect 8453 1333 8467 1347
rect 8453 1293 8467 1307
rect 8473 1173 8487 1187
rect 8393 1093 8407 1107
rect 8413 1093 8427 1107
rect 8453 1093 8467 1107
rect 8133 833 8147 847
rect 8153 833 8167 847
rect 8233 833 8247 847
rect 8173 813 8187 827
rect 8073 773 8087 787
rect 8193 673 8207 687
rect 8153 633 8167 647
rect 8213 633 8227 647
rect 8173 613 8187 627
rect 8113 573 8127 587
rect 8213 573 8227 587
rect 8233 573 8247 587
rect 8033 453 8047 467
rect 7993 373 8007 387
rect 7913 333 7927 347
rect 8113 393 8127 407
rect 8073 353 8087 367
rect 8093 333 8107 347
rect 8133 293 8147 307
rect 8113 253 8127 267
rect 7913 173 7927 187
rect 8073 173 8087 187
rect 7793 113 7807 127
rect 7913 133 7927 147
rect 7513 93 7527 107
rect 7853 113 7867 127
rect 7873 113 7887 127
rect 8293 1073 8307 1087
rect 8293 913 8307 927
rect 8313 893 8327 907
rect 8333 833 8347 847
rect 8373 833 8387 847
rect 8473 933 8487 947
rect 8293 653 8307 667
rect 8313 653 8327 667
rect 8393 793 8407 807
rect 8353 753 8367 767
rect 8393 753 8407 767
rect 8373 633 8387 647
rect 8273 613 8287 627
rect 8333 613 8347 627
rect 8273 533 8287 547
rect 8333 433 8347 447
rect 8293 373 8307 387
rect 8413 653 8427 667
rect 8393 413 8407 427
rect 8593 2213 8607 2227
rect 8573 1973 8587 1987
rect 8573 1873 8587 1887
rect 8593 1853 8607 1867
rect 8533 1773 8547 1787
rect 8553 1773 8567 1787
rect 8673 2353 8687 2367
rect 8633 2313 8647 2327
rect 8673 2253 8687 2267
rect 8753 2753 8767 2767
rect 8793 2753 8807 2767
rect 8773 2733 8787 2747
rect 8733 2713 8747 2727
rect 8713 2533 8727 2547
rect 8853 2713 8867 2727
rect 8793 2693 8807 2707
rect 8833 2653 8847 2667
rect 8813 2573 8827 2587
rect 8773 2533 8787 2547
rect 8773 2453 8787 2467
rect 8733 2333 8747 2347
rect 8753 2333 8767 2347
rect 8733 2293 8747 2307
rect 8753 2293 8767 2307
rect 8713 2273 8727 2287
rect 8733 2253 8747 2267
rect 8753 2173 8767 2187
rect 8733 2113 8747 2127
rect 8693 2093 8707 2107
rect 8653 2073 8667 2087
rect 8633 2053 8647 2067
rect 8673 2053 8687 2067
rect 8713 1953 8727 1967
rect 8733 1953 8747 1967
rect 8633 1873 8647 1887
rect 8513 1753 8527 1767
rect 8553 1753 8567 1767
rect 8533 1673 8547 1687
rect 8513 1153 8527 1167
rect 8693 1853 8707 1867
rect 8713 1853 8727 1867
rect 8713 1793 8727 1807
rect 8693 1753 8707 1767
rect 8733 1753 8747 1767
rect 8953 3973 8967 3987
rect 8913 3953 8927 3967
rect 8913 3713 8927 3727
rect 9053 4213 9067 4227
rect 9033 4193 9047 4207
rect 9053 4013 9067 4027
rect 9013 3973 9027 3987
rect 8993 3953 9007 3967
rect 9193 4713 9207 4727
rect 9453 6073 9467 6087
rect 9433 5933 9447 5947
rect 9353 5573 9367 5587
rect 9473 5913 9487 5927
rect 9533 5933 9547 5947
rect 9493 5893 9507 5907
rect 9493 5873 9507 5887
rect 9673 6133 9687 6147
rect 9813 6133 9827 6147
rect 10033 6553 10047 6567
rect 10173 6553 10187 6567
rect 9993 6413 10007 6427
rect 9973 6393 9987 6407
rect 9933 6373 9947 6387
rect 9913 6353 9927 6367
rect 9973 6333 9987 6347
rect 9953 6153 9967 6167
rect 9893 6113 9907 6127
rect 9773 6093 9787 6107
rect 9813 6093 9827 6107
rect 9633 6073 9647 6087
rect 9653 6073 9667 6087
rect 9673 6053 9687 6067
rect 9813 6033 9827 6047
rect 9713 5933 9727 5947
rect 9653 5873 9667 5887
rect 9693 5873 9707 5887
rect 9573 5853 9587 5867
rect 9593 5853 9607 5867
rect 9533 5713 9547 5727
rect 9573 5633 9587 5647
rect 9773 5893 9787 5907
rect 9733 5853 9747 5867
rect 9773 5713 9787 5727
rect 9933 5913 9947 5927
rect 9913 5893 9927 5907
rect 9933 5873 9947 5887
rect 9893 5693 9907 5707
rect 9933 5693 9947 5707
rect 9993 6093 10007 6107
rect 9513 5613 9527 5627
rect 9433 5473 9447 5487
rect 9413 5453 9427 5467
rect 9353 5433 9367 5447
rect 9373 5433 9387 5447
rect 9333 5413 9347 5427
rect 9553 5453 9567 5467
rect 9653 5613 9667 5627
rect 9733 5613 9747 5627
rect 9813 5613 9827 5627
rect 9713 5493 9727 5507
rect 9793 5493 9807 5507
rect 9813 5473 9827 5487
rect 9713 5413 9727 5427
rect 9393 5393 9407 5407
rect 9613 5393 9627 5407
rect 9713 5393 9727 5407
rect 9793 5433 9807 5447
rect 9773 5413 9787 5427
rect 10133 6433 10147 6447
rect 10073 6413 10087 6427
rect 10113 6413 10127 6427
rect 10093 6373 10107 6387
rect 10193 6393 10207 6407
rect 10113 6093 10127 6107
rect 10133 6053 10147 6067
rect 10113 5913 10127 5927
rect 10153 5913 10167 5927
rect 10093 5893 10107 5907
rect 10293 6393 10307 6407
rect 10253 6333 10267 6347
rect 10273 6333 10287 6347
rect 10493 7073 10507 7087
rect 10593 7373 10607 7387
rect 10573 7333 10587 7347
rect 10673 7473 10687 7487
rect 10633 7333 10647 7347
rect 10633 7293 10647 7307
rect 10613 7193 10627 7207
rect 10833 7533 10847 7547
rect 10853 7493 10867 7507
rect 10933 7933 10947 7947
rect 10933 7813 10947 7827
rect 10913 7453 10927 7467
rect 10913 7393 10927 7407
rect 10773 7373 10787 7387
rect 10753 7333 10767 7347
rect 10793 7333 10807 7347
rect 10733 7273 10747 7287
rect 10913 7313 10927 7327
rect 10953 7773 10967 7787
rect 10993 7973 11007 7987
rect 11053 7713 11067 7727
rect 11053 7573 11067 7587
rect 11293 9473 11307 9487
rect 11233 8853 11247 8867
rect 11253 8853 11267 8867
rect 11273 8833 11287 8847
rect 11273 8813 11287 8827
rect 11353 10453 11367 10467
rect 11333 10113 11347 10127
rect 11333 9933 11347 9947
rect 11333 9773 11347 9787
rect 11473 10973 11487 10987
rect 11453 10873 11467 10887
rect 11413 10813 11427 10827
rect 11473 10793 11487 10807
rect 11453 10773 11467 10787
rect 11513 11433 11527 11447
rect 11553 11593 11567 11607
rect 11553 11493 11567 11507
rect 11533 11413 11547 11427
rect 11533 11313 11547 11327
rect 11513 11233 11527 11247
rect 11533 11193 11547 11207
rect 11533 11113 11547 11127
rect 11533 11033 11547 11047
rect 11513 10973 11527 10987
rect 11513 10953 11527 10967
rect 11413 10753 11427 10767
rect 11393 10553 11407 10567
rect 11373 10413 11387 10427
rect 11393 10413 11407 10427
rect 11373 10393 11387 10407
rect 11393 10293 11407 10307
rect 11373 10213 11387 10227
rect 11433 10713 11447 10727
rect 11433 10653 11447 10667
rect 11633 11833 11647 11847
rect 11613 11773 11627 11787
rect 11593 11613 11607 11627
rect 11573 11433 11587 11447
rect 11573 11413 11587 11427
rect 11553 10953 11567 10967
rect 11533 10873 11547 10887
rect 11513 10753 11527 10767
rect 11493 10733 11507 10747
rect 11573 10893 11587 10907
rect 11573 10793 11587 10807
rect 11533 10713 11547 10727
rect 11553 10713 11567 10727
rect 11473 10613 11487 10627
rect 11553 10693 11567 10707
rect 11533 10533 11547 10547
rect 11513 10513 11527 10527
rect 11513 10493 11527 10507
rect 11453 10453 11467 10467
rect 11453 10433 11467 10447
rect 11433 10413 11447 10427
rect 11473 10413 11487 10427
rect 11493 10413 11507 10427
rect 11413 10253 11427 10267
rect 11473 10253 11487 10267
rect 11433 10233 11447 10247
rect 11433 10213 11447 10227
rect 11393 10193 11407 10207
rect 11453 10193 11467 10207
rect 11413 10173 11427 10187
rect 11373 10013 11387 10027
rect 11433 10113 11447 10127
rect 11413 9913 11427 9927
rect 11393 9893 11407 9907
rect 11413 9893 11427 9907
rect 11373 9853 11387 9867
rect 11453 9933 11467 9947
rect 11453 9913 11467 9927
rect 11433 9873 11447 9887
rect 11413 9813 11427 9827
rect 11393 9793 11407 9807
rect 11433 9753 11447 9767
rect 11373 9633 11387 9647
rect 11353 9533 11367 9547
rect 11433 9533 11447 9547
rect 11353 9513 11367 9527
rect 11413 9513 11427 9527
rect 11393 9453 11407 9467
rect 11373 9433 11387 9447
rect 11333 9393 11347 9407
rect 11333 9313 11347 9327
rect 11313 9273 11327 9287
rect 11373 9293 11387 9307
rect 11393 9293 11407 9307
rect 11393 9273 11407 9287
rect 11313 9253 11327 9267
rect 11313 9133 11327 9147
rect 11313 8993 11327 9007
rect 11393 9013 11407 9027
rect 11373 8993 11387 9007
rect 11333 8913 11347 8927
rect 11293 8793 11307 8807
rect 11213 8773 11227 8787
rect 11253 8773 11267 8787
rect 11133 8533 11147 8547
rect 11153 8513 11167 8527
rect 11113 8453 11127 8467
rect 11113 8433 11127 8447
rect 11093 8333 11107 8347
rect 11133 8393 11147 8407
rect 11113 8313 11127 8327
rect 11113 8293 11127 8307
rect 11113 8113 11127 8127
rect 11233 8533 11247 8547
rect 11213 8393 11227 8407
rect 11153 8333 11167 8347
rect 11153 8253 11167 8267
rect 11253 8473 11267 8487
rect 11313 8533 11327 8547
rect 11313 8493 11327 8507
rect 11213 8293 11227 8307
rect 11193 8273 11207 8287
rect 11193 8253 11207 8267
rect 11193 8233 11207 8247
rect 11133 8093 11147 8107
rect 11093 8073 11107 8087
rect 11093 8053 11107 8067
rect 11153 8053 11167 8067
rect 11113 8033 11127 8047
rect 11173 8013 11187 8027
rect 11233 8213 11247 8227
rect 11213 8113 11227 8127
rect 11133 7993 11147 8007
rect 11193 7993 11207 8007
rect 11233 8093 11247 8107
rect 11173 7953 11187 7967
rect 11213 7953 11227 7967
rect 11133 7853 11147 7867
rect 11113 7793 11127 7807
rect 11153 7793 11167 7807
rect 11093 7673 11107 7687
rect 11293 8453 11307 8467
rect 11273 8033 11287 8047
rect 11273 7973 11287 7987
rect 11373 8853 11387 8867
rect 11353 8493 11367 8507
rect 11353 8473 11367 8487
rect 11433 8933 11447 8947
rect 11433 8873 11447 8887
rect 11493 10213 11507 10227
rect 11493 9753 11507 9767
rect 11493 9733 11507 9747
rect 11493 9573 11507 9587
rect 11473 9513 11487 9527
rect 11473 9493 11487 9507
rect 11453 8813 11467 8827
rect 11753 11873 11767 11887
rect 11913 11853 11927 11867
rect 11813 11753 11827 11767
rect 11713 11713 11727 11727
rect 11893 11653 11907 11667
rect 11653 11553 11667 11567
rect 11693 11553 11707 11567
rect 11733 11553 11747 11567
rect 11633 11433 11647 11447
rect 11613 11293 11627 11307
rect 11673 11413 11687 11427
rect 11713 11413 11727 11427
rect 11693 11393 11707 11407
rect 11653 11333 11667 11347
rect 11633 11233 11647 11247
rect 11613 11193 11627 11207
rect 11693 11233 11707 11247
rect 11633 11133 11647 11147
rect 11613 10993 11627 11007
rect 11613 10933 11627 10947
rect 11633 10753 11647 10767
rect 11613 10733 11627 10747
rect 11633 10713 11647 10727
rect 11613 10673 11627 10687
rect 11613 10553 11627 10567
rect 11673 11093 11687 11107
rect 11713 11093 11727 11107
rect 11693 10773 11707 10787
rect 11653 10693 11667 10707
rect 11633 10513 11647 10527
rect 11613 10493 11627 10507
rect 11593 10393 11607 10407
rect 11813 11533 11827 11547
rect 11773 11453 11787 11467
rect 11793 11413 11807 11427
rect 11853 11473 11867 11487
rect 11833 11413 11847 11427
rect 11813 11393 11827 11407
rect 11793 11373 11807 11387
rect 11833 11333 11847 11347
rect 11773 11033 11787 11047
rect 11993 11893 12007 11907
rect 11973 11853 11987 11867
rect 11993 11753 12007 11767
rect 11933 11573 11947 11587
rect 11973 11553 11987 11567
rect 12013 11733 12027 11747
rect 11993 11473 12007 11487
rect 11913 11453 11927 11467
rect 11873 11413 11887 11427
rect 11893 11393 11907 11407
rect 11933 11373 11947 11387
rect 11873 11353 11887 11367
rect 11913 11353 11927 11367
rect 12033 11373 12047 11387
rect 12013 11133 12027 11147
rect 11993 11033 12007 11047
rect 11813 11013 11827 11027
rect 11853 11013 11867 11027
rect 11733 10733 11747 10747
rect 11773 10733 11787 10747
rect 11753 10713 11767 10727
rect 11753 10673 11767 10687
rect 11733 10653 11747 10667
rect 11733 10513 11747 10527
rect 11673 10473 11687 10487
rect 11653 10453 11667 10467
rect 11713 10453 11727 10467
rect 11693 10433 11707 10447
rect 11673 10413 11687 10427
rect 11673 10393 11687 10407
rect 11653 10353 11667 10367
rect 11633 10273 11647 10287
rect 11633 10253 11647 10267
rect 11553 10213 11567 10227
rect 11553 10193 11567 10207
rect 11633 10153 11647 10167
rect 11573 9993 11587 10007
rect 11573 9953 11587 9967
rect 11553 9933 11567 9947
rect 11533 9833 11547 9847
rect 11613 9913 11627 9927
rect 11613 9893 11627 9907
rect 11573 9853 11587 9867
rect 11573 9773 11587 9787
rect 11593 9733 11607 9747
rect 11593 9533 11607 9547
rect 11513 9493 11527 9507
rect 11553 9493 11567 9507
rect 11593 9493 11607 9507
rect 11533 9473 11547 9487
rect 11513 9453 11527 9467
rect 11553 9453 11567 9467
rect 11673 10153 11687 10167
rect 11713 10353 11727 10367
rect 11713 10293 11727 10307
rect 11713 10193 11727 10207
rect 11653 10073 11667 10087
rect 11633 9873 11647 9887
rect 11633 9833 11647 9847
rect 11613 9473 11627 9487
rect 11593 9453 11607 9467
rect 11573 9433 11587 9447
rect 11613 9373 11627 9387
rect 11493 9273 11507 9287
rect 11553 9253 11567 9267
rect 11513 9233 11527 9247
rect 11493 9153 11507 9167
rect 11493 8993 11507 9007
rect 11473 8793 11487 8807
rect 11413 8773 11427 8787
rect 11453 8733 11467 8747
rect 11393 8553 11407 8567
rect 11433 8553 11447 8567
rect 11413 8513 11427 8527
rect 11373 8353 11387 8367
rect 11393 8333 11407 8347
rect 11413 8333 11427 8347
rect 11413 8313 11427 8327
rect 11333 8213 11347 8227
rect 11313 8193 11327 8207
rect 11313 8153 11327 8167
rect 11293 7873 11307 7887
rect 11273 7853 11287 7867
rect 11253 7813 11267 7827
rect 11293 7813 11307 7827
rect 11333 8073 11347 8087
rect 11353 8013 11367 8027
rect 11373 7993 11387 8007
rect 11393 7853 11407 7867
rect 11333 7813 11347 7827
rect 11393 7813 11407 7827
rect 11313 7793 11327 7807
rect 11373 7793 11387 7807
rect 11313 7753 11327 7767
rect 11353 7753 11367 7767
rect 11233 7593 11247 7607
rect 11173 7573 11187 7587
rect 11073 7553 11087 7567
rect 11033 7533 11047 7547
rect 11253 7573 11267 7587
rect 11273 7553 11287 7567
rect 11293 7513 11307 7527
rect 11193 7473 11207 7487
rect 11173 7433 11187 7447
rect 10973 7373 10987 7387
rect 11353 7553 11367 7567
rect 11393 7773 11407 7787
rect 11533 9033 11547 9047
rect 11573 9013 11587 9027
rect 11553 8993 11567 9007
rect 11633 9233 11647 9247
rect 11613 8973 11627 8987
rect 11753 10433 11767 10447
rect 11793 10693 11807 10707
rect 11753 10413 11767 10427
rect 11773 10413 11787 10427
rect 11793 10353 11807 10367
rect 11773 10313 11787 10327
rect 11773 10233 11787 10247
rect 11973 10973 11987 10987
rect 11833 10873 11847 10887
rect 11833 10833 11847 10847
rect 11953 10813 11967 10827
rect 11913 10753 11927 10767
rect 11893 10673 11907 10687
rect 11933 10653 11947 10667
rect 11933 10493 11947 10507
rect 11933 10433 11947 10447
rect 11853 10413 11867 10427
rect 11893 10413 11907 10427
rect 11833 10353 11847 10367
rect 11853 10333 11867 10347
rect 11773 10193 11787 10207
rect 11813 10193 11827 10207
rect 11813 10173 11827 10187
rect 11753 10013 11767 10027
rect 11733 9973 11747 9987
rect 11733 9933 11747 9947
rect 11713 9913 11727 9927
rect 11673 9893 11687 9907
rect 11693 9893 11707 9907
rect 11673 9873 11687 9887
rect 11653 8953 11667 8967
rect 11593 8933 11607 8947
rect 11553 8913 11567 8927
rect 11533 8813 11547 8827
rect 11513 8593 11527 8607
rect 11573 8853 11587 8867
rect 11573 8793 11587 8807
rect 11553 8733 11567 8747
rect 11533 8573 11547 8587
rect 11453 8353 11467 8367
rect 11453 8013 11467 8027
rect 11453 7853 11467 7867
rect 11453 7773 11467 7787
rect 11373 7533 11387 7547
rect 10953 7353 10967 7367
rect 10953 7313 10967 7327
rect 10833 7153 10847 7167
rect 10813 7133 10827 7147
rect 10473 7053 10487 7067
rect 10653 7053 10667 7067
rect 10453 7033 10467 7047
rect 10873 7073 10887 7087
rect 10673 7013 10687 7027
rect 10433 6993 10447 7007
rect 10913 7053 10927 7067
rect 10633 6933 10647 6947
rect 10853 6933 10867 6947
rect 10893 6933 10907 6947
rect 10473 6893 10487 6907
rect 10573 6893 10587 6907
rect 10613 6893 10627 6907
rect 10593 6873 10607 6887
rect 10853 6913 10867 6927
rect 10673 6893 10687 6907
rect 10573 6813 10587 6827
rect 10453 6793 10467 6807
rect 10453 6753 10467 6767
rect 10373 6613 10387 6627
rect 10393 6593 10407 6607
rect 10433 6553 10447 6567
rect 10353 6433 10367 6447
rect 10813 6873 10827 6887
rect 10873 6873 10887 6887
rect 10833 6853 10847 6867
rect 10813 6833 10827 6847
rect 10773 6773 10787 6787
rect 10773 6613 10787 6627
rect 10573 6593 10587 6607
rect 10593 6553 10607 6567
rect 10553 6533 10567 6547
rect 10473 6473 10487 6487
rect 10673 6593 10687 6607
rect 10773 6593 10787 6607
rect 10913 6853 10927 6867
rect 10873 6773 10887 6787
rect 10633 6433 10647 6447
rect 10753 6553 10767 6567
rect 10793 6453 10807 6467
rect 10813 6433 10827 6447
rect 10353 6333 10367 6347
rect 10253 5933 10267 5947
rect 10233 5913 10247 5927
rect 10173 5893 10187 5907
rect 10093 5873 10107 5887
rect 10053 5693 10067 5707
rect 10033 5613 10047 5627
rect 10133 5613 10147 5627
rect 10313 5913 10327 5927
rect 10253 5893 10267 5907
rect 10293 5893 10307 5907
rect 10353 5913 10367 5927
rect 10233 5633 10247 5647
rect 10313 5633 10327 5647
rect 10353 5633 10367 5647
rect 10413 5633 10427 5647
rect 10153 5493 10167 5507
rect 10173 5473 10187 5487
rect 9933 5453 9947 5467
rect 9953 5453 9967 5467
rect 10013 5453 10027 5467
rect 10133 5453 10147 5467
rect 10193 5453 10207 5467
rect 9953 5433 9967 5447
rect 9993 5433 10007 5447
rect 9933 5413 9947 5427
rect 9973 5413 9987 5427
rect 10053 5433 10067 5447
rect 10073 5433 10087 5447
rect 10033 5413 10047 5427
rect 9573 5373 9587 5387
rect 9733 5373 9747 5387
rect 9353 5353 9367 5367
rect 9333 5313 9347 5327
rect 9393 5313 9407 5327
rect 9353 5193 9367 5207
rect 9573 5233 9587 5247
rect 9953 5193 9967 5207
rect 9313 5153 9327 5167
rect 9373 5153 9387 5167
rect 9593 5153 9607 5167
rect 9633 5153 9647 5167
rect 9753 5153 9767 5167
rect 9793 5153 9807 5167
rect 9553 5133 9567 5147
rect 9613 5133 9627 5147
rect 10053 5393 10067 5407
rect 10153 5433 10167 5447
rect 10313 5613 10327 5627
rect 10273 5493 10287 5507
rect 10233 5433 10247 5447
rect 10173 5413 10187 5427
rect 10133 5213 10147 5227
rect 10193 5213 10207 5227
rect 10153 5193 10167 5207
rect 10113 5173 10127 5187
rect 10073 5153 10087 5167
rect 9773 5113 9787 5127
rect 9813 5113 9827 5127
rect 9573 5093 9587 5107
rect 9633 5093 9647 5107
rect 10033 5113 10047 5127
rect 9313 4993 9327 5007
rect 9333 4993 9347 5007
rect 9973 4993 9987 5007
rect 9293 4873 9307 4887
rect 9253 4693 9267 4707
rect 9233 4653 9247 4667
rect 9193 4633 9207 4647
rect 9273 4633 9287 4647
rect 9513 4973 9527 4987
rect 9613 4973 9627 4987
rect 10053 4973 10067 4987
rect 9533 4933 9547 4947
rect 9813 4953 9827 4967
rect 9993 4953 10007 4967
rect 10033 4953 10047 4967
rect 9633 4933 9647 4947
rect 9653 4933 9667 4947
rect 9853 4933 9867 4947
rect 9893 4933 9907 4947
rect 9653 4893 9667 4907
rect 9453 4713 9467 4727
rect 9413 4693 9427 4707
rect 9433 4673 9447 4687
rect 9973 4913 9987 4927
rect 10053 4913 10067 4927
rect 9673 4853 9687 4867
rect 9913 4853 9927 4867
rect 9653 4753 9667 4767
rect 9793 4733 9807 4747
rect 9713 4713 9727 4727
rect 9613 4673 9627 4687
rect 9653 4673 9667 4687
rect 9693 4673 9707 4687
rect 9353 4653 9367 4667
rect 9593 4653 9607 4667
rect 9633 4653 9647 4667
rect 9673 4653 9687 4667
rect 9313 4473 9327 4487
rect 9253 4453 9267 4467
rect 9273 4433 9287 4447
rect 9253 4273 9267 4287
rect 9233 4213 9247 4227
rect 9213 4193 9227 4207
rect 9293 4213 9307 4227
rect 9293 4193 9307 4207
rect 9833 4713 9847 4727
rect 9813 4673 9827 4687
rect 9713 4653 9727 4667
rect 9693 4613 9707 4627
rect 9433 4493 9447 4507
rect 9773 4493 9787 4507
rect 9413 4453 9427 4467
rect 9453 4453 9467 4467
rect 9593 4473 9607 4487
rect 9513 4433 9527 4447
rect 9993 4713 10007 4727
rect 10173 5033 10187 5047
rect 10193 4973 10207 4987
rect 10213 4973 10227 4987
rect 10213 4933 10227 4947
rect 10173 4913 10187 4927
rect 10233 4893 10247 4907
rect 10033 4673 10047 4687
rect 10133 4673 10147 4687
rect 10193 4673 10207 4687
rect 10493 6373 10507 6387
rect 10533 6373 10547 6387
rect 10653 6373 10667 6387
rect 10833 6413 10847 6427
rect 10873 6413 10887 6427
rect 10933 6413 10947 6427
rect 10833 6393 10847 6407
rect 10873 6393 10887 6407
rect 10853 6373 10867 6387
rect 10933 6373 10947 6387
rect 11313 7333 11327 7347
rect 11153 7293 11167 7307
rect 10993 7273 11007 7287
rect 11153 7153 11167 7167
rect 11013 7093 11027 7107
rect 11033 7053 11047 7067
rect 11293 7093 11307 7107
rect 11353 7093 11367 7107
rect 11393 7093 11407 7107
rect 11213 7053 11227 7067
rect 10973 6933 10987 6947
rect 11093 7033 11107 7047
rect 11193 7033 11207 7047
rect 11013 6873 11027 6887
rect 11033 6873 11047 6887
rect 11033 6853 11047 6867
rect 10993 6793 11007 6807
rect 11013 6593 11027 6607
rect 11053 6593 11067 6607
rect 11033 6533 11047 6547
rect 10993 6433 11007 6447
rect 10973 6393 10987 6407
rect 11053 6413 11067 6427
rect 11013 6393 11027 6407
rect 10993 6373 11007 6387
rect 10953 6353 10967 6367
rect 11033 6353 11047 6367
rect 10653 6333 10667 6347
rect 10653 6313 10667 6327
rect 10513 6113 10527 6127
rect 10453 6053 10467 6067
rect 10493 6053 10507 6067
rect 10493 5993 10507 6007
rect 10573 6113 10587 6127
rect 10553 6073 10567 6087
rect 10573 5993 10587 6007
rect 10533 5933 10547 5947
rect 10573 5933 10587 5947
rect 10533 5913 10547 5927
rect 10553 5913 10567 5927
rect 10513 5893 10527 5907
rect 10473 5713 10487 5727
rect 10433 5613 10447 5627
rect 10493 5653 10507 5667
rect 10573 5893 10587 5907
rect 10473 5593 10487 5607
rect 10513 5593 10527 5607
rect 10373 5453 10387 5467
rect 10413 5453 10427 5467
rect 10513 5433 10527 5447
rect 10393 5413 10407 5427
rect 10373 5173 10387 5187
rect 10413 5173 10427 5187
rect 10373 5153 10387 5167
rect 10353 5133 10367 5147
rect 10433 5153 10447 5167
rect 10553 5453 10567 5467
rect 10593 5433 10607 5447
rect 10533 5413 10547 5427
rect 10573 5413 10587 5427
rect 10613 5413 10627 5427
rect 10633 5393 10647 5407
rect 10333 5053 10347 5067
rect 10333 5033 10347 5047
rect 10313 4993 10327 5007
rect 10393 4973 10407 4987
rect 10353 4933 10367 4947
rect 10293 4913 10307 4927
rect 10333 4913 10347 4927
rect 10273 4793 10287 4807
rect 10373 4733 10387 4747
rect 10293 4693 10307 4707
rect 9973 4653 9987 4667
rect 10253 4653 10267 4667
rect 10213 4553 10227 4567
rect 10013 4493 10027 4507
rect 10153 4493 10167 4507
rect 10333 4473 10347 4487
rect 10533 4993 10547 5007
rect 10493 4933 10507 4947
rect 10593 5133 10607 5147
rect 10633 5133 10647 5147
rect 10593 4993 10607 5007
rect 10553 4973 10567 4987
rect 10593 4973 10607 4987
rect 10553 4953 10567 4967
rect 10473 4733 10487 4747
rect 10433 4713 10447 4727
rect 10393 4693 10407 4707
rect 10453 4673 10467 4687
rect 10413 4653 10427 4667
rect 9933 4433 9947 4447
rect 9993 4433 10007 4447
rect 10373 4453 10387 4467
rect 10413 4453 10427 4467
rect 10573 4893 10587 4907
rect 10533 4793 10547 4807
rect 10613 4793 10627 4807
rect 10533 4633 10547 4647
rect 10493 4573 10507 4587
rect 10573 4633 10587 4647
rect 10553 4553 10567 4567
rect 10593 4473 10607 4487
rect 10613 4453 10627 4467
rect 10873 6153 10887 6167
rect 10773 6133 10787 6147
rect 10913 6113 10927 6127
rect 10733 6073 10747 6087
rect 10873 6073 10887 6087
rect 10713 5993 10727 6007
rect 10733 5993 10747 6007
rect 10673 5933 10687 5947
rect 10713 5933 10727 5947
rect 10713 5913 10727 5927
rect 10873 5933 10887 5947
rect 10753 5913 10767 5927
rect 10733 5893 10747 5907
rect 10693 5713 10707 5727
rect 10833 5813 10847 5827
rect 10753 5633 10767 5647
rect 10713 5573 10727 5587
rect 10693 5433 10707 5447
rect 10773 5613 10787 5627
rect 10933 6073 10947 6087
rect 10953 6073 10967 6087
rect 10973 6073 10987 6087
rect 10893 5913 10907 5927
rect 10913 5913 10927 5927
rect 10893 5893 10907 5907
rect 10913 5873 10927 5887
rect 10893 5653 10907 5667
rect 10853 5633 10867 5647
rect 10933 5813 10947 5827
rect 10833 5593 10847 5607
rect 10833 5573 10847 5587
rect 10773 5453 10787 5467
rect 10793 5453 10807 5467
rect 10793 5433 10807 5447
rect 10833 5433 10847 5447
rect 10913 5593 10927 5607
rect 10993 5613 11007 5627
rect 10953 5473 10967 5487
rect 10953 5453 10967 5467
rect 10733 5413 10747 5427
rect 10773 5413 10787 5427
rect 10813 5413 10827 5427
rect 10853 5413 10867 5427
rect 10973 5393 10987 5407
rect 10693 5173 10707 5187
rect 10733 5173 10747 5187
rect 10913 5173 10927 5187
rect 10733 5153 10747 5167
rect 10773 5153 10787 5167
rect 10973 5133 10987 5147
rect 11013 5393 11027 5407
rect 11013 5133 11027 5147
rect 10993 5113 11007 5127
rect 10953 5093 10967 5107
rect 10813 5013 10827 5027
rect 10733 4953 10747 4967
rect 10773 4953 10787 4967
rect 10973 4993 10987 5007
rect 10933 4973 10947 4987
rect 10753 4933 10767 4947
rect 10793 4933 10807 4947
rect 10753 4913 10767 4927
rect 10853 4753 10867 4767
rect 10793 4693 10807 4707
rect 10793 4613 10807 4627
rect 10773 4513 10787 4527
rect 10753 4473 10767 4487
rect 10833 4473 10847 4487
rect 10953 4933 10967 4947
rect 10933 4693 10947 4707
rect 10953 4613 10967 4627
rect 11013 4973 11027 4987
rect 10973 4533 10987 4547
rect 10773 4453 10787 4467
rect 10813 4453 10827 4467
rect 10853 4453 10867 4467
rect 10993 4453 11007 4467
rect 10653 4373 10667 4387
rect 10473 4273 10487 4287
rect 10493 4253 10507 4267
rect 9753 4233 9767 4247
rect 10493 4233 10507 4247
rect 10733 4233 10747 4247
rect 9493 4193 9507 4207
rect 9573 4193 9587 4207
rect 10193 4213 10207 4227
rect 9793 4193 9807 4207
rect 9993 4193 10007 4207
rect 10133 4193 10147 4207
rect 9353 4173 9367 4187
rect 9233 4153 9247 4167
rect 9193 4093 9207 4107
rect 9393 4053 9407 4067
rect 9373 4013 9387 4027
rect 8973 3933 8987 3947
rect 8933 3673 8947 3687
rect 8953 3513 8967 3527
rect 8913 3473 8927 3487
rect 8913 3193 8927 3207
rect 8933 3133 8947 3147
rect 8913 3113 8927 3127
rect 8913 3013 8927 3027
rect 8933 2973 8947 2987
rect 8893 2733 8907 2747
rect 8893 2673 8907 2687
rect 9053 3913 9067 3927
rect 9013 3713 9027 3727
rect 9133 3713 9147 3727
rect 9013 3673 9027 3687
rect 8993 3613 9007 3627
rect 9013 3533 9027 3547
rect 9053 3533 9067 3547
rect 9213 3993 9227 4007
rect 9313 3993 9327 4007
rect 9433 4153 9447 4167
rect 9413 4013 9427 4027
rect 9633 4173 9647 4187
rect 9933 4173 9947 4187
rect 9713 4153 9727 4167
rect 9953 4153 9967 4167
rect 9453 4133 9467 4147
rect 9653 4113 9667 4127
rect 9473 4053 9487 4067
rect 9373 3973 9387 3987
rect 9413 3973 9427 3987
rect 9313 3953 9327 3967
rect 9413 3953 9427 3967
rect 9313 3933 9327 3947
rect 9193 3873 9207 3887
rect 9253 3753 9267 3767
rect 9273 3713 9287 3727
rect 9353 3873 9367 3887
rect 9333 3693 9347 3707
rect 9253 3673 9267 3687
rect 9293 3673 9307 3687
rect 9273 3613 9287 3627
rect 9173 3533 9187 3547
rect 9113 3513 9127 3527
rect 8993 3493 9007 3507
rect 9033 3493 9047 3507
rect 9073 3473 9087 3487
rect 9093 3433 9107 3447
rect 8973 3393 8987 3407
rect 9013 3293 9027 3307
rect 8973 3253 8987 3267
rect 9053 3233 9067 3247
rect 8973 3213 8987 3227
rect 9033 3213 9047 3227
rect 9113 3353 9127 3367
rect 9233 3513 9247 3527
rect 9173 3293 9187 3307
rect 9173 3273 9187 3287
rect 9173 3253 9187 3267
rect 9113 3193 9127 3207
rect 9153 3193 9167 3207
rect 9113 3173 9127 3187
rect 8993 3133 9007 3147
rect 8993 3053 9007 3067
rect 9073 3053 9087 3067
rect 8973 3013 8987 3027
rect 8973 2853 8987 2867
rect 9033 3013 9047 3027
rect 9013 2993 9027 3007
rect 9093 2993 9107 3007
rect 9013 2893 9027 2907
rect 8993 2773 9007 2787
rect 8953 2713 8967 2727
rect 8973 2613 8987 2627
rect 9033 2873 9047 2887
rect 9073 2773 9087 2787
rect 9033 2713 9047 2727
rect 9033 2553 9047 2567
rect 8913 2313 8927 2327
rect 9013 2533 9027 2547
rect 9053 2533 9067 2547
rect 9033 2513 9047 2527
rect 9013 2473 9027 2487
rect 8953 2293 8967 2307
rect 8973 2293 8987 2307
rect 8893 2273 8907 2287
rect 8933 2273 8947 2287
rect 8873 2113 8887 2127
rect 8873 2073 8887 2087
rect 8813 2053 8827 2067
rect 8793 1753 8807 1767
rect 8773 1693 8787 1707
rect 8633 1573 8647 1587
rect 8693 1573 8707 1587
rect 8593 1533 8607 1547
rect 8553 1513 8567 1527
rect 8813 1733 8827 1747
rect 8913 2193 8927 2207
rect 8913 2093 8927 2107
rect 8873 1953 8887 1967
rect 8853 1713 8867 1727
rect 8793 1533 8807 1547
rect 8693 1453 8707 1467
rect 8593 1433 8607 1447
rect 8553 1393 8567 1407
rect 8553 1313 8567 1327
rect 8593 1313 8607 1327
rect 8673 1313 8687 1327
rect 8533 1073 8547 1087
rect 8613 1293 8627 1307
rect 8593 1193 8607 1207
rect 8633 1093 8647 1107
rect 8793 1393 8807 1407
rect 8713 1313 8727 1327
rect 8713 1293 8727 1307
rect 8733 1253 8747 1267
rect 8693 1093 8707 1107
rect 8573 1053 8587 1067
rect 8673 1013 8687 1027
rect 8533 973 8547 987
rect 8633 973 8647 987
rect 8533 933 8547 947
rect 8593 873 8607 887
rect 8513 833 8527 847
rect 8553 833 8567 847
rect 8593 833 8607 847
rect 8573 813 8587 827
rect 8493 793 8507 807
rect 8573 793 8587 807
rect 8553 693 8567 707
rect 8473 593 8487 607
rect 8413 373 8427 387
rect 8313 353 8327 367
rect 8493 533 8507 547
rect 8593 773 8607 787
rect 8533 513 8547 527
rect 8493 393 8507 407
rect 8533 393 8547 407
rect 8493 353 8507 367
rect 8473 333 8487 347
rect 8413 273 8427 287
rect 8253 213 8267 227
rect 8233 173 8247 187
rect 8393 173 8407 187
rect 8293 153 8307 167
rect 8433 173 8447 187
rect 8693 893 8707 907
rect 8653 833 8667 847
rect 8633 733 8647 747
rect 8613 693 8627 707
rect 8613 673 8627 687
rect 8613 653 8627 667
rect 8653 633 8667 647
rect 8713 733 8727 747
rect 8713 673 8727 687
rect 8693 613 8707 627
rect 8753 1193 8767 1207
rect 8893 1733 8907 1747
rect 8933 2073 8947 2087
rect 8933 1893 8947 1907
rect 8993 2253 9007 2267
rect 8993 2153 9007 2167
rect 8973 2113 8987 2127
rect 8993 2033 9007 2047
rect 8973 1973 8987 1987
rect 8953 1793 8967 1807
rect 8993 1793 9007 1807
rect 8933 1773 8947 1787
rect 8933 1733 8947 1747
rect 8913 1693 8927 1707
rect 9053 2413 9067 2427
rect 9073 2313 9087 2327
rect 9073 2253 9087 2267
rect 9133 3033 9147 3047
rect 9133 2993 9147 3007
rect 9133 2913 9147 2927
rect 9113 2813 9127 2827
rect 9173 3053 9187 3067
rect 9173 3033 9187 3047
rect 9233 3413 9247 3427
rect 9233 3273 9247 3287
rect 9293 3453 9307 3467
rect 9313 3293 9327 3307
rect 9253 3253 9267 3267
rect 9213 3213 9227 3227
rect 9253 3173 9267 3187
rect 9273 3173 9287 3187
rect 9213 3153 9227 3167
rect 9253 3133 9267 3147
rect 9193 2893 9207 2907
rect 9233 2893 9247 2907
rect 9173 2813 9187 2827
rect 9153 2773 9167 2787
rect 9153 2713 9167 2727
rect 9153 2653 9167 2667
rect 9113 2633 9127 2647
rect 9133 2533 9147 2547
rect 9133 2493 9147 2507
rect 9233 2573 9247 2587
rect 9213 2533 9227 2547
rect 9173 2353 9187 2367
rect 9153 2293 9167 2307
rect 9113 2273 9127 2287
rect 9153 2273 9167 2287
rect 9133 2233 9147 2247
rect 9133 2113 9147 2127
rect 9093 2093 9107 2107
rect 9093 2073 9107 2087
rect 9173 2233 9187 2247
rect 9173 2073 9187 2087
rect 9113 2053 9127 2067
rect 9153 2053 9167 2067
rect 9073 1993 9087 2007
rect 9033 1853 9047 1867
rect 9033 1753 9047 1767
rect 9013 1673 9027 1687
rect 8993 1653 9007 1667
rect 8953 1613 8967 1627
rect 8973 1613 8987 1627
rect 9053 1553 9067 1567
rect 8973 1533 8987 1547
rect 9013 1533 9027 1547
rect 8953 1393 8967 1407
rect 8933 1373 8947 1387
rect 8933 1333 8947 1347
rect 8993 1513 9007 1527
rect 8993 1473 9007 1487
rect 9033 1473 9047 1487
rect 9013 1333 9027 1347
rect 8893 1233 8907 1247
rect 8813 1113 8827 1127
rect 8833 1073 8847 1087
rect 8853 1073 8867 1087
rect 8773 993 8787 1007
rect 8793 773 8807 787
rect 8813 733 8827 747
rect 8753 673 8767 687
rect 8733 653 8747 667
rect 8793 633 8807 647
rect 8733 613 8747 627
rect 8773 613 8787 627
rect 8813 613 8827 627
rect 8713 553 8727 567
rect 8673 513 8687 527
rect 8613 433 8627 447
rect 8593 353 8607 367
rect 8653 373 8667 387
rect 8813 493 8827 507
rect 8733 373 8747 387
rect 8633 333 8647 347
rect 8693 333 8707 347
rect 8733 333 8747 347
rect 8673 253 8687 267
rect 8773 173 8787 187
rect 8873 1053 8887 1067
rect 8973 1153 8987 1167
rect 9013 1113 9027 1127
rect 8993 1093 9007 1107
rect 9053 1353 9067 1367
rect 9053 1313 9067 1327
rect 9113 1933 9127 1947
rect 9093 1853 9107 1867
rect 9113 1853 9127 1867
rect 9133 1793 9147 1807
rect 9113 1753 9127 1767
rect 9113 1713 9127 1727
rect 9093 1673 9107 1687
rect 9093 1653 9107 1667
rect 9073 1253 9087 1267
rect 9073 1233 9087 1247
rect 8953 1073 8967 1087
rect 8913 873 8927 887
rect 8933 833 8947 847
rect 8973 833 8987 847
rect 9013 833 9027 847
rect 8873 633 8887 647
rect 8933 793 8947 807
rect 8953 793 8967 807
rect 8913 733 8927 747
rect 9213 2093 9227 2107
rect 9213 1993 9227 2007
rect 9293 3133 9307 3147
rect 9293 3033 9307 3047
rect 9333 3073 9347 3087
rect 9333 3013 9347 3027
rect 9313 2893 9327 2907
rect 9293 2873 9307 2887
rect 9313 2873 9327 2887
rect 9293 2853 9307 2867
rect 9413 3853 9427 3867
rect 9373 3613 9387 3627
rect 9393 3533 9407 3547
rect 9373 3393 9387 3407
rect 9433 3533 9447 3547
rect 9493 4013 9507 4027
rect 9593 4013 9607 4027
rect 9473 3973 9487 3987
rect 9453 3513 9467 3527
rect 9393 3333 9407 3347
rect 9393 3253 9407 3267
rect 9373 3193 9387 3207
rect 9413 3193 9427 3207
rect 9413 3093 9427 3107
rect 9433 3093 9447 3107
rect 9373 3053 9387 3067
rect 9393 2853 9407 2867
rect 9353 2833 9367 2847
rect 9393 2793 9407 2807
rect 9353 2753 9367 2767
rect 9393 2753 9407 2767
rect 9333 2713 9347 2727
rect 9333 2633 9347 2647
rect 9353 2633 9367 2647
rect 9313 2553 9327 2567
rect 9273 2473 9287 2487
rect 9333 2533 9347 2547
rect 9333 2453 9347 2467
rect 9253 2293 9267 2307
rect 9273 2273 9287 2287
rect 9253 2253 9267 2267
rect 9233 1873 9247 1887
rect 9213 1793 9227 1807
rect 9193 1753 9207 1767
rect 9213 1753 9227 1767
rect 9173 1713 9187 1727
rect 9193 1593 9207 1607
rect 9273 2133 9287 2147
rect 9373 2573 9387 2587
rect 9373 2553 9387 2567
rect 9373 2413 9387 2427
rect 9353 2153 9367 2167
rect 9293 2113 9307 2127
rect 9353 2113 9367 2127
rect 9313 2093 9327 2107
rect 9293 2053 9307 2067
rect 9333 2033 9347 2047
rect 9293 1973 9307 1987
rect 9253 1813 9267 1827
rect 9293 1653 9307 1667
rect 9213 1573 9227 1587
rect 9273 1573 9287 1587
rect 9253 1553 9267 1567
rect 9153 1533 9167 1547
rect 9233 1533 9247 1547
rect 9133 1473 9147 1487
rect 9153 1333 9167 1347
rect 9173 1313 9187 1327
rect 9113 1293 9127 1307
rect 9193 1293 9207 1307
rect 9253 1433 9267 1447
rect 9253 1333 9267 1347
rect 9213 1233 9227 1247
rect 9233 1233 9247 1247
rect 9273 1273 9287 1287
rect 9273 1253 9287 1267
rect 9113 1153 9127 1167
rect 9213 1153 9227 1167
rect 9253 1153 9267 1167
rect 9093 1113 9107 1127
rect 9073 813 9087 827
rect 9013 793 9027 807
rect 8993 753 9007 767
rect 9033 693 9047 707
rect 8993 673 9007 687
rect 8893 613 8907 627
rect 8893 573 8907 587
rect 8973 613 8987 627
rect 8873 553 8887 567
rect 8933 553 8947 567
rect 8853 473 8867 487
rect 8893 413 8907 427
rect 8913 333 8927 347
rect 8873 293 8887 307
rect 8853 273 8867 287
rect 8973 233 8987 247
rect 8933 173 8947 187
rect 8633 133 8647 147
rect 8833 133 8847 147
rect 8953 133 8967 147
rect 9213 1093 9227 1107
rect 9233 1073 9247 1087
rect 9153 833 9167 847
rect 9253 853 9267 867
rect 9133 813 9147 827
rect 9113 673 9127 687
rect 9173 673 9187 687
rect 9133 633 9147 647
rect 9153 593 9167 607
rect 9073 533 9087 547
rect 9213 653 9227 667
rect 9093 513 9107 527
rect 9193 513 9207 527
rect 9033 373 9047 387
rect 9053 353 9067 367
rect 9153 353 9167 367
rect 9073 333 9087 347
rect 9113 333 9127 347
rect 9013 253 9027 267
rect 9233 573 9247 587
rect 9273 653 9287 667
rect 9273 633 9287 647
rect 9253 493 9267 507
rect 9253 353 9267 367
rect 9213 313 9227 327
rect 9213 173 9227 187
rect 9013 133 9027 147
rect 9313 1593 9327 1607
rect 9313 1393 9327 1407
rect 9353 1813 9367 1827
rect 9453 3053 9467 3067
rect 9453 2753 9467 2767
rect 9433 2473 9447 2487
rect 9573 3973 9587 3987
rect 9533 3933 9547 3947
rect 9533 3733 9547 3747
rect 9633 3733 9647 3747
rect 9693 4033 9707 4047
rect 9993 4153 10007 4167
rect 9973 4113 9987 4127
rect 9813 4073 9827 4087
rect 9753 4053 9767 4067
rect 9733 3993 9747 4007
rect 9793 3993 9807 4007
rect 9693 3973 9707 3987
rect 9713 3973 9727 3987
rect 9693 3733 9707 3747
rect 9673 3633 9687 3647
rect 9653 3613 9667 3627
rect 9573 3513 9587 3527
rect 9613 3513 9627 3527
rect 9493 3373 9507 3387
rect 9573 3373 9587 3387
rect 9553 3233 9567 3247
rect 9553 3153 9567 3167
rect 9553 3073 9567 3087
rect 9633 3353 9647 3367
rect 9653 3293 9667 3307
rect 9693 3293 9707 3307
rect 9593 3033 9607 3047
rect 9513 2993 9527 3007
rect 9573 2793 9587 2807
rect 9493 2753 9507 2767
rect 9533 2753 9547 2767
rect 9593 2753 9607 2767
rect 9513 2673 9527 2687
rect 9513 2613 9527 2627
rect 9473 2593 9487 2607
rect 9453 2453 9467 2467
rect 9433 2433 9447 2447
rect 9453 2433 9467 2447
rect 9393 2393 9407 2407
rect 9493 2573 9507 2587
rect 9493 2533 9507 2547
rect 9413 2333 9427 2347
rect 9433 2333 9447 2347
rect 9473 2333 9487 2347
rect 9413 2233 9427 2247
rect 9413 2133 9427 2147
rect 9413 2053 9427 2067
rect 9613 2733 9627 2747
rect 9653 3153 9667 3167
rect 9653 2913 9667 2927
rect 9633 2713 9647 2727
rect 9613 2693 9627 2707
rect 9553 2573 9567 2587
rect 9593 2573 9607 2587
rect 9593 2553 9607 2567
rect 9533 2533 9547 2547
rect 9573 2513 9587 2527
rect 9453 2253 9467 2267
rect 9513 2293 9527 2307
rect 9493 2113 9507 2127
rect 9453 2073 9467 2087
rect 9553 2273 9567 2287
rect 9533 2073 9547 2087
rect 9513 2053 9527 2067
rect 9433 2033 9447 2047
rect 9473 2033 9487 2047
rect 9393 1933 9407 1947
rect 9373 1733 9387 1747
rect 9373 1653 9387 1667
rect 9353 1613 9367 1627
rect 9393 1593 9407 1607
rect 9493 1993 9507 2007
rect 9433 1853 9447 1867
rect 9473 1853 9487 1867
rect 9413 1573 9427 1587
rect 9413 1533 9427 1547
rect 9333 1333 9347 1347
rect 9353 1333 9367 1347
rect 9313 1313 9327 1327
rect 9393 1313 9407 1327
rect 9313 1213 9327 1227
rect 9393 1253 9407 1267
rect 9453 1813 9467 1827
rect 9633 2553 9647 2567
rect 9613 2273 9627 2287
rect 9573 2253 9587 2267
rect 9593 2253 9607 2267
rect 9573 2053 9587 2067
rect 9553 1973 9567 1987
rect 9533 1873 9547 1887
rect 9513 1853 9527 1867
rect 9473 1793 9487 1807
rect 9453 1733 9467 1747
rect 9413 1173 9427 1187
rect 9433 1173 9447 1187
rect 9553 1853 9567 1867
rect 9693 3193 9707 3207
rect 9773 3973 9787 3987
rect 10113 4073 10127 4087
rect 10173 4173 10187 4187
rect 10153 4033 10167 4047
rect 9853 3993 9867 4007
rect 9993 3993 10007 4007
rect 10033 3993 10047 4007
rect 9773 3933 9787 3947
rect 9733 3913 9747 3927
rect 9753 3493 9767 3507
rect 9813 3493 9827 3507
rect 9833 3473 9847 3487
rect 9753 3433 9767 3447
rect 9833 3433 9847 3447
rect 9833 3273 9847 3287
rect 9953 3973 9967 3987
rect 9973 3953 9987 3967
rect 10313 4093 10327 4107
rect 10453 4173 10467 4187
rect 10513 4173 10527 4187
rect 10393 4013 10407 4027
rect 10233 3993 10247 4007
rect 10353 3993 10367 4007
rect 10213 3973 10227 3987
rect 10153 3953 10167 3967
rect 9953 3933 9967 3947
rect 10033 3933 10047 3947
rect 9913 3713 9927 3727
rect 9873 3693 9887 3707
rect 9893 3693 9907 3707
rect 10033 3733 10047 3747
rect 9973 3713 9987 3727
rect 9893 3653 9907 3667
rect 10013 3553 10027 3567
rect 9913 3533 9927 3547
rect 9973 3533 9987 3547
rect 9893 3473 9907 3487
rect 9893 3273 9907 3287
rect 9713 3173 9727 3187
rect 9733 3173 9747 3187
rect 9693 3073 9707 3087
rect 9733 3053 9747 3067
rect 9853 3213 9867 3227
rect 9853 3173 9867 3187
rect 9813 3153 9827 3167
rect 9833 3153 9847 3167
rect 9693 3013 9707 3027
rect 9753 3013 9767 3027
rect 9793 2973 9807 2987
rect 9713 2913 9727 2927
rect 9773 2773 9787 2787
rect 9713 2753 9727 2767
rect 9753 2753 9767 2767
rect 9733 2733 9747 2747
rect 9693 2713 9707 2727
rect 9673 2653 9687 2667
rect 9673 2593 9687 2607
rect 9653 2413 9667 2427
rect 9713 2693 9727 2707
rect 9753 2693 9767 2707
rect 9733 2613 9747 2627
rect 9713 2573 9727 2587
rect 9693 2513 9707 2527
rect 9673 2393 9687 2407
rect 9833 2793 9847 2807
rect 9793 2693 9807 2707
rect 9753 2513 9767 2527
rect 9733 2393 9747 2407
rect 9713 2333 9727 2347
rect 9713 2273 9727 2287
rect 9653 2253 9667 2267
rect 9613 2113 9627 2127
rect 9633 2073 9647 2087
rect 9693 2153 9707 2167
rect 9693 2113 9707 2127
rect 9673 2053 9687 2067
rect 9653 1993 9667 2007
rect 9733 1993 9747 2007
rect 9713 1973 9727 1987
rect 9633 1953 9647 1967
rect 9693 1953 9707 1967
rect 9613 1853 9627 1867
rect 9673 1813 9687 1827
rect 9593 1773 9607 1787
rect 9633 1793 9647 1807
rect 9653 1793 9667 1807
rect 9653 1773 9667 1787
rect 9613 1733 9627 1747
rect 9573 1673 9587 1687
rect 9593 1653 9607 1667
rect 9553 1613 9567 1627
rect 9553 1593 9567 1607
rect 9633 1593 9647 1607
rect 9573 1573 9587 1587
rect 9613 1553 9627 1567
rect 9673 1753 9687 1767
rect 9653 1433 9667 1447
rect 9533 1353 9547 1367
rect 9593 1353 9607 1367
rect 9513 1333 9527 1347
rect 9513 1313 9527 1327
rect 9513 1253 9527 1267
rect 9613 1293 9627 1307
rect 9553 1233 9567 1247
rect 9453 1153 9467 1167
rect 9693 1713 9707 1727
rect 9693 1613 9707 1627
rect 9833 2533 9847 2547
rect 9813 2473 9827 2487
rect 9773 2333 9787 2347
rect 9813 2313 9827 2327
rect 9813 2253 9827 2267
rect 9793 2153 9807 2167
rect 9773 2073 9787 2087
rect 9793 2073 9807 2087
rect 9793 2053 9807 2067
rect 9773 1993 9787 2007
rect 9753 1953 9767 1967
rect 9753 1893 9767 1907
rect 9753 1793 9767 1807
rect 9753 1773 9767 1787
rect 9893 3213 9907 3227
rect 9893 3013 9907 3027
rect 9893 2793 9907 2807
rect 9993 3493 10007 3507
rect 10073 3713 10087 3727
rect 10093 3653 10107 3667
rect 10133 3673 10147 3687
rect 10113 3533 10127 3547
rect 10113 3513 10127 3527
rect 10033 3413 10047 3427
rect 9993 3333 10007 3347
rect 9993 3233 10007 3247
rect 10073 3233 10087 3247
rect 9953 3153 9967 3167
rect 10053 3193 10067 3207
rect 10013 3133 10027 3147
rect 10093 3133 10107 3147
rect 9993 3033 10007 3047
rect 9953 3013 9967 3027
rect 9973 3013 9987 3027
rect 9933 2973 9947 2987
rect 9973 2793 9987 2807
rect 9913 2773 9927 2787
rect 9973 2753 9987 2767
rect 9913 2733 9927 2747
rect 9953 2733 9967 2747
rect 9993 2733 10007 2747
rect 9933 2713 9947 2727
rect 9893 2693 9907 2707
rect 9913 2693 9927 2707
rect 9873 2533 9887 2547
rect 9913 2673 9927 2687
rect 9953 2693 9967 2707
rect 10053 2993 10067 3007
rect 10033 2973 10047 2987
rect 10013 2633 10027 2647
rect 9933 2533 9947 2547
rect 9973 2533 9987 2547
rect 9913 2433 9927 2447
rect 9973 2333 9987 2347
rect 9893 2293 9907 2307
rect 9853 2273 9867 2287
rect 9933 2273 9947 2287
rect 9873 2253 9887 2267
rect 9973 2233 9987 2247
rect 9993 2233 10007 2247
rect 9973 2213 9987 2227
rect 9913 2153 9927 2167
rect 9873 2113 9887 2127
rect 9933 2113 9947 2127
rect 9913 2073 9927 2087
rect 9893 2053 9907 2067
rect 9953 2073 9967 2087
rect 9833 2033 9847 2047
rect 9893 2033 9907 2047
rect 9933 2033 9947 2047
rect 9813 1953 9827 1967
rect 9793 1933 9807 1947
rect 9793 1893 9807 1907
rect 9753 1613 9767 1627
rect 9833 1793 9847 1807
rect 9993 2173 10007 2187
rect 9973 2053 9987 2067
rect 9953 1993 9967 2007
rect 9933 1893 9947 1907
rect 9953 1893 9967 1907
rect 9853 1773 9867 1787
rect 9853 1713 9867 1727
rect 9833 1613 9847 1627
rect 9753 1593 9767 1607
rect 9733 1573 9747 1587
rect 9713 1533 9727 1547
rect 9753 1513 9767 1527
rect 9713 1433 9727 1447
rect 9713 1293 9727 1307
rect 9773 1233 9787 1247
rect 9753 1213 9767 1227
rect 9733 1173 9747 1187
rect 9693 1153 9707 1167
rect 9693 1133 9707 1147
rect 9533 1113 9547 1127
rect 9573 1113 9587 1127
rect 9633 1113 9647 1127
rect 9673 1113 9687 1127
rect 9553 1093 9567 1107
rect 9533 1073 9547 1087
rect 9453 1053 9467 1067
rect 9333 953 9347 967
rect 9373 953 9387 967
rect 9433 953 9447 967
rect 9393 853 9407 867
rect 9313 673 9327 687
rect 9373 813 9387 827
rect 9353 653 9367 667
rect 9473 953 9487 967
rect 9473 893 9487 907
rect 9453 733 9467 747
rect 9433 693 9447 707
rect 9553 813 9567 827
rect 9613 953 9627 967
rect 9593 833 9607 847
rect 9673 1073 9687 1087
rect 9693 1073 9707 1087
rect 9673 1013 9687 1027
rect 9653 833 9667 847
rect 9573 793 9587 807
rect 9633 793 9647 807
rect 9473 653 9487 667
rect 9513 653 9527 667
rect 9573 653 9587 667
rect 9593 653 9607 667
rect 9333 633 9347 647
rect 9373 633 9387 647
rect 9413 633 9427 647
rect 9313 613 9327 627
rect 9353 613 9367 627
rect 9553 633 9567 647
rect 9413 593 9427 607
rect 9553 573 9567 587
rect 9513 533 9527 547
rect 9433 453 9447 467
rect 9453 353 9467 367
rect 9593 613 9607 627
rect 9593 593 9607 607
rect 9573 353 9587 367
rect 9353 213 9367 227
rect 9473 213 9487 227
rect 9553 213 9567 227
rect 9513 173 9527 187
rect 9393 153 9407 167
rect 9653 573 9667 587
rect 9773 1153 9787 1167
rect 9813 1113 9827 1127
rect 9753 1053 9767 1067
rect 9913 1693 9927 1707
rect 9873 1653 9887 1667
rect 9853 1133 9867 1147
rect 9753 893 9767 907
rect 9833 893 9847 907
rect 9733 793 9747 807
rect 9713 653 9727 667
rect 9793 853 9807 867
rect 9793 833 9807 847
rect 9833 833 9847 847
rect 9773 813 9787 827
rect 9973 1853 9987 1867
rect 10373 3953 10387 3967
rect 10413 3953 10427 3967
rect 10333 3933 10347 3947
rect 10353 3933 10367 3947
rect 10333 3913 10347 3927
rect 10173 3893 10187 3907
rect 10353 3893 10367 3907
rect 10193 3733 10207 3747
rect 10273 3733 10287 3747
rect 10153 3653 10167 3667
rect 10313 3713 10327 3727
rect 10293 3693 10307 3707
rect 10333 3653 10347 3667
rect 10293 3633 10307 3647
rect 10233 3593 10247 3607
rect 10273 3553 10287 3567
rect 10153 3353 10167 3367
rect 10173 3353 10187 3367
rect 10153 3313 10167 3327
rect 10133 3153 10147 3167
rect 10133 3013 10147 3027
rect 10253 3433 10267 3447
rect 10253 3393 10267 3407
rect 10213 3273 10227 3287
rect 10273 3273 10287 3287
rect 10133 2893 10147 2907
rect 10093 2853 10107 2867
rect 10173 2953 10187 2967
rect 10153 2733 10167 2747
rect 10113 2713 10127 2727
rect 10113 2573 10127 2587
rect 10073 2393 10087 2407
rect 10053 2353 10067 2367
rect 10053 2313 10067 2327
rect 10053 2293 10067 2307
rect 10033 2153 10047 2167
rect 10013 1993 10027 2007
rect 10133 2553 10147 2567
rect 10233 3233 10247 3247
rect 10213 3153 10227 3167
rect 10193 2613 10207 2627
rect 10253 3053 10267 3067
rect 10333 3333 10347 3347
rect 10293 3253 10307 3267
rect 10333 3253 10347 3267
rect 10333 3193 10347 3207
rect 10293 3153 10307 3167
rect 10293 3073 10307 3087
rect 10673 4153 10687 4167
rect 10693 4153 10707 4167
rect 10653 4113 10667 4127
rect 10573 4093 10587 4107
rect 10533 4033 10547 4047
rect 10653 4073 10667 4087
rect 10693 4053 10707 4067
rect 10593 4033 10607 4047
rect 10653 4033 10667 4047
rect 10573 3993 10587 4007
rect 10633 4013 10647 4027
rect 10613 3973 10627 3987
rect 10553 3913 10567 3927
rect 10533 3713 10547 3727
rect 10493 3693 10507 3707
rect 10473 3633 10487 3647
rect 10453 3613 10467 3627
rect 10533 3593 10547 3607
rect 10453 3533 10467 3547
rect 10493 3533 10507 3547
rect 10413 3513 10427 3527
rect 10513 3513 10527 3527
rect 10433 3333 10447 3347
rect 10453 3333 10467 3347
rect 10373 3273 10387 3287
rect 10393 3193 10407 3207
rect 10433 3193 10447 3207
rect 10393 3153 10407 3167
rect 10333 3053 10347 3067
rect 10353 3053 10367 3067
rect 10313 2993 10327 3007
rect 10273 2893 10287 2907
rect 10333 2853 10347 2867
rect 10293 2773 10307 2787
rect 10253 2753 10267 2767
rect 10313 2753 10327 2767
rect 10273 2593 10287 2607
rect 10213 2573 10227 2587
rect 10273 2573 10287 2587
rect 10193 2533 10207 2547
rect 10133 2353 10147 2367
rect 10093 2273 10107 2287
rect 10113 2273 10127 2287
rect 10153 2273 10167 2287
rect 10073 2253 10087 2267
rect 10113 2213 10127 2227
rect 10053 1973 10067 1987
rect 10133 2013 10147 2027
rect 10113 1973 10127 1987
rect 10093 1933 10107 1947
rect 10013 1833 10027 1847
rect 10033 1813 10047 1827
rect 10073 1813 10087 1827
rect 10053 1773 10067 1787
rect 10073 1713 10087 1727
rect 10013 1593 10027 1607
rect 9973 1553 9987 1567
rect 9913 1493 9927 1507
rect 9913 1293 9927 1307
rect 9973 1313 9987 1327
rect 9953 1293 9967 1307
rect 10113 1713 10127 1727
rect 10113 1653 10127 1667
rect 10093 1593 10107 1607
rect 10093 1553 10107 1567
rect 10133 1553 10147 1567
rect 10073 1313 10087 1327
rect 10073 1273 10087 1287
rect 10033 1233 10047 1247
rect 9893 1193 9907 1207
rect 9933 1193 9947 1207
rect 9773 633 9787 647
rect 9733 613 9747 627
rect 9693 593 9707 607
rect 9673 353 9687 367
rect 9653 333 9667 347
rect 9733 373 9747 387
rect 9693 233 9707 247
rect 9713 173 9727 187
rect 9853 713 9867 727
rect 9813 573 9827 587
rect 9873 613 9887 627
rect 9853 553 9867 567
rect 9873 393 9887 407
rect 9773 353 9787 367
rect 9833 353 9847 367
rect 10073 1173 10087 1187
rect 10033 1153 10047 1167
rect 9953 1133 9967 1147
rect 9973 1133 9987 1147
rect 9993 1133 10007 1147
rect 9933 1093 9947 1107
rect 9973 1053 9987 1067
rect 9913 893 9927 907
rect 9933 873 9947 887
rect 9913 773 9927 787
rect 10033 1053 10047 1067
rect 10013 853 10027 867
rect 9993 833 10007 847
rect 10033 813 10047 827
rect 9993 793 10007 807
rect 9973 733 9987 747
rect 9933 713 9947 727
rect 9933 653 9947 667
rect 9913 633 9927 647
rect 9993 673 10007 687
rect 10053 653 10067 667
rect 9953 613 9967 627
rect 9993 613 10007 627
rect 10013 513 10027 527
rect 9893 373 9907 387
rect 9993 353 10007 367
rect 10213 2313 10227 2327
rect 10193 2293 10207 2307
rect 10213 2253 10227 2267
rect 10213 2233 10227 2247
rect 10253 2553 10267 2567
rect 10253 2493 10267 2507
rect 10293 2553 10307 2567
rect 10353 2833 10367 2847
rect 10433 3033 10447 3047
rect 10693 3993 10707 4007
rect 10693 3873 10707 3887
rect 10693 3753 10707 3767
rect 10633 3693 10647 3707
rect 10633 3553 10647 3567
rect 10533 3493 10547 3507
rect 10553 3493 10567 3507
rect 10673 3513 10687 3527
rect 10613 3493 10627 3507
rect 10653 3493 10667 3507
rect 10613 3453 10627 3467
rect 10513 3253 10527 3267
rect 10533 3253 10547 3267
rect 10573 3253 10587 3267
rect 10473 3173 10487 3187
rect 10493 3033 10507 3047
rect 10573 3233 10587 3247
rect 10713 3553 10727 3567
rect 10593 3193 10607 3207
rect 10633 3193 10647 3207
rect 10553 3073 10567 3087
rect 10573 3033 10587 3047
rect 10593 3033 10607 3047
rect 10473 3013 10487 3027
rect 10513 3013 10527 3027
rect 10433 2913 10447 2927
rect 10393 2633 10407 2647
rect 10413 2593 10427 2607
rect 10373 2573 10387 2587
rect 10333 2533 10347 2547
rect 10393 2493 10407 2507
rect 10453 2733 10467 2747
rect 10453 2653 10467 2667
rect 10293 2453 10307 2467
rect 10313 2453 10327 2467
rect 10273 2373 10287 2387
rect 10373 2413 10387 2427
rect 10333 2393 10347 2407
rect 10293 2313 10307 2327
rect 10253 2253 10267 2267
rect 10293 2253 10307 2267
rect 10313 2233 10327 2247
rect 10253 2213 10267 2227
rect 10233 2153 10247 2167
rect 10213 2113 10227 2127
rect 10193 2033 10207 2047
rect 10193 1953 10207 1967
rect 10213 1893 10227 1907
rect 10273 2133 10287 2147
rect 10313 2073 10327 2087
rect 10293 2033 10307 2047
rect 10233 1873 10247 1887
rect 10233 1813 10247 1827
rect 10273 1793 10287 1807
rect 10353 2273 10367 2287
rect 10333 1773 10347 1787
rect 10293 1713 10307 1727
rect 10253 1633 10267 1647
rect 10373 1833 10387 1847
rect 10173 1553 10187 1567
rect 10193 1553 10207 1567
rect 10353 1613 10367 1627
rect 10293 1573 10307 1587
rect 10273 1513 10287 1527
rect 10253 1453 10267 1467
rect 10193 1433 10207 1447
rect 10213 1433 10227 1447
rect 10153 1373 10167 1387
rect 10133 1293 10147 1307
rect 10213 1293 10227 1307
rect 10153 1273 10167 1287
rect 10113 1213 10127 1227
rect 10133 1093 10147 1107
rect 10153 1093 10167 1107
rect 10313 1313 10327 1327
rect 10353 1313 10367 1327
rect 10333 1293 10347 1307
rect 10293 1273 10307 1287
rect 10293 1233 10307 1247
rect 10353 1233 10367 1247
rect 10273 1033 10287 1047
rect 10233 1013 10247 1027
rect 10233 993 10247 1007
rect 10193 853 10207 867
rect 10253 833 10267 847
rect 10253 753 10267 767
rect 10233 693 10247 707
rect 10093 653 10107 667
rect 10113 653 10127 667
rect 10153 653 10167 667
rect 10073 633 10087 647
rect 10093 633 10107 647
rect 10133 633 10147 647
rect 10113 613 10127 627
rect 10173 633 10187 647
rect 10213 633 10227 647
rect 10173 553 10187 567
rect 10113 393 10127 407
rect 10053 353 10067 367
rect 10113 353 10127 367
rect 9893 293 9907 307
rect 9853 273 9867 287
rect 9873 253 9887 267
rect 9913 193 9927 207
rect 9333 133 9347 147
rect 9573 133 9587 147
rect 10013 313 10027 327
rect 10033 313 10047 327
rect 10073 273 10087 287
rect 10133 273 10147 287
rect 10073 173 10087 187
rect 10113 153 10127 167
rect 10253 673 10267 687
rect 10253 613 10267 627
rect 10513 2993 10527 3007
rect 10493 2573 10507 2587
rect 10473 2493 10487 2507
rect 10453 2433 10467 2447
rect 10433 2313 10447 2327
rect 10433 2133 10447 2147
rect 10593 2993 10607 3007
rect 10693 3073 10707 3087
rect 10633 2893 10647 2907
rect 10593 2813 10607 2827
rect 10653 2813 10667 2827
rect 10613 2773 10627 2787
rect 10593 2733 10607 2747
rect 10573 2673 10587 2687
rect 10633 2673 10647 2687
rect 10553 2573 10567 2587
rect 10613 2633 10627 2647
rect 10533 2553 10547 2567
rect 10553 2533 10567 2547
rect 10593 2513 10607 2527
rect 10553 2393 10567 2407
rect 10533 2313 10547 2327
rect 10493 2273 10507 2287
rect 10513 2273 10527 2287
rect 10513 2233 10527 2247
rect 10493 2133 10507 2147
rect 10473 2073 10487 2087
rect 10453 2053 10467 2067
rect 10413 2013 10427 2027
rect 10533 2073 10547 2087
rect 10513 1833 10527 1847
rect 10453 1753 10467 1767
rect 10453 1633 10467 1647
rect 10493 1773 10507 1787
rect 10493 1753 10507 1767
rect 10493 1633 10507 1647
rect 10493 1573 10507 1587
rect 10453 1393 10467 1407
rect 10433 1373 10447 1387
rect 10413 1293 10427 1307
rect 10393 1173 10407 1187
rect 10633 2553 10647 2567
rect 10653 2333 10667 2347
rect 10833 4193 10847 4207
rect 10873 4193 10887 4207
rect 10913 4193 10927 4207
rect 10813 4093 10827 4107
rect 10753 4033 10767 4047
rect 10773 4013 10787 4027
rect 10793 3993 10807 4007
rect 10753 3953 10767 3967
rect 10793 3853 10807 3867
rect 10893 4153 10907 4167
rect 10993 4093 11007 4107
rect 10853 3973 10867 3987
rect 11013 3973 11027 3987
rect 10973 3913 10987 3927
rect 10933 3853 10947 3867
rect 11133 6913 11147 6927
rect 11113 6813 11127 6827
rect 11173 6893 11187 6907
rect 11213 6893 11227 6907
rect 11193 6853 11207 6867
rect 11373 7053 11387 7067
rect 11333 6913 11347 6927
rect 11313 6873 11327 6887
rect 11373 6893 11387 6907
rect 11393 6873 11407 6887
rect 11293 6753 11307 6767
rect 11393 6853 11407 6867
rect 11353 6813 11367 6827
rect 11433 7573 11447 7587
rect 11453 7513 11467 7527
rect 11453 7373 11467 7387
rect 11433 7353 11447 7367
rect 11413 6633 11427 6647
rect 11313 6593 11327 6607
rect 11353 6593 11367 6607
rect 11393 6593 11407 6607
rect 11113 6553 11127 6567
rect 11153 6553 11167 6567
rect 11233 6433 11247 6447
rect 11193 6413 11207 6427
rect 11213 6393 11227 6407
rect 11193 6373 11207 6387
rect 11373 6573 11387 6587
rect 11413 6573 11427 6587
rect 11413 6553 11427 6567
rect 11413 6533 11427 6547
rect 11373 6433 11387 6447
rect 11353 6393 11367 6407
rect 11153 6333 11167 6347
rect 11093 6313 11107 6327
rect 11093 6153 11107 6167
rect 11153 6133 11167 6147
rect 11133 6113 11147 6127
rect 11113 6093 11127 6107
rect 11073 6073 11087 6087
rect 11093 5993 11107 6007
rect 11353 6113 11367 6127
rect 11153 6093 11167 6107
rect 11333 6093 11347 6107
rect 11153 6073 11167 6087
rect 11253 6073 11267 6087
rect 11293 6073 11307 6087
rect 11093 5933 11107 5947
rect 11133 5933 11147 5947
rect 11113 5913 11127 5927
rect 11173 6013 11187 6027
rect 11193 5933 11207 5947
rect 11133 5893 11147 5907
rect 11173 5893 11187 5907
rect 11073 5633 11087 5647
rect 11113 5613 11127 5627
rect 11093 5473 11107 5487
rect 11353 6033 11367 6047
rect 11293 6013 11307 6027
rect 11333 5913 11347 5927
rect 11313 5893 11327 5907
rect 11313 5653 11327 5667
rect 11413 6413 11427 6427
rect 11513 8513 11527 8527
rect 11493 8493 11507 8507
rect 11493 8433 11507 8447
rect 11493 8313 11507 8327
rect 11613 8833 11627 8847
rect 11633 8813 11647 8827
rect 11653 8793 11667 8807
rect 11653 8633 11667 8647
rect 11633 8593 11647 8607
rect 11593 8373 11607 8387
rect 11573 8053 11587 8067
rect 11533 8013 11547 8027
rect 11573 8013 11587 8027
rect 11513 7973 11527 7987
rect 11553 7973 11567 7987
rect 11513 7853 11527 7867
rect 11493 7833 11507 7847
rect 11573 7893 11587 7907
rect 11493 7793 11507 7807
rect 11533 7793 11547 7807
rect 11533 7773 11547 7787
rect 11473 7353 11487 7367
rect 11493 7333 11507 7347
rect 11573 7793 11587 7807
rect 11553 7553 11567 7567
rect 11693 9753 11707 9767
rect 11693 9713 11707 9727
rect 11753 9793 11767 9807
rect 11733 9753 11747 9767
rect 11733 9733 11747 9747
rect 11773 9733 11787 9747
rect 11713 9653 11727 9667
rect 11753 9713 11767 9727
rect 11793 9713 11807 9727
rect 11733 9613 11747 9627
rect 11753 9513 11767 9527
rect 11693 9493 11707 9507
rect 11733 9473 11747 9487
rect 11773 9473 11787 9487
rect 11713 9433 11727 9447
rect 11753 9433 11767 9447
rect 11693 9293 11707 9307
rect 11693 9273 11707 9287
rect 11753 9273 11767 9287
rect 11813 9613 11827 9627
rect 11793 9453 11807 9467
rect 11813 9273 11827 9287
rect 11733 9253 11747 9267
rect 11773 9253 11787 9267
rect 11793 9193 11807 9207
rect 11773 9013 11787 9027
rect 11753 8973 11767 8987
rect 11713 8933 11727 8947
rect 11733 8893 11747 8907
rect 11753 8893 11767 8907
rect 11813 8953 11827 8967
rect 11733 8873 11747 8887
rect 11793 8873 11807 8887
rect 11713 8813 11727 8827
rect 11713 8653 11727 8667
rect 11793 8853 11807 8867
rect 11773 8833 11787 8847
rect 11753 8793 11767 8807
rect 11813 8793 11827 8807
rect 11733 8533 11747 8547
rect 11693 8493 11707 8507
rect 11733 8493 11747 8507
rect 11813 8753 11827 8767
rect 11773 8613 11787 8627
rect 11793 8533 11807 8547
rect 11773 8493 11787 8507
rect 11713 8413 11727 8427
rect 11673 8393 11687 8407
rect 11673 8333 11687 8347
rect 11713 8333 11727 8347
rect 11753 8333 11767 8347
rect 11773 8313 11787 8327
rect 11733 8253 11747 8267
rect 11713 8133 11727 8147
rect 11673 8093 11687 8107
rect 11693 8053 11707 8067
rect 11653 8033 11667 8047
rect 11713 8033 11727 8047
rect 11633 8013 11647 8027
rect 11733 7893 11747 7907
rect 11773 7873 11787 7887
rect 11713 7793 11727 7807
rect 11733 7773 11747 7787
rect 11653 7633 11667 7647
rect 11613 7613 11627 7627
rect 11673 7613 11687 7627
rect 11633 7553 11647 7567
rect 11613 7533 11627 7547
rect 11733 7393 11747 7407
rect 11473 7313 11487 7327
rect 11533 7313 11547 7327
rect 11613 7313 11627 7327
rect 11533 7273 11547 7287
rect 11553 7073 11567 7087
rect 11513 7053 11527 7067
rect 11593 7033 11607 7047
rect 11573 6933 11587 6947
rect 11533 6913 11547 6927
rect 11613 6813 11627 6827
rect 11473 6633 11487 6647
rect 11453 6593 11467 6607
rect 11453 6513 11467 6527
rect 11393 6393 11407 6407
rect 11433 6393 11447 6407
rect 11413 6153 11427 6167
rect 11193 5613 11207 5627
rect 11133 5453 11147 5467
rect 11153 5453 11167 5467
rect 11253 5453 11267 5467
rect 11113 5433 11127 5447
rect 11193 5433 11207 5447
rect 11213 5433 11227 5447
rect 11133 5413 11147 5427
rect 11173 5393 11187 5407
rect 11213 5173 11227 5187
rect 11093 5153 11107 5167
rect 11153 5153 11167 5167
rect 11173 5113 11187 5127
rect 11133 5033 11147 5047
rect 11193 5033 11207 5047
rect 11113 5013 11127 5027
rect 11133 5013 11147 5027
rect 11093 4973 11107 4987
rect 11173 4953 11187 4967
rect 11093 4933 11107 4947
rect 11153 4933 11167 4947
rect 11233 4953 11247 4967
rect 11053 4673 11067 4687
rect 11213 4673 11227 4687
rect 11133 4653 11147 4667
rect 11373 5453 11387 5467
rect 11373 5433 11387 5447
rect 11393 5433 11407 5447
rect 11273 5413 11287 5427
rect 11353 5413 11367 5427
rect 11273 5253 11287 5267
rect 11293 5173 11307 5187
rect 11273 5153 11287 5167
rect 11313 5153 11327 5167
rect 11373 5173 11387 5187
rect 11353 5133 11367 5147
rect 11393 4973 11407 4987
rect 11353 4753 11367 4767
rect 11273 4713 11287 4727
rect 11313 4673 11327 4687
rect 11293 4653 11307 4667
rect 11233 4613 11247 4627
rect 11093 4573 11107 4587
rect 11133 4553 11147 4567
rect 11193 4493 11207 4507
rect 11333 4573 11347 4587
rect 11153 4473 11167 4487
rect 11313 4473 11327 4487
rect 11053 4453 11067 4467
rect 11133 4453 11147 4467
rect 11173 4453 11187 4467
rect 11213 4453 11227 4467
rect 11213 4433 11227 4447
rect 11393 4633 11407 4647
rect 11353 4553 11367 4567
rect 11373 4453 11387 4467
rect 11393 4433 11407 4447
rect 11053 4213 11067 4227
rect 11153 4213 11167 4227
rect 11233 4213 11247 4227
rect 11073 4193 11087 4207
rect 11093 4193 11107 4207
rect 11033 3793 11047 3807
rect 10893 3733 10907 3747
rect 11013 3733 11027 3747
rect 10853 3713 10867 3727
rect 10833 3653 10847 3667
rect 10853 3633 10867 3647
rect 10913 3693 10927 3707
rect 10893 3653 10907 3667
rect 10873 3613 10887 3627
rect 10833 3533 10847 3547
rect 10813 3513 10827 3527
rect 10793 3493 10807 3507
rect 10873 3493 10887 3507
rect 10773 3273 10787 3287
rect 10753 3173 10767 3187
rect 10733 3153 10747 3167
rect 10733 3113 10747 3127
rect 10933 3573 10947 3587
rect 10913 3513 10927 3527
rect 10913 3393 10927 3407
rect 10893 3353 10907 3367
rect 10773 3073 10787 3087
rect 10873 3213 10887 3227
rect 10833 3133 10847 3147
rect 10833 3113 10847 3127
rect 10793 3033 10807 3047
rect 10753 2993 10767 3007
rect 10753 2973 10767 2987
rect 10733 2773 10747 2787
rect 10793 2793 10807 2807
rect 11053 3693 11067 3707
rect 11013 3553 11027 3567
rect 11053 3513 11067 3527
rect 11113 4153 11127 4167
rect 11253 4193 11267 4207
rect 11293 4193 11307 4207
rect 11393 4193 11407 4207
rect 11273 4173 11287 4187
rect 11273 4113 11287 4127
rect 11253 4033 11267 4047
rect 11313 4013 11327 4027
rect 11333 4013 11347 4027
rect 11173 3993 11187 4007
rect 11213 3993 11227 4007
rect 11253 3993 11267 4007
rect 11193 3973 11207 3987
rect 11133 3953 11147 3967
rect 11113 3693 11127 3707
rect 11273 3673 11287 3687
rect 11093 3653 11107 3667
rect 11073 3373 11087 3387
rect 11033 3353 11047 3367
rect 10993 3313 11007 3327
rect 10953 3293 10967 3307
rect 11033 3273 11047 3287
rect 10933 3113 10947 3127
rect 10913 3073 10927 3087
rect 10993 3153 11007 3167
rect 10933 3033 10947 3047
rect 10973 3033 10987 3047
rect 10973 3013 10987 3027
rect 10913 2993 10927 3007
rect 10953 2993 10967 3007
rect 10873 2893 10887 2907
rect 10873 2813 10887 2827
rect 10833 2753 10847 2767
rect 11013 3033 11027 3047
rect 11013 2853 11027 2867
rect 11273 3573 11287 3587
rect 11193 3513 11207 3527
rect 11233 3513 11247 3527
rect 11213 3493 11227 3507
rect 11253 3493 11267 3507
rect 11233 3473 11247 3487
rect 11193 3453 11207 3467
rect 11213 3373 11227 3387
rect 11173 3273 11187 3287
rect 11133 3233 11147 3247
rect 11153 3193 11167 3207
rect 11093 3113 11107 3127
rect 11133 3113 11147 3127
rect 11073 3073 11087 3087
rect 11053 3013 11067 3027
rect 10893 2753 10907 2767
rect 10753 2653 10767 2667
rect 10733 2633 10747 2647
rect 10773 2593 10787 2607
rect 10773 2573 10787 2587
rect 10733 2553 10747 2567
rect 10693 2533 10707 2547
rect 10713 2513 10727 2527
rect 10753 2513 10767 2527
rect 10773 2493 10787 2507
rect 10753 2353 10767 2367
rect 10673 2313 10687 2327
rect 10653 2253 10667 2267
rect 10713 2273 10727 2287
rect 10693 2253 10707 2267
rect 10733 2253 10747 2267
rect 10673 2173 10687 2187
rect 10653 2153 10667 2167
rect 10613 2093 10627 2107
rect 10693 2093 10707 2107
rect 10553 2053 10567 2067
rect 10533 1493 10547 1507
rect 10553 1413 10567 1427
rect 10473 1373 10487 1387
rect 10513 1373 10527 1387
rect 10453 1313 10467 1327
rect 10393 1133 10407 1147
rect 10433 1133 10447 1147
rect 10333 1093 10347 1107
rect 10313 973 10327 987
rect 10293 813 10307 827
rect 10353 933 10367 947
rect 10293 733 10307 747
rect 10373 813 10387 827
rect 10333 633 10347 647
rect 10353 633 10367 647
rect 10313 613 10327 627
rect 10493 1333 10507 1347
rect 10513 1313 10527 1327
rect 10553 1293 10567 1307
rect 10633 2053 10647 2067
rect 10593 2013 10607 2027
rect 10573 1213 10587 1227
rect 10573 1193 10587 1207
rect 10533 1153 10547 1167
rect 10573 1133 10587 1147
rect 10513 1093 10527 1107
rect 10673 1993 10687 2007
rect 10653 1793 10667 1807
rect 10613 1613 10627 1627
rect 10713 1833 10727 1847
rect 10693 1813 10707 1827
rect 10693 1733 10707 1747
rect 10673 1613 10687 1627
rect 10633 1573 10647 1587
rect 10613 1493 10627 1507
rect 10593 813 10607 827
rect 10513 713 10527 727
rect 10533 713 10547 727
rect 10553 693 10567 707
rect 10653 1453 10667 1467
rect 10633 1373 10647 1387
rect 10633 1133 10647 1147
rect 10633 933 10647 947
rect 10733 1513 10747 1527
rect 10713 1293 10727 1307
rect 10733 1293 10747 1307
rect 10673 1273 10687 1287
rect 10653 793 10667 807
rect 10713 1233 10727 1247
rect 10713 1113 10727 1127
rect 10693 1053 10707 1067
rect 10733 1033 10747 1047
rect 10733 1013 10747 1027
rect 10693 993 10707 1007
rect 10693 913 10707 927
rect 10833 2693 10847 2707
rect 10953 2573 10967 2587
rect 10853 2533 10867 2547
rect 10833 2513 10847 2527
rect 10913 2533 10927 2547
rect 10853 2473 10867 2487
rect 10853 2313 10867 2327
rect 10913 2473 10927 2487
rect 10813 2293 10827 2307
rect 10893 2293 10907 2307
rect 10833 2273 10847 2287
rect 10873 2273 10887 2287
rect 10933 2273 10947 2287
rect 10853 2253 10867 2267
rect 10893 2213 10907 2227
rect 10833 2173 10847 2187
rect 10953 2133 10967 2147
rect 10913 2113 10927 2127
rect 10933 2113 10947 2127
rect 10813 2093 10827 2107
rect 10893 2093 10907 2107
rect 10813 2053 10827 2067
rect 10833 2053 10847 2067
rect 10793 1793 10807 1807
rect 10853 1913 10867 1927
rect 10913 1833 10927 1847
rect 10873 1793 10887 1807
rect 10893 1793 10907 1807
rect 10913 1653 10927 1667
rect 10873 1553 10887 1567
rect 10833 1333 10847 1347
rect 11093 3053 11107 3067
rect 11073 2953 11087 2967
rect 11073 2933 11087 2947
rect 11073 2853 11087 2867
rect 11053 2753 11067 2767
rect 11093 2813 11107 2827
rect 11033 2713 11047 2727
rect 11073 2713 11087 2727
rect 10993 2673 11007 2687
rect 11033 2673 11047 2687
rect 10993 2633 11007 2647
rect 11013 2253 11027 2267
rect 11013 2193 11027 2207
rect 10973 2093 10987 2107
rect 10993 2093 11007 2107
rect 10973 2073 10987 2087
rect 11073 2633 11087 2647
rect 11113 2753 11127 2767
rect 11153 3073 11167 3087
rect 11173 3053 11187 3067
rect 11193 2973 11207 2987
rect 11153 2953 11167 2967
rect 11213 2773 11227 2787
rect 11213 2733 11227 2747
rect 11193 2713 11207 2727
rect 11153 2613 11167 2627
rect 11213 2613 11227 2627
rect 11133 2593 11147 2607
rect 11093 2573 11107 2587
rect 11113 2573 11127 2587
rect 11113 2553 11127 2567
rect 11173 2593 11187 2607
rect 11093 2513 11107 2527
rect 11133 2433 11147 2447
rect 11093 2353 11107 2367
rect 11113 2293 11127 2307
rect 11073 2273 11087 2287
rect 11053 2253 11067 2267
rect 11153 2213 11167 2227
rect 11093 2193 11107 2207
rect 11093 2153 11107 2167
rect 11093 2093 11107 2107
rect 11213 2573 11227 2587
rect 11173 2113 11187 2127
rect 11373 3993 11387 4007
rect 11353 3973 11367 3987
rect 11573 6613 11587 6627
rect 11513 6573 11527 6587
rect 11593 6573 11607 6587
rect 11553 6513 11567 6527
rect 11533 6453 11547 6467
rect 11513 6393 11527 6407
rect 11473 6153 11487 6167
rect 11553 6413 11567 6427
rect 11533 6353 11547 6367
rect 11473 6133 11487 6147
rect 11513 6133 11527 6147
rect 11493 6113 11507 6127
rect 11473 6053 11487 6067
rect 11453 5973 11467 5987
rect 11513 5973 11527 5987
rect 11493 5953 11507 5967
rect 11573 6393 11587 6407
rect 11673 7353 11687 7367
rect 11693 7313 11707 7327
rect 11673 7213 11687 7227
rect 11793 7853 11807 7867
rect 11813 7773 11827 7787
rect 11913 10373 11927 10387
rect 11893 10353 11907 10367
rect 11873 10193 11887 10207
rect 11893 10173 11907 10187
rect 11953 10373 11967 10387
rect 11933 10313 11947 10327
rect 11953 10293 11967 10307
rect 11933 10273 11947 10287
rect 12013 10913 12027 10927
rect 12013 10893 12027 10907
rect 12053 11313 12067 11327
rect 12053 11253 12067 11267
rect 12053 11213 12067 11227
rect 12053 11133 12067 11147
rect 12193 11813 12207 11827
rect 12093 11793 12107 11807
rect 12153 11693 12167 11707
rect 12133 11673 12147 11687
rect 12173 11653 12187 11667
rect 12153 11513 12167 11527
rect 12113 11493 12127 11507
rect 12093 11413 12107 11427
rect 12133 11413 12147 11427
rect 12113 11353 12127 11367
rect 12113 10993 12127 11007
rect 12093 10913 12107 10927
rect 12073 10893 12087 10907
rect 12053 10813 12067 10827
rect 12033 10713 12047 10727
rect 12133 10973 12147 10987
rect 12033 10693 12047 10707
rect 12013 10633 12027 10647
rect 12053 10673 12067 10687
rect 12133 10693 12147 10707
rect 12093 10653 12107 10667
rect 12113 10633 12127 10647
rect 12053 10473 12067 10487
rect 12093 10473 12107 10487
rect 12033 10453 12047 10467
rect 12033 10433 12047 10447
rect 11993 10333 12007 10347
rect 11973 10273 11987 10287
rect 11993 10273 12007 10287
rect 11973 10233 11987 10247
rect 11973 10153 11987 10167
rect 11913 10133 11927 10147
rect 11933 9913 11947 9927
rect 11893 9773 11907 9787
rect 11873 9673 11887 9687
rect 12053 10413 12067 10427
rect 12133 10593 12147 10607
rect 12013 10253 12027 10267
rect 12033 10253 12047 10267
rect 12013 10133 12027 10147
rect 11993 9893 12007 9907
rect 11993 9773 12007 9787
rect 11993 9753 12007 9767
rect 11933 9733 11947 9747
rect 11973 9733 11987 9747
rect 11913 9713 11927 9727
rect 11953 9713 11967 9727
rect 11933 9673 11947 9687
rect 11913 9513 11927 9527
rect 11873 9493 11887 9507
rect 11913 9493 11927 9507
rect 11873 9453 11887 9467
rect 11853 9273 11867 9287
rect 11893 9433 11907 9447
rect 11893 9293 11907 9307
rect 11993 9413 12007 9427
rect 11933 9213 11947 9227
rect 11933 9013 11947 9027
rect 11893 8973 11907 8987
rect 11873 8753 11887 8767
rect 12133 10253 12147 10267
rect 12173 11253 12187 11267
rect 12173 10953 12187 10967
rect 12173 10913 12187 10927
rect 12173 10573 12187 10587
rect 12153 10233 12167 10247
rect 12113 10213 12127 10227
rect 12153 10213 12167 10227
rect 12033 9933 12047 9947
rect 12073 9913 12087 9927
rect 12053 9793 12067 9807
rect 12133 9773 12147 9787
rect 12073 9693 12087 9707
rect 12093 9533 12107 9547
rect 12053 9493 12067 9507
rect 12033 9433 12047 9447
rect 11973 9273 11987 9287
rect 12013 9273 12027 9287
rect 11993 9253 12007 9267
rect 11953 8933 11967 8947
rect 11953 8913 11967 8927
rect 11933 8893 11947 8907
rect 11913 8833 11927 8847
rect 11893 8613 11907 8627
rect 11973 8793 11987 8807
rect 12013 9013 12027 9027
rect 11953 8773 11967 8787
rect 11993 8773 12007 8787
rect 11913 8553 11927 8567
rect 11853 8533 11867 8547
rect 11933 8533 11947 8547
rect 11873 8493 11887 8507
rect 11973 8553 11987 8567
rect 11953 8493 11967 8507
rect 11853 8473 11867 8487
rect 11853 8253 11867 8267
rect 11913 8393 11927 8407
rect 11913 8333 11927 8347
rect 12153 9713 12167 9727
rect 12073 9373 12087 9387
rect 12073 9273 12087 9287
rect 12053 9233 12067 9247
rect 12113 9273 12127 9287
rect 12173 9273 12187 9287
rect 12093 9213 12107 9227
rect 12033 8973 12047 8987
rect 12033 8953 12047 8967
rect 12153 9253 12167 9267
rect 12133 9233 12147 9247
rect 12173 9213 12187 9227
rect 12113 9013 12127 9027
rect 12073 8953 12087 8967
rect 12053 8793 12067 8807
rect 12113 8833 12127 8847
rect 12133 8813 12147 8827
rect 12153 8793 12167 8807
rect 12093 8773 12107 8787
rect 12133 8773 12147 8787
rect 12113 8533 12127 8547
rect 12033 8513 12047 8527
rect 12073 8473 12087 8487
rect 12013 8433 12027 8447
rect 11953 8333 11967 8347
rect 12073 8333 12087 8347
rect 12113 8333 12127 8347
rect 11893 8313 11907 8327
rect 11933 8313 11947 8327
rect 12093 8313 12107 8327
rect 11913 8293 11927 8307
rect 11953 8293 11967 8307
rect 11873 8233 11887 8247
rect 11853 8093 11867 8107
rect 11873 8093 11887 8107
rect 11893 7993 11907 8007
rect 11913 7813 11927 7827
rect 11853 7793 11867 7807
rect 11893 7793 11907 7807
rect 11933 7793 11947 7807
rect 11793 7573 11807 7587
rect 11833 7573 11847 7587
rect 11773 7213 11787 7227
rect 11773 7193 11787 7207
rect 11753 7173 11767 7187
rect 11713 7053 11727 7067
rect 11733 7033 11747 7047
rect 11693 6913 11707 6927
rect 11733 6873 11747 6887
rect 11713 6853 11727 6867
rect 11753 6853 11767 6867
rect 11813 7553 11827 7567
rect 11893 7573 11907 7587
rect 11833 7533 11847 7547
rect 12033 8193 12047 8207
rect 12013 8053 12027 8067
rect 11973 7853 11987 7867
rect 11993 7853 12007 7867
rect 11973 7793 11987 7807
rect 11973 7653 11987 7667
rect 12093 8013 12107 8027
rect 12053 7893 12067 7907
rect 12013 7793 12027 7807
rect 11993 7573 12007 7587
rect 12133 7913 12147 7927
rect 12113 7893 12127 7907
rect 12093 7853 12107 7867
rect 12093 7833 12107 7847
rect 12073 7793 12087 7807
rect 11933 7553 11947 7567
rect 11953 7553 11967 7567
rect 11973 7553 11987 7567
rect 12013 7553 12027 7567
rect 11793 6633 11807 6647
rect 11753 6593 11767 6607
rect 11773 6573 11787 6587
rect 11733 6553 11747 6567
rect 11793 6473 11807 6487
rect 11793 6413 11807 6427
rect 11713 6373 11727 6387
rect 11753 6373 11767 6387
rect 11873 7473 11887 7487
rect 11893 7393 11907 7407
rect 12033 7473 12047 7487
rect 11953 7453 11967 7467
rect 11933 7373 11947 7387
rect 11913 7333 11927 7347
rect 11873 7233 11887 7247
rect 12013 7373 12027 7387
rect 12013 7313 12027 7327
rect 12073 7473 12087 7487
rect 12073 7453 12087 7467
rect 12053 7433 12067 7447
rect 12053 7353 12067 7367
rect 12093 7313 12107 7327
rect 11833 6633 11847 6647
rect 11673 6333 11687 6347
rect 11753 6333 11767 6347
rect 11773 6333 11787 6347
rect 11813 6333 11827 6347
rect 11613 6133 11627 6147
rect 11653 6133 11667 6147
rect 11593 6093 11607 6107
rect 11633 6113 11647 6127
rect 11673 6113 11687 6127
rect 11613 6073 11627 6087
rect 11693 6093 11707 6107
rect 11653 6073 11667 6087
rect 11633 6053 11647 6067
rect 11713 6033 11727 6047
rect 11593 5973 11607 5987
rect 11553 5933 11567 5947
rect 11513 5913 11527 5927
rect 11533 5893 11547 5907
rect 11473 5773 11487 5787
rect 11573 5713 11587 5727
rect 11493 5653 11507 5667
rect 11533 5653 11547 5667
rect 11553 5633 11567 5647
rect 11673 5953 11687 5967
rect 11653 5913 11667 5927
rect 11713 5933 11727 5947
rect 11733 5913 11747 5927
rect 11593 5653 11607 5667
rect 11513 5613 11527 5627
rect 11573 5613 11587 5627
rect 11693 5893 11707 5907
rect 11673 5693 11687 5707
rect 11713 5673 11727 5687
rect 11693 5633 11707 5647
rect 11653 5573 11667 5587
rect 11713 5573 11727 5587
rect 11473 5453 11487 5467
rect 11653 5453 11667 5467
rect 11453 5393 11467 5407
rect 11553 5433 11567 5447
rect 11533 5413 11547 5427
rect 11493 5393 11507 5407
rect 11573 5393 11587 5407
rect 11473 5173 11487 5187
rect 11633 5413 11647 5427
rect 11553 5353 11567 5367
rect 11613 5353 11627 5367
rect 11613 5193 11627 5207
rect 11473 5113 11487 5127
rect 11513 4993 11527 5007
rect 11553 4993 11567 5007
rect 11493 4973 11507 4987
rect 11533 4973 11547 4987
rect 11533 4953 11547 4967
rect 11453 4933 11467 4947
rect 11513 4933 11527 4947
rect 11733 5413 11747 5427
rect 11713 5233 11727 5247
rect 11653 5193 11667 5207
rect 11693 5153 11707 5167
rect 11673 4993 11687 5007
rect 11653 4953 11667 4967
rect 11633 4933 11647 4947
rect 11653 4933 11667 4947
rect 11613 4733 11627 4747
rect 11613 4713 11627 4727
rect 11513 4673 11527 4687
rect 11453 4633 11467 4647
rect 11533 4533 11547 4547
rect 11513 4473 11527 4487
rect 11553 4513 11567 4527
rect 11573 4433 11587 4447
rect 11713 4933 11727 4947
rect 11733 4913 11747 4927
rect 11693 4673 11707 4687
rect 11733 4673 11747 4687
rect 11633 4653 11647 4667
rect 11673 4653 11687 4667
rect 11673 4513 11687 4527
rect 11713 4493 11727 4507
rect 11733 4433 11747 4447
rect 11613 4413 11627 4427
rect 11533 4393 11547 4407
rect 11433 4213 11447 4227
rect 11493 4213 11507 4227
rect 11473 4153 11487 4167
rect 11473 4133 11487 4147
rect 11433 3973 11447 3987
rect 11353 3553 11367 3567
rect 11373 3513 11387 3527
rect 11353 3493 11367 3507
rect 11313 3453 11327 3467
rect 11253 3293 11267 3307
rect 11273 3253 11287 3267
rect 11253 3193 11267 3207
rect 11253 3133 11267 3147
rect 11233 2513 11247 2527
rect 11293 3153 11307 3167
rect 11453 3653 11467 3667
rect 11473 3653 11487 3667
rect 11413 3573 11427 3587
rect 11433 3513 11447 3527
rect 11413 3493 11427 3507
rect 11433 3473 11447 3487
rect 11373 3333 11387 3347
rect 11393 3333 11407 3347
rect 11393 3293 11407 3307
rect 11333 3213 11347 3227
rect 11353 3173 11367 3187
rect 11393 3173 11407 3187
rect 11313 3113 11327 3127
rect 11373 3113 11387 3127
rect 11333 3053 11347 3067
rect 11293 3033 11307 3047
rect 11353 3033 11367 3047
rect 11373 3013 11387 3027
rect 11293 2993 11307 3007
rect 11313 2993 11327 3007
rect 11273 2853 11287 2867
rect 11273 2773 11287 2787
rect 11373 2893 11387 2907
rect 11413 3033 11427 3047
rect 11453 3453 11467 3467
rect 11473 3273 11487 3287
rect 11453 3033 11467 3047
rect 11433 2973 11447 2987
rect 11413 2873 11427 2887
rect 11413 2813 11427 2827
rect 11393 2773 11407 2787
rect 11393 2733 11407 2747
rect 11433 2733 11447 2747
rect 11373 2693 11387 2707
rect 11313 2593 11327 2607
rect 11293 2573 11307 2587
rect 11273 2553 11287 2567
rect 11293 2553 11307 2567
rect 11253 2493 11267 2507
rect 11213 2433 11227 2447
rect 11213 2413 11227 2427
rect 10953 2053 10967 2067
rect 10993 2053 11007 2067
rect 11033 2053 11047 2067
rect 11093 2053 11107 2067
rect 11193 2073 11207 2087
rect 11153 2053 11167 2067
rect 11193 2053 11207 2067
rect 10993 2033 11007 2047
rect 11113 2033 11127 2047
rect 10973 1813 10987 1827
rect 10933 1373 10947 1387
rect 10933 1333 10947 1347
rect 10873 1293 10887 1307
rect 11073 1893 11087 1907
rect 11033 1813 11047 1827
rect 11253 2313 11267 2327
rect 11233 2013 11247 2027
rect 11213 1853 11227 1867
rect 11133 1833 11147 1847
rect 11053 1793 11067 1807
rect 11353 2533 11367 2547
rect 11313 2493 11327 2507
rect 11353 2453 11367 2467
rect 11313 2273 11327 2287
rect 11293 2253 11307 2267
rect 11273 2233 11287 2247
rect 11313 2233 11327 2247
rect 11333 2233 11347 2247
rect 11293 2073 11307 2087
rect 11273 1793 11287 1807
rect 11193 1773 11207 1787
rect 11213 1773 11227 1787
rect 11133 1693 11147 1707
rect 11073 1673 11087 1687
rect 11033 1613 11047 1627
rect 11013 1593 11027 1607
rect 11093 1593 11107 1607
rect 11053 1573 11067 1587
rect 10973 1253 10987 1267
rect 10913 1193 10927 1207
rect 10953 1193 10967 1207
rect 10773 913 10787 927
rect 10933 1093 10947 1107
rect 10893 1013 10907 1027
rect 10913 993 10927 1007
rect 10953 993 10967 1007
rect 10773 853 10787 867
rect 10853 853 10867 867
rect 10753 793 10767 807
rect 10733 733 10747 747
rect 10693 673 10707 687
rect 10673 653 10687 667
rect 10473 613 10487 627
rect 10533 613 10547 627
rect 10573 613 10587 627
rect 10613 613 10627 627
rect 10453 573 10467 587
rect 10373 413 10387 427
rect 10273 373 10287 387
rect 10253 353 10267 367
rect 10213 253 10227 267
rect 10373 373 10387 387
rect 10413 353 10427 367
rect 10553 433 10567 447
rect 10533 373 10547 387
rect 10433 333 10447 347
rect 10473 333 10487 347
rect 10533 333 10547 347
rect 10473 313 10487 327
rect 10473 213 10487 227
rect 10393 173 10407 187
rect 10433 173 10447 187
rect 10513 173 10527 187
rect 9993 133 10007 147
rect 10053 133 10067 147
rect 10093 133 10107 147
rect 10133 133 10147 147
rect 10453 133 10467 147
rect 10713 433 10727 447
rect 10673 393 10687 407
rect 10573 353 10587 367
rect 10633 353 10647 367
rect 10653 333 10667 347
rect 10693 333 10707 347
rect 10613 313 10627 327
rect 10613 193 10627 207
rect 10653 173 10667 187
rect 10953 873 10967 887
rect 10993 833 11007 847
rect 10913 793 10927 807
rect 10813 713 10827 727
rect 10873 713 10887 727
rect 10913 693 10927 707
rect 10953 793 10967 807
rect 10933 653 10947 667
rect 10893 613 10907 627
rect 10973 773 10987 787
rect 10973 713 10987 727
rect 10813 593 10827 607
rect 10893 593 10907 607
rect 10953 593 10967 607
rect 10853 373 10867 387
rect 10793 333 10807 347
rect 10813 333 10827 347
rect 10813 173 10827 187
rect 10533 133 10547 147
rect 10553 133 10567 147
rect 10633 133 10647 147
rect 10673 133 10687 147
rect 10813 133 10827 147
rect 11073 1413 11087 1427
rect 11033 1313 11047 1327
rect 11013 713 11027 727
rect 11053 1273 11067 1287
rect 11253 1673 11267 1687
rect 11233 1593 11247 1607
rect 11253 1593 11267 1607
rect 11213 1573 11227 1587
rect 11353 2213 11367 2227
rect 11353 2193 11367 2207
rect 11333 2053 11347 2067
rect 11313 1773 11327 1787
rect 11353 2033 11367 2047
rect 11433 2593 11447 2607
rect 11413 2573 11427 2587
rect 11393 2533 11407 2547
rect 11413 2533 11427 2547
rect 11433 2513 11447 2527
rect 11413 2433 11427 2447
rect 11393 2153 11407 2167
rect 11393 2113 11407 2127
rect 11393 1853 11407 1867
rect 11373 1813 11387 1827
rect 11433 2413 11447 2427
rect 11513 4173 11527 4187
rect 11513 3493 11527 3507
rect 11613 4173 11627 4187
rect 11653 4173 11667 4187
rect 11553 4013 11567 4027
rect 11593 3993 11607 4007
rect 11633 3953 11647 3967
rect 11573 3793 11587 3807
rect 11553 3693 11567 3707
rect 11553 3493 11567 3507
rect 11533 3473 11547 3487
rect 11593 3713 11607 3727
rect 11793 6133 11807 6147
rect 11773 4393 11787 4407
rect 11773 4173 11787 4187
rect 11673 3973 11687 3987
rect 11733 3973 11747 3987
rect 11673 3893 11687 3907
rect 11653 3793 11667 3807
rect 11613 3693 11627 3707
rect 11753 3953 11767 3967
rect 11713 3933 11727 3947
rect 11653 3653 11667 3667
rect 11693 3653 11707 3667
rect 11673 3613 11687 3627
rect 11633 3593 11647 3607
rect 11593 3533 11607 3547
rect 11613 3493 11627 3507
rect 11633 3473 11647 3487
rect 11553 3213 11567 3227
rect 11573 3173 11587 3187
rect 11513 3133 11527 3147
rect 11513 3073 11527 3087
rect 11493 3033 11507 3047
rect 11493 3013 11507 3027
rect 11533 3013 11547 3027
rect 11493 2973 11507 2987
rect 11513 2913 11527 2927
rect 11593 2913 11607 2927
rect 11493 2673 11507 2687
rect 11553 2833 11567 2847
rect 11733 3573 11747 3587
rect 11713 3473 11727 3487
rect 11773 3933 11787 3947
rect 11813 5933 11827 5947
rect 11813 5693 11827 5707
rect 11813 5233 11827 5247
rect 11813 4913 11827 4927
rect 11813 4893 11827 4907
rect 11813 4693 11827 4707
rect 11813 4633 11827 4647
rect 11813 4173 11827 4187
rect 11813 3953 11827 3967
rect 11793 3713 11807 3727
rect 11773 3693 11787 3707
rect 11793 3613 11807 3627
rect 11813 3553 11827 3567
rect 11773 3533 11787 3547
rect 11753 3473 11767 3487
rect 11733 3453 11747 3467
rect 11753 3333 11767 3347
rect 11673 3313 11687 3327
rect 11653 3173 11667 3187
rect 11653 3153 11667 3167
rect 11713 3213 11727 3227
rect 11693 3193 11707 3207
rect 11713 3173 11727 3187
rect 11913 6873 11927 6887
rect 11973 6873 11987 6887
rect 11893 6433 11907 6447
rect 12113 6913 12127 6927
rect 12073 6813 12087 6827
rect 11993 6613 12007 6627
rect 12033 6613 12047 6627
rect 11993 6593 12007 6607
rect 11953 6573 11967 6587
rect 12133 6853 12147 6867
rect 12093 6593 12107 6607
rect 11933 6413 11947 6427
rect 11853 6393 11867 6407
rect 11873 6373 11887 6387
rect 11913 6373 11927 6387
rect 11853 6353 11867 6367
rect 11893 6353 11907 6367
rect 11933 6353 11947 6367
rect 11913 6333 11927 6347
rect 12093 6573 12107 6587
rect 12133 6573 12147 6587
rect 12013 6473 12027 6487
rect 12013 6393 12027 6407
rect 11973 6353 11987 6367
rect 11973 6133 11987 6147
rect 11853 6093 11867 6107
rect 11953 6113 11967 6127
rect 11913 6093 11927 6107
rect 11893 5973 11907 5987
rect 11933 5873 11947 5887
rect 11893 5713 11907 5727
rect 11873 5693 11887 5707
rect 11973 5693 11987 5707
rect 11853 5653 11867 5667
rect 12113 6393 12127 6407
rect 12173 6473 12187 6487
rect 12133 6373 12147 6387
rect 12033 6113 12047 6127
rect 12093 6133 12107 6147
rect 12073 6093 12087 6107
rect 12213 11673 12227 11687
rect 12053 5933 12067 5947
rect 12073 5933 12087 5947
rect 12033 5873 12047 5887
rect 12093 5873 12107 5887
rect 12013 5673 12027 5687
rect 11913 5653 11927 5667
rect 11933 5653 11947 5667
rect 11893 5453 11907 5467
rect 12073 5673 12087 5687
rect 12033 5653 12047 5667
rect 12093 5653 12107 5667
rect 12053 5633 12067 5647
rect 12013 5473 12027 5487
rect 12073 5473 12087 5487
rect 12053 5433 12067 5447
rect 11913 5413 11927 5427
rect 11953 5413 11967 5427
rect 12013 5413 12027 5427
rect 11873 5233 11887 5247
rect 12133 5433 12147 5447
rect 11913 5173 11927 5187
rect 11953 5173 11967 5187
rect 11913 5153 11927 5167
rect 12073 5153 12087 5167
rect 11893 5133 11907 5147
rect 11953 5133 11967 5147
rect 12053 5133 12067 5147
rect 11873 5033 11887 5047
rect 11913 5033 11927 5047
rect 11873 4973 11887 4987
rect 12013 4933 12027 4947
rect 12053 4933 12067 4947
rect 11893 4913 11907 4927
rect 11913 4913 11927 4927
rect 11853 4773 11867 4787
rect 11893 4753 11907 4767
rect 11873 4733 11887 4747
rect 11853 4693 11867 4707
rect 12033 4913 12047 4927
rect 12073 4893 12087 4907
rect 12013 4693 12027 4707
rect 12053 4693 12067 4707
rect 12113 4973 12127 4987
rect 12073 4673 12087 4687
rect 11913 4653 11927 4667
rect 11873 4633 11887 4647
rect 11853 4613 11867 4627
rect 11993 4473 12007 4487
rect 11893 4453 11907 4467
rect 11913 4413 11927 4427
rect 11973 4173 11987 4187
rect 11873 4153 11887 4167
rect 11793 3513 11807 3527
rect 11833 3513 11847 3527
rect 11753 3193 11767 3207
rect 11773 3193 11787 3207
rect 11733 3153 11747 3167
rect 11673 3033 11687 3047
rect 11713 3033 11727 3047
rect 11733 2993 11747 3007
rect 11773 3093 11787 3107
rect 11773 3053 11787 3067
rect 11693 2973 11707 2987
rect 11753 2973 11767 2987
rect 11693 2853 11707 2867
rect 11633 2793 11647 2807
rect 11533 2773 11547 2787
rect 11553 2773 11567 2787
rect 11553 2713 11567 2727
rect 11593 2713 11607 2727
rect 11633 2713 11647 2727
rect 11533 2693 11547 2707
rect 11513 2653 11527 2667
rect 11513 2573 11527 2587
rect 11533 2573 11547 2587
rect 11513 2533 11527 2547
rect 11593 2673 11607 2687
rect 11573 2653 11587 2667
rect 11473 2473 11487 2487
rect 11493 2313 11507 2327
rect 11553 2313 11567 2327
rect 11453 2293 11467 2307
rect 11453 2273 11467 2287
rect 11533 2293 11547 2307
rect 11433 2253 11447 2267
rect 11473 2253 11487 2267
rect 11513 2233 11527 2247
rect 11453 2213 11467 2227
rect 11513 2213 11527 2227
rect 11533 2213 11547 2227
rect 11433 2153 11447 2167
rect 11473 2193 11487 2207
rect 11453 1913 11467 1927
rect 11493 2093 11507 2107
rect 11433 1853 11447 1867
rect 11473 1853 11487 1867
rect 11413 1833 11427 1847
rect 11433 1813 11447 1827
rect 11473 1813 11487 1827
rect 11393 1773 11407 1787
rect 11333 1593 11347 1607
rect 11293 1573 11307 1587
rect 11293 1453 11307 1467
rect 11173 1313 11187 1327
rect 11153 1273 11167 1287
rect 11273 1353 11287 1367
rect 11213 1333 11227 1347
rect 11193 1233 11207 1247
rect 11113 1173 11127 1187
rect 11073 1133 11087 1147
rect 11113 1133 11127 1147
rect 11073 1113 11087 1127
rect 11093 1073 11107 1087
rect 11153 1073 11167 1087
rect 11133 1013 11147 1027
rect 11093 853 11107 867
rect 11153 853 11167 867
rect 11053 833 11067 847
rect 11053 673 11067 687
rect 10993 593 11007 607
rect 11073 653 11087 667
rect 11053 613 11067 627
rect 11193 813 11207 827
rect 11153 653 11167 667
rect 11093 613 11107 627
rect 11133 593 11147 607
rect 11033 433 11047 447
rect 11113 413 11127 427
rect 11093 393 11107 407
rect 10993 353 11007 367
rect 11033 353 11047 367
rect 11073 353 11087 367
rect 11153 393 11167 407
rect 11273 1293 11287 1307
rect 11253 1273 11267 1287
rect 11253 1113 11267 1127
rect 11373 1553 11387 1567
rect 11413 1553 11427 1567
rect 11373 1413 11387 1427
rect 11353 1333 11367 1347
rect 11313 1293 11327 1307
rect 11353 1273 11367 1287
rect 11413 1273 11427 1287
rect 11333 1233 11347 1247
rect 11453 1773 11467 1787
rect 11553 2193 11567 2207
rect 11553 2153 11567 2167
rect 11533 2093 11547 2107
rect 11613 2633 11627 2647
rect 11593 2233 11607 2247
rect 11573 2113 11587 2127
rect 11593 2093 11607 2107
rect 11573 2053 11587 2067
rect 11533 2033 11547 2047
rect 11553 1913 11567 1927
rect 11533 1853 11547 1867
rect 11513 1833 11527 1847
rect 11493 1553 11507 1567
rect 11473 1373 11487 1387
rect 11453 1213 11467 1227
rect 11433 1133 11447 1147
rect 11593 1753 11607 1767
rect 11593 1633 11607 1647
rect 11673 2653 11687 2667
rect 11673 2573 11687 2587
rect 11653 2493 11667 2507
rect 11733 2813 11747 2827
rect 11773 2813 11787 2827
rect 11713 2633 11727 2647
rect 11773 2793 11787 2807
rect 11833 3493 11847 3507
rect 11813 3473 11827 3487
rect 11853 3453 11867 3467
rect 11813 3293 11827 3307
rect 11893 3993 11907 4007
rect 11973 3993 11987 4007
rect 11893 3553 11907 3567
rect 11893 3493 11907 3507
rect 11893 3253 11907 3267
rect 11873 3193 11887 3207
rect 11833 3173 11847 3187
rect 11873 3173 11887 3187
rect 11893 3173 11907 3187
rect 12093 4473 12107 4487
rect 12073 4233 12087 4247
rect 12133 4233 12147 4247
rect 12013 4153 12027 4167
rect 12053 3993 12067 4007
rect 12093 3993 12107 4007
rect 12033 3873 12047 3887
rect 11933 3713 11947 3727
rect 11933 3253 11947 3267
rect 11933 3213 11947 3227
rect 11953 3133 11967 3147
rect 11913 3053 11927 3067
rect 11933 3053 11947 3067
rect 11913 3033 11927 3047
rect 11833 2993 11847 3007
rect 11853 2973 11867 2987
rect 11813 2853 11827 2867
rect 11813 2773 11827 2787
rect 11793 2753 11807 2767
rect 11833 2753 11847 2767
rect 11753 2713 11767 2727
rect 11793 2693 11807 2707
rect 11713 2553 11727 2567
rect 11733 2553 11747 2567
rect 11693 2313 11707 2327
rect 11633 2273 11647 2287
rect 11653 2273 11667 2287
rect 11653 2253 11667 2267
rect 11673 2253 11687 2267
rect 11713 2253 11727 2267
rect 11633 2193 11647 2207
rect 11633 2053 11647 2067
rect 11653 2013 11667 2027
rect 11753 2313 11767 2327
rect 11813 2653 11827 2667
rect 11813 2533 11827 2547
rect 11813 2333 11827 2347
rect 11793 2253 11807 2267
rect 11813 2253 11827 2267
rect 11753 2193 11767 2207
rect 11793 2173 11807 2187
rect 11753 2153 11767 2167
rect 11693 1893 11707 1907
rect 11653 1793 11667 1807
rect 11633 1773 11647 1787
rect 11693 1773 11707 1787
rect 11653 1633 11667 1647
rect 11673 1633 11687 1647
rect 11653 1613 11667 1627
rect 11553 1433 11567 1447
rect 11533 1373 11547 1387
rect 11513 1333 11527 1347
rect 11513 1313 11527 1327
rect 11613 1553 11627 1567
rect 11573 1313 11587 1327
rect 11593 1313 11607 1327
rect 11493 1193 11507 1207
rect 11413 1073 11427 1087
rect 11593 1273 11607 1287
rect 11533 1253 11547 1267
rect 11653 1553 11667 1567
rect 11693 1593 11707 1607
rect 11693 1573 11707 1587
rect 11673 1333 11687 1347
rect 11913 2873 11927 2887
rect 11893 2833 11907 2847
rect 11873 2773 11887 2787
rect 11853 2733 11867 2747
rect 11873 2713 11887 2727
rect 11853 2633 11867 2647
rect 11893 2633 11907 2647
rect 11893 2573 11907 2587
rect 11853 2553 11867 2567
rect 11993 3653 12007 3667
rect 12093 3693 12107 3707
rect 12153 3693 12167 3707
rect 12053 3533 12067 3547
rect 12033 3513 12047 3527
rect 12073 3513 12087 3527
rect 12013 3473 12027 3487
rect 12073 3293 12087 3307
rect 12173 3673 12187 3687
rect 12193 3673 12207 3687
rect 12093 3273 12107 3287
rect 12013 3253 12027 3267
rect 12053 3253 12067 3267
rect 11933 2733 11947 2747
rect 11953 2713 11967 2727
rect 11873 2533 11887 2547
rect 11933 2493 11947 2507
rect 11973 2493 11987 2507
rect 11953 2293 11967 2307
rect 11853 2273 11867 2287
rect 11893 2273 11907 2287
rect 11873 2253 11887 2267
rect 11913 2233 11927 2247
rect 11933 2133 11947 2147
rect 11893 2113 11907 2127
rect 11873 2093 11887 2107
rect 11833 1833 11847 1847
rect 11733 1773 11747 1787
rect 11793 1793 11807 1807
rect 11773 1773 11787 1787
rect 11753 1753 11767 1767
rect 11813 1753 11827 1767
rect 11833 1693 11847 1707
rect 11753 1633 11767 1647
rect 11793 1593 11807 1607
rect 11773 1573 11787 1587
rect 11813 1573 11827 1587
rect 11733 1553 11747 1567
rect 11793 1373 11807 1387
rect 11653 1313 11667 1327
rect 11633 1253 11647 1267
rect 11613 1233 11627 1247
rect 11573 1193 11587 1207
rect 11513 1093 11527 1107
rect 11453 1033 11467 1047
rect 11333 933 11347 947
rect 11473 933 11487 947
rect 11453 833 11467 847
rect 11353 733 11367 747
rect 11393 733 11407 747
rect 11253 653 11267 667
rect 11353 653 11367 667
rect 11313 613 11327 627
rect 11333 593 11347 607
rect 11293 573 11307 587
rect 11293 393 11307 407
rect 11253 373 11267 387
rect 11113 353 11127 367
rect 11133 353 11147 367
rect 11213 353 11227 367
rect 11013 333 11027 347
rect 11053 333 11067 347
rect 11093 333 11107 347
rect 10993 313 11007 327
rect 10973 273 10987 287
rect 11053 273 11067 287
rect 10873 213 10887 227
rect 10913 213 10927 227
rect 10873 153 10887 167
rect 10893 133 10907 147
rect 11073 153 11087 167
rect 11093 133 11107 147
rect 11273 313 11287 327
rect 11233 293 11247 307
rect 11213 193 11227 207
rect 11373 633 11387 647
rect 11373 593 11387 607
rect 11353 573 11367 587
rect 11373 573 11387 587
rect 11473 713 11487 727
rect 11533 713 11547 727
rect 11493 673 11507 687
rect 11533 653 11547 667
rect 11453 573 11467 587
rect 11513 573 11527 587
rect 11433 373 11447 387
rect 11473 353 11487 367
rect 11633 1113 11647 1127
rect 11613 1093 11627 1107
rect 11673 1293 11687 1307
rect 11693 1273 11707 1287
rect 11713 1253 11727 1267
rect 11673 1113 11687 1127
rect 11753 1333 11767 1347
rect 11653 1093 11667 1107
rect 11673 1093 11687 1107
rect 11653 1073 11667 1087
rect 11693 1073 11707 1087
rect 11733 1093 11747 1107
rect 11773 1213 11787 1227
rect 11753 1073 11767 1087
rect 11733 1033 11747 1047
rect 11793 1073 11807 1087
rect 11793 1053 11807 1067
rect 11773 873 11787 887
rect 11713 833 11727 847
rect 11673 813 11687 827
rect 11693 813 11707 827
rect 11653 713 11667 727
rect 11613 613 11627 627
rect 11633 613 11647 627
rect 11613 593 11627 607
rect 11633 573 11647 587
rect 11773 853 11787 867
rect 11753 653 11767 667
rect 11733 633 11747 647
rect 11693 613 11707 627
rect 11673 593 11687 607
rect 11713 593 11727 607
rect 11753 593 11767 607
rect 11713 373 11727 387
rect 11633 353 11647 367
rect 11673 353 11687 367
rect 11373 313 11387 327
rect 11573 333 11587 347
rect 11633 333 11647 347
rect 11653 333 11667 347
rect 11793 333 11807 347
rect 11273 173 11287 187
rect 11333 173 11347 187
rect 11233 153 11247 167
rect 11333 153 11347 167
rect 11473 193 11487 207
rect 11493 193 11507 207
rect 11873 1413 11887 1427
rect 11913 2073 11927 2087
rect 11953 2093 11967 2107
rect 11973 2093 11987 2107
rect 12053 3213 12067 3227
rect 12033 3193 12047 3207
rect 12113 3213 12127 3227
rect 12073 3053 12087 3067
rect 12133 2993 12147 3007
rect 12053 2793 12067 2807
rect 12073 2793 12087 2807
rect 12053 2393 12067 2407
rect 12033 2293 12047 2307
rect 12093 2553 12107 2567
rect 12073 2293 12087 2307
rect 12093 2273 12107 2287
rect 12073 2253 12087 2267
rect 12033 2213 12047 2227
rect 12013 2113 12027 2127
rect 12013 2093 12027 2107
rect 11993 2073 12007 2087
rect 11893 1393 11907 1407
rect 11993 2053 12007 2067
rect 11953 2033 11967 2047
rect 11933 1833 11947 1847
rect 12093 2053 12107 2067
rect 12053 2013 12067 2027
rect 11933 1613 11947 1627
rect 11973 1613 11987 1627
rect 12033 1733 12047 1747
rect 12153 2733 12167 2747
rect 12213 2033 12227 2047
rect 12113 1713 12127 1727
rect 12073 1693 12087 1707
rect 12033 1613 12047 1627
rect 11993 1593 12007 1607
rect 11953 1573 11967 1587
rect 11973 1413 11987 1427
rect 11913 1353 11927 1367
rect 11953 1353 11967 1367
rect 11853 1313 11867 1327
rect 11833 1233 11847 1247
rect 11913 1333 11927 1347
rect 11893 1273 11907 1287
rect 11873 1213 11887 1227
rect 11933 1213 11947 1227
rect 11873 1173 11887 1187
rect 11853 1073 11867 1087
rect 11893 1073 11907 1087
rect 12033 1553 12047 1567
rect 12033 1393 12047 1407
rect 12013 1273 12027 1287
rect 11993 1233 12007 1247
rect 11973 1213 11987 1227
rect 11973 1133 11987 1147
rect 11973 1113 11987 1127
rect 11953 1073 11967 1087
rect 11933 893 11947 907
rect 11933 873 11947 887
rect 11873 853 11887 867
rect 11893 813 11907 827
rect 11853 713 11867 727
rect 11913 713 11927 727
rect 11853 693 11867 707
rect 11893 633 11907 647
rect 12053 1373 12067 1387
rect 12093 1313 12107 1327
rect 12113 1273 12127 1287
rect 12073 1233 12087 1247
rect 12013 1113 12027 1127
rect 11993 1093 12007 1107
rect 12033 1093 12047 1107
rect 12033 873 12047 887
rect 12093 813 12107 827
rect 12053 753 12067 767
rect 12073 753 12087 767
rect 11973 633 11987 647
rect 11873 593 11887 607
rect 11953 593 11967 607
rect 12033 593 12047 607
rect 11833 373 11847 387
rect 12013 393 12027 407
rect 12053 373 12067 387
rect 12033 353 12047 367
rect 11853 333 11867 347
rect 11953 333 11967 347
rect 12033 333 12047 347
rect 12073 333 12087 347
rect 11813 233 11827 247
rect 11833 233 11847 247
rect 11793 193 11807 207
rect 11813 173 11827 187
rect 11853 153 11867 167
rect 11213 133 11227 147
rect 11293 133 11307 147
rect 11453 133 11467 147
rect 11493 133 11507 147
rect 11653 133 11667 147
rect 8053 113 8067 127
rect 8273 113 8287 127
rect 8393 113 8407 127
rect 9293 113 9307 127
rect 9373 113 9387 127
rect 10293 113 10307 127
rect 11133 113 11147 127
rect 11253 113 11267 127
rect 8013 93 8027 107
rect 12033 153 12047 167
<< metal3 >>
rect 507 12016 1213 12024
rect 1227 12016 5993 12024
rect 6007 12016 6213 12024
rect 1527 11936 1673 11944
rect 1687 11936 5793 11944
rect 207 11916 733 11924
rect 747 11916 873 11924
rect 2267 11916 2613 11924
rect 2627 11916 2933 11924
rect 2947 11916 3813 11924
rect 4767 11916 5133 11924
rect 5147 11916 5773 11924
rect 6107 11916 6833 11924
rect 7587 11916 8233 11924
rect 8247 11916 8833 11924
rect 10567 11916 10613 11924
rect 11307 11916 12073 11924
rect 307 11896 513 11904
rect 567 11896 793 11904
rect 807 11896 1053 11904
rect 2047 11896 2424 11904
rect 2416 11887 2424 11896
rect 2447 11896 2553 11904
rect 2927 11896 2973 11904
rect 3707 11896 3773 11904
rect 3827 11896 4133 11904
rect 4156 11896 4893 11904
rect 4156 11887 4164 11896
rect 4907 11896 4973 11904
rect 5467 11896 6013 11904
rect 6807 11896 6913 11904
rect 7147 11896 7653 11904
rect 8147 11896 8253 11904
rect 8647 11896 8693 11904
rect 9247 11896 9433 11904
rect 10607 11896 10893 11904
rect 10907 11896 11153 11904
rect 11707 11896 11993 11904
rect 167 11876 253 11884
rect 547 11876 693 11884
rect 1087 11876 1153 11884
rect 1267 11876 1393 11884
rect 1827 11876 2024 11884
rect 2016 11867 2024 11876
rect 4176 11876 4493 11884
rect 107 11856 133 11864
rect 367 11856 893 11864
rect 907 11856 953 11864
rect 1427 11856 1613 11864
rect 2216 11864 2224 11873
rect 2216 11856 3153 11864
rect 3307 11856 3793 11864
rect 4176 11864 4184 11876
rect 4547 11876 4573 11884
rect 4947 11876 5113 11884
rect 5247 11876 5313 11884
rect 6367 11876 6753 11884
rect 6887 11876 7013 11884
rect 7027 11876 7093 11884
rect 7107 11876 7313 11884
rect 7367 11876 7453 11884
rect 7927 11876 7953 11884
rect 8247 11876 8273 11884
rect 8327 11876 8453 11884
rect 8687 11876 9393 11884
rect 9976 11884 9984 11893
rect 9547 11876 10653 11884
rect 11067 11876 11093 11884
rect 11407 11876 11753 11884
rect 3807 11856 4184 11864
rect 4327 11856 4393 11864
rect 4567 11856 4693 11864
rect 4747 11856 4913 11864
rect 5347 11856 5473 11864
rect 6536 11856 7073 11864
rect 6536 11847 6544 11856
rect 7127 11856 7493 11864
rect 7507 11856 7693 11864
rect 8087 11856 8864 11864
rect 267 11836 333 11844
rect 767 11836 793 11844
rect 1247 11836 1273 11844
rect 1647 11836 1833 11844
rect 2767 11836 2953 11844
rect 4207 11836 4333 11844
rect 4347 11836 5073 11844
rect 5307 11836 5313 11844
rect 5327 11836 5453 11844
rect 6067 11836 6093 11844
rect 6947 11836 7153 11844
rect 7167 11836 7373 11844
rect 7727 11836 8833 11844
rect 8856 11844 8864 11856
rect 8887 11856 8933 11864
rect 9067 11856 9233 11864
rect 9467 11856 10893 11864
rect 11467 11856 11913 11864
rect 11927 11856 11973 11864
rect 8856 11836 8993 11844
rect 9047 11836 9193 11844
rect 9427 11836 9653 11844
rect 10327 11836 10853 11844
rect 10927 11836 11073 11844
rect 11387 11836 11433 11844
rect 11587 11836 11633 11844
rect 187 11816 353 11824
rect 787 11816 933 11824
rect 947 11816 1113 11824
rect 1487 11816 1973 11824
rect 1987 11816 2193 11824
rect 2387 11816 3613 11824
rect 3627 11816 4753 11824
rect 5127 11816 5253 11824
rect 5267 11816 6513 11824
rect 6527 11816 6673 11824
rect 6727 11816 7053 11824
rect 7347 11816 7713 11824
rect 8107 11816 8593 11824
rect 8927 11816 9873 11824
rect 10727 11816 12193 11824
rect 2347 11796 3113 11804
rect 3127 11796 4513 11804
rect 4527 11796 4553 11804
rect 4587 11796 4873 11804
rect 4887 11796 5233 11804
rect 5247 11796 5893 11804
rect 5907 11796 5973 11804
rect 5987 11796 6073 11804
rect 6087 11796 6553 11804
rect 6567 11796 7893 11804
rect 8827 11796 9173 11804
rect 9187 11796 10533 11804
rect 10587 11796 10833 11804
rect 11207 11796 12093 11804
rect 1267 11776 2053 11784
rect 2067 11776 3493 11784
rect 4007 11776 4133 11784
rect 4147 11776 4493 11784
rect 4987 11776 5513 11784
rect 5527 11776 5713 11784
rect 5727 11776 5853 11784
rect 5887 11776 7293 11784
rect 7387 11776 8133 11784
rect 8327 11776 9313 11784
rect 9427 11776 9833 11784
rect 9847 11776 10313 11784
rect 10387 11776 11344 11784
rect 2567 11756 2613 11764
rect 2627 11756 2873 11764
rect 3467 11756 3573 11764
rect 3767 11756 4593 11764
rect 4727 11756 4873 11764
rect 5087 11756 6313 11764
rect 6907 11756 7513 11764
rect 7947 11756 8093 11764
rect 8107 11756 9333 11764
rect 9407 11756 9533 11764
rect 9647 11756 10693 11764
rect 11336 11764 11344 11776
rect 11367 11776 11613 11784
rect 11336 11756 11473 11764
rect 11827 11756 11993 11764
rect 2807 11736 2993 11744
rect 3007 11736 3253 11744
rect 3267 11736 5433 11744
rect 5707 11736 8353 11744
rect 8507 11736 8713 11744
rect 9047 11736 11053 11744
rect 11287 11736 12013 11744
rect 727 11716 1593 11724
rect 1707 11716 2133 11724
rect 2147 11716 3073 11724
rect 3087 11716 3193 11724
rect 3207 11716 4293 11724
rect 4987 11716 6733 11724
rect 7767 11716 8533 11724
rect 8707 11716 10933 11724
rect 11347 11716 11713 11724
rect 647 11696 913 11704
rect 1347 11696 1953 11704
rect 1967 11696 2173 11704
rect 2707 11696 2773 11704
rect 2787 11696 2833 11704
rect 3427 11696 3453 11704
rect 4307 11696 4433 11704
rect 4907 11696 5413 11704
rect 5447 11696 6393 11704
rect 6447 11696 6613 11704
rect 6767 11696 7473 11704
rect 7587 11696 7693 11704
rect 7887 11696 8053 11704
rect 8147 11696 8213 11704
rect 8247 11696 8273 11704
rect 8307 11696 8433 11704
rect 8607 11696 8653 11704
rect 9227 11696 10013 11704
rect 10027 11696 10133 11704
rect 11047 11696 12153 11704
rect 227 11676 313 11684
rect 496 11676 673 11684
rect 136 11664 144 11673
rect 136 11656 153 11664
rect 167 11656 373 11664
rect 496 11664 504 11676
rect 807 11676 1093 11684
rect 1147 11676 1273 11684
rect 1927 11676 2273 11684
rect 2667 11676 2713 11684
rect 3327 11676 3433 11684
rect 3896 11676 3973 11684
rect 387 11656 504 11664
rect 907 11656 933 11664
rect 987 11656 1073 11664
rect 1087 11656 1113 11664
rect 1547 11656 1593 11664
rect 1607 11656 2013 11664
rect 1287 11636 1313 11644
rect 1496 11644 1504 11653
rect 1716 11647 1724 11656
rect 2287 11656 2313 11664
rect 2456 11664 2464 11673
rect 2456 11656 2633 11664
rect 2867 11656 2933 11664
rect 2967 11656 3033 11664
rect 3247 11656 3313 11664
rect 3647 11656 3733 11664
rect 3896 11664 3904 11676
rect 4027 11676 4073 11684
rect 4087 11676 4113 11684
rect 4347 11676 4373 11684
rect 4547 11676 4673 11684
rect 4747 11676 4913 11684
rect 4967 11676 5113 11684
rect 5127 11676 5653 11684
rect 3787 11656 3904 11664
rect 3927 11656 3953 11664
rect 3967 11656 4293 11664
rect 4367 11656 4613 11664
rect 5287 11656 5333 11664
rect 5376 11664 5384 11676
rect 5947 11676 6033 11684
rect 6087 11676 6213 11684
rect 6247 11676 6413 11684
rect 6436 11676 6684 11684
rect 5376 11656 5493 11664
rect 5516 11656 5553 11664
rect 1367 11636 1673 11644
rect 2087 11636 2153 11644
rect 2607 11636 2693 11644
rect 3067 11636 3253 11644
rect 3447 11636 3873 11644
rect 3887 11636 4353 11644
rect 4387 11636 4513 11644
rect 5516 11644 5524 11656
rect 5607 11656 5693 11664
rect 5887 11656 6233 11664
rect 6436 11664 6444 11676
rect 6287 11656 6444 11664
rect 6507 11656 6653 11664
rect 6676 11664 6684 11676
rect 6727 11676 6813 11684
rect 6867 11676 6893 11684
rect 7967 11676 8473 11684
rect 8527 11676 8573 11684
rect 9027 11676 9173 11684
rect 9187 11676 9793 11684
rect 9847 11676 9873 11684
rect 9887 11676 9993 11684
rect 10047 11676 10273 11684
rect 10307 11676 10673 11684
rect 10947 11676 11053 11684
rect 11127 11676 11293 11684
rect 11507 11676 11533 11684
rect 12147 11676 12213 11684
rect 6676 11656 7064 11664
rect 4536 11636 5524 11644
rect 5536 11636 5673 11644
rect 2187 11616 2253 11624
rect 2267 11616 2673 11624
rect 2687 11616 3433 11624
rect 4536 11624 4544 11636
rect 3487 11616 4544 11624
rect 4947 11616 4973 11624
rect 5536 11624 5544 11636
rect 5687 11636 5933 11644
rect 6307 11636 6453 11644
rect 6567 11636 6633 11644
rect 6707 11636 7033 11644
rect 7056 11644 7064 11656
rect 7127 11656 7173 11664
rect 8287 11656 8873 11664
rect 8887 11656 9073 11664
rect 9127 11656 9273 11664
rect 9287 11656 9433 11664
rect 9487 11656 9673 11664
rect 9707 11656 10333 11664
rect 10367 11656 10393 11664
rect 10407 11656 10493 11664
rect 10736 11664 10744 11673
rect 10736 11656 11253 11664
rect 11907 11656 12173 11664
rect 7056 11636 8253 11644
rect 8607 11636 8653 11644
rect 8827 11636 8853 11644
rect 9007 11636 9053 11644
rect 9107 11636 9153 11644
rect 9307 11636 9324 11644
rect 9316 11627 9324 11636
rect 9347 11636 9453 11644
rect 10127 11636 10153 11644
rect 10287 11636 10313 11644
rect 10467 11636 10513 11644
rect 10536 11636 11273 11644
rect 5107 11616 5544 11624
rect 5567 11616 5893 11624
rect 5947 11616 6573 11624
rect 6687 11616 6713 11624
rect 6747 11616 6833 11624
rect 7007 11616 8073 11624
rect 8087 11616 8233 11624
rect 9347 11616 9493 11624
rect 10536 11624 10544 11636
rect 9867 11616 10544 11624
rect 10627 11616 10713 11624
rect 10887 11616 11093 11624
rect 11427 11616 11593 11624
rect 1867 11596 2193 11604
rect 2207 11596 2393 11604
rect 2407 11596 2653 11604
rect 4267 11596 4573 11604
rect 4607 11596 5624 11604
rect 1927 11576 3253 11584
rect 3267 11576 3593 11584
rect 3607 11576 4313 11584
rect 5347 11576 5593 11584
rect 5616 11584 5624 11596
rect 5727 11596 6293 11604
rect 6907 11596 8633 11604
rect 8727 11596 9693 11604
rect 10667 11596 11173 11604
rect 11187 11596 11553 11604
rect 5616 11576 5853 11584
rect 5907 11576 6693 11584
rect 8947 11576 10293 11584
rect 10427 11576 10533 11584
rect 10747 11576 11393 11584
rect 11467 11576 11933 11584
rect 3627 11556 3813 11564
rect 3827 11556 4173 11564
rect 4196 11556 4413 11564
rect 2307 11536 2913 11544
rect 3047 11536 3533 11544
rect 3607 11536 3913 11544
rect 3947 11536 3953 11544
rect 4196 11544 4204 11556
rect 4427 11556 4473 11564
rect 4547 11556 4713 11564
rect 4727 11556 6773 11564
rect 9447 11556 10413 11564
rect 11667 11556 11693 11564
rect 11747 11556 11973 11564
rect 3967 11536 4204 11544
rect 4287 11536 6553 11544
rect 7527 11536 11813 11544
rect 3467 11516 4284 11524
rect 2507 11496 3373 11504
rect 3387 11496 3993 11504
rect 4007 11496 4253 11504
rect 4276 11504 4284 11516
rect 4307 11516 8513 11524
rect 8547 11516 9793 11524
rect 11247 11516 12153 11524
rect 4276 11496 4353 11504
rect 4587 11496 5293 11504
rect 5307 11496 5433 11504
rect 5467 11496 5713 11504
rect 8467 11496 11073 11504
rect 11087 11496 11433 11504
rect 11567 11496 12113 11504
rect 2007 11476 2753 11484
rect 3027 11476 3053 11484
rect 3547 11476 3644 11484
rect 2127 11456 2393 11464
rect 2407 11456 2513 11464
rect 2527 11456 3553 11464
rect 3636 11464 3644 11476
rect 3667 11476 3773 11484
rect 4367 11476 6053 11484
rect 7087 11476 7864 11484
rect 3636 11456 4093 11464
rect 4347 11456 4553 11464
rect 4567 11456 5633 11464
rect 5647 11456 7833 11464
rect 7856 11464 7864 11476
rect 8307 11476 9073 11484
rect 9327 11476 9933 11484
rect 9947 11476 10453 11484
rect 11867 11476 11993 11484
rect 7856 11456 10653 11464
rect 11787 11456 11913 11464
rect 1007 11436 1473 11444
rect 1887 11436 2073 11444
rect 2447 11436 2573 11444
rect 2647 11436 3153 11444
rect 3167 11436 4113 11444
rect 4127 11436 4733 11444
rect 4747 11436 6113 11444
rect 6127 11436 7313 11444
rect 7507 11436 8113 11444
rect 8587 11436 9713 11444
rect 10267 11436 11013 11444
rect 11107 11436 11513 11444
rect 11587 11436 11633 11444
rect 227 11416 633 11424
rect 647 11416 753 11424
rect 1467 11416 1513 11424
rect 1527 11416 1873 11424
rect 1987 11416 2033 11424
rect 2056 11416 2433 11424
rect 2056 11407 2064 11416
rect 2487 11416 2833 11424
rect 2847 11416 2953 11424
rect 2967 11416 3333 11424
rect 3567 11416 3833 11424
rect 4247 11416 4313 11424
rect 4327 11416 4813 11424
rect 5507 11416 5573 11424
rect 5647 11416 5733 11424
rect 5807 11416 5913 11424
rect 5927 11416 6073 11424
rect 7087 11416 7213 11424
rect 7227 11416 7393 11424
rect 7407 11416 7573 11424
rect 7847 11416 7913 11424
rect 7967 11416 8033 11424
rect 8247 11416 8313 11424
rect 8927 11416 9013 11424
rect 9067 11416 9153 11424
rect 9167 11416 9313 11424
rect 9387 11416 9473 11424
rect 9496 11416 9864 11424
rect 407 11396 424 11404
rect 107 11376 373 11384
rect 416 11384 424 11396
rect 447 11396 833 11404
rect 847 11396 933 11404
rect 1167 11396 1364 11404
rect 416 11376 604 11384
rect 596 11367 604 11376
rect 827 11376 913 11384
rect 967 11376 993 11384
rect 1207 11376 1313 11384
rect 1327 11376 1333 11384
rect 1356 11384 1364 11396
rect 2427 11396 2573 11404
rect 2627 11396 2693 11404
rect 2807 11396 2924 11404
rect 1356 11376 1653 11384
rect 1667 11376 1864 11384
rect 367 11356 413 11364
rect 427 11356 573 11364
rect 787 11356 973 11364
rect 1127 11356 1573 11364
rect 1587 11356 1833 11364
rect 1856 11364 1864 11376
rect 2147 11376 2253 11384
rect 2327 11376 2413 11384
rect 2427 11376 2553 11384
rect 2607 11376 2733 11384
rect 2916 11384 2924 11396
rect 2947 11396 2973 11404
rect 3067 11396 3213 11404
rect 3327 11396 3764 11404
rect 3756 11387 3764 11396
rect 3887 11396 4493 11404
rect 5147 11396 5893 11404
rect 5947 11396 5973 11404
rect 6207 11396 6293 11404
rect 6436 11396 6613 11404
rect 2916 11376 2993 11384
rect 3167 11376 3213 11384
rect 3507 11376 3713 11384
rect 3767 11376 3893 11384
rect 4247 11376 4273 11384
rect 4447 11376 4873 11384
rect 4887 11376 5053 11384
rect 5067 11376 5193 11384
rect 5587 11376 5633 11384
rect 5727 11376 5753 11384
rect 6067 11376 6293 11384
rect 6436 11384 6444 11396
rect 6667 11396 6953 11404
rect 7107 11396 7133 11404
rect 7387 11396 7533 11404
rect 7587 11396 7673 11404
rect 7687 11396 7893 11404
rect 7927 11396 7933 11404
rect 7947 11396 8133 11404
rect 8187 11396 8293 11404
rect 8567 11396 8893 11404
rect 9496 11404 9504 11416
rect 9307 11396 9504 11404
rect 9856 11404 9864 11416
rect 10027 11416 10393 11424
rect 10467 11416 10573 11424
rect 10627 11416 10813 11424
rect 10827 11416 10893 11424
rect 11007 11416 11324 11424
rect 11316 11407 11324 11416
rect 11547 11416 11564 11424
rect 9856 11396 10064 11404
rect 6307 11376 6444 11384
rect 6647 11376 6733 11384
rect 6787 11376 6813 11384
rect 6987 11376 7153 11384
rect 7287 11376 7553 11384
rect 7607 11376 7713 11384
rect 7747 11376 7833 11384
rect 7856 11376 8113 11384
rect 1856 11356 2393 11364
rect 2687 11356 3113 11364
rect 3387 11356 3733 11364
rect 3747 11356 3953 11364
rect 4187 11356 4473 11364
rect 4707 11356 4753 11364
rect 5047 11356 5093 11364
rect 5427 11356 5593 11364
rect 6456 11364 6464 11373
rect 5767 11356 6464 11364
rect 6847 11356 6913 11364
rect 6967 11356 7753 11364
rect 7856 11364 7864 11376
rect 8167 11376 9093 11384
rect 9107 11376 9253 11384
rect 9267 11376 9373 11384
rect 9507 11376 9633 11384
rect 9707 11376 9853 11384
rect 9887 11376 10033 11384
rect 10056 11384 10064 11396
rect 10607 11396 10653 11404
rect 10927 11396 10953 11404
rect 11147 11396 11293 11404
rect 10056 11376 10213 11384
rect 10807 11376 10933 11384
rect 10987 11376 11013 11384
rect 11336 11384 11344 11413
rect 11556 11404 11564 11416
rect 11587 11416 11673 11424
rect 11727 11416 11793 11424
rect 11847 11416 11873 11424
rect 12107 11416 12133 11424
rect 11556 11396 11693 11404
rect 11827 11396 11893 11404
rect 11327 11376 11344 11384
rect 11807 11376 11933 11384
rect 11947 11376 12033 11384
rect 7767 11356 7864 11364
rect 7947 11356 9193 11364
rect 9607 11356 10073 11364
rect 10567 11356 11873 11364
rect 11927 11356 12113 11364
rect 1367 11336 1533 11344
rect 1547 11336 1593 11344
rect 1627 11336 1693 11344
rect 1707 11336 2793 11344
rect 2927 11336 3153 11344
rect 3356 11344 3364 11353
rect 3247 11336 3873 11344
rect 3887 11336 3913 11344
rect 3947 11336 4793 11344
rect 4807 11336 4953 11344
rect 4967 11336 5233 11344
rect 5247 11336 5253 11344
rect 5267 11336 5373 11344
rect 5747 11336 6133 11344
rect 6487 11336 6793 11344
rect 8347 11336 9484 11344
rect 1567 11316 1833 11324
rect 1847 11316 2213 11324
rect 2247 11316 2273 11324
rect 2667 11316 3933 11324
rect 3956 11316 5013 11324
rect 2107 11296 2673 11304
rect 2727 11296 2993 11304
rect 3147 11296 3393 11304
rect 3956 11304 3964 11316
rect 5407 11316 7333 11324
rect 7987 11316 8193 11324
rect 8447 11316 8733 11324
rect 8767 11316 9453 11324
rect 9476 11324 9484 11336
rect 9647 11336 11193 11344
rect 11667 11336 11833 11344
rect 9476 11316 10453 11324
rect 11547 11316 12053 11324
rect 3447 11296 3964 11304
rect 4187 11296 4293 11304
rect 4867 11296 7913 11304
rect 8207 11296 8853 11304
rect 9007 11296 9593 11304
rect 9747 11296 9833 11304
rect 10027 11296 11033 11304
rect 11287 11296 11613 11304
rect 1527 11276 2113 11284
rect 2247 11276 2673 11284
rect 2687 11276 3133 11284
rect 3747 11276 4073 11284
rect 4087 11276 4133 11284
rect 4167 11276 6093 11284
rect 6187 11276 6653 11284
rect 7787 11276 8253 11284
rect 8267 11276 8313 11284
rect 8327 11276 8493 11284
rect 9127 11276 10653 11284
rect 10867 11276 11133 11284
rect 1907 11256 2373 11264
rect 2407 11256 3433 11264
rect 3647 11256 4313 11264
rect 5027 11256 5733 11264
rect 6167 11256 7353 11264
rect 8047 11256 8553 11264
rect 8607 11256 8713 11264
rect 8827 11256 11473 11264
rect 12067 11256 12173 11264
rect 947 11236 2153 11244
rect 2527 11236 2553 11244
rect 2807 11236 3153 11244
rect 3167 11236 3733 11244
rect 4507 11236 4653 11244
rect 4667 11236 5493 11244
rect 6447 11236 7893 11244
rect 8367 11236 9913 11244
rect 11467 11236 11513 11244
rect 11647 11236 11693 11244
rect 167 11216 373 11224
rect 1327 11216 1353 11224
rect 1547 11216 1693 11224
rect 2347 11216 2573 11224
rect 2887 11216 3053 11224
rect 3067 11216 3713 11224
rect 3727 11216 3753 11224
rect 4087 11216 4153 11224
rect 4827 11216 4993 11224
rect 5227 11216 5333 11224
rect 5447 11216 5693 11224
rect 5727 11216 5753 11224
rect 6587 11216 7013 11224
rect 7567 11216 8113 11224
rect 8407 11216 8453 11224
rect 8567 11216 8713 11224
rect 9207 11216 9553 11224
rect 9607 11216 9953 11224
rect 10067 11216 10833 11224
rect 11147 11216 12053 11224
rect 147 11196 233 11204
rect 767 11196 1113 11204
rect 1247 11196 1293 11204
rect 1347 11196 1473 11204
rect 1707 11196 1753 11204
rect 1787 11196 2113 11204
rect 2267 11196 2293 11204
rect 2527 11196 2604 11204
rect 356 11184 364 11193
rect 227 11176 564 11184
rect 556 11167 564 11176
rect 587 11176 733 11184
rect 1167 11176 1253 11184
rect 1287 11176 1313 11184
rect 1667 11176 1713 11184
rect 1727 11176 1913 11184
rect 1936 11176 2073 11184
rect 1936 11167 1944 11176
rect 2167 11176 2433 11184
rect 2447 11176 2493 11184
rect 2547 11176 2573 11184
rect 2596 11184 2604 11196
rect 2847 11196 2913 11204
rect 3327 11196 3433 11204
rect 3527 11196 3633 11204
rect 3707 11196 3913 11204
rect 4307 11196 4353 11204
rect 4387 11196 4393 11204
rect 4407 11196 4833 11204
rect 4847 11196 4933 11204
rect 5047 11196 5053 11204
rect 5067 11196 5193 11204
rect 5207 11196 5473 11204
rect 5487 11196 5513 11204
rect 5547 11196 5893 11204
rect 5947 11196 6013 11204
rect 6347 11196 6993 11204
rect 7067 11196 7204 11204
rect 2596 11176 2893 11184
rect 3707 11176 3864 11184
rect 967 11156 1093 11164
rect 1107 11156 1133 11164
rect 1747 11156 1773 11164
rect 2147 11156 2313 11164
rect 2367 11156 3193 11164
rect 3587 11156 3673 11164
rect 3856 11164 3864 11176
rect 3887 11176 4133 11184
rect 4187 11176 4233 11184
rect 4287 11176 4333 11184
rect 4407 11176 4453 11184
rect 5007 11176 5073 11184
rect 5507 11176 5553 11184
rect 5927 11176 6113 11184
rect 6136 11184 6144 11193
rect 7196 11187 7204 11196
rect 7327 11196 7533 11204
rect 8167 11196 8564 11204
rect 6136 11176 6313 11184
rect 7047 11176 7073 11184
rect 7367 11176 8333 11184
rect 8556 11184 8564 11196
rect 8787 11196 8953 11204
rect 8967 11196 9313 11204
rect 9387 11196 9433 11204
rect 9927 11196 10193 11204
rect 10327 11196 10513 11204
rect 10547 11196 10633 11204
rect 10867 11196 11004 11204
rect 10996 11187 11004 11196
rect 11316 11196 11333 11204
rect 11316 11187 11324 11196
rect 11547 11196 11613 11204
rect 8527 11176 8544 11184
rect 8556 11176 9533 11184
rect 3856 11156 5213 11164
rect 5367 11156 5913 11164
rect 6356 11164 6364 11173
rect 5967 11156 6364 11164
rect 6807 11156 6833 11164
rect 6847 11156 7153 11164
rect 7707 11156 7913 11164
rect 8536 11164 8544 11176
rect 8536 11156 8693 11164
rect 8707 11156 8753 11164
rect 8847 11156 8933 11164
rect 9336 11164 9344 11176
rect 9567 11176 10084 11184
rect 9167 11156 9344 11164
rect 9367 11156 10053 11164
rect 10076 11164 10084 11176
rect 10107 11176 10133 11184
rect 10487 11176 10573 11184
rect 11347 11176 11433 11184
rect 10076 11156 10113 11164
rect 10507 11156 10513 11164
rect 10527 11156 11113 11164
rect 11187 11156 11453 11164
rect 1027 11136 1173 11144
rect 1187 11136 1273 11144
rect 1287 11136 1853 11144
rect 2727 11136 3073 11144
rect 3087 11136 3273 11144
rect 3407 11136 3893 11144
rect 4447 11136 4673 11144
rect 6367 11136 6413 11144
rect 6567 11136 8193 11144
rect 10907 11136 11633 11144
rect 12027 11136 12053 11144
rect 2107 11116 2253 11124
rect 2327 11116 2413 11124
rect 3147 11116 3193 11124
rect 3207 11116 3673 11124
rect 3907 11116 5133 11124
rect 5187 11116 5533 11124
rect 5767 11116 7373 11124
rect 7387 11116 8093 11124
rect 8947 11116 9653 11124
rect 10147 11116 11533 11124
rect 1627 11096 2313 11104
rect 3187 11096 3613 11104
rect 3667 11096 5173 11104
rect 6027 11096 6813 11104
rect 8387 11096 8493 11104
rect 8507 11096 8893 11104
rect 11467 11096 11673 11104
rect 11687 11096 11713 11104
rect 207 11076 773 11084
rect 1487 11076 3913 11084
rect 4087 11076 4393 11084
rect 4447 11076 4473 11084
rect 4547 11076 6173 11084
rect 7407 11076 7593 11084
rect 7607 11076 7733 11084
rect 7747 11076 7773 11084
rect 11047 11076 11133 11084
rect 11147 11076 11353 11084
rect 1147 11056 1833 11064
rect 2007 11056 2133 11064
rect 2747 11056 3013 11064
rect 3087 11056 3553 11064
rect 4667 11056 4973 11064
rect 5147 11056 7133 11064
rect 7727 11056 7933 11064
rect 11167 11056 11253 11064
rect 11427 11056 11453 11064
rect 1767 11036 4193 11044
rect 4467 11036 5313 11044
rect 6947 11036 7053 11044
rect 7647 11036 9393 11044
rect 9907 11036 11533 11044
rect 11787 11036 11993 11044
rect 1187 11016 1213 11024
rect 1487 11016 1653 11024
rect 1667 11016 2773 11024
rect 2787 11016 4053 11024
rect 4367 11016 4413 11024
rect 4427 11016 6253 11024
rect 6747 11016 9933 11024
rect 11827 11016 11853 11024
rect 1087 10996 1213 11004
rect 1707 10996 2453 11004
rect 2467 10996 4473 11004
rect 6907 10996 8933 11004
rect 10767 10996 11293 11004
rect 11627 10996 12113 11004
rect 387 10976 953 10984
rect 967 10976 1573 10984
rect 1767 10976 1793 10984
rect 2027 10976 2633 10984
rect 2987 10976 3633 10984
rect 3687 10976 4293 10984
rect 4307 10976 5593 10984
rect 5887 10976 7033 10984
rect 9027 10976 9573 10984
rect 9587 10976 10313 10984
rect 11487 10976 11513 10984
rect 11987 10976 12133 10984
rect 1167 10956 2384 10964
rect 347 10936 413 10944
rect 427 10936 553 10944
rect 747 10936 1033 10944
rect 1327 10936 1553 10944
rect 1596 10936 2193 10944
rect 367 10916 513 10924
rect 607 10916 693 10924
rect 707 10916 813 10924
rect 827 10916 993 10924
rect 1127 10916 1153 10924
rect 1596 10924 1604 10936
rect 2207 10936 2353 10944
rect 2376 10944 2384 10956
rect 3327 10956 3373 10964
rect 4527 10956 5793 10964
rect 6867 10956 7173 10964
rect 7187 10956 7393 10964
rect 8967 10956 9173 10964
rect 9407 10956 9553 10964
rect 11087 10956 11433 10964
rect 11527 10956 11553 10964
rect 12016 10956 12173 10964
rect 2376 10936 2473 10944
rect 2667 10936 2913 10944
rect 3336 10936 3513 10944
rect 3336 10927 3344 10936
rect 3847 10936 4373 10944
rect 5087 10936 5853 10944
rect 5867 10936 5933 10944
rect 5967 10936 6084 10944
rect 6076 10927 6084 10936
rect 6987 10936 7013 10944
rect 7227 10936 7553 10944
rect 8607 10936 8853 10944
rect 8867 10936 9113 10944
rect 9176 10936 9513 10944
rect 1307 10916 1604 10924
rect 2007 10916 2193 10924
rect 2567 10916 2713 10924
rect 2927 10916 3113 10924
rect 3167 10916 3193 10924
rect 3887 10916 4113 10924
rect 4147 10916 4213 10924
rect 4227 10916 4373 10924
rect 5027 10916 5053 10924
rect 5807 10916 6033 10924
rect 6107 10916 6233 10924
rect 6307 10916 6373 10924
rect 6767 10916 7073 10924
rect 7247 10916 7353 10924
rect 7927 10916 8033 10924
rect 8727 10916 8753 10924
rect 8947 10916 8973 10924
rect 9047 10916 9153 10924
rect 247 10896 373 10904
rect 767 10896 913 10904
rect 947 10896 1013 10904
rect 1847 10896 2873 10904
rect 2947 10896 2973 10904
rect 3147 10896 3173 10904
rect 3267 10896 3313 10904
rect 3787 10896 4193 10904
rect 4207 10896 4433 10904
rect 4827 10896 4993 10904
rect 5007 10896 5153 10904
rect 5516 10904 5524 10913
rect 9176 10907 9184 10936
rect 9527 10936 9673 10944
rect 10127 10936 10173 10944
rect 10207 10936 10273 10944
rect 11167 10936 11213 10944
rect 11407 10936 11613 10944
rect 12016 10927 12024 10956
rect 9547 10916 9853 10924
rect 9927 10916 9973 10924
rect 10267 10916 10293 10924
rect 11036 10916 11173 10924
rect 5516 10896 6213 10904
rect 6687 10896 6773 10904
rect 7047 10896 7113 10904
rect 7127 10896 7333 10904
rect 7527 10896 7653 10904
rect 8187 10896 8253 10904
rect 8787 10896 8993 10904
rect 187 10876 413 10884
rect 587 10876 713 10884
rect 1507 10876 1613 10884
rect 1667 10876 1793 10884
rect 1807 10876 1953 10884
rect 2387 10876 2453 10884
rect 2487 10876 2533 10884
rect 2607 10876 2893 10884
rect 2907 10876 3093 10884
rect 3127 10876 3373 10884
rect 3707 10876 3853 10884
rect 4167 10876 4593 10884
rect 4627 10876 4793 10884
rect 4807 10876 5493 10884
rect 5547 10876 5693 10884
rect 5707 10876 7013 10884
rect 7387 10876 7773 10884
rect 8427 10876 8733 10884
rect 9196 10884 9204 10913
rect 9376 10904 9384 10913
rect 9227 10896 9384 10904
rect 9747 10896 10133 10904
rect 10656 10904 10664 10913
rect 11036 10907 11044 10916
rect 12107 10916 12173 10924
rect 10487 10896 10664 10904
rect 10867 10896 10993 10904
rect 11056 10896 11573 10904
rect 8747 10876 9204 10884
rect 10187 10876 10493 10884
rect 10707 10876 10833 10884
rect 11056 10884 11064 10896
rect 12027 10896 12073 10904
rect 11027 10876 11064 10884
rect 11387 10876 11453 10884
rect 11547 10876 11833 10884
rect 547 10856 573 10864
rect 1707 10856 2953 10864
rect 2967 10856 3213 10864
rect 3227 10856 3833 10864
rect 3887 10856 4033 10864
rect 4247 10856 4513 10864
rect 4647 10856 6853 10864
rect 7687 10856 7773 10864
rect 7967 10856 9413 10864
rect 2407 10836 3333 10844
rect 3467 10836 3713 10844
rect 3747 10836 3873 10844
rect 4427 10836 4833 10844
rect 4847 10836 5333 10844
rect 5347 10836 5593 10844
rect 5667 10836 5953 10844
rect 6067 10836 6133 10844
rect 6267 10836 6493 10844
rect 8247 10836 11233 10844
rect 11327 10836 11833 10844
rect 2747 10816 6093 10824
rect 6367 10816 6593 10824
rect 6787 10816 6993 10824
rect 7007 10816 7033 10824
rect 7047 10816 7473 10824
rect 7487 10816 7953 10824
rect 8467 10816 8933 10824
rect 9247 10816 11413 10824
rect 11967 10816 12053 10824
rect 1047 10796 2593 10804
rect 3207 10796 3793 10804
rect 4767 10796 7233 10804
rect 7427 10796 7853 10804
rect 8507 10796 9513 10804
rect 11487 10796 11573 10804
rect 2507 10776 2793 10784
rect 2887 10776 3633 10784
rect 4127 10776 5193 10784
rect 6007 10776 7573 10784
rect 7587 10776 7733 10784
rect 7747 10776 8393 10784
rect 8627 10776 8873 10784
rect 8907 10776 9353 10784
rect 9367 10776 10973 10784
rect 11467 10776 11693 10784
rect 1247 10756 1513 10764
rect 1527 10756 1633 10764
rect 2287 10756 3233 10764
rect 3287 10756 3733 10764
rect 3747 10756 3993 10764
rect 6147 10756 6613 10764
rect 7167 10756 7293 10764
rect 8927 10756 9013 10764
rect 10187 10756 10613 10764
rect 10767 10756 10813 10764
rect 11427 10756 11513 10764
rect 11647 10756 11913 10764
rect 1327 10736 1433 10744
rect 1447 10736 1813 10744
rect 1907 10736 1953 10744
rect 2007 10736 2073 10744
rect 2087 10736 2873 10744
rect 3147 10736 3233 10744
rect 3256 10736 3293 10744
rect 387 10716 493 10724
rect 507 10716 613 10724
rect 876 10724 884 10733
rect 707 10716 1464 10724
rect 1456 10707 1464 10716
rect 1487 10716 1524 10724
rect 727 10696 853 10704
rect 987 10696 1293 10704
rect 1516 10704 1524 10716
rect 2036 10716 2233 10724
rect 1516 10696 1873 10704
rect 2036 10704 2044 10716
rect 2527 10716 2813 10724
rect 2867 10716 2893 10724
rect 3256 10724 3264 10736
rect 3387 10736 3433 10744
rect 3547 10736 3653 10744
rect 4407 10736 4733 10744
rect 5267 10736 5373 10744
rect 5767 10736 5993 10744
rect 6287 10736 6393 10744
rect 7087 10736 7153 10744
rect 8067 10736 8233 10744
rect 8607 10736 8693 10744
rect 8727 10736 8773 10744
rect 8807 10736 8844 10744
rect 2987 10716 3264 10724
rect 3216 10707 3224 10716
rect 3307 10716 3393 10724
rect 3467 10716 3473 10724
rect 3487 10716 3613 10724
rect 4047 10716 4173 10724
rect 4187 10716 4253 10724
rect 4267 10716 4373 10724
rect 4427 10716 4473 10724
rect 4707 10716 6553 10724
rect 6607 10716 7113 10724
rect 7127 10716 7633 10724
rect 7687 10716 8013 10724
rect 8836 10724 8844 10736
rect 8867 10736 9013 10744
rect 9547 10736 9713 10744
rect 9887 10736 9913 10744
rect 9947 10736 10033 10744
rect 10047 10736 10233 10744
rect 10807 10736 11333 10744
rect 11507 10736 11613 10744
rect 11747 10736 11773 10744
rect 8327 10716 8984 10724
rect 1907 10696 2044 10704
rect 2067 10696 2213 10704
rect 2267 10696 2293 10704
rect 2307 10696 2693 10704
rect 2767 10696 3013 10704
rect 3276 10704 3284 10713
rect 8976 10707 8984 10716
rect 9007 10716 9133 10724
rect 9187 10716 9353 10724
rect 9376 10716 9393 10724
rect 3276 10696 3573 10704
rect 4027 10696 4113 10704
rect 4587 10696 4753 10704
rect 5316 10696 5353 10704
rect 1496 10684 1504 10693
rect 1496 10676 1673 10684
rect 1827 10676 1913 10684
rect 2447 10676 2893 10684
rect 3047 10676 3293 10684
rect 4216 10684 4224 10693
rect 3427 10676 4224 10684
rect 5316 10684 5324 10696
rect 5567 10696 5733 10704
rect 5867 10696 6173 10704
rect 6967 10696 7093 10704
rect 7187 10696 7273 10704
rect 7567 10696 7593 10704
rect 7607 10696 7793 10704
rect 7827 10696 8073 10704
rect 8207 10696 8253 10704
rect 8276 10696 8893 10704
rect 4247 10676 5324 10684
rect 5347 10676 5473 10684
rect 5487 10676 5533 10684
rect 5667 10676 5773 10684
rect 5787 10676 6373 10684
rect 8276 10684 8284 10696
rect 9376 10704 9384 10716
rect 9567 10716 9713 10724
rect 9767 10716 9893 10724
rect 10167 10716 10193 10724
rect 10807 10716 10873 10724
rect 10907 10716 11013 10724
rect 11047 10716 11193 10724
rect 11447 10716 11533 10724
rect 11567 10716 11633 10724
rect 11767 10716 12033 10724
rect 9327 10696 9384 10704
rect 10627 10696 10773 10704
rect 11227 10696 11553 10704
rect 11667 10696 11793 10704
rect 12047 10696 12133 10704
rect 8047 10676 8284 10684
rect 8447 10676 8713 10684
rect 9447 10676 9693 10684
rect 9747 10676 10053 10684
rect 10687 10676 11193 10684
rect 11207 10676 11313 10684
rect 11627 10676 11753 10684
rect 11767 10676 11893 10684
rect 11907 10676 12053 10684
rect 2847 10656 3073 10664
rect 3927 10656 3973 10664
rect 3987 10656 4313 10664
rect 5167 10656 5393 10664
rect 5827 10656 6413 10664
rect 7087 10656 7673 10664
rect 8747 10656 9473 10664
rect 9487 10656 10593 10664
rect 10647 10656 10853 10664
rect 11367 10656 11433 10664
rect 11447 10656 11733 10664
rect 11947 10656 12093 10664
rect 2367 10636 3253 10644
rect 3267 10636 3813 10644
rect 3827 10636 4633 10644
rect 7627 10636 8293 10644
rect 8307 10636 10593 10644
rect 12027 10636 12113 10644
rect 3007 10616 3133 10624
rect 10407 10616 10953 10624
rect 11147 10616 11193 10624
rect 11347 10616 11473 10624
rect 2287 10596 2393 10604
rect 10567 10596 12133 10604
rect 8347 10576 9053 10584
rect 10727 10576 10813 10584
rect 11147 10576 12173 10584
rect 7487 10556 8853 10564
rect 9507 10556 9533 10564
rect 11127 10556 11313 10564
rect 11327 10556 11393 10564
rect 11407 10556 11613 10564
rect 127 10536 173 10544
rect 4987 10536 5653 10544
rect 8167 10536 8453 10544
rect 8467 10536 8573 10544
rect 8987 10536 10073 10544
rect 11267 10536 11533 10544
rect 447 10516 1533 10524
rect 1547 10516 1973 10524
rect 3767 10516 4853 10524
rect 7967 10516 8373 10524
rect 8687 10516 9053 10524
rect 9467 10516 9713 10524
rect 10007 10516 10413 10524
rect 10607 10516 11513 10524
rect 11647 10516 11733 10524
rect 787 10496 2013 10504
rect 7687 10496 7833 10504
rect 7847 10496 8753 10504
rect 9187 10496 10113 10504
rect 10987 10496 11053 10504
rect 11307 10496 11513 10504
rect 11627 10496 11933 10504
rect 67 10476 433 10484
rect 847 10476 873 10484
rect 1187 10476 1833 10484
rect 3187 10476 3753 10484
rect 5047 10476 5393 10484
rect 6027 10476 7073 10484
rect 7927 10476 8013 10484
rect 8187 10476 8353 10484
rect 8827 10476 8873 10484
rect 8887 10476 9093 10484
rect 9107 10476 10893 10484
rect 11616 10476 11673 10484
rect -24 10456 113 10464
rect 287 10456 453 10464
rect 807 10456 1013 10464
rect 1027 10456 1173 10464
rect 2067 10456 2133 10464
rect 2147 10456 2353 10464
rect 2707 10456 2773 10464
rect 2787 10456 2933 10464
rect 2947 10456 3073 10464
rect 3087 10456 3253 10464
rect 3267 10456 3473 10464
rect 4367 10456 4893 10464
rect 5127 10456 5333 10464
rect 6387 10456 6633 10464
rect 7527 10456 7593 10464
rect 7616 10456 7744 10464
rect 147 10436 313 10444
rect 367 10436 384 10444
rect 376 10424 384 10436
rect 407 10436 473 10444
rect 847 10436 853 10444
rect 867 10436 973 10444
rect 987 10436 993 10444
rect 1047 10436 1093 10444
rect 1507 10436 1633 10444
rect 1896 10436 2313 10444
rect 376 10416 1793 10424
rect 1896 10424 1904 10436
rect 2327 10436 2473 10444
rect 2907 10436 3093 10444
rect 3627 10436 3793 10444
rect 4887 10436 5073 10444
rect 5087 10436 5293 10444
rect 5827 10436 5913 10444
rect 5947 10436 5973 10444
rect 6147 10436 6193 10444
rect 6207 10436 6333 10444
rect 6507 10436 6533 10444
rect 6547 10436 6733 10444
rect 6747 10436 6913 10444
rect 7616 10444 7624 10456
rect 7307 10436 7624 10444
rect 7676 10436 7713 10444
rect 1867 10416 1904 10424
rect 1927 10416 2073 10424
rect 2516 10424 2524 10433
rect 2387 10416 2524 10424
rect 2647 10416 2913 10424
rect 3527 10416 3633 10424
rect 3647 10416 3813 10424
rect 4647 10416 4713 10424
rect 4727 10416 4813 10424
rect 4827 10416 5033 10424
rect 5367 10416 5933 10424
rect 6307 10416 6753 10424
rect 6987 10416 6993 10424
rect 7007 10416 7353 10424
rect 7547 10416 7633 10424
rect 7676 10407 7684 10436
rect 7736 10444 7744 10456
rect 7907 10456 7973 10464
rect 8287 10456 8373 10464
rect 8667 10456 9273 10464
rect 9347 10456 9493 10464
rect 10076 10456 10093 10464
rect 7736 10436 7933 10444
rect 8047 10436 8093 10444
rect 8207 10436 8553 10444
rect 9267 10436 9333 10444
rect 9707 10436 9893 10444
rect 7747 10416 7813 10424
rect 7927 10416 7953 10424
rect 8127 10416 8213 10424
rect 8527 10416 8713 10424
rect 8787 10416 8893 10424
rect 8907 10416 8953 10424
rect 9287 10416 9453 10424
rect 9527 10416 9693 10424
rect 10076 10407 10084 10456
rect 10207 10456 10433 10464
rect 10547 10456 10613 10464
rect 11036 10456 11084 10464
rect 10307 10436 10433 10444
rect 10507 10436 10533 10444
rect 10676 10427 10684 10453
rect 10787 10436 10853 10444
rect 11036 10444 11044 10456
rect 10907 10436 11044 10444
rect 10127 10416 10453 10424
rect 187 10396 373 10404
rect 387 10396 433 10404
rect 2187 10396 2293 10404
rect 2447 10396 2533 10404
rect 2547 10396 3113 10404
rect 3687 10396 3913 10404
rect 4667 10396 4713 10404
rect 4967 10396 5093 10404
rect 5327 10396 5553 10404
rect 5927 10396 5953 10404
rect 6187 10396 6553 10404
rect 6967 10396 7013 10404
rect 7467 10396 7573 10404
rect 7747 10396 7933 10404
rect 7987 10396 8293 10404
rect 8307 10396 8333 10404
rect 8387 10396 8573 10404
rect 8587 10396 8673 10404
rect 8687 10396 9113 10404
rect 9147 10396 9293 10404
rect 9307 10396 9853 10404
rect 9967 10396 10053 10404
rect 10696 10404 10704 10433
rect 10727 10416 10833 10424
rect 10847 10416 10953 10424
rect 10447 10396 10704 10404
rect 11056 10404 11064 10433
rect 11076 10427 11084 10456
rect 11367 10456 11453 10464
rect 11616 10464 11624 10476
rect 12067 10476 12093 10484
rect 11596 10456 11624 10464
rect 11267 10436 11304 10444
rect 11296 10427 11304 10436
rect 11596 10444 11604 10456
rect 11667 10456 11713 10464
rect 12047 10456 12064 10464
rect 11476 10436 11604 10444
rect 11227 10416 11273 10424
rect 11327 10416 11373 10424
rect 11407 10416 11433 10424
rect 11056 10396 11213 10404
rect 11456 10404 11464 10433
rect 11476 10427 11484 10436
rect 11707 10436 11753 10444
rect 11947 10436 12033 10444
rect 12056 10427 12064 10456
rect 11507 10416 11673 10424
rect 11767 10416 11773 10424
rect 11787 10416 11853 10424
rect 11387 10396 11464 10404
rect 11607 10396 11673 10404
rect 2487 10376 2673 10384
rect 4427 10376 4513 10384
rect 4527 10376 5053 10384
rect 5747 10376 5853 10384
rect 6527 10376 6713 10384
rect 6727 10376 6973 10384
rect 7087 10376 7593 10384
rect 7607 10376 7693 10384
rect 8027 10376 8153 10384
rect 8607 10376 8713 10384
rect 9207 10376 9653 10384
rect 9887 10376 10473 10384
rect 10507 10376 10653 10384
rect 10707 10376 10733 10384
rect 10887 10376 11153 10384
rect 11896 10384 11904 10413
rect 11287 10376 11904 10384
rect 11927 10376 11953 10384
rect 2127 10356 2393 10364
rect 3567 10356 4673 10364
rect 5067 10356 6313 10364
rect 7367 10356 8133 10364
rect 8547 10356 9133 10364
rect 9867 10356 10533 10364
rect 10547 10356 10773 10364
rect 11667 10356 11713 10364
rect 11727 10356 11793 10364
rect 11847 10356 11893 10364
rect 207 10336 333 10344
rect 1387 10336 1713 10344
rect 2167 10336 2333 10344
rect 4547 10336 4753 10344
rect 4767 10336 5273 10344
rect 5667 10336 7133 10344
rect 7147 10336 7313 10344
rect 7327 10336 8813 10344
rect 9447 10336 10273 10344
rect 10327 10336 10513 10344
rect 10527 10336 10633 10344
rect 10687 10336 10933 10344
rect 11867 10336 11993 10344
rect 807 10316 1513 10324
rect 1547 10316 1953 10324
rect 2327 10316 2653 10324
rect 3407 10316 3773 10324
rect 5287 10316 6113 10324
rect 7347 10316 7453 10324
rect 7467 10316 7953 10324
rect 7967 10316 8073 10324
rect 8707 10316 9193 10324
rect 9227 10316 10153 10324
rect 10167 10316 10313 10324
rect 10347 10316 10493 10324
rect 10587 10316 10893 10324
rect 11787 10316 11933 10324
rect 1147 10296 1333 10304
rect 1607 10296 1613 10304
rect 1627 10296 1733 10304
rect 1947 10296 3053 10304
rect 3267 10296 3533 10304
rect 3707 10296 3973 10304
rect 4167 10296 4213 10304
rect 5247 10296 5273 10304
rect 5407 10296 5433 10304
rect 5687 10296 6153 10304
rect 6327 10296 6413 10304
rect 6927 10296 8393 10304
rect 8527 10296 8633 10304
rect 8767 10296 10793 10304
rect 11067 10296 11133 10304
rect 11407 10296 11713 10304
rect 11727 10296 11953 10304
rect 1207 10276 2333 10284
rect 2347 10276 2793 10284
rect 2807 10276 2813 10284
rect 2827 10276 4093 10284
rect 4107 10276 4993 10284
rect 5007 10276 5173 10284
rect 5187 10276 5353 10284
rect 5367 10276 5853 10284
rect 5867 10276 6133 10284
rect 6347 10276 7033 10284
rect 7107 10276 7173 10284
rect 7247 10276 7493 10284
rect 7887 10276 7913 10284
rect 7927 10276 7993 10284
rect 8007 10276 9013 10284
rect 9027 10276 9113 10284
rect 9507 10276 9673 10284
rect 9687 10276 9733 10284
rect 10007 10276 10873 10284
rect 11047 10276 11633 10284
rect 11947 10276 11973 10284
rect 11987 10276 11993 10284
rect 1087 10256 1173 10264
rect 1607 10256 1673 10264
rect 1696 10256 2053 10264
rect 687 10236 833 10244
rect 847 10236 1133 10244
rect 1356 10236 1653 10244
rect 1356 10227 1364 10236
rect 1667 10236 1673 10244
rect 1696 10227 1704 10256
rect 2927 10256 3033 10264
rect 3467 10256 3633 10264
rect 3687 10256 3933 10264
rect 4007 10256 4153 10264
rect 4187 10256 4353 10264
rect 4587 10256 4813 10264
rect 5147 10256 5173 10264
rect 5236 10256 5433 10264
rect 1967 10236 3153 10244
rect 3327 10236 3433 10244
rect 3487 10236 3693 10244
rect 3827 10236 3873 10244
rect 3947 10236 4133 10244
rect 4147 10236 4253 10244
rect 4327 10236 4373 10244
rect 5236 10244 5244 10256
rect 6167 10256 6353 10264
rect 6447 10256 6553 10264
rect 6907 10256 7053 10264
rect 7067 10256 7193 10264
rect 7207 10256 7273 10264
rect 7287 10256 7513 10264
rect 7527 10256 7693 10264
rect 7707 10256 7753 10264
rect 7827 10256 8193 10264
rect 8607 10256 8653 10264
rect 8807 10256 8833 10264
rect 8867 10256 8953 10264
rect 8967 10256 9453 10264
rect 9587 10256 9833 10264
rect 10147 10256 10253 10264
rect 10327 10256 10393 10264
rect 10627 10256 10713 10264
rect 10767 10256 10793 10264
rect 10927 10256 10953 10264
rect 11107 10256 11113 10264
rect 11127 10256 11233 10264
rect 11427 10256 11473 10264
rect 11647 10256 12013 10264
rect 12047 10256 12133 10264
rect 4607 10236 5244 10244
rect 5487 10236 6513 10244
rect 6747 10236 6893 10244
rect 6967 10236 7073 10244
rect 7087 10236 7213 10244
rect 7907 10236 7933 10244
rect 8067 10236 8133 10244
rect 8567 10236 8633 10244
rect 8647 10236 8673 10244
rect 8807 10236 8913 10244
rect 8927 10236 9213 10244
rect 9567 10236 9653 10244
rect 9687 10236 10073 10244
rect 10356 10236 10493 10244
rect 387 10216 393 10224
rect 407 10216 493 10224
rect 647 10216 773 10224
rect 947 10216 993 10224
rect 1067 10216 1193 10224
rect 1747 10216 1853 10224
rect 2967 10216 3053 10224
rect 3067 10216 3073 10224
rect 3107 10216 3413 10224
rect 3667 10216 3793 10224
rect 3807 10216 3953 10224
rect 3967 10216 4153 10224
rect 4207 10216 4233 10224
rect 4347 10216 4393 10224
rect 4407 10216 4553 10224
rect 5256 10224 5264 10233
rect 5087 10216 5413 10224
rect 5947 10216 6593 10224
rect 6787 10216 6933 10224
rect 6947 10216 7153 10224
rect 7856 10224 7864 10233
rect 7327 10216 7973 10224
rect 8187 10216 8213 10224
rect 8396 10224 8404 10233
rect 10356 10227 10364 10236
rect 10507 10236 11213 10244
rect 11447 10236 11773 10244
rect 11987 10236 12153 10244
rect 8396 10216 8573 10224
rect 9007 10216 9253 10224
rect 9427 10216 9873 10224
rect 10547 10216 10693 10224
rect 11067 10216 11373 10224
rect 11416 10216 11433 10224
rect 427 10196 973 10204
rect 1027 10196 1153 10204
rect 1167 10196 1433 10204
rect 1567 10196 1593 10204
rect 2007 10196 2473 10204
rect 3247 10196 3453 10204
rect 5047 10196 5513 10204
rect 5527 10196 5653 10204
rect 5667 10196 5833 10204
rect 5847 10196 5993 10204
rect 6007 10196 6453 10204
rect 6467 10196 6653 10204
rect 6727 10196 7453 10204
rect 7767 10196 8013 10204
rect 8036 10204 8044 10213
rect 8036 10196 8213 10204
rect 8467 10196 9133 10204
rect 9467 10196 10513 10204
rect 10767 10196 10893 10204
rect 11267 10196 11393 10204
rect 11416 10187 11424 10216
rect 11507 10216 11553 10224
rect 12127 10216 12153 10224
rect 11467 10196 11553 10204
rect 11727 10196 11773 10204
rect 11827 10196 11873 10204
rect 3387 10176 3633 10184
rect 4247 10176 5053 10184
rect 5067 10176 5193 10184
rect 5947 10176 6493 10184
rect 8027 10176 8773 10184
rect 8887 10176 9693 10184
rect 9987 10176 10393 10184
rect 10707 10176 11213 10184
rect 11227 10176 11233 10184
rect 11827 10176 11893 10184
rect 4607 10156 4793 10164
rect 8067 10156 9033 10164
rect 9267 10156 9493 10164
rect 10827 10156 11633 10164
rect 11687 10156 11973 10164
rect 2296 10124 2304 10153
rect 5287 10136 5753 10144
rect 8427 10136 8473 10144
rect 8487 10136 9173 10144
rect 9187 10136 9764 10144
rect 2267 10116 2304 10124
rect 7467 10116 8733 10124
rect 9067 10116 9453 10124
rect 9756 10124 9764 10136
rect 9827 10136 10553 10144
rect 10567 10136 10773 10144
rect 11927 10136 12013 10144
rect 9756 10116 10113 10124
rect 10127 10116 10533 10124
rect 10747 10116 10913 10124
rect 11047 10116 11153 10124
rect 11347 10116 11433 10124
rect 5467 10096 5933 10104
rect 6407 10096 6573 10104
rect 6587 10096 10313 10104
rect 1807 10076 6493 10084
rect 8307 10076 8613 10084
rect 9147 10076 9333 10084
rect 9547 10076 9573 10084
rect 9667 10076 11653 10084
rect 627 10056 653 10064
rect 1947 10056 2293 10064
rect 2307 10056 2373 10064
rect 2387 10056 2573 10064
rect 2587 10056 3233 10064
rect 6807 10056 6853 10064
rect 7887 10056 8484 10064
rect 587 10036 3553 10044
rect 7847 10036 8093 10044
rect 8127 10036 8453 10044
rect 8476 10044 8484 10056
rect 8587 10056 9233 10064
rect 9256 10056 9833 10064
rect 9256 10044 9264 10056
rect 10887 10056 11013 10064
rect 11027 10056 11093 10064
rect 8476 10036 9264 10044
rect 9347 10036 9873 10044
rect 10427 10036 11253 10044
rect 11267 10036 11273 10044
rect 3327 10016 3453 10024
rect 7727 10016 8013 10024
rect 8027 10016 8844 10024
rect 447 9996 613 10004
rect 627 9996 1293 10004
rect 2227 9996 2473 10004
rect 2487 9996 2673 10004
rect 2687 9996 3173 10004
rect 4167 9996 4373 10004
rect 7987 9996 8073 10004
rect 8287 9996 8813 10004
rect 8836 10004 8844 10016
rect 9207 10016 9293 10024
rect 9307 10016 10093 10024
rect 10107 10016 10693 10024
rect 10947 10016 11073 10024
rect 11387 10016 11753 10024
rect 8836 9996 9933 10004
rect 10087 9996 10153 10004
rect 10167 9996 10393 10004
rect 10907 9996 10973 10004
rect 11207 9996 11273 10004
rect 607 9976 1853 9984
rect 3587 9976 3673 9984
rect 6467 9976 6713 9984
rect 7127 9976 7153 9984
rect 7607 9976 7653 9984
rect 8007 9976 8053 9984
rect 8067 9976 8393 9984
rect 8447 9976 8493 9984
rect 9087 9976 9153 9984
rect 9467 9976 9553 9984
rect 10127 9976 10593 9984
rect 10787 9976 10953 9984
rect 10967 9976 11004 9984
rect 87 9956 733 9964
rect 796 9956 913 9964
rect 796 9947 804 9956
rect 927 9956 993 9964
rect 1287 9956 1353 9964
rect 1367 9956 1393 9964
rect 1427 9956 1493 9964
rect 1547 9956 1593 9964
rect 1687 9956 1713 9964
rect 2107 9956 2133 9964
rect 2447 9956 2533 9964
rect 2647 9956 2713 9964
rect 3107 9956 3213 9964
rect 3667 9956 3853 9964
rect 4427 9956 4513 9964
rect 4567 9956 4713 9964
rect 4727 9956 4933 9964
rect 5456 9956 5613 9964
rect 67 9936 373 9944
rect 1027 9936 1033 9944
rect 1047 9936 1133 9944
rect 1756 9944 1764 9953
rect 1487 9936 1813 9944
rect 1827 9936 1953 9944
rect 1967 9936 2073 9944
rect 2507 9936 2613 9944
rect 3027 9936 3493 9944
rect 3507 9936 3533 9944
rect 3747 9936 3793 9944
rect 4267 9936 4353 9944
rect 4367 9936 4413 9944
rect 4427 9936 4753 9944
rect 5456 9944 5464 9956
rect 5627 9956 5733 9964
rect 6427 9956 6553 9964
rect 6767 9956 6873 9964
rect 7307 9956 7333 9964
rect 7427 9956 7673 9964
rect 7687 9956 7753 9964
rect 8227 9956 8413 9964
rect 8427 9956 8593 9964
rect 8647 9956 9273 9964
rect 9387 9956 9493 9964
rect 9547 9956 10604 9964
rect 5007 9936 5464 9944
rect 6687 9936 7333 9944
rect 7487 9936 7693 9944
rect 7707 9936 7833 9944
rect 8047 9936 8233 9944
rect 8267 9936 8613 9944
rect 8747 9936 8953 9944
rect 9727 9936 9833 9944
rect 9947 9936 10073 9944
rect 10087 9936 10293 9944
rect 10596 9944 10604 9956
rect 10627 9956 10773 9964
rect 10996 9964 11004 9976
rect 11027 9976 11113 9984
rect 11576 9967 11584 9993
rect 11596 9976 11733 9984
rect 10996 9956 11113 9964
rect 11167 9956 11213 9964
rect 10596 9936 10633 9944
rect 10827 9936 10973 9944
rect 11087 9936 11173 9944
rect 11267 9936 11333 9944
rect 11467 9936 11484 9944
rect 487 9916 633 9924
rect 1107 9916 1333 9924
rect 1647 9916 1693 9924
rect 1907 9916 1933 9924
rect 2467 9916 2693 9924
rect 2847 9916 2993 9924
rect 3327 9916 3473 9924
rect 3607 9916 3873 9924
rect 3987 9916 4313 9924
rect 4407 9916 4573 9924
rect 4627 9916 4693 9924
rect 4927 9916 5073 9924
rect 5487 9916 5493 9924
rect 5507 9916 5593 9924
rect 5867 9916 5973 9924
rect 6647 9916 6873 9924
rect 7167 9916 7273 9924
rect 7347 9916 7433 9924
rect 7847 9916 8653 9924
rect 8667 9916 8733 9924
rect 8747 9916 8773 9924
rect 8807 9916 8833 9924
rect 9367 9916 9613 9924
rect 9767 9916 9853 9924
rect 9867 9916 9913 9924
rect 10167 9916 10253 9924
rect 10287 9916 10433 9924
rect 10667 9916 10753 9924
rect 10767 9916 10833 9924
rect 11147 9916 11413 9924
rect 11427 9916 11453 9924
rect 1527 9896 1673 9904
rect 1867 9896 1913 9904
rect 2607 9896 2973 9904
rect 4967 9896 5193 9904
rect 5927 9896 5973 9904
rect 6307 9896 6513 9904
rect 7667 9896 7993 9904
rect 8087 9896 9173 9904
rect 9327 9896 10293 9904
rect 10307 9896 10413 9904
rect 10507 9896 10733 9904
rect 11247 9896 11393 9904
rect 11476 9904 11484 9936
rect 11596 9944 11604 9976
rect 11567 9936 11604 9944
rect 11747 9936 12033 9944
rect 11627 9916 11713 9924
rect 11947 9916 12073 9924
rect 11427 9896 11484 9904
rect 11627 9896 11673 9904
rect 11707 9896 11993 9904
rect 987 9876 1113 9884
rect 1227 9876 1513 9884
rect 2127 9876 2633 9884
rect 2787 9876 3013 9884
rect 3547 9876 4153 9884
rect 4167 9876 4193 9884
rect 4807 9876 5673 9884
rect 7507 9876 7653 9884
rect 8227 9876 8273 9884
rect 9007 9876 9813 9884
rect 10867 9876 10913 9884
rect 10927 9876 11033 9884
rect 11187 9876 11433 9884
rect 11647 9876 11673 9884
rect 1387 9856 1793 9864
rect 3307 9856 3333 9864
rect 3367 9856 3453 9864
rect 3627 9856 5113 9864
rect 5307 9856 5353 9864
rect 5967 9856 6213 9864
rect 6967 9856 7253 9864
rect 7267 9856 8293 9864
rect 8607 9856 8833 9864
rect 9447 9856 9733 9864
rect 9787 9856 9873 9864
rect 10427 9856 11193 9864
rect 11387 9856 11573 9864
rect 647 9836 1633 9844
rect 1947 9836 7853 9844
rect 7947 9836 8113 9844
rect 8367 9836 11053 9844
rect 11067 9836 11233 9844
rect 11547 9836 11633 9844
rect 707 9816 1153 9824
rect 1167 9816 1433 9824
rect 1647 9816 2133 9824
rect 3787 9816 4253 9824
rect 5187 9816 5313 9824
rect 5827 9816 5953 9824
rect 7207 9816 9773 9824
rect 10507 9816 11413 9824
rect 1007 9796 1853 9804
rect 1867 9796 1953 9804
rect 3727 9796 3773 9804
rect 5827 9796 5873 9804
rect 5887 9796 6073 9804
rect 7007 9796 7173 9804
rect 7187 9796 7273 9804
rect 7287 9796 7313 9804
rect 7527 9796 7633 9804
rect 8107 9796 8524 9804
rect 167 9776 333 9784
rect 347 9776 353 9784
rect 367 9776 573 9784
rect 927 9776 993 9784
rect 1607 9776 2553 9784
rect 3227 9776 3253 9784
rect 3727 9776 3793 9784
rect 3827 9776 3913 9784
rect 4027 9776 4453 9784
rect 5487 9776 5884 9784
rect 87 9756 193 9764
rect 407 9756 593 9764
rect 607 9756 693 9764
rect 747 9756 953 9764
rect 1187 9756 1233 9764
rect 1247 9756 1413 9764
rect 2047 9756 2113 9764
rect 2156 9756 2293 9764
rect 2156 9747 2164 9756
rect 3787 9756 3993 9764
rect 4387 9756 4413 9764
rect 4887 9756 5293 9764
rect 5876 9764 5884 9776
rect 5907 9776 6053 9784
rect 6067 9776 6533 9784
rect 6787 9776 6973 9784
rect 6987 9776 7553 9784
rect 7587 9776 7853 9784
rect 7927 9776 7953 9784
rect 8516 9784 8524 9796
rect 8627 9796 8693 9804
rect 8807 9796 8973 9804
rect 9047 9796 9133 9804
rect 9207 9796 10173 9804
rect 10467 9796 11213 9804
rect 11407 9796 11753 9804
rect 11767 9796 12053 9804
rect 8516 9776 8673 9784
rect 8767 9776 8813 9784
rect 8967 9776 8993 9784
rect 9007 9776 9033 9784
rect 9187 9776 9393 9784
rect 9627 9776 9893 9784
rect 9927 9776 10364 9784
rect 5876 9756 6013 9764
rect 6227 9756 6384 9764
rect 627 9736 653 9744
rect 667 9736 753 9744
rect 827 9736 1013 9744
rect 1407 9736 1573 9744
rect 1587 9736 1733 9744
rect 2267 9736 2393 9744
rect 2587 9736 2773 9744
rect 3107 9736 3213 9744
rect 3227 9736 3233 9744
rect 3767 9736 3893 9744
rect 3927 9736 4433 9744
rect 4476 9744 4484 9753
rect 6376 9747 6384 9756
rect 6407 9756 6453 9764
rect 6667 9756 6813 9764
rect 7507 9756 7653 9764
rect 7727 9756 7893 9764
rect 8087 9756 8433 9764
rect 8647 9756 8653 9764
rect 8667 9756 8773 9764
rect 8827 9756 8993 9764
rect 9247 9756 9413 9764
rect 9807 9756 10333 9764
rect 10356 9764 10364 9776
rect 10387 9776 10713 9784
rect 10727 9776 10753 9784
rect 11207 9776 11273 9784
rect 11347 9776 11573 9784
rect 11587 9776 11893 9784
rect 12007 9776 12133 9784
rect 10356 9756 10893 9764
rect 10967 9756 11013 9764
rect 11447 9756 11493 9764
rect 11707 9756 11733 9764
rect 11916 9756 11993 9764
rect 4447 9736 4484 9744
rect 4527 9736 4953 9744
rect 4967 9736 5133 9744
rect 5927 9736 5993 9744
rect 807 9716 973 9724
rect 1287 9716 1413 9724
rect 1627 9716 1773 9724
rect 3627 9716 5073 9724
rect 6027 9716 6333 9724
rect 6616 9724 6624 9753
rect 6847 9736 6873 9744
rect 7587 9736 7644 9744
rect 6587 9716 6624 9724
rect 6807 9716 7033 9724
rect 7187 9716 7393 9724
rect 7636 9724 7644 9736
rect 7847 9736 7873 9744
rect 7887 9736 7973 9744
rect 8287 9736 8373 9744
rect 8707 9736 8853 9744
rect 8987 9736 9153 9744
rect 9307 9736 9333 9744
rect 9427 9736 9653 9744
rect 9667 9736 9973 9744
rect 10607 9736 10904 9744
rect 7636 9716 8213 9724
rect 8276 9716 8873 9724
rect 1307 9696 1373 9704
rect 1567 9696 2273 9704
rect 3627 9696 3833 9704
rect 3847 9696 3853 9704
rect 3867 9696 4533 9704
rect 6467 9696 6633 9704
rect 7547 9696 7913 9704
rect 8276 9704 8284 9716
rect 9027 9716 9293 9724
rect 10487 9716 10553 9724
rect 10567 9716 10693 9724
rect 10896 9724 10904 9736
rect 10927 9736 11013 9744
rect 11067 9736 11153 9744
rect 11507 9736 11593 9744
rect 11747 9736 11773 9744
rect 11916 9727 11924 9756
rect 11947 9736 11973 9744
rect 10896 9716 11073 9724
rect 11707 9716 11753 9724
rect 11807 9716 11913 9724
rect 11967 9716 12153 9724
rect 7927 9696 8284 9704
rect 8307 9696 8553 9704
rect 8567 9696 8773 9704
rect 9127 9696 9453 9704
rect 10507 9696 10573 9704
rect 10727 9696 12073 9704
rect 1887 9676 2233 9684
rect 4587 9676 6473 9684
rect 6487 9676 6953 9684
rect 7507 9676 8053 9684
rect 8396 9676 9213 9684
rect 4267 9656 6153 9664
rect 6607 9656 7173 9664
rect 7227 9656 7673 9664
rect 8396 9664 8404 9676
rect 9387 9676 10993 9684
rect 11887 9676 11933 9684
rect 7767 9656 8404 9664
rect 8427 9656 8853 9664
rect 9087 9656 9953 9664
rect 10047 9656 11713 9664
rect 87 9636 1993 9644
rect 2207 9636 2353 9644
rect 3727 9636 3933 9644
rect 6447 9636 6973 9644
rect 7047 9636 7493 9644
rect 7527 9636 9633 9644
rect 11007 9636 11373 9644
rect 3707 9616 5113 9624
rect 8747 9616 8913 9624
rect 8927 9616 8993 9624
rect 10767 9616 11733 9624
rect 11747 9616 11813 9624
rect 227 9596 513 9604
rect 527 9596 1053 9604
rect 1347 9596 1573 9604
rect 4007 9596 4713 9604
rect 5787 9596 7213 9604
rect 7867 9596 8433 9604
rect 8887 9596 9893 9604
rect 9907 9596 9933 9604
rect 10847 9596 11253 9604
rect 447 9576 973 9584
rect 987 9576 1193 9584
rect 1667 9576 1973 9584
rect 3147 9576 3373 9584
rect 3687 9576 3953 9584
rect 6427 9576 7413 9584
rect 8027 9576 8193 9584
rect 9127 9576 9913 9584
rect 9927 9576 10433 9584
rect 10447 9576 11493 9584
rect 1907 9556 3973 9564
rect 3987 9556 5893 9564
rect 7347 9556 8393 9564
rect 8407 9556 9513 9564
rect 9567 9556 10653 9564
rect 1667 9536 1833 9544
rect 1847 9536 2913 9544
rect 3087 9536 5633 9544
rect 6167 9536 9173 9544
rect 9527 9536 9733 9544
rect 9747 9536 10013 9544
rect 10787 9536 10853 9544
rect 11207 9536 11233 9544
rect 11367 9536 11433 9544
rect 11607 9536 12093 9544
rect 3387 9516 3573 9524
rect 3587 9516 3613 9524
rect 4287 9516 4513 9524
rect 4527 9516 4633 9524
rect 4687 9516 4933 9524
rect 5127 9516 6013 9524
rect 7287 9516 7333 9524
rect 8147 9516 8193 9524
rect 8327 9516 8373 9524
rect 8827 9516 9113 9524
rect 9167 9516 9573 9524
rect 9967 9516 10573 9524
rect 10587 9516 10713 9524
rect 10767 9516 10793 9524
rect 11207 9516 11273 9524
rect 11287 9516 11353 9524
rect 11427 9516 11473 9524
rect 11767 9516 11913 9524
rect 1907 9496 1993 9504
rect 2287 9496 2313 9504
rect 2387 9496 2453 9504
rect 2467 9496 3313 9504
rect 3327 9496 3513 9504
rect 4167 9496 4293 9504
rect 4387 9496 4553 9504
rect 4567 9496 4673 9504
rect 4847 9496 4893 9504
rect 5227 9496 5713 9504
rect 5727 9496 5793 9504
rect 5847 9496 5873 9504
rect 6327 9496 6353 9504
rect 7027 9496 7473 9504
rect 7567 9496 7733 9504
rect 8147 9496 8333 9504
rect 8467 9496 8813 9504
rect 8867 9496 9213 9504
rect 9227 9496 9393 9504
rect 9407 9496 10033 9504
rect 10247 9496 10313 9504
rect 10687 9496 10713 9504
rect 10847 9496 10873 9504
rect 11487 9496 11513 9504
rect 11567 9496 11593 9504
rect 11707 9496 11873 9504
rect 11927 9496 12053 9504
rect 567 9476 593 9484
rect 807 9476 1004 9484
rect 996 9467 1004 9476
rect 1407 9476 1433 9484
rect 1487 9476 1613 9484
rect 1727 9476 2033 9484
rect 2547 9476 2613 9484
rect 3107 9476 3233 9484
rect 3287 9476 3353 9484
rect 3487 9476 3633 9484
rect 3747 9476 3873 9484
rect 4207 9476 4353 9484
rect 4507 9476 4533 9484
rect 4767 9476 4913 9484
rect 5087 9476 5213 9484
rect 5227 9476 5304 9484
rect 5296 9467 5304 9476
rect 5407 9476 5473 9484
rect 5827 9476 5893 9484
rect 5927 9476 6173 9484
rect 6227 9476 6373 9484
rect 6747 9476 6833 9484
rect 6887 9476 6933 9484
rect 6987 9476 7033 9484
rect 7056 9476 7153 9484
rect -24 9456 113 9464
rect 187 9456 813 9464
rect 1007 9456 1373 9464
rect 1607 9456 1873 9464
rect 1976 9456 2093 9464
rect 967 9436 1093 9444
rect 1447 9436 1633 9444
rect 1647 9436 1673 9444
rect 1867 9436 1913 9444
rect 1976 9444 1984 9456
rect 2667 9456 3053 9464
rect 3347 9456 3433 9464
rect 4287 9456 4733 9464
rect 5067 9456 5253 9464
rect 5447 9456 5493 9464
rect 5627 9456 5673 9464
rect 6167 9456 6413 9464
rect 6607 9456 6713 9464
rect 7056 9464 7064 9476
rect 7207 9476 7364 9484
rect 7356 9467 7364 9476
rect 7487 9476 7533 9484
rect 7607 9476 7713 9484
rect 8047 9476 8073 9484
rect 8127 9476 8413 9484
rect 9027 9476 9493 9484
rect 9907 9476 9933 9484
rect 10647 9476 10753 9484
rect 10767 9476 10813 9484
rect 11007 9476 11024 9484
rect 6967 9456 7064 9464
rect 7587 9456 7613 9464
rect 7756 9464 7764 9473
rect 7736 9456 7764 9464
rect 1927 9436 1984 9444
rect 2007 9436 2073 9444
rect 2467 9436 2593 9444
rect 3027 9436 3113 9444
rect 3127 9436 3593 9444
rect 3747 9436 4173 9444
rect 4227 9436 5413 9444
rect 5427 9436 6213 9444
rect 6527 9436 6753 9444
rect 6847 9436 7133 9444
rect 7347 9436 7553 9444
rect 7736 9444 7744 9456
rect 7867 9456 7893 9464
rect 8036 9456 8053 9464
rect 7707 9436 7744 9444
rect 7767 9436 7913 9444
rect 7967 9436 7993 9444
rect 8036 9444 8044 9456
rect 8227 9456 8273 9464
rect 8287 9456 8293 9464
rect 8527 9456 8593 9464
rect 8647 9456 8673 9464
rect 8867 9456 8933 9464
rect 9207 9456 9333 9464
rect 9667 9456 9713 9464
rect 9967 9456 9993 9464
rect 10667 9456 10773 9464
rect 10847 9456 10893 9464
rect 10907 9456 10973 9464
rect 11016 9447 11024 9476
rect 11047 9476 11193 9484
rect 11307 9476 11533 9484
rect 11627 9476 11733 9484
rect 11747 9476 11773 9484
rect 11407 9456 11513 9464
rect 11567 9456 11593 9464
rect 11807 9456 11873 9464
rect 8007 9436 8044 9444
rect 8067 9436 8253 9444
rect 8327 9436 8633 9444
rect 8667 9436 8773 9444
rect 8867 9436 9073 9444
rect 9127 9436 9233 9444
rect 9607 9436 9613 9444
rect 9627 9436 9733 9444
rect 10127 9436 10253 9444
rect 10356 9436 10413 9444
rect 2187 9416 3073 9424
rect 4307 9416 4933 9424
rect 6047 9416 6193 9424
rect 6567 9416 6773 9424
rect 7947 9416 8313 9424
rect 8347 9416 8473 9424
rect 8507 9416 8793 9424
rect 10356 9424 10364 9436
rect 10427 9436 10613 9444
rect 10627 9436 10633 9444
rect 10787 9436 10913 9444
rect 11167 9436 11193 9444
rect 11387 9436 11573 9444
rect 11727 9436 11753 9444
rect 11907 9436 12033 9444
rect 8947 9416 10364 9424
rect 10407 9416 10873 9424
rect 10887 9416 11213 9424
rect 11227 9416 11993 9424
rect 2167 9396 4133 9404
rect 4147 9396 5653 9404
rect 5947 9396 6973 9404
rect 7287 9396 8093 9404
rect 8327 9396 8353 9404
rect 8427 9396 10113 9404
rect 11187 9396 11333 9404
rect 667 9376 1113 9384
rect 1127 9376 1313 9384
rect 2447 9376 2773 9384
rect 3247 9376 6013 9384
rect 7047 9376 7133 9384
rect 7147 9376 7173 9384
rect 7387 9376 9053 9384
rect 9367 9376 9413 9384
rect 10367 9376 11613 9384
rect 11627 9376 12073 9384
rect 887 9356 1133 9364
rect 1547 9356 2373 9364
rect 2727 9356 3133 9364
rect 3267 9356 3853 9364
rect 4027 9356 4313 9364
rect 4327 9356 4613 9364
rect 6467 9356 6873 9364
rect 7647 9356 8033 9364
rect 8487 9356 9313 9364
rect 9467 9356 9913 9364
rect 10087 9356 10193 9364
rect 11147 9356 11213 9364
rect 907 9336 1033 9344
rect 1467 9336 1693 9344
rect 2487 9336 2533 9344
rect 3167 9336 3293 9344
rect 3327 9336 3553 9344
rect 5887 9336 6433 9344
rect 6627 9336 7473 9344
rect 8647 9336 10133 9344
rect 10607 9336 10773 9344
rect 10947 9336 10993 9344
rect 727 9316 1433 9324
rect 2027 9316 2333 9324
rect 3507 9316 3633 9324
rect 4647 9316 4873 9324
rect 5267 9316 5353 9324
rect 6087 9316 6413 9324
rect 6427 9316 6753 9324
rect 6767 9316 7473 9324
rect 7487 9316 7593 9324
rect 8047 9316 8093 9324
rect 8447 9316 9753 9324
rect 10207 9316 10273 9324
rect 10827 9316 10953 9324
rect 11247 9316 11333 9324
rect 167 9296 393 9304
rect 407 9296 553 9304
rect 567 9296 733 9304
rect 747 9296 773 9304
rect 847 9296 913 9304
rect 1167 9296 1493 9304
rect 1507 9296 1553 9304
rect 1727 9296 2013 9304
rect 2267 9296 2973 9304
rect 4687 9296 4853 9304
rect 5487 9296 5913 9304
rect 6107 9296 6173 9304
rect 6287 9296 6593 9304
rect 6807 9296 6833 9304
rect 7007 9296 7513 9304
rect 7587 9296 7644 9304
rect 387 9276 513 9284
rect 887 9276 1173 9284
rect 1227 9276 1453 9284
rect 1847 9276 1973 9284
rect 2047 9276 2173 9284
rect 2607 9276 2793 9284
rect 2807 9276 3333 9284
rect 3347 9276 3813 9284
rect 3827 9276 3913 9284
rect 3927 9276 4453 9284
rect 4467 9276 4653 9284
rect 347 9256 493 9264
rect 747 9256 933 9264
rect 947 9256 1153 9264
rect 1267 9256 1293 9264
rect 1487 9256 1533 9264
rect 1547 9256 1633 9264
rect 1807 9256 2193 9264
rect 156 9244 164 9253
rect 2216 9247 2224 9273
rect 2247 9256 2413 9264
rect 2456 9264 2464 9273
rect 5276 9267 5284 9293
rect 5307 9276 5333 9284
rect 5476 9276 5513 9284
rect 2456 9256 2513 9264
rect 3527 9256 3613 9264
rect 3907 9256 4013 9264
rect 4727 9256 5033 9264
rect 5087 9256 5113 9264
rect 156 9236 313 9244
rect 367 9236 393 9244
rect 547 9236 593 9244
rect 607 9236 1093 9244
rect 1207 9236 1233 9244
rect 2947 9236 2993 9244
rect 3007 9236 3373 9244
rect 3387 9236 3473 9244
rect 3547 9236 4053 9244
rect 4067 9236 4273 9244
rect 4647 9236 4733 9244
rect 4927 9236 5093 9244
rect 5436 9244 5444 9273
rect 5476 9264 5484 9276
rect 5547 9276 5733 9284
rect 5747 9276 5813 9284
rect 6267 9276 6373 9284
rect 6587 9276 7073 9284
rect 7107 9276 7413 9284
rect 7427 9276 7553 9284
rect 7636 9284 7644 9296
rect 7727 9296 7753 9304
rect 7787 9296 8073 9304
rect 8287 9296 8673 9304
rect 9027 9296 9193 9304
rect 9667 9296 9813 9304
rect 10007 9296 10353 9304
rect 10867 9296 10953 9304
rect 11167 9296 11373 9304
rect 11387 9296 11393 9304
rect 11707 9296 11893 9304
rect 7636 9276 7853 9284
rect 8087 9276 8233 9284
rect 8667 9276 8973 9284
rect 10227 9276 10293 9284
rect 10307 9276 10313 9284
rect 10447 9276 10913 9284
rect 10927 9276 11093 9284
rect 11327 9276 11393 9284
rect 11507 9276 11693 9284
rect 11767 9276 11813 9284
rect 11867 9276 11973 9284
rect 12027 9276 12073 9284
rect 12127 9276 12173 9284
rect 5467 9256 5484 9264
rect 5507 9256 5673 9264
rect 6447 9256 6493 9264
rect 6507 9256 6733 9264
rect 6827 9256 6853 9264
rect 7187 9256 7353 9264
rect 7507 9256 7593 9264
rect 5436 9236 5453 9244
rect 5476 9236 6933 9244
rect 1887 9216 1993 9224
rect 2007 9216 2493 9224
rect 3487 9216 4113 9224
rect 5476 9224 5484 9236
rect 7167 9236 7233 9244
rect 7616 9244 7624 9273
rect 7687 9256 7913 9264
rect 8187 9256 8413 9264
rect 8656 9264 8664 9273
rect 8447 9256 8664 9264
rect 8967 9256 9013 9264
rect 9036 9264 9044 9273
rect 9036 9256 9253 9264
rect 9447 9256 9573 9264
rect 9627 9256 9713 9264
rect 10047 9256 10193 9264
rect 10287 9256 10373 9264
rect 10527 9256 10573 9264
rect 10627 9256 10653 9264
rect 11027 9256 11113 9264
rect 11136 9264 11144 9273
rect 11136 9256 11313 9264
rect 11567 9256 11733 9264
rect 11747 9256 11773 9264
rect 12007 9256 12153 9264
rect 7547 9236 7624 9244
rect 7867 9236 7953 9244
rect 8187 9236 8573 9244
rect 8876 9244 8884 9253
rect 8876 9236 9113 9244
rect 9427 9236 9513 9244
rect 9787 9236 9973 9244
rect 10467 9236 10533 9244
rect 10976 9244 10984 9253
rect 10967 9236 10984 9244
rect 11127 9236 11173 9244
rect 11527 9236 11633 9244
rect 12067 9236 12133 9244
rect 5127 9216 5484 9224
rect 5707 9216 5773 9224
rect 6227 9216 6313 9224
rect 6947 9216 7193 9224
rect 7747 9216 7873 9224
rect 7887 9216 8373 9224
rect 8847 9216 8913 9224
rect 9047 9216 9353 9224
rect 9587 9216 9973 9224
rect 10167 9216 10353 9224
rect 10367 9216 10933 9224
rect 10947 9216 11933 9224
rect 12107 9216 12173 9224
rect 5347 9196 5513 9204
rect 6587 9196 7313 9204
rect 7447 9196 7893 9204
rect 8467 9196 8873 9204
rect 8987 9196 9593 9204
rect 10147 9196 10433 9204
rect 10507 9196 10613 9204
rect 10767 9196 11793 9204
rect 1747 9176 3233 9184
rect 3387 9176 4253 9184
rect 4287 9176 5433 9184
rect 5467 9176 5613 9184
rect 5627 9176 5653 9184
rect 5667 9176 6133 9184
rect 6887 9176 8933 9184
rect 9267 9176 10553 9184
rect 10667 9176 10773 9184
rect 11147 9176 11213 9184
rect 1767 9156 5333 9164
rect 6787 9156 7273 9164
rect 7827 9156 8393 9164
rect 8447 9156 9453 9164
rect 10247 9156 11493 9164
rect 2147 9136 2633 9144
rect 3967 9136 5453 9144
rect 6127 9136 6153 9144
rect 6947 9136 7453 9144
rect 7887 9136 8553 9144
rect 9287 9136 9593 9144
rect 10047 9136 11313 9144
rect 1587 9116 2233 9124
rect 3007 9116 3113 9124
rect 3187 9116 6833 9124
rect 7467 9116 7633 9124
rect 7767 9116 10973 9124
rect 1567 9096 1793 9104
rect 1967 9096 2193 9104
rect 2967 9096 6633 9104
rect 6747 9096 7813 9104
rect 8007 9096 8464 9104
rect 8456 9087 8464 9096
rect 9547 9096 9693 9104
rect 9707 9096 10573 9104
rect 10607 9096 11033 9104
rect 1287 9076 1773 9084
rect 1787 9076 1853 9084
rect 2507 9076 2773 9084
rect 2787 9076 2953 9084
rect 2987 9076 6213 9084
rect 7087 9076 8433 9084
rect 8667 9076 8693 9084
rect 8727 9076 9553 9084
rect 9867 9076 10553 9084
rect 407 9056 1073 9064
rect 1747 9056 3513 9064
rect 4907 9056 5293 9064
rect 5316 9056 6013 9064
rect 547 9036 693 9044
rect 1087 9036 1833 9044
rect 3887 9036 4013 9044
rect 5316 9044 5324 9056
rect 7267 9056 7313 9064
rect 7407 9056 7473 9064
rect 7567 9056 7933 9064
rect 7956 9056 8284 9064
rect 5187 9036 5324 9044
rect 5447 9036 7173 9044
rect 7956 9044 7964 9056
rect 7267 9036 7964 9044
rect 7987 9036 8004 9044
rect 187 9016 253 9024
rect 667 9016 684 9024
rect 187 8996 233 9004
rect 127 8976 153 8984
rect 336 8984 344 8993
rect 207 8976 473 8984
rect 676 8967 684 9016
rect 847 9016 893 9024
rect 1607 9016 1733 9024
rect 2816 9016 2993 9024
rect 2816 9007 2824 9016
rect 3007 9016 3093 9024
rect 3947 9016 4053 9024
rect 4107 9016 4413 9024
rect 4547 9016 4833 9024
rect 4847 9016 4853 9024
rect 4867 9016 5113 9024
rect 5127 9016 5153 9024
rect 5467 9016 5573 9024
rect 6187 9016 6433 9024
rect 6447 9016 6773 9024
rect 6827 9016 6873 9024
rect 7007 9016 7293 9024
rect 7307 9016 7613 9024
rect 7767 9016 7953 9024
rect 7996 9024 8004 9036
rect 8027 9036 8053 9044
rect 8276 9044 8284 9056
rect 8307 9056 8693 9064
rect 9387 9056 10033 9064
rect 10387 9056 11013 9064
rect 8276 9036 8933 9044
rect 9887 9036 10713 9044
rect 11167 9036 11193 9044
rect 11247 9036 11253 9044
rect 11267 9036 11533 9044
rect 7996 9016 8064 9024
rect 907 8996 933 9004
rect 1687 8996 2173 9004
rect 2267 8996 2293 9004
rect 2427 8996 2473 9004
rect 3587 8996 3713 9004
rect 3747 8996 3813 9004
rect 3907 8996 3953 9004
rect 4087 8996 4373 9004
rect 4387 8996 4473 9004
rect 4887 8996 5033 9004
rect 5087 8996 5233 9004
rect 5416 8996 5773 9004
rect 1007 8976 1093 8984
rect 1387 8976 1513 8984
rect 1527 8976 1553 8984
rect 1567 8976 2404 8984
rect 2396 8967 2404 8976
rect 2447 8976 2493 8984
rect 2547 8976 2753 8984
rect 3107 8976 3193 8984
rect 4707 8976 5053 8984
rect 5236 8984 5244 8993
rect 5416 8987 5424 8996
rect 5796 8996 5973 9004
rect 5796 8987 5804 8996
rect 5236 8976 5373 8984
rect 5996 8967 6004 9013
rect 6467 8996 6653 9004
rect 6707 8996 6893 9004
rect 6907 8996 7033 9004
rect 7427 8996 7453 9004
rect 7587 8996 7933 9004
rect 7987 8996 8033 9004
rect 8056 9004 8064 9016
rect 8087 9016 8153 9024
rect 8767 9016 8853 9024
rect 8907 9016 8953 9024
rect 9007 9016 9073 9024
rect 9207 9016 9373 9024
rect 9387 9016 9613 9024
rect 9947 9016 10053 9024
rect 10567 9016 10704 9024
rect 8056 8996 8093 9004
rect 8247 8996 8533 9004
rect 8956 8996 8973 9004
rect 6087 8976 6353 8984
rect 6687 8976 6853 8984
rect 7247 8976 7393 8984
rect 7507 8976 7593 8984
rect 7647 8976 7773 8984
rect 7787 8976 7853 8984
rect 7927 8976 7993 8984
rect 8427 8976 8473 8984
rect 8587 8976 8673 8984
rect 8687 8976 8753 8984
rect 8956 8984 8964 8996
rect 9307 8996 9353 9004
rect 9727 8996 10093 9004
rect 10147 8996 10173 9004
rect 10316 8996 10473 9004
rect 10316 8987 10324 8996
rect 10527 8996 10573 9004
rect 10696 8987 10704 9016
rect 10787 9016 11173 9024
rect 11227 9016 11393 9024
rect 11407 9016 11573 9024
rect 11787 9016 11933 9024
rect 12027 9016 12113 9024
rect 10727 8996 11193 9004
rect 11327 8996 11373 9004
rect 11507 8996 11553 9004
rect 8827 8976 8964 8984
rect 8987 8976 9033 8984
rect 9087 8976 9213 8984
rect 9227 8976 9293 8984
rect 9316 8976 10093 8984
rect 507 8956 533 8964
rect 887 8956 1053 8964
rect 1187 8956 1253 8964
rect 1287 8956 1413 8964
rect 2407 8956 2653 8964
rect 3027 8956 3153 8964
rect 3607 8956 4573 8964
rect 5147 8956 5593 8964
rect 5607 8956 5753 8964
rect 6387 8956 6673 8964
rect 7087 8956 7213 8964
rect 7607 8956 7833 8964
rect 8147 8956 8173 8964
rect 8307 8956 8333 8964
rect 8427 8956 8793 8964
rect 9316 8964 9324 8976
rect 10107 8976 10153 8984
rect 10347 8976 10373 8984
rect 10387 8976 10453 8984
rect 10507 8976 10553 8984
rect 10607 8976 10653 8984
rect 10827 8976 10893 8984
rect 10907 8976 11053 8984
rect 11627 8976 11753 8984
rect 11907 8976 12033 8984
rect 8887 8956 9324 8964
rect 9887 8956 9953 8964
rect 10207 8956 10453 8964
rect 10847 8956 11013 8964
rect 11087 8956 11653 8964
rect 11827 8956 12033 8964
rect 12047 8956 12073 8964
rect 367 8936 653 8944
rect 667 8936 1573 8944
rect 2327 8936 2413 8944
rect 2487 8936 2593 8944
rect 2607 8936 3353 8944
rect 3427 8936 3753 8944
rect 4187 8936 5933 8944
rect 5967 8936 6173 8944
rect 6367 8936 8513 8944
rect 8907 8936 9153 8944
rect 9167 8936 9313 8944
rect 9327 8936 9393 8944
rect 9407 8936 9553 8944
rect 9627 8936 9893 8944
rect 10167 8936 11113 8944
rect 11447 8936 11593 8944
rect 11727 8936 11953 8944
rect 247 8916 693 8924
rect 947 8916 1393 8924
rect 1407 8916 1553 8924
rect 2287 8916 2973 8924
rect 5227 8916 5273 8924
rect 5287 8916 5713 8924
rect 5787 8916 5973 8924
rect 7067 8916 7873 8924
rect 7947 8916 9024 8924
rect 5047 8896 5133 8904
rect 5367 8896 5533 8904
rect 6547 8896 7133 8904
rect 7147 8896 7373 8904
rect 7527 8896 7653 8904
rect 7727 8896 7813 8904
rect 7887 8896 8153 8904
rect 8267 8896 8313 8904
rect 8636 8896 8713 8904
rect 927 8876 1433 8884
rect 1447 8876 1933 8884
rect 2347 8876 3413 8884
rect 4507 8876 5233 8884
rect 5247 8876 5573 8884
rect 5587 8876 6053 8884
rect 7387 8876 7553 8884
rect 8636 8884 8644 8896
rect 9016 8904 9024 8916
rect 9047 8916 9093 8924
rect 9107 8916 9733 8924
rect 10307 8916 10873 8924
rect 10927 8916 11333 8924
rect 11567 8916 11953 8924
rect 9016 8896 9253 8904
rect 9367 8896 9613 8904
rect 9907 8896 11733 8904
rect 11767 8896 11933 8904
rect 8007 8876 8644 8884
rect 8667 8876 9353 8884
rect 9567 8876 9673 8884
rect 9747 8876 10153 8884
rect 10287 8876 10393 8884
rect 10867 8876 10913 8884
rect 11167 8876 11433 8884
rect 11747 8876 11793 8884
rect 1767 8856 1813 8864
rect 3767 8856 4193 8864
rect 4447 8856 5013 8864
rect 6367 8856 6773 8864
rect 7447 8856 7533 8864
rect 7547 8856 7613 8864
rect 7627 8856 7633 8864
rect 7647 8856 8373 8864
rect 8947 8856 9573 8864
rect 10227 8856 10673 8864
rect 10907 8856 11233 8864
rect 11267 8856 11373 8864
rect 11587 8856 11793 8864
rect 807 8836 853 8844
rect 867 8836 1233 8844
rect 1547 8836 2253 8844
rect 3447 8836 3813 8844
rect 6047 8836 6753 8844
rect 7207 8836 7273 8844
rect 7287 8836 7333 8844
rect 7507 8836 7593 8844
rect 7667 8836 8933 8844
rect 9067 8836 9093 8844
rect 9107 8836 10273 8844
rect 10287 8836 11273 8844
rect 11627 8836 11773 8844
rect 11787 8836 11913 8844
rect 11927 8836 12113 8844
rect 167 8816 273 8824
rect 567 8816 753 8824
rect 767 8816 773 8824
rect 1067 8816 1173 8824
rect 1367 8816 1433 8824
rect 1807 8816 2033 8824
rect 2167 8816 2353 8824
rect 2367 8816 2873 8824
rect 3087 8816 3313 8824
rect 3327 8816 3753 8824
rect 3887 8816 3953 8824
rect 5827 8816 6033 8824
rect 6207 8816 6353 8824
rect 6707 8816 6793 8824
rect 6907 8816 7024 8824
rect 627 8796 633 8804
rect 647 8796 813 8804
rect 827 8796 873 8804
rect 896 8796 973 8804
rect 327 8776 493 8784
rect 507 8776 513 8784
rect 896 8784 904 8796
rect 1087 8796 1184 8804
rect 587 8776 904 8784
rect 927 8776 953 8784
rect 1127 8776 1153 8784
rect 1176 8784 1184 8796
rect 1227 8796 1393 8804
rect 1787 8796 1953 8804
rect 2527 8796 2833 8804
rect 2867 8796 2893 8804
rect 2967 8796 2993 8804
rect 3207 8796 3273 8804
rect 3487 8796 3593 8804
rect 3616 8796 3724 8804
rect 1176 8776 1193 8784
rect 1247 8776 1333 8784
rect 1596 8784 1604 8793
rect 1567 8776 1604 8784
rect 1736 8784 1744 8793
rect 1736 8776 1893 8784
rect 2336 8784 2344 8793
rect 2027 8776 2453 8784
rect 2547 8776 2613 8784
rect 2767 8776 3193 8784
rect 3247 8776 3493 8784
rect 3616 8784 3624 8796
rect 3547 8776 3624 8784
rect 3667 8776 3693 8784
rect 3716 8784 3724 8796
rect 3787 8796 3853 8804
rect 3887 8796 4053 8804
rect 4067 8796 4153 8804
rect 4247 8796 4333 8804
rect 4356 8796 4953 8804
rect 3716 8776 3873 8784
rect 4356 8784 4364 8796
rect 5267 8796 5353 8804
rect 5407 8796 5473 8804
rect 5767 8796 5813 8804
rect 5907 8796 5953 8804
rect 6076 8796 6153 8804
rect 4267 8776 4364 8784
rect 4867 8776 4893 8784
rect 5327 8776 5373 8784
rect 5427 8776 5513 8784
rect 5587 8776 5733 8784
rect 6076 8784 6084 8796
rect 6207 8796 6393 8804
rect 6487 8796 6533 8804
rect 7016 8804 7024 8816
rect 7047 8816 7733 8824
rect 8127 8816 8233 8824
rect 8287 8816 8313 8824
rect 8467 8816 8533 8824
rect 8547 8816 8653 8824
rect 8827 8816 8853 8824
rect 9687 8816 9793 8824
rect 9827 8816 9993 8824
rect 10687 8816 10753 8824
rect 11287 8816 11453 8824
rect 11547 8816 11633 8824
rect 11727 8816 12133 8824
rect 6727 8796 6884 8804
rect 7016 8796 7193 8804
rect 6876 8787 6884 8796
rect 7227 8796 7273 8804
rect 7467 8796 7573 8804
rect 7587 8796 7653 8804
rect 7987 8796 8164 8804
rect 8156 8787 8164 8796
rect 8407 8796 8493 8804
rect 8647 8796 8853 8804
rect 8967 8796 9053 8804
rect 9127 8796 9233 8804
rect 9247 8796 9313 8804
rect 9356 8796 9433 8804
rect 5947 8776 6084 8784
rect 6107 8776 6133 8784
rect 6187 8776 6373 8784
rect 7687 8776 7733 8784
rect 8247 8776 8653 8784
rect 8847 8776 8973 8784
rect 8987 8776 8993 8784
rect 9356 8784 9364 8796
rect 9447 8796 9633 8804
rect 9647 8796 9913 8804
rect 10027 8796 10213 8804
rect 11027 8796 11073 8804
rect 11096 8804 11104 8813
rect 11096 8796 11293 8804
rect 11487 8796 11573 8804
rect 11667 8796 11753 8804
rect 11827 8796 11964 8804
rect 11956 8787 11964 8796
rect 11987 8796 12053 8804
rect 12067 8796 12153 8804
rect 9087 8776 9364 8784
rect 9387 8776 9453 8784
rect 9607 8776 9693 8784
rect 10056 8776 10173 8784
rect 267 8756 293 8764
rect 316 8756 333 8764
rect 316 8744 324 8756
rect 887 8756 1753 8764
rect 1947 8756 2693 8764
rect 2747 8756 2824 8764
rect 147 8736 324 8744
rect 1707 8736 1953 8744
rect 2587 8736 2713 8744
rect 2816 8744 2824 8756
rect 2847 8756 2913 8764
rect 3647 8756 3973 8764
rect 4127 8756 4313 8764
rect 4787 8756 6584 8764
rect 2816 8736 3093 8744
rect 3547 8736 3713 8744
rect 3727 8736 4773 8744
rect 4967 8736 5053 8744
rect 5067 8736 5833 8744
rect 5927 8736 5953 8744
rect 5987 8736 6113 8744
rect 6127 8736 6513 8744
rect 6527 8736 6553 8744
rect 6576 8744 6584 8756
rect 6887 8756 6993 8764
rect 8147 8756 8213 8764
rect 8627 8756 8733 8764
rect 8887 8756 9413 8764
rect 10056 8764 10064 8776
rect 10187 8776 10353 8784
rect 10427 8776 10513 8784
rect 10847 8776 10933 8784
rect 11227 8776 11253 8784
rect 11267 8776 11413 8784
rect 11967 8776 11993 8784
rect 12107 8776 12133 8784
rect 9587 8756 10064 8764
rect 10107 8756 10193 8764
rect 10607 8756 10773 8764
rect 10807 8756 11073 8764
rect 11827 8756 11873 8764
rect 6576 8736 8133 8744
rect 9047 8736 9813 8744
rect 9827 8736 10333 8744
rect 10567 8736 11453 8744
rect 11467 8736 11553 8744
rect 3467 8716 3833 8724
rect 3847 8716 4213 8724
rect 4227 8716 5713 8724
rect 5727 8716 8593 8724
rect 8607 8716 8793 8724
rect 8807 8716 10233 8724
rect 10447 8716 10793 8724
rect 3667 8696 3693 8704
rect 4747 8696 5173 8704
rect 5187 8696 5793 8704
rect 5827 8696 7013 8704
rect 7387 8696 10933 8704
rect 10947 8696 10953 8704
rect 3347 8676 4033 8684
rect 4047 8676 7913 8684
rect 8027 8676 9173 8684
rect 9267 8676 10693 8684
rect 3067 8656 4093 8664
rect 7667 8656 7693 8664
rect 7707 8656 8233 8664
rect 8507 8656 8533 8664
rect 8647 8656 9313 8664
rect 9336 8656 10433 8664
rect 1327 8636 1633 8644
rect 2867 8636 4173 8644
rect 4427 8636 6364 8644
rect 1047 8616 2693 8624
rect 3007 8616 4593 8624
rect 4887 8616 5053 8624
rect 6356 8624 6364 8636
rect 6387 8636 6673 8644
rect 6687 8636 7193 8644
rect 8187 8636 8373 8644
rect 8687 8636 9113 8644
rect 9336 8644 9344 8656
rect 10447 8656 11713 8664
rect 9127 8636 9344 8644
rect 9367 8636 10593 8644
rect 10627 8636 10873 8644
rect 10987 8636 11653 8644
rect 6356 8616 6813 8624
rect 6867 8616 9453 8624
rect 9507 8616 9573 8624
rect 9587 8616 11033 8624
rect 11787 8616 11893 8624
rect 1427 8596 1653 8604
rect 3687 8596 3773 8604
rect 3787 8596 4553 8604
rect 4727 8596 6073 8604
rect 6427 8596 6633 8604
rect 6647 8596 6833 8604
rect 6847 8596 7393 8604
rect 7707 8596 7913 8604
rect 8207 8596 8313 8604
rect 8367 8596 9073 8604
rect 9387 8596 10213 8604
rect 11527 8596 11633 8604
rect 1507 8576 1573 8584
rect 1647 8576 3144 8584
rect 127 8556 233 8564
rect 1247 8556 1593 8564
rect 1627 8556 2813 8564
rect 3136 8564 3144 8576
rect 3167 8576 4033 8584
rect 4067 8576 5873 8584
rect 5887 8576 6313 8584
rect 6327 8576 7233 8584
rect 7567 8576 9013 8584
rect 9067 8576 9373 8584
rect 9847 8576 9873 8584
rect 10896 8576 11533 8584
rect 2927 8556 2964 8564
rect 3136 8556 3473 8564
rect 2956 8547 2964 8556
rect 4387 8556 4613 8564
rect 4627 8556 4973 8564
rect 5087 8556 5253 8564
rect 5267 8556 5553 8564
rect 5967 8556 6273 8564
rect 6347 8556 6573 8564
rect 6827 8556 8133 8564
rect 8167 8556 8513 8564
rect 8176 8547 8184 8556
rect 8747 8556 8933 8564
rect 9047 8556 9133 8564
rect 9887 8556 9933 8564
rect 10896 8564 10904 8576
rect 10227 8556 10904 8564
rect 10927 8556 10993 8564
rect 11407 8556 11433 8564
rect 11927 8556 11973 8564
rect 167 8536 673 8544
rect 1107 8536 1173 8544
rect 1367 8536 1833 8544
rect 1987 8536 2024 8544
rect 147 8516 313 8524
rect 527 8516 653 8524
rect 707 8516 724 8524
rect 287 8496 493 8504
rect 547 8496 593 8504
rect 607 8496 693 8504
rect 716 8504 724 8516
rect 1056 8524 1064 8533
rect 1047 8516 1064 8524
rect 1087 8516 1193 8524
rect 1507 8516 1553 8524
rect 1707 8516 1753 8524
rect 1767 8516 1853 8524
rect 1927 8516 1993 8524
rect 716 8496 853 8504
rect 907 8496 1433 8504
rect 1447 8496 1473 8504
rect 1607 8496 1673 8504
rect 1947 8496 1973 8504
rect 2016 8504 2024 8536
rect 2387 8536 2913 8544
rect 3567 8536 3693 8544
rect 3747 8536 3853 8544
rect 4327 8536 5113 8544
rect 5167 8536 5393 8544
rect 5487 8536 6344 8544
rect 2047 8516 2193 8524
rect 2427 8516 2493 8524
rect 2507 8516 2924 8524
rect 1996 8496 2024 8504
rect 1996 8487 2004 8496
rect 2047 8496 2213 8504
rect 2247 8496 2513 8504
rect 2527 8496 2533 8504
rect 2707 8496 2773 8504
rect 2787 8496 2853 8504
rect 2916 8504 2924 8516
rect 2947 8516 2993 8524
rect 3047 8516 3153 8524
rect 3516 8516 4453 8524
rect 2916 8496 3113 8504
rect 3516 8504 3524 8516
rect 4647 8516 5084 8524
rect 3467 8496 3524 8504
rect 3807 8496 3913 8504
rect 4047 8496 4053 8504
rect 4067 8496 4713 8504
rect 4727 8496 4753 8504
rect 4827 8496 4893 8504
rect 4927 8496 5033 8504
rect 5076 8504 5084 8516
rect 5107 8516 5193 8524
rect 5247 8516 5413 8524
rect 5527 8516 5573 8524
rect 6067 8516 6164 8524
rect 6156 8507 6164 8516
rect 6187 8516 6313 8524
rect 6336 8524 6344 8536
rect 7127 8536 7413 8544
rect 7487 8536 7753 8544
rect 8027 8536 8164 8544
rect 8156 8527 8164 8536
rect 8227 8536 8353 8544
rect 8487 8536 8533 8544
rect 8556 8527 8564 8553
rect 8767 8536 8893 8544
rect 9707 8536 9864 8544
rect 6336 8516 6713 8524
rect 6827 8516 6873 8524
rect 7407 8516 7573 8524
rect 7596 8516 7613 8524
rect 5076 8496 5213 8504
rect 5787 8496 5893 8504
rect 5907 8496 6113 8504
rect 6527 8496 6693 8504
rect 6747 8496 6893 8504
rect 7207 8496 7253 8504
rect 7267 8496 7433 8504
rect 7596 8504 7604 8516
rect 7807 8516 7933 8524
rect 8587 8516 8864 8524
rect 7487 8496 7604 8504
rect 7867 8496 7973 8504
rect 8147 8496 8473 8504
rect 8527 8496 8773 8504
rect 8787 8496 8813 8504
rect 8856 8504 8864 8516
rect 8887 8516 8933 8524
rect 8987 8516 9053 8524
rect 9156 8516 9333 8524
rect 8856 8496 8953 8504
rect 9156 8504 9164 8516
rect 9856 8524 9864 8536
rect 10847 8536 11133 8544
rect 11156 8536 11233 8544
rect 11156 8527 11164 8536
rect 11247 8536 11313 8544
rect 11747 8536 11793 8544
rect 11867 8536 11933 8544
rect 11947 8536 12113 8544
rect 9856 8516 9933 8524
rect 9987 8516 10064 8524
rect 8996 8496 9164 8504
rect 347 8476 573 8484
rect 847 8476 873 8484
rect 1307 8476 1453 8484
rect 1707 8476 1813 8484
rect 2187 8476 2333 8484
rect 2347 8476 2553 8484
rect 2987 8476 3013 8484
rect 3027 8476 3193 8484
rect 3767 8476 4033 8484
rect 4056 8476 4433 8484
rect 167 8456 213 8464
rect 487 8456 1213 8464
rect 1867 8456 2013 8464
rect 4056 8464 4064 8476
rect 4467 8476 4813 8484
rect 4887 8476 7453 8484
rect 7467 8476 7513 8484
rect 7527 8476 7613 8484
rect 7687 8476 7773 8484
rect 7847 8476 8024 8484
rect 2687 8456 4064 8464
rect 4087 8456 4213 8464
rect 4747 8456 4793 8464
rect 4927 8456 4993 8464
rect 5067 8456 5733 8464
rect 6247 8456 6913 8464
rect 7127 8456 7253 8464
rect 7447 8456 7493 8464
rect 7747 8456 7993 8464
rect 8016 8464 8024 8476
rect 8047 8476 8193 8484
rect 8216 8476 8273 8484
rect 8016 8456 8033 8464
rect 8216 8464 8224 8476
rect 8996 8484 9004 8496
rect 9187 8496 9513 8504
rect 9667 8496 10033 8504
rect 10056 8504 10064 8516
rect 10087 8516 10113 8524
rect 10427 8516 10453 8524
rect 11427 8516 11513 8524
rect 11696 8516 12033 8524
rect 11696 8507 11704 8516
rect 10056 8496 10253 8504
rect 10847 8496 10993 8504
rect 11047 8496 11313 8504
rect 11367 8496 11493 8504
rect 11747 8496 11773 8504
rect 11887 8496 11953 8504
rect 8407 8476 9004 8484
rect 9027 8476 9113 8484
rect 9127 8476 9233 8484
rect 9687 8476 10073 8484
rect 10087 8476 10113 8484
rect 10127 8476 10153 8484
rect 10827 8476 11253 8484
rect 11267 8476 11353 8484
rect 11867 8476 12073 8484
rect 8207 8456 8224 8464
rect 8247 8456 8533 8464
rect 8587 8456 8593 8464
rect 8607 8456 9153 8464
rect 9227 8456 9793 8464
rect 10107 8456 10313 8464
rect 10327 8456 10333 8464
rect 10487 8456 10633 8464
rect 10707 8456 10973 8464
rect 11127 8456 11293 8464
rect 787 8436 1253 8444
rect 1467 8436 2353 8444
rect 2607 8436 2933 8444
rect 3007 8436 3173 8444
rect 3187 8436 3513 8444
rect 3527 8436 3833 8444
rect 3847 8436 4873 8444
rect 4907 8436 5173 8444
rect 5467 8436 5753 8444
rect 5847 8436 6513 8444
rect 6767 8436 6873 8444
rect 6967 8436 7733 8444
rect 7767 8436 7873 8444
rect 7907 8436 8413 8444
rect 9467 8436 9573 8444
rect 10247 8436 10693 8444
rect 10727 8436 10953 8444
rect 10967 8436 11113 8444
rect 11507 8436 12013 8444
rect 187 8416 233 8424
rect 247 8416 733 8424
rect 747 8416 793 8424
rect 1687 8416 1733 8424
rect 2667 8416 4893 8424
rect 4967 8416 5153 8424
rect 5507 8416 5933 8424
rect 5956 8416 6353 8424
rect 1227 8396 3333 8404
rect 3756 8396 3933 8404
rect 1587 8376 1653 8384
rect 2247 8376 2393 8384
rect 2627 8376 2833 8384
rect 3756 8384 3764 8396
rect 5956 8404 5964 8416
rect 7587 8416 10673 8424
rect 10827 8416 11713 8424
rect 5187 8396 5964 8404
rect 5987 8396 6493 8404
rect 6516 8396 6953 8404
rect 3187 8376 3764 8384
rect 3776 8376 4513 8384
rect 427 8356 633 8364
rect 1727 8356 1773 8364
rect 1787 8356 2173 8364
rect 2767 8356 2793 8364
rect 3776 8364 3784 8376
rect 5547 8376 5953 8384
rect 6516 8384 6524 8396
rect 7267 8396 7893 8404
rect 7967 8396 8473 8404
rect 8487 8396 9473 8404
rect 9487 8396 10193 8404
rect 11147 8396 11213 8404
rect 11687 8396 11913 8404
rect 6367 8376 6524 8384
rect 6627 8376 7273 8384
rect 7287 8376 7393 8384
rect 7667 8376 7713 8384
rect 7727 8376 7773 8384
rect 7787 8376 9293 8384
rect 9387 8376 10073 8384
rect 10987 8376 11593 8384
rect 3547 8356 3784 8364
rect 3967 8356 4073 8364
rect 5847 8356 5973 8364
rect 6267 8356 7133 8364
rect 7147 8356 7373 8364
rect 7827 8356 7853 8364
rect 7867 8356 8333 8364
rect 8567 8356 8613 8364
rect 8747 8356 8893 8364
rect 9307 8356 9713 8364
rect 10247 8356 10293 8364
rect 11387 8356 11453 8364
rect 327 8336 784 8344
rect 207 8316 313 8324
rect 367 8316 573 8324
rect 776 8324 784 8336
rect 1027 8336 1113 8344
rect 1207 8336 1233 8344
rect 1247 8336 1273 8344
rect 1356 8336 1593 8344
rect 1356 8324 1364 8336
rect 1767 8336 2193 8344
rect 2307 8336 2373 8344
rect 2387 8336 2593 8344
rect 2747 8336 2973 8344
rect 3307 8336 3373 8344
rect 3427 8336 3753 8344
rect 3827 8336 4004 8344
rect 776 8316 1364 8324
rect 1376 8316 1433 8324
rect 607 8296 753 8304
rect 767 8296 993 8304
rect 1376 8304 1384 8316
rect 1447 8316 1453 8324
rect 1467 8316 1553 8324
rect 1747 8316 1813 8324
rect 1947 8316 2173 8324
rect 2187 8316 2553 8324
rect 2567 8316 2653 8324
rect 2796 8316 2813 8324
rect 2796 8307 2804 8316
rect 2967 8316 3033 8324
rect 3047 8316 3484 8324
rect 1187 8296 1384 8304
rect 1627 8296 1693 8304
rect 1767 8296 1793 8304
rect 2327 8296 2353 8304
rect 2627 8296 2693 8304
rect 3476 8304 3484 8316
rect 3507 8316 3553 8324
rect 3587 8316 3873 8324
rect 3996 8324 4004 8336
rect 4027 8336 4153 8344
rect 4167 8336 4213 8344
rect 4267 8336 5913 8344
rect 5936 8336 5993 8344
rect 3996 8316 4193 8324
rect 4247 8316 4313 8324
rect 4587 8316 4673 8324
rect 4687 8316 5093 8324
rect 5107 8316 5313 8324
rect 5936 8324 5944 8336
rect 6007 8336 6193 8344
rect 6547 8336 6753 8344
rect 6867 8336 6913 8344
rect 6927 8336 6933 8344
rect 7427 8336 7953 8344
rect 8087 8336 8173 8344
rect 8267 8336 8373 8344
rect 8607 8336 8693 8344
rect 8787 8336 8833 8344
rect 8867 8336 8913 8344
rect 9567 8336 9613 8344
rect 10087 8336 10244 8344
rect 5867 8316 5944 8324
rect 6187 8316 6344 8324
rect 3167 8296 3464 8304
rect 3476 8296 3533 8304
rect 167 8276 373 8284
rect 387 8276 773 8284
rect 827 8276 973 8284
rect 987 8276 1253 8284
rect 1407 8276 1573 8284
rect 1587 8276 1733 8284
rect 1827 8276 1893 8284
rect 1927 8276 2233 8284
rect 2247 8276 2573 8284
rect 2587 8276 3293 8284
rect 3456 8284 3464 8296
rect 4087 8296 4133 8304
rect 4227 8296 4293 8304
rect 4367 8296 4493 8304
rect 4547 8296 4693 8304
rect 4747 8296 5053 8304
rect 5067 8296 5233 8304
rect 5527 8296 5613 8304
rect 6227 8296 6253 8304
rect 6336 8304 6344 8316
rect 6407 8316 6493 8324
rect 6567 8316 6613 8324
rect 6787 8316 7093 8324
rect 7327 8316 7353 8324
rect 7487 8316 8084 8324
rect 6336 8296 6373 8304
rect 6547 8296 6573 8304
rect 7047 8296 7473 8304
rect 7747 8296 7873 8304
rect 7896 8296 8053 8304
rect 7896 8287 7904 8296
rect 8076 8304 8084 8316
rect 8407 8316 8504 8324
rect 8496 8307 8504 8316
rect 8667 8316 8833 8324
rect 8967 8316 9033 8324
rect 9367 8316 9393 8324
rect 9447 8316 9693 8324
rect 9727 8316 10213 8324
rect 10236 8324 10244 8336
rect 10267 8336 10313 8344
rect 10996 8336 11013 8344
rect 10236 8316 10673 8324
rect 10687 8316 10813 8324
rect 10847 8316 10893 8324
rect 10907 8316 10973 8324
rect 10996 8307 11004 8336
rect 11067 8336 11093 8344
rect 11167 8336 11393 8344
rect 11407 8336 11413 8344
rect 11427 8336 11673 8344
rect 11727 8336 11753 8344
rect 11927 8336 11953 8344
rect 12087 8336 12113 8344
rect 11027 8316 11053 8324
rect 11127 8316 11413 8324
rect 11427 8316 11493 8324
rect 11787 8316 11893 8324
rect 11947 8316 12093 8324
rect 8076 8296 8093 8304
rect 8547 8296 8913 8304
rect 9007 8296 9033 8304
rect 9056 8296 9333 8304
rect 3456 8276 3493 8284
rect 3727 8276 3773 8284
rect 4407 8276 4473 8284
rect 4607 8276 5773 8284
rect 5807 8276 6073 8284
rect 6427 8276 6813 8284
rect 6827 8276 7053 8284
rect 7127 8276 7273 8284
rect 7387 8276 7793 8284
rect 8307 8276 8433 8284
rect 8456 8284 8464 8293
rect 9056 8287 9064 8296
rect 9347 8296 9373 8304
rect 9387 8296 9513 8304
rect 9696 8296 9733 8304
rect 8456 8276 8613 8284
rect 9696 8284 9704 8296
rect 10507 8296 10633 8304
rect 11047 8296 11113 8304
rect 11127 8296 11213 8304
rect 11927 8296 11953 8304
rect 9267 8276 9704 8284
rect 9727 8276 10113 8284
rect 10227 8276 10433 8284
rect 10487 8276 10853 8284
rect 10927 8276 11193 8284
rect 667 8256 1213 8264
rect 1227 8256 1353 8264
rect 2027 8256 2433 8264
rect 2667 8256 3853 8264
rect 3887 8256 4213 8264
rect 4796 8256 7373 8264
rect 887 8236 1013 8244
rect 1027 8236 2053 8244
rect 4796 8244 4804 8256
rect 7467 8256 7573 8264
rect 8247 8256 8413 8264
rect 9747 8256 9833 8264
rect 9867 8256 9953 8264
rect 9967 8256 10233 8264
rect 10527 8256 10613 8264
rect 10627 8256 11013 8264
rect 11027 8256 11153 8264
rect 11207 8256 11733 8264
rect 11747 8256 11853 8264
rect 2367 8236 4804 8244
rect 5127 8236 5613 8244
rect 5996 8236 6593 8244
rect 2467 8216 2553 8224
rect 2607 8216 2733 8224
rect 2787 8216 2853 8224
rect 2887 8216 2993 8224
rect 3167 8216 3813 8224
rect 3967 8216 4053 8224
rect 4187 8216 5093 8224
rect 5996 8224 6004 8236
rect 6987 8236 7013 8244
rect 7427 8236 7493 8244
rect 7507 8236 7713 8244
rect 8627 8236 9253 8244
rect 9507 8236 9753 8244
rect 9767 8236 10053 8244
rect 10067 8236 11193 8244
rect 11207 8236 11873 8244
rect 5107 8216 6004 8224
rect 6047 8216 7113 8224
rect 7187 8216 8013 8224
rect 8867 8216 9653 8224
rect 9767 8216 9813 8224
rect 10847 8216 11233 8224
rect 11247 8216 11333 8224
rect 2527 8196 2973 8204
rect 3407 8196 3753 8204
rect 3927 8196 4133 8204
rect 4987 8196 5133 8204
rect 5147 8196 5353 8204
rect 5587 8196 6933 8204
rect 7147 8196 8413 8204
rect 9027 8196 9073 8204
rect 9087 8196 9133 8204
rect 9427 8196 9453 8204
rect 9467 8196 10553 8204
rect 11327 8196 12033 8204
rect 1547 8176 2413 8184
rect 2467 8176 3453 8184
rect 3547 8176 3733 8184
rect 3767 8176 6473 8184
rect 6587 8176 6793 8184
rect 7747 8176 7793 8184
rect 8427 8176 9673 8184
rect 9707 8176 10393 8184
rect 10407 8176 10913 8184
rect 1147 8156 1753 8164
rect 2507 8156 2613 8164
rect 2667 8156 3153 8164
rect 3327 8156 3373 8164
rect 3527 8156 3533 8164
rect 3747 8156 7633 8164
rect 7647 8156 7653 8164
rect 8787 8156 11313 8164
rect 707 8136 853 8144
rect 1707 8136 1833 8144
rect 1847 8136 2073 8144
rect 2407 8136 3133 8144
rect 3167 8136 3413 8144
rect 3547 8136 3593 8144
rect 3727 8136 3953 8144
rect 4907 8136 5513 8144
rect 5787 8136 6273 8144
rect 6387 8136 6413 8144
rect 6467 8136 7293 8144
rect 7407 8136 7633 8144
rect 7727 8136 9173 8144
rect 9827 8136 9913 8144
rect 9927 8136 11713 8144
rect 1947 8116 1993 8124
rect 2027 8116 2093 8124
rect 2127 8116 2653 8124
rect 2747 8116 4273 8124
rect 4427 8116 5193 8124
rect 5347 8116 6633 8124
rect 6827 8116 7193 8124
rect 7207 8116 10533 8124
rect 10547 8116 10593 8124
rect 11127 8116 11213 8124
rect 1747 8096 2013 8104
rect 2027 8096 2453 8104
rect 2527 8096 4544 8104
rect 147 8076 253 8084
rect 347 8076 1393 8084
rect 1667 8076 2673 8084
rect 2707 8076 2913 8084
rect 3207 8076 4093 8084
rect 4247 8076 4313 8084
rect 4536 8084 4544 8096
rect 4567 8096 4593 8104
rect 5007 8096 5153 8104
rect 5287 8096 5393 8104
rect 5427 8096 6113 8104
rect 6127 8096 6753 8104
rect 7207 8096 7753 8104
rect 7947 8096 8153 8104
rect 8227 8096 8893 8104
rect 9267 8096 9493 8104
rect 9807 8096 9973 8104
rect 10247 8096 10373 8104
rect 10387 8096 10833 8104
rect 11147 8096 11233 8104
rect 11687 8096 11853 8104
rect 11867 8096 11873 8104
rect 4536 8076 4944 8084
rect 187 8056 233 8064
rect 407 8056 693 8064
rect 1187 8056 1493 8064
rect 1507 8056 1793 8064
rect 1927 8056 1953 8064
rect 2487 8056 2593 8064
rect 2687 8056 2764 8064
rect 207 8036 213 8044
rect 227 8036 333 8044
rect 987 8036 1033 8044
rect 1107 8036 1133 8044
rect 1427 8036 1533 8044
rect 1547 8036 2113 8044
rect 2147 8036 2304 8044
rect 936 8016 1053 8024
rect 367 7996 393 8004
rect 407 7996 413 8004
rect 936 8004 944 8016
rect 1336 8024 1344 8033
rect 2296 8027 2304 8036
rect 2427 8036 2493 8044
rect 2667 8036 2733 8044
rect 2756 8044 2764 8056
rect 2807 8056 2833 8064
rect 2856 8056 3033 8064
rect 2856 8044 2864 8056
rect 3047 8056 3633 8064
rect 3907 8056 3944 8064
rect 2756 8036 2864 8044
rect 2907 8036 3013 8044
rect 3227 8036 3353 8044
rect 3936 8044 3944 8056
rect 4527 8056 4753 8064
rect 4767 8056 4893 8064
rect 4936 8064 4944 8076
rect 4967 8076 5073 8084
rect 5216 8076 5573 8084
rect 5216 8064 5224 8076
rect 5627 8076 5933 8084
rect 6167 8076 6453 8084
rect 7167 8076 7204 8084
rect 4936 8056 5224 8064
rect 5247 8056 5373 8064
rect 5667 8056 5853 8064
rect 5867 8056 6093 8064
rect 6207 8056 6333 8064
rect 6427 8056 6493 8064
rect 6607 8056 6693 8064
rect 7196 8064 7204 8076
rect 7767 8076 7833 8084
rect 8327 8076 8713 8084
rect 8787 8076 8813 8084
rect 9787 8076 10413 8084
rect 11107 8076 11333 8084
rect 7196 8056 7733 8064
rect 7747 8056 7853 8064
rect 8107 8056 8533 8064
rect 8587 8056 8853 8064
rect 9067 8056 9573 8064
rect 9636 8056 9773 8064
rect 3936 8036 4073 8044
rect 4207 8036 4833 8044
rect 4867 8036 4933 8044
rect 5436 8044 5444 8053
rect 9636 8047 9644 8056
rect 9807 8056 9853 8064
rect 9867 8056 10353 8064
rect 10367 8056 10613 8064
rect 10647 8056 10793 8064
rect 10807 8056 10993 8064
rect 11107 8056 11153 8064
rect 11587 8056 11693 8064
rect 11707 8056 12013 8064
rect 5287 8036 5444 8044
rect 5507 8036 5613 8044
rect 5807 8036 5833 8044
rect 5856 8036 6053 8044
rect 1207 8016 1473 8024
rect 1527 8016 1573 8024
rect 1816 8016 1873 8024
rect 567 7996 944 8004
rect 967 7996 1093 8004
rect 1367 7996 1773 8004
rect 1816 8004 1824 8016
rect 1947 8016 1993 8024
rect 2667 8016 3804 8024
rect 1787 7996 1824 8004
rect 1847 7996 2093 8004
rect 2247 7996 2253 8004
rect 2267 7996 2893 8004
rect 3367 7996 3673 8004
rect 3796 8004 3804 8016
rect 3887 8016 4013 8024
rect 4047 8016 4093 8024
rect 5067 8016 5453 8024
rect 5467 8016 5593 8024
rect 5856 8024 5864 8036
rect 6067 8036 6373 8044
rect 6447 8036 6813 8044
rect 7676 8036 7944 8044
rect 5787 8016 5864 8024
rect 6087 8016 6153 8024
rect 6196 8016 6413 8024
rect 3796 7996 3953 8004
rect 3967 7996 4193 8004
rect 4747 7996 5253 8004
rect 5356 7996 5593 8004
rect 787 7976 1813 7984
rect 1827 7976 2513 7984
rect 2676 7976 3493 7984
rect 1167 7956 1353 7964
rect 1847 7956 2033 7964
rect 2676 7964 2684 7976
rect 3687 7976 3753 7984
rect 3847 7976 3893 7984
rect 5356 7984 5364 7996
rect 5627 7996 6033 8004
rect 6196 8004 6204 8016
rect 6467 8016 6533 8024
rect 6627 8016 6753 8024
rect 6807 8016 6953 8024
rect 7676 8024 7684 8036
rect 7227 8016 7684 8024
rect 7707 8016 7873 8024
rect 7936 8024 7944 8036
rect 7967 8036 8073 8044
rect 8127 8036 8433 8044
rect 8787 8036 8813 8044
rect 8907 8036 9004 8044
rect 7936 8016 8193 8024
rect 8207 8016 8273 8024
rect 8427 8016 8833 8024
rect 8887 8016 8933 8024
rect 8996 8024 9004 8036
rect 9027 8036 9513 8044
rect 9687 8036 9773 8044
rect 9787 8036 9833 8044
rect 10167 8036 10193 8044
rect 10227 8036 10373 8044
rect 10387 8036 10553 8044
rect 11027 8036 11113 8044
rect 11287 8036 11584 8044
rect 11576 8027 11584 8036
rect 11667 8036 11713 8044
rect 8996 8016 9033 8024
rect 9187 8016 9213 8024
rect 9427 8016 9613 8024
rect 9627 8016 9793 8024
rect 9927 8016 10224 8024
rect 10216 8007 10224 8016
rect 10627 8016 10713 8024
rect 10787 8016 10953 8024
rect 11187 8016 11353 8024
rect 11467 8016 11533 8024
rect 11647 8016 12093 8024
rect 6087 7996 6204 8004
rect 6227 7996 6433 8004
rect 6947 7996 6973 8004
rect 7007 7996 7133 8004
rect 7207 7996 7353 8004
rect 7407 7996 7453 8004
rect 7467 7996 7533 8004
rect 7947 7996 8193 8004
rect 8207 7996 8804 8004
rect 4027 7976 5364 7984
rect 5387 7976 5633 7984
rect 5756 7976 5953 7984
rect 2067 7956 2684 7964
rect 2867 7956 3513 7964
rect 3667 7956 4113 7964
rect 4167 7956 4513 7964
rect 5327 7956 5473 7964
rect 5756 7964 5764 7976
rect 5987 7976 6013 7984
rect 6267 7976 6833 7984
rect 6847 7976 7693 7984
rect 7847 7976 7893 7984
rect 7947 7976 8573 7984
rect 8796 7984 8804 7996
rect 8947 7996 9073 8004
rect 9207 7996 9273 8004
rect 10067 7996 10173 8004
rect 10247 7996 10313 8004
rect 11147 7996 11193 8004
rect 11387 7996 11893 8004
rect 8796 7976 8893 7984
rect 9287 7976 9433 7984
rect 9947 7976 10633 7984
rect 11007 7976 11273 7984
rect 11527 7976 11553 7984
rect 5647 7956 5764 7964
rect 5927 7956 7153 7964
rect 7507 7956 7573 7964
rect 8827 7956 10093 7964
rect 10587 7956 10633 7964
rect 11187 7956 11213 7964
rect 1827 7936 4673 7944
rect 4727 7936 5144 7944
rect 747 7916 1053 7924
rect 1407 7916 1993 7924
rect 2007 7916 2073 7924
rect 2127 7916 2213 7924
rect 3387 7916 3433 7924
rect 3487 7916 3873 7924
rect 3887 7916 4053 7924
rect 4067 7916 4153 7924
rect 4747 7916 4873 7924
rect 4887 7916 5013 7924
rect 5136 7924 5144 7936
rect 5807 7936 5873 7944
rect 6276 7936 6673 7944
rect 5136 7916 5273 7924
rect 5367 7916 5613 7924
rect 6276 7924 6284 7936
rect 7027 7936 7753 7944
rect 7887 7936 7953 7944
rect 7967 7936 8053 7944
rect 8307 7936 8393 7944
rect 8407 7936 8873 7944
rect 8927 7936 9173 7944
rect 9207 7936 10933 7944
rect 5947 7916 6284 7924
rect 6307 7916 7173 7924
rect 7347 7916 7713 7924
rect 7847 7916 8093 7924
rect 8687 7916 8813 7924
rect 8867 7916 9633 7924
rect 10007 7916 12133 7924
rect 847 7896 1693 7904
rect 1767 7896 2833 7904
rect 3247 7896 3393 7904
rect 3747 7896 3853 7904
rect 3947 7896 4164 7904
rect 407 7876 573 7884
rect 627 7876 1293 7884
rect 1367 7876 1493 7884
rect 1707 7876 1793 7884
rect 1807 7876 1853 7884
rect 2287 7876 2313 7884
rect 2707 7876 2853 7884
rect 2867 7876 2913 7884
rect 3087 7876 4073 7884
rect 4156 7884 4164 7896
rect 4867 7896 5293 7904
rect 5307 7896 5373 7904
rect 5487 7896 5513 7904
rect 5607 7896 6073 7904
rect 6107 7896 7013 7904
rect 7527 7896 8553 7904
rect 8567 7896 8633 7904
rect 8647 7896 9024 7904
rect 4156 7876 5553 7884
rect 5676 7876 6293 7884
rect 487 7856 673 7864
rect 687 7856 773 7864
rect 1267 7856 1533 7864
rect 1927 7856 1953 7864
rect 1976 7856 2033 7864
rect 127 7836 153 7844
rect 467 7836 613 7844
rect 167 7816 353 7824
rect 427 7816 473 7824
rect 636 7824 644 7833
rect 876 7827 884 7853
rect 1467 7836 1873 7844
rect 1896 7844 1904 7853
rect 1976 7844 1984 7856
rect 2047 7856 2333 7864
rect 2347 7856 2633 7864
rect 2887 7856 3113 7864
rect 3167 7856 3253 7864
rect 3787 7856 3964 7864
rect 1896 7836 1984 7844
rect 2147 7836 2273 7844
rect 2287 7836 2473 7844
rect 2567 7836 2733 7844
rect 2947 7836 3093 7844
rect 3167 7836 3233 7844
rect 3307 7836 3333 7844
rect 3507 7836 3933 7844
rect 3956 7844 3964 7856
rect 4307 7856 4633 7864
rect 4767 7856 4953 7864
rect 4967 7856 5073 7864
rect 5676 7864 5684 7876
rect 6427 7876 7493 7884
rect 7547 7876 7593 7884
rect 7647 7876 8313 7884
rect 8487 7876 8513 7884
rect 8647 7876 8693 7884
rect 8727 7876 8973 7884
rect 9016 7884 9024 7896
rect 9047 7896 9113 7904
rect 9127 7896 10333 7904
rect 10627 7896 10773 7904
rect 11587 7896 11733 7904
rect 12067 7896 12113 7904
rect 9016 7876 9193 7884
rect 9327 7876 9413 7884
rect 9427 7876 9993 7884
rect 10027 7876 10213 7884
rect 10227 7876 10753 7884
rect 11307 7876 11773 7884
rect 5167 7856 5684 7864
rect 6007 7856 6333 7864
rect 6527 7856 6913 7864
rect 6927 7856 6993 7864
rect 7727 7856 8613 7864
rect 8667 7856 8693 7864
rect 8907 7856 9053 7864
rect 9067 7856 9093 7864
rect 9307 7856 9593 7864
rect 9647 7856 9713 7864
rect 9727 7856 9853 7864
rect 9967 7856 10153 7864
rect 10347 7856 10413 7864
rect 10567 7856 10593 7864
rect 10747 7856 10764 7864
rect 3956 7836 4173 7844
rect 4227 7836 4813 7844
rect 4927 7836 5013 7844
rect 5047 7836 5113 7844
rect 5696 7844 5704 7853
rect 5387 7836 5704 7844
rect 607 7816 644 7824
rect 1107 7816 1133 7824
rect 1287 7816 1713 7824
rect 1727 7816 1813 7824
rect 1867 7816 1933 7824
rect 1947 7816 1973 7824
rect 2427 7816 2673 7824
rect 2827 7816 2873 7824
rect 2887 7816 3133 7824
rect 3356 7824 3364 7833
rect 3356 7816 3413 7824
rect 4047 7816 4213 7824
rect 4547 7816 5133 7824
rect 5156 7816 5293 7824
rect 147 7796 233 7804
rect 487 7796 533 7804
rect 587 7796 653 7804
rect 1327 7796 1513 7804
rect 1527 7796 1873 7804
rect 2127 7796 2453 7804
rect 2467 7796 2493 7804
rect 3267 7796 3313 7804
rect 3527 7796 3973 7804
rect 4007 7796 4193 7804
rect 4347 7796 4393 7804
rect 4467 7796 4513 7804
rect 4567 7796 4593 7804
rect 4907 7796 4913 7804
rect 4927 7796 4973 7804
rect 5156 7804 5164 7816
rect 5527 7816 5593 7824
rect 5696 7824 5704 7836
rect 5867 7836 6293 7844
rect 6387 7836 6593 7844
rect 6747 7836 6784 7844
rect 5696 7816 5733 7824
rect 6007 7816 6173 7824
rect 6776 7824 6784 7836
rect 7227 7836 7333 7844
rect 7387 7836 7433 7844
rect 7447 7836 7553 7844
rect 7747 7836 7773 7844
rect 8107 7836 8133 7844
rect 8367 7836 8553 7844
rect 8567 7836 8673 7844
rect 8727 7836 8833 7844
rect 8847 7836 8893 7844
rect 8947 7836 9253 7844
rect 9267 7836 9313 7844
rect 9827 7836 9873 7844
rect 10407 7836 10573 7844
rect 6367 7816 6564 7824
rect 6776 7816 6893 7824
rect 6556 7807 6564 7816
rect 7156 7824 7164 7833
rect 6947 7816 7164 7824
rect 7187 7816 7313 7824
rect 7367 7816 7493 7824
rect 7607 7816 7713 7824
rect 7727 7816 7873 7824
rect 5027 7796 5164 7804
rect 5287 7796 5413 7804
rect 5447 7796 5493 7804
rect 5687 7796 5853 7804
rect 6327 7796 6393 7804
rect 6527 7796 6544 7804
rect 1747 7776 2133 7784
rect 2407 7776 2533 7784
rect 2787 7776 2873 7784
rect 2927 7776 2933 7784
rect 2947 7776 2953 7784
rect 3087 7776 3233 7784
rect 3427 7776 3524 7784
rect 3387 7756 3453 7764
rect 3516 7764 3524 7776
rect 3547 7776 4033 7784
rect 4267 7776 4333 7784
rect 4387 7776 4793 7784
rect 4827 7776 4893 7784
rect 5087 7776 5533 7784
rect 5607 7776 6373 7784
rect 6536 7784 6544 7796
rect 6607 7796 6713 7804
rect 6867 7796 6893 7804
rect 7007 7796 7093 7804
rect 7107 7796 7373 7804
rect 7527 7796 7813 7804
rect 7896 7804 7904 7833
rect 10756 7827 10764 7856
rect 10807 7856 10853 7864
rect 11147 7856 11273 7864
rect 11287 7856 11393 7864
rect 11467 7856 11513 7864
rect 11807 7856 11973 7864
rect 12007 7856 12093 7864
rect 10867 7836 11493 7844
rect 11507 7836 12093 7844
rect 7927 7816 7953 7824
rect 8127 7816 8273 7824
rect 8307 7816 8373 7824
rect 8487 7816 8513 7824
rect 8827 7816 8913 7824
rect 9047 7816 9073 7824
rect 9127 7816 9273 7824
rect 9347 7816 9393 7824
rect 9587 7816 9833 7824
rect 9847 7816 9933 7824
rect 10107 7816 10373 7824
rect 10467 7816 10753 7824
rect 10887 7816 10933 7824
rect 11267 7816 11293 7824
rect 11347 7816 11393 7824
rect 11836 7816 11913 7824
rect 7896 7796 7913 7804
rect 8087 7796 8193 7804
rect 8447 7796 10593 7804
rect 10907 7796 11113 7804
rect 11327 7796 11373 7804
rect 11507 7796 11533 7804
rect 11587 7796 11713 7804
rect 11836 7804 11844 7816
rect 11727 7796 11844 7804
rect 11867 7796 11893 7804
rect 11947 7796 11973 7804
rect 12027 7796 12073 7804
rect 6536 7776 6973 7784
rect 7807 7776 7953 7784
rect 7987 7776 8073 7784
rect 8347 7776 8893 7784
rect 9647 7776 9733 7784
rect 11156 7784 11164 7793
rect 10967 7776 11393 7784
rect 11467 7776 11533 7784
rect 11747 7776 11813 7784
rect 3516 7756 3913 7764
rect 3967 7756 4073 7764
rect 4247 7756 5213 7764
rect 5587 7756 5673 7764
rect 6156 7756 6813 7764
rect 6156 7744 6164 7756
rect 7007 7756 8113 7764
rect 8847 7756 9433 7764
rect 10607 7756 11313 7764
rect 11327 7756 11353 7764
rect 2647 7736 6164 7744
rect 7107 7736 7213 7744
rect 7287 7736 8053 7744
rect 8087 7736 9413 7744
rect 10707 7736 10733 7744
rect 947 7716 1033 7724
rect 1047 7716 2053 7724
rect 2647 7716 5233 7724
rect 5247 7716 5973 7724
rect 6887 7716 9153 7724
rect 9167 7716 9353 7724
rect 10727 7716 11053 7724
rect 187 7696 213 7704
rect 2187 7696 2633 7704
rect 3227 7696 3313 7704
rect 3367 7696 4413 7704
rect 4767 7696 5913 7704
rect 5927 7696 8133 7704
rect 8147 7696 8433 7704
rect 8707 7696 9133 7704
rect 2507 7676 4573 7684
rect 4847 7676 4933 7684
rect 5167 7676 5553 7684
rect 5607 7676 5753 7684
rect 5767 7676 5953 7684
rect 5987 7676 6733 7684
rect 6987 7676 7073 7684
rect 8007 7676 8933 7684
rect 9527 7676 11093 7684
rect 987 7656 1213 7664
rect 1567 7656 2553 7664
rect 2867 7656 3573 7664
rect 3587 7656 6033 7664
rect 6047 7656 7033 7664
rect 7147 7656 7773 7664
rect 8627 7656 8913 7664
rect 9007 7656 9613 7664
rect 9887 7656 9993 7664
rect 10347 7656 11973 7664
rect 727 7636 793 7644
rect 807 7636 993 7644
rect 1787 7636 7193 7644
rect 7247 7636 7313 7644
rect 7587 7636 7613 7644
rect 7887 7636 11653 7644
rect 167 7616 413 7624
rect 427 7616 2153 7624
rect 2307 7616 2493 7624
rect 2567 7616 3353 7624
rect 3387 7616 3833 7624
rect 3847 7616 3873 7624
rect 3916 7616 3993 7624
rect 2227 7596 3033 7604
rect 3207 7596 3293 7604
rect 3367 7596 3433 7604
rect 3916 7604 3924 7616
rect 4087 7616 4373 7624
rect 4787 7616 5653 7624
rect 5667 7616 6153 7624
rect 6167 7616 6613 7624
rect 6627 7616 6633 7624
rect 6647 7616 7493 7624
rect 8187 7616 8333 7624
rect 8687 7616 9013 7624
rect 9187 7616 9353 7624
rect 9367 7616 10453 7624
rect 11627 7616 11673 7624
rect 3547 7596 3924 7604
rect 3987 7596 4484 7604
rect 467 7576 493 7584
rect 607 7576 693 7584
rect 1787 7576 2373 7584
rect 2387 7576 2473 7584
rect 3207 7576 3253 7584
rect 3467 7576 3593 7584
rect 4247 7576 4393 7584
rect 4476 7584 4484 7596
rect 4507 7596 4953 7604
rect 4967 7596 5053 7604
rect 5147 7596 5173 7604
rect 5547 7596 6693 7604
rect 7027 7596 7353 7604
rect 7627 7596 7653 7604
rect 8107 7596 8233 7604
rect 8267 7596 8613 7604
rect 8727 7596 8773 7604
rect 9067 7596 9193 7604
rect 9207 7596 9553 7604
rect 11247 7596 11264 7604
rect 4476 7576 4533 7584
rect 4607 7576 4813 7584
rect 4827 7576 5153 7584
rect 5207 7576 5393 7584
rect 5416 7576 5513 7584
rect 207 7556 373 7564
rect 387 7556 493 7564
rect 547 7556 713 7564
rect 736 7564 744 7573
rect 736 7556 893 7564
rect 1427 7556 1533 7564
rect 1567 7556 1733 7564
rect 1936 7556 1993 7564
rect 1936 7547 1944 7556
rect 2187 7556 2533 7564
rect 2396 7547 2404 7556
rect 2607 7556 2653 7564
rect 2667 7556 2693 7564
rect 2747 7556 2893 7564
rect 2967 7556 3073 7564
rect 3087 7556 3264 7564
rect 3256 7547 3264 7556
rect 3327 7556 3433 7564
rect 3567 7556 3633 7564
rect 4107 7556 4273 7564
rect 4296 7556 4353 7564
rect 147 7536 333 7544
rect 407 7536 1753 7544
rect 1987 7536 2353 7544
rect 2467 7536 2713 7544
rect 2736 7536 2984 7544
rect 187 7516 233 7524
rect 247 7516 393 7524
rect 687 7516 953 7524
rect 967 7516 1293 7524
rect 1607 7516 1793 7524
rect 1967 7516 2113 7524
rect 2736 7524 2744 7536
rect 2587 7516 2744 7524
rect 2927 7516 2953 7524
rect 2976 7524 2984 7536
rect 3407 7536 3433 7544
rect 4036 7536 4213 7544
rect 2976 7516 3093 7524
rect 3247 7516 3333 7524
rect 3816 7524 3824 7533
rect 4036 7524 4044 7536
rect 4296 7544 4304 7556
rect 4467 7556 4984 7564
rect 4267 7536 4304 7544
rect 4356 7536 4753 7544
rect 3667 7516 4044 7524
rect 4067 7516 4173 7524
rect 4267 7516 4293 7524
rect 4356 7524 4364 7536
rect 4976 7544 4984 7556
rect 5416 7564 5424 7576
rect 5907 7576 5933 7584
rect 5987 7576 6213 7584
rect 7427 7576 7833 7584
rect 8027 7576 8153 7584
rect 8387 7576 8753 7584
rect 8796 7567 8804 7593
rect 11256 7587 11264 7596
rect 8987 7576 9013 7584
rect 9167 7576 9244 7584
rect 5007 7556 5424 7564
rect 5967 7556 6113 7564
rect 6167 7556 6833 7564
rect 6887 7556 7013 7564
rect 7067 7556 7213 7564
rect 7227 7556 7244 7564
rect 4976 7536 5153 7544
rect 5187 7536 5253 7544
rect 5347 7536 5453 7544
rect 5667 7536 5704 7544
rect 4307 7516 4364 7524
rect 4387 7516 4413 7524
rect 4447 7516 4473 7524
rect 4647 7516 4873 7524
rect 5027 7516 5133 7524
rect 5147 7516 5653 7524
rect 5696 7524 5704 7536
rect 5807 7536 5884 7544
rect 5696 7516 5853 7524
rect 5876 7524 5884 7536
rect 5907 7536 6013 7544
rect 6027 7536 6173 7544
rect 6196 7536 7073 7544
rect 6196 7524 6204 7536
rect 7236 7544 7244 7556
rect 7267 7556 7433 7564
rect 7687 7556 8173 7564
rect 8227 7556 8273 7564
rect 8287 7556 8373 7564
rect 8527 7556 8553 7564
rect 8587 7556 8673 7564
rect 8896 7556 9193 7564
rect 7236 7536 7833 7544
rect 7867 7536 8013 7544
rect 8067 7536 8233 7544
rect 8247 7536 8353 7544
rect 8407 7536 8493 7544
rect 8607 7536 8633 7544
rect 8896 7544 8904 7556
rect 9207 7556 9213 7564
rect 9236 7564 9244 7576
rect 9267 7576 9753 7584
rect 11067 7576 11173 7584
rect 11336 7576 11433 7584
rect 9236 7556 9393 7564
rect 9487 7556 10493 7564
rect 11087 7556 11273 7564
rect 11336 7564 11344 7576
rect 11807 7576 11833 7584
rect 11907 7576 11993 7584
rect 11287 7556 11344 7564
rect 11367 7556 11553 7564
rect 11567 7556 11633 7564
rect 11827 7556 11933 7564
rect 11947 7556 11953 7564
rect 11987 7556 12013 7564
rect 8767 7536 8904 7544
rect 8927 7536 8973 7544
rect 9247 7536 9733 7544
rect 9887 7536 9893 7544
rect 9907 7536 9913 7544
rect 9967 7536 10013 7544
rect 10647 7536 10653 7544
rect 10667 7536 10833 7544
rect 11047 7536 11373 7544
rect 11627 7536 11833 7544
rect 5876 7516 6204 7524
rect 7307 7516 7793 7524
rect 7987 7516 8544 7524
rect 887 7496 913 7504
rect 1007 7496 1053 7504
rect 1067 7496 1333 7504
rect 1347 7496 1673 7504
rect 1967 7496 2013 7504
rect 2027 7496 2193 7504
rect 2307 7496 3173 7504
rect 3187 7496 3473 7504
rect 3487 7496 5833 7504
rect 5847 7496 6273 7504
rect 6287 7496 6293 7504
rect 6307 7496 7113 7504
rect 7127 7496 8513 7504
rect 8536 7504 8544 7516
rect 8567 7516 8653 7524
rect 8747 7516 8813 7524
rect 9387 7516 9533 7524
rect 9727 7516 9793 7524
rect 9947 7516 10073 7524
rect 10127 7516 10633 7524
rect 11307 7516 11453 7524
rect 8536 7496 8953 7504
rect 9127 7496 9573 7504
rect 9587 7496 9653 7504
rect 9807 7496 10253 7504
rect 10267 7496 10433 7504
rect 10527 7496 10853 7504
rect 2347 7476 2753 7484
rect 3287 7476 3613 7484
rect 3647 7476 4093 7484
rect 4207 7476 4293 7484
rect 4347 7476 4793 7484
rect 4947 7476 5113 7484
rect 5167 7476 6053 7484
rect 6127 7476 6193 7484
rect 6867 7476 7793 7484
rect 7967 7476 8613 7484
rect 9767 7476 10033 7484
rect 10567 7476 10673 7484
rect 10896 7476 11193 7484
rect 367 7456 1233 7464
rect 1947 7456 3473 7464
rect 3487 7456 3973 7464
rect 4036 7456 4633 7464
rect 867 7436 1193 7444
rect 2247 7436 2493 7444
rect 4036 7444 4044 7456
rect 4667 7456 5153 7464
rect 5227 7456 5633 7464
rect 5667 7456 6073 7464
rect 6107 7456 6453 7464
rect 6887 7456 6953 7464
rect 7087 7456 7193 7464
rect 7207 7456 7293 7464
rect 7416 7456 7553 7464
rect 2587 7436 4044 7444
rect 4067 7436 4113 7444
rect 4187 7436 4993 7444
rect 5007 7436 5753 7444
rect 6147 7436 6473 7444
rect 7416 7444 7424 7456
rect 7667 7456 7993 7464
rect 8127 7456 8813 7464
rect 8827 7456 9133 7464
rect 10896 7464 10904 7476
rect 11887 7476 12033 7484
rect 12047 7476 12073 7484
rect 9567 7456 10904 7464
rect 10927 7456 11953 7464
rect 11967 7456 12073 7464
rect 6807 7436 7424 7444
rect 7447 7436 8113 7444
rect 8227 7436 8273 7444
rect 8467 7436 8533 7444
rect 8687 7436 9513 7444
rect 9547 7436 9833 7444
rect 11187 7436 12053 7444
rect 1687 7416 2293 7424
rect 3007 7416 3333 7424
rect 3347 7416 3453 7424
rect 3467 7416 3533 7424
rect 3707 7416 3873 7424
rect 3887 7416 4493 7424
rect 4507 7416 6233 7424
rect 6247 7416 6293 7424
rect 6647 7416 7173 7424
rect 7447 7416 7473 7424
rect 7627 7416 7713 7424
rect 7867 7416 10173 7424
rect 10187 7416 10413 7424
rect 667 7396 713 7404
rect 1107 7396 2573 7404
rect 2767 7396 2993 7404
rect 3127 7396 3733 7404
rect 3987 7396 4913 7404
rect 5016 7396 7133 7404
rect 587 7376 813 7384
rect 1787 7376 1933 7384
rect 2547 7376 2713 7384
rect 2787 7376 2933 7384
rect 2947 7376 3093 7384
rect 3147 7376 3673 7384
rect 3747 7376 3784 7384
rect 187 7356 313 7364
rect 367 7356 533 7364
rect 556 7356 613 7364
rect 227 7336 273 7344
rect 287 7336 333 7344
rect 556 7344 564 7356
rect 627 7356 673 7364
rect 1167 7356 1253 7364
rect 2907 7356 3053 7364
rect 3107 7356 3284 7364
rect 387 7336 564 7344
rect 647 7336 693 7344
rect 1287 7336 1793 7344
rect 1867 7336 2133 7344
rect 2407 7336 2513 7344
rect 2747 7336 2773 7344
rect 2827 7336 2913 7344
rect 2967 7336 2993 7344
rect 3276 7344 3284 7356
rect 3307 7356 3344 7364
rect 3276 7336 3313 7344
rect 3336 7344 3344 7356
rect 3427 7356 3513 7364
rect 3627 7356 3693 7364
rect 3776 7364 3784 7376
rect 3967 7376 3993 7384
rect 4047 7376 4113 7384
rect 4147 7376 4313 7384
rect 5016 7384 5024 7396
rect 7187 7396 7233 7404
rect 7687 7396 7833 7404
rect 7847 7396 8093 7404
rect 8107 7396 8673 7404
rect 8696 7396 8873 7404
rect 4367 7376 5024 7384
rect 5047 7376 5353 7384
rect 5407 7376 5773 7384
rect 6047 7376 6133 7384
rect 6187 7376 6633 7384
rect 6727 7376 6753 7384
rect 6767 7376 6993 7384
rect 7387 7376 7593 7384
rect 7667 7376 7733 7384
rect 7907 7376 7933 7384
rect 8327 7376 8453 7384
rect 8696 7384 8704 7396
rect 8887 7396 9533 7404
rect 10927 7396 11733 7404
rect 11747 7396 11893 7404
rect 8487 7376 8704 7384
rect 8727 7376 8793 7384
rect 8947 7376 8973 7384
rect 9187 7376 9313 7384
rect 9467 7376 9533 7384
rect 9867 7376 9893 7384
rect 10027 7376 10053 7384
rect 10087 7376 10233 7384
rect 10247 7376 10293 7384
rect 10507 7376 10593 7384
rect 10787 7376 10973 7384
rect 11467 7376 11684 7384
rect 11676 7367 11684 7376
rect 11947 7376 12013 7384
rect 3776 7356 3793 7364
rect 3807 7356 3953 7364
rect 4107 7356 4213 7364
rect 4347 7356 4453 7364
rect 4647 7356 4673 7364
rect 4727 7356 4773 7364
rect 4967 7356 5133 7364
rect 5156 7356 5193 7364
rect 3336 7336 3533 7344
rect 3567 7336 3713 7344
rect 3907 7336 4173 7344
rect 4387 7336 4513 7344
rect 4587 7336 4733 7344
rect 4907 7336 4973 7344
rect 5156 7344 5164 7356
rect 5207 7356 5213 7364
rect 5287 7356 5393 7364
rect 5587 7356 5613 7364
rect 5767 7356 5833 7364
rect 5847 7356 6893 7364
rect 6907 7356 6913 7364
rect 6936 7356 6973 7364
rect 6936 7347 6944 7356
rect 6987 7356 7073 7364
rect 7296 7356 7753 7364
rect 5127 7336 5164 7344
rect 5387 7336 5413 7344
rect 5476 7336 5653 7344
rect 127 7316 553 7324
rect 667 7316 793 7324
rect 807 7316 1333 7324
rect 1347 7316 1973 7324
rect 2567 7316 2613 7324
rect 2707 7316 2813 7324
rect 2827 7316 3153 7324
rect 3467 7316 3493 7324
rect 4027 7316 4533 7324
rect 4707 7316 4933 7324
rect 4947 7316 5333 7324
rect 5476 7324 5484 7336
rect 5687 7336 5973 7344
rect 6067 7336 6873 7344
rect 7296 7344 7304 7356
rect 7847 7356 7953 7364
rect 7967 7356 8253 7364
rect 8627 7356 8673 7364
rect 9347 7356 9513 7364
rect 10007 7356 10193 7364
rect 10467 7356 10784 7364
rect 7167 7336 7304 7344
rect 7327 7336 7373 7344
rect 7396 7336 7533 7344
rect 5347 7316 5484 7324
rect 6127 7316 6193 7324
rect 6947 7316 7093 7324
rect 7396 7324 7404 7336
rect 7587 7336 7693 7344
rect 7756 7336 7773 7344
rect 7756 7327 7764 7336
rect 8067 7336 8253 7344
rect 8267 7336 8724 7344
rect 7347 7316 7404 7324
rect 7607 7316 7633 7324
rect 7907 7316 7953 7324
rect 8047 7316 8693 7324
rect 8716 7324 8724 7336
rect 9007 7336 9113 7344
rect 9167 7336 9253 7344
rect 9367 7336 10164 7344
rect 8716 7316 8753 7324
rect 8907 7316 9073 7324
rect 9087 7316 9313 7324
rect 10156 7324 10164 7336
rect 10187 7336 10573 7344
rect 10647 7336 10753 7344
rect 10776 7344 10784 7356
rect 11447 7356 11473 7364
rect 10776 7336 10793 7344
rect 10956 7327 10964 7353
rect 11327 7336 11493 7344
rect 12056 7344 12064 7353
rect 11927 7336 12064 7344
rect 10156 7316 10913 7324
rect 11487 7316 11533 7324
rect 11627 7316 11693 7324
rect 12027 7316 12093 7324
rect 267 7296 333 7304
rect 1647 7296 1933 7304
rect 2687 7296 3213 7304
rect 3227 7296 3453 7304
rect 4327 7296 4393 7304
rect 4407 7296 5273 7304
rect 5527 7296 6213 7304
rect 7147 7296 7273 7304
rect 7367 7296 7413 7304
rect 7487 7296 7573 7304
rect 8287 7296 8313 7304
rect 8507 7296 9333 7304
rect 9907 7296 10273 7304
rect 10387 7296 10633 7304
rect 10647 7296 11153 7304
rect 2607 7276 3304 7284
rect 3296 7264 3304 7276
rect 3487 7276 3824 7284
rect 3296 7256 3633 7264
rect 3816 7264 3824 7276
rect 4287 7276 4713 7284
rect 4727 7276 5353 7284
rect 5367 7276 6773 7284
rect 6787 7276 8233 7284
rect 10747 7276 10993 7284
rect 11007 7276 11533 7284
rect 3816 7256 3893 7264
rect 3907 7256 4433 7264
rect 4447 7256 4573 7264
rect 4587 7256 7233 7264
rect 7247 7256 7873 7264
rect 8207 7256 8473 7264
rect 1567 7236 1833 7244
rect 1887 7236 4353 7244
rect 5167 7236 5553 7244
rect 5567 7236 5933 7244
rect 5947 7236 6153 7244
rect 6227 7236 6493 7244
rect 6507 7236 11873 7244
rect 887 7216 1653 7224
rect 1827 7216 2893 7224
rect 3087 7216 3473 7224
rect 3527 7216 3713 7224
rect 3727 7216 4113 7224
rect 4527 7216 4953 7224
rect 5067 7216 5413 7224
rect 5547 7216 5613 7224
rect 5667 7216 6713 7224
rect 6787 7216 7253 7224
rect 8167 7216 9233 7224
rect 11687 7216 11773 7224
rect 3727 7196 3793 7204
rect 3947 7196 4033 7204
rect 4047 7196 4353 7204
rect 4627 7196 7033 7204
rect 7087 7196 7733 7204
rect 7747 7196 8633 7204
rect 8647 7196 9273 7204
rect 10627 7196 11773 7204
rect 1907 7176 3133 7184
rect 3367 7176 3633 7184
rect 4007 7176 4313 7184
rect 4327 7176 4933 7184
rect 4987 7176 5393 7184
rect 5467 7176 5873 7184
rect 5887 7176 6173 7184
rect 6567 7176 6593 7184
rect 6707 7176 7773 7184
rect 8187 7176 11753 7184
rect 1347 7156 1393 7164
rect 1907 7156 2073 7164
rect 2087 7156 2433 7164
rect 2487 7156 2573 7164
rect 2727 7156 2793 7164
rect 3127 7156 3193 7164
rect 3627 7156 3653 7164
rect 3687 7156 3793 7164
rect 3807 7156 4413 7164
rect 4607 7156 4773 7164
rect 5467 7156 5933 7164
rect 6087 7156 6433 7164
rect 6467 7156 7993 7164
rect 10847 7156 11153 7164
rect 2047 7136 2233 7144
rect 2247 7136 2413 7144
rect 2427 7136 2613 7144
rect 3307 7136 3693 7144
rect 3796 7136 4193 7144
rect 607 7116 2113 7124
rect 2127 7116 2533 7124
rect 2987 7116 3184 7124
rect 167 7096 753 7104
rect 767 7096 933 7104
rect 1347 7096 1713 7104
rect 1767 7096 2273 7104
rect 2287 7096 2593 7104
rect 2636 7096 2933 7104
rect 147 7076 193 7084
rect 216 7076 293 7084
rect 216 7064 224 7076
rect 347 7076 684 7084
rect 187 7056 224 7064
rect 287 7056 493 7064
rect 676 7064 684 7076
rect 707 7076 1093 7084
rect 1527 7076 1984 7084
rect 676 7056 733 7064
rect 1127 7056 1293 7064
rect 1327 7056 1453 7064
rect 1547 7056 1653 7064
rect 1676 7064 1684 7076
rect 1676 7056 1693 7064
rect 1727 7056 1833 7064
rect 1847 7056 1913 7064
rect 1976 7064 1984 7076
rect 2636 7084 2644 7096
rect 2987 7096 3153 7104
rect 3176 7104 3184 7116
rect 3267 7116 3393 7124
rect 3407 7116 3473 7124
rect 3796 7124 3804 7136
rect 4207 7136 4513 7144
rect 5207 7136 5273 7144
rect 5847 7136 7673 7144
rect 8147 7136 10333 7144
rect 10347 7136 10813 7144
rect 3487 7116 3804 7124
rect 3847 7116 4293 7124
rect 4807 7116 5593 7124
rect 5767 7116 6013 7124
rect 6207 7116 6533 7124
rect 7047 7116 7484 7124
rect 3176 7096 3193 7104
rect 3767 7096 4053 7104
rect 4136 7096 4173 7104
rect 2047 7076 2644 7084
rect 2667 7076 2753 7084
rect 3227 7076 3253 7084
rect 3327 7076 3373 7084
rect 3427 7076 3533 7084
rect 3767 7076 3833 7084
rect 4136 7084 4144 7096
rect 4367 7096 4673 7104
rect 4807 7096 5273 7104
rect 5316 7096 5684 7104
rect 3967 7076 4144 7084
rect 4167 7076 4333 7084
rect 4356 7076 4773 7084
rect 1976 7056 2684 7064
rect 167 7036 353 7044
rect 367 7036 533 7044
rect 967 7036 1053 7044
rect 1147 7036 1313 7044
rect 1327 7036 1353 7044
rect 1367 7036 1573 7044
rect 1667 7036 1853 7044
rect 2267 7036 2353 7044
rect 2676 7044 2684 7056
rect 2747 7056 2833 7064
rect 3187 7056 3293 7064
rect 3367 7056 3553 7064
rect 3607 7056 3653 7064
rect 3707 7056 3733 7064
rect 4356 7064 4364 7076
rect 5316 7084 5324 7096
rect 4967 7076 5324 7084
rect 5336 7076 5453 7084
rect 3927 7056 4364 7064
rect 4667 7056 4693 7064
rect 4767 7056 4913 7064
rect 4936 7064 4944 7073
rect 5336 7067 5344 7076
rect 5587 7076 5653 7084
rect 5676 7084 5684 7096
rect 5707 7096 5833 7104
rect 5867 7096 5893 7104
rect 5907 7096 6373 7104
rect 6447 7096 6553 7104
rect 6887 7096 6913 7104
rect 7476 7104 7484 7116
rect 7507 7116 8153 7124
rect 8607 7116 8913 7124
rect 9047 7116 9133 7124
rect 7127 7096 7164 7104
rect 7476 7096 7544 7104
rect 7156 7087 7164 7096
rect 5676 7076 5713 7084
rect 5727 7076 5873 7084
rect 5956 7076 6113 7084
rect 5956 7067 5964 7076
rect 6247 7076 6513 7084
rect 6627 7076 6673 7084
rect 7467 7076 7513 7084
rect 7536 7084 7544 7096
rect 7567 7096 7693 7104
rect 7707 7096 8873 7104
rect 8936 7096 9093 7104
rect 8936 7087 8944 7096
rect 10027 7096 10093 7104
rect 10307 7096 11013 7104
rect 11307 7096 11353 7104
rect 11407 7096 11564 7104
rect 11556 7087 11564 7096
rect 7536 7076 7564 7084
rect 4936 7056 5133 7064
rect 5267 7056 5313 7064
rect 5387 7056 5473 7064
rect 5487 7056 5493 7064
rect 5727 7056 5944 7064
rect 2676 7036 2773 7044
rect 2807 7036 3373 7044
rect 3407 7036 3573 7044
rect 3787 7036 3873 7044
rect 3887 7036 4033 7044
rect 4147 7036 4213 7044
rect 4307 7036 4733 7044
rect 4847 7036 5113 7044
rect 5307 7036 5333 7044
rect 5407 7036 5604 7044
rect 547 7016 1493 7024
rect 2647 7016 2933 7024
rect 3007 7016 3073 7024
rect 3367 7016 3933 7024
rect 4727 7016 4813 7024
rect 4967 7016 5193 7024
rect 5207 7016 5553 7024
rect 5596 7024 5604 7036
rect 5667 7036 5773 7044
rect 5936 7044 5944 7056
rect 6067 7056 6133 7064
rect 6156 7056 6813 7064
rect 6156 7044 6164 7056
rect 7016 7064 7024 7073
rect 6847 7056 7453 7064
rect 7556 7064 7564 7076
rect 7587 7076 7653 7084
rect 7927 7076 8173 7084
rect 8096 7067 8104 7076
rect 8587 7076 8713 7084
rect 8727 7076 8833 7084
rect 8847 7076 8893 7084
rect 9087 7076 9113 7084
rect 9207 7076 9273 7084
rect 9347 7076 9653 7084
rect 9707 7076 9853 7084
rect 10127 7076 10493 7084
rect 7556 7056 7893 7064
rect 7947 7056 8033 7064
rect 8047 7056 8053 7064
rect 8187 7056 8693 7064
rect 8787 7056 9313 7064
rect 9427 7056 9513 7064
rect 9727 7056 9833 7064
rect 10087 7056 10253 7064
rect 10487 7056 10653 7064
rect 10876 7064 10884 7073
rect 10876 7056 10913 7064
rect 10927 7056 11033 7064
rect 11227 7056 11373 7064
rect 11527 7056 11713 7064
rect 5787 7036 5924 7044
rect 5936 7036 6164 7044
rect 5596 7016 5613 7024
rect 5707 7016 5893 7024
rect 5916 7024 5924 7036
rect 6587 7036 6693 7044
rect 6927 7036 7033 7044
rect 7047 7036 7093 7044
rect 7316 7036 7333 7044
rect 5916 7016 6073 7024
rect 6187 7016 6833 7024
rect 1067 6996 1473 7004
rect 1487 6996 2053 7004
rect 3087 6996 4533 7004
rect 4767 6996 5753 7004
rect 5807 6996 6173 7004
rect 6267 6996 6333 7004
rect 6567 6996 7193 7004
rect 7316 7004 7324 7036
rect 7827 7036 8073 7044
rect 8687 7036 8733 7044
rect 9507 7036 10293 7044
rect 10327 7036 10453 7044
rect 11107 7036 11193 7044
rect 11607 7036 11733 7044
rect 7347 7016 7573 7024
rect 7807 7016 7873 7024
rect 7887 7016 7933 7024
rect 8487 7016 9893 7024
rect 10167 7016 10673 7024
rect 7296 6996 7324 7004
rect 7296 6987 7304 6996
rect 7407 6996 7453 7004
rect 7467 6996 7633 7004
rect 7707 6996 8453 7004
rect 8467 6996 8713 7004
rect 9227 6996 10433 7004
rect 687 6976 733 6984
rect 747 6976 1133 6984
rect 1367 6976 1953 6984
rect 2387 6976 4433 6984
rect 4447 6976 6653 6984
rect 6727 6976 7033 6984
rect 7587 6976 7833 6984
rect 8007 6976 8373 6984
rect 8887 6976 10033 6984
rect 947 6956 1673 6964
rect 1807 6956 7013 6964
rect 7227 6956 7373 6964
rect 7427 6956 7473 6964
rect 7867 6956 7993 6964
rect 8327 6956 8673 6964
rect 9207 6956 9473 6964
rect 1827 6936 2033 6944
rect 2047 6936 6244 6944
rect 107 6916 693 6924
rect 707 6916 1893 6924
rect 2247 6916 2613 6924
rect 2647 6916 3353 6924
rect 3447 6916 4333 6924
rect 4427 6916 4793 6924
rect 4807 6916 4813 6924
rect 4887 6916 4993 6924
rect 5047 6916 5173 6924
rect 5227 6916 5453 6924
rect 5487 6916 5733 6924
rect 5827 6916 5973 6924
rect 6236 6924 6244 6936
rect 6267 6936 6513 6944
rect 6547 6936 7133 6944
rect 7267 6936 7533 6944
rect 7547 6936 7693 6944
rect 7867 6936 8253 6944
rect 8327 6936 9453 6944
rect 10647 6936 10853 6944
rect 10907 6936 10973 6944
rect 10987 6936 11573 6944
rect 6236 6916 6344 6924
rect 187 6896 553 6904
rect 567 6896 653 6904
rect 1667 6896 1833 6904
rect 2207 6896 2393 6904
rect 2787 6896 2973 6904
rect 3487 6896 3593 6904
rect 3847 6896 3953 6904
rect 4187 6896 4413 6904
rect 4507 6896 4753 6904
rect 4787 6896 5133 6904
rect 5187 6896 5253 6904
rect 5287 6896 5313 6904
rect 5327 6896 5693 6904
rect 5736 6896 5913 6904
rect 347 6876 473 6884
rect 487 6876 1013 6884
rect 1247 6876 1613 6884
rect 1927 6876 1993 6884
rect 2287 6876 2573 6884
rect 2596 6867 2604 6893
rect 3007 6876 3153 6884
rect 3227 6876 3373 6884
rect 3547 6876 3633 6884
rect 3987 6876 4013 6884
rect 4067 6876 4633 6884
rect 4707 6876 4733 6884
rect 4787 6876 4824 6884
rect 147 6856 333 6864
rect 807 6856 893 6864
rect 947 6856 1073 6864
rect 1227 6856 1273 6864
rect 1447 6856 1633 6864
rect 1996 6856 2233 6864
rect 167 6836 193 6844
rect 207 6836 353 6844
rect 576 6844 584 6853
rect 536 6836 584 6844
rect 536 6827 544 6836
rect 727 6836 1253 6844
rect 1327 6836 1413 6844
rect 1887 6836 1973 6844
rect 1996 6844 2004 6856
rect 2707 6856 2793 6864
rect 2927 6856 3053 6864
rect 3067 6856 3393 6864
rect 3787 6856 3833 6864
rect 4167 6856 4213 6864
rect 4336 6856 4473 6864
rect 4336 6847 4344 6856
rect 4487 6856 4593 6864
rect 4647 6856 4753 6864
rect 4776 6856 4793 6864
rect 1987 6836 2004 6844
rect 2027 6836 2033 6844
rect 2047 6836 2213 6844
rect 3147 6836 4133 6844
rect 4407 6836 4613 6844
rect 4727 6836 4753 6844
rect 1267 6816 2173 6824
rect 2907 6816 3393 6824
rect 3667 6816 3773 6824
rect 3867 6816 3973 6824
rect 4027 6816 4113 6824
rect 4167 6816 4233 6824
rect 4356 6824 4364 6833
rect 4327 6816 4364 6824
rect 4776 6824 4784 6856
rect 4816 6864 4824 6876
rect 4867 6876 4973 6884
rect 5027 6876 5053 6884
rect 5087 6876 5273 6884
rect 5307 6876 5373 6884
rect 5736 6884 5744 6896
rect 6027 6896 6313 6904
rect 6336 6904 6344 6916
rect 6367 6916 6533 6924
rect 6567 6916 6773 6924
rect 6927 6916 6993 6924
rect 7047 6916 7493 6924
rect 7507 6916 8073 6924
rect 8447 6916 8533 6924
rect 9027 6916 9233 6924
rect 10867 6916 11133 6924
rect 11147 6916 11333 6924
rect 11347 6916 11533 6924
rect 11547 6916 11693 6924
rect 11707 6916 12113 6924
rect 6336 6896 6713 6904
rect 6787 6896 7213 6904
rect 7247 6896 7524 6904
rect 5567 6876 5744 6884
rect 5856 6876 5933 6884
rect 4816 6856 4953 6864
rect 5127 6856 5193 6864
rect 5327 6856 5353 6864
rect 5607 6856 5713 6864
rect 5856 6864 5864 6876
rect 6296 6876 6573 6884
rect 5747 6856 5864 6864
rect 5887 6856 5913 6864
rect 5967 6856 6013 6864
rect 6296 6864 6304 6876
rect 6707 6876 6833 6884
rect 6867 6876 7304 6884
rect 6207 6856 6304 6864
rect 6327 6856 6433 6864
rect 7087 6856 7273 6864
rect 7296 6864 7304 6876
rect 7327 6876 7453 6884
rect 7516 6884 7524 6896
rect 7547 6896 7893 6904
rect 9227 6896 9333 6904
rect 9407 6896 9713 6904
rect 10067 6896 10473 6904
rect 10487 6896 10573 6904
rect 10627 6896 10673 6904
rect 11187 6896 11213 6904
rect 11227 6896 11373 6904
rect 7516 6876 7553 6884
rect 7727 6876 7793 6884
rect 7907 6876 8033 6884
rect 8096 6876 8313 6884
rect 8096 6867 8104 6876
rect 8347 6876 8493 6884
rect 9127 6876 9533 6884
rect 9587 6876 9613 6884
rect 9627 6876 9693 6884
rect 9707 6876 9873 6884
rect 10207 6876 10593 6884
rect 10887 6876 11013 6884
rect 11047 6876 11313 6884
rect 11327 6876 11393 6884
rect 11747 6876 11913 6884
rect 7296 6856 7533 6864
rect 7567 6856 7653 6864
rect 7687 6856 7713 6864
rect 7747 6856 7873 6864
rect 7887 6856 8053 6864
rect 8527 6856 8653 6864
rect 8707 6856 8853 6864
rect 9387 6856 9473 6864
rect 9727 6856 9924 6864
rect 4807 6836 4833 6844
rect 5067 6836 5133 6844
rect 5556 6827 5564 6853
rect 5627 6836 5953 6844
rect 6136 6844 6144 6853
rect 6027 6836 6144 6844
rect 6287 6836 6384 6844
rect 4687 6816 5073 6824
rect 5107 6816 5213 6824
rect 5707 6816 5933 6824
rect 6056 6816 6193 6824
rect 1467 6796 1913 6804
rect 2007 6796 2373 6804
rect 2387 6796 3433 6804
rect 3467 6796 3473 6804
rect 3487 6796 4813 6804
rect 4907 6796 5173 6804
rect 5187 6796 5613 6804
rect 5647 6796 5693 6804
rect 6056 6804 6064 6816
rect 6376 6824 6384 6836
rect 6587 6836 7264 6844
rect 6376 6816 6453 6824
rect 6527 6816 6804 6824
rect 5747 6796 6064 6804
rect 6087 6796 6553 6804
rect 6676 6796 6773 6804
rect 2107 6776 2413 6784
rect 2427 6776 3073 6784
rect 3667 6776 4933 6784
rect 4967 6776 5113 6784
rect 5287 6776 5513 6784
rect 5527 6776 6113 6784
rect 6676 6784 6684 6796
rect 6796 6804 6804 6816
rect 6907 6816 7113 6824
rect 7256 6824 7264 6836
rect 7287 6836 7393 6844
rect 7467 6836 7633 6844
rect 7687 6836 7833 6844
rect 8027 6836 8133 6844
rect 8147 6836 8273 6844
rect 8307 6836 8473 6844
rect 8867 6836 9013 6844
rect 9687 6836 9773 6844
rect 9916 6844 9924 6856
rect 9947 6856 10033 6864
rect 10107 6856 10264 6864
rect 9916 6836 10113 6844
rect 10256 6844 10264 6856
rect 10287 6856 10313 6864
rect 10816 6847 10824 6873
rect 10847 6856 10913 6864
rect 11047 6856 11193 6864
rect 11407 6856 11713 6864
rect 11976 6864 11984 6873
rect 11767 6856 12133 6864
rect 10256 6836 10293 6844
rect 7256 6816 7553 6824
rect 7607 6816 7693 6824
rect 10047 6816 10073 6824
rect 10587 6816 11113 6824
rect 11127 6816 11353 6824
rect 11627 6816 12073 6824
rect 6796 6796 7213 6804
rect 7287 6796 8333 6804
rect 8767 6796 8993 6804
rect 9747 6796 9753 6804
rect 9767 6796 10453 6804
rect 10467 6796 10993 6804
rect 6127 6776 6684 6784
rect 6707 6776 8253 6784
rect 8267 6776 8413 6784
rect 8747 6776 8973 6784
rect 8987 6776 9053 6784
rect 10787 6776 10873 6784
rect 1167 6756 2393 6764
rect 2807 6756 4253 6764
rect 4567 6756 5533 6764
rect 5987 6756 5993 6764
rect 6007 6756 6253 6764
rect 6376 6756 6633 6764
rect 1607 6736 2273 6744
rect 2987 6736 3113 6744
rect 3187 6736 3733 6744
rect 4047 6736 4133 6744
rect 4247 6736 4564 6744
rect 2587 6716 3653 6724
rect 3687 6716 3793 6724
rect 3807 6716 3913 6724
rect 4307 6716 4373 6724
rect 4556 6724 4564 6736
rect 4587 6736 4673 6744
rect 4756 6736 5393 6744
rect 4756 6724 4764 6736
rect 6376 6744 6384 6756
rect 6687 6756 7333 6764
rect 7727 6756 9273 6764
rect 9287 6756 9953 6764
rect 9967 6756 10053 6764
rect 10467 6756 11293 6764
rect 5907 6736 6384 6744
rect 6407 6736 7273 6744
rect 7387 6736 8713 6744
rect 4556 6716 4764 6724
rect 4787 6716 5053 6724
rect 5207 6716 5253 6724
rect 5467 6716 6293 6724
rect 6427 6716 6893 6724
rect 6967 6716 7113 6724
rect 7387 6716 7873 6724
rect 8067 6716 8193 6724
rect 9307 6716 9813 6724
rect 3207 6696 3233 6704
rect 3827 6696 3933 6704
rect 4087 6696 4873 6704
rect 4887 6696 4993 6704
rect 5127 6696 6393 6704
rect 6467 6696 6533 6704
rect 6647 6696 6704 6704
rect 2407 6676 6633 6684
rect 6696 6684 6704 6696
rect 6727 6696 6773 6704
rect 6787 6696 7233 6704
rect 7547 6696 7753 6704
rect 6696 6676 6953 6684
rect 7047 6676 7573 6684
rect 7627 6676 9973 6684
rect 527 6656 2373 6664
rect 3527 6656 3693 6664
rect 4027 6656 4093 6664
rect 4127 6656 4584 6664
rect 407 6636 693 6644
rect 1167 6636 2193 6644
rect 2247 6636 2433 6644
rect 2447 6636 2653 6644
rect 2847 6636 3284 6644
rect 167 6616 393 6624
rect 407 6616 433 6624
rect 1487 6616 1693 6624
rect 1707 6616 1793 6624
rect 1847 6616 2033 6624
rect 3276 6624 3284 6636
rect 3307 6636 3453 6644
rect 3887 6636 4553 6644
rect 4576 6644 4584 6656
rect 4687 6656 7053 6664
rect 7067 6656 7153 6664
rect 7767 6656 7933 6664
rect 4576 6636 4893 6644
rect 4987 6636 5173 6644
rect 5696 6636 6013 6644
rect 2307 6616 2884 6624
rect 3276 6616 3753 6624
rect 176 6596 353 6604
rect 176 6587 184 6596
rect 1287 6596 1304 6604
rect 347 6576 493 6584
rect 527 6576 553 6584
rect 607 6576 744 6584
rect 736 6567 744 6576
rect 767 6576 913 6584
rect 927 6576 973 6584
rect 1227 6576 1253 6584
rect 1296 6584 1304 6596
rect 1327 6596 1613 6604
rect 1667 6596 1864 6604
rect 1856 6587 1864 6596
rect 1887 6596 1993 6604
rect 2047 6596 2593 6604
rect 2876 6604 2884 6616
rect 3927 6616 4713 6624
rect 4827 6616 5153 6624
rect 5167 6616 5293 6624
rect 5367 6616 5453 6624
rect 5696 6624 5704 6636
rect 6187 6636 6333 6644
rect 6947 6636 6973 6644
rect 7367 6636 7413 6644
rect 7467 6636 7593 6644
rect 9047 6636 9893 6644
rect 11427 6636 11473 6644
rect 11807 6636 11833 6644
rect 5567 6616 5704 6624
rect 2647 6596 2684 6604
rect 2876 6596 2993 6604
rect 2676 6587 2684 6596
rect 3307 6596 3373 6604
rect 3467 6596 3553 6604
rect 3727 6596 3833 6604
rect 3847 6596 3953 6604
rect 3967 6596 4053 6604
rect 4247 6596 4313 6604
rect 4627 6596 4673 6604
rect 4807 6596 4973 6604
rect 5007 6596 5233 6604
rect 5296 6596 5373 6604
rect 1296 6576 1633 6584
rect 2207 6576 2253 6584
rect 2387 6576 2453 6584
rect 2547 6576 2613 6584
rect 2967 6576 2993 6584
rect 3547 6576 3693 6584
rect 3767 6576 3853 6584
rect 3907 6576 4113 6584
rect 4247 6576 4293 6584
rect 4476 6567 4484 6593
rect 4707 6576 4773 6584
rect 4947 6576 5264 6584
rect 5256 6567 5264 6576
rect 5296 6584 5304 6596
rect 5547 6596 5613 6604
rect 5636 6604 5644 6616
rect 5727 6616 6653 6624
rect 6767 6616 6953 6624
rect 6967 6616 7493 6624
rect 7507 6616 7613 6624
rect 8127 6616 8593 6624
rect 8836 6616 9233 6624
rect 8836 6607 8844 6616
rect 9247 6616 9293 6624
rect 9547 6616 9573 6624
rect 9667 6616 9913 6624
rect 9927 6616 10013 6624
rect 10387 6616 10773 6624
rect 11376 6616 11573 6624
rect 5636 6596 5653 6604
rect 5767 6596 5833 6604
rect 6027 6596 6113 6604
rect 6376 6596 6564 6604
rect 5287 6576 5304 6584
rect 5476 6584 5484 6593
rect 5327 6576 5484 6584
rect 5667 6576 5693 6584
rect 6376 6584 6384 6596
rect 6556 6587 6564 6596
rect 6687 6596 6733 6604
rect 7127 6596 7573 6604
rect 7627 6596 7933 6604
rect 7947 6596 8173 6604
rect 8207 6596 8273 6604
rect 8327 6596 8433 6604
rect 8447 6596 8593 6604
rect 8647 6596 8673 6604
rect 8867 6596 9073 6604
rect 9267 6596 9973 6604
rect 9987 6596 10153 6604
rect 10207 6596 10253 6604
rect 10327 6596 10393 6604
rect 10587 6596 10673 6604
rect 10687 6596 10773 6604
rect 11027 6596 11053 6604
rect 11327 6596 11353 6604
rect 6227 6576 6384 6584
rect 6407 6576 6513 6584
rect 6667 6576 6793 6584
rect 6936 6584 6944 6593
rect 11376 6587 11384 6616
rect 12007 6616 12033 6624
rect 11407 6596 11453 6604
rect 11736 6596 11753 6604
rect 6936 6576 6973 6584
rect 7207 6576 7864 6584
rect 427 6556 713 6564
rect 947 6556 1093 6564
rect 1467 6556 1493 6564
rect 1947 6556 2213 6564
rect 2667 6556 2953 6564
rect 3027 6556 3913 6564
rect 4087 6556 4213 6564
rect 4307 6556 4353 6564
rect 4527 6556 4724 6564
rect 547 6536 573 6544
rect 707 6536 1113 6544
rect 2027 6536 2153 6544
rect 2287 6536 2813 6544
rect 2947 6536 3653 6544
rect 3927 6536 3973 6544
rect 4147 6536 4653 6544
rect 4716 6544 4724 6556
rect 4747 6556 4793 6564
rect 4927 6556 5093 6564
rect 5127 6556 5213 6564
rect 5287 6556 6153 6564
rect 6387 6556 6433 6564
rect 6527 6556 6613 6564
rect 6827 6556 6933 6564
rect 6947 6556 7053 6564
rect 7856 6564 7864 6576
rect 7907 6576 7953 6584
rect 8007 6576 8053 6584
rect 8107 6576 8153 6584
rect 8467 6576 8573 6584
rect 8807 6576 9013 6584
rect 9387 6576 9673 6584
rect 9687 6576 9733 6584
rect 9907 6576 9953 6584
rect 11427 6576 11513 6584
rect 11736 6584 11744 6596
rect 11767 6596 11993 6604
rect 12007 6596 12093 6604
rect 12107 6596 12144 6604
rect 12136 6587 12144 6596
rect 11607 6576 11744 6584
rect 11787 6576 11953 6584
rect 11967 6576 12093 6584
rect 7067 6556 7364 6564
rect 7856 6556 8453 6564
rect 4716 6536 4893 6544
rect 5007 6536 5453 6544
rect 5487 6536 5533 6544
rect 5927 6536 5993 6544
rect 6127 6536 6193 6544
rect 6367 6536 6413 6544
rect 6607 6536 6733 6544
rect 6787 6536 7253 6544
rect 7356 6544 7364 6556
rect 9607 6556 9653 6564
rect 9807 6556 10033 6564
rect 10047 6556 10173 6564
rect 10447 6556 10593 6564
rect 10607 6556 10753 6564
rect 11127 6556 11153 6564
rect 11427 6556 11733 6564
rect 7356 6536 7473 6544
rect 7567 6536 8333 6544
rect 8347 6536 8393 6544
rect 8667 6536 10553 6544
rect 11047 6536 11413 6544
rect 587 6516 953 6524
rect 967 6516 2084 6524
rect 387 6496 893 6504
rect 1687 6496 2053 6504
rect 2076 6504 2084 6516
rect 2727 6516 2833 6524
rect 3047 6516 4733 6524
rect 4847 6516 5713 6524
rect 6207 6516 6553 6524
rect 6767 6516 8853 6524
rect 8867 6516 9393 6524
rect 9407 6516 11453 6524
rect 11467 6516 11553 6524
rect 2076 6496 3653 6504
rect 3727 6496 5333 6504
rect 5467 6496 6393 6504
rect 6447 6496 6813 6504
rect 7376 6496 8593 6504
rect 1627 6476 1813 6484
rect 2327 6476 2513 6484
rect 2527 6476 2793 6484
rect 2887 6476 3473 6484
rect 3507 6476 3553 6484
rect 3707 6476 3853 6484
rect 4027 6476 4073 6484
rect 4267 6476 4573 6484
rect 4607 6476 4673 6484
rect 4747 6476 4993 6484
rect 5047 6476 5093 6484
rect 5187 6476 5353 6484
rect 5407 6476 5773 6484
rect 7376 6484 7384 6496
rect 8607 6496 8913 6504
rect 9007 6496 10784 6504
rect 6167 6476 7384 6484
rect 7467 6476 7813 6484
rect 7847 6476 7913 6484
rect 8387 6476 8413 6484
rect 8687 6476 10473 6484
rect 10776 6484 10784 6496
rect 10776 6476 11793 6484
rect 11807 6476 12013 6484
rect 12027 6476 12173 6484
rect 2147 6456 2233 6464
rect 3667 6456 3753 6464
rect 3767 6456 4113 6464
rect 4367 6456 5953 6464
rect 5967 6456 8213 6464
rect 8887 6456 9253 6464
rect 9287 6456 9393 6464
rect 10807 6456 11533 6464
rect 147 6436 493 6444
rect 2007 6436 2433 6444
rect 2607 6436 3053 6444
rect 3167 6436 3273 6444
rect 3527 6436 3573 6444
rect 3627 6436 3813 6444
rect 3827 6436 4084 6444
rect 27 6416 173 6424
rect 296 6416 313 6424
rect -24 6396 133 6404
rect -24 6356 -16 6396
rect 296 6364 304 6416
rect 1187 6416 1333 6424
rect 1347 6416 1533 6424
rect 1587 6416 1753 6424
rect 2287 6416 2593 6424
rect 2747 6416 3113 6424
rect 3487 6416 3553 6424
rect 3567 6416 4013 6424
rect 4076 6424 4084 6436
rect 4107 6436 5533 6444
rect 5887 6436 6473 6444
rect 6667 6436 6853 6444
rect 6927 6436 6953 6444
rect 7587 6436 7693 6444
rect 7727 6436 7853 6444
rect 8847 6436 9373 6444
rect 9607 6436 10133 6444
rect 10147 6436 10353 6444
rect 10647 6436 10813 6444
rect 10827 6436 10993 6444
rect 11007 6436 11233 6444
rect 11387 6436 11893 6444
rect 4076 6416 4533 6424
rect 4556 6416 4573 6424
rect 4587 6416 4593 6424
rect 4947 6416 4973 6424
rect 5447 6416 5513 6424
rect 6187 6416 6233 6424
rect 6287 6416 6613 6424
rect 6687 6416 6853 6424
rect 6887 6416 7133 6424
rect 7227 6416 7564 6424
rect 327 6396 353 6404
rect 2487 6396 2624 6404
rect 2616 6387 2624 6396
rect 2936 6396 3033 6404
rect 2936 6387 2944 6396
rect 3047 6396 3073 6404
rect 3147 6396 3293 6404
rect 3647 6396 3733 6404
rect 4567 6396 4653 6404
rect 4667 6396 4713 6404
rect 4747 6396 4773 6404
rect 4796 6404 4804 6413
rect 4796 6396 4953 6404
rect 5007 6396 5193 6404
rect 5247 6396 5313 6404
rect 6007 6396 6193 6404
rect 6447 6396 6493 6404
rect 6707 6396 6733 6404
rect 6807 6396 6913 6404
rect 6987 6396 7173 6404
rect 7287 6396 7333 6404
rect 7467 6396 7533 6404
rect 7556 6404 7564 6416
rect 7667 6416 7733 6424
rect 7947 6416 8073 6424
rect 8267 6416 8433 6424
rect 8547 6416 8613 6424
rect 9087 6416 9633 6424
rect 10007 6416 10073 6424
rect 10127 6416 10833 6424
rect 10847 6416 10873 6424
rect 10947 6416 11053 6424
rect 11067 6416 11193 6424
rect 11427 6416 11553 6424
rect 11807 6416 11933 6424
rect 7556 6396 7793 6404
rect 7907 6396 8033 6404
rect 8467 6396 8633 6404
rect 8807 6396 8853 6404
rect 8907 6396 8953 6404
rect 9016 6396 9213 6404
rect 9016 6387 9024 6396
rect 9267 6396 9553 6404
rect 9987 6396 10193 6404
rect 10207 6396 10293 6404
rect 10496 6396 10833 6404
rect 10496 6387 10504 6396
rect 10887 6396 10973 6404
rect 10987 6396 11013 6404
rect 11227 6396 11344 6404
rect 727 6376 1313 6384
rect 1387 6376 1473 6384
rect 1627 6376 2173 6384
rect 2187 6376 2293 6384
rect 2627 6376 2904 6384
rect 296 6356 333 6364
rect 547 6356 733 6364
rect 1407 6356 1833 6364
rect 2687 6356 2793 6364
rect 2896 6364 2904 6376
rect 3067 6376 3613 6384
rect 3667 6376 3873 6384
rect 4207 6376 4313 6384
rect 4327 6376 4413 6384
rect 4447 6376 4484 6384
rect 2896 6356 3433 6364
rect 3487 6356 3533 6364
rect 4227 6356 4253 6364
rect 4427 6356 4453 6364
rect 1707 6336 2333 6344
rect 3107 6336 3273 6344
rect 3567 6336 3673 6344
rect 4476 6344 4484 6376
rect 4547 6376 4613 6384
rect 4667 6376 4753 6384
rect 4907 6376 5153 6384
rect 5307 6376 5433 6384
rect 5567 6376 5804 6384
rect 5087 6356 5233 6364
rect 5287 6356 5333 6364
rect 5587 6356 5753 6364
rect 5796 6364 5804 6376
rect 5827 6376 5973 6384
rect 5987 6376 6273 6384
rect 6387 6376 6713 6384
rect 6827 6376 7113 6384
rect 7567 6376 7613 6384
rect 7647 6376 7713 6384
rect 8227 6376 8273 6384
rect 8627 6376 8773 6384
rect 8787 6376 8973 6384
rect 9247 6376 9273 6384
rect 9767 6376 9793 6384
rect 9947 6376 10093 6384
rect 10547 6376 10653 6384
rect 10867 6376 10933 6384
rect 11007 6376 11193 6384
rect 11336 6384 11344 6396
rect 11367 6396 11393 6404
rect 11447 6396 11513 6404
rect 11527 6396 11573 6404
rect 11867 6396 12004 6404
rect 11336 6376 11713 6384
rect 11767 6376 11873 6384
rect 11996 6384 12004 6396
rect 12027 6396 12113 6404
rect 11996 6376 12133 6384
rect 5796 6356 5893 6364
rect 5947 6356 5973 6364
rect 6247 6356 6353 6364
rect 6467 6356 6873 6364
rect 6887 6356 7544 6364
rect 4047 6336 5333 6344
rect 5647 6336 5733 6344
rect 6567 6336 6593 6344
rect 6607 6336 6813 6344
rect 6867 6336 6953 6344
rect 7327 6336 7473 6344
rect 7536 6344 7544 6356
rect 7607 6356 7733 6364
rect 8107 6356 8233 6364
rect 8767 6356 8793 6364
rect 8827 6356 9213 6364
rect 9787 6356 9913 6364
rect 10967 6356 11033 6364
rect 11547 6356 11853 6364
rect 11867 6356 11893 6364
rect 11916 6347 11924 6373
rect 11947 6356 11973 6364
rect 7536 6336 7833 6344
rect 8847 6336 8873 6344
rect 9107 6336 9333 6344
rect 9347 6336 9613 6344
rect 9627 6336 9973 6344
rect 9987 6336 10253 6344
rect 10267 6336 10273 6344
rect 10287 6336 10353 6344
rect 10667 6336 11153 6344
rect 11687 6336 11753 6344
rect 11787 6336 11813 6344
rect 1787 6316 1813 6324
rect 2187 6316 2773 6324
rect 2907 6316 3013 6324
rect 3327 6316 4093 6324
rect 4327 6316 4453 6324
rect 4747 6316 4973 6324
rect 4987 6316 5573 6324
rect 5587 6316 6873 6324
rect 6887 6316 7153 6324
rect 7167 6316 8553 6324
rect 10667 6316 11093 6324
rect 2967 6296 3633 6304
rect 3687 6296 3833 6304
rect 4047 6296 4373 6304
rect 4727 6296 5393 6304
rect 5707 6296 5993 6304
rect 6147 6296 6393 6304
rect 6447 6296 6753 6304
rect 6847 6296 9433 6304
rect 1827 6276 5633 6284
rect 5647 6276 6193 6284
rect 6287 6276 6593 6284
rect 6627 6276 7133 6284
rect 7267 6276 9533 6284
rect 9547 6276 9713 6284
rect 847 6256 1053 6264
rect 1607 6256 1633 6264
rect 1987 6256 2013 6264
rect 2347 6256 2453 6264
rect 2467 6256 3093 6264
rect 3187 6256 3693 6264
rect 3787 6256 3953 6264
rect 4007 6256 4353 6264
rect 4947 6256 5013 6264
rect 5047 6256 5133 6264
rect 5147 6256 5813 6264
rect 5947 6256 6173 6264
rect 6707 6256 6733 6264
rect 6827 6256 6993 6264
rect 7167 6256 7453 6264
rect 2787 6236 5433 6244
rect 5447 6236 6913 6244
rect 7067 6236 7173 6244
rect 7207 6236 7973 6244
rect 907 6216 1373 6224
rect 2227 6216 3333 6224
rect 3407 6216 3873 6224
rect 3947 6216 4213 6224
rect 4227 6216 4573 6224
rect 4587 6216 4673 6224
rect 4687 6216 4693 6224
rect 4707 6216 5533 6224
rect 5547 6216 7033 6224
rect 7367 6216 7413 6224
rect 8527 6216 8553 6224
rect 3707 6196 4153 6204
rect 4547 6196 4873 6204
rect 5407 6196 5613 6204
rect 5627 6196 6213 6204
rect 6227 6196 6413 6204
rect 6427 6196 7213 6204
rect 7287 6196 7413 6204
rect 1767 6176 1793 6184
rect 1807 6176 1813 6184
rect 1847 6176 2413 6184
rect 3287 6176 4053 6184
rect 4067 6176 4173 6184
rect 4447 6176 5113 6184
rect 5427 6176 5513 6184
rect 5527 6176 5933 6184
rect 6127 6176 6433 6184
rect 6447 6176 6553 6184
rect 6607 6176 7433 6184
rect 7507 6176 8073 6184
rect 8087 6176 8193 6184
rect 467 6156 653 6164
rect 2827 6156 3193 6164
rect 3427 6156 3433 6164
rect 3447 6156 3893 6164
rect 3907 6156 3993 6164
rect 4367 6156 4393 6164
rect 4416 6156 4533 6164
rect 467 6136 513 6144
rect 1047 6136 1173 6144
rect 1687 6136 1793 6144
rect 1807 6136 1984 6144
rect -24 6104 -16 6124
rect 567 6116 973 6124
rect 987 6116 1213 6124
rect 1976 6107 1984 6136
rect 2287 6136 2333 6144
rect 2387 6136 2433 6144
rect 2927 6136 2973 6144
rect 3627 6136 4093 6144
rect 4416 6144 4424 6156
rect 4727 6156 4773 6164
rect 4827 6156 5233 6164
rect 5327 6156 5664 6164
rect 4327 6136 4424 6144
rect 5136 6136 5224 6144
rect 2007 6116 2133 6124
rect 2307 6116 2353 6124
rect 2407 6116 2453 6124
rect 3007 6116 3053 6124
rect 3187 6116 3233 6124
rect 3436 6116 3644 6124
rect -24 6096 1093 6104
rect 1827 6096 1933 6104
rect 2867 6096 3013 6104
rect 3436 6104 3444 6116
rect 3636 6107 3644 6116
rect 3847 6116 3993 6124
rect 4187 6116 4253 6124
rect 4267 6116 4293 6124
rect 4307 6116 4444 6124
rect 3047 6096 3444 6104
rect 3796 6087 3804 6113
rect 3867 6096 4313 6104
rect 4436 6104 4444 6116
rect 4627 6116 4813 6124
rect 4887 6116 4933 6124
rect 5136 6124 5144 6136
rect 5027 6116 5144 6124
rect 5216 6124 5224 6136
rect 5307 6136 5373 6144
rect 5656 6144 5664 6156
rect 5767 6156 5793 6164
rect 6316 6156 6393 6164
rect 5656 6136 5713 6144
rect 5807 6136 6093 6144
rect 6107 6136 6213 6144
rect 6316 6144 6324 6156
rect 6427 6156 6473 6164
rect 6496 6156 6853 6164
rect 6496 6144 6504 6156
rect 7047 6156 7233 6164
rect 7547 6156 7673 6164
rect 7787 6156 7873 6164
rect 7907 6156 8093 6164
rect 8107 6156 8273 6164
rect 8287 6156 8373 6164
rect 8907 6156 9173 6164
rect 9447 6156 9953 6164
rect 9967 6156 10873 6164
rect 10887 6156 11093 6164
rect 11427 6156 11473 6164
rect 6267 6136 6324 6144
rect 6436 6136 6504 6144
rect 5187 6116 5204 6124
rect 5216 6116 5353 6124
rect 4327 6096 4384 6104
rect 4436 6096 4533 6104
rect 1967 6076 2113 6084
rect 2587 6076 2733 6084
rect 2887 6076 2973 6084
rect 2987 6076 3753 6084
rect 4207 6076 4313 6084
rect 4327 6076 4333 6084
rect 4376 6084 4384 6096
rect 4556 6096 4733 6104
rect 4556 6087 4564 6096
rect 4767 6096 4893 6104
rect 5007 6096 5033 6104
rect 5067 6096 5153 6104
rect 5196 6104 5204 6116
rect 5556 6124 5564 6133
rect 6436 6127 6444 6136
rect 6947 6136 7013 6144
rect 7207 6136 7273 6144
rect 7296 6136 7473 6144
rect 5556 6116 5644 6124
rect 5196 6096 5373 6104
rect 5567 6096 5613 6104
rect 5636 6104 5644 6116
rect 5696 6116 5753 6124
rect 5696 6107 5704 6116
rect 6096 6116 6433 6124
rect 5636 6096 5653 6104
rect 5776 6104 5784 6113
rect 6096 6104 6104 6116
rect 6487 6116 6653 6124
rect 6967 6116 6993 6124
rect 7087 6116 7113 6124
rect 7296 6124 7304 6136
rect 7527 6136 7593 6144
rect 7647 6136 7973 6144
rect 8227 6136 8253 6144
rect 8947 6136 9053 6144
rect 9587 6136 9673 6144
rect 9827 6136 10773 6144
rect 10787 6136 11153 6144
rect 11487 6136 11513 6144
rect 11527 6136 11613 6144
rect 11667 6136 11793 6144
rect 11987 6136 12093 6144
rect 7267 6116 7304 6124
rect 7316 6116 7433 6124
rect 5776 6096 6104 6104
rect 6227 6096 6273 6104
rect 6447 6096 6513 6104
rect 6627 6096 6693 6104
rect 6947 6096 6973 6104
rect 4376 6076 4413 6084
rect 5127 6076 5513 6084
rect 5667 6076 5753 6084
rect 6176 6076 6253 6084
rect 3047 6056 3153 6064
rect 3427 6056 3573 6064
rect 3787 6056 3813 6064
rect 3987 6056 3993 6064
rect 4107 6056 4153 6064
rect 4247 6056 4333 6064
rect 4387 6056 5013 6064
rect 5047 6056 5793 6064
rect 6176 6064 6184 6076
rect 6267 6076 6333 6084
rect 6347 6076 6573 6084
rect 6627 6076 6733 6084
rect 6847 6076 6893 6084
rect 7036 6084 7044 6113
rect 7067 6096 7073 6104
rect 7087 6096 7133 6104
rect 7316 6104 7324 6116
rect 7627 6116 7673 6124
rect 7816 6116 8033 6124
rect 7816 6107 7824 6116
rect 8247 6116 8353 6124
rect 8667 6116 8753 6124
rect 8927 6116 8993 6124
rect 9407 6116 9593 6124
rect 9607 6116 9893 6124
rect 10527 6116 10573 6124
rect 11147 6116 11353 6124
rect 11507 6116 11624 6124
rect 7247 6096 7324 6104
rect 7467 6096 7513 6104
rect 7727 6096 7773 6104
rect 7987 6096 8013 6104
rect 8536 6087 8544 6113
rect 9327 6096 9373 6104
rect 9787 6096 9813 6104
rect 9827 6096 9993 6104
rect 10007 6096 10113 6104
rect 10916 6104 10924 6113
rect 10916 6096 11113 6104
rect 11167 6096 11333 6104
rect 11347 6096 11593 6104
rect 11616 6104 11624 6116
rect 11647 6116 11673 6124
rect 11967 6116 12033 6124
rect 11616 6096 11693 6104
rect 11867 6096 11913 6104
rect 11927 6096 12073 6104
rect 7036 6076 7053 6084
rect 7427 6076 7893 6084
rect 8067 6076 8093 6084
rect 9127 6076 9453 6084
rect 9467 6076 9633 6084
rect 9647 6076 9653 6084
rect 10567 6076 10733 6084
rect 10887 6076 10933 6084
rect 10967 6076 10973 6084
rect 10987 6076 11073 6084
rect 11087 6076 11153 6084
rect 11167 6076 11253 6084
rect 11267 6076 11293 6084
rect 11627 6076 11653 6084
rect 5927 6056 6184 6064
rect 6287 6056 6313 6064
rect 7027 6056 9673 6064
rect 9687 6056 10133 6064
rect 10147 6056 10453 6064
rect 10467 6056 10493 6064
rect 11487 6056 11633 6064
rect 1147 6036 3013 6044
rect 3067 6036 3273 6044
rect 3287 6036 5133 6044
rect 5207 6036 5273 6044
rect 5347 6036 6473 6044
rect 6547 6036 6633 6044
rect 6687 6036 6713 6044
rect 6747 6036 7013 6044
rect 7207 6036 7253 6044
rect 7267 6036 7853 6044
rect 8607 6036 9033 6044
rect 9047 6036 9293 6044
rect 9307 6036 9813 6044
rect 11367 6036 11713 6044
rect 2047 6016 2153 6024
rect 3207 6016 4433 6024
rect 4527 6016 4553 6024
rect 4587 6016 4953 6024
rect 5027 6016 5113 6024
rect 5227 6016 5313 6024
rect 5367 6016 5993 6024
rect 6007 6016 6133 6024
rect 6167 6016 6853 6024
rect 6987 6016 9013 6024
rect 9027 6016 9233 6024
rect 9247 6016 11173 6024
rect 11187 6016 11293 6024
rect 2227 5996 2533 6004
rect 2547 5996 2753 6004
rect 3027 5996 3213 6004
rect 3587 5996 4053 6004
rect 4787 5996 5333 6004
rect 5427 5996 6413 6004
rect 6467 5996 6493 6004
rect 6567 5996 6673 6004
rect 6907 5996 7073 6004
rect 7107 5996 7153 6004
rect 7187 5996 7513 6004
rect 8347 5996 8413 6004
rect 8647 5996 8733 6004
rect 10507 5996 10573 6004
rect 10587 5996 10713 6004
rect 10747 5996 11093 6004
rect 987 5976 1093 5984
rect 1407 5976 1513 5984
rect 1827 5976 1993 5984
rect 3067 5976 3493 5984
rect 3527 5976 3613 5984
rect 3767 5976 4913 5984
rect 5107 5976 6133 5984
rect 6187 5976 6293 5984
rect 6547 5976 6933 5984
rect 7156 5976 7493 5984
rect 547 5956 693 5964
rect 707 5956 1033 5964
rect 3407 5956 3653 5964
rect 4187 5956 4253 5964
rect 4547 5956 4853 5964
rect 4927 5956 5593 5964
rect 5607 5956 6733 5964
rect 6767 5956 7093 5964
rect 7156 5964 7164 5976
rect 7647 5976 8113 5984
rect 11467 5976 11513 5984
rect 11607 5976 11893 5984
rect 7107 5956 7164 5964
rect 7367 5956 7393 5964
rect 8747 5956 11493 5964
rect 11507 5956 11673 5964
rect 327 5936 364 5944
rect 307 5916 333 5924
rect 356 5907 364 5936
rect 1647 5936 2353 5944
rect 2447 5936 2473 5944
rect 2767 5936 3233 5944
rect 3467 5936 3853 5944
rect 4047 5936 4573 5944
rect 4807 5936 4833 5944
rect 4847 5936 4933 5944
rect 4947 5936 5133 5944
rect 5207 5936 5353 5944
rect 5387 5936 5533 5944
rect 5947 5936 6033 5944
rect 6147 5936 6373 5944
rect 6607 5936 6793 5944
rect 6827 5936 6953 5944
rect 7187 5936 7353 5944
rect 7367 5936 7433 5944
rect 7727 5936 7833 5944
rect 7847 5936 7873 5944
rect 8187 5936 8393 5944
rect 8787 5936 8873 5944
rect 9187 5936 9433 5944
rect 9447 5936 9533 5944
rect 9727 5936 10253 5944
rect 10547 5936 10573 5944
rect 10687 5936 10713 5944
rect 10727 5936 10873 5944
rect 11107 5936 11133 5944
rect 11207 5936 11553 5944
rect 11727 5936 11813 5944
rect 11827 5936 12053 5944
rect 12067 5936 12073 5944
rect 387 5916 433 5924
rect 667 5916 713 5924
rect 1527 5916 2213 5924
rect 2407 5916 2473 5924
rect 2507 5916 2844 5924
rect 2836 5907 2844 5916
rect 3376 5916 3393 5924
rect 167 5896 313 5904
rect 527 5896 573 5904
rect 867 5896 893 5904
rect 1007 5896 1393 5904
rect 1487 5896 1613 5904
rect 2627 5896 2653 5904
rect 2867 5896 2913 5904
rect 3376 5904 3384 5916
rect 3547 5916 4153 5924
rect 3676 5907 3684 5916
rect 4247 5916 4613 5924
rect 4827 5916 4893 5924
rect 4987 5916 5113 5924
rect 5187 5916 5393 5924
rect 5527 5916 5593 5924
rect 6067 5916 6313 5924
rect 6367 5916 6493 5924
rect 6527 5916 6573 5924
rect 6707 5916 6764 5924
rect 3327 5896 3384 5904
rect 3407 5896 3513 5904
rect 3527 5896 3553 5904
rect 3827 5896 3913 5904
rect 4007 5896 4373 5904
rect 4427 5896 4453 5904
rect 4467 5896 4753 5904
rect 4807 5896 4873 5904
rect 5047 5896 5153 5904
rect 5467 5896 5573 5904
rect 5736 5887 5744 5913
rect 5956 5904 5964 5913
rect 5927 5896 5964 5904
rect 6307 5896 6713 5904
rect 6727 5896 6733 5904
rect 6756 5904 6764 5916
rect 7376 5916 7864 5924
rect 6756 5896 6773 5904
rect 7007 5896 7053 5904
rect 7376 5904 7384 5916
rect 7856 5907 7864 5916
rect 7887 5916 8053 5924
rect 8756 5916 8953 5924
rect 8756 5907 8764 5916
rect 9007 5916 9113 5924
rect 9287 5916 9473 5924
rect 9496 5916 9933 5924
rect 9496 5907 9504 5916
rect 10127 5916 10153 5924
rect 10247 5916 10313 5924
rect 10367 5916 10533 5924
rect 10567 5916 10713 5924
rect 10767 5916 10893 5924
rect 11127 5916 11324 5924
rect 7087 5896 7384 5904
rect 7447 5896 7513 5904
rect 8667 5896 8713 5904
rect 8987 5896 9013 5904
rect 9067 5896 9133 5904
rect 9787 5896 9913 5904
rect 10107 5896 10173 5904
rect 10267 5896 10293 5904
rect 10527 5896 10573 5904
rect 10747 5896 10893 5904
rect 10916 5887 10924 5913
rect 11316 5907 11324 5916
rect 11347 5916 11504 5924
rect 11147 5896 11173 5904
rect 11496 5904 11504 5916
rect 11527 5916 11653 5924
rect 11667 5916 11733 5924
rect 11496 5896 11533 5904
rect 11547 5896 11693 5904
rect 147 5876 433 5884
rect 447 5876 733 5884
rect 1847 5876 2193 5884
rect 2647 5876 3353 5884
rect 3527 5876 3713 5884
rect 3887 5876 3973 5884
rect 4287 5876 4593 5884
rect 4607 5876 4953 5884
rect 5767 5876 5813 5884
rect 5827 5876 5893 5884
rect 5927 5876 6093 5884
rect 6167 5876 6413 5884
rect 6467 5876 7133 5884
rect 7167 5876 7253 5884
rect 7347 5876 7453 5884
rect 7487 5876 7513 5884
rect 7887 5876 7993 5884
rect 8547 5876 8553 5884
rect 8567 5876 8673 5884
rect 9167 5876 9273 5884
rect 9287 5876 9293 5884
rect 9347 5876 9493 5884
rect 9667 5876 9693 5884
rect 9947 5876 10093 5884
rect 11947 5876 12033 5884
rect 12047 5876 12093 5884
rect 67 5856 173 5864
rect 187 5856 473 5864
rect 667 5856 2393 5864
rect 3607 5856 3973 5864
rect 4067 5856 5673 5864
rect 5867 5856 5993 5864
rect 6076 5856 6513 5864
rect 2427 5836 3773 5844
rect 3947 5836 4353 5844
rect 4527 5836 5053 5844
rect 5407 5836 5853 5844
rect 6076 5844 6084 5856
rect 6556 5856 6813 5864
rect 5907 5836 6084 5844
rect 6187 5836 6333 5844
rect 6556 5844 6564 5856
rect 6827 5856 6953 5864
rect 6967 5856 7073 5864
rect 7507 5856 7573 5864
rect 7867 5856 8193 5864
rect 9587 5856 9593 5864
rect 9607 5856 9733 5864
rect 6347 5836 6564 5844
rect 6587 5836 6653 5844
rect 6847 5836 6933 5844
rect 7007 5836 7893 5844
rect 8227 5836 8253 5844
rect 1547 5816 3513 5824
rect 3567 5816 3833 5824
rect 3847 5816 4013 5824
rect 4327 5816 5773 5824
rect 5787 5816 6153 5824
rect 6167 5816 6173 5824
rect 6507 5816 8553 5824
rect 8567 5816 9113 5824
rect 9127 5816 10833 5824
rect 10847 5816 10933 5824
rect 2767 5796 2853 5804
rect 2987 5796 3033 5804
rect 3067 5796 3573 5804
rect 3627 5796 4213 5804
rect 4227 5796 4713 5804
rect 4727 5796 5873 5804
rect 6836 5796 8833 5804
rect 327 5776 413 5784
rect 2247 5776 3993 5784
rect 4007 5776 5273 5784
rect 5407 5776 5753 5784
rect 6836 5784 6844 5796
rect 5867 5776 6844 5784
rect 6867 5776 8353 5784
rect 8367 5776 8953 5784
rect 8967 5776 11473 5784
rect 3387 5756 4233 5764
rect 4367 5756 4653 5764
rect 4947 5756 5013 5764
rect 5447 5756 5573 5764
rect 5687 5756 6073 5764
rect 6107 5756 6233 5764
rect 6247 5756 7213 5764
rect 8167 5756 8373 5764
rect 347 5736 473 5744
rect 487 5736 533 5744
rect 1447 5736 1553 5744
rect 2407 5736 3333 5744
rect 4027 5736 5053 5744
rect 5507 5736 5813 5744
rect 5907 5736 6113 5744
rect 6147 5736 6373 5744
rect 6387 5736 6993 5744
rect 8187 5736 8233 5744
rect 9307 5736 9353 5744
rect 2467 5716 2793 5724
rect 2807 5716 3793 5724
rect 3807 5716 4473 5724
rect 4487 5716 5473 5724
rect 5487 5716 6553 5724
rect 6567 5716 7293 5724
rect 7307 5716 7433 5724
rect 7447 5716 7473 5724
rect 8067 5716 9533 5724
rect 9547 5716 9773 5724
rect 9787 5716 10473 5724
rect 10487 5716 10693 5724
rect 11587 5716 11893 5724
rect 2367 5696 5093 5704
rect 5227 5696 6613 5704
rect 6627 5696 6793 5704
rect 7007 5696 7973 5704
rect 7987 5696 9893 5704
rect 9907 5696 9933 5704
rect 9947 5696 10053 5704
rect 11687 5696 11813 5704
rect 11887 5696 11973 5704
rect 1047 5676 1373 5684
rect 2647 5676 3933 5684
rect 4067 5676 4093 5684
rect 4207 5676 4433 5684
rect 4447 5676 4693 5684
rect 4707 5676 4984 5684
rect 147 5656 633 5664
rect 647 5656 853 5664
rect 907 5656 1313 5664
rect 2287 5656 2433 5664
rect 2507 5656 2633 5664
rect 2687 5656 2733 5664
rect 2747 5656 3013 5664
rect 3027 5656 3113 5664
rect 3747 5656 3773 5664
rect 3936 5656 4133 5664
rect 3936 5647 3944 5656
rect 4147 5656 4473 5664
rect 4487 5656 4773 5664
rect 4827 5656 4953 5664
rect 4976 5664 4984 5676
rect 5127 5676 9153 5684
rect 11727 5676 12013 5684
rect 12027 5676 12073 5684
rect 4976 5656 5893 5664
rect 5987 5656 6153 5664
rect 6247 5656 6333 5664
rect 6767 5656 6913 5664
rect 6927 5656 7373 5664
rect 7567 5656 7613 5664
rect 8087 5656 8173 5664
rect 8507 5656 8573 5664
rect 9007 5656 9093 5664
rect 10507 5656 10893 5664
rect 11327 5656 11493 5664
rect 11547 5656 11593 5664
rect 11607 5656 11853 5664
rect 11947 5656 12033 5664
rect 12047 5656 12093 5664
rect 127 5636 273 5644
rect 287 5636 304 5644
rect 296 5624 304 5636
rect 327 5636 373 5644
rect 867 5636 913 5644
rect 1407 5636 1513 5644
rect 1527 5636 1713 5644
rect 1767 5636 1793 5644
rect 2327 5636 2473 5644
rect 2627 5636 2653 5644
rect 2707 5636 2873 5644
rect 2887 5636 3153 5644
rect 3367 5636 3453 5644
rect 3547 5636 3653 5644
rect 3707 5636 3893 5644
rect 4087 5636 4113 5644
rect 4467 5636 4613 5644
rect 4767 5636 4793 5644
rect 4847 5636 5213 5644
rect 5267 5636 5313 5644
rect 5487 5636 5513 5644
rect 5567 5636 5724 5644
rect 296 5616 393 5624
rect 407 5616 673 5624
rect 687 5616 833 5624
rect 887 5616 1053 5624
rect 1076 5624 1084 5633
rect 1076 5616 1113 5624
rect 1847 5616 1973 5624
rect 1987 5616 2093 5624
rect 2116 5624 2124 5633
rect 2116 5616 2253 5624
rect 2447 5616 2853 5624
rect 3927 5616 4593 5624
rect 5027 5616 5333 5624
rect 5356 5624 5364 5633
rect 5716 5627 5724 5636
rect 5767 5636 5913 5644
rect 5967 5636 6033 5644
rect 6147 5636 6293 5644
rect 6487 5636 6813 5644
rect 7067 5636 7133 5644
rect 7147 5636 7273 5644
rect 7407 5636 7693 5644
rect 8007 5636 8133 5644
rect 8516 5636 8593 5644
rect 8516 5627 8524 5636
rect 8927 5636 9153 5644
rect 9167 5636 9573 5644
rect 10247 5636 10313 5644
rect 10367 5636 10413 5644
rect 10767 5636 10853 5644
rect 10867 5636 11073 5644
rect 11567 5636 11693 5644
rect 11916 5644 11924 5653
rect 11916 5636 12053 5644
rect 5356 5616 5404 5624
rect 787 5596 1133 5604
rect 1907 5596 1933 5604
rect 1947 5596 4013 5604
rect 4267 5596 4373 5604
rect 4687 5596 4793 5604
rect 5067 5596 5224 5604
rect 507 5576 1293 5584
rect 2147 5576 2673 5584
rect 2687 5576 3253 5584
rect 3307 5576 3593 5584
rect 4067 5576 5173 5584
rect 5187 5576 5193 5584
rect 5216 5584 5224 5596
rect 5247 5596 5373 5604
rect 5396 5604 5404 5616
rect 5507 5616 5573 5624
rect 5827 5616 5893 5624
rect 6047 5616 6693 5624
rect 6707 5616 6813 5624
rect 6887 5616 6913 5624
rect 7007 5616 7033 5624
rect 7127 5616 7453 5624
rect 7667 5616 7793 5624
rect 7807 5616 8073 5624
rect 8167 5616 8233 5624
rect 8407 5616 8513 5624
rect 8567 5616 8613 5624
rect 8747 5616 8893 5624
rect 8987 5616 9093 5624
rect 9107 5616 9513 5624
rect 9527 5616 9653 5624
rect 9747 5616 9813 5624
rect 10047 5616 10133 5624
rect 10327 5616 10433 5624
rect 10787 5616 10993 5624
rect 11007 5616 11113 5624
rect 11127 5616 11193 5624
rect 11527 5616 11573 5624
rect 5396 5596 5533 5604
rect 5547 5596 5753 5604
rect 5907 5596 6233 5604
rect 6247 5596 6253 5604
rect 6287 5596 6333 5604
rect 6407 5596 6893 5604
rect 6907 5596 7073 5604
rect 7227 5596 8033 5604
rect 8047 5596 8193 5604
rect 8347 5596 8693 5604
rect 8707 5596 8753 5604
rect 9187 5596 9213 5604
rect 10487 5596 10513 5604
rect 10847 5596 10913 5604
rect 5216 5576 6033 5584
rect 6647 5576 6673 5584
rect 6947 5576 7033 5584
rect 7067 5576 7553 5584
rect 7567 5576 7833 5584
rect 7847 5576 8633 5584
rect 8647 5576 8693 5584
rect 8747 5576 8793 5584
rect 9367 5576 10713 5584
rect 10727 5576 10833 5584
rect 11667 5576 11713 5584
rect 1107 5556 1273 5564
rect 1387 5556 2653 5564
rect 3767 5556 4153 5564
rect 4647 5556 5073 5564
rect 5527 5556 5673 5564
rect 5767 5556 5993 5564
rect 6027 5556 6153 5564
rect 6467 5556 6553 5564
rect 7116 5556 7233 5564
rect 2087 5536 4253 5544
rect 4807 5536 5453 5544
rect 5707 5536 5773 5544
rect 5787 5536 6353 5544
rect 7116 5544 7124 5556
rect 7447 5556 7513 5564
rect 7667 5556 7733 5564
rect 6507 5536 7124 5544
rect 7767 5536 7833 5544
rect 1347 5516 1373 5524
rect 2307 5516 2433 5524
rect 2607 5516 2813 5524
rect 3267 5516 4693 5524
rect 4707 5516 5153 5524
rect 5167 5516 5413 5524
rect 5627 5516 5753 5524
rect 5807 5516 6053 5524
rect 6327 5516 6353 5524
rect 6947 5516 7233 5524
rect 7247 5516 7933 5524
rect 1147 5496 1613 5504
rect 2027 5496 2813 5504
rect 3407 5496 3713 5504
rect 3727 5496 3913 5504
rect 3967 5496 4613 5504
rect 4627 5496 6133 5504
rect 6147 5496 6433 5504
rect 6667 5496 7013 5504
rect 7176 5496 7253 5504
rect 1207 5476 2173 5484
rect 2787 5476 3253 5484
rect 4307 5476 5033 5484
rect 5247 5476 5293 5484
rect 5487 5476 5693 5484
rect 5716 5476 6273 5484
rect 847 5456 913 5464
rect 1807 5456 2033 5464
rect 2627 5456 3004 5464
rect -24 5436 613 5444
rect -24 5396 -16 5436
rect 707 5436 773 5444
rect 816 5427 824 5453
rect 1667 5436 2213 5444
rect 2436 5436 2613 5444
rect 2436 5427 2444 5436
rect 2867 5436 2933 5444
rect 2996 5444 3004 5456
rect 3067 5456 3213 5464
rect 3467 5456 3873 5464
rect 3927 5456 4073 5464
rect 4427 5456 4553 5464
rect 4636 5456 4793 5464
rect 2996 5436 3433 5444
rect 3447 5436 3633 5444
rect 3747 5436 3784 5444
rect 856 5416 973 5424
rect 856 5404 864 5416
rect 1107 5416 1213 5424
rect 1847 5416 2013 5424
rect 2267 5416 2313 5424
rect 2807 5416 2833 5424
rect 2887 5416 3033 5424
rect 3087 5416 3193 5424
rect 3247 5416 3273 5424
rect 3727 5416 3753 5424
rect 3776 5424 3784 5436
rect 4416 5436 4453 5444
rect 3776 5416 3893 5424
rect 3947 5416 4313 5424
rect 4416 5424 4424 5436
rect 4636 5427 4644 5456
rect 4887 5456 5033 5464
rect 5087 5456 5253 5464
rect 5307 5456 5393 5464
rect 5716 5464 5724 5476
rect 7176 5484 7184 5496
rect 7547 5496 8113 5504
rect 9727 5496 9793 5504
rect 10167 5496 10273 5504
rect 6827 5476 7184 5484
rect 7287 5476 7773 5484
rect 8867 5476 9433 5484
rect 9447 5476 9813 5484
rect 9827 5476 10173 5484
rect 10967 5476 11093 5484
rect 12027 5476 12073 5484
rect 5687 5456 5724 5464
rect 5747 5456 5833 5464
rect 5847 5456 6033 5464
rect 6047 5456 6433 5464
rect 6627 5456 6833 5464
rect 6847 5456 6973 5464
rect 7767 5456 7784 5464
rect 4867 5436 4973 5444
rect 5067 5436 5433 5444
rect 4327 5416 4424 5424
rect 4447 5416 4493 5424
rect 787 5396 864 5404
rect 1607 5396 1633 5404
rect 1647 5396 1693 5404
rect 2287 5396 2913 5404
rect 2927 5396 3293 5404
rect 3667 5396 3753 5404
rect 4147 5396 4233 5404
rect 4656 5404 4664 5433
rect 4687 5416 4753 5424
rect 4927 5416 4953 5424
rect 5016 5424 5024 5433
rect 5456 5427 5464 5453
rect 5667 5436 5713 5444
rect 5867 5436 5913 5444
rect 6087 5436 6213 5444
rect 6387 5436 6473 5444
rect 7027 5436 7173 5444
rect 7207 5436 7333 5444
rect 7527 5436 7553 5444
rect 7607 5436 7733 5444
rect 7776 5444 7784 5456
rect 7807 5456 7933 5464
rect 8327 5456 8473 5464
rect 8587 5456 9253 5464
rect 9287 5456 9413 5464
rect 9567 5456 9933 5464
rect 9967 5456 10013 5464
rect 10147 5456 10193 5464
rect 10387 5456 10413 5464
rect 10427 5456 10553 5464
rect 10567 5456 10773 5464
rect 10807 5456 10953 5464
rect 11167 5456 11253 5464
rect 11387 5456 11473 5464
rect 11667 5456 11893 5464
rect 7776 5436 7913 5444
rect 7987 5436 8073 5444
rect 8847 5436 8993 5444
rect 9047 5436 9353 5444
rect 9807 5436 9953 5444
rect 10007 5436 10053 5444
rect 10087 5436 10153 5444
rect 10167 5436 10233 5444
rect 10527 5436 10593 5444
rect 10707 5436 10793 5444
rect 10847 5436 11113 5444
rect 5016 5416 5033 5424
rect 5147 5416 5213 5424
rect 5267 5416 5313 5424
rect 5507 5416 5633 5424
rect 5707 5416 5833 5424
rect 5947 5416 6053 5424
rect 6327 5416 6413 5424
rect 6427 5416 6493 5424
rect 6867 5416 6993 5424
rect 7587 5416 7813 5424
rect 8136 5424 8144 5433
rect 7967 5416 8293 5424
rect 8767 5416 8813 5424
rect 8947 5416 9013 5424
rect 9376 5424 9384 5433
rect 11136 5427 11144 5453
rect 11207 5436 11213 5444
rect 11227 5436 11373 5444
rect 11407 5436 11553 5444
rect 12067 5436 12133 5444
rect 9347 5416 9384 5424
rect 9727 5416 9773 5424
rect 9947 5416 9973 5424
rect 10047 5416 10173 5424
rect 10187 5416 10393 5424
rect 10547 5416 10573 5424
rect 10747 5416 10773 5424
rect 10827 5416 10853 5424
rect 11287 5416 11353 5424
rect 11547 5416 11633 5424
rect 11747 5416 11913 5424
rect 11967 5416 12013 5424
rect 4507 5396 4664 5404
rect 4767 5396 5413 5404
rect 5467 5396 5873 5404
rect 5927 5396 6144 5404
rect 1007 5376 1853 5384
rect 1887 5376 1993 5384
rect 2007 5376 2273 5384
rect 2587 5376 2913 5384
rect 2947 5376 3193 5384
rect 3607 5376 3633 5384
rect 4787 5376 4873 5384
rect 4987 5376 6113 5384
rect 6136 5384 6144 5396
rect 6267 5396 6373 5404
rect 6487 5396 6533 5404
rect 6707 5396 6853 5404
rect 7367 5396 7793 5404
rect 8227 5396 8393 5404
rect 8407 5396 8453 5404
rect 8687 5396 8973 5404
rect 9267 5396 9393 5404
rect 9627 5396 9713 5404
rect 10616 5404 10624 5413
rect 10067 5396 10633 5404
rect 10987 5396 11013 5404
rect 11027 5396 11173 5404
rect 11467 5396 11493 5404
rect 11507 5396 11573 5404
rect 6136 5376 6633 5384
rect 7267 5376 7313 5384
rect 7687 5376 7813 5384
rect 8087 5376 8313 5384
rect 9587 5376 9733 5384
rect 1487 5356 1813 5364
rect 3027 5356 3053 5364
rect 3227 5356 5293 5364
rect 5327 5356 5693 5364
rect 5847 5356 6673 5364
rect 6687 5356 6893 5364
rect 7387 5356 7493 5364
rect 9367 5356 11553 5364
rect 11567 5356 11613 5364
rect 1687 5336 1973 5344
rect 2987 5336 3013 5344
rect 3327 5336 5353 5344
rect 5427 5336 7113 5344
rect 7127 5336 7213 5344
rect 3447 5316 3533 5324
rect 3567 5316 3673 5324
rect 4707 5316 9193 5324
rect 9207 5316 9333 5324
rect 9347 5316 9393 5324
rect 767 5296 1033 5304
rect 1047 5296 1233 5304
rect 3447 5296 3853 5304
rect 3927 5296 4193 5304
rect 5427 5296 5513 5304
rect 5627 5296 5713 5304
rect 6127 5296 8633 5304
rect 8647 5296 8773 5304
rect 2907 5276 4093 5284
rect 4127 5276 4933 5284
rect 5787 5276 5853 5284
rect 5987 5276 6793 5284
rect 6827 5276 7633 5284
rect 8207 5276 8293 5284
rect 2727 5256 3233 5264
rect 3807 5256 4673 5264
rect 5167 5256 5653 5264
rect 5667 5256 5773 5264
rect 6087 5256 6573 5264
rect 6587 5256 6673 5264
rect 6727 5256 6833 5264
rect 6847 5256 7853 5264
rect 8227 5256 11273 5264
rect 5367 5236 5973 5244
rect 6007 5236 7073 5244
rect 7087 5236 7093 5244
rect 7347 5236 9013 5244
rect 9027 5236 9573 5244
rect 11727 5236 11813 5244
rect 11827 5236 11873 5244
rect 1407 5216 1433 5224
rect 1447 5216 1713 5224
rect 2107 5216 2613 5224
rect 3107 5216 3593 5224
rect 5307 5216 5873 5224
rect 6367 5216 7333 5224
rect 7387 5216 8933 5224
rect 10147 5216 10193 5224
rect 267 5196 313 5204
rect 656 5204 664 5213
rect 656 5196 793 5204
rect 1307 5196 1333 5204
rect 1347 5196 1373 5204
rect 1547 5196 1653 5204
rect 2327 5196 2793 5204
rect 2907 5196 3833 5204
rect 3887 5196 4753 5204
rect 4767 5196 5033 5204
rect 5167 5196 5693 5204
rect 6127 5196 6713 5204
rect 8507 5196 8593 5204
rect 8987 5196 9353 5204
rect 9967 5196 10153 5204
rect 11627 5196 11653 5204
rect 307 5176 513 5184
rect 527 5176 573 5184
rect 607 5176 713 5184
rect 1487 5176 1513 5184
rect 1747 5176 2033 5184
rect 2047 5176 2133 5184
rect 2147 5176 2193 5184
rect 3307 5176 3353 5184
rect 3487 5176 3693 5184
rect 3947 5176 3993 5184
rect 4007 5176 4073 5184
rect 4527 5176 4613 5184
rect 4967 5176 5313 5184
rect 267 5156 324 5164
rect 136 5144 144 5153
rect 316 5147 324 5156
rect 347 5156 493 5164
rect 647 5156 793 5164
rect 927 5156 1093 5164
rect 1387 5156 1533 5164
rect 1767 5156 1833 5164
rect 2367 5156 2513 5164
rect 3076 5147 3084 5173
rect 5116 5167 5124 5176
rect 5387 5176 5533 5184
rect 5707 5176 5833 5184
rect 6447 5176 6513 5184
rect 6527 5176 6593 5184
rect 7167 5176 7293 5184
rect 7807 5176 7973 5184
rect 7987 5176 8273 5184
rect 8287 5176 8533 5184
rect 8647 5176 8873 5184
rect 9147 5176 9213 5184
rect 9756 5176 10113 5184
rect 9756 5167 9764 5176
rect 10127 5176 10373 5184
rect 10427 5176 10693 5184
rect 10747 5176 10784 5184
rect 10776 5167 10784 5176
rect 10927 5176 11213 5184
rect 11307 5176 11344 5184
rect 3327 5156 3473 5164
rect 3527 5156 3553 5164
rect 3667 5156 3693 5164
rect 3747 5156 3913 5164
rect 3927 5156 3953 5164
rect 4227 5156 4293 5164
rect 4467 5156 4573 5164
rect 4667 5156 4793 5164
rect 5347 5156 5444 5164
rect 136 5136 273 5144
rect 467 5136 713 5144
rect 1227 5136 1353 5144
rect 1447 5136 1693 5144
rect 1747 5136 1793 5144
rect 1987 5136 2033 5144
rect 2187 5136 2293 5144
rect 2687 5136 2873 5144
rect 3147 5136 3293 5144
rect 3347 5136 3433 5144
rect 3607 5136 3673 5144
rect 4147 5136 4193 5144
rect 4447 5136 4493 5144
rect 4607 5136 4693 5144
rect 4727 5136 4773 5144
rect 4827 5136 5173 5144
rect 5187 5136 5193 5144
rect 5436 5144 5444 5156
rect 5467 5156 5513 5164
rect 5607 5156 5833 5164
rect 6287 5156 6633 5164
rect 6807 5156 6933 5164
rect 7007 5156 7113 5164
rect 7767 5156 7913 5164
rect 8627 5156 8793 5164
rect 8847 5156 8893 5164
rect 9007 5156 9173 5164
rect 9327 5156 9373 5164
rect 9607 5156 9633 5164
rect 9807 5156 10073 5164
rect 10387 5156 10433 5164
rect 10447 5156 10733 5164
rect 11107 5156 11153 5164
rect 11287 5156 11313 5164
rect 11336 5164 11344 5176
rect 11387 5176 11473 5184
rect 11927 5176 11953 5184
rect 11336 5156 11693 5164
rect 11927 5156 12073 5164
rect 5436 5136 5673 5144
rect 5727 5136 6053 5144
rect 6267 5136 6353 5144
rect 6667 5136 6873 5144
rect 6896 5136 6953 5144
rect 47 5116 113 5124
rect 127 5116 473 5124
rect 647 5116 693 5124
rect 736 5116 813 5124
rect 736 5104 744 5116
rect 827 5116 1313 5124
rect 1327 5116 1373 5124
rect 1387 5116 1573 5124
rect 1607 5116 1933 5124
rect 1947 5116 2093 5124
rect 2547 5116 2693 5124
rect 2947 5116 3493 5124
rect 3647 5116 3673 5124
rect 3727 5116 3793 5124
rect 3827 5116 3873 5124
rect 4207 5116 4533 5124
rect 4807 5116 4933 5124
rect 5547 5116 5893 5124
rect 6047 5116 6093 5124
rect 6896 5124 6904 5136
rect 6967 5136 7273 5144
rect 7467 5136 7933 5144
rect 8407 5136 8433 5144
rect 9187 5136 9553 5144
rect 9627 5136 10353 5144
rect 10607 5136 10633 5144
rect 10987 5136 11013 5144
rect 11367 5136 11893 5144
rect 11967 5136 12053 5144
rect 6456 5116 6904 5124
rect 687 5096 744 5104
rect 1567 5096 1853 5104
rect 1867 5096 1953 5104
rect 3287 5096 3413 5104
rect 3767 5096 3793 5104
rect 4067 5096 4893 5104
rect 4907 5096 5233 5104
rect 5647 5096 5813 5104
rect 6456 5104 6464 5116
rect 6927 5116 6993 5124
rect 8287 5116 8373 5124
rect 8907 5116 9773 5124
rect 9827 5116 10033 5124
rect 11007 5116 11173 5124
rect 11187 5116 11473 5124
rect 5827 5096 6464 5104
rect 6647 5096 6693 5104
rect 7647 5096 9573 5104
rect 9647 5096 10953 5104
rect 787 5076 873 5084
rect 916 5076 2333 5084
rect 187 5056 433 5064
rect 916 5064 924 5076
rect 2347 5076 3133 5084
rect 4427 5076 4453 5084
rect 4687 5076 5353 5084
rect 5367 5076 5913 5084
rect 6067 5076 6153 5084
rect 7507 5076 7733 5084
rect 8127 5076 8333 5084
rect 8447 5076 8553 5084
rect 447 5056 924 5064
rect 947 5056 4533 5064
rect 4567 5056 6853 5064
rect 7567 5056 7833 5064
rect 7887 5056 8053 5064
rect 8087 5056 8733 5064
rect 8967 5056 10333 5064
rect 687 5036 1773 5044
rect 1787 5036 2153 5044
rect 2767 5036 3213 5044
rect 3647 5036 3653 5044
rect 3667 5036 4393 5044
rect 4547 5036 5613 5044
rect 5927 5036 6093 5044
rect 6507 5036 6693 5044
rect 7667 5036 8033 5044
rect 10187 5036 10333 5044
rect 11147 5036 11193 5044
rect 11887 5036 11913 5044
rect 1247 5016 1533 5024
rect 1587 5016 2653 5024
rect 2667 5016 2733 5024
rect 2767 5016 4553 5024
rect 4707 5016 4733 5024
rect 5307 5016 6013 5024
rect 6027 5016 6433 5024
rect 6647 5016 7053 5024
rect 7147 5016 7433 5024
rect 7447 5016 7573 5024
rect 8307 5016 8953 5024
rect 9207 5016 10813 5024
rect 10827 5016 11113 5024
rect 11127 5016 11133 5024
rect 927 4996 1253 5004
rect 1307 4996 1613 5004
rect 1967 4996 2933 5004
rect 4067 4996 4173 5004
rect 4287 4996 4513 5004
rect 4587 4996 5533 5004
rect 5547 4996 5653 5004
rect 5667 4996 6453 5004
rect 6467 4996 6553 5004
rect 6567 4996 6913 5004
rect 6927 4996 7153 5004
rect 7487 4996 7513 5004
rect 7947 4996 8253 5004
rect 8267 4996 8453 5004
rect 8467 4996 8493 5004
rect 8507 4996 9313 5004
rect 9327 4996 9333 5004
rect 9987 4996 10313 5004
rect 10327 4996 10533 5004
rect 10607 4996 10973 5004
rect 11527 4996 11553 5004
rect 11567 4996 11673 5004
rect 727 4976 893 4984
rect 907 4976 1233 4984
rect 1367 4976 1453 4984
rect 2267 4976 2693 4984
rect 2827 4976 3073 4984
rect 3127 4976 3233 4984
rect 3247 4976 3733 4984
rect 4147 4976 4413 4984
rect 4427 4976 4573 4984
rect 5087 4976 5153 4984
rect 5947 4976 6053 4984
rect 6107 4976 6353 4984
rect 6767 4976 7193 4984
rect 7467 4976 7613 4984
rect 7807 4976 8133 4984
rect 8687 4976 8813 4984
rect 9527 4976 9613 4984
rect 10067 4976 10193 4984
rect 10227 4976 10393 4984
rect 10567 4976 10593 4984
rect 10756 4976 10933 4984
rect -24 4956 133 4964
rect -24 4916 -16 4956
rect 567 4956 673 4964
rect 1027 4956 1053 4964
rect 1107 4956 1113 4964
rect 1127 4956 1133 4964
rect 1207 4956 1433 4964
rect 1687 4956 1853 4964
rect 1987 4956 3273 4964
rect 3667 4956 3773 4964
rect 3787 4956 3853 4964
rect 3907 4956 3973 4964
rect 3987 4956 4213 4964
rect 4267 4956 4373 4964
rect 5047 4956 5073 4964
rect 5227 4956 5253 4964
rect 5447 4956 5473 4964
rect 127 4936 313 4944
rect 516 4944 524 4953
rect 516 4936 893 4944
rect 1287 4936 1353 4944
rect 1607 4936 1633 4944
rect 2087 4936 2133 4944
rect 2727 4936 2873 4944
rect 3227 4936 3253 4944
rect 3656 4944 3664 4953
rect 5496 4947 5504 4973
rect 5527 4956 5793 4964
rect 5847 4956 5873 4964
rect 6547 4956 6573 4964
rect 6967 4956 6993 4964
rect 7387 4956 7453 4964
rect 8127 4956 8253 4964
rect 8316 4956 8373 4964
rect 8316 4947 8324 4956
rect 8416 4956 8473 4964
rect 8416 4947 8424 4956
rect 8707 4956 9233 4964
rect 9827 4956 9993 4964
rect 10047 4956 10553 4964
rect 3467 4936 3664 4944
rect 3847 4936 3993 4944
rect 4167 4936 4273 4944
rect 4407 4936 4553 4944
rect 4567 4936 4833 4944
rect 4907 4936 5053 4944
rect 5147 4936 5273 4944
rect 5607 4936 5673 4944
rect 6047 4936 6073 4944
rect 6247 4936 6553 4944
rect 6867 4936 6893 4944
rect 6947 4936 7104 4944
rect 307 4916 453 4924
rect 487 4916 533 4924
rect 1327 4916 1493 4924
rect 2067 4916 2153 4924
rect 2747 4916 2893 4924
rect 2927 4916 3093 4924
rect 3107 4916 3713 4924
rect 3827 4916 4133 4924
rect 4227 4916 4424 4924
rect 187 4896 333 4904
rect 347 4896 693 4904
rect 707 4896 1113 4904
rect 1147 4896 1433 4904
rect 2007 4896 2093 4904
rect 2687 4896 2813 4904
rect 2847 4896 2953 4904
rect 3847 4896 3933 4904
rect 4027 4896 4113 4904
rect 4187 4896 4233 4904
rect 4347 4896 4393 4904
rect 4416 4904 4424 4916
rect 5107 4916 5493 4924
rect 5967 4916 6033 4924
rect 6347 4916 6593 4924
rect 7047 4916 7073 4924
rect 7096 4924 7104 4936
rect 7127 4936 7173 4944
rect 7287 4936 7433 4944
rect 7487 4936 7513 4944
rect 8167 4936 8213 4944
rect 8436 4936 8993 4944
rect 7096 4916 7413 4924
rect 8436 4924 8444 4936
rect 9547 4936 9633 4944
rect 9667 4936 9853 4944
rect 9907 4936 10213 4944
rect 10367 4936 10493 4944
rect 8387 4916 8444 4924
rect 8547 4916 8833 4924
rect 8847 4916 8853 4924
rect 8947 4916 9153 4924
rect 9987 4916 10053 4924
rect 10187 4916 10293 4924
rect 10307 4916 10333 4924
rect 10736 4924 10744 4953
rect 10756 4947 10764 4976
rect 11027 4976 11093 4984
rect 11407 4976 11493 4984
rect 11507 4976 11533 4984
rect 11796 4976 11873 4984
rect 11187 4956 11233 4964
rect 11547 4956 11653 4964
rect 11796 4964 11804 4976
rect 11887 4976 12113 4984
rect 11667 4956 11804 4964
rect 10736 4916 10753 4924
rect 4416 4896 5733 4904
rect 6127 4896 6413 4904
rect 6907 4896 7253 4904
rect 9027 4896 9653 4904
rect 10247 4896 10573 4904
rect 10776 4904 10784 4953
rect 10807 4936 10953 4944
rect 11107 4936 11153 4944
rect 11467 4936 11513 4944
rect 11647 4936 11653 4944
rect 11667 4936 11713 4944
rect 12027 4936 12053 4944
rect 11747 4916 11813 4924
rect 11907 4916 11913 4924
rect 11927 4916 12033 4924
rect 10587 4896 10784 4904
rect 11827 4896 12073 4904
rect 1007 4876 3173 4884
rect 3187 4876 6513 4884
rect 9167 4876 9293 4884
rect 467 4856 1973 4864
rect 2527 4856 2853 4864
rect 2867 4856 2893 4864
rect 3527 4856 4233 4864
rect 4307 4856 4633 4864
rect 5047 4856 5093 4864
rect 5627 4856 5833 4864
rect 5907 4856 5973 4864
rect 6307 4856 6773 4864
rect 6787 4856 7093 4864
rect 7107 4856 8413 4864
rect 8427 4856 8433 4864
rect 8867 4856 9673 4864
rect 9687 4856 9913 4864
rect 3427 4836 4693 4844
rect 5327 4836 5393 4844
rect 5407 4836 6113 4844
rect 6147 4836 6713 4844
rect 4147 4816 5213 4824
rect 5587 4816 5653 4824
rect 5767 4816 6273 4824
rect 7447 4816 7453 4824
rect 1887 4796 2013 4804
rect 2027 4796 2433 4804
rect 3747 4796 4973 4804
rect 10287 4796 10533 4804
rect 10547 4796 10613 4804
rect 3327 4776 4953 4784
rect 5087 4776 6253 4784
rect 8127 4776 8513 4784
rect 8747 4776 11853 4784
rect 3147 4756 4433 4764
rect 4687 4756 5413 4764
rect 5747 4756 7533 4764
rect 7816 4764 7824 4773
rect 7547 4756 8133 4764
rect 9667 4756 10853 4764
rect 11367 4756 11893 4764
rect 1087 4736 1553 4744
rect 1967 4736 2293 4744
rect 4107 4736 4333 4744
rect 6107 4736 9793 4744
rect 9807 4736 10373 4744
rect 10487 4736 11613 4744
rect 11627 4736 11873 4744
rect 847 4716 893 4724
rect 1447 4716 2353 4724
rect 2367 4716 2473 4724
rect 3187 4716 3333 4724
rect 3347 4716 3653 4724
rect 3767 4716 4213 4724
rect 4227 4716 4813 4724
rect 5007 4716 5333 4724
rect 6347 4716 6533 4724
rect 6547 4716 6633 4724
rect 6967 4716 7953 4724
rect 8187 4716 8193 4724
rect 8207 4716 8873 4724
rect 9207 4716 9453 4724
rect 9467 4716 9713 4724
rect 9727 4716 9833 4724
rect 10007 4716 10433 4724
rect 10447 4716 10964 4724
rect 727 4696 773 4704
rect 787 4696 1033 4704
rect 1247 4696 2153 4704
rect 2167 4696 2213 4704
rect 2867 4696 3073 4704
rect 3207 4696 3493 4704
rect 3507 4696 3893 4704
rect 3916 4696 4124 4704
rect 336 4676 513 4684
rect 336 4664 344 4676
rect 1887 4676 2073 4684
rect 2327 4676 2493 4684
rect 2556 4684 2564 4693
rect 3916 4687 3924 4696
rect 2556 4676 2693 4684
rect 2727 4676 2913 4684
rect 3067 4676 3213 4684
rect 3967 4676 4093 4684
rect 4116 4684 4124 4696
rect 4207 4696 4473 4704
rect 4487 4696 4833 4704
rect 5227 4696 5293 4704
rect 5587 4696 5764 4704
rect 5756 4687 5764 4696
rect 5947 4696 6093 4704
rect 6147 4696 6213 4704
rect 6227 4696 6293 4704
rect 6567 4696 6633 4704
rect 6687 4696 6844 4704
rect 6836 4687 6844 4696
rect 6867 4696 6913 4704
rect 7167 4696 7513 4704
rect 7527 4696 7993 4704
rect 8007 4696 8013 4704
rect 8327 4696 8393 4704
rect 8407 4696 8473 4704
rect 8496 4696 8533 4704
rect 4116 4676 4133 4684
rect 4167 4676 4293 4684
rect 4467 4676 4793 4684
rect 4847 4676 4913 4684
rect 5047 4676 5204 4684
rect 207 4656 344 4664
rect 367 4656 693 4664
rect 1287 4656 1453 4664
rect 1927 4656 2373 4664
rect 2487 4656 3013 4664
rect 3027 4656 3093 4664
rect 3107 4656 3233 4664
rect 3867 4656 4073 4664
rect 4096 4664 4104 4673
rect 5196 4667 5204 4676
rect 5916 4676 5933 4684
rect 5916 4667 5924 4676
rect 7007 4676 7853 4684
rect 7967 4676 8093 4684
rect 8167 4676 8253 4684
rect 8496 4684 8504 4696
rect 8547 4696 8773 4704
rect 9267 4696 9413 4704
rect 10307 4696 10393 4704
rect 10807 4696 10933 4704
rect 10956 4704 10964 4716
rect 11287 4716 11613 4724
rect 10956 4696 11664 4704
rect 8387 4676 8504 4684
rect 8527 4676 8693 4684
rect 9447 4676 9613 4684
rect 9667 4676 9693 4684
rect 9827 4676 10033 4684
rect 10147 4676 10193 4684
rect 10467 4676 11053 4684
rect 11227 4676 11313 4684
rect 11527 4676 11644 4684
rect 11636 4667 11644 4676
rect 4096 4656 4133 4664
rect 4147 4656 4193 4664
rect 4787 4656 4853 4664
rect 4967 4656 5013 4664
rect 5307 4656 5373 4664
rect 5387 4656 5593 4664
rect 5967 4656 5973 4664
rect 5987 4656 6473 4664
rect 6487 4656 6593 4664
rect 7147 4656 7473 4664
rect 8947 4656 9053 4664
rect 9067 4656 9233 4664
rect 9247 4656 9353 4664
rect 9607 4656 9633 4664
rect 9687 4656 9713 4664
rect 9727 4656 9973 4664
rect 10267 4656 10413 4664
rect 11147 4656 11293 4664
rect 11656 4664 11664 4696
rect 11827 4696 11853 4704
rect 12027 4696 12053 4704
rect 11747 4676 12073 4684
rect 11656 4656 11673 4664
rect 11696 4664 11704 4673
rect 11696 4656 11913 4664
rect 87 4636 173 4644
rect 547 4636 833 4644
rect 1707 4636 2133 4644
rect 2427 4636 2473 4644
rect 3627 4636 3733 4644
rect 4087 4636 4173 4644
rect 4667 4636 4733 4644
rect 4827 4636 4893 4644
rect 5067 4636 5393 4644
rect 5807 4636 5933 4644
rect 5947 4636 6053 4644
rect 6407 4636 7173 4644
rect 7187 4636 7633 4644
rect 7647 4636 7653 4644
rect 8767 4636 8773 4644
rect 8787 4636 9093 4644
rect 9207 4636 9273 4644
rect 10547 4636 10573 4644
rect 11407 4636 11453 4644
rect 11827 4636 11873 4644
rect 167 4616 193 4624
rect 827 4616 1013 4624
rect 1027 4616 1413 4624
rect 1427 4616 1913 4624
rect 2127 4616 2333 4624
rect 2427 4616 2773 4624
rect 4047 4616 4093 4624
rect 4127 4616 4413 4624
rect 4927 4616 4993 4624
rect 5267 4616 5413 4624
rect 5427 4616 5893 4624
rect 5976 4616 6553 4624
rect 1667 4596 2233 4604
rect 2247 4596 2533 4604
rect 2547 4596 3053 4604
rect 3067 4596 3133 4604
rect 3167 4596 3273 4604
rect 3747 4596 3833 4604
rect 5976 4604 5984 4616
rect 6567 4616 8053 4624
rect 8067 4616 8433 4624
rect 8507 4616 9073 4624
rect 9707 4616 10793 4624
rect 10967 4616 11233 4624
rect 11247 4616 11853 4624
rect 5167 4596 5984 4604
rect 7147 4596 7353 4604
rect 1127 4576 1253 4584
rect 1647 4576 1933 4584
rect 1947 4576 2513 4584
rect 2527 4576 2853 4584
rect 2967 4576 3613 4584
rect 4347 4576 5033 4584
rect 5767 4576 5813 4584
rect 5827 4576 5953 4584
rect 6987 4576 7433 4584
rect 7707 4576 8193 4584
rect 10507 4576 11093 4584
rect 11107 4576 11333 4584
rect 587 4556 953 4564
rect 967 4556 1313 4564
rect 1807 4556 2053 4564
rect 2067 4556 2713 4564
rect 6327 4556 6733 4564
rect 6747 4556 7693 4564
rect 7807 4556 7833 4564
rect 10227 4556 10553 4564
rect 11147 4556 11353 4564
rect 1027 4536 1393 4544
rect 1407 4536 1433 4544
rect 2087 4536 2133 4544
rect 2147 4536 2453 4544
rect 2947 4536 3113 4544
rect 3347 4536 4173 4544
rect 5367 4536 5713 4544
rect 5947 4536 6193 4544
rect 6507 4536 6913 4544
rect 6927 4536 7253 4544
rect 7327 4536 8473 4544
rect 10987 4536 11533 4544
rect 607 4516 1524 4524
rect 507 4496 1013 4504
rect 1127 4496 1213 4504
rect 1516 4504 1524 4516
rect 1907 4516 2333 4524
rect 2367 4516 2533 4524
rect 2967 4516 2993 4524
rect 3167 4516 3473 4524
rect 5467 4516 5533 4524
rect 5727 4516 6073 4524
rect 6127 4516 6393 4524
rect 7127 4516 7833 4524
rect 7867 4516 7893 4524
rect 7907 4516 8313 4524
rect 8467 4516 8513 4524
rect 8527 4516 8533 4524
rect 9127 4516 10184 4524
rect 1516 4496 3644 4504
rect 587 4476 633 4484
rect 1407 4476 2073 4484
rect 2187 4476 2293 4484
rect 2307 4476 2673 4484
rect 2687 4476 2784 4484
rect 467 4456 533 4464
rect 887 4456 893 4464
rect 907 4456 1413 4464
rect 1427 4456 1653 4464
rect 1707 4456 1773 4464
rect 2167 4456 2553 4464
rect 2567 4456 2733 4464
rect 2776 4464 2784 4476
rect 2807 4476 2973 4484
rect 3636 4484 3644 4496
rect 3667 4496 3813 4504
rect 3827 4496 3933 4504
rect 4007 4496 4153 4504
rect 4247 4496 4633 4504
rect 4647 4496 4813 4504
rect 5227 4496 5533 4504
rect 5567 4496 5733 4504
rect 5747 4496 5793 4504
rect 5987 4496 6233 4504
rect 7027 4496 7093 4504
rect 7207 4496 7653 4504
rect 7867 4496 8033 4504
rect 8367 4496 8393 4504
rect 9447 4496 9773 4504
rect 10027 4496 10153 4504
rect 10176 4504 10184 4516
rect 10787 4516 11553 4524
rect 11567 4516 11673 4524
rect 10176 4496 11193 4504
rect 11207 4496 11713 4504
rect 2987 4476 3124 4484
rect 3636 4476 3753 4484
rect 2776 4456 3093 4464
rect 3116 4464 3124 4476
rect 3767 4476 3773 4484
rect 3847 4476 4233 4484
rect 4247 4476 4293 4484
rect 4327 4476 4424 4484
rect 4416 4467 4424 4476
rect 5487 4476 5513 4484
rect 6107 4476 6133 4484
rect 6367 4476 7144 4484
rect 3116 4456 3213 4464
rect 3947 4456 4124 4464
rect 47 4436 53 4444
rect 67 4436 573 4444
rect 807 4436 973 4444
rect 1067 4436 1513 4444
rect 2727 4436 2833 4444
rect 3007 4436 3133 4444
rect 3807 4436 3973 4444
rect 4116 4444 4124 4456
rect 4147 4456 4193 4464
rect 5147 4456 5173 4464
rect 4116 4436 4213 4444
rect 4227 4436 4253 4444
rect 4687 4436 4733 4444
rect 5196 4444 5204 4473
rect 5787 4456 5873 4464
rect 5967 4456 6573 4464
rect 6767 4456 6933 4464
rect 7047 4456 7113 4464
rect 7136 4464 7144 4476
rect 7227 4476 7293 4484
rect 7527 4476 7573 4484
rect 7676 4484 7684 4493
rect 7627 4476 7684 4484
rect 8247 4476 8373 4484
rect 8427 4476 8733 4484
rect 8827 4476 9053 4484
rect 9327 4476 9593 4484
rect 9607 4476 10333 4484
rect 10607 4476 10753 4484
rect 10847 4476 11153 4484
rect 11327 4476 11513 4484
rect 12007 4476 12093 4484
rect 7136 4456 7313 4464
rect 7387 4456 7493 4464
rect 7807 4456 7873 4464
rect 8347 4456 9033 4464
rect 9087 4456 9113 4464
rect 9267 4456 9413 4464
rect 9467 4456 10024 4464
rect 5187 4436 5204 4444
rect 5927 4436 6113 4444
rect 6147 4436 6253 4444
rect 6267 4436 6413 4444
rect 6627 4436 6693 4444
rect 6707 4436 7073 4444
rect 7287 4436 8213 4444
rect 8747 4436 9273 4444
rect 9287 4436 9513 4444
rect 9947 4436 9993 4444
rect 10016 4444 10024 4456
rect 10387 4456 10413 4464
rect 10627 4456 10773 4464
rect 10827 4456 10853 4464
rect 11007 4456 11053 4464
rect 11147 4456 11173 4464
rect 11227 4456 11373 4464
rect 11736 4456 11893 4464
rect 11736 4447 11744 4456
rect 10016 4436 11213 4444
rect 11407 4436 11573 4444
rect 347 4416 373 4424
rect 867 4416 1053 4424
rect 1636 4424 1644 4433
rect 1067 4416 1644 4424
rect 2567 4416 2613 4424
rect 4107 4416 4253 4424
rect 5147 4416 5373 4424
rect 6167 4416 6213 4424
rect 6607 4416 6773 4424
rect 11627 4416 11913 4424
rect 2647 4396 2973 4404
rect 6407 4396 8073 4404
rect 11547 4396 11773 4404
rect 1607 4376 2313 4384
rect 2327 4376 2633 4384
rect 3887 4376 4493 4384
rect 6267 4376 6893 4384
rect 7407 4376 10653 4384
rect 347 4356 373 4364
rect 2507 4356 4073 4364
rect 6887 4356 7453 4364
rect 1747 4336 1813 4344
rect 2707 4336 2753 4344
rect 4247 4336 5373 4344
rect 1587 4316 1673 4324
rect 1767 4316 4033 4324
rect 4047 4316 6973 4324
rect 107 4296 173 4304
rect 307 4296 393 4304
rect 667 4296 713 4304
rect 6387 4296 7653 4304
rect 367 4276 393 4284
rect 2387 4276 2833 4284
rect 6187 4276 8273 4284
rect 8287 4276 8453 4284
rect 8467 4276 9013 4284
rect 9267 4276 10473 4284
rect 1087 4256 1373 4264
rect 1407 4256 1553 4264
rect 2547 4256 2593 4264
rect 3067 4256 3373 4264
rect 4567 4256 4713 4264
rect 6147 4256 6173 4264
rect 8407 4256 10493 4264
rect 547 4236 613 4244
rect 967 4236 993 4244
rect 1127 4236 1153 4244
rect 1167 4236 1193 4244
rect 1207 4236 1453 4244
rect 2227 4236 2693 4244
rect 2707 4236 3013 4244
rect 3167 4236 3213 4244
rect 6007 4236 6233 4244
rect 6467 4236 6533 4244
rect 8027 4236 8173 4244
rect 8987 4236 9753 4244
rect 10507 4236 10733 4244
rect 10747 4236 12073 4244
rect 12087 4236 12133 4244
rect 1007 4216 1333 4224
rect 1347 4216 1513 4224
rect 1536 4216 1713 4224
rect 1536 4207 1544 4216
rect 2327 4216 2413 4224
rect 2867 4216 3293 4224
rect 3307 4216 3413 4224
rect 3567 4216 3613 4224
rect 3667 4216 3693 4224
rect 4636 4224 4644 4233
rect 4616 4216 4644 4224
rect 4616 4207 4624 4216
rect 5767 4216 5793 4224
rect 5847 4216 5873 4224
rect 6027 4216 6104 4224
rect -24 4184 -16 4204
rect 387 4196 513 4204
rect 747 4196 973 4204
rect 1207 4196 1353 4204
rect 1667 4196 1693 4204
rect 2247 4196 2373 4204
rect 2387 4196 2393 4204
rect 2447 4196 2513 4204
rect 2536 4196 2593 4204
rect -24 4176 133 4184
rect 467 4176 553 4184
rect 567 4176 613 4184
rect 1087 4176 1133 4184
rect 1687 4176 1853 4184
rect 2536 4184 2544 4196
rect 2647 4196 2673 4204
rect 2747 4196 2793 4204
rect 3267 4196 3353 4204
rect 3367 4196 3393 4204
rect 3487 4196 3773 4204
rect 4007 4196 4153 4204
rect 4207 4196 4353 4204
rect 4647 4196 4693 4204
rect 5007 4196 5153 4204
rect 5647 4196 5673 4204
rect 5727 4196 5773 4204
rect 5787 4196 5813 4204
rect 6096 4204 6104 4216
rect 6127 4216 6173 4224
rect 6347 4216 6433 4224
rect 6507 4216 6624 4224
rect 6096 4196 6153 4204
rect 6407 4196 6473 4204
rect 6527 4196 6593 4204
rect 6616 4204 6624 4216
rect 7107 4216 7513 4224
rect 7527 4216 8353 4224
rect 8887 4216 8913 4224
rect 9067 4216 9233 4224
rect 9247 4216 9293 4224
rect 10207 4216 11053 4224
rect 11167 4216 11233 4224
rect 11447 4216 11493 4224
rect 6616 4196 7053 4204
rect 7067 4196 7104 4204
rect 2427 4176 2544 4184
rect 2767 4176 2853 4184
rect 2876 4176 2993 4184
rect 367 4156 393 4164
rect 747 4156 1173 4164
rect 1987 4156 2593 4164
rect 2627 4156 2653 4164
rect 2876 4164 2884 4176
rect 3067 4176 3233 4184
rect 3387 4176 3433 4184
rect 3647 4176 3793 4184
rect 4147 4176 4573 4184
rect 4876 4184 4884 4193
rect 4876 4176 4993 4184
rect 5047 4176 5093 4184
rect 5607 4176 5873 4184
rect 5887 4176 5993 4184
rect 6127 4176 6453 4184
rect 6747 4176 6853 4184
rect 7007 4176 7073 4184
rect 7096 4184 7104 4196
rect 7727 4196 7873 4204
rect 8147 4196 8213 4204
rect 9047 4196 9213 4204
rect 9307 4196 9493 4204
rect 9507 4196 9573 4204
rect 9636 4196 9793 4204
rect 7096 4176 7213 4184
rect 7227 4176 7233 4184
rect 7436 4184 7444 4193
rect 9636 4187 9644 4196
rect 10007 4196 10133 4204
rect 10847 4196 10873 4204
rect 10927 4196 11073 4204
rect 11107 4196 11253 4204
rect 11307 4196 11393 4204
rect 7287 4176 7444 4184
rect 7707 4176 7733 4184
rect 7847 4176 8513 4184
rect 9367 4176 9633 4184
rect 9656 4176 9933 4184
rect 2667 4156 3213 4164
rect 3427 4156 4053 4164
rect 4347 4156 4393 4164
rect 5127 4156 5393 4164
rect 5407 4156 5453 4164
rect 5467 4156 5513 4164
rect 5587 4156 5753 4164
rect 6607 4156 7013 4164
rect 7027 4156 7433 4164
rect 7467 4156 7653 4164
rect 7667 4156 8033 4164
rect 8727 4156 9233 4164
rect 9656 4164 9664 4176
rect 9947 4176 10173 4184
rect 10187 4176 10453 4184
rect 10467 4176 10513 4184
rect 11287 4176 11513 4184
rect 11527 4176 11613 4184
rect 11667 4176 11773 4184
rect 11827 4176 11973 4184
rect 9447 4156 9664 4164
rect 9727 4156 9953 4164
rect 10007 4156 10673 4164
rect 10707 4156 10893 4164
rect 10907 4156 11113 4164
rect 11487 4156 11873 4164
rect 11887 4156 12013 4164
rect 947 4136 993 4144
rect 1967 4136 2353 4144
rect 2367 4136 2453 4144
rect 2467 4136 3173 4144
rect 3187 4136 3193 4144
rect 3407 4136 3493 4144
rect 4287 4136 4333 4144
rect 4747 4136 5213 4144
rect 5707 4136 6013 4144
rect 6447 4136 8013 4144
rect 9467 4136 11473 4144
rect 207 4116 313 4124
rect 2827 4116 3813 4124
rect 3847 4116 4533 4124
rect 4987 4116 5253 4124
rect 6767 4116 6893 4124
rect 6907 4116 7233 4124
rect 9667 4116 9973 4124
rect 9987 4116 10653 4124
rect 10667 4116 11273 4124
rect 1467 4096 2784 4104
rect 307 4076 373 4084
rect 667 4076 713 4084
rect 2776 4084 2784 4096
rect 2807 4096 2933 4104
rect 4427 4096 4573 4104
rect 6207 4096 8373 4104
rect 9207 4096 10313 4104
rect 10587 4096 10813 4104
rect 10827 4096 10993 4104
rect 2776 4076 4404 4084
rect 4396 4064 4404 4076
rect 4987 4076 6953 4084
rect 7227 4076 7473 4084
rect 7487 4076 7613 4084
rect 9827 4076 10113 4084
rect 10127 4076 10653 4084
rect 4396 4056 6633 4064
rect 6707 4056 6873 4064
rect 8907 4056 9393 4064
rect 9487 4056 9753 4064
rect 9767 4056 10693 4064
rect 1527 4036 1913 4044
rect 2167 4036 2573 4044
rect 2667 4036 2773 4044
rect 3647 4036 3973 4044
rect 5267 4036 6053 4044
rect 6067 4036 6393 4044
rect 6507 4036 6673 4044
rect 8707 4036 8813 4044
rect 9707 4036 10153 4044
rect 10547 4036 10593 4044
rect 10667 4036 10753 4044
rect 10767 4036 11253 4044
rect 687 4016 1093 4024
rect 1227 4016 1293 4024
rect 1387 4016 1493 4024
rect 1707 4016 1733 4024
rect 2447 4016 2753 4024
rect 3507 4016 3693 4024
rect 3727 4016 4173 4024
rect 4187 4016 4353 4024
rect 5227 4016 5333 4024
rect 5567 4016 5633 4024
rect 5947 4016 6093 4024
rect 6647 4016 6853 4024
rect 6907 4016 7053 4024
rect 7147 4016 8153 4024
rect 8407 4016 9053 4024
rect 9387 4016 9413 4024
rect 9507 4016 9593 4024
rect 10407 4016 10633 4024
rect 10647 4016 10773 4024
rect 11327 4016 11333 4024
rect 11347 4016 11553 4024
rect 387 3996 473 4004
rect 487 3996 853 4004
rect 867 3996 913 4004
rect 927 3996 1033 4004
rect 1096 3996 1273 4004
rect 467 3976 493 3984
rect 1096 3984 1104 3996
rect 1287 3996 1653 4004
rect 1747 3996 1793 4004
rect 1887 3996 1953 4004
rect 2807 3996 2833 4004
rect 3327 3996 3773 4004
rect 4947 3996 5313 4004
rect 5407 3996 5473 4004
rect 5487 3996 6813 4004
rect 5736 3987 5744 3996
rect 6827 3996 7033 4004
rect 7087 3996 7253 4004
rect 7447 3996 7813 4004
rect 7676 3987 7684 3996
rect 8147 3996 8193 4004
rect 9227 3996 9313 4004
rect 9747 3996 9793 4004
rect 9867 3996 9993 4004
rect 10047 3996 10233 4004
rect 10367 3996 10573 4004
rect 10707 3996 10793 4004
rect 11227 3996 11253 4004
rect 11336 3996 11373 4004
rect 947 3976 1104 3984
rect 1127 3976 1213 3984
rect 1447 3976 1673 3984
rect 1727 3976 1893 3984
rect 2047 3976 2133 3984
rect 2607 3976 2653 3984
rect 2787 3976 3193 3984
rect 3287 3976 3353 3984
rect 3467 3976 3653 3984
rect 3687 3976 3973 3984
rect 4367 3976 4533 3984
rect 4547 3976 4693 3984
rect 4727 3976 4773 3984
rect 4827 3976 5493 3984
rect 5547 3976 5573 3984
rect 5867 3976 6073 3984
rect 6227 3976 6273 3984
rect 6287 3976 6553 3984
rect 6747 3976 6833 3984
rect 6887 3976 6993 3984
rect 7767 3976 7813 3984
rect 8027 3976 8113 3984
rect 8187 3976 8373 3984
rect 8447 3976 8473 3984
rect 8967 3976 9013 3984
rect 9387 3976 9404 3984
rect 67 3956 513 3964
rect 1687 3956 1773 3964
rect 2336 3964 2344 3973
rect 2336 3956 2773 3964
rect 2867 3956 4133 3964
rect 4147 3956 4193 3964
rect 5007 3956 5113 3964
rect 5347 3956 5773 3964
rect 6327 3956 6633 3964
rect 7187 3956 7633 3964
rect 7647 3956 7993 3964
rect 8867 3956 8913 3964
rect 9007 3956 9313 3964
rect 9396 3964 9404 3976
rect 9427 3976 9473 3984
rect 9587 3976 9693 3984
rect 9727 3976 9773 3984
rect 10227 3976 10424 3984
rect 9396 3956 9413 3964
rect 9956 3947 9964 3973
rect 10416 3967 10424 3976
rect 10627 3976 10853 3984
rect 11176 3984 11184 3993
rect 11027 3976 11184 3984
rect 11336 3984 11344 3996
rect 11607 3996 11893 4004
rect 11987 3996 12053 4004
rect 12067 3996 12093 4004
rect 11207 3976 11344 3984
rect 11367 3976 11433 3984
rect 11687 3976 11733 3984
rect 9987 3956 10153 3964
rect 10767 3956 11133 3964
rect 11647 3956 11753 3964
rect 11767 3956 11813 3964
rect 1007 3936 1153 3944
rect 1167 3936 1333 3944
rect 1347 3936 2633 3944
rect 2647 3936 2833 3944
rect 3167 3936 3193 3944
rect 3227 3936 3613 3944
rect 3627 3936 5913 3944
rect 7487 3936 7793 3944
rect 7887 3936 8033 3944
rect 8047 3936 8973 3944
rect 9327 3936 9533 3944
rect 9547 3936 9773 3944
rect 10047 3936 10333 3944
rect 10376 3944 10384 3953
rect 10367 3936 10384 3944
rect 11727 3936 11773 3944
rect 567 3916 1813 3924
rect 1827 3916 1933 3924
rect 2887 3916 3353 3924
rect 3367 3916 3433 3924
rect 3447 3916 3573 3924
rect 3627 3916 3833 3924
rect 5447 3916 6093 3924
rect 9067 3916 9733 3924
rect 10347 3916 10553 3924
rect 10567 3916 10973 3924
rect 187 3896 3413 3904
rect 8027 3896 10173 3904
rect 10367 3896 11673 3904
rect 1027 3876 1833 3884
rect 1847 3876 1993 3884
rect 2207 3876 2513 3884
rect 3467 3876 4153 3884
rect 7227 3876 9193 3884
rect 9367 3876 10693 3884
rect 10707 3876 12033 3884
rect 5067 3856 6393 3864
rect 7847 3856 7933 3864
rect 7947 3856 9413 3864
rect 10807 3856 10933 3864
rect 367 3836 393 3844
rect 1476 3844 1484 3853
rect 407 3836 1593 3844
rect 2267 3836 2473 3844
rect 3087 3836 4913 3844
rect 987 3816 1693 3824
rect 1947 3816 2193 3824
rect 3247 3816 3293 3824
rect 4407 3816 4613 3824
rect 527 3796 1013 3804
rect 1787 3796 2393 3804
rect 2407 3796 2733 3804
rect 8887 3796 11033 3804
rect 11047 3796 11573 3804
rect 11587 3796 11653 3804
rect 727 3776 953 3784
rect 1447 3776 1713 3784
rect 1807 3776 1933 3784
rect 2167 3776 4813 3784
rect 5547 3776 7053 3784
rect 7067 3776 7073 3784
rect 7087 3776 7153 3784
rect 7767 3776 8553 3784
rect 956 3756 1053 3764
rect 956 3747 964 3756
rect 1067 3756 2044 3764
rect 2036 3747 2044 3756
rect 3316 3756 3373 3764
rect 507 3736 533 3744
rect 876 3736 913 3744
rect -24 3704 -16 3724
rect 367 3716 413 3724
rect 876 3724 884 3736
rect 3247 3736 3293 3744
rect 3316 3727 3324 3756
rect 3547 3756 4673 3764
rect 4687 3756 5093 3764
rect 6547 3756 6913 3764
rect 7807 3756 8293 3764
rect 9267 3756 10693 3764
rect 3747 3736 3953 3744
rect 4127 3736 4253 3744
rect 4727 3736 4833 3744
rect 4847 3736 5013 3744
rect 5027 3736 5533 3744
rect 6747 3736 7553 3744
rect 7567 3736 7793 3744
rect 8087 3736 8153 3744
rect 9547 3736 9633 3744
rect 9647 3736 9693 3744
rect 9707 3736 10033 3744
rect 10207 3736 10273 3744
rect 10907 3736 11013 3744
rect 787 3716 884 3724
rect 907 3716 933 3724
rect 1047 3716 1353 3724
rect 1427 3716 2013 3724
rect 2247 3716 2433 3724
rect 2447 3716 2713 3724
rect 3107 3716 3173 3724
rect 3336 3724 3344 3733
rect 3336 3716 3473 3724
rect 3667 3716 3873 3724
rect 4087 3716 4233 3724
rect 4687 3716 4753 3724
rect 6407 3716 7373 3724
rect 7647 3716 7673 3724
rect 7907 3716 7973 3724
rect 8147 3716 8173 3724
rect 8367 3716 8584 3724
rect 8576 3707 8584 3716
rect 8607 3716 8653 3724
rect 8787 3716 8913 3724
rect 9027 3716 9133 3724
rect 9147 3716 9273 3724
rect 9927 3716 9973 3724
rect 9987 3716 10073 3724
rect 10096 3716 10313 3724
rect -24 3696 133 3704
rect 327 3696 533 3704
rect 887 3696 1053 3704
rect 1647 3696 1813 3704
rect 1987 3696 2073 3704
rect 2427 3696 3513 3704
rect 3767 3696 5073 3704
rect 6027 3696 6113 3704
rect 6187 3696 6333 3704
rect 7247 3696 7333 3704
rect 7427 3696 7813 3704
rect 8227 3696 8533 3704
rect 9347 3696 9873 3704
rect 10096 3704 10104 3716
rect 10476 3716 10533 3724
rect 9907 3696 10104 3704
rect 10476 3704 10484 3716
rect 10867 3716 11593 3724
rect 11807 3716 11933 3724
rect 10307 3696 10484 3704
rect 10507 3696 10633 3704
rect 10927 3696 11053 3704
rect 11067 3696 11113 3704
rect 11567 3696 11613 3704
rect 11787 3696 12093 3704
rect 12107 3696 12153 3704
rect 1347 3676 1473 3684
rect 2367 3676 2433 3684
rect 2687 3676 2713 3684
rect 3127 3676 3553 3684
rect 4907 3676 4933 3684
rect 5867 3676 6153 3684
rect 6167 3676 7413 3684
rect 7587 3676 7613 3684
rect 8947 3676 9013 3684
rect 9267 3676 9293 3684
rect 9816 3676 10133 3684
rect 427 3656 873 3664
rect 1187 3656 1373 3664
rect 1587 3656 1653 3664
rect 2227 3656 2613 3664
rect 2647 3656 2973 3664
rect 3267 3656 4053 3664
rect 4067 3656 4553 3664
rect 4907 3656 5193 3664
rect 6247 3656 6333 3664
rect 6347 3656 7773 3664
rect 9816 3664 9824 3676
rect 10147 3676 11273 3684
rect 11287 3676 12173 3684
rect 12187 3676 12193 3684
rect 7827 3656 9824 3664
rect 9907 3656 10093 3664
rect 10167 3656 10333 3664
rect 10847 3656 10893 3664
rect 11107 3656 11453 3664
rect 11487 3656 11653 3664
rect 11667 3656 11693 3664
rect 11707 3656 11993 3664
rect 667 3636 953 3644
rect 1947 3636 2453 3644
rect 2567 3636 3053 3644
rect 5647 3636 5673 3644
rect 7387 3636 7453 3644
rect 8207 3636 8453 3644
rect 8627 3636 9673 3644
rect 10307 3636 10473 3644
rect 10487 3636 10853 3644
rect 207 3616 333 3624
rect 667 3616 1933 3624
rect 2427 3616 2493 3624
rect 2747 3616 2873 3624
rect 2947 3616 2993 3624
rect 3907 3616 4333 3624
rect 4347 3616 4513 3624
rect 5187 3616 5313 3624
rect 5327 3616 5893 3624
rect 6747 3616 6873 3624
rect 7107 3616 7953 3624
rect 8007 3616 8233 3624
rect 8247 3616 8393 3624
rect 8407 3616 8993 3624
rect 9287 3616 9373 3624
rect 9387 3616 9653 3624
rect 10467 3616 10873 3624
rect 11687 3616 11793 3624
rect 1267 3596 1393 3604
rect 1467 3596 1613 3604
rect 2767 3596 3773 3604
rect 3787 3596 3933 3604
rect 3947 3596 4373 3604
rect 4387 3596 4413 3604
rect 6247 3596 10233 3604
rect 10547 3596 11633 3604
rect 587 3576 1073 3584
rect 1087 3576 1853 3584
rect 1867 3576 2173 3584
rect 2187 3576 2273 3584
rect 2567 3576 2733 3584
rect 2847 3576 3273 3584
rect 3567 3576 3693 3584
rect 5707 3576 5753 3584
rect 6087 3576 6133 3584
rect 7787 3576 8213 3584
rect 10947 3576 11273 3584
rect 11287 3576 11413 3584
rect 11427 3576 11733 3584
rect 767 3556 1213 3564
rect 1747 3556 1793 3564
rect 2727 3556 2953 3564
rect 2967 3556 3033 3564
rect 5267 3556 5653 3564
rect 5667 3556 5733 3564
rect 6107 3556 6513 3564
rect 6587 3556 7873 3564
rect 8107 3556 10013 3564
rect 10287 3556 10633 3564
rect 10727 3556 11013 3564
rect 11027 3556 11353 3564
rect 11827 3556 11893 3564
rect 627 3536 733 3544
rect 827 3536 1033 3544
rect 1907 3536 2113 3544
rect 2227 3536 2313 3544
rect 2367 3536 3193 3544
rect 447 3516 573 3524
rect 847 3516 913 3524
rect 956 3516 1773 3524
rect 387 3496 393 3504
rect 407 3496 473 3504
rect 956 3504 964 3516
rect 1807 3516 1924 3524
rect 1916 3507 1924 3516
rect 2187 3516 2313 3524
rect 2747 3516 2993 3524
rect 3176 3507 3184 3536
rect 3247 3536 3753 3544
rect 4587 3536 4693 3544
rect 5207 3536 5353 3544
rect 5367 3536 5593 3544
rect 5607 3536 5773 3544
rect 5787 3536 5973 3544
rect 5987 3536 6153 3544
rect 6547 3536 7673 3544
rect 7687 3536 7853 3544
rect 8287 3536 8333 3544
rect 8487 3536 9013 3544
rect 9067 3536 9173 3544
rect 9407 3536 9433 3544
rect 9927 3536 9973 3544
rect 10127 3536 10453 3544
rect 10507 3536 10833 3544
rect 11036 3536 11593 3544
rect 4107 3516 4153 3524
rect 4987 3516 5553 3524
rect 5847 3516 5933 3524
rect 6047 3516 6053 3524
rect 6067 3516 6113 3524
rect 6727 3516 7393 3524
rect 7887 3516 7893 3524
rect 7907 3516 8113 3524
rect 8127 3516 8133 3524
rect 8307 3516 8413 3524
rect 8427 3516 8504 3524
rect 607 3496 964 3504
rect 1787 3496 1873 3504
rect 2067 3496 2233 3504
rect 2247 3496 2333 3504
rect 3027 3496 3164 3504
rect 467 3476 513 3484
rect 527 3476 633 3484
rect 1167 3476 1193 3484
rect 1987 3476 2093 3484
rect 2116 3476 2693 3484
rect 2116 3467 2124 3476
rect 2707 3476 2973 3484
rect 3156 3484 3164 3496
rect 3196 3484 3204 3513
rect 3227 3496 3273 3504
rect 4187 3496 4373 3504
rect 4687 3496 5013 3504
rect 5027 3496 5053 3504
rect 5136 3496 5373 3504
rect 5136 3487 5144 3496
rect 5587 3496 5693 3504
rect 5967 3496 6073 3504
rect 6367 3496 6513 3504
rect 6556 3504 6564 3513
rect 6556 3496 6613 3504
rect 7327 3496 7833 3504
rect 8496 3504 8504 3516
rect 8527 3516 8613 3524
rect 8627 3516 8833 3524
rect 8967 3516 9113 3524
rect 9127 3516 9233 3524
rect 9467 3516 9573 3524
rect 10127 3516 10413 3524
rect 10527 3516 10673 3524
rect 10827 3516 10913 3524
rect 11036 3524 11044 3536
rect 11787 3536 12053 3544
rect 10927 3516 11044 3524
rect 11207 3516 11233 3524
rect 11387 3516 11433 3524
rect 11807 3516 11833 3524
rect 12047 3516 12073 3524
rect 8496 3496 8633 3504
rect 9007 3496 9033 3504
rect 9616 3504 9624 3513
rect 9056 3496 9624 3504
rect 3156 3476 3204 3484
rect 3547 3476 3573 3484
rect 5747 3476 6053 3484
rect 7047 3476 7073 3484
rect 7087 3476 7733 3484
rect 7927 3476 8433 3484
rect 8447 3476 8913 3484
rect 9056 3484 9064 3496
rect 9767 3496 9813 3504
rect 10007 3496 10533 3504
rect 10567 3496 10613 3504
rect 10667 3496 10793 3504
rect 11056 3504 11064 3513
rect 10887 3496 11064 3504
rect 11267 3496 11353 3504
rect 11427 3496 11513 3504
rect 11567 3496 11613 3504
rect 11847 3496 11893 3504
rect 8927 3476 9064 3484
rect 9087 3476 9824 3484
rect 1187 3456 1293 3464
rect 2307 3456 2353 3464
rect 2467 3456 3373 3464
rect 3567 3456 3593 3464
rect 6507 3456 7273 3464
rect 7287 3456 7773 3464
rect 7907 3456 9293 3464
rect 9816 3464 9824 3476
rect 9847 3476 9893 3484
rect 11216 3484 11224 3493
rect 10556 3476 11233 3484
rect 10556 3464 10564 3476
rect 11447 3476 11533 3484
rect 11647 3476 11713 3484
rect 11767 3476 11813 3484
rect 11827 3476 12013 3484
rect 9816 3456 10564 3464
rect 10627 3456 11193 3464
rect 11327 3456 11453 3464
rect 11747 3456 11853 3464
rect 907 3436 6473 3444
rect 6956 3436 8853 3444
rect 867 3416 2113 3424
rect 3427 3416 3493 3424
rect 3507 3416 4013 3424
rect 6956 3424 6964 3436
rect 9107 3436 9753 3444
rect 9847 3436 10253 3444
rect 5707 3416 6964 3424
rect 7167 3416 8053 3424
rect 8147 3416 9233 3424
rect 10047 3416 10284 3424
rect 1707 3396 6273 3404
rect 6807 3396 8973 3404
rect 9387 3396 10253 3404
rect 10276 3404 10284 3416
rect 10276 3396 10913 3404
rect 587 3376 773 3384
rect 1067 3376 2293 3384
rect 3187 3376 4713 3384
rect 8007 3376 8744 3384
rect 2547 3356 2673 3364
rect 5507 3356 5753 3364
rect 8736 3364 8744 3376
rect 8847 3376 9493 3384
rect 9587 3376 11073 3384
rect 11087 3376 11213 3384
rect 8736 3356 9113 3364
rect 9127 3356 9633 3364
rect 9647 3356 10153 3364
rect 10187 3356 10893 3364
rect 10907 3356 11033 3364
rect 1267 3336 1953 3344
rect 2507 3336 2793 3344
rect 2867 3336 5213 3344
rect 8347 3336 9393 3344
rect 10007 3336 10333 3344
rect 10347 3336 10433 3344
rect 10467 3336 11373 3344
rect 11407 3336 11753 3344
rect 6687 3316 8613 3324
rect 10167 3316 10993 3324
rect 11007 3316 11673 3324
rect 2907 3296 3033 3304
rect 3047 3296 3173 3304
rect 3787 3296 4033 3304
rect 7367 3296 7953 3304
rect 7967 3296 8513 3304
rect 8547 3296 9013 3304
rect 9187 3296 9313 3304
rect 9667 3296 9693 3304
rect 10967 3296 11253 3304
rect 11267 3296 11393 3304
rect 11827 3296 12073 3304
rect 1087 3276 1173 3284
rect 1187 3276 1993 3284
rect 3067 3276 3753 3284
rect 3767 3276 3853 3284
rect 3867 3276 4093 3284
rect 6947 3276 8153 3284
rect 8167 3276 8233 3284
rect 8707 3276 9173 3284
rect 9247 3276 9833 3284
rect 9907 3276 10213 3284
rect 10287 3276 10373 3284
rect 10787 3276 11033 3284
rect 11047 3276 11173 3284
rect 11187 3276 11473 3284
rect 11487 3276 12093 3284
rect 47 3256 513 3264
rect 1107 3256 1233 3264
rect 1547 3256 1913 3264
rect 2007 3256 2393 3264
rect 2407 3256 2813 3264
rect 2827 3256 3113 3264
rect 3147 3256 3353 3264
rect 3647 3256 3713 3264
rect 3876 3256 4233 3264
rect 3876 3247 3884 3256
rect 4567 3256 4833 3264
rect 4847 3256 5313 3264
rect 6067 3256 6313 3264
rect 7567 3256 7593 3264
rect 7647 3256 7793 3264
rect 7847 3256 8373 3264
rect 8687 3256 8713 3264
rect 8807 3256 8973 3264
rect 9187 3256 9253 3264
rect 9407 3256 10293 3264
rect 10347 3256 10513 3264
rect 10547 3256 10573 3264
rect 11287 3256 11893 3264
rect 11947 3256 12013 3264
rect 12067 3256 12264 3264
rect 407 3236 853 3244
rect 1067 3236 1213 3244
rect 1607 3236 1833 3244
rect 1127 3216 1173 3224
rect 1527 3216 1613 3224
rect 1776 3224 1784 3236
rect 1947 3236 1973 3244
rect 3027 3236 3113 3244
rect 3227 3236 3393 3244
rect 3747 3236 3773 3244
rect 3947 3236 4133 3244
rect 4227 3236 4413 3244
rect 4907 3236 5173 3244
rect 5187 3236 5653 3244
rect 5676 3236 5873 3244
rect 1776 3216 1793 3224
rect 3207 3216 3233 3224
rect 3987 3216 4013 3224
rect 4027 3216 4053 3224
rect 5676 3224 5684 3236
rect 5887 3236 6273 3244
rect 6327 3236 6593 3244
rect 6876 3244 6884 3253
rect 6647 3236 6884 3244
rect 7047 3236 7204 3244
rect 4107 3216 5684 3224
rect 6087 3216 6433 3224
rect 6847 3216 7153 3224
rect 7196 3224 7204 3236
rect 7236 3244 7244 3253
rect 7227 3236 7244 3244
rect 7267 3236 7293 3244
rect 8047 3236 8093 3244
rect 8116 3236 8173 3244
rect 7196 3216 7233 3224
rect 7387 3216 7393 3224
rect 7407 3216 7453 3224
rect 7607 3216 7673 3224
rect 7996 3224 8004 3233
rect 7687 3216 8004 3224
rect 8116 3224 8124 3236
rect 8227 3236 8393 3244
rect 8447 3236 8824 3244
rect 8816 3227 8824 3236
rect 8836 3236 8873 3244
rect 8027 3216 8124 3224
rect 8247 3216 8533 3224
rect 8667 3216 8793 3224
rect 8836 3207 8844 3236
rect 9067 3236 9224 3244
rect 9216 3227 9224 3236
rect 9567 3236 9993 3244
rect 10087 3236 10233 3244
rect 10247 3236 10573 3244
rect 11147 3236 11164 3244
rect 8987 3216 9033 3224
rect 9867 3216 9893 3224
rect 10296 3216 10873 3224
rect 687 3196 913 3204
rect 3127 3196 3533 3204
rect 3587 3196 3933 3204
rect 5487 3196 5833 3204
rect 5907 3196 6693 3204
rect 6707 3196 6813 3204
rect 6867 3196 7053 3204
rect 7447 3196 7573 3204
rect 7587 3196 8033 3204
rect 8047 3196 8193 3204
rect 8387 3196 8493 3204
rect 8887 3196 8913 3204
rect 9127 3196 9153 3204
rect 9387 3196 9413 3204
rect 9707 3196 10053 3204
rect 10296 3204 10304 3216
rect 11156 3224 11164 3236
rect 11156 3216 11333 3224
rect 11347 3216 11553 3224
rect 11567 3216 11713 3224
rect 11947 3216 12053 3224
rect 12127 3216 12264 3224
rect 10067 3196 10304 3204
rect 10347 3196 10393 3204
rect 10447 3196 10593 3204
rect 10647 3196 11124 3204
rect 567 3176 2413 3184
rect 3007 3176 3953 3184
rect 3967 3176 4393 3184
rect 5347 3176 6653 3184
rect 6827 3176 7213 3184
rect 7227 3176 7413 3184
rect 7627 3176 8413 3184
rect 9127 3176 9253 3184
rect 9287 3176 9713 3184
rect 9747 3176 9853 3184
rect 9867 3176 10473 3184
rect 10487 3176 10753 3184
rect 11116 3184 11124 3196
rect 11167 3196 11253 3204
rect 11707 3196 11753 3204
rect 11767 3196 11773 3204
rect 11887 3196 12033 3204
rect 11116 3176 11353 3184
rect 11367 3176 11393 3184
rect 11587 3176 11653 3184
rect 11727 3176 11833 3184
rect 11847 3176 11873 3184
rect 11887 3176 11893 3184
rect 147 3156 193 3164
rect 2027 3156 2133 3164
rect 3587 3156 6253 3164
rect 6507 3156 7333 3164
rect 8727 3156 9213 3164
rect 9227 3156 9553 3164
rect 9667 3156 9813 3164
rect 9847 3156 9953 3164
rect 10147 3156 10213 3164
rect 10307 3156 10393 3164
rect 10747 3156 10993 3164
rect 11307 3156 11653 3164
rect 11667 3156 11733 3164
rect 207 3136 893 3144
rect 1467 3136 1653 3144
rect 1667 3136 1793 3144
rect 1807 3136 2093 3144
rect 2107 3136 3344 3144
rect 347 3116 993 3124
rect 1007 3116 1753 3124
rect 1767 3116 1833 3124
rect 1847 3116 2313 3124
rect 2647 3116 2893 3124
rect 2987 3116 3133 3124
rect 3336 3124 3344 3136
rect 3367 3136 3993 3144
rect 4387 3136 4653 3144
rect 6287 3136 6293 3144
rect 6307 3136 7653 3144
rect 7667 3136 8933 3144
rect 9007 3136 9253 3144
rect 9307 3136 10013 3144
rect 10107 3136 10833 3144
rect 11267 3136 11513 3144
rect 11527 3136 11953 3144
rect 3336 3116 4853 3124
rect 5667 3116 5713 3124
rect 5727 3116 6713 3124
rect 6736 3116 8213 3124
rect 267 3096 493 3104
rect 1527 3096 2193 3104
rect 2207 3096 2473 3104
rect 2827 3096 3333 3104
rect 3347 3096 3893 3104
rect 4767 3096 4913 3104
rect 4927 3096 6253 3104
rect 6736 3104 6744 3116
rect 8927 3116 10733 3124
rect 10847 3116 10933 3124
rect 11107 3116 11133 3124
rect 11327 3116 11373 3124
rect 6267 3096 6744 3104
rect 7267 3096 7293 3104
rect 7887 3096 9404 3104
rect 187 3076 313 3084
rect 327 3076 1844 3084
rect 127 3056 353 3064
rect 767 3056 1193 3064
rect 1247 3056 1433 3064
rect 1447 3056 1613 3064
rect 1836 3064 1844 3076
rect 2607 3076 2653 3084
rect 2747 3076 2813 3084
rect 2987 3076 3653 3084
rect 4827 3076 5153 3084
rect 6707 3076 7033 3084
rect 7227 3076 7433 3084
rect 7447 3076 8093 3084
rect 8467 3076 8613 3084
rect 8867 3076 9333 3084
rect 9396 3084 9404 3096
rect 9427 3096 9433 3104
rect 9447 3096 11773 3104
rect 9396 3076 9553 3084
rect 9707 3076 10293 3084
rect 10567 3076 10693 3084
rect 10707 3076 10773 3084
rect 10927 3076 11073 3084
rect 11087 3076 11153 3084
rect 11167 3076 11513 3084
rect 1836 3056 3353 3064
rect 3547 3056 3853 3064
rect 3887 3056 4033 3064
rect 4187 3056 4233 3064
rect 4247 3056 4393 3064
rect 4567 3056 4633 3064
rect 4707 3056 4893 3064
rect 4907 3056 4973 3064
rect 5827 3056 5933 3064
rect 6147 3056 6473 3064
rect 6667 3056 6713 3064
rect 7087 3056 7273 3064
rect 7427 3056 7893 3064
rect 8267 3056 8353 3064
rect 8367 3056 8473 3064
rect 8487 3056 8653 3064
rect 9007 3056 9073 3064
rect 9087 3056 9173 3064
rect 9187 3056 9373 3064
rect 9467 3056 9733 3064
rect 9756 3056 10253 3064
rect 387 3036 433 3044
rect 467 3036 513 3044
rect 907 3036 1184 3044
rect 127 3016 153 3024
rect 336 3024 344 3033
rect 207 3016 344 3024
rect 507 3016 633 3024
rect 947 3016 973 3024
rect 1027 3016 1153 3024
rect 1176 3024 1184 3036
rect 1347 3036 1753 3044
rect 1776 3027 1784 3053
rect 2847 3036 3693 3044
rect 3847 3036 4093 3044
rect 4447 3036 4493 3044
rect 4667 3036 4713 3044
rect 4727 3036 4804 3044
rect 4796 3027 4804 3036
rect 6307 3036 6333 3044
rect 6467 3036 6473 3044
rect 6487 3036 6633 3044
rect 7127 3036 7233 3044
rect 7287 3036 7393 3044
rect 7667 3036 7733 3044
rect 8087 3036 8413 3044
rect 8707 3036 8793 3044
rect 8807 3036 8813 3044
rect 9147 3036 9173 3044
rect 9307 3036 9593 3044
rect 9756 3044 9764 3056
rect 10267 3056 10333 3064
rect 10347 3056 10353 3064
rect 10416 3056 11093 3064
rect 9607 3036 9764 3044
rect 9776 3036 9993 3044
rect 1176 3016 1213 3024
rect 1387 3016 1404 3024
rect -24 2996 453 3004
rect 1247 2996 1353 3004
rect 1396 3004 1404 3016
rect 1427 3016 1453 3024
rect 1476 3016 1573 3024
rect 1476 3004 1484 3016
rect 2247 3016 2273 3024
rect 2327 3016 2653 3024
rect 3007 3016 3073 3024
rect 3307 3016 3333 3024
rect 3527 3016 3653 3024
rect 3667 3016 4073 3024
rect 6687 3016 6793 3024
rect 6856 3024 6864 3033
rect 6856 3016 7053 3024
rect 7636 3024 7644 3033
rect 7636 3016 7813 3024
rect 8027 3016 8333 3024
rect 8436 3024 8444 3033
rect 8436 3016 8633 3024
rect 8687 3016 8913 3024
rect 8987 3016 9033 3024
rect 9347 3016 9693 3024
rect 9776 3024 9784 3036
rect 10416 3044 10424 3056
rect 11187 3056 11333 3064
rect 11787 3056 11913 3064
rect 11947 3056 12073 3064
rect 10116 3036 10424 3044
rect 9767 3016 9784 3024
rect 9907 3016 9953 3024
rect 10116 3024 10124 3036
rect 10447 3036 10493 3044
rect 10587 3036 10593 3044
rect 10607 3036 10793 3044
rect 10947 3036 10973 3044
rect 11027 3036 11293 3044
rect 11367 3036 11413 3044
rect 11467 3036 11493 3044
rect 11687 3036 11713 3044
rect 11876 3036 11913 3044
rect 9987 3016 10124 3024
rect 10487 3016 10513 3024
rect 10987 3016 11053 3024
rect 11387 3016 11493 3024
rect 11516 3016 11533 3024
rect 1396 2996 1484 3004
rect 1867 2996 1993 3004
rect 2187 2996 3053 3004
rect 3067 2996 3113 3004
rect 3327 2996 3473 3004
rect 3527 2996 3673 3004
rect 3987 2996 4093 3004
rect 4836 3004 4844 3013
rect 4507 2996 4844 3004
rect 5267 2996 5373 3004
rect 7107 2996 7193 3004
rect 7287 2996 7413 3004
rect 7467 2996 7513 3004
rect 7627 2996 7753 3004
rect 8587 2996 8773 3004
rect 8807 2996 9013 3004
rect 9107 2996 9133 3004
rect 9527 2996 10053 3004
rect 10136 3004 10144 3013
rect 10067 2996 10144 3004
rect 10327 2996 10513 3004
rect 10527 2996 10593 3004
rect 10767 2996 10913 3004
rect 10967 2996 11293 3004
rect 11516 3004 11524 3016
rect 11876 3024 11884 3036
rect 11547 3016 11884 3024
rect 11327 2996 11524 3004
rect 11747 2996 11833 3004
rect 12147 2996 12264 3004
rect 27 2976 3293 2984
rect 3307 2976 3573 2984
rect 3727 2976 4413 2984
rect 4767 2976 5953 2984
rect 6847 2976 6913 2984
rect 8467 2976 8853 2984
rect 8867 2976 8873 2984
rect 8947 2976 9793 2984
rect 9947 2976 10033 2984
rect 10767 2976 11193 2984
rect 11447 2976 11493 2984
rect 11707 2976 11753 2984
rect 11767 2976 11853 2984
rect 2347 2956 2613 2964
rect 3507 2956 4013 2964
rect 4307 2956 4473 2964
rect 4487 2956 4893 2964
rect 7127 2956 10173 2964
rect 11087 2956 11153 2964
rect 2247 2936 3453 2944
rect 5707 2936 7553 2944
rect 8107 2936 11073 2944
rect 87 2916 273 2924
rect 2967 2916 3173 2924
rect 5147 2916 5913 2924
rect 6667 2916 8013 2924
rect 8407 2916 9133 2924
rect 9147 2916 9653 2924
rect 9727 2916 10433 2924
rect 11527 2916 11593 2924
rect 1987 2896 2853 2904
rect 3887 2896 4253 2904
rect 7447 2896 7653 2904
rect 7667 2896 7913 2904
rect 9027 2896 9193 2904
rect 9247 2896 9313 2904
rect 10147 2896 10273 2904
rect 10336 2896 10633 2904
rect 407 2876 2253 2884
rect 2267 2876 3393 2884
rect 5887 2876 7173 2884
rect 7347 2876 8413 2884
rect 9047 2876 9293 2884
rect 10336 2884 10344 2896
rect 10887 2896 11373 2904
rect 9327 2876 10344 2884
rect 11427 2876 11913 2884
rect 1527 2856 1553 2864
rect 5447 2856 6113 2864
rect 7427 2856 8013 2864
rect 8107 2856 8973 2864
rect 8987 2856 9293 2864
rect 9407 2856 10093 2864
rect 10347 2856 11013 2864
rect 11087 2856 11273 2864
rect 11707 2856 11813 2864
rect 47 2836 93 2844
rect 107 2836 2993 2844
rect 5287 2836 5353 2844
rect 5407 2836 6193 2844
rect 6887 2836 7113 2844
rect 7127 2836 7733 2844
rect 7747 2836 8093 2844
rect 8687 2836 9353 2844
rect 10367 2836 11553 2844
rect 11716 2836 11893 2844
rect 6047 2816 7513 2824
rect 7807 2816 8453 2824
rect 8867 2816 9113 2824
rect 9187 2816 10593 2824
rect 10667 2816 10873 2824
rect 11107 2816 11413 2824
rect 11716 2824 11724 2836
rect 11427 2816 11724 2824
rect 11747 2816 11773 2824
rect 2687 2796 2773 2804
rect 3167 2796 3233 2804
rect 3487 2796 3513 2804
rect 4187 2796 5153 2804
rect 5987 2796 6713 2804
rect 6887 2796 7133 2804
rect 7787 2796 7893 2804
rect 7947 2796 7993 2804
rect 8247 2796 9393 2804
rect 9587 2796 9833 2804
rect 9907 2796 9973 2804
rect 10807 2796 11633 2804
rect 11647 2796 11773 2804
rect 11787 2796 12053 2804
rect 12067 2796 12073 2804
rect 607 2776 613 2784
rect 627 2776 1073 2784
rect 2707 2776 2873 2784
rect 3147 2776 3313 2784
rect 3567 2776 3593 2784
rect 3807 2776 3873 2784
rect 3896 2776 4253 2784
rect -24 2744 -16 2764
rect 567 2756 753 2764
rect 1687 2756 1873 2764
rect 1927 2756 2093 2764
rect 2127 2756 2273 2764
rect 2327 2756 2373 2764
rect 2727 2756 2793 2764
rect 3027 2756 3773 2764
rect 3896 2764 3904 2776
rect 4267 2776 4293 2784
rect 4416 2776 4593 2784
rect 3827 2756 3904 2764
rect 4047 2756 4233 2764
rect 4416 2764 4424 2776
rect 4607 2776 4753 2784
rect 4767 2776 4933 2784
rect 5387 2776 6333 2784
rect 6347 2776 6553 2784
rect 6567 2776 6813 2784
rect 7647 2776 7913 2784
rect 8027 2776 8993 2784
rect 9087 2776 9153 2784
rect 9787 2776 9913 2784
rect 10307 2776 10613 2784
rect 10627 2776 10733 2784
rect 11227 2776 11273 2784
rect 11407 2776 11533 2784
rect 11567 2776 11813 2784
rect 11827 2776 11873 2784
rect 4287 2756 4424 2764
rect 4447 2756 4513 2764
rect 4647 2756 4733 2764
rect 4827 2756 4973 2764
rect 5027 2756 5513 2764
rect 5607 2756 5913 2764
rect 5956 2756 6133 2764
rect 5956 2747 5964 2756
rect 6187 2756 6384 2764
rect 6376 2747 6384 2756
rect 6407 2756 6453 2764
rect 6727 2756 6753 2764
rect 6807 2756 6944 2764
rect -24 2736 133 2744
rect 527 2736 653 2744
rect 1407 2736 1893 2744
rect 1907 2736 1973 2744
rect 2227 2736 2293 2744
rect 2496 2736 2673 2744
rect 2496 2727 2504 2736
rect 2967 2736 3213 2744
rect 4007 2736 4173 2744
rect 4207 2736 4413 2744
rect 4507 2736 4553 2744
rect 5187 2736 5353 2744
rect 5547 2736 5573 2744
rect 6007 2736 6033 2744
rect 6127 2736 6333 2744
rect 6447 2736 6613 2744
rect 6627 2736 6913 2744
rect 6936 2744 6944 2756
rect 6987 2756 7113 2764
rect 7136 2756 7353 2764
rect 6936 2736 6993 2744
rect 7136 2744 7144 2756
rect 7367 2756 7393 2764
rect 7607 2756 7693 2764
rect 7747 2756 7773 2764
rect 7787 2756 8033 2764
rect 8267 2756 8293 2764
rect 8316 2756 8493 2764
rect 8316 2747 8324 2756
rect 8547 2756 8653 2764
rect 8767 2756 8793 2764
rect 9367 2756 9393 2764
rect 9467 2756 9493 2764
rect 9547 2756 9593 2764
rect 9727 2756 9753 2764
rect 9916 2756 9973 2764
rect 9916 2747 9924 2756
rect 10267 2756 10313 2764
rect 10847 2756 10893 2764
rect 11067 2756 11113 2764
rect 11807 2756 11833 2764
rect 7007 2736 7144 2744
rect 7187 2736 7213 2744
rect 7327 2736 7573 2744
rect 7767 2736 7793 2744
rect 7827 2736 7993 2744
rect 8007 2736 8153 2744
rect 8527 2736 8593 2744
rect 8787 2736 8893 2744
rect 9627 2736 9733 2744
rect 9967 2736 9993 2744
rect 10007 2736 10153 2744
rect 10167 2736 10453 2744
rect 10607 2736 11204 2744
rect 11196 2727 11204 2736
rect 11227 2736 11393 2744
rect 11447 2736 11853 2744
rect 11867 2736 11933 2744
rect 12256 2744 12264 2764
rect 12167 2736 12264 2744
rect 1707 2716 1933 2724
rect 2067 2716 2173 2724
rect 2647 2716 2853 2724
rect 2867 2716 3053 2724
rect 4147 2716 4453 2724
rect 4727 2716 4773 2724
rect 5427 2716 5733 2724
rect 5747 2716 6533 2724
rect 6587 2716 6853 2724
rect 6887 2716 6953 2724
rect 7267 2716 7333 2724
rect 7547 2716 7593 2724
rect 8147 2716 8273 2724
rect 8747 2716 8853 2724
rect 8967 2716 9033 2724
rect 9167 2716 9333 2724
rect 9647 2716 9693 2724
rect 9707 2716 9933 2724
rect 9947 2716 10113 2724
rect 11047 2716 11073 2724
rect 11567 2716 11593 2724
rect 11647 2716 11753 2724
rect 11887 2716 11953 2724
rect 587 2696 1393 2704
rect 1747 2696 2053 2704
rect 2467 2696 2493 2704
rect 3527 2696 3593 2704
rect 3607 2696 4313 2704
rect 4427 2696 4813 2704
rect 5527 2696 5933 2704
rect 6587 2696 7013 2704
rect 7247 2696 7773 2704
rect 7967 2696 8053 2704
rect 8087 2696 8453 2704
rect 8807 2696 9613 2704
rect 9727 2696 9753 2704
rect 9807 2696 9893 2704
rect 9927 2696 9953 2704
rect 10847 2696 11373 2704
rect 11547 2696 11793 2704
rect 1067 2676 1713 2684
rect 1947 2676 2333 2684
rect 2887 2676 3933 2684
rect 4747 2676 4953 2684
rect 5927 2676 6153 2684
rect 6467 2676 6733 2684
rect 8907 2676 9513 2684
rect 9927 2676 10573 2684
rect 10587 2676 10633 2684
rect 11007 2676 11033 2684
rect 11507 2676 11593 2684
rect 967 2656 1433 2664
rect 1447 2656 1553 2664
rect 1667 2656 2073 2664
rect 3947 2656 4113 2664
rect 5947 2656 6233 2664
rect 6927 2656 8833 2664
rect 8847 2656 9144 2664
rect 647 2636 2533 2644
rect 2547 2636 2633 2644
rect 6047 2636 6953 2644
rect 7387 2636 7673 2644
rect 8667 2636 9113 2644
rect 9136 2644 9144 2656
rect 9167 2656 9673 2664
rect 9687 2656 10453 2664
rect 10467 2656 10753 2664
rect 11527 2656 11573 2664
rect 11687 2656 11813 2664
rect 9136 2636 9333 2644
rect 9367 2636 10013 2644
rect 10407 2636 10613 2644
rect 10747 2636 10993 2644
rect 11007 2636 11073 2644
rect 11627 2636 11713 2644
rect 11867 2636 11893 2644
rect 947 2616 2473 2624
rect 2487 2616 3533 2624
rect 5607 2616 5613 2624
rect 5627 2616 5953 2624
rect 5967 2616 6173 2624
rect 6187 2616 6413 2624
rect 6787 2616 7433 2624
rect 8207 2616 8973 2624
rect 8987 2616 9513 2624
rect 9527 2616 9733 2624
rect 9747 2616 10193 2624
rect 11167 2616 11213 2624
rect 1187 2596 2213 2604
rect 3047 2596 3093 2604
rect 3107 2596 3353 2604
rect 3927 2596 3953 2604
rect 5187 2596 5213 2604
rect 5747 2596 5773 2604
rect 6207 2596 8253 2604
rect 8427 2596 9473 2604
rect 9687 2596 10273 2604
rect 10427 2596 10773 2604
rect 11147 2596 11173 2604
rect 11327 2596 11433 2604
rect 307 2576 433 2584
rect 447 2576 673 2584
rect 687 2576 893 2584
rect 907 2576 953 2584
rect 1147 2576 1373 2584
rect 2147 2576 2253 2584
rect 2267 2576 2713 2584
rect 3007 2576 3193 2584
rect 3527 2576 3553 2584
rect 3867 2576 3893 2584
rect 3907 2576 4373 2584
rect 4647 2576 4873 2584
rect 5287 2576 6353 2584
rect 6627 2576 6813 2584
rect 6947 2576 6993 2584
rect 7567 2576 7633 2584
rect 7647 2576 7713 2584
rect 7807 2576 8073 2584
rect 8247 2576 8433 2584
rect 8687 2576 8813 2584
rect 8976 2576 9233 2584
rect 187 2556 393 2564
rect 427 2556 633 2564
rect 2307 2556 2433 2564
rect 2587 2556 2833 2564
rect 3227 2556 3493 2564
rect 3536 2556 3693 2564
rect 3536 2547 3544 2556
rect 3767 2556 3924 2564
rect 3916 2547 3924 2556
rect 4327 2556 4693 2564
rect 5067 2556 5193 2564
rect 5247 2556 5273 2564
rect 5307 2556 5373 2564
rect 5387 2556 5584 2564
rect 5576 2547 5584 2556
rect 5687 2556 5773 2564
rect 6427 2556 6473 2564
rect 7107 2556 7133 2564
rect 7307 2556 7833 2564
rect 8567 2556 8633 2564
rect 147 2536 293 2544
rect 1207 2536 1253 2544
rect 1847 2536 2453 2544
rect 2667 2536 2793 2544
rect 3387 2536 3473 2544
rect 3747 2536 3773 2544
rect 4407 2536 4513 2544
rect 4627 2536 4653 2544
rect 5767 2536 5784 2544
rect 1087 2516 1213 2524
rect 2707 2516 2813 2524
rect 3347 2516 3713 2524
rect 4507 2516 4553 2524
rect 5776 2524 5784 2536
rect 5996 2544 6004 2553
rect 5807 2536 6004 2544
rect 6196 2544 6204 2553
rect 6027 2536 6204 2544
rect 6396 2544 6404 2553
rect 6396 2536 6593 2544
rect 6787 2536 6913 2544
rect 6987 2536 7253 2544
rect 7287 2536 7353 2544
rect 7467 2536 7533 2544
rect 7747 2536 7873 2544
rect 7907 2536 7933 2544
rect 7967 2536 8253 2544
rect 8267 2536 8713 2544
rect 8976 2544 8984 2576
rect 9247 2576 9373 2584
rect 9507 2576 9553 2584
rect 9607 2576 9713 2584
rect 10127 2576 10213 2584
rect 10287 2576 10373 2584
rect 10507 2576 10553 2584
rect 10787 2576 10953 2584
rect 10967 2576 11093 2584
rect 11127 2576 11213 2584
rect 11307 2576 11413 2584
rect 11496 2576 11513 2584
rect 11527 2576 11533 2584
rect 11687 2576 11893 2584
rect 8787 2536 8984 2544
rect 8996 2556 9033 2564
rect 5776 2516 5893 2524
rect 6776 2524 6784 2533
rect 6227 2516 6784 2524
rect 7187 2516 7373 2524
rect 7447 2516 7513 2524
rect 7567 2516 7813 2524
rect 7927 2516 7993 2524
rect 8007 2516 8373 2524
rect 8996 2524 9004 2556
rect 9327 2556 9373 2564
rect 9607 2556 9633 2564
rect 10147 2556 10253 2564
rect 10307 2556 10533 2564
rect 10647 2556 10733 2564
rect 11127 2556 11273 2564
rect 11307 2556 11713 2564
rect 11727 2556 11733 2564
rect 11867 2556 12093 2564
rect 9027 2536 9053 2544
rect 9147 2536 9213 2544
rect 9347 2536 9493 2544
rect 9547 2536 9833 2544
rect 9847 2536 9873 2544
rect 9947 2536 9973 2544
rect 10207 2536 10333 2544
rect 10567 2536 10693 2544
rect 10867 2536 10913 2544
rect 11407 2536 11413 2544
rect 11427 2536 11513 2544
rect 11827 2536 11873 2544
rect 8996 2516 9033 2524
rect 9587 2516 9693 2524
rect 9716 2516 9753 2524
rect 1567 2496 2733 2504
rect 2816 2504 2824 2513
rect 2807 2496 2824 2504
rect 3147 2496 3973 2504
rect 3987 2496 4033 2504
rect 4047 2496 5033 2504
rect 5047 2496 5253 2504
rect 5587 2496 6373 2504
rect 6387 2496 6433 2504
rect 6447 2496 6753 2504
rect 6827 2496 7173 2504
rect 7307 2496 7973 2504
rect 8327 2496 9133 2504
rect 9716 2504 9724 2516
rect 10607 2516 10713 2524
rect 10767 2516 10833 2524
rect 11107 2516 11233 2524
rect 11356 2524 11364 2533
rect 11356 2516 11433 2524
rect 9147 2496 9724 2504
rect 10267 2496 10393 2504
rect 10407 2496 10473 2504
rect 10787 2496 11253 2504
rect 11327 2496 11653 2504
rect 11667 2496 11933 2504
rect 11947 2496 11973 2504
rect 4707 2476 4733 2484
rect 5687 2476 5773 2484
rect 6647 2476 6673 2484
rect 6707 2476 6773 2484
rect 7547 2476 7573 2484
rect 7707 2476 8213 2484
rect 9027 2476 9273 2484
rect 9447 2476 9804 2484
rect 2367 2456 2513 2464
rect 2527 2456 2913 2464
rect 5747 2456 7233 2464
rect 7527 2456 8193 2464
rect 8356 2456 8773 2464
rect 7027 2436 7393 2444
rect 8356 2444 8364 2456
rect 9347 2456 9453 2464
rect 9796 2464 9804 2476
rect 9827 2476 10853 2484
rect 10927 2476 11473 2484
rect 9796 2456 10293 2464
rect 10327 2456 11353 2464
rect 7447 2436 8364 2444
rect 8667 2436 9433 2444
rect 9467 2436 9913 2444
rect 10467 2436 11133 2444
rect 11227 2436 11413 2444
rect 6747 2416 7573 2424
rect 7587 2416 9053 2424
rect 9387 2416 9653 2424
rect 9667 2416 10373 2424
rect 11227 2416 11433 2424
rect 6527 2396 7713 2404
rect 7867 2396 8593 2404
rect 8607 2396 8613 2404
rect 9407 2396 9673 2404
rect 9687 2396 9733 2404
rect 10087 2396 10333 2404
rect 10567 2396 12053 2404
rect 3207 2376 3233 2384
rect 6587 2376 7093 2384
rect 7227 2376 7333 2384
rect 7347 2376 8233 2384
rect 8367 2376 8533 2384
rect 8587 2376 10273 2384
rect 6867 2356 7624 2364
rect -24 2336 33 2344
rect 287 2336 1433 2344
rect 1447 2336 3813 2344
rect 3827 2336 4673 2344
rect 7027 2336 7153 2344
rect 7287 2336 7593 2344
rect 7616 2344 7624 2356
rect 7987 2356 8553 2364
rect 8567 2356 8673 2364
rect 9187 2356 10053 2364
rect 10147 2356 10744 2364
rect 7616 2336 8273 2344
rect 8607 2336 8733 2344
rect 8767 2336 9413 2344
rect 9447 2336 9473 2344
rect 9727 2336 9773 2344
rect 9987 2336 10653 2344
rect 10736 2344 10744 2356
rect 10767 2356 11093 2364
rect 10736 2336 11813 2344
rect 147 2316 193 2324
rect 207 2316 413 2324
rect 1887 2316 2353 2324
rect 2927 2316 2953 2324
rect 2967 2316 3433 2324
rect 3447 2316 3733 2324
rect 3747 2316 3773 2324
rect 5187 2316 5233 2324
rect 5747 2316 5813 2324
rect 5987 2316 6053 2324
rect 6767 2316 6813 2324
rect 7047 2316 7133 2324
rect 7387 2316 7933 2324
rect 8187 2316 8253 2324
rect 8387 2316 8573 2324
rect 8647 2316 8913 2324
rect 9087 2316 9813 2324
rect 10067 2316 10213 2324
rect 10307 2316 10433 2324
rect 10547 2316 10673 2324
rect 10867 2316 11253 2324
rect 11507 2316 11553 2324
rect 11707 2316 11753 2324
rect 187 2296 393 2304
rect 407 2296 513 2304
rect 687 2296 1073 2304
rect 1087 2296 1313 2304
rect 1587 2296 1993 2304
rect 2007 2296 2013 2304
rect 3027 2296 3053 2304
rect 3567 2296 3913 2304
rect 3927 2296 4093 2304
rect 5227 2296 5833 2304
rect 6367 2296 6513 2304
rect 6547 2296 6633 2304
rect 7007 2296 7093 2304
rect 7136 2296 7293 2304
rect -24 2276 1064 2284
rect 527 2256 633 2264
rect 707 2256 813 2264
rect 827 2256 853 2264
rect 907 2256 1033 2264
rect 1056 2264 1064 2276
rect 1827 2276 1933 2284
rect 2167 2276 2293 2284
rect 3047 2276 3173 2284
rect 3487 2276 3593 2284
rect 3907 2276 3953 2284
rect 4076 2276 4253 2284
rect 1056 2256 1253 2264
rect 1736 2264 1744 2273
rect 1736 2256 1893 2264
rect 2116 2264 2124 2273
rect 1967 2256 2124 2264
rect 2347 2256 2413 2264
rect 2676 2264 2684 2273
rect 4076 2267 4084 2276
rect 4267 2276 4453 2284
rect 4547 2276 5173 2284
rect 5187 2276 5293 2284
rect 5707 2276 5733 2284
rect 6116 2284 6124 2293
rect 5987 2276 6124 2284
rect 6316 2284 6324 2293
rect 6147 2276 6324 2284
rect 6347 2276 6724 2284
rect 6716 2267 6724 2276
rect 6747 2276 6853 2284
rect 7136 2284 7144 2296
rect 7327 2296 7373 2304
rect 7887 2296 8733 2304
rect 8767 2296 8953 2304
rect 8987 2296 9153 2304
rect 9267 2296 9513 2304
rect 9907 2296 10053 2304
rect 10207 2296 10813 2304
rect 10907 2296 11113 2304
rect 11467 2296 11533 2304
rect 11967 2296 12033 2304
rect 12087 2296 12104 2304
rect 12096 2287 12104 2296
rect 7096 2276 7144 2284
rect 7156 2276 7273 2284
rect 2676 2256 2833 2264
rect 2907 2256 2973 2264
rect 3047 2256 3113 2264
rect 3767 2256 3853 2264
rect 4127 2256 4233 2264
rect 4247 2256 4613 2264
rect 4647 2256 4673 2264
rect 4907 2256 5133 2264
rect 5147 2256 5153 2264
rect 5267 2256 5273 2264
rect 5287 2256 5373 2264
rect 5607 2256 5733 2264
rect 5747 2256 5853 2264
rect 5927 2256 6173 2264
rect 6187 2256 6533 2264
rect 6827 2256 6893 2264
rect 6907 2256 6993 2264
rect 7096 2264 7104 2276
rect 7087 2256 7104 2264
rect 7156 2264 7164 2276
rect 7296 2276 7493 2284
rect 7127 2256 7164 2264
rect 7296 2264 7304 2276
rect 8167 2276 8313 2284
rect 8447 2276 8713 2284
rect 8727 2276 8764 2284
rect 7267 2256 7304 2264
rect 7527 2256 7753 2264
rect 7807 2256 7913 2264
rect 8156 2264 8164 2273
rect 8127 2256 8164 2264
rect 8187 2256 8193 2264
rect 8207 2256 8293 2264
rect 8387 2256 8513 2264
rect 8687 2256 8733 2264
rect 8756 2264 8764 2276
rect 8907 2276 8933 2284
rect 8947 2276 9104 2284
rect 8756 2256 8993 2264
rect 9007 2256 9073 2264
rect 9096 2264 9104 2276
rect 9127 2276 9153 2284
rect 9287 2276 9553 2284
rect 9567 2276 9613 2284
rect 9727 2276 9853 2284
rect 9947 2276 10084 2284
rect 10076 2267 10084 2276
rect 10127 2276 10153 2284
rect 10296 2276 10353 2284
rect 9096 2256 9253 2264
rect 9467 2256 9573 2264
rect 9607 2256 9653 2264
rect 9827 2256 9873 2264
rect 27 2236 193 2244
rect 207 2236 293 2244
rect 727 2236 753 2244
rect 767 2236 833 2244
rect 847 2236 1193 2244
rect 1307 2236 1713 2244
rect 1727 2236 2233 2244
rect 2527 2236 2573 2244
rect 3027 2236 3073 2244
rect 3527 2236 3553 2244
rect 3887 2236 3913 2244
rect 4307 2236 4473 2244
rect 4867 2236 5053 2244
rect 5187 2236 5753 2244
rect 6167 2236 6373 2244
rect 6687 2236 6733 2244
rect 6927 2236 7033 2244
rect 7207 2236 7293 2244
rect 7307 2236 7473 2244
rect 7907 2236 7933 2244
rect 8147 2236 8193 2244
rect 9147 2236 9173 2244
rect 9427 2236 9973 2244
rect 10096 2244 10104 2273
rect 10296 2267 10304 2276
rect 10367 2276 10493 2284
rect 10727 2276 10833 2284
rect 10887 2276 10933 2284
rect 11087 2276 11313 2284
rect 11467 2276 11633 2284
rect 11647 2276 11653 2284
rect 11676 2276 11853 2284
rect 10227 2256 10253 2264
rect 10516 2247 10524 2273
rect 11676 2267 11684 2276
rect 11907 2276 12084 2284
rect 12076 2267 12084 2276
rect 10667 2256 10693 2264
rect 10747 2256 10853 2264
rect 11027 2256 11053 2264
rect 11307 2256 11433 2264
rect 11487 2256 11653 2264
rect 11727 2256 11793 2264
rect 11827 2256 11873 2264
rect 10007 2236 10104 2244
rect 10227 2236 10313 2244
rect 11287 2236 11313 2244
rect 11347 2236 11513 2244
rect 11607 2236 11913 2244
rect 2507 2216 2533 2224
rect 2547 2216 2933 2224
rect 2947 2216 3153 2224
rect 3647 2216 3793 2224
rect 4287 2216 4353 2224
rect 5847 2216 6153 2224
rect 6307 2216 7873 2224
rect 7967 2216 8353 2224
rect 8487 2216 8593 2224
rect 8607 2216 9973 2224
rect 9987 2216 10113 2224
rect 10127 2216 10253 2224
rect 10907 2216 11153 2224
rect 11367 2216 11453 2224
rect 11467 2216 11513 2224
rect 11547 2216 12033 2224
rect 3107 2196 3633 2204
rect 3967 2196 4653 2204
rect 5847 2196 7453 2204
rect 7467 2196 8093 2204
rect 8307 2196 8333 2204
rect 8567 2196 8913 2204
rect 8927 2196 11013 2204
rect 11107 2196 11353 2204
rect 11487 2196 11553 2204
rect 11647 2196 11753 2204
rect 2567 2176 3053 2184
rect 3067 2176 3873 2184
rect 6707 2176 6864 2184
rect 2887 2156 3053 2164
rect 6247 2156 6273 2164
rect 6527 2156 6753 2164
rect 6856 2164 6864 2176
rect 6887 2176 6933 2184
rect 8047 2176 8753 2184
rect 8767 2176 9993 2184
rect 10007 2176 10673 2184
rect 10847 2176 11793 2184
rect 6856 2156 7333 2164
rect 7387 2156 7513 2164
rect 7707 2156 8473 2164
rect 9007 2156 9353 2164
rect 9707 2156 9793 2164
rect 9927 2156 10033 2164
rect 10247 2156 10653 2164
rect 10667 2156 11093 2164
rect 11407 2156 11433 2164
rect 11567 2156 11753 2164
rect 4527 2136 4833 2144
rect 6707 2136 6953 2144
rect 7167 2136 7333 2144
rect 7347 2136 7493 2144
rect 8027 2136 8233 2144
rect 8247 2136 8293 2144
rect 8427 2136 9273 2144
rect 9427 2136 10273 2144
rect 10447 2136 10493 2144
rect 10967 2136 11933 2144
rect 1527 2116 2553 2124
rect 3887 2116 4533 2124
rect 5007 2116 5953 2124
rect 6567 2116 6713 2124
rect 6767 2116 6993 2124
rect 7007 2116 7033 2124
rect 7667 2116 7713 2124
rect 7787 2116 7873 2124
rect 8087 2116 8153 2124
rect 8187 2116 8253 2124
rect 8287 2116 8733 2124
rect 8887 2116 8973 2124
rect 8987 2116 9133 2124
rect 9307 2116 9353 2124
rect 9507 2116 9613 2124
rect 9627 2116 9693 2124
rect 9887 2116 9933 2124
rect 10227 2116 10913 2124
rect 10947 2116 11173 2124
rect 11407 2116 11573 2124
rect 11907 2116 12013 2124
rect 407 2096 593 2104
rect 707 2096 1013 2104
rect 1027 2096 1133 2104
rect 1187 2096 1233 2104
rect 1267 2096 2413 2104
rect 3647 2096 3833 2104
rect 4407 2096 4953 2104
rect 4967 2096 5213 2104
rect 5487 2096 5673 2104
rect 5967 2096 6073 2104
rect 6127 2096 6253 2104
rect 6267 2096 6313 2104
rect 6327 2096 6393 2104
rect 6407 2096 6513 2104
rect 6607 2096 6673 2104
rect 6847 2096 6953 2104
rect 6967 2096 7233 2104
rect 7487 2096 7613 2104
rect 7627 2096 7853 2104
rect 7867 2096 8093 2104
rect 8147 2096 8273 2104
rect 8407 2096 8544 2104
rect 587 2076 853 2084
rect 867 2076 1153 2084
rect 1207 2076 1473 2084
rect 2367 2076 2393 2084
rect 2607 2076 2793 2084
rect 3427 2076 3593 2084
rect 3607 2076 3833 2084
rect 4487 2076 4493 2084
rect 4507 2076 4613 2084
rect 5687 2076 5833 2084
rect 6287 2076 6433 2084
rect 6447 2076 6473 2084
rect 6527 2076 6553 2084
rect 6667 2076 6913 2084
rect 7067 2076 7133 2084
rect 7247 2076 7413 2084
rect 7667 2076 7833 2084
rect 7927 2076 8024 2084
rect 127 2056 273 2064
rect 487 2056 813 2064
rect 1367 2056 1813 2064
rect 2007 2056 2033 2064
rect 2127 2056 2473 2064
rect 2767 2056 2873 2064
rect 2887 2056 3233 2064
rect 3307 2056 3453 2064
rect 3827 2056 4093 2064
rect 4247 2056 4293 2064
rect 4396 2064 4404 2073
rect 4307 2056 4404 2064
rect 5467 2056 5653 2064
rect 5667 2056 5933 2064
rect 6067 2056 6264 2064
rect 6256 2047 6264 2056
rect 6507 2056 6593 2064
rect 6847 2056 7213 2064
rect 7456 2064 7464 2073
rect 7456 2056 7633 2064
rect 7807 2056 7853 2064
rect 7907 2056 7973 2064
rect 8016 2064 8024 2076
rect 8047 2076 8213 2084
rect 8247 2076 8513 2084
rect 8536 2084 8544 2096
rect 8567 2096 8693 2104
rect 8927 2096 9093 2104
rect 9227 2096 9313 2104
rect 10627 2096 10693 2104
rect 10827 2096 10893 2104
rect 10916 2096 10973 2104
rect 8536 2076 8653 2084
rect 8887 2076 8933 2084
rect 9107 2076 9173 2084
rect 9467 2076 9533 2084
rect 9647 2076 9773 2084
rect 9807 2076 9824 2084
rect 8016 2056 8413 2064
rect 8507 2056 8553 2064
rect 8647 2056 8673 2064
rect 8687 2056 8813 2064
rect 9127 2056 9153 2064
rect 9307 2056 9413 2064
rect 9527 2056 9573 2064
rect 9687 2056 9793 2064
rect 9816 2064 9824 2076
rect 9927 2076 9953 2084
rect 10327 2076 10464 2084
rect 10456 2067 10464 2076
rect 10487 2076 10533 2084
rect 10916 2084 10924 2096
rect 11007 2096 11093 2104
rect 11507 2096 11533 2104
rect 11547 2096 11593 2104
rect 11887 2096 11953 2104
rect 11987 2096 12013 2104
rect 10816 2076 10924 2084
rect 10816 2067 10824 2076
rect 11207 2076 11293 2084
rect 11927 2076 11993 2084
rect 9816 2056 9893 2064
rect 9916 2056 9973 2064
rect 427 2036 633 2044
rect 847 2036 993 2044
rect 1247 2036 1373 2044
rect 2367 2036 3753 2044
rect 4067 2036 4873 2044
rect 5547 2036 5893 2044
rect 5927 2036 6093 2044
rect 6276 2036 6293 2044
rect 1147 2016 1393 2024
rect 1407 2016 1413 2024
rect 2707 2016 3313 2024
rect 3327 2016 3433 2024
rect 6276 2024 6284 2036
rect 6456 2044 6464 2053
rect 6456 2036 6473 2044
rect 6787 2036 6853 2044
rect 6927 2036 7073 2044
rect 7087 2036 7173 2044
rect 7187 2036 7233 2044
rect 7456 2036 7553 2044
rect 5707 2016 6284 2024
rect 6807 2016 6833 2024
rect 7087 2016 7133 2024
rect 7456 2024 7464 2036
rect 7587 2036 7613 2044
rect 7747 2036 8133 2044
rect 8187 2036 8253 2044
rect 8507 2036 8993 2044
rect 9347 2036 9433 2044
rect 9487 2036 9833 2044
rect 9916 2044 9924 2056
rect 10567 2056 10633 2064
rect 10847 2056 10953 2064
rect 9907 2036 9924 2044
rect 9947 2036 10193 2044
rect 10207 2036 10293 2044
rect 10976 2044 10984 2073
rect 11007 2056 11033 2064
rect 11107 2056 11153 2064
rect 11207 2056 11333 2064
rect 11587 2056 11633 2064
rect 12007 2056 12093 2064
rect 10976 2036 10993 2044
rect 11127 2036 11353 2044
rect 11367 2036 11533 2044
rect 11967 2036 12213 2044
rect 7147 2016 7464 2024
rect 7487 2016 7593 2024
rect 7607 2016 7853 2024
rect 8067 2016 8213 2024
rect 8267 2016 10133 2024
rect 10147 2016 10413 2024
rect 10427 2016 10593 2024
rect 10607 2016 11233 2024
rect 11667 2016 12053 2024
rect 2467 1996 3513 2004
rect 3527 1996 4333 2004
rect 7407 1996 7493 2004
rect 7567 1996 7673 2004
rect 7787 1996 7833 2004
rect 7907 1996 7933 2004
rect 8007 1996 8233 2004
rect 9087 1996 9213 2004
rect 9227 1996 9493 2004
rect 9667 1996 9733 2004
rect 9787 1996 9953 2004
rect 10027 1996 10673 2004
rect 2387 1976 2413 1984
rect 5427 1976 5453 1984
rect 5467 1976 6473 1984
rect 7207 1976 7733 1984
rect 7807 1976 8373 1984
rect 8467 1976 8573 1984
rect 8987 1976 9293 1984
rect 9567 1976 9713 1984
rect 10067 1976 10113 1984
rect 1667 1956 1673 1964
rect 1687 1956 2393 1964
rect 2407 1956 2893 1964
rect 2907 1956 3033 1964
rect 3047 1956 3093 1964
rect 6747 1956 8713 1964
rect 8747 1956 8873 1964
rect 8887 1956 9633 1964
rect 9707 1956 9753 1964
rect 9827 1956 10193 1964
rect 4387 1936 7673 1944
rect 8167 1936 8253 1944
rect 8367 1936 9113 1944
rect 9407 1936 9793 1944
rect 9807 1936 10093 1944
rect 2087 1916 2133 1924
rect 2147 1916 5133 1924
rect 7447 1916 8433 1924
rect 8916 1916 10853 1924
rect 7587 1896 7993 1904
rect 8916 1904 8924 1916
rect 11467 1916 11553 1924
rect 8147 1896 8924 1904
rect 8947 1896 9753 1904
rect 9807 1896 9933 1904
rect 9967 1896 10213 1904
rect 11087 1896 11693 1904
rect 6247 1876 6273 1884
rect 6527 1876 6613 1884
rect 7407 1876 7713 1884
rect 7747 1876 8153 1884
rect 8587 1876 8633 1884
rect 9247 1876 9533 1884
rect 9547 1876 10233 1884
rect 1827 1856 2893 1864
rect 3407 1856 3433 1864
rect 6247 1856 7873 1864
rect 7947 1856 8113 1864
rect 8607 1856 8693 1864
rect 8727 1856 9033 1864
rect 9047 1856 9093 1864
rect 9127 1856 9433 1864
rect 9487 1856 9513 1864
rect 9567 1856 9613 1864
rect 9987 1856 11213 1864
rect 11407 1856 11433 1864
rect 11487 1856 11533 1864
rect 2107 1836 3113 1844
rect 5607 1836 5633 1844
rect 5747 1836 7213 1844
rect 7327 1836 7953 1844
rect 8207 1836 10013 1844
rect 10387 1836 10513 1844
rect 10527 1836 10713 1844
rect 10927 1836 11133 1844
rect 11427 1836 11513 1844
rect 11847 1836 11933 1844
rect 327 1816 593 1824
rect 747 1816 793 1824
rect 1827 1816 2153 1824
rect 2967 1816 3053 1824
rect 3667 1816 3713 1824
rect 5347 1816 5593 1824
rect 5627 1816 5673 1824
rect 5767 1816 5793 1824
rect 6207 1816 6933 1824
rect 6947 1816 7033 1824
rect 7167 1816 7433 1824
rect 7827 1816 8073 1824
rect 8107 1816 8173 1824
rect 8287 1816 8333 1824
rect 8487 1816 9253 1824
rect 9367 1816 9453 1824
rect 9687 1816 10033 1824
rect 10087 1816 10233 1824
rect 10707 1816 10973 1824
rect 10987 1816 11033 1824
rect 11387 1816 11433 1824
rect 347 1796 493 1804
rect 867 1796 1213 1804
rect 1587 1796 1713 1804
rect 2107 1796 2193 1804
rect 2387 1796 2433 1804
rect 2827 1796 2913 1804
rect 3467 1796 3513 1804
rect 3676 1796 4173 1804
rect 156 1784 164 1793
rect 3676 1787 3684 1796
rect 4836 1796 5373 1804
rect 147 1776 164 1784
rect 527 1776 673 1784
rect 727 1776 873 1784
rect 2047 1776 2233 1784
rect 2247 1776 2733 1784
rect 2747 1776 2873 1784
rect 2947 1776 3133 1784
rect 3727 1776 3753 1784
rect 3907 1776 4233 1784
rect 4327 1776 4553 1784
rect 4607 1776 4813 1784
rect 4836 1784 4844 1796
rect 5387 1796 5553 1804
rect 5567 1796 5693 1804
rect 5847 1796 6004 1804
rect 5996 1787 6004 1796
rect 6027 1796 6184 1804
rect 6176 1787 6184 1796
rect 6407 1796 6564 1804
rect 6556 1787 6564 1796
rect 6807 1796 6953 1804
rect 7107 1796 7133 1804
rect 7987 1796 8473 1804
rect 8556 1796 8713 1804
rect 8556 1787 8564 1796
rect 9007 1796 9133 1804
rect 9147 1796 9213 1804
rect 9487 1796 9633 1804
rect 9667 1796 9753 1804
rect 9776 1796 9833 1804
rect 4827 1776 4844 1784
rect 4867 1776 4913 1784
rect 5027 1776 5173 1784
rect 5187 1776 5473 1784
rect 5507 1776 5533 1784
rect 5587 1776 5633 1784
rect 6627 1776 6773 1784
rect 6907 1776 7153 1784
rect 7227 1776 7333 1784
rect 7387 1776 7533 1784
rect 7547 1776 7713 1784
rect 7767 1776 7793 1784
rect 7887 1776 7953 1784
rect 7967 1776 8273 1784
rect 8367 1776 8533 1784
rect 8956 1784 8964 1793
rect 8947 1776 8964 1784
rect 9607 1776 9653 1784
rect 9776 1784 9784 1796
rect 10287 1796 10653 1804
rect 10807 1796 10873 1804
rect 10907 1796 11053 1804
rect 11476 1804 11484 1813
rect 11287 1796 11484 1804
rect 11667 1796 11793 1804
rect 9767 1776 9784 1784
rect 9867 1776 10053 1784
rect 10347 1776 10493 1784
rect 11207 1776 11213 1784
rect 11227 1776 11313 1784
rect 11407 1776 11453 1784
rect 11647 1776 11693 1784
rect 11707 1776 11733 1784
rect 11747 1776 11773 1784
rect 367 1756 853 1764
rect 907 1756 1013 1764
rect 1307 1756 1613 1764
rect 2567 1756 3013 1764
rect 4207 1756 4453 1764
rect 5407 1756 5453 1764
rect 5707 1756 6033 1764
rect 6047 1756 6193 1764
rect 6467 1756 6573 1764
rect 6707 1756 6753 1764
rect 6947 1756 7293 1764
rect 7447 1756 7553 1764
rect 7727 1756 8313 1764
rect 8527 1756 8553 1764
rect 8707 1756 8733 1764
rect 8807 1756 9033 1764
rect 9127 1756 9193 1764
rect 9227 1756 9673 1764
rect 9687 1756 10453 1764
rect 10507 1756 11593 1764
rect 11767 1756 11813 1764
rect 467 1736 893 1744
rect 2287 1736 3493 1744
rect 4987 1736 5713 1744
rect 6427 1736 6513 1744
rect 6607 1736 6973 1744
rect 7587 1736 7613 1744
rect 7767 1736 7833 1744
rect 7907 1736 7933 1744
rect 8087 1736 8413 1744
rect 8447 1736 8813 1744
rect 8827 1736 8893 1744
rect 8947 1736 9373 1744
rect 9467 1736 9613 1744
rect 10707 1736 12033 1744
rect 547 1716 1073 1724
rect 3087 1716 3993 1724
rect 6207 1716 6673 1724
rect 7007 1716 8313 1724
rect 8347 1716 8853 1724
rect 9127 1716 9173 1724
rect 9707 1716 9853 1724
rect 10087 1716 10113 1724
rect 10127 1716 10293 1724
rect 10307 1716 12113 1724
rect 927 1696 1853 1704
rect 3507 1696 3993 1704
rect 5967 1696 8773 1704
rect 8787 1696 8913 1704
rect 8927 1696 9913 1704
rect 11147 1696 11833 1704
rect 11847 1696 12073 1704
rect 2547 1676 2613 1684
rect 5587 1676 5733 1684
rect 6147 1676 7413 1684
rect 7607 1676 7644 1684
rect 167 1656 373 1664
rect 387 1656 1313 1664
rect 1467 1656 2033 1664
rect 2427 1656 2473 1664
rect 3767 1656 4173 1664
rect 4567 1656 5033 1664
rect 5047 1656 5273 1664
rect 5627 1656 5733 1664
rect 5747 1656 7173 1664
rect 7187 1656 7613 1664
rect 7636 1664 7644 1676
rect 7816 1676 7913 1684
rect 7816 1664 7824 1676
rect 8007 1676 8533 1684
rect 8547 1676 9013 1684
rect 9107 1676 9573 1684
rect 11087 1676 11253 1684
rect 7636 1656 7824 1664
rect 7867 1656 8273 1664
rect 8327 1656 8993 1664
rect 9007 1656 9093 1664
rect 9307 1656 9373 1664
rect 9607 1656 9873 1664
rect 10127 1656 10913 1664
rect 807 1636 1613 1644
rect 1627 1636 2013 1644
rect 2027 1636 2113 1644
rect 2227 1636 2413 1644
rect 3707 1636 3893 1644
rect 4567 1636 5173 1644
rect 5247 1636 5533 1644
rect 5547 1636 6213 1644
rect 6907 1636 6993 1644
rect 7196 1636 7664 1644
rect 667 1616 773 1624
rect 947 1616 1033 1624
rect 1607 1616 1813 1624
rect 1827 1616 2133 1624
rect 2147 1616 2213 1624
rect 2407 1616 2433 1624
rect 2647 1616 2713 1624
rect 2727 1616 2753 1624
rect 2787 1616 2833 1624
rect 2927 1616 3013 1624
rect 3347 1616 3413 1624
rect 3427 1616 3613 1624
rect 3887 1616 3933 1624
rect 4167 1616 4373 1624
rect 4407 1616 4873 1624
rect 4887 1616 4933 1624
rect 5067 1616 5373 1624
rect 5387 1616 5693 1624
rect 7196 1624 7204 1636
rect 6367 1616 7204 1624
rect 7227 1616 7273 1624
rect 7656 1624 7664 1636
rect 7687 1636 10253 1644
rect 10467 1636 10493 1644
rect 11607 1636 11653 1644
rect 11687 1636 11753 1644
rect 7656 1616 8953 1624
rect 8987 1616 9353 1624
rect 9567 1616 9693 1624
rect 9767 1616 9833 1624
rect 10367 1616 10613 1624
rect 10687 1616 11033 1624
rect 11667 1616 11933 1624
rect 11987 1616 12033 1624
rect 967 1596 1064 1604
rect 47 1576 113 1584
rect 287 1576 373 1584
rect 387 1576 553 1584
rect 627 1576 793 1584
rect 1056 1584 1064 1596
rect 1087 1596 1273 1604
rect 1496 1596 1633 1604
rect 1496 1587 1504 1596
rect 1707 1596 1953 1604
rect 2236 1604 2244 1613
rect 2067 1596 2244 1604
rect 2607 1596 2673 1604
rect 3476 1596 3633 1604
rect 3476 1587 3484 1596
rect 3707 1596 3864 1604
rect 3856 1587 3864 1596
rect 4607 1596 4693 1604
rect 4767 1596 4904 1604
rect 4896 1587 4904 1596
rect 5287 1596 5393 1604
rect 5547 1596 5673 1604
rect 5807 1596 5913 1604
rect 5927 1596 5993 1604
rect 6007 1596 6293 1604
rect 6507 1596 6573 1604
rect 6747 1596 6773 1604
rect 6787 1596 6913 1604
rect 7087 1596 7244 1604
rect 1056 1576 1113 1584
rect 1596 1576 2393 1584
rect 607 1556 953 1564
rect 1147 1556 1293 1564
rect 1596 1564 1604 1576
rect 2947 1576 2973 1584
rect 5487 1576 5713 1584
rect 6316 1584 6324 1593
rect 6127 1576 6324 1584
rect 6347 1576 6373 1584
rect 6527 1576 6593 1584
rect 6696 1584 6704 1593
rect 6696 1576 7053 1584
rect 7107 1576 7213 1584
rect 7236 1584 7244 1596
rect 7307 1596 7393 1604
rect 7507 1596 7593 1604
rect 7707 1596 7733 1604
rect 7907 1596 7953 1604
rect 9207 1596 9313 1604
rect 9327 1596 9393 1604
rect 9407 1596 9544 1604
rect 7236 1576 7333 1584
rect 7407 1576 7453 1584
rect 7656 1584 7664 1593
rect 7487 1576 7664 1584
rect 7787 1576 7833 1584
rect 7887 1576 8053 1584
rect 8067 1576 8133 1584
rect 8187 1576 8333 1584
rect 8376 1584 8384 1593
rect 8376 1576 8633 1584
rect 8647 1576 8693 1584
rect 9227 1576 9273 1584
rect 9287 1576 9413 1584
rect 9536 1584 9544 1596
rect 9567 1596 9624 1604
rect 9536 1576 9573 1584
rect 9616 1584 9624 1596
rect 9647 1596 9753 1604
rect 10027 1596 10093 1604
rect 11027 1596 11093 1604
rect 11196 1596 11233 1604
rect 9616 1576 9733 1584
rect 10116 1576 10293 1584
rect 1307 1556 1604 1564
rect 1627 1556 1673 1564
rect 3267 1556 3653 1564
rect 4327 1556 4453 1564
rect 4467 1556 4713 1564
rect 4727 1556 4953 1564
rect 5107 1556 5793 1564
rect 6507 1556 6573 1564
rect 6587 1556 6713 1564
rect 6727 1556 6833 1564
rect 7207 1556 7293 1564
rect 7747 1556 7853 1564
rect 7887 1556 8013 1564
rect 8147 1556 8393 1564
rect 9067 1556 9253 1564
rect 9627 1556 9973 1564
rect 10116 1564 10124 1576
rect 10507 1576 10633 1584
rect 11196 1584 11204 1596
rect 11267 1596 11333 1604
rect 11347 1596 11693 1604
rect 11807 1596 11993 1604
rect 11067 1576 11204 1584
rect 11227 1576 11293 1584
rect 11707 1576 11773 1584
rect 11827 1576 11953 1584
rect 10107 1556 10124 1564
rect 10147 1556 10173 1564
rect 10207 1556 10873 1564
rect 10887 1556 11373 1564
rect 11427 1556 11493 1564
rect 11627 1556 11653 1564
rect 11747 1556 12033 1564
rect 107 1536 153 1544
rect 167 1536 213 1544
rect 227 1536 893 1544
rect 1667 1536 1873 1544
rect 1887 1536 2273 1544
rect 3047 1536 3313 1544
rect 6407 1536 6473 1544
rect 6487 1536 6533 1544
rect 6547 1536 7233 1544
rect 7367 1536 8033 1544
rect 8047 1536 8213 1544
rect 8487 1536 8593 1544
rect 8807 1536 8973 1544
rect 9027 1536 9153 1544
rect 9167 1536 9233 1544
rect 9427 1536 9713 1544
rect 6716 1516 7733 1524
rect 6716 1504 6724 1516
rect 7767 1516 7893 1524
rect 7947 1516 8073 1524
rect 8087 1516 8313 1524
rect 8347 1516 8553 1524
rect 9007 1516 9753 1524
rect 10287 1516 10733 1524
rect 6187 1496 6733 1504
rect 7287 1496 9913 1504
rect 10547 1496 10613 1504
rect 1347 1476 1553 1484
rect 6667 1476 7153 1484
rect 7267 1476 7513 1484
rect 7687 1476 8993 1484
rect 9047 1476 9133 1484
rect 3067 1456 3133 1464
rect 5847 1456 7453 1464
rect 7487 1456 7773 1464
rect 7867 1456 8053 1464
rect 8707 1456 10253 1464
rect 10267 1456 10653 1464
rect 10667 1456 11293 1464
rect 47 1436 473 1444
rect 6027 1436 6053 1444
rect 6607 1436 7473 1444
rect 7927 1436 7933 1444
rect 7947 1436 8293 1444
rect 8307 1436 8593 1444
rect 9267 1436 9653 1444
rect 9667 1436 9713 1444
rect 9727 1436 10193 1444
rect 10227 1436 11553 1444
rect 2707 1416 3833 1424
rect 5987 1416 6533 1424
rect 7247 1416 8193 1424
rect 8227 1416 10553 1424
rect 10567 1416 11073 1424
rect 11087 1416 11373 1424
rect 11887 1416 11973 1424
rect 4467 1396 5273 1404
rect 5287 1396 5353 1404
rect 5827 1396 6373 1404
rect 7407 1396 7493 1404
rect 7807 1396 7973 1404
rect 8567 1396 8793 1404
rect 8807 1396 8953 1404
rect 9327 1396 10453 1404
rect 11907 1396 12033 1404
rect 1067 1376 2413 1384
rect 2447 1376 2573 1384
rect 2587 1376 3093 1384
rect 3107 1376 3193 1384
rect 3207 1376 3733 1384
rect 3747 1376 4453 1384
rect 4687 1376 4713 1384
rect 5887 1376 6173 1384
rect 6527 1376 6633 1384
rect 6767 1376 6913 1384
rect 7467 1376 7693 1384
rect 8027 1376 8933 1384
rect 10167 1376 10433 1384
rect 10487 1376 10513 1384
rect 10647 1376 10933 1384
rect 11487 1376 11533 1384
rect 11807 1376 12053 1384
rect 907 1356 1433 1364
rect 2287 1356 2633 1364
rect 3127 1356 3233 1364
rect 3267 1356 4533 1364
rect 4887 1356 5053 1364
rect 5207 1356 5253 1364
rect 5347 1356 5853 1364
rect 5987 1356 6593 1364
rect 6827 1356 7453 1364
rect 9067 1356 9533 1364
rect 9547 1356 9593 1364
rect 11287 1356 11904 1364
rect 1047 1336 1793 1344
rect 1967 1336 2093 1344
rect 2467 1336 3153 1344
rect 3187 1336 3233 1344
rect 4207 1336 4273 1344
rect 4967 1336 5013 1344
rect 5087 1336 5493 1344
rect 6087 1336 6113 1344
rect 6436 1336 6633 1344
rect 187 1316 613 1324
rect 667 1316 693 1324
rect 727 1316 1493 1324
rect 2027 1316 2133 1324
rect 2367 1316 2384 1324
rect 2376 1307 2384 1316
rect 2507 1316 2533 1324
rect 3287 1316 3353 1324
rect 3607 1316 3693 1324
rect 3787 1316 4073 1324
rect 4167 1316 4253 1324
rect 4607 1316 4653 1324
rect 4907 1316 4993 1324
rect 5296 1316 5433 1324
rect 367 1296 633 1304
rect 807 1296 933 1304
rect 1607 1296 1973 1304
rect 2287 1296 2333 1304
rect 2487 1296 2553 1304
rect 2607 1296 2693 1304
rect 3127 1296 3173 1304
rect 3227 1296 3253 1304
rect 3727 1296 3793 1304
rect 4096 1296 5073 1304
rect 4096 1287 4104 1296
rect 687 1276 873 1284
rect 927 1276 1733 1284
rect 2147 1276 2353 1284
rect 3147 1276 3173 1284
rect 3196 1276 3393 1284
rect 1827 1256 2173 1264
rect 2347 1256 2493 1264
rect 2627 1256 2633 1264
rect 2647 1256 2753 1264
rect 3196 1264 3204 1276
rect 3407 1276 3473 1284
rect 4127 1276 4433 1284
rect 4487 1276 5213 1284
rect 5236 1284 5244 1313
rect 5296 1307 5304 1316
rect 6036 1324 6044 1333
rect 5887 1316 6044 1324
rect 6107 1316 6153 1324
rect 6167 1316 6273 1324
rect 6436 1324 6444 1336
rect 6707 1336 6773 1344
rect 7427 1336 7533 1344
rect 7787 1336 7893 1344
rect 8127 1336 8424 1344
rect 6427 1316 6444 1324
rect 6467 1316 6504 1324
rect 5407 1296 5573 1304
rect 5627 1296 5853 1304
rect 6387 1296 6433 1304
rect 6496 1287 6504 1316
rect 6687 1316 6753 1324
rect 7016 1316 7193 1324
rect 7016 1307 7024 1316
rect 7236 1324 7244 1333
rect 7236 1316 7604 1324
rect 6547 1296 6613 1304
rect 6847 1296 6953 1304
rect 6967 1296 6973 1304
rect 7187 1296 7253 1304
rect 7447 1296 7513 1304
rect 7527 1296 7573 1304
rect 7596 1304 7604 1316
rect 7627 1316 8193 1324
rect 8247 1316 8353 1324
rect 8416 1324 8424 1336
rect 8467 1336 8933 1344
rect 9027 1336 9153 1344
rect 9267 1336 9333 1344
rect 9367 1336 9513 1344
rect 10436 1336 10493 1344
rect 8416 1316 8553 1324
rect 8607 1316 8673 1324
rect 8727 1316 9053 1324
rect 9187 1316 9313 1324
rect 9407 1316 9513 1324
rect 9987 1316 10073 1324
rect 10087 1316 10313 1324
rect 10436 1324 10444 1336
rect 10507 1336 10833 1344
rect 10847 1336 10933 1344
rect 11227 1336 11353 1344
rect 11527 1336 11664 1344
rect 11656 1327 11664 1336
rect 11687 1336 11753 1344
rect 11896 1344 11904 1356
rect 11927 1356 11953 1364
rect 11896 1336 11913 1344
rect 10367 1316 10444 1324
rect 10467 1316 10513 1324
rect 11047 1316 11173 1324
rect 11187 1316 11324 1324
rect 11316 1307 11324 1316
rect 11527 1316 11573 1324
rect 11587 1316 11593 1324
rect 11667 1316 11853 1324
rect 7596 1296 7753 1304
rect 7867 1296 7913 1304
rect 8167 1296 8333 1304
rect 8387 1296 8453 1304
rect 8627 1296 8713 1304
rect 9127 1296 9193 1304
rect 9627 1296 9713 1304
rect 9927 1296 9953 1304
rect 10147 1296 10213 1304
rect 10347 1296 10413 1304
rect 10567 1296 10713 1304
rect 10747 1296 10873 1304
rect 10887 1296 11273 1304
rect 11576 1296 11673 1304
rect 5236 1276 5293 1284
rect 5327 1276 5413 1284
rect 5827 1276 6093 1284
rect 6787 1276 7033 1284
rect 7047 1276 7433 1284
rect 7507 1276 7593 1284
rect 7707 1276 7793 1284
rect 7867 1276 7953 1284
rect 7967 1276 8093 1284
rect 8147 1276 8173 1284
rect 8207 1276 9273 1284
rect 10087 1276 10153 1284
rect 10307 1276 10673 1284
rect 11067 1276 11153 1284
rect 11267 1276 11353 1284
rect 11367 1276 11413 1284
rect 11576 1284 11584 1296
rect 12096 1304 12104 1313
rect 11687 1296 12104 1304
rect 11427 1276 11584 1284
rect 11607 1276 11693 1284
rect 11907 1276 12013 1284
rect 12027 1276 12113 1284
rect 3007 1256 3204 1264
rect 3387 1256 3433 1264
rect 3447 1256 3873 1264
rect 4707 1256 5033 1264
rect 5047 1256 5233 1264
rect 5267 1256 5333 1264
rect 5967 1256 6373 1264
rect 6387 1256 6633 1264
rect 6707 1256 7233 1264
rect 7347 1256 7413 1264
rect 7907 1256 8033 1264
rect 8596 1256 8733 1264
rect 1547 1236 4613 1244
rect 5907 1236 6213 1244
rect 6267 1236 6653 1244
rect 6667 1236 7273 1244
rect 7807 1236 7873 1244
rect 8596 1244 8604 1256
rect 8747 1256 9073 1264
rect 9287 1256 9393 1264
rect 9527 1256 10973 1264
rect 10987 1256 11533 1264
rect 11647 1256 11713 1264
rect 8067 1236 8604 1244
rect 8907 1236 9073 1244
rect 9087 1236 9213 1244
rect 9247 1236 9553 1244
rect 9567 1236 9773 1244
rect 9787 1236 10033 1244
rect 10307 1236 10353 1244
rect 10727 1236 11193 1244
rect 11347 1236 11613 1244
rect 11627 1236 11833 1244
rect 11847 1236 11993 1244
rect 12007 1236 12073 1244
rect 1467 1216 4053 1224
rect 6367 1216 9313 1224
rect 9327 1216 9753 1224
rect 9767 1216 10113 1224
rect 10587 1216 11444 1224
rect 1787 1196 4833 1204
rect 5727 1196 5853 1204
rect 5867 1196 5893 1204
rect 5907 1196 6333 1204
rect 6767 1196 6853 1204
rect 7027 1196 7373 1204
rect 7647 1196 8273 1204
rect 8287 1196 8593 1204
rect 8607 1196 8753 1204
rect 9907 1196 9933 1204
rect 9947 1196 10573 1204
rect 10927 1196 10953 1204
rect 11436 1204 11444 1216
rect 11467 1216 11773 1224
rect 11787 1216 11873 1224
rect 11947 1216 11973 1224
rect 11436 1196 11493 1204
rect 11507 1196 11573 1204
rect 1587 1176 1973 1184
rect 2087 1176 2993 1184
rect 3487 1176 3553 1184
rect 3567 1176 4953 1184
rect 5207 1176 5953 1184
rect 6147 1176 7393 1184
rect 7467 1176 7733 1184
rect 7847 1176 7913 1184
rect 8487 1176 9413 1184
rect 9447 1176 9733 1184
rect 10087 1176 10393 1184
rect 11127 1176 11873 1184
rect 147 1156 193 1164
rect 1347 1156 1453 1164
rect 2667 1156 2713 1164
rect 3367 1156 3673 1164
rect 4227 1156 4273 1164
rect 6187 1156 6453 1164
rect 6467 1156 6533 1164
rect 6547 1156 6813 1164
rect 6887 1156 7213 1164
rect 7247 1156 8513 1164
rect 8987 1156 9113 1164
rect 9227 1156 9253 1164
rect 9267 1156 9453 1164
rect 9707 1156 9773 1164
rect 10047 1156 10533 1164
rect 187 1136 233 1144
rect 907 1136 1033 1144
rect 1247 1136 1513 1144
rect 1527 1136 1853 1144
rect 1867 1136 1873 1144
rect 2167 1136 2293 1144
rect 2487 1136 2513 1144
rect 3667 1136 3713 1144
rect 3927 1136 3953 1144
rect 4207 1136 4433 1144
rect 4447 1136 4533 1144
rect 4627 1136 4673 1144
rect 4807 1136 4833 1144
rect 4867 1136 5073 1144
rect 5387 1136 5433 1144
rect 5687 1136 6273 1144
rect 6287 1136 6693 1144
rect 6707 1136 7093 1144
rect 7107 1136 7133 1144
rect 7727 1136 7753 1144
rect 7787 1136 7913 1144
rect 8327 1136 9693 1144
rect 9867 1136 9953 1144
rect 9987 1136 9993 1144
rect 10007 1136 10024 1144
rect 10407 1136 10433 1144
rect 10587 1136 10633 1144
rect 11087 1136 11113 1144
rect 11447 1136 11973 1144
rect 707 1116 793 1124
rect 807 1116 913 1124
rect 1007 1116 1113 1124
rect 1227 1116 1293 1124
rect 1347 1116 1533 1124
rect 2067 1116 2133 1124
rect 2907 1116 3753 1124
rect 3927 1116 4153 1124
rect 4416 1116 4553 1124
rect 4416 1107 4424 1116
rect 4567 1116 4753 1124
rect 5036 1116 5213 1124
rect 5036 1107 5044 1116
rect 5407 1116 5633 1124
rect 5647 1116 5753 1124
rect 5927 1116 6084 1124
rect 107 1096 153 1104
rect 207 1096 333 1104
rect 387 1096 473 1104
rect 527 1096 733 1104
rect 767 1096 853 1104
rect 967 1096 1313 1104
rect 1967 1096 2153 1104
rect 2527 1096 2564 1104
rect 747 1076 1053 1084
rect 1107 1076 1473 1084
rect 2556 1084 2564 1096
rect 2727 1096 2913 1104
rect 2927 1096 3033 1104
rect 3047 1096 3113 1104
rect 3147 1096 3313 1104
rect 3507 1096 3633 1104
rect 3687 1096 3813 1104
rect 4027 1096 4253 1104
rect 5387 1096 5933 1104
rect 5947 1096 5973 1104
rect 6076 1104 6084 1116
rect 6107 1116 6233 1124
rect 6307 1116 6384 1124
rect 6076 1096 6173 1104
rect 6327 1096 6353 1104
rect 6376 1104 6384 1116
rect 6907 1116 7053 1124
rect 7287 1116 7333 1124
rect 7507 1116 7673 1124
rect 8007 1116 8093 1124
rect 8147 1116 8253 1124
rect 9107 1116 9533 1124
rect 9587 1116 9633 1124
rect 9687 1116 9813 1124
rect 9836 1116 10713 1124
rect 6376 1096 6433 1104
rect 6607 1096 6653 1104
rect 6836 1104 6844 1113
rect 6667 1096 6844 1104
rect 7047 1096 7073 1104
rect 7407 1096 7513 1104
rect 7707 1096 7773 1104
rect 7876 1104 7884 1113
rect 7876 1096 8033 1104
rect 8087 1096 8393 1104
rect 8427 1096 8453 1104
rect 8647 1096 8693 1104
rect 8816 1104 8824 1113
rect 8816 1096 8993 1104
rect 9016 1104 9024 1113
rect 9016 1096 9213 1104
rect 9836 1104 9844 1116
rect 11087 1116 11253 1124
rect 11647 1116 11673 1124
rect 11987 1116 12013 1124
rect 9567 1096 9844 1104
rect 9947 1096 10133 1104
rect 10167 1096 10333 1104
rect 10347 1096 10513 1104
rect 10947 1096 11513 1104
rect 11627 1096 11653 1104
rect 11687 1096 11733 1104
rect 12007 1096 12033 1104
rect 2556 1076 2693 1084
rect 2747 1076 2773 1084
rect 2787 1076 2933 1084
rect 2947 1076 3133 1084
rect 3147 1076 3193 1084
rect 3307 1076 3413 1084
rect 3627 1076 3653 1084
rect 3907 1076 4973 1084
rect 5047 1076 5553 1084
rect 6827 1076 6853 1084
rect 7127 1076 8204 1084
rect 507 1056 533 1064
rect 547 1056 593 1064
rect 867 1056 1013 1064
rect 1027 1056 1253 1064
rect 2536 1064 2544 1073
rect 2536 1056 2713 1064
rect 3127 1056 3173 1064
rect 3247 1056 3313 1064
rect 4227 1056 4593 1064
rect 4607 1056 4813 1064
rect 4827 1056 4853 1064
rect 5007 1056 5273 1064
rect 7367 1056 7453 1064
rect 8196 1064 8204 1076
rect 8227 1076 8293 1084
rect 8547 1076 8833 1084
rect 8867 1076 8953 1084
rect 9247 1076 9524 1084
rect 8196 1056 8573 1064
rect 8887 1056 9453 1064
rect 9516 1064 9524 1076
rect 9547 1076 9673 1084
rect 9707 1076 11093 1084
rect 11107 1076 11153 1084
rect 11167 1076 11413 1084
rect 11707 1076 11753 1084
rect 11807 1076 11853 1084
rect 11907 1076 11953 1084
rect 9516 1056 9753 1064
rect 9987 1056 10033 1064
rect 11656 1064 11664 1073
rect 10707 1056 11793 1064
rect 547 1036 693 1044
rect 1127 1036 1233 1044
rect 1447 1036 1533 1044
rect 3947 1036 4213 1044
rect 4547 1036 5313 1044
rect 5327 1036 5433 1044
rect 7747 1036 8193 1044
rect 8476 1036 10273 1044
rect 3207 1016 3613 1024
rect 7187 1016 8073 1024
rect 8476 1024 8484 1036
rect 10747 1036 11453 1044
rect 11467 1036 11733 1044
rect 8107 1016 8484 1024
rect 8687 1016 9673 1024
rect 9687 1016 10233 1024
rect 10747 1016 10893 1024
rect 10907 1016 11133 1024
rect 1807 996 2113 1004
rect 2587 996 3253 1004
rect 7907 996 8773 1004
rect 8787 996 10233 1004
rect 10247 996 10693 1004
rect 10927 996 10953 1004
rect 7507 976 7533 984
rect 7547 976 8533 984
rect 8647 976 10313 984
rect 947 956 1073 964
rect 1087 956 1213 964
rect 7427 956 7533 964
rect 8027 956 9333 964
rect 9387 956 9433 964
rect 9487 956 9613 964
rect 1767 936 1853 944
rect 5467 936 6833 944
rect 6847 936 8473 944
rect 8547 936 10353 944
rect 10647 936 11333 944
rect 11347 936 11473 944
rect 5167 916 7713 924
rect 8307 916 10693 924
rect 10707 916 10773 924
rect 3047 896 3493 904
rect 3507 896 3813 904
rect 4867 896 5213 904
rect 7847 896 8313 904
rect 8707 896 9473 904
rect 9767 896 9833 904
rect 9927 896 11933 904
rect 3467 876 3513 884
rect 3587 876 3873 884
rect 3987 876 4013 884
rect 4267 876 4473 884
rect 4487 876 5264 884
rect 267 856 753 864
rect 987 856 1033 864
rect 1307 856 1633 864
rect 1647 856 1733 864
rect 1747 856 2033 864
rect 2287 856 2333 864
rect 2347 856 2473 864
rect 2787 856 2913 864
rect 2936 856 3033 864
rect 167 836 393 844
rect 587 836 744 844
rect 736 827 744 836
rect 967 836 993 844
rect 1407 836 1453 844
rect 1467 836 1473 844
rect 1567 836 1793 844
rect 2056 844 2064 853
rect 2936 847 2944 856
rect 3336 856 3513 864
rect 3336 847 3344 856
rect 3567 856 3613 864
rect 3627 856 3893 864
rect 4007 856 4033 864
rect 4167 856 4253 864
rect 4267 856 4293 864
rect 4347 856 4513 864
rect 4527 856 4613 864
rect 4667 856 4713 864
rect 4907 856 5053 864
rect 5256 864 5264 876
rect 5287 876 5713 884
rect 7387 876 7473 884
rect 7647 876 8013 884
rect 8187 876 8593 884
rect 8927 876 9933 884
rect 10967 876 11773 884
rect 11947 876 12033 884
rect 5107 856 5244 864
rect 5256 856 5473 864
rect 5236 847 5244 856
rect 5787 856 7513 864
rect 7527 856 7973 864
rect 7987 856 8093 864
rect 9267 856 9393 864
rect 9807 856 10013 864
rect 10207 856 10773 864
rect 10787 856 10853 864
rect 11107 856 11153 864
rect 11787 856 11873 864
rect 2007 836 2064 844
rect 2327 836 2373 844
rect 2387 836 2433 844
rect 2487 836 2533 844
rect 2767 836 2893 844
rect 2987 836 3133 844
rect 3507 836 3533 844
rect 3587 836 3993 844
rect 4847 836 4913 844
rect 6427 836 7013 844
rect 7067 836 7193 844
rect 7327 836 7433 844
rect 7807 836 7893 844
rect 8007 836 8133 844
rect 8167 836 8233 844
rect 8347 836 8373 844
rect 8527 836 8553 844
rect 8607 836 8653 844
rect 8676 836 8933 844
rect 1587 816 1613 824
rect 1687 816 2013 824
rect 2196 824 2204 833
rect 2067 816 2204 824
rect 2407 816 2453 824
rect 2607 816 3053 824
rect 3187 816 3253 824
rect 3267 816 3373 824
rect 3787 816 3853 824
rect 3927 816 4253 824
rect 4267 816 4593 824
rect 4607 816 4673 824
rect 4727 816 4813 824
rect 4827 816 5033 824
rect 5047 816 5053 824
rect 5567 816 5613 824
rect 5667 816 5713 824
rect 5767 816 5793 824
rect 6047 816 6073 824
rect 6307 816 6513 824
rect 6647 816 6773 824
rect 6787 816 6793 824
rect 7347 816 7373 824
rect 7467 816 7493 824
rect 7827 816 8173 824
rect 8676 824 8684 836
rect 8956 836 8973 844
rect 8956 824 8964 836
rect 9027 836 9153 844
rect 9667 836 9793 844
rect 9847 836 9984 844
rect 8587 816 8684 824
rect 8936 816 8964 824
rect 8936 807 8944 816
rect 9087 816 9133 824
rect 9387 816 9553 824
rect 9596 824 9604 833
rect 9596 816 9773 824
rect 9976 824 9984 836
rect 10007 836 10253 844
rect 11007 836 11053 844
rect 11467 836 11713 844
rect 9976 816 10033 824
rect 10307 816 10373 824
rect 10607 816 11193 824
rect 11687 816 11693 824
rect 11707 816 11893 824
rect 11907 816 12093 824
rect 187 796 233 804
rect 247 796 333 804
rect 367 796 393 804
rect 407 796 513 804
rect 787 796 853 804
rect 1787 796 2073 804
rect 2187 796 2733 804
rect 2747 796 3133 804
rect 3167 796 3233 804
rect 3387 796 4053 804
rect 4887 796 4993 804
rect 6067 796 6253 804
rect 6507 796 6813 804
rect 6867 796 7024 804
rect 487 776 893 784
rect 907 776 1093 784
rect 1607 776 1813 784
rect 1867 776 2353 784
rect 3047 776 3593 784
rect 4947 776 5073 784
rect 6127 776 6993 784
rect 7016 784 7024 796
rect 7047 796 7353 804
rect 7567 796 7653 804
rect 7907 796 8393 804
rect 8507 796 8573 804
rect 8967 796 9013 804
rect 9587 796 9633 804
rect 9747 796 9993 804
rect 10667 796 10753 804
rect 10927 796 10953 804
rect 7016 776 7613 784
rect 8087 776 8593 784
rect 8807 776 9913 784
rect 10236 776 10973 784
rect 567 756 653 764
rect 867 756 2553 764
rect 6267 756 6653 764
rect 7067 756 7253 764
rect 7427 756 7513 764
rect 8367 756 8393 764
rect 10236 764 10244 776
rect 9007 756 10244 764
rect 10267 756 12053 764
rect 12067 756 12073 764
rect 1187 736 1293 744
rect 6607 736 6913 744
rect 6927 736 7173 744
rect 7187 736 8633 744
rect 8727 736 8813 744
rect 8827 736 8913 744
rect 9467 736 9973 744
rect 9987 736 10293 744
rect 10307 736 10733 744
rect 10747 736 11353 744
rect 11367 736 11393 744
rect 327 716 593 724
rect 1667 716 1713 724
rect 3027 716 3973 724
rect 3987 716 4233 724
rect 6007 716 6853 724
rect 6867 716 6913 724
rect 7267 716 7453 724
rect 7467 716 7593 724
rect 7607 716 7633 724
rect 7847 716 9853 724
rect 9947 716 10513 724
rect 10547 716 10813 724
rect 10827 716 10873 724
rect 10987 716 11013 724
rect 11487 716 11533 724
rect 11547 716 11653 724
rect 11667 716 11853 724
rect 11867 716 11913 724
rect 2227 696 2253 704
rect 4707 696 4813 704
rect 5167 696 5753 704
rect 5767 696 6273 704
rect 6627 696 8553 704
rect 8627 696 9024 704
rect 287 676 373 684
rect 387 676 493 684
rect 507 676 873 684
rect 887 676 1013 684
rect 1027 676 1373 684
rect 2227 676 2633 684
rect 3027 676 3173 684
rect 3887 676 4453 684
rect 4467 676 5393 684
rect 6467 676 7553 684
rect 7627 676 7733 684
rect 7787 676 8193 684
rect 8207 676 8613 684
rect 8727 676 8753 684
rect 9016 684 9024 696
rect 9047 696 9433 704
rect 9447 696 10233 704
rect 10567 696 10913 704
rect 11036 696 11853 704
rect 9007 676 9113 684
rect 9187 676 9313 684
rect 10007 676 10253 684
rect 11036 684 11044 696
rect 10707 676 11044 684
rect 11067 676 11493 684
rect 167 656 253 664
rect 1007 656 1033 664
rect 1087 656 1313 664
rect 2387 656 2533 664
rect 2787 656 2833 664
rect 3007 656 3493 664
rect 3507 656 3713 664
rect 3747 656 3884 664
rect 107 636 193 644
rect 1287 636 1333 644
rect 1387 636 1433 644
rect 1447 636 1773 644
rect 1967 636 2013 644
rect 2587 636 2724 644
rect 1047 616 1133 624
rect 1767 616 2133 624
rect 2367 616 2433 624
rect 2447 616 2553 624
rect 2716 624 2724 636
rect 2747 636 2933 644
rect 3527 636 3753 644
rect 3876 644 3884 656
rect 3907 656 3973 664
rect 4127 656 4273 664
rect 4307 656 4913 664
rect 4927 656 4973 664
rect 5007 656 5293 664
rect 5427 656 5473 664
rect 6387 656 6453 664
rect 6847 656 7013 664
rect 7547 656 7633 664
rect 7727 656 7813 664
rect 7827 656 8293 664
rect 8327 656 8413 664
rect 8627 656 8733 664
rect 9227 656 9273 664
rect 9367 656 9473 664
rect 9527 656 9573 664
rect 9607 656 9713 664
rect 9727 656 9933 664
rect 10067 656 10093 664
rect 10167 656 10673 664
rect 10687 656 10933 664
rect 10947 656 11073 664
rect 11087 656 11153 664
rect 11167 656 11253 664
rect 11367 656 11533 664
rect 11547 656 11753 664
rect 3876 636 4093 644
rect 4107 636 4173 644
rect 4267 636 4313 644
rect 4627 636 4793 644
rect 4807 636 5533 644
rect 5547 636 5633 644
rect 5807 636 6033 644
rect 6427 636 6533 644
rect 6547 636 6873 644
rect 7216 636 7373 644
rect 2716 616 2753 624
rect 2887 616 2973 624
rect 4147 616 4433 624
rect 4607 616 4773 624
rect 5627 616 5813 624
rect 6167 616 6253 624
rect 6407 616 6573 624
rect 6667 616 6733 624
rect 6827 616 6973 624
rect 7216 624 7224 636
rect 7007 616 7224 624
rect 827 596 1053 604
rect 1067 596 1393 604
rect 1407 596 1813 604
rect 2567 596 2793 604
rect 3007 596 3433 604
rect 4447 596 4593 604
rect 4847 596 5033 604
rect 5367 596 5593 604
rect 5647 596 5673 604
rect 6067 596 6193 604
rect 6247 596 6593 604
rect 6647 596 6793 604
rect 6887 596 7033 604
rect 7056 604 7064 616
rect 7247 616 7393 624
rect 7436 624 7444 653
rect 7587 636 7693 644
rect 7707 636 7773 644
rect 7787 636 7853 644
rect 7887 636 7933 644
rect 8167 636 8204 644
rect 7427 616 7444 624
rect 7627 616 7653 624
rect 7967 616 8173 624
rect 8196 624 8204 636
rect 8227 636 8373 644
rect 8667 636 8793 644
rect 8196 616 8273 624
rect 8676 624 8684 636
rect 8807 636 8873 644
rect 9287 636 9333 644
rect 9387 636 9413 644
rect 9567 636 9773 644
rect 9927 636 10073 644
rect 10087 636 10093 644
rect 8347 616 8684 624
rect 8707 616 8733 624
rect 8787 616 8813 624
rect 8907 616 8973 624
rect 9136 624 9144 633
rect 10116 627 10124 653
rect 10147 636 10173 644
rect 10227 636 10333 644
rect 10367 636 11344 644
rect 9136 616 9313 624
rect 9367 616 9593 624
rect 9747 616 9873 624
rect 9967 616 9993 624
rect 10267 616 10313 624
rect 10487 616 10533 624
rect 10587 616 10613 624
rect 10907 616 11053 624
rect 11107 616 11313 624
rect 11336 624 11344 636
rect 11387 636 11733 644
rect 11747 636 11893 644
rect 11907 636 11973 644
rect 11336 616 11613 624
rect 11647 616 11693 624
rect 7056 596 7173 604
rect 7227 596 7833 604
rect 7867 596 7933 604
rect 8487 596 9153 604
rect 9427 596 9593 604
rect 9607 596 9693 604
rect 9707 596 10813 604
rect 10907 596 10953 604
rect 11007 596 11133 604
rect 11347 596 11373 604
rect 11627 596 11673 604
rect 11727 596 11753 604
rect 11887 596 11953 604
rect 11967 596 12033 604
rect 187 576 213 584
rect 227 576 793 584
rect 807 576 953 584
rect 967 576 1353 584
rect 1367 576 1393 584
rect 2487 576 2513 584
rect 2527 576 2953 584
rect 3367 576 3473 584
rect 5867 576 6433 584
rect 6447 576 6493 584
rect 7407 576 8113 584
rect 8127 576 8213 584
rect 8227 576 8233 584
rect 8247 576 8893 584
rect 8907 576 9233 584
rect 9567 576 9653 584
rect 9827 576 10453 584
rect 11307 576 11353 584
rect 11387 576 11453 584
rect 11527 576 11633 584
rect 187 556 373 564
rect 387 556 393 564
rect 1727 556 1753 564
rect 2847 556 6133 564
rect 7747 556 7793 564
rect 7807 556 7973 564
rect 7987 556 8713 564
rect 8887 556 8933 564
rect 9867 556 10173 564
rect 3887 536 3953 544
rect 6487 536 7733 544
rect 8287 536 8493 544
rect 9087 536 9513 544
rect 3567 516 5453 524
rect 8547 516 8673 524
rect 8687 516 9093 524
rect 9207 516 10013 524
rect 3207 496 3953 504
rect 4087 496 4193 504
rect 7667 496 8813 504
rect 8827 496 9253 504
rect 7827 476 8853 484
rect 3867 456 4113 464
rect 6747 456 7413 464
rect 7427 456 7673 464
rect 8047 456 9433 464
rect 3687 436 4093 444
rect 7667 436 8333 444
rect 8627 436 10553 444
rect 10727 436 11033 444
rect 1567 416 2433 424
rect 2447 416 2593 424
rect 2967 416 3153 424
rect 3167 416 4413 424
rect 4927 416 5733 424
rect 6547 416 7893 424
rect 8407 416 8893 424
rect 10387 416 11113 424
rect 527 396 1153 404
rect 2147 396 2653 404
rect 2667 396 2913 404
rect 2947 396 3993 404
rect 4187 396 4253 404
rect 4267 396 4893 404
rect 4907 396 5013 404
rect 5027 396 5513 404
rect 6027 396 7053 404
rect 7487 396 7613 404
rect 7687 396 8113 404
rect 8507 396 8533 404
rect 9887 396 10113 404
rect 10687 396 11093 404
rect 11167 396 11293 404
rect 11307 396 12013 404
rect 167 376 273 384
rect 647 376 853 384
rect 1827 376 1873 384
rect 2427 376 2753 384
rect 2807 376 2993 384
rect 3007 376 3193 384
rect 3407 376 3533 384
rect 3987 376 4273 384
rect 4407 376 4853 384
rect 5487 376 5573 384
rect 5947 376 6013 384
rect 6767 376 6853 384
rect 7307 376 7653 384
rect 7676 376 7833 384
rect -24 356 93 364
rect 147 356 253 364
rect 567 356 893 364
rect 1407 356 1553 364
rect 1727 356 1853 364
rect 2247 356 2373 364
rect 2387 356 2393 364
rect 2827 356 2933 364
rect 3247 356 3373 364
rect 3447 356 3573 364
rect 3847 356 3913 364
rect 3936 356 4013 364
rect 787 336 873 344
rect 996 344 1004 353
rect 3936 347 3944 356
rect 4107 356 4133 364
rect 4267 356 4333 364
rect 4536 356 4724 364
rect 4536 347 4544 356
rect 996 336 1133 344
rect 1207 336 1373 344
rect 1427 336 1433 344
rect 1447 336 1533 344
rect 1587 336 1613 344
rect 2527 336 2613 344
rect 3427 336 3753 344
rect 3867 336 3893 344
rect 4007 336 4393 344
rect 4647 336 4693 344
rect 4716 344 4724 356
rect 4867 356 5033 364
rect 5227 356 5373 364
rect 5607 356 5773 364
rect 5827 356 5973 364
rect 6787 356 6833 364
rect 6896 364 6904 373
rect 6896 356 7073 364
rect 7676 364 7684 376
rect 8007 376 8293 384
rect 8427 376 8653 384
rect 8747 376 9033 384
rect 9747 376 9893 384
rect 10287 376 10373 384
rect 10547 376 10853 384
rect 11267 376 11433 384
rect 11447 376 11644 384
rect 11636 367 11644 376
rect 11727 376 11833 384
rect 11847 376 12053 384
rect 7127 356 7684 364
rect 7727 356 8073 364
rect 8327 356 8493 364
rect 8607 356 9053 364
rect 9067 356 9153 364
rect 9267 356 9453 364
rect 9587 356 9673 364
rect 9787 356 9833 364
rect 10007 356 10053 364
rect 10127 356 10253 364
rect 10427 356 10564 364
rect 4716 336 4733 344
rect 4747 336 4913 344
rect 4967 336 5033 344
rect 5287 336 5393 344
rect 5416 344 5424 353
rect 5416 336 5633 344
rect 5967 336 5993 344
rect 6267 336 6433 344
rect 6487 336 6533 344
rect 6567 336 7113 344
rect 7507 336 7533 344
rect 7827 336 7853 344
rect 7927 336 8093 344
rect 8487 336 8633 344
rect 8707 336 8733 344
rect 8927 336 9073 344
rect 9127 336 9653 344
rect 10016 336 10433 344
rect 10016 327 10024 336
rect 10487 336 10533 344
rect 10556 344 10564 356
rect 10587 356 10633 364
rect 11007 356 11033 364
rect 11087 356 11113 364
rect 11147 356 11213 364
rect 11227 356 11473 364
rect 11687 356 12033 364
rect 10556 336 10653 344
rect 10707 336 10793 344
rect 10827 336 11013 344
rect 11067 336 11093 344
rect 11587 336 11633 344
rect 11647 336 11653 344
rect 11807 336 11853 344
rect 11967 336 12033 344
rect 12047 336 12073 344
rect 1007 316 1353 324
rect 1547 316 2453 324
rect 2467 316 2573 324
rect 2647 316 3013 324
rect 3027 316 3173 324
rect 3227 316 3833 324
rect 3987 316 4024 324
rect 727 296 1173 304
rect 2167 296 2413 304
rect 3487 296 3993 304
rect 4016 304 4024 316
rect 4327 316 4513 324
rect 4727 316 4933 324
rect 4947 316 5073 324
rect 5967 316 6013 324
rect 6187 316 6673 324
rect 6887 316 7233 324
rect 7627 316 7653 324
rect 7747 316 9213 324
rect 10047 316 10473 324
rect 10627 316 10993 324
rect 11287 316 11373 324
rect 4016 296 6273 304
rect 6727 296 7013 304
rect 7056 296 7313 304
rect 967 276 1073 284
rect 1367 276 2973 284
rect 4227 276 4513 284
rect 7056 284 7064 296
rect 7327 296 7633 304
rect 8147 296 8873 304
rect 9907 296 11233 304
rect 6927 276 7064 284
rect 7087 276 8413 284
rect 8867 276 9853 284
rect 10087 276 10133 284
rect 10987 276 11053 284
rect 607 256 673 264
rect 2567 256 2613 264
rect 2807 256 5913 264
rect 7107 256 7453 264
rect 8127 256 8673 264
rect 9027 256 9873 264
rect 9887 256 10213 264
rect 507 236 813 244
rect 1607 236 2833 244
rect 2867 236 2893 244
rect 7267 236 8973 244
rect 9707 236 11813 244
rect 11827 236 11833 244
rect 1747 216 2073 224
rect 2087 216 2333 224
rect 2607 216 2673 224
rect 3807 216 3833 224
rect 5467 216 5693 224
rect 6987 216 8253 224
rect 9367 216 9473 224
rect 9567 216 10473 224
rect 10487 216 10873 224
rect 10887 216 10913 224
rect 1987 196 2133 204
rect 3147 196 3173 204
rect 4427 196 4873 204
rect 4887 196 5873 204
rect 6307 196 9904 204
rect 387 176 473 184
rect 1207 176 1633 184
rect 1807 176 1833 184
rect 1967 176 1993 184
rect 2507 176 2733 184
rect 3447 176 3473 184
rect 3547 176 3713 184
rect 3727 176 3953 184
rect 3967 176 4373 184
rect 4387 176 4693 184
rect 5147 176 5153 184
rect 5167 176 5333 184
rect 5587 176 5913 184
rect 6587 176 7073 184
rect 7147 176 7613 184
rect 7707 176 7913 184
rect 8087 176 8233 184
rect 8407 176 8433 184
rect 8787 176 8933 184
rect 9227 176 9513 184
rect 9896 184 9904 196
rect 9927 196 10613 204
rect 11227 196 11473 204
rect 11507 196 11793 204
rect 9896 176 10073 184
rect 10407 176 10433 184
rect 10527 176 10653 184
rect 10827 176 11273 184
rect 11347 176 11813 184
rect -24 156 133 164
rect -24 116 -16 156
rect 296 156 433 164
rect 296 147 304 156
rect 1687 156 1824 164
rect 1816 147 1824 156
rect 1956 156 2093 164
rect 1956 147 1964 156
rect 2316 156 2453 164
rect 2316 147 2324 156
rect 3327 156 3344 164
rect 467 136 513 144
rect 907 136 1373 144
rect 1467 136 1593 144
rect 1667 136 1733 144
rect 2087 136 2113 144
rect 2347 136 2473 144
rect 2727 136 3313 144
rect 247 116 553 124
rect 567 116 1033 124
rect 1887 116 2573 124
rect 3167 116 3293 124
rect 3336 107 3344 156
rect 4447 156 4473 164
rect 4627 156 4653 164
rect 5307 156 5533 164
rect 6116 164 6124 173
rect 5747 156 5904 164
rect 6116 156 6173 164
rect 5896 147 5904 156
rect 7067 156 7233 164
rect 7667 156 7813 164
rect 8307 156 9393 164
rect 9716 164 9724 173
rect 9407 156 9724 164
rect 10127 156 10873 164
rect 11247 156 11333 164
rect 11456 156 11624 164
rect 3367 136 3493 144
rect 3607 136 3653 144
rect 4167 136 4653 144
rect 5367 136 5493 144
rect 5647 136 5713 144
rect 7047 136 7133 144
rect 7167 136 7213 144
rect 7487 136 7533 144
rect 7627 136 7673 144
rect 7836 144 7844 153
rect 7687 136 7844 144
rect 7927 136 8633 144
rect 8647 136 8833 144
rect 8967 136 9013 144
rect 9347 136 9573 144
rect 10007 136 10053 144
rect 10107 136 10133 144
rect 10467 136 10533 144
rect 10567 136 10633 144
rect 10687 136 10813 144
rect 11076 144 11084 153
rect 11456 147 11464 156
rect 10907 136 11084 144
rect 11107 136 11213 144
rect 11307 136 11453 144
rect 11476 136 11493 144
rect 3367 116 3533 124
rect 4027 116 4133 124
rect 4647 116 4833 124
rect 5787 116 6113 124
rect 7807 116 7853 124
rect 7887 116 8053 124
rect 8287 116 8393 124
rect 9307 116 9373 124
rect 10307 116 11133 124
rect 11476 124 11484 136
rect 11616 144 11624 156
rect 11867 156 12033 164
rect 11616 136 11653 144
rect 11267 116 11484 124
rect 7527 96 8013 104
rect 267 16 293 24
rect 967 16 993 24
rect 2127 16 2253 24
rect 2287 16 2313 24
rect 2827 16 2893 24
rect 3467 16 3493 24
rect 3787 16 3813 24
rect 4107 16 4133 24
rect 4687 16 4753 24
rect 4807 16 4833 24
rect 6127 16 6153 24
use BUFX2  _2478_
timestamp 0
transform -1 0 190 0 1 3610
box -6 -8 86 248
use BUFX2  _2479_
timestamp 0
transform -1 0 190 0 1 2650
box -6 -8 86 248
use BUFX2  _2480_
timestamp 0
transform 1 0 1970 0 -1 730
box -6 -8 86 248
use BUFX2  _2481_
timestamp 0
transform 1 0 2790 0 -1 2170
box -6 -8 86 248
use BUFX2  _2482_
timestamp 0
transform -1 0 190 0 -1 5050
box -6 -8 86 248
use BUFX2  _2483_
timestamp 0
transform -1 0 670 0 -1 5530
box -6 -8 86 248
use BUFX2  _2484_
timestamp 0
transform -1 0 2230 0 -1 730
box -6 -8 86 248
use BUFX2  _2485_
timestamp 0
transform 1 0 3990 0 -1 1690
box -6 -8 86 248
use BUFX2  _2486_
timestamp 0
transform 1 0 12110 0 1 2650
box -6 -8 86 248
use BUFX2  _2487_
timestamp 0
transform -1 0 6750 0 -1 250
box -6 -8 86 248
use BUFX2  _2488_
timestamp 0
transform -1 0 6910 0 -1 250
box -6 -8 86 248
use BUFX2  _2489_
timestamp 0
transform 1 0 12070 0 -1 3130
box -6 -8 86 248
use BUFX2  _2490_
timestamp 0
transform 1 0 12070 0 1 3130
box -6 -8 86 248
use BUFX2  _2491_
timestamp 0
transform 1 0 6490 0 -1 250
box -6 -8 86 248
use BUFX2  _2492_
timestamp 0
transform 1 0 11890 0 1 3130
box -6 -8 86 248
use BUFX2  _2493_
timestamp 0
transform -1 0 12050 0 -1 250
box -6 -8 86 248
use BUFX2  _2494_
timestamp 0
transform -1 0 1150 0 1 6010
box -6 -8 86 248
use BUFX2  _2495_
timestamp 0
transform -1 0 1310 0 1 2170
box -6 -8 86 248
use BUFX2  _2496_
timestamp 0
transform -1 0 190 0 1 4090
box -6 -8 86 248
use BUFX2  _2497_
timestamp 0
transform -1 0 4530 0 -1 250
box -6 -8 86 248
use BUFX2  _2498_
timestamp 0
transform 1 0 4510 0 -1 3610
box -6 -8 86 248
use BUFX2  _2499_
timestamp 0
transform -1 0 3390 0 -1 730
box -6 -8 86 248
use BUFX2  _2500_
timestamp 0
transform -1 0 570 0 -1 3130
box -6 -8 86 248
use BUFX2  _2501_
timestamp 0
transform -1 0 3770 0 1 2170
box -6 -8 86 248
use BUFX2  _2502_
timestamp 0
transform -1 0 190 0 -1 6490
box -6 -8 86 248
use BUFX2  _2503_
timestamp 0
transform -1 0 190 0 -1 250
box -6 -8 86 248
use BUFX2  _2504_
timestamp 0
transform 1 0 4610 0 -1 2170
box -6 -8 86 248
use BUFX2  _2505_
timestamp 0
transform 1 0 5150 0 -1 250
box -6 -8 86 248
use BUFX2  _2506_
timestamp 0
transform -1 0 2650 0 -1 1690
box -6 -8 86 248
use BUFX2  _2507_
timestamp 0
transform 1 0 3870 0 1 1210
box -6 -8 86 248
use BUFX2  _2508_
timestamp 0
transform 1 0 3470 0 1 1210
box -6 -8 86 248
use BUFX2  _2509_
timestamp 0
transform 1 0 4270 0 -1 250
box -6 -8 86 248
use BUFX2  _2510_
timestamp 0
transform 1 0 3130 0 -1 730
box -6 -8 86 248
use BUFX2  _2511_
timestamp 0
transform -1 0 5050 0 -1 250
box -6 -8 86 248
use DFFPOSX1  _2512_
timestamp 0
transform -1 0 6390 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _2513_
timestamp 0
transform -1 0 5710 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _2514_
timestamp 0
transform -1 0 4450 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _2515_
timestamp 0
transform -1 0 5890 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _2516_
timestamp 0
transform -1 0 6570 0 1 250
box -6 -8 246 248
use DFFPOSX1  _2517_
timestamp 0
transform -1 0 5410 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _2518_
timestamp 0
transform 1 0 5090 0 -1 2170
box -6 -8 246 248
use OAI21X1  _2519_
timestamp 0
transform -1 0 5810 0 1 2170
box -6 -8 106 248
use NAND3X1  _2520_
timestamp 0
transform -1 0 7670 0 1 3130
box -6 -8 106 248
use NAND3X1  _2521_
timestamp 0
transform -1 0 7870 0 1 3130
box -6 -8 106 248
use OAI22X1  _2522_
timestamp 0
transform 1 0 7790 0 -1 3130
box -6 -8 126 248
use NOR2X1  _2523_
timestamp 0
transform 1 0 9530 0 -1 3130
box -6 -8 86 248
use AOI21X1  _2524_
timestamp 0
transform -1 0 7930 0 -1 2650
box -6 -8 106 248
use OAI21X1  _2525_
timestamp 0
transform 1 0 7590 0 -1 3130
box -6 -8 106 248
use OAI21X1  _2526_
timestamp 0
transform 1 0 8330 0 1 3610
box -6 -8 106 248
use AOI22X1  _2527_
timestamp 0
transform 1 0 8530 0 1 3610
box -6 -8 126 248
use AND2X2  _2528_
timestamp 0
transform -1 0 9750 0 1 3610
box -6 -8 106 248
use OAI21X1  _2529_
timestamp 0
transform 1 0 8610 0 -1 3610
box -6 -8 106 248
use NOR2X1  _2530_
timestamp 0
transform -1 0 8310 0 -1 3610
box -6 -8 86 248
use OAI21X1  _2531_
timestamp 0
transform -1 0 8470 0 1 3130
box -6 -8 106 248
use AOI21X1  _2532_
timestamp 0
transform -1 0 8890 0 1 3130
box -6 -8 106 248
use OAI21X1  _2533_
timestamp 0
transform 1 0 9550 0 -1 4090
box -6 -8 106 248
use OAI21X1  _2534_
timestamp 0
transform 1 0 10110 0 1 4090
box -6 -8 106 248
use AOI21X1  _2535_
timestamp 0
transform -1 0 10370 0 -1 3130
box -6 -8 106 248
use OAI21X1  _2536_
timestamp 0
transform -1 0 8890 0 -1 3130
box -6 -8 106 248
use AOI21X1  _2537_
timestamp 0
transform -1 0 8690 0 -1 3130
box -6 -8 106 248
use OAI21X1  _2538_
timestamp 0
transform -1 0 8490 0 -1 3130
box -6 -8 106 248
use AOI21X1  _2539_
timestamp 0
transform 1 0 8010 0 -1 3130
box -6 -8 106 248
use OAI21X1  _2540_
timestamp 0
transform -1 0 10790 0 -1 3130
box -6 -8 106 248
use NAND3X1  _2541_
timestamp 0
transform -1 0 10990 0 -1 3130
box -6 -8 106 248
use NAND2X1  _2542_
timestamp 0
transform 1 0 10950 0 1 3130
box -6 -8 86 248
use OAI21X1  _2543_
timestamp 0
transform -1 0 10730 0 1 3610
box -6 -8 106 248
use OAI21X1  _2544_
timestamp 0
transform -1 0 5830 0 -1 2650
box -6 -8 106 248
use OAI22X1  _2545_
timestamp 0
transform -1 0 6050 0 -1 2650
box -6 -8 126 248
use OAI21X1  _2546_
timestamp 0
transform -1 0 6250 0 -1 2650
box -6 -8 106 248
use OAI21X1  _2547_
timestamp 0
transform -1 0 6130 0 -1 2170
box -6 -8 106 248
use NAND3X1  _2548_
timestamp 0
transform -1 0 6330 0 -1 2170
box -6 -8 106 248
use NAND3X1  _2549_
timestamp 0
transform 1 0 5630 0 -1 2170
box -6 -8 106 248
use AND2X2  _2550_
timestamp 0
transform 1 0 5830 0 -1 2170
box -6 -8 106 248
use AOI21X1  _2551_
timestamp 0
transform -1 0 7030 0 -1 2650
box -6 -8 106 248
use OAI21X1  _2552_
timestamp 0
transform -1 0 7390 0 1 2650
box -6 -8 106 248
use AOI21X1  _2553_
timestamp 0
transform -1 0 5850 0 1 1690
box -6 -8 106 248
use OAI21X1  _2554_
timestamp 0
transform -1 0 6490 0 1 1210
box -6 -8 106 248
use AOI21X1  _2555_
timestamp 0
transform 1 0 6430 0 -1 1210
box -6 -8 106 248
use OAI21X1  _2556_
timestamp 0
transform -1 0 6870 0 1 730
box -6 -8 106 248
use OAI21X1  _2557_
timestamp 0
transform -1 0 6350 0 -1 1210
box -6 -8 106 248
use NOR2X1  _2558_
timestamp 0
transform 1 0 6550 0 1 1690
box -6 -8 86 248
use OAI21X1  _2559_
timestamp 0
transform 1 0 6930 0 1 1690
box -6 -8 106 248
use OAI21X1  _2560_
timestamp 0
transform -1 0 6050 0 1 1690
box -6 -8 106 248
use AOI21X1  _2561_
timestamp 0
transform -1 0 6690 0 1 1210
box -6 -8 106 248
use NOR2X1  _2562_
timestamp 0
transform 1 0 6790 0 1 1210
box -6 -8 86 248
use AOI21X1  _2563_
timestamp 0
transform -1 0 6250 0 1 1690
box -6 -8 106 248
use MUX2X1  _2564_
timestamp 0
transform 1 0 7830 0 1 250
box -6 -8 126 248
use AOI22X1  _2565_
timestamp 0
transform 1 0 8050 0 1 250
box -6 -8 126 248
use AOI21X1  _2566_
timestamp 0
transform 1 0 7630 0 1 250
box -6 -8 106 248
use OAI22X1  _2567_
timestamp 0
transform 1 0 7030 0 -1 1690
box -6 -8 126 248
use OAI21X1  _2568_
timestamp 0
transform -1 0 6750 0 -1 1690
box -6 -8 106 248
use NOR2X1  _2569_
timestamp 0
transform 1 0 7250 0 -1 1690
box -6 -8 86 248
use NAND3X1  _2570_
timestamp 0
transform -1 0 9510 0 1 250
box -6 -8 106 248
use OAI21X1  _2571_
timestamp 0
transform -1 0 9410 0 -1 250
box -6 -8 106 248
use NOR2X1  _2572_
timestamp 0
transform 1 0 9350 0 -1 1690
box -6 -8 86 248
use NAND2X1  _2573_
timestamp 0
transform 1 0 9230 0 1 250
box -6 -8 86 248
use OAI21X1  _2574_
timestamp 0
transform -1 0 9390 0 -1 730
box -6 -8 106 248
use OAI21X1  _2575_
timestamp 0
transform -1 0 9190 0 -1 730
box -6 -8 106 248
use OAI21X1  _2576_
timestamp 0
transform -1 0 8930 0 1 250
box -6 -8 106 248
use OAI21X1  _2577_
timestamp 0
transform -1 0 9130 0 1 250
box -6 -8 106 248
use OAI21X1  _2578_
timestamp 0
transform 1 0 9610 0 1 250
box -6 -8 106 248
use OAI21X1  _2579_
timestamp 0
transform -1 0 9630 0 1 1210
box -6 -8 106 248
use AOI21X1  _2580_
timestamp 0
transform -1 0 8430 0 1 730
box -6 -8 106 248
use OAI21X1  _2581_
timestamp 0
transform 1 0 8310 0 -1 730
box -6 -8 106 248
use INVX1  _2582_
timestamp 0
transform 1 0 8430 0 -1 1210
box -6 -8 66 248
use OAI21X1  _2583_
timestamp 0
transform -1 0 9910 0 1 250
box -6 -8 106 248
use AOI21X1  _2584_
timestamp 0
transform 1 0 9490 0 -1 730
box -6 -8 106 248
use AOI21X1  _2585_
timestamp 0
transform -1 0 11310 0 1 250
box -6 -8 106 248
use AOI22X1  _2586_
timestamp 0
transform 1 0 8910 0 1 1210
box -6 -8 126 248
use AOI21X1  _2587_
timestamp 0
transform 1 0 8710 0 1 1690
box -6 -8 106 248
use OAI21X1  _2588_
timestamp 0
transform -1 0 8610 0 1 1690
box -6 -8 106 248
use OAI21X1  _2589_
timestamp 0
transform 1 0 8570 0 -1 1690
box -6 -8 106 248
use OAI21X1  _2590_
timestamp 0
transform 1 0 8310 0 1 1690
box -6 -8 106 248
use AOI21X1  _2591_
timestamp 0
transform -1 0 8730 0 -1 2170
box -6 -8 106 248
use OAI21X1  _2592_
timestamp 0
transform 1 0 7910 0 1 1690
box -6 -8 106 248
use NAND3X1  _2593_
timestamp 0
transform -1 0 9230 0 1 1210
box -6 -8 106 248
use AOI22X1  _2594_
timestamp 0
transform -1 0 9150 0 -1 2170
box -6 -8 126 248
use INVX1  _2595_
timestamp 0
transform -1 0 9330 0 1 1690
box -6 -8 66 248
use NAND2X1  _2596_
timestamp 0
transform 1 0 10490 0 1 1210
box -6 -8 86 248
use OAI21X1  _2597_
timestamp 0
transform 1 0 10670 0 1 1210
box -6 -8 106 248
use AOI21X1  _2598_
timestamp 0
transform -1 0 10590 0 -1 730
box -6 -8 106 248
use OAI21X1  _2599_
timestamp 0
transform 1 0 10870 0 -1 730
box -6 -8 106 248
use OAI21X1  _2600_
timestamp 0
transform -1 0 11550 0 -1 730
box -6 -8 106 248
use OAI21X1  _2601_
timestamp 0
transform 1 0 8330 0 1 1210
box -6 -8 106 248
use AOI21X1  _2602_
timestamp 0
transform -1 0 8210 0 1 1690
box -6 -8 106 248
use NAND3X1  _2603_
timestamp 0
transform 1 0 7130 0 1 1690
box -6 -8 106 248
use OAI21X1  _2604_
timestamp 0
transform 1 0 8290 0 1 2170
box -6 -8 106 248
use NOR2X1  _2605_
timestamp 0
transform -1 0 8230 0 1 730
box -6 -8 86 248
use OAI22X1  _2606_
timestamp 0
transform -1 0 7870 0 1 730
box -6 -8 126 248
use OAI21X1  _2607_
timestamp 0
transform -1 0 6710 0 1 3130
box -6 -8 106 248
use NAND3X1  _2608_
timestamp 0
transform 1 0 6810 0 1 3130
box -6 -8 106 248
use OAI21X1  _2609_
timestamp 0
transform 1 0 7010 0 1 3130
box -6 -8 106 248
use AOI21X1  _2610_
timestamp 0
transform -1 0 8030 0 1 3610
box -6 -8 106 248
use NAND3X1  _2611_
timestamp 0
transform -1 0 10250 0 -1 4090
box -6 -8 106 248
use NAND3X1  _2612_
timestamp 0
transform 1 0 9950 0 -1 4090
box -6 -8 106 248
use NAND3X1  _2613_
timestamp 0
transform 1 0 10350 0 -1 4090
box -6 -8 106 248
use NAND3X1  _2614_
timestamp 0
transform -1 0 11130 0 1 4090
box -6 -8 106 248
use OAI21X1  _2615_
timestamp 0
transform -1 0 7290 0 1 3130
box -6 -8 106 248
use OAI21X1  _2616_
timestamp 0
transform 1 0 8370 0 -1 1690
box -6 -8 106 248
use NOR2X1  _2617_
timestamp 0
transform -1 0 7290 0 -1 3130
box -6 -8 86 248
use AOI21X1  _2618_
timestamp 0
transform -1 0 6650 0 -1 2650
box -6 -8 106 248
use OAI21X1  _2619_
timestamp 0
transform 1 0 6350 0 -1 2650
box -6 -8 106 248
use NAND3X1  _2620_
timestamp 0
transform -1 0 8130 0 -1 3610
box -6 -8 106 248
use NAND3X1  _2621_
timestamp 0
transform -1 0 8230 0 1 3610
box -6 -8 106 248
use OAI21X1  _2622_
timestamp 0
transform 1 0 8410 0 -1 3610
box -6 -8 106 248
use AOI21X1  _2623_
timestamp 0
transform -1 0 9090 0 -1 3610
box -6 -8 106 248
use OAI21X1  _2624_
timestamp 0
transform 1 0 8150 0 -1 4090
box -6 -8 106 248
use OAI21X1  _2625_
timestamp 0
transform 1 0 6910 0 1 2650
box -6 -8 106 248
use INVX1  _2626_
timestamp 0
transform -1 0 8410 0 -1 4090
box -6 -8 66 248
use OAI21X1  _2627_
timestamp 0
transform 1 0 9970 0 -1 3610
box -6 -8 106 248
use OAI22X1  _2628_
timestamp 0
transform 1 0 11590 0 -1 3610
box -6 -8 126 248
use NAND3X1  _2629_
timestamp 0
transform 1 0 11490 0 -1 3130
box -6 -8 106 248
use NOR2X1  _2630_
timestamp 0
transform 1 0 11770 0 1 3610
box -6 -8 86 248
use OAI21X1  _2631_
timestamp 0
transform -1 0 11670 0 1 3610
box -6 -8 106 248
use AOI21X1  _2632_
timestamp 0
transform 1 0 9490 0 1 2650
box -6 -8 106 248
use MUX2X1  _2633_
timestamp 0
transform -1 0 8690 0 1 3130
box -6 -8 126 248
use AOI22X1  _2634_
timestamp 0
transform 1 0 8990 0 1 3130
box -6 -8 126 248
use AOI21X1  _2635_
timestamp 0
transform -1 0 9290 0 1 3130
box -6 -8 106 248
use AOI21X1  _2636_
timestamp 0
transform -1 0 10090 0 1 3130
box -6 -8 106 248
use OAI21X1  _2637_
timestamp 0
transform -1 0 8790 0 1 2650
box -6 -8 106 248
use NAND2X1  _2638_
timestamp 0
transform 1 0 9790 0 -1 3610
box -6 -8 86 248
use OAI21X1  _2639_
timestamp 0
transform 1 0 10050 0 1 3610
box -6 -8 106 248
use AOI21X1  _2640_
timestamp 0
transform 1 0 8170 0 1 3130
box -6 -8 106 248
use OAI21X1  _2641_
timestamp 0
transform 1 0 7970 0 1 3130
box -6 -8 106 248
use NAND3X1  _2642_
timestamp 0
transform 1 0 9450 0 1 2170
box -6 -8 106 248
use OAI21X1  _2643_
timestamp 0
transform 1 0 9450 0 -1 2170
box -6 -8 106 248
use AOI22X1  _2644_
timestamp 0
transform 1 0 8470 0 1 2650
box -6 -8 126 248
use AOI21X1  _2645_
timestamp 0
transform 1 0 7690 0 1 2650
box -6 -8 106 248
use OAI21X1  _2646_
timestamp 0
transform 1 0 7490 0 1 2650
box -6 -8 106 248
use OAI21X1  _2647_
timestamp 0
transform 1 0 8270 0 1 2650
box -6 -8 106 248
use NOR2X1  _2648_
timestamp 0
transform -1 0 8170 0 1 2650
box -6 -8 86 248
use AOI21X1  _2649_
timestamp 0
transform -1 0 9190 0 1 2650
box -6 -8 106 248
use NOR2X1  _2650_
timestamp 0
transform 1 0 11170 0 1 2650
box -6 -8 86 248
use OAI21X1  _2651_
timestamp 0
transform -1 0 9390 0 1 2650
box -6 -8 106 248
use OAI21X1  _2652_
timestamp 0
transform -1 0 8690 0 -1 2650
box -6 -8 106 248
use NOR2X1  _2653_
timestamp 0
transform 1 0 8790 0 -1 2650
box -6 -8 86 248
use OAI21X1  _2654_
timestamp 0
transform 1 0 5910 0 1 2170
box -6 -8 106 248
use NAND3X1  _2655_
timestamp 0
transform -1 0 6190 0 1 2170
box -6 -8 106 248
use NAND3X1  _2656_
timestamp 0
transform -1 0 6390 0 1 2170
box -6 -8 106 248
use NAND3X1  _2657_
timestamp 0
transform -1 0 7790 0 1 2170
box -6 -8 106 248
use AOI22X1  _2658_
timestamp 0
transform 1 0 7470 0 1 2170
box -6 -8 126 248
use NOR2X1  _2659_
timestamp 0
transform -1 0 7290 0 -1 2170
box -6 -8 86 248
use NOR2X1  _2660_
timestamp 0
transform -1 0 7470 0 1 3130
box -6 -8 86 248
use NAND3X1  _2661_
timestamp 0
transform -1 0 10930 0 1 1690
box -6 -8 106 248
use NAND2X1  _2662_
timestamp 0
transform 1 0 11030 0 1 1690
box -6 -8 86 248
use NAND2X1  _2663_
timestamp 0
transform 1 0 10090 0 -1 1690
box -6 -8 86 248
use INVX1  _2664_
timestamp 0
transform 1 0 10270 0 -1 1690
box -6 -8 66 248
use OAI21X1  _2665_
timestamp 0
transform -1 0 6770 0 1 2170
box -6 -8 106 248
use AOI21X1  _2666_
timestamp 0
transform 1 0 7270 0 1 2170
box -6 -8 106 248
use AOI22X1  _2667_
timestamp 0
transform -1 0 7170 0 1 2170
box -6 -8 126 248
use NOR2X1  _2668_
timestamp 0
transform -1 0 6950 0 1 2170
box -6 -8 86 248
use OAI21X1  _2669_
timestamp 0
transform 1 0 6810 0 -1 2170
box -6 -8 106 248
use OAI21X1  _2670_
timestamp 0
transform -1 0 10750 0 1 2170
box -6 -8 106 248
use AOI21X1  _2671_
timestamp 0
transform 1 0 11730 0 -1 2170
box -6 -8 106 248
use OAI21X1  _2672_
timestamp 0
transform 1 0 11770 0 1 1690
box -6 -8 106 248
use NAND2X1  _2673_
timestamp 0
transform -1 0 11630 0 -1 1690
box -6 -8 86 248
use OAI22X1  _2674_
timestamp 0
transform 1 0 11510 0 -1 2170
box -6 -8 126 248
use AOI21X1  _2675_
timestamp 0
transform -1 0 10930 0 1 2170
box -6 -8 106 248
use OAI21X1  _2676_
timestamp 0
transform 1 0 11490 0 -1 2650
box -6 -8 106 248
use NOR2X1  _2677_
timestamp 0
transform -1 0 11630 0 1 2650
box -6 -8 86 248
use AOI22X1  _2678_
timestamp 0
transform -1 0 10290 0 -1 3610
box -6 -8 126 248
use AOI21X1  _2679_
timestamp 0
transform 1 0 9790 0 1 3130
box -6 -8 106 248
use AOI21X1  _2680_
timestamp 0
transform 1 0 9710 0 -1 3130
box -6 -8 106 248
use AOI21X1  _2681_
timestamp 0
transform 1 0 9390 0 1 3130
box -6 -8 106 248
use OAI21X1  _2682_
timestamp 0
transform -1 0 9690 0 1 3130
box -6 -8 106 248
use NAND3X1  _2683_
timestamp 0
transform -1 0 10350 0 1 3610
box -6 -8 106 248
use OAI21X1  _2684_
timestamp 0
transform -1 0 10650 0 -1 4090
box -6 -8 106 248
use AOI21X1  _2685_
timestamp 0
transform -1 0 10930 0 1 4090
box -6 -8 106 248
use NOR2X1  _2686_
timestamp 0
transform 1 0 10750 0 -1 4090
box -6 -8 86 248
use OAI21X1  _2687_
timestamp 0
transform -1 0 9950 0 1 3610
box -6 -8 106 248
use AOI21X1  _2688_
timestamp 0
transform 1 0 9270 0 1 3610
box -6 -8 106 248
use AOI22X1  _2689_
timestamp 0
transform 1 0 10590 0 -1 3610
box -6 -8 126 248
use AOI21X1  _2690_
timestamp 0
transform -1 0 11030 0 -1 4090
box -6 -8 106 248
use OAI21X1  _2691_
timestamp 0
transform -1 0 11230 0 -1 4090
box -6 -8 106 248
use OAI21X1  _2692_
timestamp 0
transform 1 0 11330 0 -1 4090
box -6 -8 106 248
use AOI22X1  _2693_
timestamp 0
transform -1 0 10590 0 -1 3130
box -6 -8 126 248
use NOR2X1  _2694_
timestamp 0
transform 1 0 9690 0 1 2650
box -6 -8 86 248
use OAI21X1  _2695_
timestamp 0
transform -1 0 10670 0 -1 2170
box -6 -8 106 248
use NAND2X1  _2696_
timestamp 0
transform 1 0 10370 0 1 3130
box -6 -8 86 248
use AOI22X1  _2697_
timestamp 0
transform 1 0 10030 0 -1 250
box -6 -8 126 248
use AOI21X1  _2698_
timestamp 0
transform 1 0 10010 0 1 250
box -6 -8 106 248
use OAI21X1  _2699_
timestamp 0
transform 1 0 9130 0 1 730
box -6 -8 106 248
use OAI22X1  _2700_
timestamp 0
transform 1 0 8910 0 1 730
box -6 -8 126 248
use OAI21X1  _2701_
timestamp 0
transform -1 0 8630 0 1 730
box -6 -8 106 248
use OAI21X1  _2702_
timestamp 0
transform 1 0 8910 0 -1 730
box -6 -8 106 248
use OAI21X1  _2703_
timestamp 0
transform 1 0 10930 0 1 730
box -6 -8 106 248
use NAND3X1  _2704_
timestamp 0
transform -1 0 9270 0 -1 1210
box -6 -8 106 248
use NAND3X1  _2705_
timestamp 0
transform -1 0 9830 0 -1 1210
box -6 -8 106 248
use OAI21X1  _2706_
timestamp 0
transform -1 0 10230 0 -1 1210
box -6 -8 106 248
use OAI21X1  _2707_
timestamp 0
transform -1 0 9750 0 -1 2170
box -6 -8 106 248
use OAI21X1  _2708_
timestamp 0
transform 1 0 8970 0 -1 1210
box -6 -8 106 248
use AOI21X1  _2709_
timestamp 0
transform 1 0 9090 0 1 1690
box -6 -8 106 248
use OAI21X1  _2710_
timestamp 0
transform -1 0 8870 0 -1 1210
box -6 -8 106 248
use OAI21X1  _2711_
timestamp 0
transform -1 0 10930 0 -1 250
box -6 -8 106 248
use AOI21X1  _2712_
timestamp 0
transform -1 0 10910 0 1 250
box -6 -8 106 248
use AOI22X1  _2713_
timestamp 0
transform 1 0 10870 0 1 1210
box -6 -8 126 248
use OAI21X1  _2714_
timestamp 0
transform 1 0 10870 0 -1 1210
box -6 -8 106 248
use AOI21X1  _2715_
timestamp 0
transform -1 0 11570 0 1 1210
box -6 -8 106 248
use NOR2X1  _2716_
timestamp 0
transform 1 0 11670 0 1 1210
box -6 -8 86 248
use INVX1  _2717_
timestamp 0
transform -1 0 10830 0 -1 2170
box -6 -8 66 248
use OAI21X1  _2718_
timestamp 0
transform 1 0 11130 0 -1 2170
box -6 -8 106 248
use NAND3X1  _2719_
timestamp 0
transform 1 0 11850 0 1 1210
box -6 -8 106 248
use OAI21X1  _2720_
timestamp 0
transform -1 0 11130 0 -1 250
box -6 -8 106 248
use OAI21X1  _2721_
timestamp 0
transform -1 0 11030 0 -1 2170
box -6 -8 106 248
use AOI21X1  _2722_
timestamp 0
transform -1 0 11070 0 1 2650
box -6 -8 106 248
use OAI21X1  _2723_
timestamp 0
transform 1 0 11430 0 -1 250
box -6 -8 106 248
use OAI21X1  _2724_
timestamp 0
transform 1 0 11410 0 1 250
box -6 -8 106 248
use AOI22X1  _2725_
timestamp 0
transform 1 0 10390 0 1 250
box -6 -8 126 248
use AOI22X1  _2726_
timestamp 0
transform -1 0 9870 0 1 730
box -6 -8 126 248
use AOI21X1  _2727_
timestamp 0
transform 1 0 9970 0 1 730
box -6 -8 106 248
use OAI21X1  _2728_
timestamp 0
transform -1 0 10030 0 -1 1210
box -6 -8 106 248
use AOI22X1  _2729_
timestamp 0
transform -1 0 9650 0 -1 1690
box -6 -8 126 248
use OAI21X1  _2730_
timestamp 0
transform 1 0 11290 0 -1 2650
box -6 -8 106 248
use AOI21X1  _2731_
timestamp 0
transform 1 0 9530 0 -1 2650
box -6 -8 106 248
use NAND2X1  _2732_
timestamp 0
transform 1 0 6750 0 -1 2650
box -6 -8 86 248
use OAI21X1  _2733_
timestamp 0
transform -1 0 9250 0 -1 1690
box -6 -8 106 248
use MUX2X1  _2734_
timestamp 0
transform 1 0 9530 0 1 730
box -6 -8 126 248
use OAI21X1  _2735_
timestamp 0
transform 1 0 9530 0 -1 1210
box -6 -8 106 248
use OAI21X1  _2736_
timestamp 0
transform -1 0 9050 0 -1 1690
box -6 -8 106 248
use OAI21X1  _2737_
timestamp 0
transform -1 0 9430 0 1 730
box -6 -8 106 248
use AOI21X1  _2738_
timestamp 0
transform -1 0 10510 0 -1 250
box -6 -8 106 248
use AOI22X1  _2739_
timestamp 0
transform 1 0 10610 0 -1 250
box -6 -8 126 248
use OAI21X1  _2740_
timestamp 0
transform 1 0 11230 0 -1 250
box -6 -8 106 248
use INVX1  _2741_
timestamp 0
transform 1 0 11630 0 -1 250
box -6 -8 66 248
use OAI21X1  _2742_
timestamp 0
transform -1 0 10710 0 1 250
box -6 -8 106 248
use AOI21X1  _2743_
timestamp 0
transform -1 0 10550 0 1 2170
box -6 -8 106 248
use OAI22X1  _2744_
timestamp 0
transform 1 0 10550 0 1 3130
box -6 -8 126 248
use OAI21X1  _2745_
timestamp 0
transform -1 0 11290 0 -1 3610
box -6 -8 106 248
use NAND2X1  _2746_
timestamp 0
transform -1 0 10270 0 1 3130
box -6 -8 86 248
use OAI21X1  _2747_
timestamp 0
transform 1 0 11010 0 1 250
box -6 -8 106 248
use INVX1  _2748_
timestamp 0
transform 1 0 9870 0 -1 250
box -6 -8 66 248
use AOI21X1  _2749_
timestamp 0
transform 1 0 10730 0 1 730
box -6 -8 106 248
use NAND3X1  _2750_
timestamp 0
transform 1 0 11070 0 -1 1210
box -6 -8 106 248
use INVX1  _2751_
timestamp 0
transform -1 0 10230 0 1 730
box -6 -8 66 248
use OAI21X1  _2752_
timestamp 0
transform 1 0 5810 0 1 1210
box -6 -8 106 248
use NAND3X1  _2753_
timestamp 0
transform -1 0 6110 0 1 1210
box -6 -8 106 248
use NAND3X1  _2754_
timestamp 0
transform -1 0 6170 0 -1 1690
box -6 -8 106 248
use NAND3X1  _2755_
timestamp 0
transform -1 0 7510 0 -1 1690
box -6 -8 106 248
use OAI21X1  _2756_
timestamp 0
transform -1 0 7650 0 1 1210
box -6 -8 106 248
use INVX1  _2757_
timestamp 0
transform 1 0 8170 0 1 1210
box -6 -8 66 248
use OAI21X1  _2758_
timestamp 0
transform -1 0 7710 0 -1 1690
box -6 -8 106 248
use INVX1  _2759_
timestamp 0
transform -1 0 9810 0 -1 1690
box -6 -8 66 248
use OAI21X1  _2760_
timestamp 0
transform -1 0 6370 0 -1 1690
box -6 -8 106 248
use NOR2X1  _2761_
timestamp 0
transform -1 0 8990 0 1 1690
box -6 -8 86 248
use AOI22X1  _2762_
timestamp 0
transform -1 0 9010 0 1 2170
box -6 -8 126 248
use AOI21X1  _2763_
timestamp 0
transform -1 0 6450 0 1 1690
box -6 -8 106 248
use OAI21X1  _2764_
timestamp 0
transform -1 0 6530 0 -1 2170
box -6 -8 106 248
use NOR2X1  _2765_
timestamp 0
transform -1 0 9470 0 -1 3610
box -6 -8 86 248
use OAI21X1  _2766_
timestamp 0
transform -1 0 6830 0 1 1690
box -6 -8 106 248
use AOI21X1  _2767_
timestamp 0
transform 1 0 8970 0 -1 2650
box -6 -8 106 248
use OAI21X1  _2768_
timestamp 0
transform -1 0 6130 0 1 730
box -6 -8 106 248
use AOI21X1  _2769_
timestamp 0
transform -1 0 7070 0 1 730
box -6 -8 106 248
use NAND2X1  _2770_
timestamp 0
transform 1 0 7170 0 -1 730
box -6 -8 86 248
use OAI21X1  _2771_
timestamp 0
transform 1 0 10090 0 -1 730
box -6 -8 106 248
use NAND3X1  _2772_
timestamp 0
transform -1 0 7530 0 -1 1210
box -6 -8 106 248
use OAI21X1  _2773_
timestamp 0
transform -1 0 7730 0 -1 1210
box -6 -8 106 248
use NOR2X1  _2774_
timestamp 0
transform -1 0 6150 0 -1 1210
box -6 -8 86 248
use OAI21X1  _2775_
timestamp 0
transform -1 0 7450 0 1 1210
box -6 -8 106 248
use NOR2X1  _2776_
timestamp 0
transform 1 0 6210 0 1 1210
box -6 -8 86 248
use OAI21X1  _2777_
timestamp 0
transform -1 0 10010 0 1 1210
box -6 -8 106 248
use AOI22X1  _2778_
timestamp 0
transform 1 0 7750 0 1 1210
box -6 -8 126 248
use AOI21X1  _2779_
timestamp 0
transform 1 0 7970 0 1 1210
box -6 -8 106 248
use AOI21X1  _2780_
timestamp 0
transform 1 0 8030 0 -1 1210
box -6 -8 106 248
use OAI21X1  _2781_
timestamp 0
transform -1 0 7930 0 -1 1210
box -6 -8 106 248
use OAI21X1  _2782_
timestamp 0
transform 1 0 7710 0 1 1690
box -6 -8 106 248
use AOI21X1  _2783_
timestamp 0
transform -1 0 8590 0 1 2170
box -6 -8 106 248
use AOI21X1  _2784_
timestamp 0
transform -1 0 11130 0 1 2170
box -6 -8 106 248
use OAI22X1  _2785_
timestamp 0
transform 1 0 9570 0 -1 3610
box -6 -8 126 248
use AOI22X1  _2786_
timestamp 0
transform -1 0 7930 0 -1 2170
box -6 -8 126 248
use AOI21X1  _2787_
timestamp 0
transform -1 0 9350 0 -1 2170
box -6 -8 106 248
use OAI21X1  _2788_
timestamp 0
transform -1 0 10330 0 -1 2170
box -6 -8 106 248
use INVX1  _2789_
timestamp 0
transform 1 0 10430 0 -1 2170
box -6 -8 66 248
use OAI21X1  _2790_
timestamp 0
transform 1 0 8030 0 -1 2170
box -6 -8 106 248
use OAI21X1  _2791_
timestamp 0
transform 1 0 8230 0 -1 2170
box -6 -8 106 248
use INVX1  _2792_
timestamp 0
transform -1 0 7730 0 -1 2650
box -6 -8 66 248
use NAND3X1  _2793_
timestamp 0
transform -1 0 7990 0 1 2650
box -6 -8 106 248
use AOI21X1  _2794_
timestamp 0
transform -1 0 7990 0 1 2170
box -6 -8 106 248
use OAI22X1  _2795_
timestamp 0
transform -1 0 7710 0 -1 2170
box -6 -8 126 248
use OAI21X1  _2796_
timestamp 0
transform -1 0 7110 0 -1 2170
box -6 -8 106 248
use OAI21X1  _2797_
timestamp 0
transform -1 0 8530 0 -1 2170
box -6 -8 106 248
use OAI21X1  _2798_
timestamp 0
transform 1 0 11990 0 -1 3610
box -6 -8 106 248
use OAI22X1  _2799_
timestamp 0
transform -1 0 7510 0 -1 2170
box -6 -8 126 248
use OAI21X1  _2800_
timestamp 0
transform -1 0 7610 0 1 1690
box -6 -8 106 248
use NAND3X1  _2801_
timestamp 0
transform 1 0 7170 0 1 1210
box -6 -8 106 248
use OAI21X1  _2802_
timestamp 0
transform 1 0 6830 0 -1 1210
box -6 -8 106 248
use AOI21X1  _2803_
timestamp 0
transform -1 0 7130 0 -1 1210
box -6 -8 106 248
use OAI21X1  _2804_
timestamp 0
transform -1 0 8630 0 1 1210
box -6 -8 106 248
use OAI21X1  _2805_
timestamp 0
transform 1 0 6970 0 1 1210
box -6 -8 106 248
use NOR2X1  _2806_
timestamp 0
transform -1 0 6930 0 -1 1690
box -6 -8 86 248
use NOR2X1  _2807_
timestamp 0
transform -1 0 7190 0 1 2650
box -6 -8 86 248
use AOI22X1  _2808_
timestamp 0
transform 1 0 10210 0 1 1690
box -6 -8 126 248
use MUX2X1  _2809_
timestamp 0
transform -1 0 10730 0 1 1690
box -6 -8 126 248
use OAI21X1  _2810_
timestamp 0
transform 1 0 10610 0 -1 1690
box -6 -8 106 248
use NOR2X1  _2811_
timestamp 0
transform 1 0 10430 0 -1 1690
box -6 -8 86 248
use OAI21X1  _2812_
timestamp 0
transform 1 0 10290 0 1 1210
box -6 -8 106 248
use NOR2X1  _2813_
timestamp 0
transform -1 0 10190 0 1 1210
box -6 -8 86 248
use AOI21X1  _2814_
timestamp 0
transform -1 0 10610 0 -1 2650
box -6 -8 106 248
use NAND3X1  _2815_
timestamp 0
transform -1 0 10790 0 -1 2650
box -6 -8 106 248
use OAI21X1  _2816_
timestamp 0
transform 1 0 10250 0 1 2170
box -6 -8 106 248
use NAND2X1  _2817_
timestamp 0
transform -1 0 10410 0 -1 2650
box -6 -8 86 248
use OAI21X1  _2818_
timestamp 0
transform -1 0 11090 0 -1 1690
box -6 -8 106 248
use AOI21X1  _2819_
timestamp 0
transform -1 0 11190 0 1 1210
box -6 -8 106 248
use AOI21X1  _2820_
timestamp 0
transform -1 0 11390 0 1 1210
box -6 -8 106 248
use NAND3X1  _2821_
timestamp 0
transform 1 0 11070 0 -1 730
box -6 -8 106 248
use NAND3X1  _2822_
timestamp 0
transform -1 0 12090 0 1 250
box -6 -8 106 248
use OAI21X1  _2823_
timestamp 0
transform 1 0 11190 0 -1 1690
box -6 -8 106 248
use NAND2X1  _2824_
timestamp 0
transform 1 0 10690 0 -1 1210
box -6 -8 86 248
use OAI21X1  _2825_
timestamp 0
transform 1 0 11210 0 1 1690
box -6 -8 106 248
use NAND3X1  _2826_
timestamp 0
transform 1 0 11410 0 1 1690
box -6 -8 106 248
use NAND3X1  _2827_
timestamp 0
transform -1 0 11950 0 1 730
box -6 -8 106 248
use OAI22X1  _2828_
timestamp 0
transform -1 0 12090 0 1 1690
box -6 -8 126 248
use AOI22X1  _2829_
timestamp 0
transform -1 0 11530 0 1 2170
box -6 -8 126 248
use AOI22X1  _2830_
timestamp 0
transform 1 0 11070 0 -1 2650
box -6 -8 126 248
use AOI21X1  _2831_
timestamp 0
transform 1 0 11130 0 1 3130
box -6 -8 106 248
use OAI21X1  _2832_
timestamp 0
transform -1 0 11450 0 1 2650
box -6 -8 106 248
use OAI21X1  _2833_
timestamp 0
transform 1 0 11430 0 -1 1210
box -6 -8 106 248
use OAI21X1  _2834_
timestamp 0
transform 1 0 11930 0 -1 2170
box -6 -8 106 248
use OAI21X1  _2835_
timestamp 0
transform 1 0 12090 0 -1 11770
box -6 -8 106 248
use AOI21X1  _2836_
timestamp 0
transform 1 0 11730 0 -1 1690
box -6 -8 106 248
use OAI21X1  _2837_
timestamp 0
transform 1 0 11930 0 -1 1690
box -6 -8 106 248
use AOI21X1  _2838_
timestamp 0
transform 1 0 12050 0 1 1210
box -6 -8 106 248
use NAND3X1  _2839_
timestamp 0
transform 1 0 11630 0 -1 1210
box -6 -8 106 248
use NAND2X1  _2840_
timestamp 0
transform -1 0 11890 0 1 250
box -6 -8 86 248
use NAND2X1  _2841_
timestamp 0
transform -1 0 11750 0 1 730
box -6 -8 86 248
use AOI21X1  _2842_
timestamp 0
transform -1 0 9950 0 1 2170
box -6 -8 106 248
use AOI21X1  _2843_
timestamp 0
transform -1 0 10150 0 1 2170
box -6 -8 106 248
use OAI21X1  _2844_
timestamp 0
transform -1 0 11930 0 1 2170
box -6 -8 106 248
use OAI21X1  _2845_
timestamp 0
transform 1 0 12030 0 1 2170
box -6 -8 106 248
use NOR2X1  _2846_
timestamp 0
transform 1 0 11590 0 1 11770
box -6 -8 86 248
use OAI21X1  _2847_
timestamp 0
transform 1 0 12010 0 -1 1210
box -6 -8 106 248
use OAI21X1  _2848_
timestamp 0
transform -1 0 11730 0 1 2170
box -6 -8 106 248
use AOI21X1  _2849_
timestamp 0
transform -1 0 11830 0 1 2650
box -6 -8 106 248
use NOR2X1  _2850_
timestamp 0
transform 1 0 11930 0 1 2650
box -6 -8 86 248
use NAND3X1  _2851_
timestamp 0
transform -1 0 10010 0 -1 3130
box -6 -8 106 248
use OR2X2  _2852_
timestamp 0
transform -1 0 11190 0 -1 3130
box -6 -8 106 248
use OAI21X1  _2853_
timestamp 0
transform 1 0 11290 0 -1 3130
box -6 -8 106 248
use OAI21X1  _2854_
timestamp 0
transform 1 0 11870 0 -1 3130
box -6 -8 106 248
use OAI21X1  _2855_
timestamp 0
transform 1 0 11850 0 -1 2650
box -6 -8 106 248
use OAI21X1  _2856_
timestamp 0
transform -1 0 9970 0 1 2650
box -6 -8 106 248
use AOI21X1  _2857_
timestamp 0
transform -1 0 10030 0 -1 2650
box -6 -8 106 248
use OAI21X1  _2858_
timestamp 0
transform -1 0 8190 0 1 2170
box -6 -8 106 248
use OAI21X1  _2859_
timestamp 0
transform 1 0 9730 0 -1 2650
box -6 -8 106 248
use NAND2X1  _2860_
timestamp 0
transform -1 0 9250 0 -1 2650
box -6 -8 86 248
use NAND3X1  _2861_
timestamp 0
transform 1 0 10010 0 1 1690
box -6 -8 106 248
use NAND3X1  _2862_
timestamp 0
transform 1 0 9610 0 1 1690
box -6 -8 106 248
use OAI21X1  _2863_
timestamp 0
transform 1 0 8830 0 -1 2170
box -6 -8 106 248
use OAI21X1  _2864_
timestamp 0
transform -1 0 7910 0 -1 1690
box -6 -8 106 248
use NAND2X1  _2865_
timestamp 0
transform -1 0 6550 0 -1 1690
box -6 -8 86 248
use OAI21X1  _2866_
timestamp 0
transform -1 0 8990 0 1 2650
box -6 -8 106 248
use NAND2X1  _2867_
timestamp 0
transform -1 0 9510 0 1 1690
box -6 -8 86 248
use OAI21X1  _2868_
timestamp 0
transform 1 0 9250 0 1 2170
box -6 -8 106 248
use NAND2X1  _2869_
timestamp 0
transform -1 0 10670 0 1 2650
box -6 -8 86 248
use OAI21X1  _2870_
timestamp 0
transform -1 0 9450 0 -1 4090
box -6 -8 106 248
use INVX2  _2871_
timestamp 0
transform -1 0 8650 0 -1 250
box -6 -8 66 248
use OAI21X1  _2872_
timestamp 0
transform 1 0 9810 0 1 1690
box -6 -8 106 248
use AOI21X1  _2873_
timestamp 0
transform 1 0 9850 0 -1 2170
box -6 -8 106 248
use OAI21X1  _2874_
timestamp 0
transform 1 0 9650 0 1 2170
box -6 -8 106 248
use NAND3X1  _2875_
timestamp 0
transform -1 0 11310 0 1 4090
box -6 -8 106 248
use INVX2  _2876_
timestamp 0
transform 1 0 10250 0 1 2650
box -6 -8 66 248
use OAI21X1  _2877_
timestamp 0
transform -1 0 10870 0 1 2650
box -6 -8 106 248
use AOI21X1  _2878_
timestamp 0
transform 1 0 9690 0 -1 730
box -6 -8 106 248
use OAI21X1  _2879_
timestamp 0
transform -1 0 9990 0 -1 730
box -6 -8 106 248
use NAND2X1  _2880_
timestamp 0
transform -1 0 10290 0 1 250
box -6 -8 86 248
use NAND2X1  _2881_
timestamp 0
transform -1 0 6070 0 -1 730
box -6 -8 86 248
use NAND3X1  _2882_
timestamp 0
transform -1 0 6270 0 -1 730
box -6 -8 106 248
use OAI21X1  _2883_
timestamp 0
transform -1 0 5630 0 1 2650
box -6 -8 106 248
use AOI21X1  _2884_
timestamp 0
transform -1 0 5630 0 -1 2650
box -6 -8 106 248
use AOI22X1  _2885_
timestamp 0
transform 1 0 5530 0 1 1690
box -6 -8 126 248
use AOI21X1  _2886_
timestamp 0
transform -1 0 5430 0 1 1690
box -6 -8 106 248
use OAI21X1  _2887_
timestamp 0
transform 1 0 5690 0 -1 1690
box -6 -8 106 248
use OAI22X1  _2888_
timestamp 0
transform 1 0 6110 0 1 2650
box -6 -8 126 248
use OAI21X1  _2889_
timestamp 0
transform -1 0 6430 0 1 2650
box -6 -8 106 248
use AOI21X1  _2890_
timestamp 0
transform -1 0 6810 0 1 2650
box -6 -8 106 248
use AOI21X1  _2891_
timestamp 0
transform 1 0 8210 0 -1 2650
box -6 -8 106 248
use NAND3X1  _2892_
timestamp 0
transform -1 0 7410 0 -1 2650
box -6 -8 106 248
use OAI21X1  _2893_
timestamp 0
transform -1 0 6010 0 1 2650
box -6 -8 106 248
use NAND3X1  _2894_
timestamp 0
transform 1 0 5430 0 -1 2170
box -6 -8 106 248
use NAND2X1  _2895_
timestamp 0
transform -1 0 7570 0 -1 2650
box -6 -8 86 248
use NOR2X1  _2896_
timestamp 0
transform -1 0 6710 0 -1 2170
box -6 -8 86 248
use NAND3X1  _2897_
timestamp 0
transform 1 0 7390 0 -1 3130
box -6 -8 106 248
use NAND2X1  _2898_
timestamp 0
transform 1 0 11810 0 -1 3610
box -6 -8 86 248
use NAND3X1  _2899_
timestamp 0
transform -1 0 6670 0 -1 730
box -6 -8 106 248
use NAND3X1  _2900_
timestamp 0
transform -1 0 6870 0 -1 730
box -6 -8 106 248
use OAI21X1  _2901_
timestamp 0
transform -1 0 8310 0 -1 250
box -6 -8 106 248
use NOR2X1  _2902_
timestamp 0
transform 1 0 9690 0 -1 250
box -6 -8 86 248
use OAI21X1  _2903_
timestamp 0
transform -1 0 11710 0 1 250
box -6 -8 106 248
use NOR2X1  _2904_
timestamp 0
transform 1 0 8410 0 -1 250
box -6 -8 86 248
use OAI21X1  _2905_
timestamp 0
transform -1 0 7070 0 -1 730
box -6 -8 106 248
use AOI21X1  _2906_
timestamp 0
transform -1 0 7450 0 -1 730
box -6 -8 106 248
use OAI21X1  _2907_
timestamp 0
transform -1 0 6470 0 -1 730
box -6 -8 106 248
use OAI21X1  _2908_
timestamp 0
transform 1 0 8510 0 -1 730
box -6 -8 106 248
use AOI21X1  _2909_
timestamp 0
transform -1 0 10490 0 -1 3610
box -6 -8 106 248
use NOR2X1  _2910_
timestamp 0
transform 1 0 10810 0 -1 3610
box -6 -8 86 248
use AOI21X1  _2911_
timestamp 0
transform 1 0 10990 0 -1 3610
box -6 -8 106 248
use OAI21X1  _2912_
timestamp 0
transform -1 0 10930 0 1 3610
box -6 -8 106 248
use OAI21X1  _2913_
timestamp 0
transform -1 0 8810 0 -1 730
box -6 -8 106 248
use NAND2X1  _2914_
timestamp 0
transform -1 0 8670 0 -1 1210
box -6 -8 86 248
use NAND2X1  _2915_
timestamp 0
transform -1 0 11330 0 -1 1210
box -6 -8 86 248
use NAND2X1  _2916_
timestamp 0
transform -1 0 8090 0 -1 1690
box -6 -8 86 248
use NAND3X1  _2917_
timestamp 0
transform -1 0 7130 0 1 250
box -6 -8 106 248
use NAND3X1  _2918_
timestamp 0
transform 1 0 6830 0 1 250
box -6 -8 106 248
use NAND3X1  _2919_
timestamp 0
transform -1 0 7330 0 1 250
box -6 -8 106 248
use NAND3X1  _2920_
timestamp 0
transform 1 0 7210 0 -1 250
box -6 -8 106 248
use OAI21X1  _2921_
timestamp 0
transform 1 0 7010 0 -1 250
box -6 -8 106 248
use INVX1  _2922_
timestamp 0
transform 1 0 6670 0 1 250
box -6 -8 66 248
use OAI21X1  _2923_
timestamp 0
transform -1 0 5970 0 -1 1210
box -6 -8 106 248
use OAI21X1  _2924_
timestamp 0
transform 1 0 8930 0 -1 250
box -6 -8 106 248
use OAI21X1  _2925_
timestamp 0
transform 1 0 10290 0 -1 730
box -6 -8 106 248
use NAND2X1  _2926_
timestamp 0
transform 1 0 12030 0 -1 730
box -6 -8 86 248
use NOR2X1  _2927_
timestamp 0
transform 1 0 8750 0 -1 250
box -6 -8 86 248
use OR2X2  _2928_
timestamp 0
transform 1 0 7550 0 -1 730
box -6 -8 106 248
use NAND3X1  _2929_
timestamp 0
transform 1 0 8270 0 1 250
box -6 -8 106 248
use INVX1  _2930_
timestamp 0
transform -1 0 8530 0 1 250
box -6 -8 66 248
use OAI21X1  _2931_
timestamp 0
transform -1 0 8210 0 -1 730
box -6 -8 106 248
use NAND2X1  _2932_
timestamp 0
transform 1 0 7930 0 -1 730
box -6 -8 86 248
use NAND2X1  _2933_
timestamp 0
transform 1 0 7970 0 1 730
box -6 -8 86 248
use INVX2  _2934_
timestamp 0
transform -1 0 10310 0 -1 250
box -6 -8 66 248
use NAND2X1  _2935_
timestamp 0
transform 1 0 11370 0 -1 1690
box -6 -8 86 248
use NAND3X1  _2936_
timestamp 0
transform -1 0 8330 0 -1 1210
box -6 -8 106 248
use NOR2X1  _2937_
timestamp 0
transform 1 0 8730 0 1 1210
box -6 -8 86 248
use NAND2X1  _2938_
timestamp 0
transform -1 0 11910 0 -1 1210
box -6 -8 86 248
use NAND2X1  _2939_
timestamp 0
transform -1 0 11350 0 -1 730
box -6 -8 86 248
use OAI21X1  _2940_
timestamp 0
transform -1 0 6710 0 -1 3130
box -6 -8 106 248
use AOI21X1  _2941_
timestamp 0
transform 1 0 8910 0 1 3610
box -6 -8 106 248
use NAND2X1  _2942_
timestamp 0
transform 1 0 8990 0 -1 4090
box -6 -8 86 248
use OAI21X1  _2943_
timestamp 0
transform 1 0 9750 0 -1 4090
box -6 -8 106 248
use NOR2X1  _2944_
timestamp 0
transform 1 0 9930 0 1 4090
box -6 -8 86 248
use INVX1  _2945_
timestamp 0
transform 1 0 9110 0 1 3610
box -6 -8 66 248
use OAI21X1  _2946_
timestamp 0
transform -1 0 9290 0 -1 3610
box -6 -8 106 248
use INVX1  _2947_
timestamp 0
transform -1 0 8810 0 1 3610
box -6 -8 66 248
use OAI21X1  _2948_
timestamp 0
transform -1 0 8790 0 1 2170
box -6 -8 106 248
use NAND2X1  _2949_
timestamp 0
transform 1 0 10890 0 -1 2650
box -6 -8 86 248
use NAND2X1  _2950_
timestamp 0
transform 1 0 11710 0 -1 4090
box -6 -8 86 248
use AOI21X1  _2951_
timestamp 0
transform -1 0 7110 0 -1 3130
box -6 -8 106 248
use OAI21X1  _2952_
timestamp 0
transform -1 0 6910 0 -1 3130
box -6 -8 106 248
use NOR2X1  _2953_
timestamp 0
transform 1 0 11330 0 1 3130
box -6 -8 86 248
use NAND2X1  _2954_
timestamp 0
transform -1 0 9070 0 -1 3130
box -6 -8 86 248
use OAI22X1  _2955_
timestamp 0
transform -1 0 10230 0 -1 2650
box -6 -8 126 248
use OAI21X1  _2956_
timestamp 0
transform -1 0 11490 0 -1 3610
box -6 -8 106 248
use NOR2X1  _2957_
timestamp 0
transform 1 0 9730 0 1 1210
box -6 -8 86 248
use AND2X2  _2958_
timestamp 0
transform 1 0 11690 0 1 3130
box -6 -8 106 248
use INVX4  _2959_
timestamp 0
transform 1 0 5170 0 1 2170
box -6 -8 86 248
use OAI21X1  _2960_
timestamp 0
transform -1 0 7510 0 -1 250
box -6 -8 106 248
use AOI21X1  _2961_
timestamp 0
transform -1 0 8110 0 -1 250
box -6 -8 106 248
use OAI21X1  _2962_
timestamp 0
transform -1 0 7710 0 -1 250
box -6 -8 106 248
use NAND2X1  _2963_
timestamp 0
transform -1 0 6610 0 1 2650
box -6 -8 86 248
use AND2X2  _2964_
timestamp 0
transform -1 0 7910 0 -1 250
box -6 -8 106 248
use NOR2X1  _2965_
timestamp 0
transform -1 0 11870 0 -1 250
box -6 -8 86 248
use OAI21X1  _2966_
timestamp 0
transform 1 0 8630 0 1 250
box -6 -8 106 248
use OAI21X1  _2967_
timestamp 0
transform 1 0 9330 0 1 1210
box -6 -8 106 248
use NOR2X1  _2968_
timestamp 0
transform 1 0 10450 0 1 3610
box -6 -8 86 248
use NOR2X1  _2969_
timestamp 0
transform 1 0 10650 0 1 4090
box -6 -8 86 248
use INVX4  _2970_
timestamp 0
transform -1 0 11390 0 1 730
box -6 -8 86 248
use NAND2X1  _2971_
timestamp 0
transform 1 0 7790 0 -1 4090
box -6 -8 86 248
use NOR2X1  _2972_
timestamp 0
transform -1 0 9450 0 -1 1210
box -6 -8 86 248
use AND2X2  _2973_
timestamp 0
transform 1 0 7430 0 1 250
box -6 -8 106 248
use AOI22X1  _2974_
timestamp 0
transform -1 0 7470 0 1 730
box -6 -8 126 248
use INVX1  _2975_
timestamp 0
transform -1 0 9150 0 1 2170
box -6 -8 66 248
use NAND2X1  _2976_
timestamp 0
transform 1 0 10110 0 -1 3130
box -6 -8 86 248
use INVX8  _2977_
timestamp 0
transform 1 0 10510 0 1 730
box -6 -8 126 248
use NAND3X1  _2978_
timestamp 0
transform -1 0 11750 0 -1 730
box -6 -8 106 248
use INVX4  _2979_
timestamp 0
transform -1 0 11970 0 -1 4090
box -6 -8 86 248
use OAI21X1  _2980_
timestamp 0
transform 1 0 7230 0 -1 1210
box -6 -8 106 248
use OAI21X1  _2981_
timestamp 0
transform 1 0 6630 0 -1 1210
box -6 -8 106 248
use NOR2X1  _2982_
timestamp 0
transform 1 0 7570 0 1 730
box -6 -8 86 248
use INVX8  _2983_
timestamp 0
transform 1 0 11950 0 1 4090
box -6 -8 126 248
use NAND2X1  _2984_
timestamp 0
transform 1 0 11690 0 -1 3130
box -6 -8 86 248
use INVX8  _2985_
timestamp 0
transform -1 0 7290 0 -1 3610
box -6 -8 126 248
use INVX8  _2986_
timestamp 0
transform -1 0 7310 0 1 3610
box -6 -8 126 248
use INVX2  _2987_
timestamp 0
transform 1 0 5870 0 1 3130
box -6 -8 66 248
use DFFSR  _2988_
timestamp 0
transform 1 0 3070 0 1 1690
box -6 -8 486 248
use DFFSR  _2989_
timestamp 0
transform 1 0 3150 0 1 2650
box -6 -8 486 248
use DFFPOSX1  _2990_
timestamp 0
transform 1 0 4270 0 -1 2170
box -6 -8 246 248
use DFFSR  _2991_
timestamp 0
transform -1 0 5070 0 -1 2650
box -6 -8 486 248
use DFFSR  _2992_
timestamp 0
transform 1 0 3950 0 -1 2650
box -6 -8 486 248
use DFFSR  _2993_
timestamp 0
transform 1 0 2870 0 -1 2170
box -6 -8 486 248
use DFFSR  _2994_
timestamp 0
transform -1 0 5350 0 -1 3130
box -6 -8 486 248
use DFFSR  _2995_
timestamp 0
transform 1 0 1630 0 -1 2170
box -6 -8 486 248
use DFFSR  _2996_
timestamp 0
transform 1 0 1670 0 -1 2650
box -6 -8 486 248
use DFFSR  _2997_
timestamp 0
transform 1 0 3110 0 1 2170
box -6 -8 486 248
use DFFSR  _2998_
timestamp 0
transform 1 0 5350 0 -1 3130
box -6 -8 486 248
use DFFSR  _2999_
timestamp 0
transform 1 0 2370 0 1 1690
box -6 -8 486 248
use MUX2X1  _3000_
timestamp 0
transform -1 0 2370 0 1 2170
box -6 -8 126 248
use INVX1  _3001_
timestamp 0
transform 1 0 2410 0 -1 3130
box -6 -8 66 248
use INVX1  _3002_
timestamp 0
transform 1 0 2210 0 -1 2170
box -6 -8 66 248
use MUX2X1  _3003_
timestamp 0
transform -1 0 3790 0 -1 2650
box -6 -8 126 248
use INVX1  _3004_
timestamp 0
transform 1 0 3890 0 -1 2650
box -6 -8 66 248
use INVX1  _3005_
timestamp 0
transform -1 0 3570 0 -1 2650
box -6 -8 66 248
use AOI22X1  _3006_
timestamp 0
transform -1 0 4510 0 1 2650
box -6 -8 126 248
use NAND3X1  _3007_
timestamp 0
transform -1 0 4290 0 1 2650
box -6 -8 106 248
use NOR3X1  _3008_
timestamp 0
transform 1 0 3910 0 1 2650
box -6 -8 186 248
use NAND3X1  _3009_
timestamp 0
transform 1 0 4030 0 -1 3130
box -6 -8 106 248
use NOR2X1  _3010_
timestamp 0
transform -1 0 4110 0 1 3130
box -6 -8 86 248
use NOR2X1  _3011_
timestamp 0
transform 1 0 3850 0 -1 3130
box -6 -8 86 248
use NAND3X1  _3012_
timestamp 0
transform 1 0 2790 0 -1 2650
box -6 -8 106 248
use NOR2X1  _3013_
timestamp 0
transform -1 0 2550 0 1 2170
box -6 -8 86 248
use INVX1  _3014_
timestamp 0
transform 1 0 2630 0 -1 2650
box -6 -8 66 248
use NOR2X1  _3015_
timestamp 0
transform -1 0 4670 0 -1 3130
box -6 -8 86 248
use INVX1  _3016_
timestamp 0
transform 1 0 4530 0 -1 2650
box -6 -8 66 248
use OAI21X1  _3017_
timestamp 0
transform 1 0 4230 0 1 2170
box -6 -8 106 248
use OAI21X1  _3018_
timestamp 0
transform 1 0 4430 0 1 2170
box -6 -8 106 248
use OAI21X1  _3019_
timestamp 0
transform -1 0 4130 0 1 2170
box -6 -8 106 248
use MUX2X1  _3020_
timestamp 0
transform 1 0 1870 0 1 2170
box -6 -8 126 248
use INVX1  _3021_
timestamp 0
transform 1 0 1710 0 1 2170
box -6 -8 66 248
use INVX1  _3022_
timestamp 0
transform -1 0 2150 0 1 2170
box -6 -8 66 248
use INVX4  _3023_
timestamp 0
transform -1 0 3010 0 -1 3130
box -6 -8 86 248
use OAI21X1  _3024_
timestamp 0
transform 1 0 4770 0 -1 3130
box -6 -8 106 248
use OAI21X1  _3025_
timestamp 0
transform 1 0 4390 0 -1 3130
box -6 -8 106 248
use NAND3X1  _3026_
timestamp 0
transform 1 0 3650 0 -1 3130
box -6 -8 106 248
use INVX1  _3027_
timestamp 0
transform 1 0 3350 0 -1 2650
box -6 -8 66 248
use INVX1  _3028_
timestamp 0
transform -1 0 2870 0 1 2650
box -6 -8 66 248
use INVX1  _3029_
timestamp 0
transform 1 0 3490 0 -1 3130
box -6 -8 66 248
use AOI21X1  _3030_
timestamp 0
transform 1 0 4930 0 1 2650
box -6 -8 106 248
use INVX1  _3031_
timestamp 0
transform 1 0 4770 0 1 2650
box -6 -8 66 248
use INVX1  _3032_
timestamp 0
transform 1 0 5930 0 -1 3130
box -6 -8 66 248
use OAI21X1  _3033_
timestamp 0
transform -1 0 4730 0 1 2170
box -6 -8 106 248
use INVX1  _3034_
timestamp 0
transform 1 0 3870 0 1 2170
box -6 -8 66 248
use INVX1  _3035_
timestamp 0
transform -1 0 4670 0 1 2650
box -6 -8 66 248
use MUX2X1  _3036_
timestamp 0
transform -1 0 2530 0 -1 2650
box -6 -8 126 248
use INVX1  _3037_
timestamp 0
transform -1 0 3410 0 -1 3610
box -6 -8 66 248
use INVX1  _3038_
timestamp 0
transform 1 0 2250 0 -1 2650
box -6 -8 66 248
use MUX2X1  _3039_
timestamp 0
transform -1 0 3730 0 -1 1690
box -6 -8 126 248
use INVX1  _3040_
timestamp 0
transform -1 0 3890 0 -1 1690
box -6 -8 66 248
use INVX1  _3041_
timestamp 0
transform 1 0 3450 0 -1 1690
box -6 -8 66 248
use MUX2X1  _3042_
timestamp 0
transform -1 0 2930 0 1 2170
box -6 -8 126 248
use INVX1  _3043_
timestamp 0
transform -1 0 3910 0 1 3610
box -6 -8 66 248
use INVX1  _3044_
timestamp 0
transform -1 0 2710 0 1 2170
box -6 -8 66 248
use MUX2X1  _3045_
timestamp 0
transform -1 0 3070 0 1 1690
box -6 -8 126 248
use INVX1  _3046_
timestamp 0
transform -1 0 3350 0 -1 1690
box -6 -8 66 248
use INVX1  _3047_
timestamp 0
transform 1 0 2910 0 -1 1690
box -6 -8 66 248
use INVX1  _3048_
timestamp 0
transform 1 0 3430 0 -1 2170
box -6 -8 66 248
use NAND3X1  _3049_
timestamp 0
transform -1 0 3830 0 1 2650
box -6 -8 106 248
use NOR3X1  _3050_
timestamp 0
transform -1 0 3150 0 1 2650
box -6 -8 186 248
use NAND2X1  _3051_
timestamp 0
transform -1 0 3070 0 -1 2650
box -6 -8 86 248
use NOR2X1  _3052_
timestamp 0
transform 1 0 3170 0 -1 2650
box -6 -8 86 248
use NOR2X1  _3053_
timestamp 0
transform -1 0 3110 0 1 2170
box -6 -8 86 248
use NAND3X1  _3054_
timestamp 0
transform -1 0 2730 0 1 2650
box -6 -8 106 248
use NOR2X1  _3055_
timestamp 0
transform -1 0 2530 0 1 2650
box -6 -8 86 248
use INVX1  _3056_
timestamp 0
transform -1 0 2830 0 -1 3130
box -6 -8 66 248
use NAND3X1  _3057_
timestamp 0
transform -1 0 3390 0 -1 3130
box -6 -8 106 248
use INVX1  _3058_
timestamp 0
transform 1 0 4230 0 -1 3130
box -6 -8 66 248
use NAND3X1  _3059_
timestamp 0
transform -1 0 5230 0 1 2650
box -6 -8 106 248
use AND2X2  _3060_
timestamp 0
transform -1 0 5430 0 1 2650
box -6 -8 106 248
use INVX1  _3061_
timestamp 0
transform -1 0 6150 0 -1 3130
box -6 -8 66 248
use NOR2X1  _3062_
timestamp 0
transform -1 0 5230 0 1 1690
box -6 -8 86 248
use NOR2X1  _3063_
timestamp 0
transform -1 0 5250 0 -1 2650
box -6 -8 86 248
use INVX1  _3064_
timestamp 0
transform -1 0 5070 0 1 2170
box -6 -8 66 248
use DFFSR  _3065_
timestamp 0
transform -1 0 1470 0 1 730
box -6 -8 486 248
use DFFSR  _3066_
timestamp 0
transform 1 0 870 0 1 1210
box -6 -8 486 248
use DFFSR  _3067_
timestamp 0
transform 1 0 530 0 -1 250
box -6 -8 486 248
use DFFSR  _3068_
timestamp 0
transform 1 0 1010 0 -1 250
box -6 -8 486 248
use DFFSR  _3069_
timestamp 0
transform 1 0 190 0 -1 1690
box -6 -8 486 248
use DFFSR  _3070_
timestamp 0
transform -1 0 850 0 -1 730
box -6 -8 486 248
use DFFSR  _3071_
timestamp 0
transform 1 0 10 0 1 1210
box -6 -8 486 248
use DFFSR  _3072_
timestamp 0
transform 1 0 1790 0 1 250
box -6 -8 486 248
use DFFSR  _3073_
timestamp 0
transform 1 0 1390 0 -1 730
box -6 -8 486 248
use DFFSR  _3074_
timestamp 0
transform 1 0 190 0 1 250
box -6 -8 486 248
use DFFSR  _3075_
timestamp 0
transform 1 0 1510 0 -1 1210
box -6 -8 486 248
use OAI21X1  _3076_
timestamp 0
transform 1 0 1130 0 1 250
box -6 -8 106 248
use OAI21X1  _3077_
timestamp 0
transform -1 0 1430 0 1 250
box -6 -8 106 248
use INVX1  _3078_
timestamp 0
transform 1 0 970 0 1 250
box -6 -8 66 248
use AOI22X1  _3079_
timestamp 0
transform 1 0 1030 0 -1 1210
box -6 -8 126 248
use NAND2X1  _3080_
timestamp 0
transform -1 0 990 0 1 730
box -6 -8 86 248
use NOR2X1  _3081_
timestamp 0
transform 1 0 870 0 -1 1210
box -6 -8 86 248
use INVX1  _3082_
timestamp 0
transform 1 0 1450 0 -1 1210
box -6 -8 66 248
use OAI21X1  _3083_
timestamp 0
transform -1 0 1690 0 -1 250
box -6 -8 106 248
use OAI21X1  _3084_
timestamp 0
transform 1 0 1530 0 1 250
box -6 -8 106 248
use INVX1  _3085_
timestamp 0
transform -1 0 1850 0 -1 250
box -6 -8 66 248
use OAI22X1  _3086_
timestamp 0
transform -1 0 610 0 1 730
box -6 -8 126 248
use NAND3X1  _3087_
timestamp 0
transform -1 0 770 0 -1 1210
box -6 -8 106 248
use NAND2X1  _3088_
timestamp 0
transform 1 0 490 0 -1 1210
box -6 -8 86 248
use NOR3X1  _3089_
timestamp 0
transform -1 0 1630 0 1 1210
box -6 -8 186 248
use NAND3X1  _3090_
timestamp 0
transform 1 0 1270 0 -1 1690
box -6 -8 106 248
use NAND2X1  _3091_
timestamp 0
transform -1 0 2010 0 1 1210
box -6 -8 86 248
use AOI21X1  _3092_
timestamp 0
transform -1 0 810 0 1 730
box -6 -8 106 248
use OAI21X1  _3093_
timestamp 0
transform -1 0 210 0 -1 730
box -6 -8 106 248
use AOI21X1  _3094_
timestamp 0
transform -1 0 210 0 1 730
box -6 -8 106 248
use NOR2X1  _3095_
timestamp 0
transform -1 0 390 0 1 730
box -6 -8 86 248
use INVX1  _3096_
timestamp 0
transform -1 0 370 0 -1 730
box -6 -8 66 248
use OAI21X1  _3097_
timestamp 0
transform 1 0 2090 0 -1 250
box -6 -8 106 248
use OAI21X1  _3098_
timestamp 0
transform -1 0 2470 0 1 250
box -6 -8 106 248
use INVX1  _3099_
timestamp 0
transform 1 0 1930 0 -1 250
box -6 -8 66 248
use INVX4  _3100_
timestamp 0
transform 1 0 110 0 -1 1690
box -6 -8 86 248
use AOI21X1  _3101_
timestamp 0
transform -1 0 210 0 -1 1210
box -6 -8 106 248
use OAI21X1  _3102_
timestamp 0
transform -1 0 1390 0 -1 730
box -6 -8 106 248
use OAI21X1  _3103_
timestamp 0
transform -1 0 1350 0 -1 1210
box -6 -8 106 248
use NAND3X1  _3104_
timestamp 0
transform -1 0 390 0 1 1690
box -6 -8 106 248
use AND2X2  _3105_
timestamp 0
transform -1 0 1310 0 1 1690
box -6 -8 106 248
use NOR2X1  _3106_
timestamp 0
transform -1 0 2450 0 -1 2170
box -6 -8 86 248
use NOR2X1  _3107_
timestamp 0
transform -1 0 1650 0 1 1690
box -6 -8 86 248
use NOR2X1  _3108_
timestamp 0
transform -1 0 530 0 1 2170
box -6 -8 86 248
use OR2X2  _3109_
timestamp 0
transform -1 0 730 0 1 2170
box -6 -8 106 248
use NAND2X1  _3110_
timestamp 0
transform 1 0 790 0 -1 2170
box -6 -8 86 248
use INVX1  _3111_
timestamp 0
transform -1 0 1030 0 -1 2170
box -6 -8 66 248
use NOR2X1  _3112_
timestamp 0
transform -1 0 190 0 1 1690
box -6 -8 86 248
use NAND2X1  _3113_
timestamp 0
transform -1 0 190 0 1 2170
box -6 -8 86 248
use NAND3X1  _3114_
timestamp 0
transform -1 0 4710 0 1 1210
box -6 -8 106 248
use AND2X2  _3115_
timestamp 0
transform -1 0 4770 0 -1 1690
box -6 -8 106 248
use AND2X2  _3116_
timestamp 0
transform 1 0 4550 0 -1 1210
box -6 -8 106 248
use OAI22X1  _3117_
timestamp 0
transform 1 0 590 0 1 1210
box -6 -8 126 248
use NAND3X1  _3118_
timestamp 0
transform -1 0 1830 0 1 1210
box -6 -8 106 248
use NOR2X1  _3119_
timestamp 0
transform 1 0 910 0 -1 1690
box -6 -8 86 248
use NAND2X1  _3120_
timestamp 0
transform 1 0 1090 0 -1 1690
box -6 -8 86 248
use NOR2X1  _3121_
timestamp 0
transform -1 0 2470 0 -1 1690
box -6 -8 86 248
use NOR2X1  _3122_
timestamp 0
transform -1 0 570 0 1 1690
box -6 -8 86 248
use NAND3X1  _3123_
timestamp 0
transform 1 0 390 0 -1 2170
box -6 -8 106 248
use INVX1  _3124_
timestamp 0
transform 1 0 290 0 1 2170
box -6 -8 66 248
use AND2X2  _3125_
timestamp 0
transform 1 0 2110 0 1 1210
box -6 -8 106 248
use NOR2X1  _3126_
timestamp 0
transform -1 0 2390 0 1 1210
box -6 -8 86 248
use AND2X2  _3127_
timestamp 0
transform 1 0 1630 0 -1 1690
box -6 -8 106 248
use INVX1  _3128_
timestamp 0
transform 1 0 1470 0 -1 1690
box -6 -8 66 248
use NOR2X1  _3129_
timestamp 0
transform 1 0 4810 0 1 1210
box -6 -8 86 248
use NAND3X1  _3130_
timestamp 0
transform 1 0 4990 0 1 1210
box -6 -8 106 248
use NOR2X1  _3131_
timestamp 0
transform 1 0 5210 0 -1 1210
box -6 -8 86 248
use INVX1  _3132_
timestamp 0
transform 1 0 4870 0 -1 1690
box -6 -8 66 248
use NAND2X1  _3133_
timestamp 0
transform -1 0 4830 0 -1 1210
box -6 -8 86 248
use INVX1  _3134_
timestamp 0
transform -1 0 4450 0 -1 1210
box -6 -8 66 248
use INVX1  _3135_
timestamp 0
transform 1 0 770 0 -1 1690
box -6 -8 66 248
use INVX1  _3136_
timestamp 0
transform -1 0 870 0 1 1210
box -6 -8 66 248
use OAI21X1  _3137_
timestamp 0
transform 1 0 430 0 -1 250
box -6 -8 106 248
use OAI21X1  _3138_
timestamp 0
transform 1 0 770 0 1 250
box -6 -8 106 248
use INVX1  _3139_
timestamp 0
transform 1 0 270 0 -1 250
box -6 -8 66 248
use OAI21X1  _3140_
timestamp 0
transform -1 0 1670 0 1 730
box -6 -8 106 248
use OAI21X1  _3141_
timestamp 0
transform 1 0 1770 0 1 730
box -6 -8 106 248
use INVX1  _3142_
timestamp 0
transform -1 0 1790 0 1 250
box -6 -8 66 248
use OAI21X1  _3143_
timestamp 0
transform 1 0 2450 0 -1 250
box -6 -8 106 248
use OAI21X1  _3144_
timestamp 0
transform 1 0 2570 0 1 250
box -6 -8 106 248
use INVX1  _3145_
timestamp 0
transform 1 0 2290 0 -1 250
box -6 -8 66 248
use OAI21X1  _3146_
timestamp 0
transform -1 0 2070 0 1 730
box -6 -8 106 248
use OAI21X1  _3147_
timestamp 0
transform 1 0 2090 0 -1 1210
box -6 -8 106 248
use INVX2  _3148_
timestamp 0
transform 1 0 1130 0 -1 730
box -6 -8 66 248
use NOR2X1  _3149_
timestamp 0
transform -1 0 1030 0 -1 730
box -6 -8 86 248
use INVX4  _3150_
timestamp 0
transform -1 0 390 0 -1 1210
box -6 -8 86 248
use INVX4  _3151_
timestamp 0
transform 1 0 110 0 1 250
box -6 -8 86 248
use INVX1  _3152_
timestamp 0
transform -1 0 2230 0 1 730
box -6 -8 66 248
use DFFSR  _3153_
timestamp 0
transform 1 0 2870 0 -1 6010
box -6 -8 486 248
use DFFSR  _3154_
timestamp 0
transform 1 0 1710 0 -1 4570
box -6 -8 486 248
use DFFSR  _3155_
timestamp 0
transform 1 0 2250 0 -1 5530
box -6 -8 486 248
use DFFSR  _3156_
timestamp 0
transform -1 0 3550 0 1 7930
box -6 -8 486 248
use DFFSR  _3157_
timestamp 0
transform 1 0 2390 0 1 6010
box -6 -8 486 248
use DFFSR  _3158_
timestamp 0
transform 1 0 5490 0 -1 10330
box -6 -8 486 248
use DFFSR  _3159_
timestamp 0
transform -1 0 5690 0 -1 8410
box -6 -8 486 248
use DFFSR  _3160_
timestamp 0
transform 1 0 4630 0 -1 10330
box -6 -8 486 248
use DFFSR  _3161_
timestamp 0
transform 1 0 4090 0 -1 9370
box -6 -8 486 248
use DFFSR  _3162_
timestamp 0
transform 1 0 550 0 1 4090
box -6 -8 486 248
use DFFSR  _3163_
timestamp 0
transform 1 0 3130 0 1 9850
box -6 -8 486 248
use DFFSR  _3164_
timestamp 0
transform 1 0 4730 0 -1 8410
box -6 -8 486 248
use DFFSR  _3165_
timestamp 0
transform 1 0 3830 0 -1 9850
box -6 -8 486 248
use DFFSR  _3166_
timestamp 0
transform -1 0 4750 0 1 3610
box -6 -8 486 248
use DFFSR  _3167_
timestamp 0
transform 1 0 570 0 -1 3130
box -6 -8 486 248
use DFFSR  _3168_
timestamp 0
transform 1 0 3790 0 1 9850
box -6 -8 486 248
use DFFSR  _3169_
timestamp 0
transform -1 0 3170 0 -1 9850
box -6 -8 486 248
use DFFSR  _3170_
timestamp 0
transform -1 0 4170 0 -1 4090
box -6 -8 486 248
use DFFPOSX1  _3171_
timestamp 0
transform 1 0 550 0 -1 11770
box -6 -8 246 248
use DFFPOSX1  _3172_
timestamp 0
transform 1 0 10 0 1 11290
box -6 -8 246 248
use DFFPOSX1  _3173_
timestamp 0
transform 1 0 1510 0 1 9370
box -6 -8 246 248
use DFFPOSX1  _3174_
timestamp 0
transform 1 0 10 0 -1 11290
box -6 -8 246 248
use DFFSR  _3175_
timestamp 0
transform 1 0 10 0 -1 3610
box -6 -8 486 248
use DFFSR  _3176_
timestamp 0
transform 1 0 4510 0 -1 9850
box -6 -8 486 248
use DFFPOSX1  _3177_
timestamp 0
transform 1 0 10 0 -1 11770
box -6 -8 246 248
use DFFSR  _3178_
timestamp 0
transform -1 0 7770 0 -1 3610
box -6 -8 486 248
use DFFSR  _3179_
timestamp 0
transform 1 0 1150 0 1 3130
box -6 -8 486 248
use DFFSR  _3180_
timestamp 0
transform 1 0 6310 0 1 10810
box -6 -8 486 248
use DFFSR  _3181_
timestamp 0
transform 1 0 2210 0 -1 9850
box -6 -8 486 248
use DFFSR  _3182_
timestamp 0
transform -1 0 7090 0 1 3610
box -6 -8 486 248
use DFFSR  _3183_
timestamp 0
transform 1 0 1030 0 -1 5530
box -6 -8 486 248
use DFFSR  _3184_
timestamp 0
transform 1 0 3270 0 -1 5530
box -6 -8 486 248
use DFFSR  _3185_
timestamp 0
transform -1 0 8590 0 -1 6010
box -6 -8 486 248
use DFFSR  _3186_
timestamp 0
transform 1 0 2970 0 -1 9370
box -6 -8 486 248
use DFFSR  _3187_
timestamp 0
transform -1 0 4930 0 1 7930
box -6 -8 486 248
use DFFSR  _3188_
timestamp 0
transform -1 0 2970 0 -1 9370
box -6 -8 486 248
use DFFSR  _3189_
timestamp 0
transform 1 0 1510 0 1 4570
box -6 -8 486 248
use DFFSR  _3190_
timestamp 0
transform 1 0 490 0 1 6010
box -6 -8 486 248
use DFFSR  _3191_
timestamp 0
transform 1 0 5290 0 1 3130
box -6 -8 486 248
use DFFSR  _3192_
timestamp 0
transform 1 0 11530 0 -1 11770
box -6 -8 486 248
use DFFSR  _3193_
timestamp 0
transform 1 0 6630 0 -1 10810
box -6 -8 486 248
use DFFSR  _3194_
timestamp 0
transform -1 0 5670 0 -1 9850
box -6 -8 486 248
use DFFSR  _3195_
timestamp 0
transform 1 0 4290 0 -1 8890
box -6 -8 486 248
use DFFSR  _3196_
timestamp 0
transform -1 0 2850 0 1 3130
box -6 -8 486 248
use DFFSR  _3197_
timestamp 0
transform -1 0 6650 0 -1 7450
box -6 -8 486 248
use DFFSR  _3198_
timestamp 0
transform 1 0 4810 0 1 3130
box -6 -8 486 248
use DFFSR  _3199_
timestamp 0
transform 1 0 3170 0 -1 9850
box -6 -8 486 248
use DFFSR  _3200_
timestamp 0
transform -1 0 5570 0 1 3610
box -6 -8 486 248
use DFFSR  _3201_
timestamp 0
transform 1 0 1070 0 1 2650
box -6 -8 486 248
use DFFSR  _3202_
timestamp 0
transform -1 0 8030 0 1 4570
box -6 -8 486 248
use DFFSR  _3203_
timestamp 0
transform 1 0 1970 0 -1 10330
box -6 -8 486 248
use DFFSR  _3204_
timestamp 0
transform -1 0 5070 0 1 4090
box -6 -8 486 248
use DFFSR  _3205_
timestamp 0
transform 1 0 3550 0 1 9370
box -6 -8 486 248
use DFFSR  _3206_
timestamp 0
transform 1 0 3570 0 -1 3610
box -6 -8 486 248
use DFFSR  _3207_
timestamp 0
transform 1 0 3150 0 1 4570
box -6 -8 486 248
use DFFSR  _3208_
timestamp 0
transform 1 0 5970 0 -1 10330
box -6 -8 486 248
use DFFPOSX1  _3209_
timestamp 0
transform 1 0 1030 0 -1 9850
box -6 -8 246 248
use DFFPOSX1  _3210_
timestamp 0
transform 1 0 490 0 -1 10810
box -6 -8 246 248
use DFFSR  _3211_
timestamp 0
transform 1 0 11650 0 1 10810
box -6 -8 486 248
use DFFSR  _3212_
timestamp 0
transform 1 0 10 0 1 3130
box -6 -8 486 248
use DFFSR  _3213_
timestamp 0
transform 1 0 10 0 -1 10810
box -6 -8 486 248
use DFFSR  _3214_
timestamp 0
transform 1 0 9470 0 1 11770
box -6 -8 486 248
use DFFSR  _3215_
timestamp 0
transform 1 0 5010 0 1 9850
box -6 -8 486 248
use DFFSR  _3216_
timestamp 0
transform -1 0 1570 0 1 10330
box -6 -8 486 248
use DFFSR  _3217_
timestamp 0
transform 1 0 4790 0 -1 10810
box -6 -8 486 248
use DFFSR  _3218_
timestamp 0
transform 1 0 6690 0 1 9850
box -6 -8 486 248
use DFFSR  _3219_
timestamp 0
transform 1 0 3450 0 -1 9370
box -6 -8 486 248
use DFFSR  _3220_
timestamp 0
transform 1 0 11690 0 -1 11290
box -6 -8 486 248
use DFFSR  _3221_
timestamp 0
transform 1 0 7110 0 -1 10810
box -6 -8 486 248
use DFFSR  _3222_
timestamp 0
transform 1 0 9950 0 1 11770
box -6 -8 486 248
use DFFSR  _3223_
timestamp 0
transform 1 0 7590 0 1 10810
box -6 -8 486 248
use DFFSR  _3224_
timestamp 0
transform 1 0 8130 0 1 6970
box -6 -8 486 248
use DFFSR  _3225_
timestamp 0
transform -1 0 6490 0 1 9850
box -6 -8 486 248
use DFFSR  _3226_
timestamp 0
transform 1 0 1810 0 -1 6490
box -6 -8 486 248
use DFFSR  _3227_
timestamp 0
transform -1 0 490 0 1 6010
box -6 -8 486 248
use DFFSR  _3228_
timestamp 0
transform 1 0 710 0 -1 6490
box -6 -8 486 248
use DFFSR  _3229_
timestamp 0
transform 1 0 1310 0 -1 7450
box -6 -8 486 248
use DFFSR  _3230_
timestamp 0
transform 1 0 490 0 -1 4090
box -6 -8 486 248
use DFFSR  _3231_
timestamp 0
transform 1 0 630 0 -1 7450
box -6 -8 486 248
use DFFSR  _3232_
timestamp 0
transform -1 0 8210 0 1 4090
box -6 -8 486 248
use DFFSR  _3233_
timestamp 0
transform 1 0 5370 0 1 10330
box -6 -8 486 248
use DFFSR  _3234_
timestamp 0
transform 1 0 190 0 1 9370
box -6 -8 486 248
use DFFSR  _3235_
timestamp 0
transform -1 0 3670 0 -1 4570
box -6 -8 486 248
use DFFSR  _3236_
timestamp 0
transform 1 0 6390 0 -1 11290
box -6 -8 486 248
use DFFSR  _3237_
timestamp 0
transform 1 0 10 0 -1 10330
box -6 -8 486 248
use DFFSR  _3238_
timestamp 0
transform 1 0 1030 0 1 9370
box -6 -8 486 248
use DFFSR  _3239_
timestamp 0
transform 1 0 1970 0 -1 4090
box -6 -8 486 248
use DFFSR  _3240_
timestamp 0
transform 1 0 370 0 1 7930
box -6 -8 486 248
use DFFSR  _3241_
timestamp 0
transform -1 0 6190 0 -1 7930
box -6 -8 486 248
use DFFSR  _3242_
timestamp 0
transform 1 0 10 0 1 9850
box -6 -8 486 248
use DFFSR  _3243_
timestamp 0
transform -1 0 3370 0 1 6490
box -6 -8 486 248
use DFFSR  _3244_
timestamp 0
transform 1 0 970 0 1 7450
box -6 -8 486 248
use DFFSR  _3245_
timestamp 0
transform -1 0 7070 0 -1 3610
box -6 -8 486 248
use DFFSR  _3246_
timestamp 0
transform 1 0 690 0 -1 7930
box -6 -8 486 248
use DFFSR  _3247_
timestamp 0
transform 1 0 1190 0 -1 2650
box -6 -8 486 248
use DFFSR  _3248_
timestamp 0
transform 1 0 1810 0 1 8890
box -6 -8 486 248
use DFFSR  _3249_
timestamp 0
transform -1 0 3870 0 -1 7930
box -6 -8 486 248
use DFFSR  _3250_
timestamp 0
transform 1 0 1950 0 -1 7450
box -6 -8 486 248
use DFFSR  _3251_
timestamp 0
transform 1 0 4170 0 -1 4090
box -6 -8 486 248
use DFFSR  _3252_
timestamp 0
transform 1 0 1150 0 1 6010
box -6 -8 486 248
use DFFSR  _3253_
timestamp 0
transform 1 0 590 0 1 2650
box -6 -8 486 248
use DFFSR  _3254_
timestamp 0
transform 1 0 1850 0 -1 6010
box -6 -8 486 248
use DFFSR  _3255_
timestamp 0
transform -1 0 4590 0 1 3130
box -6 -8 486 248
use DFFSR  _3256_
timestamp 0
transform 1 0 2450 0 -1 10330
box -6 -8 486 248
use DFFSR  _3257_
timestamp 0
transform 1 0 990 0 1 3610
box -6 -8 486 248
use DFFSR  _3258_
timestamp 0
transform -1 0 6670 0 1 7450
box -6 -8 486 248
use DFFSR  _3259_
timestamp 0
transform 1 0 730 0 1 5050
box -6 -8 486 248
use DFFSR  _3260_
timestamp 0
transform 1 0 1030 0 -1 6010
box -6 -8 486 248
use DFFSR  _3261_
timestamp 0
transform 1 0 1790 0 1 4090
box -6 -8 486 248
use DFFSR  _3262_
timestamp 0
transform -1 0 7530 0 1 6970
box -6 -8 486 248
use DFFSR  _3263_
timestamp 0
transform 1 0 2070 0 -1 5050
box -6 -8 486 248
use DFFSR  _3264_
timestamp 0
transform 1 0 1030 0 -1 4570
box -6 -8 486 248
use DFFSR  _3265_
timestamp 0
transform 1 0 1350 0 1 5530
box -6 -8 486 248
use DFFSR  _3266_
timestamp 0
transform 1 0 2650 0 1 9850
box -6 -8 486 248
use DFFSR  _3267_
timestamp 0
transform -1 0 490 0 -1 5530
box -6 -8 486 248
use DFFSR  _3268_
timestamp 0
transform 1 0 2830 0 -1 4090
box -6 -8 486 248
use DFFSR  _3269_
timestamp 0
transform 1 0 3730 0 1 10330
box -6 -8 486 248
use DFFSR  _3270_
timestamp 0
transform 1 0 490 0 1 3130
box -6 -8 486 248
use DFFSR  _3271_
timestamp 0
transform 1 0 4230 0 -1 4570
box -6 -8 486 248
use DFFSR  _3272_
timestamp 0
transform 1 0 310 0 1 5530
box -6 -8 486 248
use DFFSR  _3273_
timestamp 0
transform 1 0 10 0 -1 4090
box -6 -8 486 248
use DFFSR  _3274_
timestamp 0
transform 1 0 7110 0 -1 11770
box -6 -8 486 248
use DFFPOSX1  _3275_
timestamp 0
transform -1 0 830 0 -1 9850
box -6 -8 246 248
use DFFSR  _3276_
timestamp 0
transform 1 0 10 0 -1 4570
box -6 -8 486 248
use DFFSR  _3277_
timestamp 0
transform 1 0 1270 0 -1 3610
box -6 -8 486 248
use DFFSR  _3278_
timestamp 0
transform 1 0 1830 0 -1 3130
box -6 -8 486 248
use DFFSR  _3279_
timestamp 0
transform 1 0 5810 0 -1 10810
box -6 -8 486 248
use DFFSR  _3280_
timestamp 0
transform -1 0 7550 0 1 4570
box -6 -8 486 248
use DFFSR  _3281_
timestamp 0
transform -1 0 3170 0 1 3610
box -6 -8 486 248
use DFFSR  _3282_
timestamp 0
transform 1 0 410 0 1 10330
box -6 -8 486 248
use DFFSR  _3283_
timestamp 0
transform -1 0 11510 0 -1 11290
box -6 -8 486 248
use OAI21X1  _3284_
timestamp 0
transform -1 0 4870 0 1 4570
box -6 -8 106 248
use NAND2X1  _3285_
timestamp 0
transform 1 0 4430 0 1 4570
box -6 -8 86 248
use OAI21X1  _3286_
timestamp 0
transform -1 0 3550 0 -1 6010
box -6 -8 106 248
use NAND2X1  _3287_
timestamp 0
transform 1 0 3330 0 1 5530
box -6 -8 86 248
use OAI21X1  _3288_
timestamp 0
transform 1 0 2250 0 1 5530
box -6 -8 106 248
use NAND2X1  _3289_
timestamp 0
transform 1 0 2450 0 1 5530
box -6 -8 86 248
use INVX1  _3290_
timestamp 0
transform -1 0 2150 0 1 5530
box -6 -8 66 248
use OAI21X1  _3291_
timestamp 0
transform 1 0 3070 0 -1 6490
box -6 -8 106 248
use NAND2X1  _3292_
timestamp 0
transform 1 0 3270 0 -1 6490
box -6 -8 86 248
use AOI22X1  _3293_
timestamp 0
transform 1 0 5890 0 1 8410
box -6 -8 126 248
use OAI21X1  _3294_
timestamp 0
transform -1 0 6010 0 -1 8890
box -6 -8 106 248
use NAND2X1  _3295_
timestamp 0
transform 1 0 5970 0 1 9370
box -6 -8 86 248
use OAI21X1  _3296_
timestamp 0
transform 1 0 6450 0 1 8410
box -6 -8 106 248
use OAI21X1  _3297_
timestamp 0
transform 1 0 6650 0 1 8410
box -6 -8 106 248
use OAI21X1  _3298_
timestamp 0
transform 1 0 5350 0 -1 8890
box -6 -8 106 248
use NAND2X1  _3299_
timestamp 0
transform 1 0 5550 0 1 8410
box -6 -8 86 248
use OAI21X1  _3300_
timestamp 0
transform 1 0 4690 0 1 9370
box -6 -8 106 248
use NAND2X1  _3301_
timestamp 0
transform 1 0 4890 0 1 9370
box -6 -8 86 248
use OAI21X1  _3302_
timestamp 0
transform -1 0 3530 0 1 10330
box -6 -8 106 248
use OAI21X1  _3303_
timestamp 0
transform -1 0 3690 0 -1 10330
box -6 -8 106 248
use AND2X2  _3304_
timestamp 0
transform -1 0 3570 0 1 10810
box -6 -8 106 248
use NAND3X1  _3305_
timestamp 0
transform -1 0 3750 0 -1 11290
box -6 -8 106 248
use OAI21X1  _3306_
timestamp 0
transform 1 0 4410 0 -1 9850
box -6 -8 106 248
use NAND2X1  _3307_
timestamp 0
transform 1 0 4510 0 1 9370
box -6 -8 86 248
use OAI21X1  _3308_
timestamp 0
transform -1 0 1250 0 -1 3130
box -6 -8 106 248
use NAND2X1  _3309_
timestamp 0
transform -1 0 1150 0 1 3130
box -6 -8 86 248
use OAI21X1  _3310_
timestamp 0
transform 1 0 2550 0 1 9850
box -6 -8 106 248
use OAI21X1  _3311_
timestamp 0
transform -1 0 2870 0 -1 10810
box -6 -8 106 248
use OAI21X1  _3312_
timestamp 0
transform 1 0 3510 0 1 11290
box -6 -8 106 248
use INVX1  _3313_
timestamp 0
transform -1 0 2470 0 1 9850
box -6 -8 66 248
use OAI21X1  _3314_
timestamp 0
transform -1 0 390 0 1 3610
box -6 -8 106 248
use OAI21X1  _3315_
timestamp 0
transform -1 0 590 0 1 3610
box -6 -8 106 248
use MUX2X1  _3316_
timestamp 0
transform -1 0 7690 0 -1 4090
box -6 -8 126 248
use OAI21X1  _3317_
timestamp 0
transform 1 0 6210 0 1 10810
box -6 -8 106 248
use OAI21X1  _3318_
timestamp 0
transform 1 0 2690 0 1 10810
box -6 -8 106 248
use OAI21X1  _3319_
timestamp 0
transform 1 0 6710 0 1 10330
box -6 -8 106 248
use INVX1  _3320_
timestamp 0
transform 1 0 5490 0 1 10810
box -6 -8 66 248
use MUX2X1  _3321_
timestamp 0
transform -1 0 6610 0 1 3610
box -6 -8 126 248
use AOI21X1  _3322_
timestamp 0
transform -1 0 3950 0 -1 5530
box -6 -8 106 248
use NOR2X1  _3323_
timestamp 0
transform -1 0 3770 0 1 5530
box -6 -8 86 248
use OAI21X1  _3324_
timestamp 0
transform 1 0 5210 0 1 7930
box -6 -8 106 248
use NAND3X1  _3325_
timestamp 0
transform -1 0 5510 0 1 7930
box -6 -8 106 248
use OAI21X1  _3326_
timestamp 0
transform -1 0 5370 0 -1 7930
box -6 -8 106 248
use OAI21X1  _3327_
timestamp 0
transform 1 0 4870 0 -1 7930
box -6 -8 106 248
use MUX2X1  _3328_
timestamp 0
transform -1 0 5430 0 1 7450
box -6 -8 126 248
use NOR2X1  _3329_
timestamp 0
transform -1 0 5810 0 -1 7450
box -6 -8 86 248
use AND2X2  _3330_
timestamp 0
transform 1 0 5590 0 1 7930
box -6 -8 106 248
use NAND2X1  _3331_
timestamp 0
transform 1 0 5030 0 1 7930
box -6 -8 86 248
use NOR2X1  _3332_
timestamp 0
transform -1 0 4770 0 -1 7930
box -6 -8 86 248
use OAI21X1  _3333_
timestamp 0
transform -1 0 6090 0 1 7930
box -6 -8 106 248
use INVX1  _3334_
timestamp 0
transform 1 0 5990 0 -1 8410
box -6 -8 66 248
use OAI21X1  _3335_
timestamp 0
transform -1 0 590 0 1 10810
box -6 -8 106 248
use NAND2X1  _3336_
timestamp 0
transform -1 0 390 0 1 10810
box -6 -8 86 248
use OAI21X1  _3337_
timestamp 0
transform -1 0 1030 0 1 9850
box -6 -8 106 248
use NAND2X1  _3338_
timestamp 0
transform -1 0 1030 0 -1 10330
box -6 -8 86 248
use AOI21X1  _3339_
timestamp 0
transform -1 0 6010 0 -1 3610
box -6 -8 106 248
use NOR2X1  _3340_
timestamp 0
transform 1 0 6110 0 -1 3610
box -6 -8 86 248
use OAI22X1  _3341_
timestamp 0
transform -1 0 5990 0 -1 11290
box -6 -8 126 248
use OAI21X1  _3342_
timestamp 0
transform -1 0 5590 0 -1 11290
box -6 -8 106 248
use OAI21X1  _3343_
timestamp 0
transform -1 0 4510 0 1 8890
box -6 -8 106 248
use AOI21X1  _3344_
timestamp 0
transform -1 0 5630 0 -1 3610
box -6 -8 106 248
use NOR2X1  _3345_
timestamp 0
transform 1 0 5730 0 -1 3610
box -6 -8 86 248
use AOI21X1  _3346_
timestamp 0
transform 1 0 5330 0 -1 3610
box -6 -8 106 248
use NOR2X1  _3347_
timestamp 0
transform 1 0 5150 0 -1 3610
box -6 -8 86 248
use AOI21X1  _3348_
timestamp 0
transform -1 0 210 0 1 11770
box -6 -8 106 248
use NOR2X1  _3349_
timestamp 0
transform 1 0 310 0 1 11770
box -6 -8 86 248
use MUX2X1  _3350_
timestamp 0
transform 1 0 7810 0 -1 4570
box -6 -8 126 248
use AOI21X1  _3351_
timestamp 0
transform -1 0 210 0 1 10810
box -6 -8 106 248
use NOR2X1  _3352_
timestamp 0
transform 1 0 350 0 -1 11290
box -6 -8 86 248
use AOI21X1  _3353_
timestamp 0
transform -1 0 1950 0 1 9370
box -6 -8 106 248
use NOR2X1  _3354_
timestamp 0
transform 1 0 2050 0 1 9370
box -6 -8 86 248
use AOI21X1  _3355_
timestamp 0
transform -1 0 450 0 1 11290
box -6 -8 106 248
use NOR2X1  _3356_
timestamp 0
transform -1 0 630 0 1 11290
box -6 -8 86 248
use AOI21X1  _3357_
timestamp 0
transform -1 0 990 0 -1 11770
box -6 -8 106 248
use NOR2X1  _3358_
timestamp 0
transform -1 0 950 0 1 11770
box -6 -8 86 248
use AOI21X1  _3359_
timestamp 0
transform -1 0 210 0 -1 3130
box -6 -8 106 248
use NOR2X1  _3360_
timestamp 0
transform -1 0 390 0 -1 3130
box -6 -8 86 248
use OAI21X1  _3361_
timestamp 0
transform -1 0 5010 0 1 9850
box -6 -8 106 248
use OAI22X1  _3362_
timestamp 0
transform -1 0 5150 0 1 10330
box -6 -8 126 248
use INVX1  _3363_
timestamp 0
transform 1 0 5370 0 -1 10810
box -6 -8 66 248
use OAI21X1  _3364_
timestamp 0
transform -1 0 3550 0 1 9370
box -6 -8 106 248
use OAI21X1  _3365_
timestamp 0
transform 1 0 3390 0 -1 10810
box -6 -8 106 248
use NAND3X1  _3366_
timestamp 0
transform 1 0 2970 0 -1 10810
box -6 -8 106 248
use AOI22X1  _3367_
timestamp 0
transform 1 0 2610 0 -1 11770
box -6 -8 126 248
use OAI21X1  _3368_
timestamp 0
transform 1 0 2410 0 -1 11770
box -6 -8 106 248
use NAND2X1  _3369_
timestamp 0
transform -1 0 4250 0 -1 10810
box -6 -8 86 248
use NOR2X1  _3370_
timestamp 0
transform -1 0 5390 0 1 10810
box -6 -8 86 248
use AOI22X1  _3371_
timestamp 0
transform -1 0 7210 0 1 10810
box -6 -8 126 248
use NOR2X1  _3372_
timestamp 0
transform 1 0 5150 0 1 10810
box -6 -8 86 248
use INVX1  _3373_
timestamp 0
transform -1 0 7590 0 1 10810
box -6 -8 66 248
use AOI22X1  _3374_
timestamp 0
transform -1 0 7430 0 1 10810
box -6 -8 126 248
use NOR2X1  _3375_
timestamp 0
transform -1 0 4790 0 -1 10810
box -6 -8 86 248
use OR2X2  _3376_
timestamp 0
transform -1 0 4850 0 1 10810
box -6 -8 106 248
use OAI21X1  _3377_
timestamp 0
transform 1 0 4950 0 1 10810
box -6 -8 106 248
use NOR2X1  _3378_
timestamp 0
transform -1 0 4430 0 -1 10810
box -6 -8 86 248
use OR2X2  _3379_
timestamp 0
transform 1 0 5810 0 1 10810
box -6 -8 106 248
use INVX1  _3380_
timestamp 0
transform -1 0 7910 0 -1 10810
box -6 -8 66 248
use OAI21X1  _3381_
timestamp 0
transform 1 0 6710 0 1 9370
box -6 -8 106 248
use NAND2X1  _3382_
timestamp 0
transform 1 0 6530 0 1 9370
box -6 -8 86 248
use AOI21X1  _3383_
timestamp 0
transform -1 0 7210 0 1 9370
box -6 -8 106 248
use OAI21X1  _3384_
timestamp 0
transform -1 0 7010 0 1 9370
box -6 -8 106 248
use OAI21X1  _3385_
timestamp 0
transform 1 0 7310 0 1 9370
box -6 -8 106 248
use OAI22X1  _3386_
timestamp 0
transform -1 0 6670 0 -1 9850
box -6 -8 126 248
use OAI21X1  _3387_
timestamp 0
transform 1 0 6350 0 -1 9850
box -6 -8 106 248
use OAI21X1  _3388_
timestamp 0
transform 1 0 6770 0 -1 9850
box -6 -8 106 248
use INVX1  _3389_
timestamp 0
transform -1 0 7210 0 -1 9850
box -6 -8 66 248
use NOR2X1  _3390_
timestamp 0
transform -1 0 9810 0 -1 9850
box -6 -8 86 248
use OAI21X1  _3391_
timestamp 0
transform -1 0 10390 0 -1 9850
box -6 -8 106 248
use OAI21X1  _3392_
timestamp 0
transform -1 0 390 0 -1 6010
box -6 -8 106 248
use AND2X2  _3393_
timestamp 0
transform 1 0 290 0 -1 6490
box -6 -8 106 248
use OAI21X1  _3394_
timestamp 0
transform -1 0 370 0 1 6970
box -6 -8 106 248
use NAND3X1  _3395_
timestamp 0
transform -1 0 390 0 -1 6970
box -6 -8 106 248
use NAND2X1  _3396_
timestamp 0
transform -1 0 190 0 -1 6010
box -6 -8 86 248
use OAI21X1  _3397_
timestamp 0
transform -1 0 1370 0 1 6970
box -6 -8 106 248
use OAI21X1  _3398_
timestamp 0
transform 1 0 1070 0 1 6970
box -6 -8 106 248
use AOI21X1  _3399_
timestamp 0
transform 1 0 1030 0 -1 6970
box -6 -8 106 248
use NOR3X1  _3400_
timestamp 0
transform -1 0 830 0 1 6970
box -6 -8 186 248
use NAND3X1  _3401_
timestamp 0
transform -1 0 210 0 1 7930
box -6 -8 106 248
use INVX1  _3402_
timestamp 0
transform -1 0 930 0 -1 6970
box -6 -8 66 248
use NOR2X1  _3403_
timestamp 0
transform 1 0 1650 0 1 6970
box -6 -8 86 248
use AOI21X1  _3404_
timestamp 0
transform -1 0 1030 0 -1 9850
box -6 -8 106 248
use NOR2X1  _3405_
timestamp 0
transform 1 0 750 0 1 9850
box -6 -8 86 248
use NOR2X1  _3406_
timestamp 0
transform -1 0 1990 0 -1 9850
box -6 -8 86 248
use OAI22X1  _3407_
timestamp 0
transform -1 0 630 0 -1 7450
box -6 -8 126 248
use OAI21X1  _3408_
timestamp 0
transform 1 0 310 0 -1 7450
box -6 -8 106 248
use AND2X2  _3409_
timestamp 0
transform -1 0 210 0 -1 7450
box -6 -8 106 248
use INVX1  _3410_
timestamp 0
transform -1 0 970 0 1 6970
box -6 -8 66 248
use OAI21X1  _3411_
timestamp 0
transform -1 0 570 0 -1 9370
box -6 -8 106 248
use NAND2X1  _3412_
timestamp 0
transform -1 0 370 0 -1 9370
box -6 -8 86 248
use NAND2X1  _3413_
timestamp 0
transform -1 0 190 0 -1 9370
box -6 -8 86 248
use NAND3X1  _3414_
timestamp 0
transform -1 0 370 0 -1 8890
box -6 -8 106 248
use INVX1  _3415_
timestamp 0
transform -1 0 170 0 -1 8890
box -6 -8 66 248
use OAI21X1  _3416_
timestamp 0
transform -1 0 210 0 1 8890
box -6 -8 106 248
use OAI21X1  _3417_
timestamp 0
transform -1 0 550 0 1 8410
box -6 -8 106 248
use OAI21X1  _3418_
timestamp 0
transform -1 0 7070 0 -1 11290
box -6 -8 106 248
use OAI21X1  _3419_
timestamp 0
transform 1 0 6290 0 -1 11290
box -6 -8 106 248
use OAI21X1  _3420_
timestamp 0
transform 1 0 6090 0 -1 11290
box -6 -8 106 248
use INVX1  _3421_
timestamp 0
transform 1 0 5330 0 -1 11290
box -6 -8 66 248
use NOR2X1  _3422_
timestamp 0
transform 1 0 5190 0 1 11290
box -6 -8 86 248
use INVX1  _3423_
timestamp 0
transform 1 0 7170 0 -1 11290
box -6 -8 66 248
use OAI21X1  _3424_
timestamp 0
transform -1 0 1510 0 -1 9370
box -6 -8 106 248
use OAI21X1  _3425_
timestamp 0
transform 1 0 670 0 -1 9370
box -6 -8 106 248
use NOR2X1  _3426_
timestamp 0
transform 1 0 470 0 1 8890
box -6 -8 86 248
use NOR3X1  _3427_
timestamp 0
transform -1 0 650 0 -1 8890
box -6 -8 186 248
use INVX1  _3428_
timestamp 0
transform -1 0 370 0 1 8890
box -6 -8 66 248
use NOR2X1  _3429_
timestamp 0
transform 1 0 650 0 1 8890
box -6 -8 86 248
use NAND3X1  _3430_
timestamp 0
transform -1 0 190 0 1 8410
box -6 -8 106 248
use INVX1  _3431_
timestamp 0
transform -1 0 350 0 1 8410
box -6 -8 66 248
use OAI21X1  _3432_
timestamp 0
transform 1 0 930 0 -1 8890
box -6 -8 106 248
use OAI21X1  _3433_
timestamp 0
transform 1 0 1530 0 -1 8890
box -6 -8 106 248
use OAI21X1  _3434_
timestamp 0
transform -1 0 1110 0 1 8410
box -6 -8 106 248
use OAI21X1  _3435_
timestamp 0
transform -1 0 1230 0 -1 8890
box -6 -8 106 248
use AOI21X1  _3436_
timestamp 0
transform 1 0 1330 0 -1 8890
box -6 -8 106 248
use AND2X2  _3437_
timestamp 0
transform -1 0 1450 0 -1 8410
box -6 -8 106 248
use NOR2X1  _3438_
timestamp 0
transform -1 0 1110 0 1 8890
box -6 -8 86 248
use OAI21X1  _3439_
timestamp 0
transform -1 0 930 0 1 8890
box -6 -8 106 248
use OAI21X1  _3440_
timestamp 0
transform -1 0 1250 0 -1 8410
box -6 -8 106 248
use OAI21X1  _3441_
timestamp 0
transform 1 0 770 0 1 9370
box -6 -8 106 248
use OAI21X1  _3442_
timestamp 0
transform 1 0 870 0 -1 9370
box -6 -8 106 248
use NOR2X1  _3443_
timestamp 0
transform -1 0 910 0 1 8410
box -6 -8 86 248
use NAND2X1  _3444_
timestamp 0
transform -1 0 730 0 1 8410
box -6 -8 86 248
use AND2X2  _3445_
timestamp 0
transform -1 0 870 0 -1 8410
box -6 -8 106 248
use OAI21X1  _3446_
timestamp 0
transform -1 0 1530 0 1 8410
box -6 -8 106 248
use NOR2X1  _3447_
timestamp 0
transform -1 0 1290 0 1 8890
box -6 -8 86 248
use NOR2X1  _3448_
timestamp 0
transform -1 0 830 0 -1 8890
box -6 -8 86 248
use NOR2X1  _3449_
timestamp 0
transform 1 0 1390 0 1 8890
box -6 -8 86 248
use NOR2X1  _3450_
timestamp 0
transform 1 0 1550 0 1 8890
box -6 -8 86 248
use NAND3X1  _3451_
timestamp 0
transform -1 0 2770 0 -1 8890
box -6 -8 106 248
use AND2X2  _3452_
timestamp 0
transform -1 0 2970 0 -1 8890
box -6 -8 106 248
use OAI21X1  _3453_
timestamp 0
transform -1 0 3190 0 1 8410
box -6 -8 106 248
use OAI21X1  _3454_
timestamp 0
transform -1 0 1310 0 -1 7450
box -6 -8 106 248
use OAI21X1  _3455_
timestamp 0
transform -1 0 410 0 1 7450
box -6 -8 106 248
use AOI21X1  _3456_
timestamp 0
transform -1 0 210 0 1 7450
box -6 -8 106 248
use OAI21X1  _3457_
timestamp 0
transform -1 0 970 0 1 7450
box -6 -8 106 248
use NAND3X1  _3458_
timestamp 0
transform 1 0 670 0 1 7450
box -6 -8 106 248
use OAI21X1  _3459_
timestamp 0
transform -1 0 690 0 -1 7930
box -6 -8 106 248
use INVX1  _3460_
timestamp 0
transform 1 0 510 0 1 7450
box -6 -8 66 248
use OAI22X1  _3461_
timestamp 0
transform -1 0 2050 0 -1 8890
box -6 -8 126 248
use OAI21X1  _3462_
timestamp 0
transform 1 0 1730 0 -1 8890
box -6 -8 106 248
use AND2X2  _3463_
timestamp 0
transform -1 0 2070 0 -1 8410
box -6 -8 106 248
use OAI22X1  _3464_
timestamp 0
transform -1 0 2210 0 1 7450
box -6 -8 126 248
use NAND2X1  _3465_
timestamp 0
transform -1 0 1750 0 1 7930
box -6 -8 86 248
use OAI21X1  _3466_
timestamp 0
transform -1 0 2150 0 -1 7930
box -6 -8 106 248
use NOR2X1  _3467_
timestamp 0
transform -1 0 1990 0 1 7450
box -6 -8 86 248
use OAI21X1  _3468_
timestamp 0
transform -1 0 2410 0 1 7450
box -6 -8 106 248
use INVX1  _3469_
timestamp 0
transform -1 0 370 0 1 7930
box -6 -8 66 248
use OAI22X1  _3470_
timestamp 0
transform -1 0 1350 0 1 6490
box -6 -8 126 248
use NAND2X1  _3471_
timestamp 0
transform -1 0 1310 0 -1 6970
box -6 -8 86 248
use AOI21X1  _3472_
timestamp 0
transform -1 0 1710 0 1 6490
box -6 -8 106 248
use OAI21X1  _3473_
timestamp 0
transform 1 0 1810 0 1 6490
box -6 -8 106 248
use OAI22X1  _3474_
timestamp 0
transform -1 0 2210 0 1 6010
box -6 -8 126 248
use NAND2X1  _3475_
timestamp 0
transform -1 0 1850 0 -1 6010
box -6 -8 86 248
use NAND2X1  _3476_
timestamp 0
transform -1 0 1810 0 1 6010
box -6 -8 86 248
use NOR2X1  _3477_
timestamp 0
transform -1 0 1990 0 1 6010
box -6 -8 86 248
use OAI21X1  _3478_
timestamp 0
transform 1 0 2010 0 1 6490
box -6 -8 106 248
use INVX1  _3479_
timestamp 0
transform -1 0 1510 0 1 6490
box -6 -8 66 248
use OAI22X1  _3480_
timestamp 0
transform -1 0 2970 0 1 10330
box -6 -8 126 248
use OAI21X1  _3481_
timestamp 0
transform -1 0 6190 0 1 7450
box -6 -8 106 248
use NAND2X1  _3482_
timestamp 0
transform -1 0 5990 0 1 7450
box -6 -8 86 248
use MUX2X1  _3483_
timestamp 0
transform 1 0 6770 0 1 7450
box -6 -8 126 248
use OAI21X1  _3484_
timestamp 0
transform -1 0 7610 0 -1 7450
box -6 -8 106 248
use NAND3X1  _3485_
timestamp 0
transform -1 0 7410 0 -1 7450
box -6 -8 106 248
use OAI21X1  _3486_
timestamp 0
transform 1 0 5790 0 -1 8410
box -6 -8 106 248
use NAND3X1  _3487_
timestamp 0
transform -1 0 5890 0 1 7930
box -6 -8 106 248
use INVX1  _3488_
timestamp 0
transform 1 0 3030 0 -1 10330
box -6 -8 66 248
use OAI21X1  _3489_
timestamp 0
transform -1 0 6250 0 -1 8410
box -6 -8 106 248
use OAI22X1  _3490_
timestamp 0
transform 1 0 1570 0 -1 6970
box -6 -8 126 248
use NAND2X1  _3491_
timestamp 0
transform 1 0 1410 0 -1 6970
box -6 -8 86 248
use NAND2X1  _3492_
timestamp 0
transform 1 0 1970 0 -1 6970
box -6 -8 86 248
use NOR2X1  _3493_
timestamp 0
transform -1 0 1870 0 -1 6970
box -6 -8 86 248
use OAI21X1  _3494_
timestamp 0
transform 1 0 7250 0 -1 6970
box -6 -8 106 248
use NAND3X1  _3495_
timestamp 0
transform -1 0 7710 0 -1 6970
box -6 -8 106 248
use NAND3X1  _3496_
timestamp 0
transform -1 0 7910 0 -1 6970
box -6 -8 106 248
use AND2X2  _3497_
timestamp 0
transform -1 0 8330 0 -1 6970
box -6 -8 106 248
use INVX1  _3498_
timestamp 0
transform -1 0 7510 0 -1 6970
box -6 -8 66 248
use OAI21X1  _3499_
timestamp 0
transform 1 0 1210 0 1 4570
box -6 -8 106 248
use OAI21X1  _3500_
timestamp 0
transform 1 0 1410 0 1 4570
box -6 -8 106 248
use AOI22X1  _3501_
timestamp 0
transform -1 0 3290 0 -1 10810
box -6 -8 126 248
use AOI21X1  _3502_
timestamp 0
transform -1 0 3870 0 -1 10810
box -6 -8 106 248
use NAND3X1  _3503_
timestamp 0
transform -1 0 3370 0 -1 11290
box -6 -8 106 248
use OAI21X1  _3504_
timestamp 0
transform 1 0 2990 0 1 4090
box -6 -8 106 248
use OAI21X1  _3505_
timestamp 0
transform 1 0 3190 0 1 4090
box -6 -8 106 248
use OAI21X1  _3506_
timestamp 0
transform -1 0 890 0 -1 3610
box -6 -8 106 248
use OAI21X1  _3507_
timestamp 0
transform -1 0 1090 0 -1 3610
box -6 -8 106 248
use MUX2X1  _3508_
timestamp 0
transform 1 0 6410 0 -1 4090
box -6 -8 126 248
use NOR2X1  _3509_
timestamp 0
transform -1 0 6710 0 -1 4090
box -6 -8 86 248
use NOR2X1  _3510_
timestamp 0
transform 1 0 6850 0 1 4090
box -6 -8 86 248
use AND2X2  _3511_
timestamp 0
transform -1 0 6770 0 1 4090
box -6 -8 106 248
use NAND2X1  _3512_
timestamp 0
transform 1 0 6630 0 1 4570
box -6 -8 86 248
use NAND2X1  _3513_
timestamp 0
transform 1 0 6810 0 1 4570
box -6 -8 86 248
use OAI21X1  _3514_
timestamp 0
transform -1 0 6630 0 -1 5050
box -6 -8 106 248
use NOR2X1  _3515_
timestamp 0
transform 1 0 7210 0 -1 4090
box -6 -8 86 248
use OAI21X1  _3516_
timestamp 0
transform -1 0 1350 0 1 5530
box -6 -8 106 248
use OAI21X1  _3517_
timestamp 0
transform 1 0 1050 0 1 5530
box -6 -8 106 248
use OAI21X1  _3518_
timestamp 0
transform -1 0 7610 0 1 11290
box -6 -8 106 248
use NAND2X1  _3519_
timestamp 0
transform -1 0 7410 0 1 11290
box -6 -8 86 248
use NOR2X1  _3520_
timestamp 0
transform 1 0 5370 0 1 11290
box -6 -8 86 248
use NAND2X1  _3521_
timestamp 0
transform -1 0 5630 0 1 11290
box -6 -8 86 248
use OAI21X1  _3522_
timestamp 0
transform -1 0 210 0 1 4570
box -6 -8 106 248
use NAND2X1  _3523_
timestamp 0
transform 1 0 290 0 -1 5050
box -6 -8 86 248
use INVX1  _3524_
timestamp 0
transform -1 0 550 0 1 4570
box -6 -8 66 248
use OAI21X1  _3525_
timestamp 0
transform 1 0 2090 0 1 3130
box -6 -8 106 248
use OAI21X1  _3526_
timestamp 0
transform 1 0 2270 0 -1 3610
box -6 -8 106 248
use AOI21X1  _3527_
timestamp 0
transform 1 0 7070 0 -1 4570
box -6 -8 106 248
use NOR2X1  _3528_
timestamp 0
transform -1 0 7070 0 1 4570
box -6 -8 86 248
use INVX8  _3529_
timestamp 0
transform -1 0 230 0 -1 9850
box -6 -8 126 248
use INVX1  _3530_
timestamp 0
transform 1 0 10130 0 -1 11770
box -6 -8 66 248
use NOR2X1  _3531_
timestamp 0
transform 1 0 6110 0 1 8410
box -6 -8 86 248
use INVX1  _3532_
timestamp 0
transform 1 0 5730 0 1 8410
box -6 -8 66 248
use NOR2X1  _3533_
timestamp 0
transform 1 0 11890 0 1 6970
box -6 -8 86 248
use NOR2X1  _3534_
timestamp 0
transform -1 0 9250 0 -1 6970
box -6 -8 86 248
use INVX1  _3535_
timestamp 0
transform 1 0 7690 0 -1 11770
box -6 -8 66 248
use INVX8  _3536_
timestamp 0
transform 1 0 6090 0 1 3610
box -6 -8 126 248
use AOI21X1  _3537_
timestamp 0
transform 1 0 5630 0 -1 5050
box -6 -8 106 248
use OAI21X1  _3538_
timestamp 0
transform 1 0 5610 0 -1 5530
box -6 -8 106 248
use AND2X2  _3539_
timestamp 0
transform 1 0 6210 0 -1 5530
box -6 -8 106 248
use AOI21X1  _3540_
timestamp 0
transform 1 0 6410 0 -1 5530
box -6 -8 106 248
use OAI21X1  _3541_
timestamp 0
transform -1 0 6370 0 1 5530
box -6 -8 106 248
use NAND2X1  _3542_
timestamp 0
transform -1 0 6170 0 1 5530
box -6 -8 86 248
use AOI21X1  _3543_
timestamp 0
transform 1 0 6010 0 -1 5530
box -6 -8 106 248
use OAI21X1  _3544_
timestamp 0
transform 1 0 5890 0 1 5530
box -6 -8 106 248
use OAI21X1  _3545_
timestamp 0
transform 1 0 5890 0 -1 6010
box -6 -8 106 248
use INVX4  _3546_
timestamp 0
transform -1 0 6330 0 1 3130
box -6 -8 86 248
use AOI21X1  _3547_
timestamp 0
transform 1 0 6430 0 1 5050
box -6 -8 106 248
use OAI21X1  _3548_
timestamp 0
transform 1 0 6530 0 -1 6010
box -6 -8 106 248
use AOI21X1  _3549_
timestamp 0
transform 1 0 6730 0 -1 6010
box -6 -8 106 248
use OAI21X1  _3550_
timestamp 0
transform 1 0 6570 0 1 6010
box -6 -8 106 248
use AOI21X1  _3551_
timestamp 0
transform -1 0 6870 0 1 6010
box -6 -8 106 248
use OAI21X1  _3552_
timestamp 0
transform 1 0 6870 0 -1 6970
box -6 -8 106 248
use OAI21X1  _3553_
timestamp 0
transform -1 0 7390 0 -1 7930
box -6 -8 106 248
use NAND3X1  _3554_
timestamp 0
transform 1 0 11270 0 1 11290
box -6 -8 106 248
use NOR2X1  _3555_
timestamp 0
transform 1 0 10930 0 1 11290
box -6 -8 86 248
use OR2X2  _3556_
timestamp 0
transform 1 0 10190 0 1 11290
box -6 -8 106 248
use NAND2X1  _3557_
timestamp 0
transform -1 0 9330 0 1 11290
box -6 -8 86 248
use NAND2X1  _3558_
timestamp 0
transform -1 0 10830 0 1 11290
box -6 -8 86 248
use NOR2X1  _3559_
timestamp 0
transform 1 0 11610 0 -1 11290
box -6 -8 86 248
use NAND2X1  _3560_
timestamp 0
transform 1 0 10070 0 -1 11290
box -6 -8 86 248
use NOR2X1  _3561_
timestamp 0
transform 1 0 10050 0 1 10330
box -6 -8 86 248
use NAND3X1  _3562_
timestamp 0
transform 1 0 9850 0 1 10330
box -6 -8 106 248
use NAND2X1  _3563_
timestamp 0
transform -1 0 9990 0 -1 10330
box -6 -8 86 248
use NAND3X1  _3564_
timestamp 0
transform -1 0 11950 0 1 11290
box -6 -8 106 248
use AND2X2  _3565_
timestamp 0
transform 1 0 12050 0 1 11290
box -6 -8 106 248
use AND2X2  _3566_
timestamp 0
transform 1 0 11470 0 1 11290
box -6 -8 106 248
use INVX1  _3567_
timestamp 0
transform 1 0 11110 0 1 11290
box -6 -8 66 248
use NAND3X1  _3568_
timestamp 0
transform 1 0 11250 0 -1 11770
box -6 -8 106 248
use NOR2X1  _3569_
timestamp 0
transform 1 0 9790 0 -1 11770
box -6 -8 86 248
use AND2X2  _3570_
timestamp 0
transform 1 0 10670 0 -1 11770
box -6 -8 106 248
use NOR2X1  _3571_
timestamp 0
transform 1 0 9610 0 -1 11770
box -6 -8 86 248
use NAND2X1  _3572_
timestamp 0
transform -1 0 9510 0 -1 11770
box -6 -8 86 248
use AND2X2  _3573_
timestamp 0
transform 1 0 11050 0 -1 11770
box -6 -8 106 248
use OAI21X1  _3574_
timestamp 0
transform -1 0 9470 0 1 11770
box -6 -8 106 248
use AND2X2  _3575_
timestamp 0
transform 1 0 8590 0 1 11770
box -6 -8 106 248
use NOR2X1  _3576_
timestamp 0
transform -1 0 8130 0 1 11770
box -6 -8 86 248
use NAND3X1  _3577_
timestamp 0
transform -1 0 9130 0 -1 11770
box -6 -8 106 248
use AND2X2  _3578_
timestamp 0
transform -1 0 9210 0 -1 11290
box -6 -8 106 248
use NAND3X1  _3579_
timestamp 0
transform -1 0 8330 0 1 11770
box -6 -8 106 248
use NOR2X1  _3580_
timestamp 0
transform -1 0 8770 0 1 11290
box -6 -8 86 248
use NAND3X1  _3581_
timestamp 0
transform 1 0 9650 0 1 10330
box -6 -8 106 248
use AND2X2  _3582_
timestamp 0
transform 1 0 9450 0 1 10330
box -6 -8 106 248
use NAND3X1  _3583_
timestamp 0
transform 1 0 8510 0 -1 11290
box -6 -8 106 248
use INVX1  _3584_
timestamp 0
transform -1 0 8490 0 1 11770
box -6 -8 66 248
use NAND3X1  _3585_
timestamp 0
transform 1 0 9170 0 1 11770
box -6 -8 106 248
use NOR2X1  _3586_
timestamp 0
transform -1 0 9070 0 1 11770
box -6 -8 86 248
use NAND3X1  _3587_
timestamp 0
transform -1 0 9330 0 -1 11770
box -6 -8 106 248
use AOI21X1  _3588_
timestamp 0
transform 1 0 8250 0 -1 11770
box -6 -8 106 248
use NAND3X1  _3589_
timestamp 0
transform -1 0 9150 0 1 11290
box -6 -8 106 248
use NOR2X1  _3590_
timestamp 0
transform -1 0 10690 0 -1 11290
box -6 -8 86 248
use NOR2X1  _3591_
timestamp 0
transform -1 0 10870 0 1 10810
box -6 -8 86 248
use MUX2X1  _3592_
timestamp 0
transform 1 0 8270 0 1 10330
box -6 -8 126 248
use NAND2X1  _3593_
timestamp 0
transform -1 0 6310 0 -1 11770
box -6 -8 86 248
use INVX1  _3594_
timestamp 0
transform -1 0 10450 0 1 11290
box -6 -8 66 248
use NAND3X1  _3595_
timestamp 0
transform -1 0 10650 0 1 11290
box -6 -8 106 248
use NAND3X1  _3596_
timestamp 0
transform 1 0 7010 0 -1 11770
box -6 -8 106 248
use INVX1  _3597_
timestamp 0
transform 1 0 6670 0 1 11770
box -6 -8 66 248
use NAND2X1  _3598_
timestamp 0
transform 1 0 11890 0 -1 10810
box -6 -8 86 248
use NAND3X1  _3599_
timestamp 0
transform -1 0 9030 0 1 10810
box -6 -8 106 248
use OAI21X1  _3600_
timestamp 0
transform 1 0 8730 0 1 10810
box -6 -8 106 248
use OR2X2  _3601_
timestamp 0
transform 1 0 8870 0 1 10330
box -6 -8 106 248
use NOR2X1  _3602_
timestamp 0
transform -1 0 10050 0 -1 11770
box -6 -8 86 248
use NAND3X1  _3603_
timestamp 0
transform -1 0 10390 0 -1 11770
box -6 -8 106 248
use NOR2X1  _3604_
timestamp 0
transform -1 0 8530 0 -1 11770
box -6 -8 86 248
use INVX1  _3605_
timestamp 0
transform -1 0 7950 0 1 11770
box -6 -8 66 248
use AOI22X1  _3606_
timestamp 0
transform -1 0 8150 0 -1 11770
box -6 -8 126 248
use NOR2X1  _3607_
timestamp 0
transform 1 0 7850 0 -1 11770
box -6 -8 86 248
use NOR2X1  _3608_
timestamp 0
transform 1 0 11450 0 -1 11770
box -6 -8 86 248
use NAND2X1  _3609_
timestamp 0
transform 1 0 11670 0 1 11290
box -6 -8 86 248
use OAI21X1  _3610_
timestamp 0
transform 1 0 11510 0 1 9370
box -6 -8 106 248
use OAI21X1  _3611_
timestamp 0
transform 1 0 11330 0 1 9370
box -6 -8 106 248
use AND2X2  _3612_
timestamp 0
transform 1 0 11690 0 -1 10810
box -6 -8 106 248
use OAI21X1  _3613_
timestamp 0
transform 1 0 11430 0 1 10330
box -6 -8 106 248
use OAI21X1  _3614_
timestamp 0
transform 1 0 11630 0 1 10330
box -6 -8 106 248
use NAND3X1  _3615_
timestamp 0
transform 1 0 11370 0 1 10810
box -6 -8 106 248
use MUX2X1  _3616_
timestamp 0
transform -1 0 8250 0 1 8890
box -6 -8 126 248
use OAI21X1  _3617_
timestamp 0
transform 1 0 12070 0 -1 10810
box -6 -8 106 248
use OAI21X1  _3618_
timestamp 0
transform 1 0 12010 0 1 10330
box -6 -8 106 248
use NOR2X1  _3619_
timestamp 0
transform -1 0 11650 0 -1 10330
box -6 -8 86 248
use NAND3X1  _3620_
timestamp 0
transform 1 0 8830 0 -1 11770
box -6 -8 106 248
use AOI21X1  _3621_
timestamp 0
transform 1 0 8210 0 -1 10810
box -6 -8 106 248
use OAI21X1  _3622_
timestamp 0
transform 1 0 8170 0 1 10810
box -6 -8 106 248
use AOI21X1  _3623_
timestamp 0
transform 1 0 11170 0 1 10810
box -6 -8 106 248
use NAND2X1  _3624_
timestamp 0
transform -1 0 11210 0 -1 10810
box -6 -8 86 248
use OAI21X1  _3625_
timestamp 0
transform 1 0 10830 0 1 10330
box -6 -8 106 248
use OAI21X1  _3626_
timestamp 0
transform 1 0 11030 0 1 10330
box -6 -8 106 248
use AND2X2  _3627_
timestamp 0
transform 1 0 10970 0 1 10810
box -6 -8 106 248
use OAI21X1  _3628_
timestamp 0
transform 1 0 8010 0 -1 10810
box -6 -8 106 248
use AOI21X1  _3629_
timestamp 0
transform 1 0 7670 0 1 10330
box -6 -8 106 248
use OAI21X1  _3630_
timestamp 0
transform 1 0 7630 0 -1 10330
box -6 -8 106 248
use NAND2X1  _3631_
timestamp 0
transform -1 0 7570 0 1 10330
box -6 -8 86 248
use NOR2X1  _3632_
timestamp 0
transform 1 0 7070 0 -1 10330
box -6 -8 86 248
use OAI21X1  _3633_
timestamp 0
transform 1 0 8070 0 1 10330
box -6 -8 106 248
use AOI21X1  _3634_
timestamp 0
transform 1 0 8750 0 -1 10810
box -6 -8 106 248
use INVX1  _3635_
timestamp 0
transform 1 0 8410 0 -1 10810
box -6 -8 66 248
use OAI21X1  _3636_
timestamp 0
transform -1 0 6970 0 -1 10330
box -6 -8 106 248
use NOR2X1  _3637_
timestamp 0
transform 1 0 8770 0 1 9850
box -6 -8 86 248
use NAND2X1  _3638_
timestamp 0
transform 1 0 10870 0 -1 11770
box -6 -8 86 248
use AOI21X1  _3639_
timestamp 0
transform 1 0 8630 0 -1 11770
box -6 -8 106 248
use NAND3X1  _3640_
timestamp 0
transform 1 0 9490 0 1 9850
box -6 -8 106 248
use NAND2X1  _3641_
timestamp 0
transform 1 0 8990 0 1 9370
box -6 -8 86 248
use OAI21X1  _3642_
timestamp 0
transform -1 0 7430 0 -1 9370
box -6 -8 106 248
use NAND2X1  _3643_
timestamp 0
transform 1 0 7150 0 -1 9370
box -6 -8 86 248
use AND2X2  _3644_
timestamp 0
transform -1 0 9450 0 -1 10330
box -6 -8 106 248
use OAI21X1  _3645_
timestamp 0
transform -1 0 10530 0 1 10330
box -6 -8 106 248
use OAI21X1  _3646_
timestamp 0
transform 1 0 9150 0 -1 10330
box -6 -8 106 248
use OAI21X1  _3647_
timestamp 0
transform 1 0 10590 0 1 9850
box -6 -8 106 248
use OAI21X1  _3648_
timestamp 0
transform 1 0 10910 0 -1 9370
box -6 -8 106 248
use NAND3X1  _3649_
timestamp 0
transform 1 0 11010 0 -1 9850
box -6 -8 106 248
use OAI21X1  _3650_
timestamp 0
transform -1 0 11490 0 -1 8890
box -6 -8 106 248
use OAI21X1  _3651_
timestamp 0
transform 1 0 6810 0 -1 11770
box -6 -8 106 248
use NAND3X1  _3652_
timestamp 0
transform 1 0 4870 0 -1 11770
box -6 -8 106 248
use AND2X2  _3653_
timestamp 0
transform 1 0 4670 0 -1 11770
box -6 -8 106 248
use AOI21X1  _3654_
timestamp 0
transform 1 0 4470 0 -1 11770
box -6 -8 106 248
use AOI21X1  _3655_
timestamp 0
transform 1 0 4270 0 -1 11770
box -6 -8 106 248
use NOR2X1  _3656_
timestamp 0
transform 1 0 5470 0 1 11770
box -6 -8 86 248
use OAI22X1  _3657_
timestamp 0
transform 1 0 5430 0 -1 11770
box -6 -8 126 248
use AOI21X1  _3658_
timestamp 0
transform 1 0 5270 0 1 11770
box -6 -8 106 248
use NOR2X1  _3659_
timestamp 0
transform 1 0 4690 0 1 11770
box -6 -8 86 248
use AOI21X1  _3660_
timestamp 0
transform 1 0 4490 0 1 11770
box -6 -8 106 248
use OAI22X1  _3661_
timestamp 0
transform 1 0 4870 0 1 11770
box -6 -8 126 248
use NAND3X1  _3662_
timestamp 0
transform 1 0 6610 0 -1 11770
box -6 -8 106 248
use AND2X2  _3663_
timestamp 0
transform 1 0 6410 0 -1 11770
box -6 -8 106 248
use NAND3X1  _3664_
timestamp 0
transform 1 0 5650 0 -1 11770
box -6 -8 106 248
use NAND2X1  _3665_
timestamp 0
transform 1 0 5250 0 -1 11770
box -6 -8 86 248
use NAND2X1  _3666_
timestamp 0
transform 1 0 5850 0 -1 11770
box -6 -8 86 248
use OAI21X1  _3667_
timestamp 0
transform -1 0 3810 0 -1 11770
box -6 -8 106 248
use NAND2X1  _3668_
timestamp 0
transform 1 0 3950 0 1 11770
box -6 -8 86 248
use NOR2X1  _3669_
timestamp 0
transform -1 0 3510 0 1 11770
box -6 -8 86 248
use NAND2X1  _3670_
timestamp 0
transform -1 0 3610 0 -1 11770
box -6 -8 86 248
use AOI22X1  _3671_
timestamp 0
transform 1 0 4210 0 -1 11290
box -6 -8 126 248
use NOR2X1  _3672_
timestamp 0
transform 1 0 4270 0 1 11290
box -6 -8 86 248
use OAI21X1  _3673_
timestamp 0
transform 1 0 6030 0 -1 11770
box -6 -8 106 248
use OAI21X1  _3674_
timestamp 0
transform -1 0 10850 0 -1 10810
box -6 -8 106 248
use NAND2X1  _3675_
timestamp 0
transform -1 0 10650 0 -1 10810
box -6 -8 86 248
use OAI21X1  _3676_
timestamp 0
transform 1 0 4190 0 1 5050
box -6 -8 106 248
use INVX1  _3677_
timestamp 0
transform -1 0 4290 0 -1 5530
box -6 -8 66 248
use OAI21X1  _3678_
timestamp 0
transform 1 0 4690 0 1 6970
box -6 -8 106 248
use AOI21X1  _3679_
timestamp 0
transform -1 0 4990 0 1 6970
box -6 -8 106 248
use OAI21X1  _3680_
timestamp 0
transform -1 0 5190 0 1 6970
box -6 -8 106 248
use NAND2X1  _3681_
timestamp 0
transform -1 0 4870 0 1 7450
box -6 -8 86 248
use INVX1  _3682_
timestamp 0
transform 1 0 1690 0 -1 7930
box -6 -8 66 248
use OAI22X1  _3683_
timestamp 0
transform 1 0 6310 0 -1 6010
box -6 -8 126 248
use OAI22X1  _3684_
timestamp 0
transform 1 0 6650 0 -1 6970
box -6 -8 126 248
use OAI22X1  _3685_
timestamp 0
transform 1 0 6930 0 -1 6010
box -6 -8 126 248
use OAI22X1  _3686_
timestamp 0
transform 1 0 6710 0 1 6490
box -6 -8 126 248
use OAI21X1  _3687_
timestamp 0
transform 1 0 4930 0 -1 6010
box -6 -8 106 248
use NOR2X1  _3688_
timestamp 0
transform -1 0 5010 0 -1 6490
box -6 -8 86 248
use OAI22X1  _3689_
timestamp 0
transform 1 0 5130 0 -1 6970
box -6 -8 126 248
use NOR2X1  _3690_
timestamp 0
transform -1 0 4830 0 -1 6490
box -6 -8 86 248
use OAI21X1  _3691_
timestamp 0
transform -1 0 4810 0 1 6010
box -6 -8 106 248
use NOR2X1  _3692_
timestamp 0
transform 1 0 4530 0 1 6010
box -6 -8 86 248
use OAI22X1  _3693_
timestamp 0
transform 1 0 4910 0 1 6010
box -6 -8 126 248
use OAI22X1  _3694_
timestamp 0
transform -1 0 6210 0 -1 6010
box -6 -8 126 248
use INVX1  _3695_
timestamp 0
transform 1 0 1750 0 -1 6490
box -6 -8 66 248
use OAI22X1  _3696_
timestamp 0
transform 1 0 7630 0 1 6970
box -6 -8 126 248
use OAI22X1  _3697_
timestamp 0
transform 1 0 7830 0 -1 6010
box -6 -8 126 248
use OAI21X1  _3698_
timestamp 0
transform 1 0 6730 0 -1 6490
box -6 -8 106 248
use NOR2X1  _3699_
timestamp 0
transform 1 0 6930 0 -1 6490
box -6 -8 86 248
use OAI22X1  _3700_
timestamp 0
transform -1 0 7230 0 -1 6490
box -6 -8 126 248
use INVX8  _3701_
timestamp 0
transform 1 0 4690 0 1 3130
box -6 -8 126 248
use AOI21X1  _3702_
timestamp 0
transform 1 0 4390 0 -1 5530
box -6 -8 106 248
use OAI21X1  _3703_
timestamp 0
transform 1 0 4450 0 1 6490
box -6 -8 106 248
use NOR2X1  _3704_
timestamp 0
transform 1 0 4870 0 1 6490
box -6 -8 86 248
use OAI21X1  _3705_
timestamp 0
transform -1 0 5030 0 -1 6970
box -6 -8 106 248
use AOI22X1  _3706_
timestamp 0
transform -1 0 4830 0 -1 6970
box -6 -8 126 248
use OAI21X1  _3707_
timestamp 0
transform -1 0 5150 0 1 6490
box -6 -8 106 248
use AOI22X1  _3708_
timestamp 0
transform 1 0 4650 0 1 6490
box -6 -8 126 248
use INVX1  _3709_
timestamp 0
transform 1 0 2510 0 1 7450
box -6 -8 66 248
use NAND3X1  _3710_
timestamp 0
transform 1 0 9810 0 1 11290
box -6 -8 106 248
use NOR2X1  _3711_
timestamp 0
transform 1 0 9710 0 -1 11290
box -6 -8 86 248
use NAND3X1  _3712_
timestamp 0
transform 1 0 9690 0 1 10810
box -6 -8 106 248
use AND2X2  _3713_
timestamp 0
transform 1 0 10070 0 1 10810
box -6 -8 106 248
use NOR2X1  _3714_
timestamp 0
transform 1 0 8770 0 -1 9850
box -6 -8 86 248
use OAI21X1  _3715_
timestamp 0
transform -1 0 9050 0 -1 9850
box -6 -8 106 248
use INVX1  _3716_
timestamp 0
transform -1 0 9610 0 1 9370
box -6 -8 66 248
use NOR2X1  _3717_
timestamp 0
transform -1 0 10530 0 1 10810
box -6 -8 86 248
use INVX1  _3718_
timestamp 0
transform 1 0 10630 0 1 10810
box -6 -8 66 248
use OAI21X1  _3719_
timestamp 0
transform -1 0 9250 0 -1 9850
box -6 -8 106 248
use OAI21X1  _3720_
timestamp 0
transform 1 0 9350 0 -1 9850
box -6 -8 106 248
use OAI21X1  _3721_
timestamp 0
transform -1 0 10770 0 -1 10330
box -6 -8 106 248
use NAND2X1  _3722_
timestamp 0
transform -1 0 10570 0 -1 10330
box -6 -8 86 248
use NAND2X1  _3723_
timestamp 0
transform 1 0 10830 0 -1 9850
box -6 -8 86 248
use NOR2X1  _3724_
timestamp 0
transform 1 0 9510 0 -1 10810
box -6 -8 86 248
use NAND3X1  _3725_
timestamp 0
transform 1 0 8370 0 1 9850
box -6 -8 106 248
use NAND2X1  _3726_
timestamp 0
transform -1 0 8310 0 -1 9850
box -6 -8 86 248
use NAND2X1  _3727_
timestamp 0
transform 1 0 9690 0 -1 10810
box -6 -8 86 248
use OAI21X1  _3728_
timestamp 0
transform -1 0 10330 0 1 10330
box -6 -8 106 248
use OAI21X1  _3729_
timestamp 0
transform 1 0 10090 0 -1 10330
box -6 -8 106 248
use INVX1  _3730_
timestamp 0
transform 1 0 10030 0 -1 10810
box -6 -8 66 248
use OAI21X1  _3731_
timestamp 0
transform 1 0 8490 0 1 11290
box -6 -8 106 248
use NAND2X1  _3732_
timestamp 0
transform 1 0 8870 0 1 11290
box -6 -8 86 248
use NAND2X1  _3733_
timestamp 0
transform -1 0 3990 0 -1 11770
box -6 -8 86 248
use NOR2X1  _3734_
timestamp 0
transform -1 0 4170 0 -1 11770
box -6 -8 86 248
use AND2X2  _3735_
timestamp 0
transform 1 0 7690 0 1 11770
box -6 -8 106 248
use AOI22X1  _3736_
timestamp 0
transform -1 0 7390 0 1 11770
box -6 -8 126 248
use NOR2X1  _3737_
timestamp 0
transform -1 0 5910 0 1 11770
box -6 -8 86 248
use AND2X2  _3738_
timestamp 0
transform 1 0 9630 0 1 11290
box -6 -8 106 248
use AND2X2  _3739_
timestamp 0
transform 1 0 9430 0 1 11290
box -6 -8 106 248
use AND2X2  _3740_
timestamp 0
transform 1 0 9310 0 -1 11290
box -6 -8 106 248
use NOR2X1  _3741_
timestamp 0
transform -1 0 10870 0 -1 11290
box -6 -8 86 248
use NAND2X1  _3742_
timestamp 0
transform 1 0 11310 0 -1 10810
box -6 -8 86 248
use OAI21X1  _3743_
timestamp 0
transform 1 0 11490 0 -1 10810
box -6 -8 106 248
use OAI21X1  _3744_
timestamp 0
transform 1 0 11230 0 1 10330
box -6 -8 106 248
use OAI21X1  _3745_
timestamp 0
transform -1 0 10730 0 1 10330
box -6 -8 106 248
use OAI21X1  _3746_
timestamp 0
transform -1 0 10390 0 -1 10330
box -6 -8 106 248
use NOR2X1  _3747_
timestamp 0
transform -1 0 10310 0 1 9850
box -6 -8 86 248
use INVX1  _3748_
timestamp 0
transform -1 0 11030 0 -1 11290
box -6 -8 66 248
use OAI21X1  _3749_
timestamp 0
transform -1 0 11390 0 -1 9370
box -6 -8 106 248
use OAI21X1  _3750_
timestamp 0
transform 1 0 11090 0 -1 9370
box -6 -8 106 248
use AOI22X1  _3751_
timestamp 0
transform -1 0 8210 0 1 11290
box -6 -8 126 248
use AOI21X1  _3752_
timestamp 0
transform -1 0 6990 0 1 10810
box -6 -8 106 248
use NOR2X1  _3753_
timestamp 0
transform -1 0 6870 0 1 11290
box -6 -8 86 248
use AOI21X1  _3754_
timestamp 0
transform 1 0 4450 0 1 11290
box -6 -8 106 248
use OAI21X1  _3755_
timestamp 0
transform 1 0 3090 0 1 10810
box -6 -8 106 248
use OAI21X1  _3756_
timestamp 0
transform 1 0 4130 0 -1 5050
box -6 -8 106 248
use NOR2X1  _3757_
timestamp 0
transform 1 0 4610 0 1 7450
box -6 -8 86 248
use OAI21X1  _3758_
timestamp 0
transform -1 0 5210 0 -1 7450
box -6 -8 106 248
use AOI22X1  _3759_
timestamp 0
transform -1 0 5010 0 -1 7450
box -6 -8 126 248
use OAI21X1  _3760_
timestamp 0
transform -1 0 4430 0 -1 5050
box -6 -8 106 248
use INVX1  _3761_
timestamp 0
transform -1 0 4410 0 -1 7930
box -6 -8 66 248
use NAND3X1  _3762_
timestamp 0
transform -1 0 4550 0 -1 8410
box -6 -8 106 248
use AOI22X1  _3763_
timestamp 0
transform -1 0 4310 0 1 7450
box -6 -8 126 248
use OAI21X1  _3764_
timestamp 0
transform -1 0 3570 0 1 8410
box -6 -8 106 248
use NAND2X1  _3765_
timestamp 0
transform -1 0 4730 0 -1 8410
box -6 -8 86 248
use OAI21X1  _3766_
timestamp 0
transform 1 0 2290 0 1 5050
box -6 -8 106 248
use INVX1  _3767_
timestamp 0
transform -1 0 2550 0 1 5050
box -6 -8 66 248
use OAI21X1  _3768_
timestamp 0
transform -1 0 2750 0 1 5050
box -6 -8 106 248
use AND2X2  _3769_
timestamp 0
transform -1 0 2950 0 1 5050
box -6 -8 106 248
use AOI21X1  _3770_
timestamp 0
transform -1 0 3930 0 1 5050
box -6 -8 106 248
use OAI21X1  _3771_
timestamp 0
transform 1 0 3450 0 1 5050
box -6 -8 106 248
use INVX1  _3772_
timestamp 0
transform -1 0 1130 0 -1 9370
box -6 -8 66 248
use INVX8  _3773_
timestamp 0
transform 1 0 5870 0 1 3610
box -6 -8 126 248
use AOI21X1  _3774_
timestamp 0
transform 1 0 5090 0 -1 4090
box -6 -8 106 248
use OAI21X1  _3775_
timestamp 0
transform -1 0 5130 0 -1 5050
box -6 -8 106 248
use INVX1  _3776_
timestamp 0
transform -1 0 4930 0 -1 5050
box -6 -8 66 248
use NAND2X1  _3777_
timestamp 0
transform 1 0 4950 0 1 5530
box -6 -8 86 248
use INVX1  _3778_
timestamp 0
transform 1 0 4790 0 1 5530
box -6 -8 66 248
use NAND3X1  _3779_
timestamp 0
transform 1 0 4590 0 1 5530
box -6 -8 106 248
use AOI22X1  _3780_
timestamp 0
transform 1 0 5270 0 -1 6490
box -6 -8 126 248
use INVX1  _3781_
timestamp 0
transform -1 0 5490 0 1 6490
box -6 -8 66 248
use NAND2X1  _3782_
timestamp 0
transform -1 0 4490 0 1 5530
box -6 -8 86 248
use OAI21X1  _3783_
timestamp 0
transform 1 0 3870 0 1 5530
box -6 -8 106 248
use OAI21X1  _3784_
timestamp 0
transform -1 0 5390 0 1 5530
box -6 -8 106 248
use INVX4  _3785_
timestamp 0
transform 1 0 7590 0 1 3610
box -6 -8 86 248
use AOI21X1  _3786_
timestamp 0
transform 1 0 7450 0 -1 4570
box -6 -8 106 248
use OAI21X1  _3787_
timestamp 0
transform -1 0 7510 0 -1 5050
box -6 -8 106 248
use INVX1  _3788_
timestamp 0
transform -1 0 7310 0 -1 5050
box -6 -8 66 248
use NAND2X1  _3789_
timestamp 0
transform -1 0 7350 0 1 5050
box -6 -8 86 248
use AOI21X1  _3790_
timestamp 0
transform -1 0 6330 0 1 5050
box -6 -8 106 248
use OAI22X1  _3791_
timestamp 0
transform -1 0 6750 0 1 5050
box -6 -8 126 248
use AOI21X1  _3792_
timestamp 0
transform 1 0 7070 0 1 5050
box -6 -8 106 248
use OAI22X1  _3793_
timestamp 0
transform -1 0 6970 0 1 5050
box -6 -8 126 248
use INVX1  _3794_
timestamp 0
transform 1 0 8030 0 -1 4570
box -6 -8 66 248
use OAI21X1  _3795_
timestamp 0
transform -1 0 9730 0 1 6970
box -6 -8 106 248
use OAI21X1  _3796_
timestamp 0
transform 1 0 8350 0 1 7450
box -6 -8 106 248
use OR2X2  _3797_
timestamp 0
transform 1 0 7730 0 -1 8890
box -6 -8 106 248
use NAND2X1  _3798_
timestamp 0
transform 1 0 7010 0 -1 8890
box -6 -8 86 248
use NOR2X1  _3799_
timestamp 0
transform -1 0 7250 0 1 8890
box -6 -8 86 248
use OAI21X1  _3800_
timestamp 0
transform -1 0 7450 0 1 8890
box -6 -8 106 248
use OAI21X1  _3801_
timestamp 0
transform 1 0 5710 0 -1 8890
box -6 -8 106 248
use OAI21X1  _3802_
timestamp 0
transform -1 0 6050 0 1 8890
box -6 -8 106 248
use OAI21X1  _3803_
timestamp 0
transform 1 0 5750 0 1 8890
box -6 -8 106 248
use OAI21X1  _3804_
timestamp 0
transform 1 0 5370 0 1 8890
box -6 -8 106 248
use OR2X2  _3805_
timestamp 0
transform 1 0 5410 0 1 9370
box -6 -8 106 248
use AOI21X1  _3806_
timestamp 0
transform 1 0 5090 0 -1 9850
box -6 -8 106 248
use INVX1  _3807_
timestamp 0
transform -1 0 5610 0 -1 8890
box -6 -8 66 248
use NAND3X1  _3808_
timestamp 0
transform -1 0 8030 0 1 8890
box -6 -8 106 248
use NOR2X1  _3809_
timestamp 0
transform -1 0 8130 0 -1 9370
box -6 -8 86 248
use OAI21X1  _3810_
timestamp 0
transform 1 0 7850 0 -1 9370
box -6 -8 106 248
use OAI21X1  _3811_
timestamp 0
transform -1 0 7630 0 -1 9370
box -6 -8 106 248
use NAND3X1  _3812_
timestamp 0
transform 1 0 10490 0 -1 11770
box -6 -8 106 248
use NOR2X1  _3813_
timestamp 0
transform -1 0 9970 0 -1 11290
box -6 -8 86 248
use NAND2X1  _3814_
timestamp 0
transform 1 0 9890 0 1 10810
box -6 -8 86 248
use NOR2X1  _3815_
timestamp 0
transform -1 0 9950 0 -1 10810
box -6 -8 86 248
use OAI21X1  _3816_
timestamp 0
transform -1 0 9810 0 -1 10330
box -6 -8 106 248
use OAI21X1  _3817_
timestamp 0
transform 1 0 9190 0 -1 9370
box -6 -8 106 248
use OAI21X1  _3818_
timestamp 0
transform -1 0 9090 0 -1 9370
box -6 -8 106 248
use OAI21X1  _3819_
timestamp 0
transform 1 0 10190 0 -1 10810
box -6 -8 106 248
use NAND2X1  _3820_
timestamp 0
transform 1 0 10270 0 1 10810
box -6 -8 86 248
use OAI21X1  _3821_
timestamp 0
transform 1 0 6590 0 1 11290
box -6 -8 106 248
use NOR2X1  _3822_
timestamp 0
transform -1 0 3450 0 -1 11770
box -6 -8 86 248
use OAI22X1  _3823_
timestamp 0
transform -1 0 8410 0 -1 11290
box -6 -8 126 248
use NAND2X1  _3824_
timestamp 0
transform 1 0 7330 0 -1 11290
box -6 -8 86 248
use NOR2X1  _3825_
timestamp 0
transform -1 0 10090 0 1 11290
box -6 -8 86 248
use NAND2X1  _3826_
timestamp 0
transform 1 0 9510 0 1 10810
box -6 -8 86 248
use NOR2X1  _3827_
timestamp 0
transform -1 0 9410 0 -1 10810
box -6 -8 86 248
use NAND2X1  _3828_
timestamp 0
transform 1 0 9150 0 -1 10810
box -6 -8 86 248
use OAI21X1  _3829_
timestamp 0
transform 1 0 8950 0 -1 10810
box -6 -8 106 248
use OAI21X1  _3830_
timestamp 0
transform 1 0 7450 0 -1 10330
box -6 -8 106 248
use INVX1  _3831_
timestamp 0
transform 1 0 7710 0 -1 9370
box -6 -8 66 248
use NOR2X1  _3832_
timestamp 0
transform 1 0 8590 0 -1 9850
box -6 -8 86 248
use MUX2X1  _3833_
timestamp 0
transform 1 0 8770 0 1 9370
box -6 -8 126 248
use MUX2X1  _3834_
timestamp 0
transform -1 0 8850 0 1 8890
box -6 -8 126 248
use NAND2X1  _3835_
timestamp 0
transform 1 0 8950 0 1 8890
box -6 -8 86 248
use NAND3X1  _3836_
timestamp 0
transform 1 0 9250 0 1 10330
box -6 -8 106 248
use OAI21X1  _3837_
timestamp 0
transform -1 0 8590 0 1 10330
box -6 -8 106 248
use NAND2X1  _3838_
timestamp 0
transform 1 0 8690 0 1 10330
box -6 -8 86 248
use MUX2X1  _3839_
timestamp 0
transform 1 0 8930 0 -1 10330
box -6 -8 126 248
use OAI21X1  _3840_
timestamp 0
transform -1 0 8650 0 -1 10330
box -6 -8 106 248
use OAI21X1  _3841_
timestamp 0
transform -1 0 8450 0 -1 10330
box -6 -8 106 248
use AOI22X1  _3842_
timestamp 0
transform 1 0 9130 0 1 10810
box -6 -8 126 248
use NOR2X1  _3843_
timestamp 0
transform -1 0 8450 0 1 10810
box -6 -8 86 248
use INVX1  _3844_
timestamp 0
transform 1 0 7690 0 -1 10810
box -6 -8 66 248
use INVX1  _3845_
timestamp 0
transform 1 0 9350 0 1 10810
box -6 -8 66 248
use NAND3X1  _3846_
timestamp 0
transform 1 0 8910 0 -1 11290
box -6 -8 106 248
use NOR2X1  _3847_
timestamp 0
transform 1 0 8190 0 1 9850
box -6 -8 86 248
use OAI21X1  _3848_
timestamp 0
transform -1 0 8130 0 -1 8410
box -6 -8 106 248
use NAND3X1  _3849_
timestamp 0
transform 1 0 7830 0 -1 8410
box -6 -8 106 248
use NAND2X1  _3850_
timestamp 0
transform 1 0 8010 0 1 9850
box -6 -8 86 248
use OAI21X1  _3851_
timestamp 0
transform 1 0 7650 0 -1 9850
box -6 -8 106 248
use OAI21X1  _3852_
timestamp 0
transform -1 0 7950 0 -1 9850
box -6 -8 106 248
use OAI21X1  _3853_
timestamp 0
transform -1 0 7710 0 1 9850
box -6 -8 106 248
use OAI21X1  _3854_
timestamp 0
transform -1 0 7570 0 -1 9850
box -6 -8 106 248
use OAI21X1  _3855_
timestamp 0
transform 1 0 7870 0 1 10330
box -6 -8 106 248
use OAI21X1  _3856_
timestamp 0
transform -1 0 7350 0 -1 10330
box -6 -8 106 248
use INVX1  _3857_
timestamp 0
transform -1 0 8410 0 1 8410
box -6 -8 66 248
use AND2X2  _3858_
timestamp 0
transform 1 0 8710 0 -1 11290
box -6 -8 106 248
use NAND3X1  _3859_
timestamp 0
transform 1 0 7890 0 1 11290
box -6 -8 106 248
use NOR2X1  _3860_
timestamp 0
transform 1 0 4830 0 1 11290
box -6 -8 86 248
use NAND2X1  _3861_
timestamp 0
transform 1 0 8570 0 -1 10810
box -6 -8 86 248
use AND2X2  _3862_
timestamp 0
transform -1 0 8890 0 1 11770
box -6 -8 106 248
use NOR2X1  _3863_
timestamp 0
transform -1 0 10330 0 -1 11290
box -6 -8 86 248
use NAND3X1  _3864_
timestamp 0
transform 1 0 9510 0 -1 11290
box -6 -8 106 248
use AOI21X1  _3865_
timestamp 0
transform 1 0 8090 0 -1 11290
box -6 -8 106 248
use NOR2X1  _3866_
timestamp 0
transform 1 0 5690 0 -1 11290
box -6 -8 86 248
use NOR2X1  _3867_
timestamp 0
transform -1 0 7590 0 -1 11290
box -6 -8 86 248
use OAI21X1  _3868_
timestamp 0
transform -1 0 8670 0 1 9850
box -6 -8 106 248
use NAND2X1  _3869_
timestamp 0
transform 1 0 8010 0 -1 10330
box -6 -8 86 248
use AOI22X1  _3870_
timestamp 0
transform -1 0 7990 0 -1 11290
box -6 -8 126 248
use NOR2X1  _3871_
timestamp 0
transform 1 0 6410 0 1 11290
box -6 -8 86 248
use NAND2X1  _3872_
timestamp 0
transform 1 0 5730 0 1 11290
box -6 -8 86 248
use AOI21X1  _3873_
timestamp 0
transform -1 0 9650 0 -1 9850
box -6 -8 106 248
use OAI21X1  _3874_
timestamp 0
transform 1 0 9910 0 -1 9850
box -6 -8 106 248
use OAI21X1  _3875_
timestamp 0
transform 1 0 6950 0 -1 9370
box -6 -8 106 248
use NAND2X1  _3876_
timestamp 0
transform 1 0 5050 0 -1 9370
box -6 -8 86 248
use NAND2X1  _3877_
timestamp 0
transform -1 0 4750 0 -1 9370
box -6 -8 86 248
use OR2X2  _3878_
timestamp 0
transform 1 0 4850 0 -1 9370
box -6 -8 106 248
use MUX2X1  _3879_
timestamp 0
transform 1 0 4610 0 1 8890
box -6 -8 126 248
use OAI21X1  _3880_
timestamp 0
transform 1 0 5170 0 1 8410
box -6 -8 106 248
use NAND2X1  _3881_
timestamp 0
transform -1 0 5450 0 1 8410
box -6 -8 86 248
use INVX1  _3882_
timestamp 0
transform -1 0 4450 0 1 7930
box -6 -8 66 248
use OAI21X1  _3883_
timestamp 0
transform -1 0 5110 0 1 8890
box -6 -8 106 248
use NAND2X1  _3884_
timestamp 0
transform -1 0 4910 0 1 8890
box -6 -8 86 248
use INVX1  _3885_
timestamp 0
transform 1 0 5210 0 1 8890
box -6 -8 66 248
use NOR2X1  _3886_
timestamp 0
transform 1 0 9710 0 1 9370
box -6 -8 86 248
use NAND3X1  _3887_
timestamp 0
transform 1 0 10430 0 -1 11290
box -6 -8 106 248
use NAND2X1  _3888_
timestamp 0
transform 1 0 10390 0 -1 10810
box -6 -8 86 248
use NAND2X1  _3889_
timestamp 0
transform -1 0 10950 0 -1 10330
box -6 -8 86 248
use NOR2X1  _3890_
timestamp 0
transform -1 0 10870 0 1 9850
box -6 -8 86 248
use NAND2X1  _3891_
timestamp 0
transform 1 0 10950 0 1 9850
box -6 -8 86 248
use NOR2X1  _3892_
timestamp 0
transform -1 0 8890 0 -1 8410
box -6 -8 86 248
use OAI21X1  _3893_
timestamp 0
transform -1 0 8710 0 -1 8410
box -6 -8 106 248
use NAND3X1  _3894_
timestamp 0
transform -1 0 11410 0 1 7930
box -6 -8 106 248
use AOI21X1  _3895_
timestamp 0
transform 1 0 11110 0 1 7930
box -6 -8 106 248
use NAND2X1  _3896_
timestamp 0
transform 1 0 11870 0 1 7930
box -6 -8 86 248
use OAI21X1  _3897_
timestamp 0
transform 1 0 11130 0 1 9850
box -6 -8 106 248
use NAND2X1  _3898_
timestamp 0
transform 1 0 8310 0 1 11290
box -6 -8 86 248
use NOR2X1  _3899_
timestamp 0
transform -1 0 5730 0 1 11770
box -6 -8 86 248
use NAND2X1  _3900_
timestamp 0
transform 1 0 4130 0 1 11770
box -6 -8 86 248
use NAND2X1  _3901_
timestamp 0
transform -1 0 5150 0 -1 11770
box -6 -8 86 248
use NOR2X1  _3902_
timestamp 0
transform 1 0 5010 0 1 11290
box -6 -8 86 248
use AND2X2  _3903_
timestamp 0
transform 1 0 7490 0 1 11770
box -6 -8 106 248
use AOI22X1  _3904_
timestamp 0
transform -1 0 7170 0 1 11770
box -6 -8 126 248
use NOR2X1  _3905_
timestamp 0
transform -1 0 6570 0 1 11770
box -6 -8 86 248
use NAND2X1  _3906_
timestamp 0
transform 1 0 5090 0 1 11770
box -6 -8 86 248
use INVX1  _3907_
timestamp 0
transform -1 0 8290 0 -1 9370
box -6 -8 66 248
use AOI22X1  _3908_
timestamp 0
transform -1 0 6950 0 1 11770
box -6 -8 126 248
use NOR2X1  _3909_
timestamp 0
transform -1 0 6090 0 1 11770
box -6 -8 86 248
use NAND2X1  _3910_
timestamp 0
transform 1 0 5910 0 1 11290
box -6 -8 86 248
use OAI21X1  _3911_
timestamp 0
transform -1 0 4650 0 1 5050
box -6 -8 106 248
use NOR2X1  _3912_
timestamp 0
transform 1 0 4390 0 1 5050
box -6 -8 86 248
use OAI22X1  _3913_
timestamp 0
transform -1 0 4710 0 -1 5530
box -6 -8 126 248
use INVX1  _3914_
timestamp 0
transform 1 0 4270 0 1 4570
box -6 -8 66 248
use OAI21X1  _3915_
timestamp 0
transform 1 0 4810 0 -1 5530
box -6 -8 106 248
use NOR2X1  _3916_
timestamp 0
transform 1 0 5010 0 -1 5530
box -6 -8 86 248
use OAI22X1  _3917_
timestamp 0
transform 1 0 5390 0 -1 5530
box -6 -8 126 248
use NOR2X1  _3918_
timestamp 0
transform -1 0 4770 0 -1 5050
box -6 -8 86 248
use INVX1  _3919_
timestamp 0
transform 1 0 4810 0 -1 4570
box -6 -8 66 248
use INVX1  _3920_
timestamp 0
transform 1 0 4530 0 -1 5050
box -6 -8 66 248
use NAND3X1  _3921_
timestamp 0
transform 1 0 850 0 -1 5050
box -6 -8 106 248
use NAND2X1  _3922_
timestamp 0
transform 1 0 950 0 -1 5530
box -6 -8 86 248
use AOI22X1  _3923_
timestamp 0
transform 1 0 470 0 -1 5050
box -6 -8 126 248
use NAND3X1  _3924_
timestamp 0
transform 1 0 830 0 1 4570
box -6 -8 106 248
use OAI21X1  _3925_
timestamp 0
transform 1 0 5130 0 -1 6010
box -6 -8 106 248
use NOR2X1  _3926_
timestamp 0
transform 1 0 5330 0 -1 6010
box -6 -8 86 248
use OAI21X1  _3927_
timestamp 0
transform -1 0 4830 0 -1 6010
box -6 -8 106 248
use NOR2X1  _3928_
timestamp 0
transform 1 0 5510 0 -1 6010
box -6 -8 86 248
use INVX1  _3929_
timestamp 0
transform -1 0 4670 0 1 4570
box -6 -8 66 248
use NAND3X1  _3930_
timestamp 0
transform 1 0 3470 0 1 3610
box -6 -8 106 248
use NAND2X1  _3931_
timestamp 0
transform 1 0 3490 0 -1 3610
box -6 -8 86 248
use AOI22X1  _3932_
timestamp 0
transform 1 0 2370 0 1 3610
box -6 -8 126 248
use NAND3X1  _3933_
timestamp 0
transform 1 0 3270 0 1 3610
box -6 -8 106 248
use OAI21X1  _3934_
timestamp 0
transform -1 0 4590 0 1 4090
box -6 -8 106 248
use INVX1  _3935_
timestamp 0
transform 1 0 3870 0 1 8410
box -6 -8 66 248
use NAND3X1  _3936_
timestamp 0
transform 1 0 3670 0 1 8410
box -6 -8 106 248
use AOI22X1  _3937_
timestamp 0
transform 1 0 4250 0 -1 7450
box -6 -8 126 248
use OAI21X1  _3938_
timestamp 0
transform -1 0 3610 0 1 8890
box -6 -8 106 248
use NAND2X1  _3939_
timestamp 0
transform 1 0 3630 0 -1 8890
box -6 -8 86 248
use INVX1  _3940_
timestamp 0
transform -1 0 4810 0 -1 4090
box -6 -8 66 248
use OAI22X1  _3941_
timestamp 0
transform 1 0 6970 0 1 6010
box -6 -8 126 248
use NAND3X1  _3942_
timestamp 0
transform -1 0 10130 0 1 6970
box -6 -8 106 248
use NOR2X1  _3943_
timestamp 0
transform -1 0 10090 0 -1 7450
box -6 -8 86 248
use OAI21X1  _3944_
timestamp 0
transform -1 0 9810 0 1 7450
box -6 -8 106 248
use AND2X2  _3945_
timestamp 0
transform -1 0 10330 0 1 6970
box -6 -8 106 248
use NOR2X1  _3946_
timestamp 0
transform 1 0 9830 0 -1 7450
box -6 -8 86 248
use NOR2X1  _3947_
timestamp 0
transform 1 0 10430 0 1 6970
box -6 -8 86 248
use OAI21X1  _3948_
timestamp 0
transform 1 0 10610 0 1 6970
box -6 -8 106 248
use INVX2  _3949_
timestamp 0
transform 1 0 7730 0 1 7930
box -6 -8 66 248
use OAI21X1  _3950_
timestamp 0
transform -1 0 7090 0 1 5530
box -6 -8 106 248
use AOI21X1  _3951_
timestamp 0
transform 1 0 6590 0 -1 5530
box -6 -8 106 248
use OAI21X1  _3952_
timestamp 0
transform -1 0 5910 0 -1 5530
box -6 -8 106 248
use OAI21X1  _3953_
timestamp 0
transform 1 0 5490 0 -1 6490
box -6 -8 106 248
use INVX1  _3954_
timestamp 0
transform -1 0 5930 0 -1 6490
box -6 -8 66 248
use OAI21X1  _3955_
timestamp 0
transform 1 0 5950 0 1 6490
box -6 -8 106 248
use NOR2X1  _3956_
timestamp 0
transform -1 0 6230 0 1 6490
box -6 -8 86 248
use OAI21X1  _3957_
timestamp 0
transform 1 0 6190 0 -1 6490
box -6 -8 106 248
use NOR2X1  _3958_
timestamp 0
transform 1 0 6390 0 -1 6490
box -6 -8 86 248
use OAI21X1  _3959_
timestamp 0
transform 1 0 6510 0 1 6490
box -6 -8 106 248
use OAI21X1  _3960_
timestamp 0
transform 1 0 2430 0 -1 6010
box -6 -8 106 248
use INVX1  _3961_
timestamp 0
transform -1 0 2870 0 -1 6010
box -6 -8 66 248
use OAI21X1  _3962_
timestamp 0
transform 1 0 2970 0 1 6010
box -6 -8 106 248
use AND2X2  _3963_
timestamp 0
transform 1 0 3570 0 1 6010
box -6 -8 106 248
use AOI21X1  _3964_
timestamp 0
transform -1 0 4230 0 1 6010
box -6 -8 106 248
use OAI21X1  _3965_
timestamp 0
transform -1 0 3470 0 1 6010
box -6 -8 106 248
use NAND3X1  _3966_
timestamp 0
transform -1 0 4430 0 -1 6010
box -6 -8 106 248
use AOI21X1  _3967_
timestamp 0
transform -1 0 5230 0 1 6010
box -6 -8 106 248
use OAI21X1  _3968_
timestamp 0
transform -1 0 5430 0 1 6010
box -6 -8 106 248
use OAI21X1  _3969_
timestamp 0
transform -1 0 4430 0 1 6010
box -6 -8 106 248
use NAND2X1  _3970_
timestamp 0
transform 1 0 3970 0 -1 6010
box -6 -8 86 248
use INVX8  _3971_
timestamp 0
transform 1 0 5650 0 1 3610
box -6 -8 126 248
use AOI21X1  _3972_
timestamp 0
transform 1 0 5490 0 -1 4090
box -6 -8 106 248
use OAI21X1  _3973_
timestamp 0
transform 1 0 5490 0 1 5530
box -6 -8 106 248
use AOI21X1  _3974_
timestamp 0
transform -1 0 5790 0 1 5530
box -6 -8 106 248
use OAI21X1  _3975_
timestamp 0
transform -1 0 5790 0 -1 6010
box -6 -8 106 248
use AOI21X1  _3976_
timestamp 0
transform -1 0 5790 0 1 6010
box -6 -8 106 248
use OAI21X1  _3977_
timestamp 0
transform 1 0 5590 0 1 6490
box -6 -8 106 248
use NAND2X1  _3978_
timestamp 0
transform 1 0 6410 0 1 6010
box -6 -8 86 248
use INVX1  _3979_
timestamp 0
transform -1 0 2810 0 -1 6490
box -6 -8 66 248
use NAND3X1  _3980_
timestamp 0
transform 1 0 2070 0 -1 3610
box -6 -8 106 248
use NAND2X1  _3981_
timestamp 0
transform 1 0 1910 0 1 3130
box -6 -8 86 248
use AOI22X1  _3982_
timestamp 0
transform 1 0 1850 0 -1 3610
box -6 -8 126 248
use NAND3X1  _3983_
timestamp 0
transform -1 0 2070 0 1 3610
box -6 -8 106 248
use INVX8  _3984_
timestamp 0
transform 1 0 8310 0 1 4090
box -6 -8 126 248
use AOI21X1  _3985_
timestamp 0
transform 1 0 6890 0 -1 5050
box -6 -8 106 248
use OAI21X1  _3986_
timestamp 0
transform -1 0 7470 0 1 5530
box -6 -8 106 248
use INVX1  _3987_
timestamp 0
transform 1 0 7670 0 -1 6010
box -6 -8 66 248
use NAND2X1  _3988_
timestamp 0
transform 1 0 7590 0 1 6010
box -6 -8 86 248
use AOI21X1  _3989_
timestamp 0
transform 1 0 7390 0 1 6010
box -6 -8 106 248
use OAI21X1  _3990_
timestamp 0
transform 1 0 7190 0 1 6010
box -6 -8 106 248
use INVX1  _3991_
timestamp 0
transform -1 0 7370 0 -1 6010
box -6 -8 66 248
use AOI21X1  _3992_
timestamp 0
transform -1 0 8090 0 1 6010
box -6 -8 106 248
use OAI22X1  _3993_
timestamp 0
transform 1 0 7770 0 1 6010
box -6 -8 126 248
use INVX1  _3994_
timestamp 0
transform -1 0 7150 0 -1 5050
box -6 -8 66 248
use NOR2X1  _3995_
timestamp 0
transform -1 0 9530 0 1 6970
box -6 -8 86 248
use OAI21X1  _3996_
timestamp 0
transform -1 0 6150 0 1 6010
box -6 -8 106 248
use INVX1  _3997_
timestamp 0
transform 1 0 6030 0 -1 6490
box -6 -8 66 248
use OAI21X1  _3998_
timestamp 0
transform -1 0 6190 0 1 6970
box -6 -8 106 248
use AOI21X1  _3999_
timestamp 0
transform 1 0 5890 0 1 6970
box -6 -8 106 248
use OAI21X1  _4000_
timestamp 0
transform -1 0 5390 0 1 6970
box -6 -8 106 248
use NAND2X1  _4001_
timestamp 0
transform -1 0 5210 0 1 7450
box -6 -8 86 248
use INVX1  _4002_
timestamp 0
transform -1 0 7050 0 1 6970
box -6 -8 66 248
use INVX1  _4003_
timestamp 0
transform -1 0 6690 0 1 5530
box -6 -8 66 248
use NAND3X1  _4004_
timestamp 0
transform 1 0 2690 0 1 4570
box -6 -8 106 248
use NAND2X1  _4005_
timestamp 0
transform 1 0 2890 0 1 4570
box -6 -8 86 248
use AOI22X1  _4006_
timestamp 0
transform -1 0 2810 0 -1 4570
box -6 -8 126 248
use NAND3X1  _4007_
timestamp 0
transform 1 0 2490 0 1 4570
box -6 -8 106 248
use OAI21X1  _4008_
timestamp 0
transform -1 0 7250 0 -1 5530
box -6 -8 106 248
use AOI21X1  _4009_
timestamp 0
transform 1 0 6950 0 -1 5530
box -6 -8 106 248
use OAI21X1  _4010_
timestamp 0
transform -1 0 6890 0 1 5530
box -6 -8 106 248
use NOR2X1  _4011_
timestamp 0
transform 1 0 8670 0 -1 7930
box -6 -8 86 248
use INVX1  _4012_
timestamp 0
transform 1 0 6790 0 -1 5530
box -6 -8 66 248
use NOR2X1  _4013_
timestamp 0
transform 1 0 6670 0 -1 8890
box -6 -8 86 248
use OAI21X1  _4014_
timestamp 0
transform 1 0 6210 0 -1 9370
box -6 -8 106 248
use NOR2X1  _4015_
timestamp 0
transform 1 0 6570 0 -1 9370
box -6 -8 86 248
use NAND3X1  _4016_
timestamp 0
transform 1 0 9390 0 -1 9370
box -6 -8 106 248
use NOR2X1  _4017_
timestamp 0
transform -1 0 9770 0 1 9850
box -6 -8 86 248
use NOR2X1  _4018_
timestamp 0
transform -1 0 9950 0 1 9850
box -6 -8 86 248
use NAND2X1  _4019_
timestamp 0
transform 1 0 10050 0 1 9850
box -6 -8 86 248
use OR2X2  _4020_
timestamp 0
transform -1 0 7610 0 1 9370
box -6 -8 106 248
use INVX1  _4021_
timestamp 0
transform -1 0 10130 0 1 9370
box -6 -8 66 248
use INVX1  _4022_
timestamp 0
transform -1 0 6910 0 -1 8890
box -6 -8 66 248
use NOR2X1  _4023_
timestamp 0
transform -1 0 7270 0 -1 8890
box -6 -8 86 248
use OAI21X1  _4024_
timestamp 0
transform 1 0 9010 0 -1 8890
box -6 -8 106 248
use INVX1  _4025_
timestamp 0
transform -1 0 7770 0 1 9370
box -6 -8 66 248
use NOR2X1  _4026_
timestamp 0
transform -1 0 7950 0 1 9370
box -6 -8 86 248
use INVX1  _4027_
timestamp 0
transform 1 0 8430 0 1 9370
box -6 -8 66 248
use NOR2X1  _4028_
timestamp 0
transform 1 0 7970 0 1 7450
box -6 -8 86 248
use INVX1  _4029_
timestamp 0
transform 1 0 11070 0 1 11770
box -6 -8 66 248
use NAND2X1  _4030_
timestamp 0
transform 1 0 10890 0 1 11770
box -6 -8 86 248
use OAI21X1  _4031_
timestamp 0
transform 1 0 9250 0 1 6970
box -6 -8 106 248
use AOI21X1  _4032_
timestamp 0
transform 1 0 8710 0 1 6970
box -6 -8 106 248
use INVX1  _4033_
timestamp 0
transform -1 0 9410 0 -1 6970
box -6 -8 66 248
use INVX1  _4034_
timestamp 0
transform 1 0 4030 0 -1 9370
box -6 -8 66 248
use OAI21X1  _4035_
timestamp 0
transform 1 0 9830 0 1 6970
box -6 -8 106 248
use INVX1  _4036_
timestamp 0
transform -1 0 9730 0 -1 7450
box -6 -8 66 248
use OAI21X1  _4037_
timestamp 0
transform -1 0 9290 0 1 7930
box -6 -8 106 248
use OAI21X1  _4038_
timestamp 0
transform -1 0 8250 0 1 7450
box -6 -8 106 248
use INVX1  _4039_
timestamp 0
transform -1 0 7150 0 -1 8410
box -6 -8 66 248
use NAND2X1  _4040_
timestamp 0
transform 1 0 12050 0 -1 7450
box -6 -8 86 248
use OAI21X1  _4041_
timestamp 0
transform 1 0 9330 0 1 7450
box -6 -8 106 248
use INVX8  _4042_
timestamp 0
transform -1 0 6150 0 1 3130
box -6 -8 126 248
use AOI21X1  _4043_
timestamp 0
transform 1 0 5370 0 1 4090
box -6 -8 106 248
use OAI21X1  _4044_
timestamp 0
transform -1 0 5530 0 -1 5050
box -6 -8 106 248
use INVX1  _4045_
timestamp 0
transform -1 0 5550 0 1 5050
box -6 -8 66 248
use NAND2X1  _4046_
timestamp 0
transform -1 0 5930 0 1 5050
box -6 -8 86 248
use AOI21X1  _4047_
timestamp 0
transform -1 0 6130 0 -1 5050
box -6 -8 106 248
use OAI22X1  _4048_
timestamp 0
transform -1 0 6150 0 1 5050
box -6 -8 126 248
use INVX2  _4049_
timestamp 0
transform 1 0 5530 0 1 6010
box -6 -8 66 248
use AOI21X1  _4050_
timestamp 0
transform -1 0 5390 0 1 5050
box -6 -8 106 248
use OAI22X1  _4051_
timestamp 0
transform 1 0 5630 0 1 5050
box -6 -8 126 248
use INVX1  _4052_
timestamp 0
transform -1 0 6310 0 -1 4090
box -6 -8 66 248
use NAND2X1  _4053_
timestamp 0
transform -1 0 8310 0 1 6490
box -6 -8 86 248
use NAND3X1  _4054_
timestamp 0
transform 1 0 3770 0 1 4090
box -6 -8 106 248
use NAND2X1  _4055_
timestamp 0
transform -1 0 3670 0 1 4090
box -6 -8 86 248
use AOI22X1  _4056_
timestamp 0
transform 1 0 2770 0 1 4090
box -6 -8 126 248
use NAND3X1  _4057_
timestamp 0
transform 1 0 3390 0 1 4090
box -6 -8 106 248
use INVX2  _4058_
timestamp 0
transform -1 0 7570 0 -1 6490
box -6 -8 66 248
use NAND3X1  _4059_
timestamp 0
transform 1 0 7390 0 1 7450
box -6 -8 106 248
use OAI21X1  _4060_
timestamp 0
transform -1 0 8150 0 1 7930
box -6 -8 106 248
use OAI21X1  _4061_
timestamp 0
transform -1 0 9090 0 1 7930
box -6 -8 106 248
use OAI21X1  _4062_
timestamp 0
transform -1 0 3270 0 1 6010
box -6 -8 106 248
use INVX1  _4063_
timestamp 0
transform 1 0 5110 0 -1 6490
box -6 -8 66 248
use NAND3X1  _4064_
timestamp 0
transform -1 0 5170 0 -1 7930
box -6 -8 106 248
use AOI22X1  _4065_
timestamp 0
transform 1 0 5310 0 -1 7450
box -6 -8 126 248
use NAND2X1  _4066_
timestamp 0
transform 1 0 4510 0 -1 7930
box -6 -8 86 248
use OAI21X1  _4067_
timestamp 0
transform -1 0 7230 0 1 7930
box -6 -8 106 248
use INVX1  _4068_
timestamp 0
transform 1 0 3170 0 1 5530
box -6 -8 66 248
use NAND3X1  _4069_
timestamp 0
transform -1 0 790 0 1 3610
box -6 -8 106 248
use NAND2X1  _4070_
timestamp 0
transform 1 0 1190 0 -1 3610
box -6 -8 86 248
use AOI22X1  _4071_
timestamp 0
transform 1 0 570 0 -1 3610
box -6 -8 126 248
use NAND3X1  _4072_
timestamp 0
transform -1 0 990 0 1 3610
box -6 -8 106 248
use OAI21X1  _4073_
timestamp 0
transform 1 0 4130 0 1 4090
box -6 -8 106 248
use INVX1  _4074_
timestamp 0
transform 1 0 4330 0 1 4090
box -6 -8 66 248
use OAI21X1  _4075_
timestamp 0
transform 1 0 4250 0 1 6490
box -6 -8 106 248
use AOI21X1  _4076_
timestamp 0
transform -1 0 5590 0 1 6970
box -6 -8 106 248
use OAI21X1  _4077_
timestamp 0
transform 1 0 5530 0 -1 7450
box -6 -8 106 248
use NAND2X1  _4078_
timestamp 0
transform -1 0 5610 0 1 7450
box -6 -8 86 248
use OAI21X1  _4079_
timestamp 0
transform 1 0 3810 0 -1 8890
box -6 -8 106 248
use INVX1  _4080_
timestamp 0
transform 1 0 5910 0 -1 7450
box -6 -8 66 248
use INVX1  _4081_
timestamp 0
transform 1 0 950 0 1 7930
box -6 -8 66 248
use OAI21X1  _4082_
timestamp 0
transform 1 0 4190 0 -1 8890
box -6 -8 106 248
use INVX1  _4083_
timestamp 0
transform -1 0 4030 0 1 4090
box -6 -8 66 248
use NAND3X1  _4084_
timestamp 0
transform 1 0 1690 0 1 4090
box -6 -8 106 248
use NAND2X1  _4085_
timestamp 0
transform 1 0 1510 0 1 4090
box -6 -8 86 248
use AOI22X1  _4086_
timestamp 0
transform 1 0 1650 0 -1 4090
box -6 -8 126 248
use NAND3X1  _4087_
timestamp 0
transform 1 0 1610 0 -1 4570
box -6 -8 106 248
use OAI21X1  _4088_
timestamp 0
transform -1 0 4630 0 -1 6010
box -6 -8 106 248
use AND2X2  _4089_
timestamp 0
transform -1 0 4590 0 1 6970
box -6 -8 106 248
use AOI21X1  _4090_
timestamp 0
transform -1 0 4090 0 1 7450
box -6 -8 106 248
use OAI22X1  _4091_
timestamp 0
transform -1 0 3530 0 -1 8890
box -6 -8 126 248
use OAI21X1  _4092_
timestamp 0
transform -1 0 5810 0 1 7450
box -6 -8 106 248
use AOI22X1  _4093_
timestamp 0
transform 1 0 4670 0 -1 7450
box -6 -8 126 248
use INVX1  _4094_
timestamp 0
transform 1 0 4250 0 1 5530
box -6 -8 66 248
use NAND3X1  _4095_
timestamp 0
transform 1 0 1990 0 -1 5530
box -6 -8 106 248
use NAND2X1  _4096_
timestamp 0
transform 1 0 1810 0 -1 5530
box -6 -8 86 248
use AOI22X1  _4097_
timestamp 0
transform 1 0 1690 0 1 5050
box -6 -8 126 248
use NAND3X1  _4098_
timestamp 0
transform 1 0 1610 0 -1 5530
box -6 -8 106 248
use OAI21X1  _4099_
timestamp 0
transform 1 0 7190 0 1 7450
box -6 -8 106 248
use INVX1  _4100_
timestamp 0
transform 1 0 8070 0 -1 7450
box -6 -8 66 248
use NAND2X1  _4101_
timestamp 0
transform 1 0 8230 0 -1 7450
box -6 -8 86 248
use NOR2X1  _4102_
timestamp 0
transform -1 0 8490 0 -1 7450
box -6 -8 86 248
use OAI21X1  _4103_
timestamp 0
transform 1 0 8050 0 -1 7930
box -6 -8 106 248
use INVX1  _4104_
timestamp 0
transform -1 0 8310 0 -1 7930
box -6 -8 66 248
use OAI21X1  _4105_
timestamp 0
transform 1 0 8710 0 1 8410
box -6 -8 106 248
use INVX1  _4106_
timestamp 0
transform 1 0 6750 0 -1 7450
box -6 -8 66 248
use INVX1  _4107_
timestamp 0
transform -1 0 1190 0 -1 2650
box -6 -8 66 248
use INVX1  _4108_
timestamp 0
transform -1 0 590 0 1 2650
box -6 -8 66 248
use OAI21X1  _4109_
timestamp 0
transform -1 0 1970 0 1 9850
box -6 -8 106 248
use OAI21X1  _4110_
timestamp 0
transform -1 0 7910 0 1 9850
box -6 -8 106 248
use NOR2X1  _4111_
timestamp 0
transform -1 0 9610 0 -1 10330
box -6 -8 86 248
use OAI21X1  _4112_
timestamp 0
transform 1 0 2950 0 -1 3610
box -6 -8 106 248
use OAI21X1  _4113_
timestamp 0
transform 1 0 3150 0 -1 3610
box -6 -8 106 248
use NOR2X1  _4114_
timestamp 0
transform 1 0 3650 0 1 7930
box -6 -8 86 248
use OAI21X1  _4115_
timestamp 0
transform 1 0 4530 0 -1 10330
box -6 -8 106 248
use OAI21X1  _4116_
timestamp 0
transform -1 0 5490 0 -1 10330
box -6 -8 106 248
use OAI22X1  _4117_
timestamp 0
transform 1 0 4950 0 1 8410
box -6 -8 126 248
use NAND2X1  _4118_
timestamp 0
transform 1 0 4870 0 -1 8890
box -6 -8 86 248
use NAND3X1  _4119_
timestamp 0
transform 1 0 4030 0 1 8890
box -6 -8 106 248
use NOR2X1  _4120_
timestamp 0
transform -1 0 3830 0 -1 9850
box -6 -8 86 248
use INVX1  _4121_
timestamp 0
transform -1 0 4650 0 1 8410
box -6 -8 66 248
use OAI21X1  _4122_
timestamp 0
transform 1 0 4750 0 1 8410
box -6 -8 106 248
use INVX1  _4123_
timestamp 0
transform 1 0 8110 0 -1 8890
box -6 -8 66 248
use NAND2X1  _4124_
timestamp 0
transform 1 0 8630 0 -1 8890
box -6 -8 86 248
use OAI21X1  _4125_
timestamp 0
transform -1 0 4430 0 -1 10330
box -6 -8 106 248
use NAND2X1  _4126_
timestamp 0
transform 1 0 4310 0 1 10330
box -6 -8 86 248
use OAI21X1  _4127_
timestamp 0
transform 1 0 4130 0 -1 10330
box -6 -8 106 248
use AOI21X1  _4128_
timestamp 0
transform 1 0 4550 0 1 9850
box -6 -8 106 248
use NAND3X1  _4129_
timestamp 0
transform -1 0 5050 0 -1 11290
box -6 -8 106 248
use INVX1  _4130_
timestamp 0
transform 1 0 6090 0 1 11290
box -6 -8 66 248
use OAI21X1  _4131_
timestamp 0
transform 1 0 4350 0 1 9850
box -6 -8 106 248
use NOR2X1  _4132_
timestamp 0
transform -1 0 4650 0 1 10810
box -6 -8 86 248
use AOI22X1  _4133_
timestamp 0
transform -1 0 2170 0 1 10330
box -6 -8 126 248
use AND2X2  _4134_
timestamp 0
transform 1 0 1850 0 1 10330
box -6 -8 106 248
use OAI21X1  _4135_
timestamp 0
transform -1 0 2290 0 -1 10810
box -6 -8 106 248
use NOR2X1  _4136_
timestamp 0
transform -1 0 2270 0 1 11290
box -6 -8 86 248
use INVX1  _4137_
timestamp 0
transform -1 0 2090 0 -1 10810
box -6 -8 66 248
use AOI21X1  _4138_
timestamp 0
transform -1 0 2370 0 -1 11290
box -6 -8 106 248
use NAND3X1  _4139_
timestamp 0
transform 1 0 2070 0 -1 11290
box -6 -8 106 248
use OAI21X1  _4140_
timestamp 0
transform -1 0 3170 0 -1 11290
box -6 -8 106 248
use NAND3X1  _4141_
timestamp 0
transform 1 0 1870 0 -1 11290
box -6 -8 106 248
use NAND3X1  _4142_
timestamp 0
transform 1 0 1670 0 -1 11290
box -6 -8 106 248
use NOR2X1  _4143_
timestamp 0
transform -1 0 1570 0 -1 11290
box -6 -8 86 248
use NOR2X1  _4144_
timestamp 0
transform 1 0 1650 0 1 11290
box -6 -8 86 248
use NAND2X1  _4145_
timestamp 0
transform -1 0 1190 0 1 11290
box -6 -8 86 248
use OAI21X1  _4146_
timestamp 0
transform 1 0 3150 0 1 11290
box -6 -8 106 248
use INVX1  _4147_
timestamp 0
transform -1 0 2130 0 1 9850
box -6 -8 66 248
use OAI21X1  _4148_
timestamp 0
transform -1 0 3350 0 1 9370
box -6 -8 106 248
use NAND2X1  _4149_
timestamp 0
transform 1 0 3250 0 1 10330
box -6 -8 86 248
use NOR2X1  _4150_
timestamp 0
transform 1 0 3250 0 1 11770
box -6 -8 86 248
use NAND2X1  _4151_
timestamp 0
transform 1 0 3770 0 1 11770
box -6 -8 86 248
use INVX1  _4152_
timestamp 0
transform -1 0 3770 0 1 8890
box -6 -8 66 248
use OAI21X1  _4153_
timestamp 0
transform -1 0 2190 0 1 4570
box -6 -8 106 248
use OAI21X1  _4154_
timestamp 0
transform -1 0 2390 0 1 4570
box -6 -8 106 248
use INVX2  _4155_
timestamp 0
transform 1 0 690 0 -1 5050
box -6 -8 66 248
use NOR2X1  _4156_
timestamp 0
transform 1 0 1050 0 -1 5050
box -6 -8 86 248
use OAI21X1  _4157_
timestamp 0
transform -1 0 6070 0 -1 9850
box -6 -8 106 248
use OAI21X1  _4158_
timestamp 0
transform 1 0 6150 0 1 9370
box -6 -8 106 248
use NAND2X1  _4159_
timestamp 0
transform 1 0 6350 0 1 9370
box -6 -8 86 248
use OAI21X1  _4160_
timestamp 0
transform 1 0 5430 0 -1 9370
box -6 -8 106 248
use NAND2X1  _4161_
timestamp 0
transform -1 0 5710 0 -1 9370
box -6 -8 86 248
use AOI21X1  _4162_
timestamp 0
transform 1 0 5230 0 -1 9370
box -6 -8 106 248
use NOR2X1  _4163_
timestamp 0
transform -1 0 5310 0 1 9370
box -6 -8 86 248
use NAND2X1  _4164_
timestamp 0
transform 1 0 5790 0 1 9370
box -6 -8 86 248
use OAI21X1  _4165_
timestamp 0
transform -1 0 5870 0 -1 9850
box -6 -8 106 248
use OAI21X1  _4166_
timestamp 0
transform 1 0 5810 0 -1 9370
box -6 -8 106 248
use INVX2  _4167_
timestamp 0
transform 1 0 6510 0 -1 8890
box -6 -8 66 248
use NOR2X1  _4168_
timestamp 0
transform -1 0 6010 0 1 9850
box -6 -8 86 248
use NAND2X1  _4169_
timestamp 0
transform 1 0 5750 0 1 9850
box -6 -8 86 248
use NOR2X1  _4170_
timestamp 0
transform 1 0 6150 0 1 8890
box -6 -8 86 248
use NAND3X1  _4171_
timestamp 0
transform 1 0 5550 0 1 8890
box -6 -8 106 248
use INVX1  _4172_
timestamp 0
transform 1 0 5190 0 -1 8890
box -6 -8 66 248
use INVX1  _4173_
timestamp 0
transform 1 0 3870 0 1 8890
box -6 -8 66 248
use INVX1  _4174_
timestamp 0
transform 1 0 5590 0 1 9850
box -6 -8 66 248
use NOR2X1  _4175_
timestamp 0
transform 1 0 5210 0 -1 10330
box -6 -8 86 248
use OAI22X1  _4176_
timestamp 0
transform -1 0 3490 0 -1 10330
box -6 -8 126 248
use NAND2X1  _4177_
timestamp 0
transform 1 0 3070 0 1 10330
box -6 -8 86 248
use AOI22X1  _4178_
timestamp 0
transform -1 0 2390 0 1 10330
box -6 -8 126 248
use AOI21X1  _4179_
timestamp 0
transform -1 0 2490 0 -1 10810
box -6 -8 106 248
use OAI21X1  _4180_
timestamp 0
transform 1 0 2870 0 -1 11290
box -6 -8 106 248
use OAI21X1  _4181_
timestamp 0
transform -1 0 2570 0 -1 11290
box -6 -8 106 248
use OAI21X1  _4182_
timestamp 0
transform 1 0 2330 0 1 10810
box -6 -8 106 248
use NAND2X1  _4183_
timestamp 0
transform -1 0 3370 0 1 10810
box -6 -8 86 248
use NOR2X1  _4184_
timestamp 0
transform 1 0 3470 0 -1 11290
box -6 -8 86 248
use OAI21X1  _4185_
timestamp 0
transform 1 0 2890 0 1 10810
box -6 -8 106 248
use INVX1  _4186_
timestamp 0
transform -1 0 2550 0 1 10330
box -6 -8 66 248
use OAI21X1  _4187_
timestamp 0
transform 1 0 4130 0 1 9370
box -6 -8 106 248
use NAND2X1  _4188_
timestamp 0
transform 1 0 4330 0 1 9370
box -6 -8 86 248
use OAI21X1  _4189_
timestamp 0
transform -1 0 4230 0 -1 4570
box -6 -8 106 248
use NAND2X1  _4190_
timestamp 0
transform -1 0 4030 0 -1 4570
box -6 -8 86 248
use NAND3X1  _4191_
timestamp 0
transform -1 0 3850 0 -1 5050
box -6 -8 106 248
use AOI21X1  _4192_
timestamp 0
transform -1 0 5330 0 -1 5050
box -6 -8 106 248
use OAI21X1  _4193_
timestamp 0
transform -1 0 5190 0 1 5050
box -6 -8 106 248
use NAND2X1  _4194_
timestamp 0
transform -1 0 4030 0 -1 5050
box -6 -8 86 248
use NAND2X1  _4195_
timestamp 0
transform 1 0 3510 0 1 5530
box -6 -8 86 248
use INVX1  _4196_
timestamp 0
transform 1 0 3810 0 -1 6010
box -6 -8 66 248
use AOI22X1  _4197_
timestamp 0
transform 1 0 1670 0 -1 10330
box -6 -8 126 248
use AOI21X1  _4198_
timestamp 0
transform -1 0 1870 0 1 11770
box -6 -8 106 248
use OAI21X1  _4199_
timestamp 0
transform -1 0 2070 0 1 11770
box -6 -8 106 248
use NAND2X1  _4200_
timestamp 0
transform -1 0 2450 0 1 11770
box -6 -8 86 248
use NOR2X1  _4201_
timestamp 0
transform -1 0 1670 0 1 11770
box -6 -8 86 248
use OAI21X1  _4202_
timestamp 0
transform -1 0 1570 0 -1 11770
box -6 -8 106 248
use NOR2X1  _4203_
timestamp 0
transform -1 0 1930 0 -1 11770
box -6 -8 86 248
use AND2X2  _4204_
timestamp 0
transform -1 0 2750 0 1 10330
box -6 -8 106 248
use OR2X2  _4205_
timestamp 0
transform 1 0 2670 0 -1 11290
box -6 -8 106 248
use OAI21X1  _4206_
timestamp 0
transform -1 0 8730 0 -1 6970
box -6 -8 106 248
use NAND2X1  _4207_
timestamp 0
transform -1 0 8050 0 -1 4090
box -6 -8 86 248
use INVX1  _4208_
timestamp 0
transform -1 0 6370 0 1 4090
box -6 -8 66 248
use AOI22X1  _4209_
timestamp 0
transform -1 0 430 0 1 6490
box -6 -8 126 248
use AOI21X1  _4210_
timestamp 0
transform 1 0 110 0 1 6490
box -6 -8 106 248
use NAND3X1  _4211_
timestamp 0
transform -1 0 190 0 -1 6970
box -6 -8 106 248
use NOR3X1  _4212_
timestamp 0
transform -1 0 670 0 -1 8410
box -6 -8 186 248
use NAND2X1  _4213_
timestamp 0
transform 1 0 970 0 -1 8410
box -6 -8 86 248
use AOI22X1  _4214_
timestamp 0
transform -1 0 1590 0 -1 7930
box -6 -8 126 248
use OAI21X1  _4215_
timestamp 0
transform 1 0 1470 0 1 7930
box -6 -8 106 248
use AOI21X1  _4216_
timestamp 0
transform -1 0 2150 0 1 7930
box -6 -8 106 248
use AOI21X1  _4217_
timestamp 0
transform -1 0 3130 0 1 7450
box -6 -8 106 248
use OAI21X1  _4218_
timestamp 0
transform -1 0 2350 0 1 7930
box -6 -8 106 248
use AOI21X1  _4219_
timestamp 0
transform 1 0 2350 0 -1 8410
box -6 -8 106 248
use OAI21X1  _4220_
timestamp 0
transform 1 0 2550 0 -1 8410
box -6 -8 106 248
use NAND2X1  _4221_
timestamp 0
transform -1 0 390 0 -1 8410
box -6 -8 86 248
use INVX1  _4222_
timestamp 0
transform -1 0 170 0 1 6970
box -6 -8 66 248
use INVX1  _4223_
timestamp 0
transform -1 0 550 0 -1 6490
box -6 -8 66 248
use NAND3X1  _4224_
timestamp 0
transform -1 0 590 0 -1 6970
box -6 -8 106 248
use NOR2X1  _4225_
timestamp 0
transform -1 0 550 0 1 6970
box -6 -8 86 248
use NAND3X1  _4226_
timestamp 0
transform 1 0 110 0 -1 7930
box -6 -8 106 248
use NOR3X1  _4227_
timestamp 0
transform -1 0 490 0 -1 7930
box -6 -8 186 248
use OAI22X1  _4228_
timestamp 0
transform -1 0 2570 0 -1 7930
box -6 -8 126 248
use OAI21X1  _4229_
timestamp 0
transform 1 0 2670 0 1 7450
box -6 -8 106 248
use INVX1  _4230_
timestamp 0
transform -1 0 2930 0 1 7450
box -6 -8 66 248
use OAI21X1  _4231_
timestamp 0
transform 1 0 3210 0 1 7450
box -6 -8 106 248
use AOI21X1  _4232_
timestamp 0
transform -1 0 3770 0 -1 7450
box -6 -8 106 248
use AND2X2  _4233_
timestamp 0
transform -1 0 2350 0 -1 7930
box -6 -8 106 248
use NAND3X1  _4234_
timestamp 0
transform -1 0 3210 0 -1 8410
box -6 -8 106 248
use AOI22X1  _4235_
timestamp 0
transform -1 0 3990 0 -1 8410
box -6 -8 126 248
use OAI21X1  _4236_
timestamp 0
transform 1 0 3970 0 -1 7930
box -6 -8 106 248
use NAND2X1  _4237_
timestamp 0
transform -1 0 4250 0 -1 7930
box -6 -8 86 248
use OAI21X1  _4238_
timestamp 0
transform 1 0 3510 0 -1 8410
box -6 -8 106 248
use AOI21X1  _4239_
timestamp 0
transform 1 0 2670 0 -1 7930
box -6 -8 106 248
use INVX2  _4240_
timestamp 0
transform 1 0 2310 0 -1 8890
box -6 -8 66 248
use NAND3X1  _4241_
timestamp 0
transform -1 0 2250 0 -1 6970
box -6 -8 106 248
use AOI22X1  _4242_
timestamp 0
transform 1 0 2350 0 -1 6970
box -6 -8 126 248
use AOI21X1  _4243_
timestamp 0
transform -1 0 4610 0 -1 6970
box -6 -8 106 248
use NAND3X1  _4244_
timestamp 0
transform -1 0 5610 0 -1 6970
box -6 -8 106 248
use NAND2X1  _4245_
timestamp 0
transform -1 0 6170 0 -1 6970
box -6 -8 86 248
use NAND2X1  _4246_
timestamp 0
transform -1 0 4290 0 1 7930
box -6 -8 86 248
use NAND2X1  _4247_
timestamp 0
transform 1 0 2630 0 1 7930
box -6 -8 86 248
use NAND2X1  _4248_
timestamp 0
transform -1 0 5770 0 -1 6490
box -6 -8 86 248
use NAND2X1  _4249_
timestamp 0
transform -1 0 2470 0 1 6970
box -6 -8 86 248
use AND2X2  _4250_
timestamp 0
transform -1 0 4410 0 -1 6970
box -6 -8 106 248
use AOI21X1  _4251_
timestamp 0
transform 1 0 5690 0 -1 6970
box -6 -8 106 248
use OAI21X1  _4252_
timestamp 0
transform -1 0 5990 0 -1 6970
box -6 -8 106 248
use OAI21X1  _4253_
timestamp 0
transform -1 0 3890 0 1 7450
box -6 -8 106 248
use NAND2X1  _4254_
timestamp 0
transform -1 0 2290 0 1 6970
box -6 -8 86 248
use OAI21X1  _4255_
timestamp 0
transform 1 0 2570 0 -1 6970
box -6 -8 106 248
use AOI21X1  _4256_
timestamp 0
transform -1 0 4010 0 1 6970
box -6 -8 106 248
use NAND3X1  _4257_
timestamp 0
transform 1 0 4110 0 1 6970
box -6 -8 106 248
use NAND2X1  _4258_
timestamp 0
transform 1 0 4310 0 1 6970
box -6 -8 86 248
use NAND2X1  _4259_
timestamp 0
transform 1 0 4070 0 -1 7450
box -6 -8 86 248
use INVX1  _4260_
timestamp 0
transform -1 0 3070 0 1 7930
box -6 -8 66 248
use NAND2X1  _4261_
timestamp 0
transform -1 0 4150 0 1 5530
box -6 -8 86 248
use INVX2  _4262_
timestamp 0
transform 1 0 1610 0 -1 6010
box -6 -8 66 248
use AOI22X1  _4263_
timestamp 0
transform -1 0 8130 0 -1 6970
box -6 -8 126 248
use AND2X2  _4264_
timestamp 0
transform 1 0 7650 0 1 6490
box -6 -8 106 248
use AOI21X1  _4265_
timestamp 0
transform 1 0 7470 0 -1 6010
box -6 -8 106 248
use NOR2X1  _4266_
timestamp 0
transform 1 0 7150 0 -1 6010
box -6 -8 86 248
use OAI21X1  _4267_
timestamp 0
transform 1 0 7590 0 1 7450
box -6 -8 106 248
use NAND2X1  _4268_
timestamp 0
transform -1 0 6890 0 1 6970
box -6 -8 86 248
use NOR2X1  _4269_
timestamp 0
transform -1 0 9570 0 -1 7450
box -6 -8 86 248
use NAND3X1  _4270_
timestamp 0
transform -1 0 11290 0 1 7450
box -6 -8 106 248
use NAND2X1  _4271_
timestamp 0
transform 1 0 11170 0 1 8890
box -6 -8 86 248
use OAI21X1  _4272_
timestamp 0
transform 1 0 9290 0 -1 7450
box -6 -8 106 248
use NAND2X1  _4273_
timestamp 0
transform 1 0 9090 0 1 6970
box -6 -8 86 248
use NAND2X1  _4274_
timestamp 0
transform -1 0 9070 0 -1 6970
box -6 -8 86 248
use INVX1  _4275_
timestamp 0
transform 1 0 8830 0 -1 6970
box -6 -8 66 248
use NAND2X1  _4276_
timestamp 0
transform 1 0 8910 0 1 6970
box -6 -8 86 248
use INVX1  _4277_
timestamp 0
transform 1 0 8930 0 -1 7450
box -6 -8 66 248
use NOR2X1  _4278_
timestamp 0
transform 1 0 7810 0 1 8410
box -6 -8 86 248
use NAND3X1  _4279_
timestamp 0
transform 1 0 10590 0 1 9370
box -6 -8 106 248
use NAND2X1  _4280_
timestamp 0
transform 1 0 10790 0 1 9370
box -6 -8 86 248
use NAND2X1  _4281_
timestamp 0
transform -1 0 10810 0 -1 9370
box -6 -8 86 248
use AND2X2  _4282_
timestamp 0
transform -1 0 1370 0 -1 7930
box -6 -8 106 248
use AOI21X1  _4283_
timestamp 0
transform -1 0 7210 0 -1 7450
box -6 -8 106 248
use OAI21X1  _4284_
timestamp 0
transform 1 0 7710 0 -1 7450
box -6 -8 106 248
use AOI21X1  _4285_
timestamp 0
transform 1 0 7450 0 1 6490
box -6 -8 106 248
use OAI21X1  _4286_
timestamp 0
transform -1 0 1210 0 1 7930
box -6 -8 106 248
use INVX1  _4287_
timestamp 0
transform -1 0 1370 0 1 7930
box -6 -8 66 248
use OAI21X1  _4288_
timestamp 0
transform -1 0 1810 0 1 7450
box -6 -8 106 248
use AOI21X1  _4289_
timestamp 0
transform -1 0 4510 0 1 7450
box -6 -8 106 248
use OAI21X1  _4290_
timestamp 0
transform 1 0 6910 0 -1 7450
box -6 -8 106 248
use AOI21X1  _4291_
timestamp 0
transform 1 0 6910 0 1 6490
box -6 -8 106 248
use INVX2  _4292_
timestamp 0
transform -1 0 2630 0 1 6970
box -6 -8 66 248
use OAI21X1  _4293_
timestamp 0
transform -1 0 1950 0 1 7930
box -6 -8 106 248
use AOI21X1  _4294_
timestamp 0
transform -1 0 7430 0 1 7930
box -6 -8 106 248
use INVX1  _4295_
timestamp 0
transform 1 0 1550 0 1 7450
box -6 -8 66 248
use AND2X2  _4296_
timestamp 0
transform -1 0 210 0 -1 8410
box -6 -8 106 248
use AOI22X1  _4297_
timestamp 0
transform 1 0 1210 0 1 8410
box -6 -8 126 248
use AOI21X1  _4298_
timestamp 0
transform -1 0 3410 0 -1 8410
box -6 -8 106 248
use NAND2X1  _4299_
timestamp 0
transform 1 0 3410 0 1 7450
box -6 -8 86 248
use OAI21X1  _4300_
timestamp 0
transform -1 0 3970 0 -1 7450
box -6 -8 106 248
use AOI21X1  _4301_
timestamp 0
transform -1 0 3690 0 1 7450
box -6 -8 106 248
use INVX1  _4302_
timestamp 0
transform -1 0 3770 0 -1 8410
box -6 -8 66 248
use OAI21X1  _4303_
timestamp 0
transform -1 0 1730 0 1 8410
box -6 -8 106 248
use NAND2X1  _4304_
timestamp 0
transform 1 0 1230 0 -1 9370
box -6 -8 86 248
use AOI21X1  _4305_
timestamp 0
transform -1 0 2430 0 1 8410
box -6 -8 106 248
use NAND3X1  _4306_
timestamp 0
transform -1 0 2990 0 1 8410
box -6 -8 106 248
use AOI21X1  _4307_
timestamp 0
transform 1 0 6270 0 -1 6970
box -6 -8 106 248
use NOR2X1  _4308_
timestamp 0
transform -1 0 6410 0 1 6490
box -6 -8 86 248
use INVX1  _4309_
timestamp 0
transform 1 0 2910 0 -1 6490
box -6 -8 66 248
use OAI21X1  _4310_
timestamp 0
transform -1 0 2570 0 -1 8890
box -6 -8 106 248
use AOI21X1  _4311_
timestamp 0
transform 1 0 2370 0 1 8890
box -6 -8 106 248
use INVX2  _4312_
timestamp 0
transform 1 0 970 0 1 9370
box -6 -8 66 248
use AOI22X1  _4313_
timestamp 0
transform 1 0 1550 0 -1 8410
box -6 -8 126 248
use NAND2X1  _4314_
timestamp 0
transform 1 0 1730 0 1 8890
box -6 -8 86 248
use NOR2X1  _4315_
timestamp 0
transform -1 0 2830 0 -1 8410
box -6 -8 86 248
use NAND3X1  _4316_
timestamp 0
transform -1 0 2910 0 1 7930
box -6 -8 106 248
use AOI21X1  _4317_
timestamp 0
transform 1 0 4470 0 -1 7450
box -6 -8 106 248
use NOR2X1  _4318_
timestamp 0
transform 1 0 4150 0 -1 6010
box -6 -8 86 248
use INVX1  _4319_
timestamp 0
transform 1 0 3650 0 -1 6010
box -6 -8 66 248
use OAI21X1  _4320_
timestamp 0
transform -1 0 3170 0 -1 7930
box -6 -8 106 248
use AOI21X1  _4321_
timestamp 0
transform 1 0 2870 0 -1 7930
box -6 -8 106 248
use INVX1  _4322_
timestamp 0
transform 1 0 1610 0 -1 9370
box -6 -8 66 248
use NOR2X1  _4323_
timestamp 0
transform -1 0 2790 0 1 8410
box -6 -8 86 248
use AOI21X1  _4324_
timestamp 0
transform -1 0 1950 0 -1 7930
box -6 -8 106 248
use NAND3X1  _4325_
timestamp 0
transform -1 0 4210 0 -1 6970
box -6 -8 106 248
use AOI22X1  _4326_
timestamp 0
transform 1 0 4030 0 1 6490
box -6 -8 126 248
use NAND2X1  _4327_
timestamp 0
transform 1 0 4170 0 -1 6490
box -6 -8 86 248
use INVX2  _4328_
timestamp 0
transform -1 0 8650 0 -1 7450
box -6 -8 66 248
use OAI21X1  _4329_
timestamp 0
transform 1 0 1770 0 -1 8410
box -6 -8 106 248
use NOR2X1  _4330_
timestamp 0
transform 1 0 2170 0 -1 8410
box -6 -8 86 248
use OAI21X1  _4331_
timestamp 0
transform -1 0 1550 0 1 6970
box -6 -8 106 248
use OAI21X1  _4332_
timestamp 0
transform -1 0 2110 0 1 6970
box -6 -8 106 248
use AOI21X1  _4333_
timestamp 0
transform -1 0 3030 0 1 6970
box -6 -8 106 248
use NAND3X1  _4334_
timestamp 0
transform -1 0 3230 0 1 6970
box -6 -8 106 248
use AOI21X1  _4335_
timestamp 0
transform -1 0 3810 0 1 6970
box -6 -8 106 248
use OAI21X1  _4336_
timestamp 0
transform 1 0 2890 0 -1 7450
box -6 -8 106 248
use AOI21X1  _4337_
timestamp 0
transform 1 0 2690 0 -1 7450
box -6 -8 106 248
use OAI21X1  _4338_
timestamp 0
transform 1 0 2730 0 1 6970
box -6 -8 106 248
use NOR2X1  _4339_
timestamp 0
transform -1 0 3410 0 1 6970
box -6 -8 86 248
use OAI21X1  _4340_
timestamp 0
transform -1 0 3610 0 1 6970
box -6 -8 106 248
use OAI21X1  _4341_
timestamp 0
transform 1 0 3470 0 -1 7450
box -6 -8 106 248
use AOI21X1  _4342_
timestamp 0
transform -1 0 3370 0 -1 7450
box -6 -8 106 248
use OAI21X1  _4343_
timestamp 0
transform 1 0 3530 0 -1 6970
box -6 -8 106 248
use NOR2X1  _4344_
timestamp 0
transform 1 0 1830 0 1 6970
box -6 -8 86 248
use NAND2X1  _4345_
timestamp 0
transform -1 0 2530 0 1 7930
box -6 -8 86 248
use NOR2X1  _4346_
timestamp 0
transform 1 0 6950 0 1 7930
box -6 -8 86 248
use OAI21X1  _4347_
timestamp 0
transform -1 0 6850 0 1 7930
box -6 -8 106 248
use INVX1  _4348_
timestamp 0
transform -1 0 710 0 -1 6490
box -6 -8 66 248
use NOR2X1  _4349_
timestamp 0
transform -1 0 1150 0 1 6490
box -6 -8 86 248
use OAI21X1  _4350_
timestamp 0
transform 1 0 2210 0 1 6490
box -6 -8 106 248
use AND2X2  _4351_
timestamp 0
transform -1 0 2890 0 1 6490
box -6 -8 106 248
use AOI22X1  _4352_
timestamp 0
transform 1 0 3810 0 1 6490
box -6 -8 126 248
use NOR2X1  _4353_
timestamp 0
transform -1 0 6270 0 1 7930
box -6 -8 86 248
use NOR2X1  _4354_
timestamp 0
transform -1 0 3550 0 1 6490
box -6 -8 86 248
use NOR2X1  _4355_
timestamp 0
transform -1 0 970 0 1 6490
box -6 -8 86 248
use NOR2X1  _4356_
timestamp 0
transform -1 0 610 0 1 6490
box -6 -8 86 248
use OAI21X1  _4357_
timestamp 0
transform 1 0 2410 0 1 6490
box -6 -8 106 248
use NOR2X1  _4358_
timestamp 0
transform -1 0 5330 0 1 6490
box -6 -8 86 248
use OAI21X1  _4359_
timestamp 0
transform 1 0 5190 0 -1 5530
box -6 -8 106 248
use INVX1  _4360_
timestamp 0
transform -1 0 5190 0 1 5530
box -6 -8 66 248
use NOR2X1  _4361_
timestamp 0
transform 1 0 3090 0 -1 7450
box -6 -8 86 248
use INVX1  _4362_
timestamp 0
transform 1 0 4930 0 1 5050
box -6 -8 66 248
use NOR2X1  _4363_
timestamp 0
transform -1 0 4830 0 1 5050
box -6 -8 86 248
use INVX1  _4364_
timestamp 0
transform 1 0 3730 0 1 4570
box -6 -8 66 248
use OAI21X1  _4365_
timestamp 0
transform -1 0 5790 0 1 6970
box -6 -8 106 248
use INVX2  _4366_
timestamp 0
transform -1 0 5950 0 1 6010
box -6 -8 66 248
use NOR2X1  _4367_
timestamp 0
transform -1 0 3010 0 -1 8410
box -6 -8 86 248
use AOI22X1  _4368_
timestamp 0
transform 1 0 7590 0 1 8410
box -6 -8 126 248
use NOR2X1  _4369_
timestamp 0
transform -1 0 7490 0 1 8410
box -6 -8 86 248
use NOR2X1  _4370_
timestamp 0
transform 1 0 710 0 1 6490
box -6 -8 86 248
use INVX1  _4371_
timestamp 0
transform -1 0 1870 0 1 8410
box -6 -8 66 248
use OAI21X1  _4372_
timestamp 0
transform 1 0 1970 0 1 8410
box -6 -8 106 248
use INVX1  _4373_
timestamp 0
transform 1 0 2170 0 1 8410
box -6 -8 66 248
use NOR2X1  _4374_
timestamp 0
transform 1 0 2530 0 1 8410
box -6 -8 86 248
use NAND3X1  _4375_
timestamp 0
transform -1 0 3930 0 1 7930
box -6 -8 106 248
use OAI21X1  _4376_
timestamp 0
transform 1 0 7530 0 1 7930
box -6 -8 106 248
use NAND3X1  _4377_
timestamp 0
transform 1 0 11590 0 1 7450
box -6 -8 106 248
use INVX1  _4378_
timestamp 0
transform -1 0 1350 0 -1 6490
box -6 -8 66 248
use OAI22X1  _4379_
timestamp 0
transform -1 0 5370 0 1 10330
box -6 -8 126 248
use NAND2X1  _4380_
timestamp 0
transform 1 0 4850 0 1 10330
box -6 -8 86 248
use INVX1  _4381_
timestamp 0
transform 1 0 5950 0 1 10330
box -6 -8 66 248
use OAI22X1  _4382_
timestamp 0
transform 1 0 290 0 1 10330
box -6 -8 126 248
use NAND2X1  _4383_
timestamp 0
transform 1 0 110 0 1 10330
box -6 -8 86 248
use OAI21X1  _4384_
timestamp 0
transform 1 0 6290 0 -1 7930
box -6 -8 106 248
use NAND3X1  _4385_
timestamp 0
transform 1 0 6490 0 -1 7930
box -6 -8 106 248
use AOI21X1  _4386_
timestamp 0
transform 1 0 6890 0 -1 7930
box -6 -8 106 248
use OAI21X1  _4387_
timestamp 0
transform 1 0 6690 0 -1 7930
box -6 -8 106 248
use NAND2X1  _4388_
timestamp 0
transform -1 0 5550 0 -1 7930
box -6 -8 86 248
use NAND2X1  _4389_
timestamp 0
transform -1 0 6650 0 1 7930
box -6 -8 86 248
use AOI21X1  _4390_
timestamp 0
transform 1 0 7090 0 -1 7930
box -6 -8 106 248
use INVX1  _4391_
timestamp 0
transform 1 0 5030 0 -1 8890
box -6 -8 66 248
use AND2X2  _4392_
timestamp 0
transform -1 0 6470 0 1 7930
box -6 -8 106 248
use NAND2X1  _4393_
timestamp 0
transform 1 0 6550 0 -1 8410
box -6 -8 86 248
use NOR2X1  _4394_
timestamp 0
transform 1 0 6730 0 -1 8410
box -6 -8 86 248
use OAI21X1  _4395_
timestamp 0
transform 1 0 6850 0 1 8410
box -6 -8 106 248
use OAI21X1  _4396_
timestamp 0
transform -1 0 6410 0 -1 8890
box -6 -8 106 248
use AOI21X1  _4397_
timestamp 0
transform 1 0 4090 0 -1 8410
box -6 -8 106 248
use NAND2X1  _4398_
timestamp 0
transform 1 0 3070 0 1 4570
box -6 -8 86 248
use INVX2  _4399_
timestamp 0
transform 1 0 2190 0 -1 5530
box -6 -8 66 248
use OAI21X1  _4400_
timestamp 0
transform -1 0 6450 0 -1 8410
box -6 -8 106 248
use INVX1  _4401_
timestamp 0
transform 1 0 6290 0 1 8410
box -6 -8 66 248
use OAI21X1  _4402_
timestamp 0
transform -1 0 6210 0 -1 8890
box -6 -8 106 248
use INVX1  _4403_
timestamp 0
transform -1 0 5710 0 -1 7930
box -6 -8 66 248
use OAI21X1  _4404_
timestamp 0
transform 1 0 1450 0 -1 4090
box -6 -8 106 248
use OAI21X1  _4405_
timestamp 0
transform -1 0 1970 0 -1 4090
box -6 -8 106 248
use OAI21X1  _4406_
timestamp 0
transform -1 0 2670 0 1 4090
box -6 -8 106 248
use OAI21X1  _4407_
timestamp 0
transform -1 0 2470 0 1 4090
box -6 -8 106 248
use OAI21X1  _4408_
timestamp 0
transform 1 0 1610 0 -1 5050
box -6 -8 106 248
use OAI21X1  _4409_
timestamp 0
transform -1 0 1910 0 -1 5050
box -6 -8 106 248
use OAI21X1  _4410_
timestamp 0
transform 1 0 3630 0 1 10330
box -6 -8 106 248
use OAI21X1  _4411_
timestamp 0
transform 1 0 3930 0 -1 10330
box -6 -8 106 248
use INVX1  _4412_
timestamp 0
transform 1 0 1790 0 1 10810
box -6 -8 66 248
use AOI21X1  _4413_
timestamp 0
transform -1 0 390 0 1 4090
box -6 -8 106 248
use NOR2X1  _4414_
timestamp 0
transform 1 0 310 0 1 4570
box -6 -8 86 248
use INVX1  _4415_
timestamp 0
transform 1 0 490 0 1 4090
box -6 -8 66 248
use OAI21X1  _4416_
timestamp 0
transform 1 0 1570 0 1 3610
box -6 -8 106 248
use OAI21X1  _4417_
timestamp 0
transform -1 0 1870 0 1 3610
box -6 -8 106 248
use OAI21X1  _4418_
timestamp 0
transform -1 0 2690 0 1 3610
box -6 -8 106 248
use OAI21X1  _4419_
timestamp 0
transform 1 0 2170 0 1 3610
box -6 -8 106 248
use OAI21X1  _4420_
timestamp 0
transform 1 0 2290 0 -1 4570
box -6 -8 106 248
use OAI21X1  _4421_
timestamp 0
transform 1 0 2490 0 -1 4570
box -6 -8 106 248
use INVX2  _4422_
timestamp 0
transform -1 0 2070 0 -1 5050
box -6 -8 66 248
use NAND2X1  _4423_
timestamp 0
transform -1 0 730 0 1 4570
box -6 -8 86 248
use AND2X2  _4424_
timestamp 0
transform 1 0 2090 0 1 5050
box -6 -8 106 248
use OAI21X1  _4425_
timestamp 0
transform 1 0 1130 0 1 4090
box -6 -8 106 248
use NAND2X1  _4426_
timestamp 0
transform 1 0 1330 0 1 4090
box -6 -8 86 248
use OAI21X1  _4427_
timestamp 0
transform 1 0 3590 0 -1 4090
box -6 -8 106 248
use NAND2X1  _4428_
timestamp 0
transform -1 0 3490 0 -1 4090
box -6 -8 86 248
use OAI21X1  _4429_
timestamp 0
transform 1 0 1310 0 1 5050
box -6 -8 106 248
use NAND2X1  _4430_
timestamp 0
transform 1 0 1510 0 1 5050
box -6 -8 86 248
use AOI21X1  _4431_
timestamp 0
transform -1 0 850 0 -1 5530
box -6 -8 106 248
use NOR2X1  _4432_
timestamp 0
transform -1 0 730 0 1 5050
box -6 -8 86 248
use INVX1  _4433_
timestamp 0
transform -1 0 950 0 1 5530
box -6 -8 66 248
use OAI21X1  _4434_
timestamp 0
transform -1 0 1450 0 -1 3130
box -6 -8 106 248
use NAND2X1  _4435_
timestamp 0
transform 1 0 1550 0 -1 3130
box -6 -8 86 248
use OAI21X1  _4436_
timestamp 0
transform 1 0 3150 0 1 3130
box -6 -8 106 248
use NAND2X1  _4437_
timestamp 0
transform -1 0 3430 0 1 3130
box -6 -8 86 248
use OAI21X1  _4438_
timestamp 0
transform -1 0 6690 0 1 9850
box -6 -8 106 248
use OAI21X1  _4439_
timestamp 0
transform 1 0 6010 0 1 10810
box -6 -8 106 248
use NOR2X1  _4440_
timestamp 0
transform -1 0 4850 0 -1 11290
box -6 -8 86 248
use OAI21X1  _4441_
timestamp 0
transform 1 0 4190 0 1 10810
box -6 -8 106 248
use AOI21X1  _4442_
timestamp 0
transform 1 0 3970 0 -1 10810
box -6 -8 106 248
use INVX1  _4443_
timestamp 0
transform 1 0 3850 0 1 10810
box -6 -8 66 248
use NAND2X1  _4444_
timestamp 0
transform 1 0 3670 0 1 10810
box -6 -8 86 248
use NOR2X1  _4445_
timestamp 0
transform 1 0 4010 0 1 10810
box -6 -8 86 248
use NAND2X1  _4446_
timestamp 0
transform 1 0 4430 0 -1 11290
box -6 -8 86 248
use INVX1  _4447_
timestamp 0
transform 1 0 4610 0 -1 11290
box -6 -8 66 248
use INVX1  _4448_
timestamp 0
transform 1 0 2530 0 1 10810
box -6 -8 66 248
use NAND2X1  _4449_
timestamp 0
transform 1 0 1090 0 1 10810
box -6 -8 86 248
use AOI21X1  _4450_
timestamp 0
transform -1 0 1930 0 -1 10810
box -6 -8 106 248
use OAI21X1  _4451_
timestamp 0
transform 1 0 1430 0 -1 10810
box -6 -8 106 248
use INVX2  _4452_
timestamp 0
transform -1 0 2290 0 1 9370
box -6 -8 66 248
use INVX1  _4453_
timestamp 0
transform 1 0 7270 0 1 9850
box -6 -8 66 248
use AOI21X1  _4454_
timestamp 0
transform -1 0 1170 0 -1 4090
box -6 -8 106 248
use AOI22X1  _4455_
timestamp 0
transform 1 0 6810 0 -1 4090
box -6 -8 126 248
use NOR2X1  _4456_
timestamp 0
transform 1 0 7030 0 -1 4090
box -6 -8 86 248
use NOR2X1  _4457_
timestamp 0
transform 1 0 7230 0 1 4090
box -6 -8 86 248
use OR2X2  _4458_
timestamp 0
transform -1 0 7510 0 1 4090
box -6 -8 106 248
use OAI21X1  _4459_
timestamp 0
transform -1 0 7130 0 1 4090
box -6 -8 106 248
use NOR2X1  _4460_
timestamp 0
transform -1 0 8430 0 -1 4570
box -6 -8 86 248
use NOR2X1  _4461_
timestamp 0
transform 1 0 7650 0 -1 4570
box -6 -8 86 248
use INVX2  _4462_
timestamp 0
transform -1 0 6790 0 -1 5050
box -6 -8 66 248
use NOR2X1  _4463_
timestamp 0
transform 1 0 1270 0 -1 4090
box -6 -8 86 248
use AOI21X1  _4464_
timestamp 0
transform -1 0 2650 0 -1 4090
box -6 -8 106 248
use INVX1  _4465_
timestamp 0
transform -1 0 5950 0 -1 4090
box -6 -8 66 248
use OAI21X1  _4466_
timestamp 0
transform 1 0 6050 0 -1 4090
box -6 -8 106 248
use NAND3X1  _4467_
timestamp 0
transform 1 0 6470 0 1 4090
box -6 -8 106 248
use NAND3X1  _4468_
timestamp 0
transform 1 0 6710 0 -1 4570
box -6 -8 106 248
use INVX1  _4469_
timestamp 0
transform 1 0 6910 0 -1 4570
box -6 -8 66 248
use INVX1  _4470_
timestamp 0
transform -1 0 6710 0 1 6970
box -6 -8 66 248
use OAI21X1  _4471_
timestamp 0
transform 1 0 7250 0 -1 4570
box -6 -8 106 248
use NOR2X1  _4472_
timestamp 0
transform -1 0 6530 0 1 4570
box -6 -8 86 248
use INVX1  _4473_
timestamp 0
transform 1 0 8190 0 -1 4570
box -6 -8 66 248
use NAND2X1  _4474_
timestamp 0
transform -1 0 6350 0 1 4570
box -6 -8 86 248
use NOR2X1  _4475_
timestamp 0
transform 1 0 2750 0 -1 4090
box -6 -8 86 248
use AOI21X1  _4476_
timestamp 0
transform -1 0 1330 0 -1 5050
box -6 -8 106 248
use OAI21X1  _4477_
timestamp 0
transform -1 0 2730 0 1 5530
box -6 -8 106 248
use NAND2X1  _4478_
timestamp 0
transform 1 0 2630 0 -1 6010
box -6 -8 86 248
use INVX2  _4479_
timestamp 0
transform 1 0 5350 0 -1 6970
box -6 -8 66 248
use NOR2X1  _4480_
timestamp 0
transform 1 0 1430 0 -1 5050
box -6 -8 86 248
use OAI21X1  _4481_
timestamp 0
transform 1 0 270 0 1 5050
box -6 -8 106 248
use NAND2X1  _4482_
timestamp 0
transform 1 0 470 0 1 5050
box -6 -8 86 248
use OAI21X1  _4483_
timestamp 0
transform 1 0 3230 0 -1 5050
box -6 -8 106 248
use OAI21X1  _4484_
timestamp 0
transform -1 0 5070 0 1 4570
box -6 -8 106 248
use NOR2X1  _4485_
timestamp 0
transform 1 0 5370 0 1 4570
box -6 -8 86 248
use AND2X2  _4486_
timestamp 0
transform -1 0 5270 0 1 4570
box -6 -8 106 248
use NAND2X1  _4487_
timestamp 0
transform -1 0 5630 0 1 4570
box -6 -8 86 248
use NAND2X1  _4488_
timestamp 0
transform 1 0 5730 0 1 4570
box -6 -8 86 248
use OAI21X1  _4489_
timestamp 0
transform -1 0 5930 0 -1 5050
box -6 -8 106 248
use INVX1  _4490_
timestamp 0
transform -1 0 5850 0 1 6490
box -6 -8 66 248
use OAI21X1  _4491_
timestamp 0
transform -1 0 5950 0 -1 4570
box -6 -8 106 248
use INVX1  _4492_
timestamp 0
transform 1 0 110 0 1 5050
box -6 -8 66 248
use OAI21X1  _4493_
timestamp 0
transform -1 0 5810 0 -1 10810
box -6 -8 106 248
use NAND2X1  _4494_
timestamp 0
transform 1 0 5530 0 -1 10810
box -6 -8 86 248
use NOR2X1  _4495_
timestamp 0
transform 1 0 4390 0 1 10810
box -6 -8 86 248
use NAND2X1  _4496_
timestamp 0
transform 1 0 3850 0 -1 11290
box -6 -8 86 248
use NAND2X1  _4497_
timestamp 0
transform -1 0 3690 0 1 11770
box -6 -8 86 248
use NOR2X1  _4498_
timestamp 0
transform -1 0 4730 0 1 11290
box -6 -8 86 248
use OAI21X1  _4499_
timestamp 0
transform 1 0 1290 0 -1 11290
box -6 -8 106 248
use INVX1  _4500_
timestamp 0
transform 1 0 6390 0 -1 10810
box -6 -8 66 248
use OAI21X1  _4501_
timestamp 0
transform 1 0 6110 0 1 10330
box -6 -8 106 248
use NAND2X1  _4502_
timestamp 0
transform -1 0 4610 0 -1 10810
box -6 -8 86 248
use OAI21X1  _4503_
timestamp 0
transform 1 0 6510 0 1 10330
box -6 -8 106 248
use AOI21X1  _4504_
timestamp 0
transform -1 0 1830 0 -1 3130
box -6 -8 106 248
use INVX1  _4505_
timestamp 0
transform -1 0 4910 0 1 3610
box -6 -8 66 248
use AOI21X1  _4506_
timestamp 0
transform -1 0 5390 0 -1 4090
box -6 -8 106 248
use AOI21X1  _4507_
timestamp 0
transform 1 0 5690 0 -1 4090
box -6 -8 106 248
use OR2X2  _4508_
timestamp 0
transform 1 0 5570 0 1 4090
box -6 -8 106 248
use NAND2X1  _4509_
timestamp 0
transform -1 0 5850 0 1 4090
box -6 -8 86 248
use NAND2X1  _4510_
timestamp 0
transform -1 0 6030 0 1 4090
box -6 -8 86 248
use NAND2X1  _4511_
timestamp 0
transform 1 0 6130 0 1 4090
box -6 -8 86 248
use NAND2X1  _4512_
timestamp 0
transform 1 0 6210 0 -1 4570
box -6 -8 86 248
use INVX2  _4513_
timestamp 0
transform 1 0 6250 0 1 6010
box -6 -8 66 248
use NOR2X1  _4514_
timestamp 0
transform -1 0 1810 0 1 3130
box -6 -8 86 248
use AOI21X1  _4515_
timestamp 0
transform -1 0 2670 0 -1 3130
box -6 -8 106 248
use INVX1  _4516_
timestamp 0
transform -1 0 4750 0 -1 3610
box -6 -8 66 248
use OAI21X1  _4517_
timestamp 0
transform -1 0 5270 0 1 4090
box -6 -8 106 248
use OAI21X1  _4518_
timestamp 0
transform 1 0 5150 0 -1 4570
box -6 -8 106 248
use NOR2X1  _4519_
timestamp 0
transform 1 0 5510 0 -1 4570
box -6 -8 86 248
use NOR2X1  _4520_
timestamp 0
transform -1 0 5770 0 -1 4570
box -6 -8 86 248
use INVX1  _4521_
timestamp 0
transform 1 0 6550 0 -1 4570
box -6 -8 66 248
use AND2X2  _4522_
timestamp 0
transform -1 0 9050 0 1 7450
box -6 -8 106 248
use INVX1  _4523_
timestamp 0
transform 1 0 5350 0 -1 4570
box -6 -8 66 248
use NOR2X1  _4524_
timestamp 0
transform 1 0 6050 0 -1 4570
box -6 -8 86 248
use NOR2X1  _4525_
timestamp 0
transform 1 0 5910 0 1 4570
box -6 -8 86 248
use NAND2X1  _4526_
timestamp 0
transform -1 0 6550 0 1 6970
box -6 -8 86 248
use INVX1  _4527_
timestamp 0
transform -1 0 5030 0 1 7450
box -6 -8 66 248
use INVX1  _4528_
timestamp 0
transform 1 0 6390 0 -1 4570
box -6 -8 66 248
use NAND2X1  _4529_
timestamp 0
transform 1 0 6090 0 1 4570
box -6 -8 86 248
use AND2X2  _4530_
timestamp 0
transform 1 0 6070 0 -1 7450
box -6 -8 106 248
use NOR2X1  _4531_
timestamp 0
transform -1 0 2370 0 1 3130
box -6 -8 86 248
use OAI22X1  _4532_
timestamp 0
transform -1 0 6410 0 1 10330
box -6 -8 126 248
use NAND2X1  _4533_
timestamp 0
transform -1 0 6330 0 1 11290
box -6 -8 86 248
use NOR2X1  _4534_
timestamp 0
transform 1 0 4310 0 1 11770
box -6 -8 86 248
use NOR2X1  _4535_
timestamp 0
transform 1 0 3710 0 1 11290
box -6 -8 86 248
use NAND2X1  _4536_
timestamp 0
transform -1 0 1190 0 -1 11290
box -6 -8 86 248
use NAND2X1  _4537_
timestamp 0
transform 1 0 4490 0 1 10330
box -6 -8 86 248
use NOR2X1  _4538_
timestamp 0
transform -1 0 7790 0 1 11290
box -6 -8 86 248
use INVX2  _4539_
timestamp 0
transform -1 0 3150 0 1 11770
box -6 -8 66 248
use INVX4  _4540_
timestamp 0
transform 1 0 7690 0 -1 11290
box -6 -8 86 248
use INVX1  _4541_
timestamp 0
transform 1 0 6550 0 -1 10330
box -6 -8 66 248
use AOI21X1  _4542_
timestamp 0
transform 1 0 3090 0 -1 4570
box -6 -8 106 248
use NOR2X1  _4543_
timestamp 0
transform -1 0 2990 0 -1 4570
box -6 -8 86 248
use AND2X2  _4544_
timestamp 0
transform -1 0 1030 0 -1 4570
box -6 -8 106 248
use AOI22X1  _4545_
timestamp 0
transform 1 0 2170 0 -1 9370
box -6 -8 126 248
use NAND2X1  _4546_
timestamp 0
transform 1 0 2950 0 1 8890
box -6 -8 86 248
use OR2X2  _4547_
timestamp 0
transform -1 0 2490 0 -1 9370
box -6 -8 106 248
use OR2X2  _4548_
timestamp 0
transform -1 0 1870 0 -1 9370
box -6 -8 106 248
use OAI21X1  _4549_
timestamp 0
transform 1 0 2650 0 -1 5050
box -6 -8 106 248
use NAND2X1  _4550_
timestamp 0
transform 1 0 2850 0 -1 5050
box -6 -8 86 248
use OAI21X1  _4551_
timestamp 0
transform -1 0 3130 0 -1 5050
box -6 -8 106 248
use NAND2X1  _4552_
timestamp 0
transform -1 0 3070 0 1 5530
box -6 -8 86 248
use INVX1  _4553_
timestamp 0
transform -1 0 6630 0 -1 6490
box -6 -8 66 248
use NAND2X1  _4554_
timestamp 0
transform 1 0 1030 0 1 4570
box -6 -8 86 248
use INVX1  _4555_
timestamp 0
transform -1 0 830 0 -1 4570
box -6 -8 66 248
use OAI21X1  _4556_
timestamp 0
transform 1 0 4390 0 1 8410
box -6 -8 106 248
use NOR2X1  _4557_
timestamp 0
transform 1 0 4210 0 1 8410
box -6 -8 86 248
use NAND2X1  _4558_
timestamp 0
transform -1 0 4110 0 1 8410
box -6 -8 86 248
use INVX2  _4559_
timestamp 0
transform 1 0 5070 0 1 9370
box -6 -8 66 248
use NAND3X1  _4560_
timestamp 0
transform -1 0 8610 0 1 8410
box -6 -8 106 248
use OAI21X1  _4561_
timestamp 0
transform -1 0 9010 0 1 8410
box -6 -8 106 248
use NOR2X1  _4562_
timestamp 0
transform 1 0 8450 0 -1 8890
box -6 -8 86 248
use INVX1  _4563_
timestamp 0
transform -1 0 6470 0 -1 9370
box -6 -8 66 248
use NOR2X1  _4564_
timestamp 0
transform -1 0 1990 0 1 5050
box -6 -8 86 248
use OAI21X1  _4565_
timestamp 0
transform 1 0 2750 0 1 8890
box -6 -8 106 248
use AOI21X1  _4566_
timestamp 0
transform 1 0 3130 0 1 8890
box -6 -8 106 248
use NAND3X1  _4567_
timestamp 0
transform -1 0 6910 0 1 8890
box -6 -8 106 248
use OAI21X1  _4568_
timestamp 0
transform 1 0 6750 0 -1 9370
box -6 -8 106 248
use OAI21X1  _4569_
timestamp 0
transform 1 0 1970 0 -1 9370
box -6 -8 106 248
use NAND3X1  _4570_
timestamp 0
transform -1 0 6710 0 1 8890
box -6 -8 106 248
use NOR3X1  _4571_
timestamp 0
transform 1 0 6330 0 1 8890
box -6 -8 186 248
use NOR2X1  _4572_
timestamp 0
transform -1 0 9610 0 -1 8410
box -6 -8 86 248
use NAND3X1  _4573_
timestamp 0
transform -1 0 10510 0 -1 8410
box -6 -8 106 248
use NAND3X1  _4574_
timestamp 0
transform -1 0 9690 0 1 7930
box -6 -8 106 248
use INVX1  _4575_
timestamp 0
transform -1 0 7070 0 1 8890
box -6 -8 66 248
use NAND3X1  _4576_
timestamp 0
transform -1 0 8630 0 1 8890
box -6 -8 106 248
use AOI21X1  _4577_
timestamp 0
transform -1 0 3150 0 1 9370
box -6 -8 106 248
use OR2X2  _4578_
timestamp 0
transform -1 0 6110 0 -1 9370
box -6 -8 106 248
use OAI21X1  _4579_
timestamp 0
transform 1 0 8050 0 1 9370
box -6 -8 106 248
use NAND2X1  _4580_
timestamp 0
transform 1 0 10230 0 1 9370
box -6 -8 86 248
use OAI21X1  _4581_
timestamp 0
transform -1 0 7650 0 1 8890
box -6 -8 106 248
use INVX1  _4582_
timestamp 0
transform 1 0 1330 0 -1 10330
box -6 -8 66 248
use OAI21X1  _4583_
timestamp 0
transform -1 0 2490 0 1 9370
box -6 -8 106 248
use NAND2X1  _4584_
timestamp 0
transform -1 0 2310 0 1 9850
box -6 -8 86 248
use OAI21X1  _4585_
timestamp 0
transform -1 0 2230 0 1 10810
box -6 -8 106 248
use NAND2X1  _4586_
timestamp 0
transform -1 0 2030 0 1 10810
box -6 -8 86 248
use NOR2X1  _4587_
timestamp 0
transform -1 0 1690 0 1 10810
box -6 -8 86 248
use INVX1  _4588_
timestamp 0
transform 1 0 3350 0 1 11290
box -6 -8 66 248
use NOR2X1  _4589_
timestamp 0
transform 1 0 3890 0 1 11290
box -6 -8 86 248
use NAND2X1  _4590_
timestamp 0
transform 1 0 1270 0 1 10810
box -6 -8 86 248
use AOI21X1  _4591_
timestamp 0
transform -1 0 1770 0 1 9850
box -6 -8 106 248
use OAI21X1  _4592_
timestamp 0
transform 1 0 1470 0 1 9850
box -6 -8 106 248
use INVX2  _4593_
timestamp 0
transform -1 0 4090 0 1 5050
box -6 -8 66 248
use NAND2X1  _4594_
timestamp 0
transform -1 0 3270 0 -1 11770
box -6 -8 86 248
use AOI21X1  _4595_
timestamp 0
transform -1 0 2850 0 1 11290
box -6 -8 106 248
use OAI21X1  _4596_
timestamp 0
transform -1 0 3050 0 1 11290
box -6 -8 106 248
use INVX1  _4597_
timestamp 0
transform 1 0 2830 0 -1 11770
box -6 -8 66 248
use NOR2X1  _4598_
timestamp 0
transform -1 0 2810 0 1 11770
box -6 -8 86 248
use NAND2X1  _4599_
timestamp 0
transform -1 0 2990 0 1 11770
box -6 -8 86 248
use OR2X2  _4600_
timestamp 0
transform -1 0 4170 0 1 11290
box -6 -8 106 248
use NAND2X1  _4601_
timestamp 0
transform -1 0 4110 0 -1 11290
box -6 -8 86 248
use INVX1  _4602_
timestamp 0
transform -1 0 1510 0 1 10810
box -6 -8 66 248
use AND2X2  _4603_
timestamp 0
transform -1 0 1490 0 1 11770
box -6 -8 106 248
use NAND3X1  _4604_
timestamp 0
transform -1 0 3090 0 -1 11770
box -6 -8 106 248
use AND2X2  _4605_
timestamp 0
transform 1 0 1830 0 1 11290
box -6 -8 106 248
use OAI21X1  _4606_
timestamp 0
transform -1 0 810 0 -1 11290
box -6 -8 106 248
use NAND2X1  _4607_
timestamp 0
transform -1 0 610 0 -1 11290
box -6 -8 86 248
use MUX2X1  _4608_
timestamp 0
transform -1 0 3390 0 -1 7930
box -6 -8 126 248
use NAND2X1  _4609_
timestamp 0
transform 1 0 1670 0 -1 11770
box -6 -8 86 248
use OAI21X1  _4610_
timestamp 0
transform 1 0 2550 0 1 11290
box -6 -8 106 248
use NAND2X1  _4611_
timestamp 0
transform -1 0 2450 0 1 11290
box -6 -8 86 248
use NAND2X1  _4612_
timestamp 0
transform -1 0 2090 0 1 11290
box -6 -8 86 248
use AND2X2  _4613_
timestamp 0
transform 1 0 2030 0 -1 11770
box -6 -8 106 248
use OAI21X1  _4614_
timestamp 0
transform -1 0 770 0 1 11770
box -6 -8 106 248
use NAND2X1  _4615_
timestamp 0
transform -1 0 570 0 1 11770
box -6 -8 86 248
use OAI21X1  _4616_
timestamp 0
transform -1 0 1950 0 1 2650
box -6 -8 106 248
use OR2X2  _4617_
timestamp 0
transform -1 0 1750 0 1 2650
box -6 -8 106 248
use NAND2X1  _4618_
timestamp 0
transform -1 0 2630 0 1 11770
box -6 -8 86 248
use NOR2X1  _4619_
timestamp 0
transform -1 0 1970 0 -1 10330
box -6 -8 86 248
use NAND2X1  _4620_
timestamp 0
transform -1 0 1570 0 -1 10330
box -6 -8 86 248
use AOI21X1  _4621_
timestamp 0
transform 1 0 2170 0 1 11770
box -6 -8 106 248
use NOR2X1  _4622_
timestamp 0
transform 1 0 2590 0 -1 10810
box -6 -8 86 248
use MUX2X1  _4623_
timestamp 0
transform 1 0 2090 0 -1 9850
box -6 -8 126 248
use INVX2  _4624_
timestamp 0
transform 1 0 1290 0 -1 10810
box -6 -8 66 248
use OAI21X1  _4625_
timestamp 0
transform 1 0 910 0 1 11290
box -6 -8 106 248
use NAND2X1  _4626_
timestamp 0
transform -1 0 810 0 1 11290
box -6 -8 86 248
use NAND2X1  _4627_
timestamp 0
transform -1 0 2310 0 -1 11770
box -6 -8 86 248
use NAND2X1  _4628_
timestamp 0
transform -1 0 1370 0 -1 11770
box -6 -8 86 248
use OAI21X1  _4629_
timestamp 0
transform 1 0 1090 0 -1 11770
box -6 -8 106 248
use NAND2X1  _4630_
timestamp 0
transform 1 0 1050 0 1 11770
box -6 -8 86 248
use AND2X2  _4631_
timestamp 0
transform 1 0 1630 0 -1 10810
box -6 -8 106 248
use OAI21X1  _4632_
timestamp 0
transform -1 0 850 0 -1 10330
box -6 -8 106 248
use NAND2X1  _4633_
timestamp 0
transform -1 0 670 0 -1 10330
box -6 -8 86 248
use MUX2X1  _4634_
timestamp 0
transform -1 0 7730 0 1 4090
box -6 -8 126 248
use OAI21X1  _4635_
timestamp 0
transform -1 0 1650 0 -1 9850
box -6 -8 106 248
use NAND2X1  _4636_
timestamp 0
transform 1 0 1370 0 -1 9850
box -6 -8 86 248
use INVX1  _4637_
timestamp 0
transform -1 0 1810 0 -1 9850
box -6 -8 66 248
use AND2X2  _4638_
timestamp 0
transform -1 0 1010 0 -1 11290
box -6 -8 106 248
use OAI21X1  _4639_
timestamp 0
transform 1 0 1130 0 -1 10330
box -6 -8 106 248
use AOI21X1  _4640_
timestamp 0
transform 1 0 990 0 1 10330
box -6 -8 106 248
use INVX1  _4641_
timestamp 0
transform -1 0 1190 0 1 9850
box -6 -8 66 248
use OAI21X1  _4642_
timestamp 0
transform -1 0 3050 0 1 3130
box -6 -8 106 248
use NAND2X1  _4643_
timestamp 0
transform 1 0 3110 0 -1 3130
box -6 -8 86 248
use INVX1  _4644_
timestamp 0
transform -1 0 3590 0 1 3130
box -6 -8 66 248
use OAI21X1  _4645_
timestamp 0
transform -1 0 990 0 1 10810
box -6 -8 106 248
use AOI21X1  _4646_
timestamp 0
transform 1 0 690 0 1 10810
box -6 -8 106 248
use OAI21X1  _4647_
timestamp 0
transform -1 0 1390 0 1 9850
box -6 -8 106 248
use INVX1  _4648_
timestamp 0
transform -1 0 1290 0 1 11770
box -6 -8 66 248
use INVX1  _4649_
timestamp 0
transform -1 0 650 0 1 9850
box -6 -8 66 248
use INVX1  _4650_
timestamp 0
transform -1 0 890 0 -1 10810
box -6 -8 66 248
use OAI21X1  _4651_
timestamp 0
transform 1 0 4150 0 -1 3610
box -6 -8 106 248
use NAND2X1  _4652_
timestamp 0
transform 1 0 3850 0 1 3130
box -6 -8 86 248
use INVX1  _4653_
timestamp 0
transform -1 0 4410 0 -1 3610
box -6 -8 66 248
use NOR2X1  _4654_
timestamp 0
transform -1 0 6990 0 1 10330
box -6 -8 86 248
use INVX1  _4655_
timestamp 0
transform 1 0 2590 0 1 9370
box -6 -8 66 248
use OAI21X1  _4656_
timestamp 0
transform -1 0 2490 0 -1 6490
box -6 -8 106 248
use NAND2X1  _4657_
timestamp 0
transform -1 0 2390 0 1 6010
box -6 -8 86 248
use OAI21X1  _4658_
timestamp 0
transform 1 0 3770 0 1 6010
box -6 -8 106 248
use INVX1  _4659_
timestamp 0
transform -1 0 4030 0 1 6010
box -6 -8 66 248
use NAND3X1  _4660_
timestamp 0
transform -1 0 4450 0 -1 6490
box -6 -8 106 248
use AOI22X1  _4661_
timestamp 0
transform 1 0 4550 0 -1 6490
box -6 -8 126 248
use INVX1  _4662_
timestamp 0
transform 1 0 4010 0 -1 6490
box -6 -8 66 248
use NOR2X1  _4663_
timestamp 0
transform 1 0 3450 0 -1 6490
box -6 -8 86 248
use INVX1  _4664_
timestamp 0
transform 1 0 2590 0 -1 6490
box -6 -8 66 248
use OAI21X1  _4665_
timestamp 0
transform -1 0 7950 0 1 6970
box -6 -8 106 248
use INVX1  _4666_
timestamp 0
transform 1 0 7770 0 1 3610
box -6 -8 66 248
use OAI21X1  _4667_
timestamp 0
transform 1 0 6290 0 -1 3610
box -6 -8 106 248
use OR2X2  _4668_
timestamp 0
transform -1 0 6590 0 -1 3610
box -6 -8 106 248
use INVX1  _4669_
timestamp 0
transform 1 0 490 0 -1 6010
box -6 -8 66 248
use OAI21X1  _4670_
timestamp 0
transform 1 0 4070 0 1 4570
box -6 -8 106 248
use NAND2X1  _4671_
timestamp 0
transform 1 0 3890 0 1 4570
box -6 -8 86 248
use OAI21X1  _4672_
timestamp 0
transform 1 0 2810 0 -1 5530
box -6 -8 106 248
use INVX1  _4673_
timestamp 0
transform -1 0 3070 0 -1 5530
box -6 -8 66 248
use OAI21X1  _4674_
timestamp 0
transform -1 0 3270 0 -1 5530
box -6 -8 106 248
use AND2X2  _4675_
timestamp 0
transform -1 0 3150 0 1 5050
box -6 -8 106 248
use AOI21X1  _4676_
timestamp 0
transform -1 0 3750 0 1 5050
box -6 -8 106 248
use NOR2X1  _4677_
timestamp 0
transform -1 0 3670 0 -1 5050
box -6 -8 86 248
use INVX1  _4678_
timestamp 0
transform 1 0 3430 0 -1 5050
box -6 -8 66 248
use OAI21X1  _4679_
timestamp 0
transform -1 0 3350 0 1 5050
box -6 -8 106 248
use OAI21X1  _4680_
timestamp 0
transform -1 0 2350 0 1 2650
box -6 -8 106 248
use OR2X2  _4681_
timestamp 0
transform 1 0 2050 0 1 2650
box -6 -8 106 248
use INVX8  _4682_
timestamp 0
transform -1 0 7210 0 1 10330
box -6 -8 126 248
use INVX1  _4683_
timestamp 0
transform -1 0 1950 0 -1 7450
box -6 -8 66 248
use OAI21X1  _4684_
timestamp 0
transform 1 0 3810 0 -1 6490
box -6 -8 106 248
use NAND2X1  _4685_
timestamp 0
transform 1 0 3630 0 -1 6490
box -6 -8 86 248
use NOR2X1  _4686_
timestamp 0
transform 1 0 11170 0 1 6970
box -6 -8 86 248
use NAND2X1  _4687_
timestamp 0
transform 1 0 11350 0 1 6970
box -6 -8 86 248
use NAND2X1  _4688_
timestamp 0
transform 1 0 11530 0 1 6970
box -6 -8 86 248
use NOR2X1  _4689_
timestamp 0
transform 1 0 11710 0 1 6970
box -6 -8 86 248
use NAND3X1  _4690_
timestamp 0
transform 1 0 10550 0 -1 7450
box -6 -8 106 248
use NOR2X1  _4691_
timestamp 0
transform 1 0 10190 0 -1 7450
box -6 -8 86 248
use OAI21X1  _4692_
timestamp 0
transform 1 0 10250 0 1 7450
box -6 -8 106 248
use OAI21X1  _4693_
timestamp 0
transform -1 0 9870 0 -1 7930
box -6 -8 106 248
use NAND2X1  _4694_
timestamp 0
transform -1 0 9870 0 1 7930
box -6 -8 86 248
use NOR2X1  _4695_
timestamp 0
transform 1 0 10650 0 1 7450
box -6 -8 86 248
use OAI21X1  _4696_
timestamp 0
transform 1 0 10970 0 -1 8410
box -6 -8 106 248
use NAND3X1  _4697_
timestamp 0
transform 1 0 11450 0 -1 7450
box -6 -8 106 248
use INVX1  _4698_
timestamp 0
transform 1 0 11290 0 -1 7450
box -6 -8 66 248
use NAND3X1  _4699_
timestamp 0
transform 1 0 11290 0 -1 7930
box -6 -8 106 248
use NAND2X1  _4700_
timestamp 0
transform 1 0 11130 0 1 8410
box -6 -8 86 248
use AND2X2  _4701_
timestamp 0
transform -1 0 11590 0 -1 7930
box -6 -8 106 248
use OAI21X1  _4702_
timestamp 0
transform 1 0 11490 0 1 8410
box -6 -8 106 248
use NOR2X1  _4703_
timestamp 0
transform 1 0 11770 0 -1 8890
box -6 -8 86 248
use AND2X2  _4704_
timestamp 0
transform -1 0 11750 0 -1 7450
box -6 -8 106 248
use OAI21X1  _4705_
timestamp 0
transform -1 0 11950 0 -1 7450
box -6 -8 106 248
use OAI21X1  _4706_
timestamp 0
transform -1 0 11890 0 1 7450
box -6 -8 106 248
use AOI21X1  _4707_
timestamp 0
transform 1 0 10750 0 -1 7450
box -6 -8 106 248
use NAND2X1  _4708_
timestamp 0
transform 1 0 10950 0 -1 7450
box -6 -8 86 248
use NOR2X1  _4709_
timestamp 0
transform -1 0 11010 0 1 7930
box -6 -8 86 248
use OAI21X1  _4710_
timestamp 0
transform -1 0 10830 0 1 7930
box -6 -8 106 248
use NOR2X1  _4711_
timestamp 0
transform 1 0 10210 0 1 8410
box -6 -8 86 248
use NAND3X1  _4712_
timestamp 0
transform -1 0 10050 0 -1 8890
box -6 -8 106 248
use NOR2X1  _4713_
timestamp 0
transform 1 0 9790 0 -1 8890
box -6 -8 86 248
use NAND3X1  _4714_
timestamp 0
transform 1 0 9590 0 -1 8890
box -6 -8 106 248
use NAND2X1  _4715_
timestamp 0
transform -1 0 9970 0 -1 8410
box -6 -8 86 248
use NAND2X1  _4716_
timestamp 0
transform 1 0 9330 0 1 8890
box -6 -8 86 248
use OR2X2  _4717_
timestamp 0
transform 1 0 9670 0 1 8410
box -6 -8 106 248
use OAI21X1  _4718_
timestamp 0
transform -1 0 8890 0 1 7930
box -6 -8 106 248
use NAND2X1  _4719_
timestamp 0
transform 1 0 11350 0 1 8890
box -6 -8 86 248
use NAND2X1  _4720_
timestamp 0
transform 1 0 10090 0 1 7450
box -6 -8 86 248
use NOR2X1  _4721_
timestamp 0
transform 1 0 9910 0 1 7450
box -6 -8 86 248
use NAND3X1  _4722_
timestamp 0
transform -1 0 10070 0 -1 7930
box -6 -8 106 248
use NOR2X1  _4723_
timestamp 0
transform -1 0 10050 0 1 7930
box -6 -8 86 248
use INVX2  _4724_
timestamp 0
transform 1 0 4290 0 -1 8410
box -6 -8 66 248
use NOR2X1  _4725_
timestamp 0
transform -1 0 10250 0 -1 7930
box -6 -8 86 248
use NOR2X1  _4726_
timestamp 0
transform -1 0 10450 0 -1 7450
box -6 -8 86 248
use INVX1  _4727_
timestamp 0
transform -1 0 11190 0 -1 7450
box -6 -8 66 248
use NOR2X1  _4728_
timestamp 0
transform 1 0 10230 0 -1 8410
box -6 -8 86 248
use AOI21X1  _4729_
timestamp 0
transform -1 0 10250 0 1 7930
box -6 -8 106 248
use NOR2X1  _4730_
timestamp 0
transform -1 0 10110 0 1 8410
box -6 -8 86 248
use NOR2X1  _4731_
timestamp 0
transform -1 0 11790 0 -1 8410
box -6 -8 86 248
use NAND2X1  _4732_
timestamp 0
transform -1 0 9930 0 1 8410
box -6 -8 86 248
use AOI21X1  _4733_
timestamp 0
transform 1 0 9870 0 1 8890
box -6 -8 106 248
use NOR2X1  _4734_
timestamp 0
transform -1 0 7910 0 -1 10330
box -6 -8 86 248
use OAI21X1  _4735_
timestamp 0
transform 1 0 9390 0 -1 8890
box -6 -8 106 248
use OAI21X1  _4736_
timestamp 0
transform -1 0 10170 0 1 8890
box -6 -8 106 248
use NAND2X1  _4737_
timestamp 0
transform 1 0 9590 0 -1 9370
box -6 -8 86 248
use NOR2X1  _4738_
timestamp 0
transform -1 0 9850 0 -1 9370
box -6 -8 86 248
use NAND3X1  _4739_
timestamp 0
transform -1 0 10050 0 -1 9370
box -6 -8 106 248
use AOI21X1  _4740_
timestamp 0
transform -1 0 10430 0 -1 9370
box -6 -8 106 248
use NOR2X1  _4741_
timestamp 0
transform -1 0 10230 0 -1 9370
box -6 -8 86 248
use NAND2X1  _4742_
timestamp 0
transform 1 0 10390 0 1 8410
box -6 -8 86 248
use OAI21X1  _4743_
timestamp 0
transform 1 0 10150 0 -1 8890
box -6 -8 106 248
use NOR2X1  _4744_
timestamp 0
transform 1 0 10650 0 1 8890
box -6 -8 86 248
use OAI21X1  _4745_
timestamp 0
transform 1 0 10970 0 1 9370
box -6 -8 106 248
use OAI21X1  _4746_
timestamp 0
transform 1 0 10450 0 1 8890
box -6 -8 106 248
use NAND3X1  _4747_
timestamp 0
transform 1 0 8390 0 -1 9370
box -6 -8 106 248
use AND2X2  _4748_
timestamp 0
transform 1 0 8590 0 -1 9370
box -6 -8 106 248
use OAI21X1  _4749_
timestamp 0
transform -1 0 8910 0 -1 8890
box -6 -8 106 248
use NOR2X1  _4750_
timestamp 0
transform 1 0 8590 0 1 9370
box -6 -8 86 248
use INVX2  _4751_
timestamp 0
transform 1 0 3790 0 -1 10330
box -6 -8 66 248
use NAND3X1  _4752_
timestamp 0
transform -1 0 9250 0 1 9370
box -6 -8 106 248
use NOR2X1  _4753_
timestamp 0
transform -1 0 8130 0 -1 9850
box -6 -8 86 248
use INVX1  _4754_
timestamp 0
transform 1 0 8190 0 -1 10330
box -6 -8 66 248
use INVX1  _4755_
timestamp 0
transform 1 0 7310 0 -1 9850
box -6 -8 66 248
use NOR2X1  _4756_
timestamp 0
transform 1 0 6970 0 -1 9850
box -6 -8 86 248
use NAND2X1  _4757_
timestamp 0
transform 1 0 8410 0 -1 9850
box -6 -8 86 248
use NAND3X1  _4758_
timestamp 0
transform -1 0 10550 0 1 7450
box -6 -8 106 248
use NOR2X1  _4759_
timestamp 0
transform 1 0 10830 0 1 7450
box -6 -8 86 248
use NAND3X1  _4760_
timestamp 0
transform -1 0 11190 0 -1 7930
box -6 -8 106 248
use AND2X2  _4761_
timestamp 0
transform 1 0 11390 0 1 7450
box -6 -8 106 248
use NAND2X1  _4762_
timestamp 0
transform -1 0 10610 0 1 11770
box -6 -8 86 248
use NOR2X1  _4763_
timestamp 0
transform 1 0 11890 0 -1 8410
box -6 -8 86 248
use INVX1  _4764_
timestamp 0
transform 1 0 10930 0 -1 7930
box -6 -8 66 248
use NAND2X1  _4765_
timestamp 0
transform -1 0 11250 0 -1 8410
box -6 -8 86 248
use OAI21X1  _4766_
timestamp 0
transform -1 0 10630 0 1 7930
box -6 -8 106 248
use NOR2X1  _4767_
timestamp 0
transform -1 0 10630 0 -1 7930
box -6 -8 86 248
use OAI21X1  _4768_
timestamp 0
transform 1 0 10350 0 -1 7930
box -6 -8 106 248
use OAI21X1  _4769_
timestamp 0
transform 1 0 10730 0 -1 7930
box -6 -8 106 248
use NAND2X1  _4770_
timestamp 0
transform 1 0 11210 0 -1 10330
box -6 -8 86 248
use NAND2X1  _4771_
timestamp 0
transform 1 0 12070 0 -1 7930
box -6 -8 86 248
use AOI21X1  _4772_
timestamp 0
transform 1 0 9390 0 -1 7930
box -6 -8 106 248
use OAI21X1  _4773_
timestamp 0
transform -1 0 8950 0 -1 7930
box -6 -8 106 248
use OAI21X1  _4774_
timestamp 0
transform 1 0 2610 0 1 6490
box -6 -8 106 248
use INVX1  _4775_
timestamp 0
transform 1 0 2770 0 -1 6970
box -6 -8 66 248
use OAI21X1  _4776_
timestamp 0
transform 1 0 2930 0 -1 6970
box -6 -8 106 248
use AND2X2  _4777_
timestamp 0
transform -1 0 3230 0 -1 6970
box -6 -8 106 248
use AOI21X1  _4778_
timestamp 0
transform -1 0 3830 0 -1 6970
box -6 -8 106 248
use NOR2X1  _4779_
timestamp 0
transform 1 0 3930 0 -1 6970
box -6 -8 86 248
use NAND3X1  _4780_
timestamp 0
transform -1 0 8890 0 -1 9370
box -6 -8 106 248
use INVX1  _4781_
timestamp 0
transform 1 0 3650 0 1 6490
box -6 -8 66 248
use OAI21X1  _4782_
timestamp 0
transform 1 0 3330 0 -1 6970
box -6 -8 106 248
use INVX4  _4783_
timestamp 0
transform 1 0 9150 0 1 7450
box -6 -8 86 248
use NOR2X1  _4784_
timestamp 0
transform 1 0 7790 0 1 7450
box -6 -8 86 248
use INVX1  _4785_
timestamp 0
transform 1 0 2150 0 -1 8890
box -6 -8 66 248
use OAI21X1  _4786_
timestamp 0
transform -1 0 4110 0 1 3610
box -6 -8 106 248
use NAND2X1  _4787_
timestamp 0
transform -1 0 3770 0 1 3130
box -6 -8 86 248
use INVX1  _4788_
timestamp 0
transform -1 0 4270 0 1 3610
box -6 -8 66 248
use NAND2X1  _4789_
timestamp 0
transform 1 0 7270 0 1 6490
box -6 -8 86 248
use NOR2X1  _4790_
timestamp 0
transform 1 0 7330 0 -1 6490
box -6 -8 86 248
use NAND3X1  _4791_
timestamp 0
transform -1 0 7950 0 1 6490
box -6 -8 106 248
use NOR2X1  _4792_
timestamp 0
transform -1 0 7970 0 -1 7450
box -6 -8 86 248
use OAI21X1  _4793_
timestamp 0
transform -1 0 7950 0 -1 7930
box -6 -8 106 248
use NOR2X1  _4794_
timestamp 0
transform -1 0 7570 0 -1 7930
box -6 -8 86 248
use NOR2X1  _4795_
timestamp 0
transform -1 0 7630 0 -1 8890
box -6 -8 86 248
use NAND2X1  _4796_
timestamp 0
transform 1 0 11870 0 1 9850
box -6 -8 86 248
use NOR2X1  _4797_
timestamp 0
transform 1 0 8610 0 1 7930
box -6 -8 86 248
use INVX1  _4798_
timestamp 0
transform 1 0 10070 0 -1 8410
box -6 -8 66 248
use NAND2X1  _4799_
timestamp 0
transform -1 0 9970 0 1 9370
box -6 -8 86 248
use NAND3X1  _4800_
timestamp 0
transform 1 0 8550 0 1 7450
box -6 -8 106 248
use NAND2X1  _4801_
timestamp 0
transform 1 0 11010 0 1 7450
box -6 -8 86 248
use NAND2X1  _4802_
timestamp 0
transform -1 0 10610 0 -1 8890
box -6 -8 86 248
use NAND2X1  _4803_
timestamp 0
transform -1 0 7510 0 -1 8410
box -6 -8 86 248
use INVX2  _4804_
timestamp 0
transform -1 0 7170 0 1 6490
box -6 -8 66 248
use OAI21X1  _4805_
timestamp 0
transform -1 0 7090 0 1 7450
box -6 -8 106 248
use OAI21X1  _4806_
timestamp 0
transform -1 0 9450 0 -1 8410
box -6 -8 106 248
use NAND2X1  _4807_
timestamp 0
transform -1 0 9210 0 1 9850
box -6 -8 86 248
use NOR2X1  _4808_
timestamp 0
transform -1 0 8830 0 -1 7450
box -6 -8 86 248
use NAND3X1  _4809_
timestamp 0
transform -1 0 8850 0 1 7450
box -6 -8 106 248
use NAND2X1  _4810_
timestamp 0
transform -1 0 9070 0 -1 8410
box -6 -8 86 248
use NAND2X1  _4811_
timestamp 0
transform 1 0 11990 0 1 7450
box -6 -8 86 248
use NOR2X1  _4812_
timestamp 0
transform 1 0 12050 0 -1 8410
box -6 -8 86 248
use NAND2X1  _4813_
timestamp 0
transform 1 0 11530 0 1 8890
box -6 -8 86 248
use NOR2X1  _4814_
timestamp 0
transform 1 0 11410 0 1 11770
box -6 -8 86 248
use OAI21X1  _4815_
timestamp 0
transform -1 0 9190 0 -1 7450
box -6 -8 106 248
use NAND2X1  _4816_
timestamp 0
transform -1 0 9610 0 1 7450
box -6 -8 86 248
use NOR2X1  _4817_
timestamp 0
transform -1 0 11670 0 -1 8890
box -6 -8 86 248
use NAND2X1  _4818_
timestamp 0
transform -1 0 11610 0 1 9850
box -6 -8 86 248
use INVX2  _4819_
timestamp 0
transform -1 0 6530 0 1 5530
box -6 -8 66 248
use NOR2X1  _4820_
timestamp 0
transform 1 0 8050 0 1 6970
box -6 -8 86 248
use NAND3X1  _4821_
timestamp 0
transform 1 0 11690 0 -1 7930
box -6 -8 106 248
use NAND2X1  _4822_
timestamp 0
transform 1 0 11890 0 -1 7930
box -6 -8 86 248
use NOR3X1  _4823_
timestamp 0
transform 1 0 11670 0 -1 9370
box -6 -8 186 248
use NOR2X1  _4824_
timestamp 0
transform -1 0 11590 0 1 7930
box -6 -8 86 248
use NOR2X1  _4825_
timestamp 0
transform 1 0 11230 0 -1 8890
box -6 -8 86 248
use NOR2X1  _4826_
timestamp 0
transform -1 0 11130 0 -1 8890
box -6 -8 86 248
use NAND2X1  _4827_
timestamp 0
transform -1 0 11830 0 -1 10330
box -6 -8 86 248
use NOR2X1  _4828_
timestamp 0
transform -1 0 11910 0 1 10330
box -6 -8 86 248
use NAND2X1  _4829_
timestamp 0
transform 1 0 11690 0 1 7930
box -6 -8 86 248
use OAI21X1  _4830_
timestamp 0
transform 1 0 9050 0 -1 7930
box -6 -8 106 248
use OAI21X1  _4831_
timestamp 0
transform -1 0 9490 0 1 7930
box -6 -8 106 248
use NOR2X1  _4832_
timestamp 0
transform 1 0 11930 0 -1 8890
box -6 -8 86 248
use AND2X2  _4833_
timestamp 0
transform 1 0 8430 0 -1 6970
box -6 -8 106 248
use NOR2X1  _4834_
timestamp 0
transform 1 0 8230 0 -1 8410
box -6 -8 86 248
use NAND3X1  _4835_
timestamp 0
transform -1 0 8510 0 -1 8410
box -6 -8 106 248
use NAND2X1  _4836_
timestamp 0
transform 1 0 9710 0 -1 8410
box -6 -8 86 248
use NOR2X1  _4837_
timestamp 0
transform -1 0 10910 0 1 8890
box -6 -8 86 248
use NOR2X1  _4838_
timestamp 0
transform 1 0 11870 0 1 8410
box -6 -8 86 248
use NAND2X1  _4839_
timestamp 0
transform 1 0 12130 0 -1 9370
box -6 -8 86 248
use NAND2X1  _4840_
timestamp 0
transform 1 0 9310 0 1 8410
box -6 -8 86 248
use NAND2X1  _4841_
timestamp 0
transform 1 0 10350 0 1 7930
box -6 -8 86 248
use NOR2X1  _4842_
timestamp 0
transform 1 0 12050 0 1 8410
box -6 -8 86 248
use NOR2X1  _4843_
timestamp 0
transform 1 0 11210 0 -1 9850
box -6 -8 86 248
use INVX1  _4844_
timestamp 0
transform -1 0 11230 0 1 9370
box -6 -8 66 248
use NOR2X1  _4845_
timestamp 0
transform -1 0 12030 0 -1 9370
box -6 -8 86 248
use NAND2X1  _4846_
timestamp 0
transform 1 0 11950 0 1 11770
box -6 -8 86 248
use NOR3X1  _4847_
timestamp 0
transform -1 0 8590 0 -1 7930
box -6 -8 186 248
use NAND2X1  _4848_
timestamp 0
transform -1 0 8510 0 1 7930
box -6 -8 86 248
use OAI21X1  _4849_
timestamp 0
transform 1 0 9110 0 1 8410
box -6 -8 106 248
use AND2X2  _4850_
timestamp 0
transform 1 0 9350 0 1 9370
box -6 -8 106 248
use AND2X2  _4851_
timestamp 0
transform 1 0 11330 0 1 9850
box -6 -8 106 248
use NOR2X1  _4852_
timestamp 0
transform 1 0 11690 0 1 9850
box -6 -8 86 248
use NOR2X1  _4853_
timestamp 0
transform 1 0 12110 0 -1 8890
box -6 -8 86 248
use NAND2X1  _4854_
timestamp 0
transform -1 0 11310 0 1 11770
box -6 -8 86 248
use NOR2X1  _4855_
timestamp 0
transform -1 0 8330 0 1 7930
box -6 -8 86 248
use NOR2X1  _4856_
timestamp 0
transform -1 0 8350 0 -1 8890
box -6 -8 86 248
use INVX4  _4857_
timestamp 0
transform -1 0 10430 0 -1 8890
box -6 -8 86 248
use NAND2X1  _4858_
timestamp 0
transform -1 0 10570 0 -1 9850
box -6 -8 86 248
use NOR2X1  _4859_
timestamp 0
transform -1 0 7310 0 1 8410
box -6 -8 86 248
use NAND2X1  _4860_
timestamp 0
transform -1 0 10490 0 1 9370
box -6 -8 86 248
use INVX1  _4861_
timestamp 0
transform -1 0 10730 0 -1 9850
box -6 -8 66 248
use NOR2X1  _4862_
timestamp 0
transform 1 0 11490 0 -1 9370
box -6 -8 86 248
use INVX8  _4863_
timestamp 0
transform -1 0 10850 0 1 8410
box -6 -8 126 248
use INVX1  _4864_
timestamp 0
transform -1 0 10630 0 1 8410
box -6 -8 66 248
use NAND2X1  _4865_
timestamp 0
transform 1 0 10610 0 -1 8410
box -6 -8 86 248
use NOR2X1  _4866_
timestamp 0
transform 1 0 11690 0 1 8410
box -6 -8 86 248
use NAND2X1  _4867_
timestamp 0
transform 1 0 11870 0 1 9370
box -6 -8 86 248
use NOR2X1  _4868_
timestamp 0
transform -1 0 11430 0 -1 8410
box -6 -8 86 248
use INVX2  _4869_
timestamp 0
transform -1 0 10950 0 -1 8890
box -6 -8 66 248
use NAND3X1  _4870_
timestamp 0
transform 1 0 8150 0 1 8410
box -6 -8 106 248
use INVX1  _4871_
timestamp 0
transform 1 0 7990 0 1 8410
box -6 -8 66 248
use NOR2X1  _4872_
timestamp 0
transform 1 0 7870 0 1 7930
box -6 -8 86 248
use NAND2X1  _4873_
timestamp 0
transform -1 0 11470 0 -1 10330
box -6 -8 86 248
use NOR2X1  _4874_
timestamp 0
transform 1 0 11930 0 -1 10330
box -6 -8 86 248
use INVX8  _4875_
timestamp 0
transform -1 0 7730 0 -1 8410
box -6 -8 126 248
use NAND3X1  _4876_
timestamp 0
transform -1 0 10630 0 -1 9370
box -6 -8 106 248
use NOR2X1  _4877_
timestamp 0
transform 1 0 10950 0 1 8410
box -6 -8 86 248
use NOR2X1  _4878_
timestamp 0
transform 1 0 11390 0 -1 9850
box -6 -8 86 248
use NOR2X1  _4879_
timestamp 0
transform 1 0 12050 0 1 9850
box -6 -8 86 248
use INVX1  _4880_
timestamp 0
transform -1 0 12150 0 -1 9850
box -6 -8 66 248
use OAI21X1  _4881_
timestamp 0
transform -1 0 9230 0 1 8890
box -6 -8 106 248
use NOR2X1  _4882_
timestamp 0
transform 1 0 12070 0 1 8890
box -6 -8 86 248
use NAND2X1  _4883_
timestamp 0
transform 1 0 11890 0 1 8890
box -6 -8 86 248
use INVX1  _4884_
timestamp 0
transform 1 0 11710 0 1 9370
box -6 -8 66 248
use NAND2X1  _4885_
timestamp 0
transform -1 0 11810 0 -1 9850
box -6 -8 86 248
use NOR2X1  _4886_
timestamp 0
transform 1 0 11010 0 1 8890
box -6 -8 86 248
use INVX1  _4887_
timestamp 0
transform 1 0 11050 0 -1 10330
box -6 -8 66 248
use NOR2X1  _4888_
timestamp 0
transform 1 0 11710 0 1 8890
box -6 -8 86 248
use NAND2X1  _4889_
timestamp 0
transform 1 0 12050 0 1 9370
box -6 -8 86 248
use INVX1  _4890_
timestamp 0
transform 1 0 11570 0 -1 9850
box -6 -8 66 248
use NAND2X1  _4891_
timestamp 0
transform 1 0 11910 0 -1 9850
box -6 -8 86 248
use INVX1  _4892_
timestamp 0
transform -1 0 12150 0 -1 10330
box -6 -8 66 248
use INVX1  _4893_
timestamp 0
transform -1 0 2590 0 -1 7450
box -6 -8 66 248
use INVX4  _4894_
timestamp 0
transform 1 0 9750 0 1 4090
box -6 -8 86 248
use NAND2X1  _4895_
timestamp 0
transform 1 0 8490 0 1 4570
box -6 -8 86 248
use INVX2  _4896_
timestamp 0
transform -1 0 9570 0 -1 6970
box -6 -8 66 248
use NAND2X1  _4897_
timestamp 0
transform 1 0 9570 0 1 6010
box -6 -8 86 248
use INVX2  _4898_
timestamp 0
transform 1 0 9750 0 1 6010
box -6 -8 66 248
use NAND2X1  _4899_
timestamp 0
transform -1 0 9290 0 1 6490
box -6 -8 86 248
use NAND2X1  _4900_
timestamp 0
transform -1 0 9630 0 1 6490
box -6 -8 86 248
use AOI22X1  _4901_
timestamp 0
transform -1 0 10050 0 1 6490
box -6 -8 126 248
use INVX2  _4902_
timestamp 0
transform 1 0 10270 0 -1 6490
box -6 -8 66 248
use INVX1  _4903_
timestamp 0
transform 1 0 9730 0 -1 6490
box -6 -8 66 248
use INVX1  _4904_
timestamp 0
transform -1 0 10490 0 -1 6970
box -6 -8 66 248
use OAI21X1  _4905_
timestamp 0
transform 1 0 9730 0 1 6490
box -6 -8 106 248
use NAND2X1  _4906_
timestamp 0
transform -1 0 9970 0 -1 6490
box -6 -8 86 248
use NAND2X1  _4907_
timestamp 0
transform -1 0 9630 0 -1 6490
box -6 -8 86 248
use OAI21X1  _4908_
timestamp 0
transform 1 0 10070 0 -1 6490
box -6 -8 106 248
use INVX2  _4909_
timestamp 0
transform 1 0 11010 0 1 6970
box -6 -8 66 248
use NOR2X1  _4910_
timestamp 0
transform -1 0 11450 0 -1 6490
box -6 -8 86 248
use OAI21X1  _4911_
timestamp 0
transform 1 0 11330 0 -1 6970
box -6 -8 106 248
use AOI21X1  _4912_
timestamp 0
transform 1 0 11130 0 1 6490
box -6 -8 106 248
use OAI21X1  _4913_
timestamp 0
transform -1 0 11050 0 1 6490
box -6 -8 106 248
use INVX1  _4914_
timestamp 0
transform 1 0 11530 0 -1 6970
box -6 -8 66 248
use OAI21X1  _4915_
timestamp 0
transform -1 0 10910 0 1 6970
box -6 -8 106 248
use NOR2X1  _4916_
timestamp 0
transform 1 0 10590 0 -1 6970
box -6 -8 86 248
use INVX1  _4917_
timestamp 0
transform -1 0 10690 0 -1 6490
box -6 -8 66 248
use NOR2X1  _4918_
timestamp 0
transform -1 0 11070 0 -1 6490
box -6 -8 86 248
use OAI21X1  _4919_
timestamp 0
transform 1 0 11170 0 -1 6490
box -6 -8 106 248
use INVX1  _4920_
timestamp 0
transform 1 0 8590 0 -1 6490
box -6 -8 66 248
use NAND3X1  _4921_
timestamp 0
transform -1 0 8890 0 1 6490
box -6 -8 106 248
use AOI22X1  _4922_
timestamp 0
transform -1 0 9110 0 1 6490
box -6 -8 126 248
use INVX1  _4923_
timestamp 0
transform 1 0 9390 0 1 6490
box -6 -8 66 248
use NOR2X1  _4924_
timestamp 0
transform 1 0 9370 0 -1 6490
box -6 -8 86 248
use OAI21X1  _4925_
timestamp 0
transform -1 0 9270 0 -1 6490
box -6 -8 106 248
use OAI22X1  _4926_
timestamp 0
transform 1 0 8950 0 -1 6490
box -6 -8 126 248
use OAI21X1  _4927_
timestamp 0
transform -1 0 11430 0 1 6490
box -6 -8 106 248
use AOI21X1  _4928_
timestamp 0
transform 1 0 11530 0 1 6490
box -6 -8 106 248
use INVX1  _4929_
timestamp 0
transform 1 0 12110 0 -1 6970
box -6 -8 66 248
use OAI21X1  _4930_
timestamp 0
transform 1 0 11690 0 -1 6970
box -6 -8 106 248
use MUX2X1  _4931_
timestamp 0
transform -1 0 12010 0 -1 6970
box -6 -8 126 248
use NAND2X1  _4932_
timestamp 0
transform -1 0 11790 0 -1 6490
box -6 -8 86 248
use INVX1  _4933_
timestamp 0
transform -1 0 11230 0 -1 6970
box -6 -8 66 248
use OAI21X1  _4934_
timestamp 0
transform 1 0 10970 0 -1 6970
box -6 -8 106 248
use OAI21X1  _4935_
timestamp 0
transform -1 0 10870 0 -1 6970
box -6 -8 106 248
use MUX2X1  _4936_
timestamp 0
transform -1 0 9790 0 -1 6970
box -6 -8 126 248
use NAND2X1  _4937_
timestamp 0
transform -1 0 9970 0 -1 6970
box -6 -8 86 248
use NAND2X1  _4938_
timestamp 0
transform 1 0 10070 0 -1 6970
box -6 -8 86 248
use AOI21X1  _4939_
timestamp 0
transform 1 0 10150 0 1 6490
box -6 -8 106 248
use NAND2X1  _4940_
timestamp 0
transform 1 0 10250 0 -1 6970
box -6 -8 86 248
use NAND3X1  _4941_
timestamp 0
transform 1 0 10350 0 1 6490
box -6 -8 106 248
use AOI22X1  _4942_
timestamp 0
transform -1 0 10850 0 1 6490
box -6 -8 126 248
use OAI21X1  _4943_
timestamp 0
transform 1 0 11730 0 1 6490
box -6 -8 106 248
use OAI21X1  _4944_
timestamp 0
transform -1 0 12030 0 1 6490
box -6 -8 106 248
use NAND2X1  _4945_
timestamp 0
transform 1 0 11890 0 -1 6490
box -6 -8 86 248
use NAND2X1  _4946_
timestamp 0
transform -1 0 11930 0 1 6010
box -6 -8 86 248
use OAI21X1  _4947_
timestamp 0
transform -1 0 8770 0 1 4570
box -6 -8 106 248
use NAND2X1  _4948_
timestamp 0
transform 1 0 9010 0 1 4090
box -6 -8 86 248
use NOR2X1  _4949_
timestamp 0
transform 1 0 12130 0 1 6490
box -6 -8 86 248
use OAI21X1  _4950_
timestamp 0
transform -1 0 12170 0 -1 6490
box -6 -8 106 248
use NAND2X1  _4951_
timestamp 0
transform -1 0 8690 0 -1 5530
box -6 -8 86 248
use NAND3X1  _4952_
timestamp 0
transform 1 0 8990 0 1 6010
box -6 -8 106 248
use AOI22X1  _4953_
timestamp 0
transform -1 0 9010 0 -1 6010
box -6 -8 126 248
use INVX1  _4954_
timestamp 0
transform -1 0 9250 0 1 6010
box -6 -8 66 248
use OAI21X1  _4955_
timestamp 0
transform -1 0 8850 0 -1 6490
box -6 -8 106 248
use NAND2X1  _4956_
timestamp 0
transform -1 0 8910 0 1 6010
box -6 -8 86 248
use OAI21X1  _4957_
timestamp 0
transform -1 0 8790 0 -1 6010
box -6 -8 106 248
use OAI21X1  _4958_
timestamp 0
transform -1 0 11170 0 -1 6010
box -6 -8 106 248
use AOI21X1  _4959_
timestamp 0
transform 1 0 11270 0 -1 6010
box -6 -8 106 248
use OAI21X1  _4960_
timestamp 0
transform -1 0 11570 0 -1 6010
box -6 -8 106 248
use OAI21X1  _4961_
timestamp 0
transform 1 0 11670 0 -1 6010
box -6 -8 106 248
use INVX1  _4962_
timestamp 0
transform 1 0 12070 0 -1 6010
box -6 -8 66 248
use NAND2X1  _4963_
timestamp 0
transform 1 0 12030 0 1 5530
box -6 -8 86 248
use NAND3X1  _4964_
timestamp 0
transform 1 0 12030 0 1 6010
box -6 -8 106 248
use NAND2X1  _4965_
timestamp 0
transform -1 0 11930 0 1 5530
box -6 -8 86 248
use OAI21X1  _4966_
timestamp 0
transform -1 0 9290 0 1 4090
box -6 -8 106 248
use NAND2X1  _4967_
timestamp 0
transform 1 0 8130 0 1 4570
box -6 -8 86 248
use INVX1  _4968_
timestamp 0
transform 1 0 11710 0 -1 5530
box -6 -8 66 248
use AND2X2  _4969_
timestamp 0
transform 1 0 12070 0 -1 5530
box -6 -8 106 248
use NAND2X1  _4970_
timestamp 0
transform 1 0 9110 0 -1 6010
box -6 -8 86 248
use AND2X2  _4971_
timestamp 0
transform -1 0 8410 0 1 5530
box -6 -8 106 248
use NAND2X1  _4972_
timestamp 0
transform -1 0 8770 0 1 5530
box -6 -8 86 248
use AOI22X1  _4973_
timestamp 0
transform -1 0 8990 0 1 5530
box -6 -8 126 248
use OAI21X1  _4974_
timestamp 0
transform 1 0 8790 0 -1 5530
box -6 -8 106 248
use OAI21X1  _4975_
timestamp 0
transform 1 0 8990 0 -1 5530
box -6 -8 106 248
use OAI21X1  _4976_
timestamp 0
transform 1 0 11650 0 1 6010
box -6 -8 106 248
use AOI21X1  _4977_
timestamp 0
transform 1 0 11450 0 1 6010
box -6 -8 106 248
use OAI21X1  _4978_
timestamp 0
transform 1 0 11470 0 1 5050
box -6 -8 106 248
use OAI21X1  _4979_
timestamp 0
transform 1 0 11490 0 -1 5050
box -6 -8 106 248
use INVX1  _4980_
timestamp 0
transform 1 0 11870 0 -1 5050
box -6 -8 66 248
use OAI21X1  _4981_
timestamp 0
transform -1 0 11950 0 1 5050
box -6 -8 106 248
use AOI21X1  _4982_
timestamp 0
transform -1 0 11970 0 -1 5530
box -6 -8 106 248
use NAND2X1  _4983_
timestamp 0
transform 1 0 11670 0 1 5050
box -6 -8 86 248
use NAND2X1  _4984_
timestamp 0
transform 1 0 11290 0 1 5050
box -6 -8 86 248
use OAI21X1  _4985_
timestamp 0
transform -1 0 8190 0 -1 5050
box -6 -8 106 248
use NAND2X1  _4986_
timestamp 0
transform 1 0 9150 0 -1 5050
box -6 -8 86 248
use NAND2X1  _4987_
timestamp 0
transform 1 0 11670 0 1 5530
box -6 -8 86 248
use NAND3X1  _4988_
timestamp 0
transform -1 0 11970 0 -1 6010
box -6 -8 106 248
use NAND3X1  _4989_
timestamp 0
transform -1 0 11570 0 1 5530
box -6 -8 106 248
use NAND2X1  _4990_
timestamp 0
transform -1 0 11370 0 1 5530
box -6 -8 86 248
use NAND2X1  _4991_
timestamp 0
transform 1 0 11690 0 -1 5050
box -6 -8 86 248
use OAI21X1  _4992_
timestamp 0
transform -1 0 11610 0 -1 5530
box -6 -8 106 248
use OAI21X1  _4993_
timestamp 0
transform 1 0 11330 0 -1 5530
box -6 -8 106 248
use NAND2X1  _4994_
timestamp 0
transform 1 0 9350 0 1 5050
box -6 -8 86 248
use AND2X2  _4995_
timestamp 0
transform -1 0 10010 0 1 6010
box -6 -8 106 248
use NAND2X1  _4996_
timestamp 0
transform 1 0 9290 0 -1 6010
box -6 -8 86 248
use AOI22X1  _4997_
timestamp 0
transform -1 0 9470 0 1 6010
box -6 -8 126 248
use OAI21X1  _4998_
timestamp 0
transform 1 0 9470 0 -1 6010
box -6 -8 106 248
use OAI21X1  _4999_
timestamp 0
transform -1 0 9410 0 1 5530
box -6 -8 106 248
use OAI21X1  _5000_
timestamp 0
transform 1 0 11070 0 1 6010
box -6 -8 106 248
use AOI21X1  _5001_
timestamp 0
transform -1 0 10970 0 1 6010
box -6 -8 106 248
use OAI21X1  _5002_
timestamp 0
transform -1 0 10790 0 1 5530
box -6 -8 106 248
use OAI21X1  _5003_
timestamp 0
transform -1 0 10850 0 -1 5530
box -6 -8 106 248
use INVX1  _5004_
timestamp 0
transform 1 0 10950 0 -1 5530
box -6 -8 66 248
use NOR2X1  _5005_
timestamp 0
transform -1 0 10990 0 1 5050
box -6 -8 86 248
use OR2X2  _5006_
timestamp 0
transform 1 0 11450 0 1 4570
box -6 -8 106 248
use OAI21X1  _5007_
timestamp 0
transform 1 0 12050 0 1 5050
box -6 -8 106 248
use NAND2X1  _5008_
timestamp 0
transform 1 0 12030 0 -1 5050
box -6 -8 86 248
use NAND2X1  _5009_
timestamp 0
transform 1 0 12050 0 1 4570
box -6 -8 86 248
use INVX1  _5010_
timestamp 0
transform -1 0 11390 0 -1 5050
box -6 -8 66 248
use AOI21X1  _5011_
timestamp 0
transform 1 0 11850 0 1 4570
box -6 -8 106 248
use AOI22X1  _5012_
timestamp 0
transform 1 0 11630 0 1 4570
box -6 -8 126 248
use OAI21X1  _5013_
timestamp 0
transform -1 0 10410 0 1 5050
box -6 -8 106 248
use OAI21X1  _5014_
timestamp 0
transform -1 0 9630 0 1 5050
box -6 -8 106 248
use NAND2X1  _5015_
timestamp 0
transform 1 0 8310 0 1 4570
box -6 -8 86 248
use OAI21X1  _5016_
timestamp 0
transform 1 0 10710 0 1 5050
box -6 -8 106 248
use NAND2X1  _5017_
timestamp 0
transform 1 0 8970 0 1 5050
box -6 -8 86 248
use AND2X2  _5018_
timestamp 0
transform 1 0 8510 0 1 5530
box -6 -8 106 248
use NAND2X1  _5019_
timestamp 0
transform 1 0 9190 0 -1 5530
box -6 -8 86 248
use AOI22X1  _5020_
timestamp 0
transform 1 0 9090 0 1 5530
box -6 -8 126 248
use OAI21X1  _5021_
timestamp 0
transform 1 0 9370 0 -1 5530
box -6 -8 106 248
use OAI21X1  _5022_
timestamp 0
transform -1 0 9250 0 1 5050
box -6 -8 106 248
use OAI21X1  _5023_
timestamp 0
transform -1 0 10970 0 -1 6010
box -6 -8 106 248
use AOI21X1  _5024_
timestamp 0
transform 1 0 10890 0 1 5530
box -6 -8 106 248
use OAI21X1  _5025_
timestamp 0
transform -1 0 11190 0 1 5050
box -6 -8 106 248
use OAI21X1  _5026_
timestamp 0
transform 1 0 11130 0 -1 5050
box -6 -8 106 248
use INVX1  _5027_
timestamp 0
transform -1 0 10970 0 1 4570
box -6 -8 66 248
use NAND2X1  _5028_
timestamp 0
transform -1 0 10810 0 1 4570
box -6 -8 86 248
use OR2X2  _5029_
timestamp 0
transform 1 0 11090 0 1 5530
box -6 -8 106 248
use AOI22X1  _5030_
timestamp 0
transform 1 0 11110 0 -1 5530
box -6 -8 126 248
use NAND2X1  _5031_
timestamp 0
transform 1 0 11870 0 -1 4570
box -6 -8 86 248
use NAND2X1  _5032_
timestamp 0
transform 1 0 11690 0 -1 4570
box -6 -8 86 248
use OAI21X1  _5033_
timestamp 0
transform -1 0 9110 0 -1 4570
box -6 -8 106 248
use NAND2X1  _5034_
timestamp 0
transform -1 0 9290 0 -1 4570
box -6 -8 86 248
use OAI21X1  _5035_
timestamp 0
transform 1 0 11250 0 1 4570
box -6 -8 106 248
use NAND2X1  _5036_
timestamp 0
transform 1 0 9930 0 1 5530
box -6 -8 86 248
use AND2X2  _5037_
timestamp 0
transform 1 0 9730 0 1 5530
box -6 -8 106 248
use NAND2X1  _5038_
timestamp 0
transform 1 0 9570 0 -1 5530
box -6 -8 86 248
use AOI22X1  _5039_
timestamp 0
transform 1 0 9510 0 1 5530
box -6 -8 126 248
use OAI21X1  _5040_
timestamp 0
transform 1 0 9750 0 -1 5530
box -6 -8 106 248
use OAI21X1  _5041_
timestamp 0
transform 1 0 9950 0 -1 5530
box -6 -8 106 248
use OAI21X1  _5042_
timestamp 0
transform 1 0 10670 0 -1 6010
box -6 -8 106 248
use AOI21X1  _5043_
timestamp 0
transform 1 0 10490 0 1 5530
box -6 -8 106 248
use OAI21X1  _5044_
timestamp 0
transform 1 0 10550 0 -1 5530
box -6 -8 106 248
use OAI21X1  _5045_
timestamp 0
transform -1 0 10610 0 1 5050
box -6 -8 106 248
use INVX1  _5046_
timestamp 0
transform 1 0 10970 0 -1 4570
box -6 -8 66 248
use NAND2X1  _5047_
timestamp 0
transform 1 0 11070 0 1 4570
box -6 -8 86 248
use NAND3X1  _5048_
timestamp 0
transform 1 0 11510 0 -1 4570
box -6 -8 106 248
use NAND2X1  _5049_
timestamp 0
transform -1 0 11410 0 -1 4570
box -6 -8 86 248
use OAI21X1  _5050_
timestamp 0
transform -1 0 9490 0 -1 4570
box -6 -8 106 248
use INVX1  _5051_
timestamp 0
transform 1 0 8410 0 1 6490
box -6 -8 66 248
use AOI21X1  _5052_
timestamp 0
transform -1 0 10630 0 1 6490
box -6 -8 106 248
use OAI21X1  _5053_
timestamp 0
transform -1 0 10890 0 -1 6490
box -6 -8 106 248
use OAI21X1  _5054_
timestamp 0
transform -1 0 10530 0 -1 6490
box -6 -8 106 248
use OAI22X1  _5055_
timestamp 0
transform 1 0 8570 0 1 6490
box -6 -8 126 248
use INVX1  _5056_
timestamp 0
transform 1 0 8190 0 1 6010
box -6 -8 66 248
use NOR2X1  _5057_
timestamp 0
transform 1 0 8410 0 -1 6490
box -6 -8 86 248
use NAND3X1  _5058_
timestamp 0
transform -1 0 8310 0 -1 6490
box -6 -8 106 248
use NOR2X1  _5059_
timestamp 0
transform 1 0 8050 0 1 6490
box -6 -8 86 248
use NOR2X1  _5060_
timestamp 0
transform -1 0 7750 0 -1 6490
box -6 -8 86 248
use NAND2X1  _5061_
timestamp 0
transform -1 0 7930 0 -1 6490
box -6 -8 86 248
use NOR2X1  _5062_
timestamp 0
transform 1 0 8030 0 -1 6490
box -6 -8 86 248
use INVX1  _5063_
timestamp 0
transform -1 0 8110 0 -1 6010
box -6 -8 66 248
use AND2X2  _5064_
timestamp 0
transform -1 0 7670 0 1 5530
box -6 -8 106 248
use NOR2X1  _5065_
timestamp 0
transform -1 0 7850 0 1 5530
box -6 -8 86 248
use NOR2X1  _5066_
timestamp 0
transform -1 0 7790 0 -1 5530
box -6 -8 86 248
use NOR2X1  _5067_
timestamp 0
transform -1 0 8490 0 1 5050
box -6 -8 86 248
use NAND2X1  _5068_
timestamp 0
transform -1 0 8510 0 -1 5530
box -6 -8 86 248
use INVX1  _5069_
timestamp 0
transform -1 0 8330 0 -1 5530
box -6 -8 66 248
use OAI21X1  _5070_
timestamp 0
transform -1 0 7990 0 -1 5530
box -6 -8 106 248
use NOR2X1  _5071_
timestamp 0
transform 1 0 8090 0 -1 5530
box -6 -8 86 248
use OAI21X1  _5072_
timestamp 0
transform -1 0 7610 0 -1 5530
box -6 -8 106 248
use NAND2X1  _5073_
timestamp 0
transform 1 0 7350 0 -1 5530
box -6 -8 86 248
use INVX4  _5074_
timestamp 0
transform 1 0 4910 0 -1 4090
box -6 -8 86 248
use NAND2X1  _5075_
timestamp 0
transform 1 0 10310 0 1 6010
box -6 -8 86 248
use AND2X2  _5076_
timestamp 0
transform 1 0 10110 0 1 6010
box -6 -8 106 248
use NAND2X1  _5077_
timestamp 0
transform 1 0 9890 0 -1 6010
box -6 -8 86 248
use AOI22X1  _5078_
timestamp 0
transform 1 0 9670 0 -1 6010
box -6 -8 126 248
use OAI21X1  _5079_
timestamp 0
transform 1 0 10070 0 -1 6010
box -6 -8 106 248
use OAI21X1  _5080_
timestamp 0
transform 1 0 10270 0 -1 6010
box -6 -8 106 248
use OAI21X1  _5081_
timestamp 0
transform 1 0 10490 0 1 6010
box -6 -8 106 248
use AOI21X1  _5082_
timestamp 0
transform 1 0 10470 0 -1 6010
box -6 -8 106 248
use OR2X2  _5083_
timestamp 0
transform -1 0 10450 0 -1 5530
box -6 -8 106 248
use OAI21X1  _5084_
timestamp 0
transform -1 0 9830 0 1 5050
box -6 -8 106 248
use NAND2X1  _5085_
timestamp 0
transform 1 0 8590 0 1 5050
box -6 -8 86 248
use OAI21X1  _5086_
timestamp 0
transform -1 0 8870 0 1 5050
box -6 -8 106 248
use OR2X2  _5087_
timestamp 0
transform -1 0 11030 0 -1 5050
box -6 -8 106 248
use AOI22X1  _5088_
timestamp 0
transform -1 0 10830 0 -1 5050
box -6 -8 126 248
use OAI21X1  _5089_
timestamp 0
transform -1 0 10610 0 -1 5050
box -6 -8 106 248
use OAI21X1  _5090_
timestamp 0
transform -1 0 10390 0 1 5530
box -6 -8 106 248
use OAI21X1  _5091_
timestamp 0
transform 1 0 10150 0 -1 5530
box -6 -8 106 248
use NAND2X1  _5092_
timestamp 0
transform 1 0 9970 0 -1 5050
box -6 -8 86 248
use INVX1  _5093_
timestamp 0
transform -1 0 10210 0 -1 5050
box -6 -8 66 248
use NAND3X1  _5094_
timestamp 0
transform 1 0 10310 0 -1 5050
box -6 -8 106 248
use NAND2X1  _5095_
timestamp 0
transform -1 0 9890 0 -1 5050
box -6 -8 86 248
use NAND2X1  _5096_
timestamp 0
transform 1 0 8970 0 -1 5050
box -6 -8 86 248
use OAI21X1  _5097_
timestamp 0
transform 1 0 8290 0 -1 5050
box -6 -8 106 248
use NAND2X1  _5098_
timestamp 0
transform 1 0 9790 0 1 4570
box -6 -8 86 248
use OAI21X1  _5099_
timestamp 0
transform 1 0 9970 0 1 4570
box -6 -8 106 248
use NAND2X1  _5100_
timestamp 0
transform 1 0 9410 0 1 4570
box -6 -8 86 248
use NOR2X1  _5101_
timestamp 0
transform -1 0 10190 0 1 5530
box -6 -8 86 248
use INVX1  _5102_
timestamp 0
transform -1 0 9990 0 1 5050
box -6 -8 66 248
use AOI22X1  _5103_
timestamp 0
transform 1 0 10090 0 1 5050
box -6 -8 126 248
use NAND2X1  _5104_
timestamp 0
transform -1 0 10450 0 1 4570
box -6 -8 86 248
use OAI21X1  _5105_
timestamp 0
transform -1 0 10270 0 1 4570
box -6 -8 106 248
use NAND2X1  _5106_
timestamp 0
transform -1 0 10630 0 1 4570
box -6 -8 86 248
use OR2X2  _5107_
timestamp 0
transform 1 0 10550 0 -1 4570
box -6 -8 106 248
use AOI21X1  _5108_
timestamp 0
transform -1 0 11230 0 -1 4570
box -6 -8 106 248
use AOI22X1  _5109_
timestamp 0
transform 1 0 10750 0 -1 4570
box -6 -8 126 248
use OAI21X1  _5110_
timestamp 0
transform -1 0 9690 0 1 4570
box -6 -8 106 248
use NAND2X1  _5111_
timestamp 0
transform -1 0 8030 0 1 5530
box -6 -8 86 248
use OAI21X1  _5112_
timestamp 0
transform -1 0 8210 0 1 5530
box -6 -8 106 248
use DFFSR  _5113_
timestamp 0
transform -1 0 8890 0 -1 4090
box -6 -8 486 248
use DFFSR  _5114_
timestamp 0
transform -1 0 8730 0 1 6010
box -6 -8 486 248
use DFFSR  _5115_
timestamp 0
transform -1 0 7990 0 -1 5050
box -6 -8 486 248
use DFFSR  _5116_
timestamp 0
transform -1 0 8870 0 -1 5050
box -6 -8 486 248
use DFFSR  _5117_
timestamp 0
transform -1 0 9970 0 -1 4570
box -6 -8 486 248
use DFFSR  _5118_
timestamp 0
transform -1 0 8310 0 1 5050
box -6 -8 486 248
use DFFSR  _5119_
timestamp 0
transform -1 0 8910 0 1 4090
box -6 -8 486 248
use DFFSR  _5120_
timestamp 0
transform 1 0 9970 0 -1 4570
box -6 -8 486 248
use DFFSR  _5121_
timestamp 0
transform -1 0 7830 0 1 5050
box -6 -8 486 248
use DFFSR  _5122_
timestamp 0
transform -1 0 9710 0 -1 5050
box -6 -8 486 248
use DFFSR  _5123_
timestamp 0
transform -1 0 8910 0 -1 4570
box -6 -8 486 248
use NAND2X1  _5124_
timestamp 0
transform 1 0 1830 0 -1 1690
box -6 -8 86 248
use NAND2X1  _5125_
timestamp 0
transform -1 0 750 0 1 1690
box -6 -8 86 248
use NOR2X1  _5126_
timestamp 0
transform -1 0 930 0 1 1690
box -6 -8 86 248
use AND2X2  _5127_
timestamp 0
transform 1 0 830 0 1 2170
box -6 -8 106 248
use AND2X2  _5128_
timestamp 0
transform 1 0 590 0 -1 2170
box -6 -8 106 248
use AND2X2  _5129_
timestamp 0
transform 1 0 1030 0 1 2170
box -6 -8 106 248
use NAND2X1  _5130_
timestamp 0
transform 1 0 1030 0 1 1690
box -6 -8 86 248
use INVX4  _5131_
timestamp 0
transform -1 0 2410 0 -1 730
box -6 -8 86 248
use NAND2X1  _5132_
timestamp 0
transform -1 0 5650 0 -1 730
box -6 -8 86 248
use INVX1  _5133_
timestamp 0
transform 1 0 5330 0 -1 250
box -6 -8 66 248
use INVX1  _5134_
timestamp 0
transform 1 0 1410 0 1 1690
box -6 -8 66 248
use NOR2X1  _5135_
timestamp 0
transform 1 0 2210 0 -1 1690
box -6 -8 86 248
use NAND3X1  _5136_
timestamp 0
transform 1 0 2010 0 -1 1690
box -6 -8 106 248
use NOR2X1  _5137_
timestamp 0
transform -1 0 1210 0 -1 2170
box -6 -8 86 248
use NAND2X1  _5138_
timestamp 0
transform -1 0 1390 0 -1 2170
box -6 -8 86 248
use NOR2X1  _5139_
timestamp 0
transform -1 0 3770 0 -1 730
box -6 -8 86 248
use INVX1  _5140_
timestamp 0
transform 1 0 4170 0 -1 1690
box -6 -8 66 248
use NOR2X1  _5141_
timestamp 0
transform -1 0 4410 0 -1 1690
box -6 -8 86 248
use NAND3X1  _5142_
timestamp 0
transform -1 0 4310 0 1 1210
box -6 -8 106 248
use INVX1  _5143_
timestamp 0
transform -1 0 4470 0 -1 730
box -6 -8 66 248
use NOR2X1  _5144_
timestamp 0
transform 1 0 5610 0 1 730
box -6 -8 86 248
use INVX1  _5145_
timestamp 0
transform -1 0 4190 0 1 730
box -6 -8 66 248
use NOR2X1  _5146_
timestamp 0
transform -1 0 4730 0 1 730
box -6 -8 86 248
use NAND3X1  _5147_
timestamp 0
transform 1 0 4770 0 -1 730
box -6 -8 106 248
use NOR2X1  _5148_
timestamp 0
transform 1 0 4970 0 -1 730
box -6 -8 86 248
use NAND3X1  _5149_
timestamp 0
transform 1 0 5490 0 -1 250
box -6 -8 106 248
use INVX1  _5150_
timestamp 0
transform -1 0 6150 0 -1 250
box -6 -8 66 248
use OR2X2  _5151_
timestamp 0
transform 1 0 3490 0 -1 730
box -6 -8 106 248
use INVX1  _5152_
timestamp 0
transform 1 0 5750 0 1 250
box -6 -8 66 248
use INVX1  _5153_
timestamp 0
transform 1 0 4230 0 -1 1210
box -6 -8 66 248
use NAND2X1  _5154_
timestamp 0
transform 1 0 5430 0 1 730
box -6 -8 86 248
use NOR2X1  _5155_
timestamp 0
transform 1 0 5390 0 -1 730
box -6 -8 86 248
use NAND3X1  _5156_
timestamp 0
transform 1 0 5550 0 1 250
box -6 -8 106 248
use OAI21X1  _5157_
timestamp 0
transform 1 0 5690 0 -1 250
box -6 -8 106 248
use NAND3X1  _5158_
timestamp 0
transform 1 0 4570 0 -1 730
box -6 -8 106 248
use NOR2X1  _5159_
timestamp 0
transform -1 0 4750 0 1 250
box -6 -8 86 248
use NAND2X1  _5160_
timestamp 0
transform 1 0 5010 0 1 250
box -6 -8 86 248
use INVX2  _5161_
timestamp 0
transform 1 0 4850 0 1 250
box -6 -8 66 248
use AOI21X1  _5162_
timestamp 0
transform 1 0 5890 0 -1 250
box -6 -8 106 248
use OAI21X1  _5163_
timestamp 0
transform -1 0 2850 0 1 250
box -6 -8 106 248
use OAI21X1  _5164_
timestamp 0
transform 1 0 5910 0 1 250
box -6 -8 106 248
use INVX1  _5165_
timestamp 0
transform -1 0 3890 0 1 1690
box -6 -8 66 248
use NAND2X1  _5166_
timestamp 0
transform 1 0 4290 0 1 730
box -6 -8 86 248
use NOR2X1  _5167_
timestamp 0
transform 1 0 4250 0 -1 730
box -6 -8 86 248
use NAND3X1  _5168_
timestamp 0
transform -1 0 4150 0 -1 730
box -6 -8 106 248
use INVX1  _5169_
timestamp 0
transform 1 0 2750 0 -1 1690
box -6 -8 66 248
use NOR2X1  _5170_
timestamp 0
transform 1 0 3870 0 -1 730
box -6 -8 86 248
use INVX1  _5171_
timestamp 0
transform -1 0 4210 0 1 1690
box -6 -8 66 248
use NOR2X1  _5172_
timestamp 0
transform -1 0 3730 0 1 1690
box -6 -8 86 248
use NOR3X1  _5173_
timestamp 0
transform -1 0 5110 0 -1 1210
box -6 -8 186 248
use NAND3X1  _5174_
timestamp 0
transform -1 0 3930 0 -1 1210
box -6 -8 106 248
use NOR3X1  _5175_
timestamp 0
transform 1 0 3690 0 1 730
box -6 -8 186 248
use NAND3X1  _5176_
timestamp 0
transform -1 0 2770 0 -1 1210
box -6 -8 106 248
use INVX1  _5177_
timestamp 0
transform 1 0 3130 0 -1 250
box -6 -8 66 248
use NAND2X1  _5178_
timestamp 0
transform 1 0 4470 0 1 730
box -6 -8 86 248
use NOR2X1  _5179_
timestamp 0
transform 1 0 4490 0 1 250
box -6 -8 86 248
use NAND3X1  _5180_
timestamp 0
transform 1 0 4290 0 1 250
box -6 -8 106 248
use NAND2X1  _5181_
timestamp 0
transform 1 0 3290 0 -1 250
box -6 -8 86 248
use NAND3X1  _5182_
timestamp 0
transform -1 0 2570 0 -1 1210
box -6 -8 106 248
use AOI21X1  _5183_
timestamp 0
transform 1 0 2270 0 -1 1210
box -6 -8 106 248
use AOI22X1  _5184_
timestamp 0
transform -1 0 2610 0 1 1210
box -6 -8 126 248
use INVX1  _5185_
timestamp 0
transform -1 0 4110 0 1 1210
box -6 -8 66 248
use INVX1  _5186_
timestamp 0
transform -1 0 3390 0 1 1210
box -6 -8 66 248
use NAND3X1  _5187_
timestamp 0
transform -1 0 3170 0 -1 1210
box -6 -8 106 248
use INVX1  _5188_
timestamp 0
transform 1 0 3790 0 -1 250
box -6 -8 66 248
use NAND2X1  _5189_
timestamp 0
transform -1 0 3790 0 1 250
box -6 -8 86 248
use NAND3X1  _5190_
timestamp 0
transform 1 0 3270 0 -1 1210
box -6 -8 106 248
use AOI21X1  _5191_
timestamp 0
transform 1 0 2950 0 1 250
box -6 -8 106 248
use AOI22X1  _5192_
timestamp 0
transform -1 0 3770 0 1 1210
box -6 -8 126 248
use INVX1  _5193_
timestamp 0
transform 1 0 6110 0 1 250
box -6 -8 66 248
use INVX1  _5194_
timestamp 0
transform -1 0 3010 0 1 1210
box -6 -8 66 248
use NAND3X1  _5195_
timestamp 0
transform -1 0 2970 0 -1 1210
box -6 -8 106 248
use INVX1  _5196_
timestamp 0
transform 1 0 3630 0 -1 250
box -6 -8 66 248
use NAND2X1  _5197_
timestamp 0
transform -1 0 3610 0 1 250
box -6 -8 86 248
use NAND3X1  _5198_
timestamp 0
transform -1 0 3030 0 -1 730
box -6 -8 106 248
use AOI21X1  _5199_
timestamp 0
transform 1 0 2510 0 -1 730
box -6 -8 106 248
use AOI22X1  _5200_
timestamp 0
transform -1 0 2830 0 -1 730
box -6 -8 126 248
use INVX1  _5201_
timestamp 0
transform -1 0 4050 0 1 1690
box -6 -8 66 248
use INVX1  _5202_
timestamp 0
transform 1 0 3970 0 1 730
box -6 -8 66 248
use NAND3X1  _5203_
timestamp 0
transform -1 0 3590 0 1 730
box -6 -8 106 248
use INVX1  _5204_
timestamp 0
transform 1 0 4110 0 -1 250
box -6 -8 66 248
use NAND2X1  _5205_
timestamp 0
transform -1 0 4030 0 -1 250
box -6 -8 86 248
use NAND3X1  _5206_
timestamp 0
transform -1 0 3390 0 1 730
box -6 -8 106 248
use AOI21X1  _5207_
timestamp 0
transform 1 0 2530 0 1 730
box -6 -8 106 248
use AOI22X1  _5208_
timestamp 0
transform 1 0 3070 0 -1 1690
box -6 -8 126 248
use INVX1  _5209_
timestamp 0
transform -1 0 4570 0 -1 1690
box -6 -8 66 248
use INVX1  _5210_
timestamp 0
transform 1 0 2730 0 1 730
box -6 -8 66 248
use NAND3X1  _5211_
timestamp 0
transform 1 0 2890 0 1 730
box -6 -8 106 248
use INVX1  _5212_
timestamp 0
transform 1 0 3470 0 -1 250
box -6 -8 66 248
use NAND2X1  _5213_
timestamp 0
transform 1 0 3350 0 1 250
box -6 -8 86 248
use NAND3X1  _5214_
timestamp 0
transform -1 0 3190 0 1 730
box -6 -8 106 248
use AOI21X1  _5215_
timestamp 0
transform 1 0 2330 0 1 730
box -6 -8 106 248
use AOI22X1  _5216_
timestamp 0
transform -1 0 3230 0 1 1210
box -6 -8 126 248
use INVX1  _5217_
timestamp 0
transform -1 0 6330 0 1 250
box -6 -8 66 248
use INVX1  _5218_
timestamp 0
transform 1 0 3470 0 -1 1210
box -6 -8 66 248
use NAND3X1  _5219_
timestamp 0
transform 1 0 3630 0 -1 1210
box -6 -8 106 248
use INVX1  _5220_
timestamp 0
transform 1 0 4810 0 -1 250
box -6 -8 66 248
use NAND2X1  _5221_
timestamp 0
transform 1 0 4630 0 -1 250
box -6 -8 86 248
use NAND3X1  _5222_
timestamp 0
transform -1 0 4190 0 1 250
box -6 -8 106 248
use AOI21X1  _5223_
timestamp 0
transform 1 0 3150 0 1 250
box -6 -8 106 248
use AOI22X1  _5224_
timestamp 0
transform -1 0 3990 0 1 250
box -6 -8 126 248
use INVX1  _5225_
timestamp 0
transform 1 0 5410 0 1 1210
box -6 -8 66 248
use INVX1  _5226_
timestamp 0
transform 1 0 5190 0 1 250
box -6 -8 66 248
use OAI21X1  _5227_
timestamp 0
transform -1 0 5450 0 1 250
box -6 -8 106 248
use INVX1  _5228_
timestamp 0
transform -1 0 4850 0 -1 2170
box -6 -8 66 248
use NAND3X1  _5229_
timestamp 0
transform -1 0 4930 0 1 730
box -6 -8 106 248
use NAND3X1  _5230_
timestamp 0
transform 1 0 5030 0 1 730
box -6 -8 106 248
use NAND3X1  _5231_
timestamp 0
transform 1 0 5230 0 1 730
box -6 -8 106 248
use OR2X2  _5232_
timestamp 0
transform 1 0 4030 0 -1 1210
box -6 -8 106 248
use AOI21X1  _5233_
timestamp 0
transform 1 0 4410 0 1 1210
box -6 -8 106 248
use AOI22X1  _5234_
timestamp 0
transform -1 0 5310 0 1 1210
box -6 -8 126 248
use DFFPOSX1  _5235_
timestamp 0
transform -1 0 4690 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _5236_
timestamp 0
transform -1 0 2690 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _5237_
timestamp 0
transform -1 0 5930 0 1 730
box -6 -8 246 248
use DFFPOSX1  _5238_
timestamp 0
transform 1 0 550 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _5239_
timestamp 0
transform 1 0 310 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _5240_
timestamp 0
transform -1 0 2850 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _5241_
timestamp 0
transform -1 0 5090 0 -1 2170
box -6 -8 246 248
use DFFSR  _5242_
timestamp 0
transform 1 0 1650 0 1 1690
box -6 -8 486 248
use DFFSR  _5243_
timestamp 0
transform 1 0 2550 0 -1 250
box -6 -8 486 248
use DFFPOSX1  _5244_
timestamp 0
transform -1 0 5530 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _5245_
timestamp 0
transform -1 0 5290 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _5246_
timestamp 0
transform -1 0 5170 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _5247_
timestamp 0
transform -1 0 3970 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _5248_
timestamp 0
transform -1 0 3730 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _5249_
timestamp 0
transform -1 0 5770 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _5250_
timestamp 0
transform -1 0 430 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _5251_
timestamp 0
transform -1 0 1630 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _5252_
timestamp 0
transform -1 0 2370 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _5253_
timestamp 0
transform -1 0 1030 0 -1 2650
box -6 -8 246 248
use DFFSR  _5254_
timestamp 0
transform 1 0 2370 0 -1 3610
box -6 -8 486 248
use BUFX2  BUFX2_insert0
timestamp 0
transform -1 0 4310 0 1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert1
timestamp 0
transform 1 0 6170 0 -1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert2
timestamp 0
transform -1 0 3410 0 1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert3
timestamp 0
transform -1 0 3790 0 1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert4
timestamp 0
transform 1 0 9510 0 1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert5
timestamp 0
transform 1 0 11310 0 1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert6
timestamp 0
transform -1 0 9570 0 1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert7
timestamp 0
transform 1 0 12050 0 1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert8
timestamp 0
transform -1 0 7270 0 1 5530
box -6 -8 86 248
use BUFX2  BUFX2_insert9
timestamp 0
transform 1 0 6690 0 -1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert10
timestamp 0
transform 1 0 8750 0 -1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert11
timestamp 0
transform 1 0 6910 0 -1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert12
timestamp 0
transform 1 0 8950 0 1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert13
timestamp 0
transform 1 0 7430 0 1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert14
timestamp 0
transform 1 0 690 0 -1 6970
box -6 -8 86 248
use BUFX2  BUFX2_insert15
timestamp 0
transform 1 0 110 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert16
timestamp 0
transform 1 0 1930 0 1 5530
box -6 -8 86 248
use BUFX2  BUFX2_insert17
timestamp 0
transform -1 0 9250 0 -1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert18
timestamp 0
transform -1 0 11610 0 -1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert19
timestamp 0
transform 1 0 10710 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert20
timestamp 0
transform -1 0 9290 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert21
timestamp 0
transform 1 0 2570 0 1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert22
timestamp 0
transform -1 0 1370 0 1 11290
box -6 -8 86 248
use BUFX2  BUFX2_insert23
timestamp 0
transform -1 0 1550 0 1 11290
box -6 -8 86 248
use BUFX2  BUFX2_insert24
timestamp 0
transform -1 0 1750 0 1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert38
timestamp 0
transform -1 0 11630 0 -1 6490
box -6 -8 86 248
use BUFX2  BUFX2_insert39
timestamp 0
transform -1 0 10770 0 1 6010
box -6 -8 86 248
use BUFX2  BUFX2_insert40
timestamp 0
transform 1 0 12070 0 1 6970
box -6 -8 86 248
use BUFX2  BUFX2_insert41
timestamp 0
transform -1 0 11350 0 1 6010
box -6 -8 86 248
use BUFX2  BUFX2_insert42
timestamp 0
transform 1 0 11490 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert43
timestamp 0
transform -1 0 11110 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert44
timestamp 0
transform -1 0 10590 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert45
timestamp 0
transform -1 0 11470 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert46
timestamp 0
transform -1 0 10850 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert47
timestamp 0
transform 1 0 6250 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert48
timestamp 0
transform -1 0 4870 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert49
timestamp 0
transform 1 0 11590 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert50
timestamp 0
transform -1 0 10510 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert51
timestamp 0
transform 1 0 8210 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert52
timestamp 0
transform 1 0 10070 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert53
timestamp 0
transform 1 0 9230 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert54
timestamp 0
transform 1 0 9050 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert55
timestamp 0
transform -1 0 9650 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert56
timestamp 0
transform -1 0 8950 0 1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert57
timestamp 0
transform 1 0 11510 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert58
timestamp 0
transform 1 0 10690 0 -1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert59
timestamp 0
transform -1 0 7830 0 -1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert60
timestamp 0
transform 1 0 11850 0 -1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert61
timestamp 0
transform 1 0 11950 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert62
timestamp 0
transform -1 0 4910 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert63
timestamp 0
transform -1 0 9430 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert64
timestamp 0
transform -1 0 11770 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert65
timestamp 0
transform -1 0 9430 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert66
timestamp 0
transform -1 0 11610 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert67
timestamp 0
transform 1 0 6970 0 1 11290
box -6 -8 86 248
use BUFX2  BUFX2_insert68
timestamp 0
transform -1 0 3270 0 -1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert69
timestamp 0
transform -1 0 5710 0 1 10810
box -6 -8 86 248
use BUFX2  BUFX2_insert70
timestamp 0
transform 1 0 5150 0 -1 11290
box -6 -8 86 248
use BUFX2  BUFX2_insert71
timestamp 0
transform -1 0 3670 0 -1 10810
box -6 -8 86 248
use BUFX2  BUFX2_insert72
timestamp 0
transform 1 0 7150 0 1 11290
box -6 -8 86 248
use BUFX2  BUFX2_insert73
timestamp 0
transform 1 0 7170 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert74
timestamp 0
transform -1 0 6570 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert75
timestamp 0
transform 1 0 7130 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert76
timestamp 0
transform 1 0 6590 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert77
timestamp 0
transform 1 0 10310 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert78
timestamp 0
transform 1 0 9170 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert79
timestamp 0
transform 1 0 10330 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert80
timestamp 0
transform -1 0 5050 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert81
timestamp 0
transform -1 0 2910 0 1 5530
box -6 -8 86 248
use BUFX2  BUFX2_insert82
timestamp 0
transform -1 0 4130 0 -1 5530
box -6 -8 86 248
use BUFX2  BUFX2_insert83
timestamp 0
transform -1 0 6390 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert84
timestamp 0
transform 1 0 7390 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert85
timestamp 0
transform -1 0 3370 0 1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert86
timestamp 0
transform 1 0 4010 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert87
timestamp 0
transform -1 0 3330 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert88
timestamp 0
transform 1 0 7930 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert89
timestamp 0
transform -1 0 4810 0 1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert90
timestamp 0
transform 1 0 5610 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert91
timestamp 0
transform 1 0 9070 0 1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert92
timestamp 0
transform -1 0 8630 0 1 10810
box -6 -8 86 248
use BUFX2  BUFX2_insert93
timestamp 0
transform -1 0 11030 0 -1 10810
box -6 -8 86 248
use BUFX2  BUFX2_insert94
timestamp 0
transform 1 0 7310 0 1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert95
timestamp 0
transform 1 0 11570 0 1 10810
box -6 -8 86 248
use BUFX2  BUFX2_insert96
timestamp 0
transform -1 0 5090 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert97
timestamp 0
transform 1 0 650 0 -1 6010
box -6 -8 86 248
use BUFX2  BUFX2_insert98
timestamp 0
transform -1 0 4110 0 1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert99
timestamp 0
transform 1 0 590 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert100
timestamp 0
transform 1 0 3070 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert101
timestamp 0
transform -1 0 590 0 -1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert102
timestamp 0
transform 1 0 3770 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert103
timestamp 0
transform -1 0 3750 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert104
timestamp 0
transform 1 0 4670 0 1 10330
box -6 -8 86 248
use BUFX2  BUFX2_insert105
timestamp 0
transform 1 0 330 0 -1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert106
timestamp 0
transform 1 0 6550 0 -1 10810
box -6 -8 86 248
use BUFX2  BUFX2_insert107
timestamp 0
transform -1 0 6310 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert108
timestamp 0
transform 1 0 5730 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert109
timestamp 0
transform 1 0 7850 0 -1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert110
timestamp 0
transform -1 0 5430 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert111
timestamp 0
transform 1 0 7330 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert112
timestamp 0
transform 1 0 10710 0 1 11770
box -6 -8 86 248
use BUFX2  BUFX2_insert113
timestamp 0
transform -1 0 12210 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert114
timestamp 0
transform -1 0 10410 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert115
timestamp 0
transform 1 0 7410 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert116
timestamp 0
transform -1 0 5610 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert117
timestamp 0
transform -1 0 5590 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert118
timestamp 0
transform -1 0 11290 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert119
timestamp 0
transform 1 0 10410 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert120
timestamp 0
transform -1 0 11210 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert121
timestamp 0
transform -1 0 8270 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert122
timestamp 0
transform 1 0 11230 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert123
timestamp 0
transform -1 0 10130 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert124
timestamp 0
transform -1 0 8110 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert125
timestamp 0
transform -1 0 5430 0 1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert126
timestamp 0
transform 1 0 12050 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert127
timestamp 0
transform 1 0 10810 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert128
timestamp 0
transform -1 0 12150 0 -1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert129
timestamp 0
transform 1 0 10470 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert130
timestamp 0
transform 1 0 12050 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert131
timestamp 0
transform -1 0 9470 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert132
timestamp 0
transform -1 0 8810 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert133
timestamp 0
transform 1 0 12050 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert134
timestamp 0
transform -1 0 11490 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert135
timestamp 0
transform -1 0 9210 0 -1 250
box -6 -8 86 248
use BUFX2  BUFX2_insert136
timestamp 0
transform 1 0 9510 0 -1 250
box -6 -8 86 248
use BUFX2  BUFX2_insert137
timestamp 0
transform -1 0 6490 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert138
timestamp 0
transform 1 0 8410 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert139
timestamp 0
transform -1 0 6510 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert140
timestamp 0
transform 1 0 9470 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert141
timestamp 0
transform -1 0 7150 0 -1 6970
box -6 -8 86 248
use BUFX2  BUFX2_insert142
timestamp 0
transform -1 0 7130 0 1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert143
timestamp 0
transform -1 0 6550 0 -1 6970
box -6 -8 86 248
use BUFX2  BUFX2_insert144
timestamp 0
transform -1 0 6370 0 1 6970
box -6 -8 86 248
use BUFX2  BUFX2_insert145
timestamp 0
transform 1 0 9590 0 -1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert146
timestamp 0
transform 1 0 9690 0 1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert147
timestamp 0
transform -1 0 7830 0 1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert148
timestamp 0
transform -1 0 7750 0 -1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert149
timestamp 0
transform -1 0 9310 0 -1 7930
box -6 -8 86 248
use BUFX2  BUFX2_insert150
timestamp 0
transform -1 0 7330 0 -1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert151
timestamp 0
transform 1 0 7370 0 -1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert152
timestamp 0
transform -1 0 8330 0 1 9370
box -6 -8 86 248
use BUFX2  BUFX2_insert153
timestamp 0
transform 1 0 10110 0 -1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert154
timestamp 0
transform 1 0 10790 0 -1 8410
box -6 -8 86 248
use BUFX2  BUFX2_insert155
timestamp 0
transform 1 0 6430 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert156
timestamp 0
transform 1 0 9170 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert157
timestamp 0
transform -1 0 5970 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert158
timestamp 0
transform 1 0 9910 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert159
timestamp 0
transform 1 0 8770 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert160
timestamp 0
transform 1 0 10410 0 1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert161
timestamp 0
transform 1 0 9310 0 1 9850
box -6 -8 86 248
use BUFX2  BUFX2_insert162
timestamp 0
transform 1 0 10270 0 1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert163
timestamp 0
transform -1 0 8430 0 1 8890
box -6 -8 86 248
use BUFX2  BUFX2_insert164
timestamp 0
transform 1 0 11770 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert165
timestamp 0
transform -1 0 8890 0 -1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert166
timestamp 0
transform -1 0 11670 0 1 4090
box -6 -8 86 248
use BUFX2  BUFX2_insert167
timestamp 0
transform 1 0 11770 0 1 11770
box -6 -8 86 248
use BUFX2  BUFX2_insert168
timestamp 0
transform -1 0 11410 0 -1 2170
box -6 -8 86 248
use BUFX2  BUFX2_insert169
timestamp 0
transform 1 0 4970 0 1 1690
box -6 -8 86 248
use CLKBUF1  CLKBUF1_insert25
timestamp 0
transform 1 0 1410 0 1 2170
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert26
timestamp 0
transform 1 0 4070 0 -1 2170
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert27
timestamp 0
transform -1 0 310 0 -1 2650
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert28
timestamp 0
transform -1 0 2950 0 1 9370
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert29
timestamp 0
transform 1 0 90 0 -1 2170
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert30
timestamp 0
transform 1 0 6230 0 -1 5050
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert31
timestamp 0
transform 1 0 830 0 -1 6010
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert32
timestamp 0
transform -1 0 5050 0 -1 3610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert33
timestamp 0
transform -1 0 1190 0 -1 10810
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert34
timestamp 0
transform 1 0 1450 0 -1 6490
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert35
timestamp 0
transform -1 0 550 0 -1 11770
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert36
timestamp 0
transform 1 0 110 0 1 5530
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert37
timestamp 0
transform 1 0 6190 0 1 11770
box -6 -8 206 248
use FILL  FILL180450x21750
timestamp 0
transform -1 0 12050 0 -1 1690
box -6 -8 26 248
use FILL  FILL180450x28950
timestamp 0
transform -1 0 12050 0 -1 2170
box -6 -8 26 248
use FILL  FILL180450x176550
timestamp 0
transform 1 0 12030 0 1 11770
box -6 -8 26 248
use FILL  FILL180750x150
timestamp 0
transform -1 0 12070 0 -1 250
box -6 -8 26 248
use FILL  FILL180750x21750
timestamp 0
transform -1 0 12070 0 -1 1690
box -6 -8 26 248
use FILL  FILL180750x28950
timestamp 0
transform -1 0 12070 0 -1 2170
box -6 -8 26 248
use FILL  FILL180750x176550
timestamp 0
transform 1 0 12050 0 1 11770
box -6 -8 26 248
use FILL  FILL181050x150
timestamp 0
transform -1 0 12090 0 -1 250
box -6 -8 26 248
use FILL  FILL181050x21750
timestamp 0
transform -1 0 12090 0 -1 1690
box -6 -8 26 248
use FILL  FILL181050x28950
timestamp 0
transform -1 0 12090 0 -1 2170
box -6 -8 26 248
use FILL  FILL181050x61350
timestamp 0
transform 1 0 12070 0 1 4090
box -6 -8 26 248
use FILL  FILL181050x111750
timestamp 0
transform 1 0 12070 0 1 7450
box -6 -8 26 248
use FILL  FILL181050x176550
timestamp 0
transform 1 0 12070 0 1 11770
box -6 -8 26 248
use FILL  FILL181350x150
timestamp 0
transform -1 0 12110 0 -1 250
box -6 -8 26 248
use FILL  FILL181350x3750
timestamp 0
transform 1 0 12090 0 1 250
box -6 -8 26 248
use FILL  FILL181350x21750
timestamp 0
transform -1 0 12110 0 -1 1690
box -6 -8 26 248
use FILL  FILL181350x25350
timestamp 0
transform 1 0 12090 0 1 1690
box -6 -8 26 248
use FILL  FILL181350x28950
timestamp 0
transform -1 0 12110 0 -1 2170
box -6 -8 26 248
use FILL  FILL181350x50550
timestamp 0
transform -1 0 12110 0 -1 3610
box -6 -8 26 248
use FILL  FILL181350x61350
timestamp 0
transform 1 0 12090 0 1 4090
box -6 -8 26 248
use FILL  FILL181350x111750
timestamp 0
transform 1 0 12090 0 1 7450
box -6 -8 26 248
use FILL  FILL181350x176550
timestamp 0
transform 1 0 12090 0 1 11770
box -6 -8 26 248
use FILL  FILL181650x150
timestamp 0
transform -1 0 12130 0 -1 250
box -6 -8 26 248
use FILL  FILL181650x3750
timestamp 0
transform 1 0 12110 0 1 250
box -6 -8 26 248
use FILL  FILL181650x7350
timestamp 0
transform -1 0 12130 0 -1 730
box -6 -8 26 248
use FILL  FILL181650x14550
timestamp 0
transform -1 0 12130 0 -1 1210
box -6 -8 26 248
use FILL  FILL181650x21750
timestamp 0
transform -1 0 12130 0 -1 1690
box -6 -8 26 248
use FILL  FILL181650x25350
timestamp 0
transform 1 0 12110 0 1 1690
box -6 -8 26 248
use FILL  FILL181650x28950
timestamp 0
transform -1 0 12130 0 -1 2170
box -6 -8 26 248
use FILL  FILL181650x50550
timestamp 0
transform -1 0 12130 0 -1 3610
box -6 -8 26 248
use FILL  FILL181650x61350
timestamp 0
transform 1 0 12110 0 1 4090
box -6 -8 26 248
use FILL  FILL181650x72150
timestamp 0
transform -1 0 12130 0 -1 5050
box -6 -8 26 248
use FILL  FILL181650x82950
timestamp 0
transform 1 0 12110 0 1 5530
box -6 -8 26 248
use FILL  FILL181650x111750
timestamp 0
transform 1 0 12110 0 1 7450
box -6 -8 26 248
use FILL  FILL181650x154950
timestamp 0
transform 1 0 12110 0 1 10330
box -6 -8 26 248
use FILL  FILL181650x176550
timestamp 0
transform 1 0 12110 0 1 11770
box -6 -8 26 248
use FILL  FILL181950x150
timestamp 0
transform -1 0 12150 0 -1 250
box -6 -8 26 248
use FILL  FILL181950x3750
timestamp 0
transform 1 0 12130 0 1 250
box -6 -8 26 248
use FILL  FILL181950x7350
timestamp 0
transform -1 0 12150 0 -1 730
box -6 -8 26 248
use FILL  FILL181950x10950
timestamp 0
transform 1 0 12130 0 1 730
box -6 -8 26 248
use FILL  FILL181950x14550
timestamp 0
transform -1 0 12150 0 -1 1210
box -6 -8 26 248
use FILL  FILL181950x21750
timestamp 0
transform -1 0 12150 0 -1 1690
box -6 -8 26 248
use FILL  FILL181950x25350
timestamp 0
transform 1 0 12130 0 1 1690
box -6 -8 26 248
use FILL  FILL181950x28950
timestamp 0
transform -1 0 12150 0 -1 2170
box -6 -8 26 248
use FILL  FILL181950x32550
timestamp 0
transform 1 0 12130 0 1 2170
box -6 -8 26 248
use FILL  FILL181950x36150
timestamp 0
transform -1 0 12150 0 -1 2650
box -6 -8 26 248
use FILL  FILL181950x50550
timestamp 0
transform -1 0 12150 0 -1 3610
box -6 -8 26 248
use FILL  FILL181950x61350
timestamp 0
transform 1 0 12130 0 1 4090
box -6 -8 26 248
use FILL  FILL181950x64950
timestamp 0
transform -1 0 12150 0 -1 4570
box -6 -8 26 248
use FILL  FILL181950x68550
timestamp 0
transform 1 0 12130 0 1 4570
box -6 -8 26 248
use FILL  FILL181950x72150
timestamp 0
transform -1 0 12150 0 -1 5050
box -6 -8 26 248
use FILL  FILL181950x82950
timestamp 0
transform 1 0 12130 0 1 5530
box -6 -8 26 248
use FILL  FILL181950x86550
timestamp 0
transform -1 0 12150 0 -1 6010
box -6 -8 26 248
use FILL  FILL181950x90150
timestamp 0
transform 1 0 12130 0 1 6010
box -6 -8 26 248
use FILL  FILL181950x108150
timestamp 0
transform -1 0 12150 0 -1 7450
box -6 -8 26 248
use FILL  FILL181950x111750
timestamp 0
transform 1 0 12130 0 1 7450
box -6 -8 26 248
use FILL  FILL181950x118950
timestamp 0
transform 1 0 12130 0 1 7930
box -6 -8 26 248
use FILL  FILL181950x122550
timestamp 0
transform -1 0 12150 0 -1 8410
box -6 -8 26 248
use FILL  FILL181950x126150
timestamp 0
transform 1 0 12130 0 1 8410
box -6 -8 26 248
use FILL  FILL181950x140550
timestamp 0
transform 1 0 12130 0 1 9370
box -6 -8 26 248
use FILL  FILL181950x147750
timestamp 0
transform 1 0 12130 0 1 9850
box -6 -8 26 248
use FILL  FILL181950x154950
timestamp 0
transform 1 0 12130 0 1 10330
box -6 -8 26 248
use FILL  FILL181950x162150
timestamp 0
transform 1 0 12130 0 1 10810
box -6 -8 26 248
use FILL  FILL181950x176550
timestamp 0
transform 1 0 12130 0 1 11770
box -6 -8 26 248
use FILL  FILL182250x150
timestamp 0
transform -1 0 12170 0 -1 250
box -6 -8 26 248
use FILL  FILL182250x3750
timestamp 0
transform 1 0 12150 0 1 250
box -6 -8 26 248
use FILL  FILL182250x7350
timestamp 0
transform -1 0 12170 0 -1 730
box -6 -8 26 248
use FILL  FILL182250x10950
timestamp 0
transform 1 0 12150 0 1 730
box -6 -8 26 248
use FILL  FILL182250x14550
timestamp 0
transform -1 0 12170 0 -1 1210
box -6 -8 26 248
use FILL  FILL182250x18150
timestamp 0
transform 1 0 12150 0 1 1210
box -6 -8 26 248
use FILL  FILL182250x21750
timestamp 0
transform -1 0 12170 0 -1 1690
box -6 -8 26 248
use FILL  FILL182250x25350
timestamp 0
transform 1 0 12150 0 1 1690
box -6 -8 26 248
use FILL  FILL182250x28950
timestamp 0
transform -1 0 12170 0 -1 2170
box -6 -8 26 248
use FILL  FILL182250x32550
timestamp 0
transform 1 0 12150 0 1 2170
box -6 -8 26 248
use FILL  FILL182250x36150
timestamp 0
transform -1 0 12170 0 -1 2650
box -6 -8 26 248
use FILL  FILL182250x43350
timestamp 0
transform -1 0 12170 0 -1 3130
box -6 -8 26 248
use FILL  FILL182250x46950
timestamp 0
transform 1 0 12150 0 1 3130
box -6 -8 26 248
use FILL  FILL182250x50550
timestamp 0
transform -1 0 12170 0 -1 3610
box -6 -8 26 248
use FILL  FILL182250x57750
timestamp 0
transform -1 0 12170 0 -1 4090
box -6 -8 26 248
use FILL  FILL182250x61350
timestamp 0
transform 1 0 12150 0 1 4090
box -6 -8 26 248
use FILL  FILL182250x64950
timestamp 0
transform -1 0 12170 0 -1 4570
box -6 -8 26 248
use FILL  FILL182250x68550
timestamp 0
transform 1 0 12150 0 1 4570
box -6 -8 26 248
use FILL  FILL182250x72150
timestamp 0
transform -1 0 12170 0 -1 5050
box -6 -8 26 248
use FILL  FILL182250x75750
timestamp 0
transform 1 0 12150 0 1 5050
box -6 -8 26 248
use FILL  FILL182250x82950
timestamp 0
transform 1 0 12150 0 1 5530
box -6 -8 26 248
use FILL  FILL182250x86550
timestamp 0
transform -1 0 12170 0 -1 6010
box -6 -8 26 248
use FILL  FILL182250x90150
timestamp 0
transform 1 0 12150 0 1 6010
box -6 -8 26 248
use FILL  FILL182250x104550
timestamp 0
transform 1 0 12150 0 1 6970
box -6 -8 26 248
use FILL  FILL182250x108150
timestamp 0
transform -1 0 12170 0 -1 7450
box -6 -8 26 248
use FILL  FILL182250x111750
timestamp 0
transform 1 0 12150 0 1 7450
box -6 -8 26 248
use FILL  FILL182250x115350
timestamp 0
transform -1 0 12170 0 -1 7930
box -6 -8 26 248
use FILL  FILL182250x118950
timestamp 0
transform 1 0 12150 0 1 7930
box -6 -8 26 248
use FILL  FILL182250x122550
timestamp 0
transform -1 0 12170 0 -1 8410
box -6 -8 26 248
use FILL  FILL182250x126150
timestamp 0
transform 1 0 12150 0 1 8410
box -6 -8 26 248
use FILL  FILL182250x133350
timestamp 0
transform 1 0 12150 0 1 8890
box -6 -8 26 248
use FILL  FILL182250x140550
timestamp 0
transform 1 0 12150 0 1 9370
box -6 -8 26 248
use FILL  FILL182250x144150
timestamp 0
transform -1 0 12170 0 -1 9850
box -6 -8 26 248
use FILL  FILL182250x147750
timestamp 0
transform 1 0 12150 0 1 9850
box -6 -8 26 248
use FILL  FILL182250x151350
timestamp 0
transform -1 0 12170 0 -1 10330
box -6 -8 26 248
use FILL  FILL182250x154950
timestamp 0
transform 1 0 12150 0 1 10330
box -6 -8 26 248
use FILL  FILL182250x162150
timestamp 0
transform 1 0 12150 0 1 10810
box -6 -8 26 248
use FILL  FILL182250x169350
timestamp 0
transform 1 0 12150 0 1 11290
box -6 -8 26 248
use FILL  FILL182250x176550
timestamp 0
transform 1 0 12150 0 1 11770
box -6 -8 26 248
use FILL  FILL182550x150
timestamp 0
transform -1 0 12190 0 -1 250
box -6 -8 26 248
use FILL  FILL182550x3750
timestamp 0
transform 1 0 12170 0 1 250
box -6 -8 26 248
use FILL  FILL182550x7350
timestamp 0
transform -1 0 12190 0 -1 730
box -6 -8 26 248
use FILL  FILL182550x10950
timestamp 0
transform 1 0 12170 0 1 730
box -6 -8 26 248
use FILL  FILL182550x14550
timestamp 0
transform -1 0 12190 0 -1 1210
box -6 -8 26 248
use FILL  FILL182550x18150
timestamp 0
transform 1 0 12170 0 1 1210
box -6 -8 26 248
use FILL  FILL182550x21750
timestamp 0
transform -1 0 12190 0 -1 1690
box -6 -8 26 248
use FILL  FILL182550x25350
timestamp 0
transform 1 0 12170 0 1 1690
box -6 -8 26 248
use FILL  FILL182550x28950
timestamp 0
transform -1 0 12190 0 -1 2170
box -6 -8 26 248
use FILL  FILL182550x32550
timestamp 0
transform 1 0 12170 0 1 2170
box -6 -8 26 248
use FILL  FILL182550x36150
timestamp 0
transform -1 0 12190 0 -1 2650
box -6 -8 26 248
use FILL  FILL182550x43350
timestamp 0
transform -1 0 12190 0 -1 3130
box -6 -8 26 248
use FILL  FILL182550x46950
timestamp 0
transform 1 0 12170 0 1 3130
box -6 -8 26 248
use FILL  FILL182550x50550
timestamp 0
transform -1 0 12190 0 -1 3610
box -6 -8 26 248
use FILL  FILL182550x57750
timestamp 0
transform -1 0 12190 0 -1 4090
box -6 -8 26 248
use FILL  FILL182550x61350
timestamp 0
transform 1 0 12170 0 1 4090
box -6 -8 26 248
use FILL  FILL182550x64950
timestamp 0
transform -1 0 12190 0 -1 4570
box -6 -8 26 248
use FILL  FILL182550x68550
timestamp 0
transform 1 0 12170 0 1 4570
box -6 -8 26 248
use FILL  FILL182550x72150
timestamp 0
transform -1 0 12190 0 -1 5050
box -6 -8 26 248
use FILL  FILL182550x75750
timestamp 0
transform 1 0 12170 0 1 5050
box -6 -8 26 248
use FILL  FILL182550x79350
timestamp 0
transform -1 0 12190 0 -1 5530
box -6 -8 26 248
use FILL  FILL182550x82950
timestamp 0
transform 1 0 12170 0 1 5530
box -6 -8 26 248
use FILL  FILL182550x86550
timestamp 0
transform -1 0 12190 0 -1 6010
box -6 -8 26 248
use FILL  FILL182550x90150
timestamp 0
transform 1 0 12170 0 1 6010
box -6 -8 26 248
use FILL  FILL182550x93750
timestamp 0
transform -1 0 12190 0 -1 6490
box -6 -8 26 248
use FILL  FILL182550x100950
timestamp 0
transform -1 0 12190 0 -1 6970
box -6 -8 26 248
use FILL  FILL182550x104550
timestamp 0
transform 1 0 12170 0 1 6970
box -6 -8 26 248
use FILL  FILL182550x108150
timestamp 0
transform -1 0 12190 0 -1 7450
box -6 -8 26 248
use FILL  FILL182550x111750
timestamp 0
transform 1 0 12170 0 1 7450
box -6 -8 26 248
use FILL  FILL182550x115350
timestamp 0
transform -1 0 12190 0 -1 7930
box -6 -8 26 248
use FILL  FILL182550x118950
timestamp 0
transform 1 0 12170 0 1 7930
box -6 -8 26 248
use FILL  FILL182550x122550
timestamp 0
transform -1 0 12190 0 -1 8410
box -6 -8 26 248
use FILL  FILL182550x126150
timestamp 0
transform 1 0 12170 0 1 8410
box -6 -8 26 248
use FILL  FILL182550x133350
timestamp 0
transform 1 0 12170 0 1 8890
box -6 -8 26 248
use FILL  FILL182550x140550
timestamp 0
transform 1 0 12170 0 1 9370
box -6 -8 26 248
use FILL  FILL182550x144150
timestamp 0
transform -1 0 12190 0 -1 9850
box -6 -8 26 248
use FILL  FILL182550x147750
timestamp 0
transform 1 0 12170 0 1 9850
box -6 -8 26 248
use FILL  FILL182550x151350
timestamp 0
transform -1 0 12190 0 -1 10330
box -6 -8 26 248
use FILL  FILL182550x154950
timestamp 0
transform 1 0 12170 0 1 10330
box -6 -8 26 248
use FILL  FILL182550x158550
timestamp 0
transform -1 0 12190 0 -1 10810
box -6 -8 26 248
use FILL  FILL182550x162150
timestamp 0
transform 1 0 12170 0 1 10810
box -6 -8 26 248
use FILL  FILL182550x165750
timestamp 0
transform -1 0 12190 0 -1 11290
box -6 -8 26 248
use FILL  FILL182550x169350
timestamp 0
transform 1 0 12170 0 1 11290
box -6 -8 26 248
use FILL  FILL182550x176550
timestamp 0
transform 1 0 12170 0 1 11770
box -6 -8 26 248
use FILL  FILL182850x150
timestamp 0
transform -1 0 12210 0 -1 250
box -6 -8 26 248
use FILL  FILL182850x3750
timestamp 0
transform 1 0 12190 0 1 250
box -6 -8 26 248
use FILL  FILL182850x7350
timestamp 0
transform -1 0 12210 0 -1 730
box -6 -8 26 248
use FILL  FILL182850x10950
timestamp 0
transform 1 0 12190 0 1 730
box -6 -8 26 248
use FILL  FILL182850x14550
timestamp 0
transform -1 0 12210 0 -1 1210
box -6 -8 26 248
use FILL  FILL182850x18150
timestamp 0
transform 1 0 12190 0 1 1210
box -6 -8 26 248
use FILL  FILL182850x21750
timestamp 0
transform -1 0 12210 0 -1 1690
box -6 -8 26 248
use FILL  FILL182850x25350
timestamp 0
transform 1 0 12190 0 1 1690
box -6 -8 26 248
use FILL  FILL182850x28950
timestamp 0
transform -1 0 12210 0 -1 2170
box -6 -8 26 248
use FILL  FILL182850x32550
timestamp 0
transform 1 0 12190 0 1 2170
box -6 -8 26 248
use FILL  FILL182850x36150
timestamp 0
transform -1 0 12210 0 -1 2650
box -6 -8 26 248
use FILL  FILL182850x39750
timestamp 0
transform 1 0 12190 0 1 2650
box -6 -8 26 248
use FILL  FILL182850x43350
timestamp 0
transform -1 0 12210 0 -1 3130
box -6 -8 26 248
use FILL  FILL182850x46950
timestamp 0
transform 1 0 12190 0 1 3130
box -6 -8 26 248
use FILL  FILL182850x50550
timestamp 0
transform -1 0 12210 0 -1 3610
box -6 -8 26 248
use FILL  FILL182850x57750
timestamp 0
transform -1 0 12210 0 -1 4090
box -6 -8 26 248
use FILL  FILL182850x61350
timestamp 0
transform 1 0 12190 0 1 4090
box -6 -8 26 248
use FILL  FILL182850x64950
timestamp 0
transform -1 0 12210 0 -1 4570
box -6 -8 26 248
use FILL  FILL182850x68550
timestamp 0
transform 1 0 12190 0 1 4570
box -6 -8 26 248
use FILL  FILL182850x72150
timestamp 0
transform -1 0 12210 0 -1 5050
box -6 -8 26 248
use FILL  FILL182850x75750
timestamp 0
transform 1 0 12190 0 1 5050
box -6 -8 26 248
use FILL  FILL182850x79350
timestamp 0
transform -1 0 12210 0 -1 5530
box -6 -8 26 248
use FILL  FILL182850x82950
timestamp 0
transform 1 0 12190 0 1 5530
box -6 -8 26 248
use FILL  FILL182850x86550
timestamp 0
transform -1 0 12210 0 -1 6010
box -6 -8 26 248
use FILL  FILL182850x90150
timestamp 0
transform 1 0 12190 0 1 6010
box -6 -8 26 248
use FILL  FILL182850x93750
timestamp 0
transform -1 0 12210 0 -1 6490
box -6 -8 26 248
use FILL  FILL182850x100950
timestamp 0
transform -1 0 12210 0 -1 6970
box -6 -8 26 248
use FILL  FILL182850x104550
timestamp 0
transform 1 0 12190 0 1 6970
box -6 -8 26 248
use FILL  FILL182850x108150
timestamp 0
transform -1 0 12210 0 -1 7450
box -6 -8 26 248
use FILL  FILL182850x111750
timestamp 0
transform 1 0 12190 0 1 7450
box -6 -8 26 248
use FILL  FILL182850x115350
timestamp 0
transform -1 0 12210 0 -1 7930
box -6 -8 26 248
use FILL  FILL182850x118950
timestamp 0
transform 1 0 12190 0 1 7930
box -6 -8 26 248
use FILL  FILL182850x122550
timestamp 0
transform -1 0 12210 0 -1 8410
box -6 -8 26 248
use FILL  FILL182850x126150
timestamp 0
transform 1 0 12190 0 1 8410
box -6 -8 26 248
use FILL  FILL182850x129750
timestamp 0
transform -1 0 12210 0 -1 8890
box -6 -8 26 248
use FILL  FILL182850x133350
timestamp 0
transform 1 0 12190 0 1 8890
box -6 -8 26 248
use FILL  FILL182850x140550
timestamp 0
transform 1 0 12190 0 1 9370
box -6 -8 26 248
use FILL  FILL182850x144150
timestamp 0
transform -1 0 12210 0 -1 9850
box -6 -8 26 248
use FILL  FILL182850x147750
timestamp 0
transform 1 0 12190 0 1 9850
box -6 -8 26 248
use FILL  FILL182850x151350
timestamp 0
transform -1 0 12210 0 -1 10330
box -6 -8 26 248
use FILL  FILL182850x154950
timestamp 0
transform 1 0 12190 0 1 10330
box -6 -8 26 248
use FILL  FILL182850x158550
timestamp 0
transform -1 0 12210 0 -1 10810
box -6 -8 26 248
use FILL  FILL182850x162150
timestamp 0
transform 1 0 12190 0 1 10810
box -6 -8 26 248
use FILL  FILL182850x165750
timestamp 0
transform -1 0 12210 0 -1 11290
box -6 -8 26 248
use FILL  FILL182850x169350
timestamp 0
transform 1 0 12190 0 1 11290
box -6 -8 26 248
use FILL  FILL182850x172950
timestamp 0
transform -1 0 12210 0 -1 11770
box -6 -8 26 248
use FILL  FILL182850x176550
timestamp 0
transform 1 0 12190 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__2478_
timestamp 0
transform -1 0 30 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2479_
timestamp 0
transform -1 0 30 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2480_
timestamp 0
transform 1 0 1870 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2481_
timestamp 0
transform 1 0 2690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2482_
timestamp 0
transform -1 0 30 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__2483_
timestamp 0
transform -1 0 510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__2484_
timestamp 0
transform -1 0 2070 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2485_
timestamp 0
transform 1 0 3890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2486_
timestamp 0
transform 1 0 12010 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2487_
timestamp 0
transform -1 0 6590 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2488_
timestamp 0
transform -1 0 6770 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2489_
timestamp 0
transform 1 0 11970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2490_
timestamp 0
transform 1 0 11970 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2491_
timestamp 0
transform 1 0 6390 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2492_
timestamp 0
transform 1 0 11790 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2493_
timestamp 0
transform -1 0 11890 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2494_
timestamp 0
transform -1 0 990 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__2495_
timestamp 0
transform -1 0 1150 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2496_
timestamp 0
transform -1 0 30 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__2497_
timestamp 0
transform -1 0 4370 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2498_
timestamp 0
transform 1 0 4410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2499_
timestamp 0
transform -1 0 3230 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2500_
timestamp 0
transform -1 0 410 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2501_
timestamp 0
transform -1 0 3610 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2502_
timestamp 0
transform -1 0 30 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__2503_
timestamp 0
transform -1 0 30 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2504_
timestamp 0
transform 1 0 4510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2505_
timestamp 0
transform 1 0 5050 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2506_
timestamp 0
transform -1 0 2490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2507_
timestamp 0
transform 1 0 3770 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2508_
timestamp 0
transform 1 0 3390 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2509_
timestamp 0
transform 1 0 4170 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2510_
timestamp 0
transform 1 0 3030 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2511_
timestamp 0
transform -1 0 4890 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2519_
timestamp 0
transform -1 0 5630 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2520_
timestamp 0
transform -1 0 7490 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2521_
timestamp 0
transform -1 0 7690 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2522_
timestamp 0
transform 1 0 7690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2523_
timestamp 0
transform 1 0 9430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2524_
timestamp 0
transform -1 0 7750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2525_
timestamp 0
transform 1 0 7490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2526_
timestamp 0
transform 1 0 8230 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2527_
timestamp 0
transform 1 0 8430 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2528_
timestamp 0
transform -1 0 9570 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2529_
timestamp 0
transform 1 0 8510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2530_
timestamp 0
transform -1 0 8150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2531_
timestamp 0
transform -1 0 8290 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2532_
timestamp 0
transform -1 0 8710 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2533_
timestamp 0
transform 1 0 9450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2534_
timestamp 0
transform 1 0 10010 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__2535_
timestamp 0
transform -1 0 10210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2536_
timestamp 0
transform -1 0 8710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2537_
timestamp 0
transform -1 0 8510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2538_
timestamp 0
transform -1 0 8310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2539_
timestamp 0
transform 1 0 7910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2540_
timestamp 0
transform -1 0 10610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2541_
timestamp 0
transform -1 0 10810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2542_
timestamp 0
transform 1 0 10850 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2543_
timestamp 0
transform -1 0 10550 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2544_
timestamp 0
transform -1 0 5650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2545_
timestamp 0
transform -1 0 5850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2546_
timestamp 0
transform -1 0 6070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2547_
timestamp 0
transform -1 0 5950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2548_
timestamp 0
transform -1 0 6150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2549_
timestamp 0
transform 1 0 5530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2550_
timestamp 0
transform 1 0 5730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2551_
timestamp 0
transform -1 0 6850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2552_
timestamp 0
transform -1 0 7210 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2553_
timestamp 0
transform -1 0 5670 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2554_
timestamp 0
transform -1 0 6310 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2555_
timestamp 0
transform 1 0 6350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2556_
timestamp 0
transform -1 0 6690 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2557_
timestamp 0
transform -1 0 6170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2558_
timestamp 0
transform 1 0 6450 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2559_
timestamp 0
transform 1 0 6830 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2560_
timestamp 0
transform -1 0 5870 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2561_
timestamp 0
transform -1 0 6510 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2562_
timestamp 0
transform 1 0 6690 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2563_
timestamp 0
transform -1 0 6070 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2564_
timestamp 0
transform 1 0 7730 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2565_
timestamp 0
transform 1 0 7950 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2566_
timestamp 0
transform 1 0 7530 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2567_
timestamp 0
transform 1 0 6930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2568_
timestamp 0
transform -1 0 6570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2569_
timestamp 0
transform 1 0 7150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2570_
timestamp 0
transform -1 0 9330 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2571_
timestamp 0
transform -1 0 9230 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2572_
timestamp 0
transform 1 0 9250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2573_
timestamp 0
transform 1 0 9130 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2574_
timestamp 0
transform -1 0 9210 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2575_
timestamp 0
transform -1 0 9030 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2576_
timestamp 0
transform -1 0 8750 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2577_
timestamp 0
transform -1 0 8950 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2578_
timestamp 0
transform 1 0 9510 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2579_
timestamp 0
transform -1 0 9450 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2580_
timestamp 0
transform -1 0 8250 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2581_
timestamp 0
transform 1 0 8210 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2582_
timestamp 0
transform 1 0 8330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2583_
timestamp 0
transform -1 0 9730 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2584_
timestamp 0
transform 1 0 9390 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2585_
timestamp 0
transform -1 0 11130 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2586_
timestamp 0
transform 1 0 8810 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2587_
timestamp 0
transform 1 0 8610 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2588_
timestamp 0
transform -1 0 8430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2589_
timestamp 0
transform 1 0 8470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2590_
timestamp 0
transform 1 0 8210 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2591_
timestamp 0
transform -1 0 8550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2592_
timestamp 0
transform 1 0 7810 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2593_
timestamp 0
transform -1 0 9050 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2594_
timestamp 0
transform -1 0 8950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2595_
timestamp 0
transform -1 0 9210 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2596_
timestamp 0
transform 1 0 10390 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2597_
timestamp 0
transform 1 0 10570 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2598_
timestamp 0
transform -1 0 10410 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2599_
timestamp 0
transform 1 0 10770 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2600_
timestamp 0
transform -1 0 11370 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2601_
timestamp 0
transform 1 0 8230 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2602_
timestamp 0
transform -1 0 8030 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2603_
timestamp 0
transform 1 0 7030 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2604_
timestamp 0
transform 1 0 8190 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2605_
timestamp 0
transform -1 0 8070 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2606_
timestamp 0
transform -1 0 7670 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2607_
timestamp 0
transform -1 0 6530 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2608_
timestamp 0
transform 1 0 6710 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2609_
timestamp 0
transform 1 0 6910 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2610_
timestamp 0
transform -1 0 7850 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2611_
timestamp 0
transform -1 0 10070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2612_
timestamp 0
transform 1 0 9850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2613_
timestamp 0
transform 1 0 10250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2614_
timestamp 0
transform -1 0 10950 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__2615_
timestamp 0
transform -1 0 7130 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2616_
timestamp 0
transform 1 0 8270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2617_
timestamp 0
transform -1 0 7130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2618_
timestamp 0
transform -1 0 6470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2619_
timestamp 0
transform 1 0 6250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2620_
timestamp 0
transform -1 0 7950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2621_
timestamp 0
transform -1 0 8050 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2622_
timestamp 0
transform 1 0 8310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2623_
timestamp 0
transform -1 0 8910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2624_
timestamp 0
transform 1 0 8050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2625_
timestamp 0
transform 1 0 6810 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2626_
timestamp 0
transform -1 0 8270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2627_
timestamp 0
transform 1 0 9870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2628_
timestamp 0
transform 1 0 11490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2629_
timestamp 0
transform 1 0 11390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2630_
timestamp 0
transform 1 0 11670 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2631_
timestamp 0
transform -1 0 11490 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2632_
timestamp 0
transform 1 0 9390 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2633_
timestamp 0
transform -1 0 8490 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2634_
timestamp 0
transform 1 0 8890 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2635_
timestamp 0
transform -1 0 9130 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2636_
timestamp 0
transform -1 0 9910 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2637_
timestamp 0
transform -1 0 8610 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2638_
timestamp 0
transform 1 0 9690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2639_
timestamp 0
transform 1 0 9950 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2640_
timestamp 0
transform 1 0 8070 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2641_
timestamp 0
transform 1 0 7870 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2642_
timestamp 0
transform 1 0 9350 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2643_
timestamp 0
transform 1 0 9350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2644_
timestamp 0
transform 1 0 8370 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2645_
timestamp 0
transform 1 0 7590 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2646_
timestamp 0
transform 1 0 7390 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2647_
timestamp 0
transform 1 0 8170 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2648_
timestamp 0
transform -1 0 8010 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2649_
timestamp 0
transform -1 0 9010 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2650_
timestamp 0
transform 1 0 11070 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2651_
timestamp 0
transform -1 0 9210 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2652_
timestamp 0
transform -1 0 8510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2653_
timestamp 0
transform 1 0 8690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2654_
timestamp 0
transform 1 0 5810 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2655_
timestamp 0
transform -1 0 6030 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2656_
timestamp 0
transform -1 0 6210 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2657_
timestamp 0
transform -1 0 7610 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2658_
timestamp 0
transform 1 0 7370 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2659_
timestamp 0
transform -1 0 7130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2660_
timestamp 0
transform -1 0 7310 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2661_
timestamp 0
transform -1 0 10750 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2662_
timestamp 0
transform 1 0 10930 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2663_
timestamp 0
transform 1 0 9990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2664_
timestamp 0
transform 1 0 10170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2665_
timestamp 0
transform -1 0 6590 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2666_
timestamp 0
transform 1 0 7170 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2667_
timestamp 0
transform -1 0 6970 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2668_
timestamp 0
transform -1 0 6790 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2669_
timestamp 0
transform 1 0 6710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2670_
timestamp 0
transform -1 0 10570 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2671_
timestamp 0
transform 1 0 11630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2672_
timestamp 0
transform 1 0 11670 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2673_
timestamp 0
transform -1 0 11470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2674_
timestamp 0
transform 1 0 11410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2675_
timestamp 0
transform -1 0 10770 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2676_
timestamp 0
transform 1 0 11390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2677_
timestamp 0
transform -1 0 11470 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2678_
timestamp 0
transform -1 0 10090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2679_
timestamp 0
transform 1 0 9690 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2680_
timestamp 0
transform 1 0 9610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2681_
timestamp 0
transform 1 0 9290 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2682_
timestamp 0
transform -1 0 9510 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2683_
timestamp 0
transform -1 0 10170 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2684_
timestamp 0
transform -1 0 10470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2685_
timestamp 0
transform -1 0 10750 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__2686_
timestamp 0
transform 1 0 10650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2687_
timestamp 0
transform -1 0 9770 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2688_
timestamp 0
transform 1 0 9170 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2689_
timestamp 0
transform 1 0 10490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2690_
timestamp 0
transform -1 0 10850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2691_
timestamp 0
transform -1 0 11050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2692_
timestamp 0
transform 1 0 11230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2693_
timestamp 0
transform -1 0 10390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2694_
timestamp 0
transform 1 0 9590 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2695_
timestamp 0
transform -1 0 10510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2696_
timestamp 0
transform 1 0 10270 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2697_
timestamp 0
transform 1 0 9930 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2698_
timestamp 0
transform 1 0 9910 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2699_
timestamp 0
transform 1 0 9030 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2700_
timestamp 0
transform 1 0 8810 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2701_
timestamp 0
transform -1 0 8450 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2702_
timestamp 0
transform 1 0 8810 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2703_
timestamp 0
transform 1 0 10830 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2704_
timestamp 0
transform -1 0 9090 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2705_
timestamp 0
transform -1 0 9650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2706_
timestamp 0
transform -1 0 10050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2707_
timestamp 0
transform -1 0 9570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2708_
timestamp 0
transform 1 0 8870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2709_
timestamp 0
transform 1 0 8990 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2710_
timestamp 0
transform -1 0 8690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2711_
timestamp 0
transform -1 0 10750 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2712_
timestamp 0
transform -1 0 10730 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2713_
timestamp 0
transform 1 0 10770 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2714_
timestamp 0
transform 1 0 10770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2715_
timestamp 0
transform -1 0 11410 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2716_
timestamp 0
transform 1 0 11570 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2717_
timestamp 0
transform -1 0 10690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2718_
timestamp 0
transform 1 0 11030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2719_
timestamp 0
transform 1 0 11750 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2720_
timestamp 0
transform -1 0 10950 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2721_
timestamp 0
transform -1 0 10850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2722_
timestamp 0
transform -1 0 10890 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2723_
timestamp 0
transform 1 0 11330 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2724_
timestamp 0
transform 1 0 11310 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2725_
timestamp 0
transform 1 0 10290 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2726_
timestamp 0
transform -1 0 9670 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2727_
timestamp 0
transform 1 0 9870 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2728_
timestamp 0
transform -1 0 9850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2729_
timestamp 0
transform -1 0 9450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2730_
timestamp 0
transform 1 0 11190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2731_
timestamp 0
transform 1 0 9430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2732_
timestamp 0
transform 1 0 6650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2733_
timestamp 0
transform -1 0 9070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2734_
timestamp 0
transform 1 0 9430 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2735_
timestamp 0
transform 1 0 9450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2736_
timestamp 0
transform -1 0 8870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2737_
timestamp 0
transform -1 0 9250 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2738_
timestamp 0
transform -1 0 10330 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2739_
timestamp 0
transform 1 0 10510 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2740_
timestamp 0
transform 1 0 11130 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2741_
timestamp 0
transform 1 0 11530 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2742_
timestamp 0
transform -1 0 10530 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2743_
timestamp 0
transform -1 0 10370 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2744_
timestamp 0
transform 1 0 10450 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2745_
timestamp 0
transform -1 0 11110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2746_
timestamp 0
transform -1 0 10110 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2747_
timestamp 0
transform 1 0 10910 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2748_
timestamp 0
transform 1 0 9770 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2749_
timestamp 0
transform 1 0 10630 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2750_
timestamp 0
transform 1 0 10970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2751_
timestamp 0
transform -1 0 10090 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2752_
timestamp 0
transform 1 0 5710 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2753_
timestamp 0
transform -1 0 5930 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2754_
timestamp 0
transform -1 0 5990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2755_
timestamp 0
transform -1 0 7350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2756_
timestamp 0
transform -1 0 7470 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2757_
timestamp 0
transform 1 0 8070 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2758_
timestamp 0
transform -1 0 7530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2759_
timestamp 0
transform -1 0 9670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2760_
timestamp 0
transform -1 0 6190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2761_
timestamp 0
transform -1 0 8830 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2762_
timestamp 0
transform -1 0 8810 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2763_
timestamp 0
transform -1 0 6270 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2764_
timestamp 0
transform -1 0 6350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2765_
timestamp 0
transform -1 0 9310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2766_
timestamp 0
transform -1 0 6650 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2767_
timestamp 0
transform 1 0 8870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2768_
timestamp 0
transform -1 0 5950 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2769_
timestamp 0
transform -1 0 6890 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2770_
timestamp 0
transform 1 0 7070 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2771_
timestamp 0
transform 1 0 9990 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2772_
timestamp 0
transform -1 0 7350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2773_
timestamp 0
transform -1 0 7550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2774_
timestamp 0
transform -1 0 5990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2775_
timestamp 0
transform -1 0 7290 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2776_
timestamp 0
transform 1 0 6110 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2777_
timestamp 0
transform -1 0 9830 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2778_
timestamp 0
transform 1 0 7650 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2779_
timestamp 0
transform 1 0 7870 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2780_
timestamp 0
transform 1 0 7930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2781_
timestamp 0
transform -1 0 7750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2782_
timestamp 0
transform 1 0 7610 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2783_
timestamp 0
transform -1 0 8410 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2784_
timestamp 0
transform -1 0 10950 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2785_
timestamp 0
transform 1 0 9470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2786_
timestamp 0
transform -1 0 7730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2787_
timestamp 0
transform -1 0 9170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2788_
timestamp 0
transform -1 0 10150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2789_
timestamp 0
transform 1 0 10330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2790_
timestamp 0
transform 1 0 7930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2791_
timestamp 0
transform 1 0 8130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2792_
timestamp 0
transform -1 0 7590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2793_
timestamp 0
transform -1 0 7810 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2794_
timestamp 0
transform -1 0 7810 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2795_
timestamp 0
transform -1 0 7530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2796_
timestamp 0
transform -1 0 6930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2797_
timestamp 0
transform -1 0 8350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2798_
timestamp 0
transform 1 0 11890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2799_
timestamp 0
transform -1 0 7310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2800_
timestamp 0
transform -1 0 7430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2801_
timestamp 0
transform 1 0 7070 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2802_
timestamp 0
transform 1 0 6730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2803_
timestamp 0
transform -1 0 6950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2804_
timestamp 0
transform -1 0 8450 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2805_
timestamp 0
transform 1 0 6870 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2806_
timestamp 0
transform -1 0 6770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2807_
timestamp 0
transform -1 0 7030 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2808_
timestamp 0
transform 1 0 10110 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2809_
timestamp 0
transform -1 0 10530 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2810_
timestamp 0
transform 1 0 10510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2811_
timestamp 0
transform 1 0 10330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2812_
timestamp 0
transform 1 0 10190 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2813_
timestamp 0
transform -1 0 10030 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2814_
timestamp 0
transform -1 0 10430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2815_
timestamp 0
transform -1 0 10630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2816_
timestamp 0
transform 1 0 10150 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2817_
timestamp 0
transform -1 0 10250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2818_
timestamp 0
transform -1 0 10910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2819_
timestamp 0
transform -1 0 11010 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2820_
timestamp 0
transform -1 0 11210 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2821_
timestamp 0
transform 1 0 10970 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2822_
timestamp 0
transform -1 0 11910 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2823_
timestamp 0
transform 1 0 11090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2824_
timestamp 0
transform 1 0 10590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2825_
timestamp 0
transform 1 0 11110 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2826_
timestamp 0
transform 1 0 11310 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2827_
timestamp 0
transform -1 0 11770 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2828_
timestamp 0
transform -1 0 11890 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2829_
timestamp 0
transform -1 0 11330 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2830_
timestamp 0
transform 1 0 10970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2831_
timestamp 0
transform 1 0 11030 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2832_
timestamp 0
transform -1 0 11270 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2833_
timestamp 0
transform 1 0 11330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2834_
timestamp 0
transform 1 0 11830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2835_
timestamp 0
transform 1 0 12010 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__2836_
timestamp 0
transform 1 0 11630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2837_
timestamp 0
transform 1 0 11830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2838_
timestamp 0
transform 1 0 11950 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2839_
timestamp 0
transform 1 0 11530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2840_
timestamp 0
transform -1 0 11730 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2841_
timestamp 0
transform -1 0 11590 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2842_
timestamp 0
transform -1 0 9770 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2843_
timestamp 0
transform -1 0 9970 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2844_
timestamp 0
transform -1 0 11750 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2845_
timestamp 0
transform 1 0 11930 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2846_
timestamp 0
transform 1 0 11490 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__2847_
timestamp 0
transform 1 0 11910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2848_
timestamp 0
transform -1 0 11550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2849_
timestamp 0
transform -1 0 11650 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2850_
timestamp 0
transform 1 0 11830 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2851_
timestamp 0
transform -1 0 9830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2852_
timestamp 0
transform -1 0 11010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2853_
timestamp 0
transform 1 0 11190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2854_
timestamp 0
transform 1 0 11770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2855_
timestamp 0
transform 1 0 11770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2856_
timestamp 0
transform -1 0 9790 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2857_
timestamp 0
transform -1 0 9850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2858_
timestamp 0
transform -1 0 8010 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2859_
timestamp 0
transform 1 0 9630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2860_
timestamp 0
transform -1 0 9090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2861_
timestamp 0
transform 1 0 9910 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2862_
timestamp 0
transform 1 0 9510 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2863_
timestamp 0
transform 1 0 8730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2864_
timestamp 0
transform -1 0 7730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2865_
timestamp 0
transform -1 0 6390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2866_
timestamp 0
transform -1 0 8810 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2867_
timestamp 0
transform -1 0 9350 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2868_
timestamp 0
transform 1 0 9150 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2869_
timestamp 0
transform -1 0 10510 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2870_
timestamp 0
transform -1 0 9270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2871_
timestamp 0
transform -1 0 8510 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2872_
timestamp 0
transform 1 0 9710 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2873_
timestamp 0
transform 1 0 9750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2874_
timestamp 0
transform 1 0 9550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2875_
timestamp 0
transform -1 0 11150 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__2876_
timestamp 0
transform 1 0 10150 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2877_
timestamp 0
transform -1 0 10690 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2878_
timestamp 0
transform 1 0 9590 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2879_
timestamp 0
transform -1 0 9810 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2880_
timestamp 0
transform -1 0 10130 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2881_
timestamp 0
transform -1 0 5910 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2882_
timestamp 0
transform -1 0 6090 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2883_
timestamp 0
transform -1 0 5450 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2884_
timestamp 0
transform -1 0 5450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2885_
timestamp 0
transform 1 0 5430 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2886_
timestamp 0
transform -1 0 5250 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__2887_
timestamp 0
transform 1 0 5590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2888_
timestamp 0
transform 1 0 6010 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2889_
timestamp 0
transform -1 0 6250 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2890_
timestamp 0
transform -1 0 6630 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2891_
timestamp 0
transform 1 0 8110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2892_
timestamp 0
transform -1 0 7230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2893_
timestamp 0
transform -1 0 5830 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2894_
timestamp 0
transform 1 0 5330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2895_
timestamp 0
transform -1 0 7430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2896_
timestamp 0
transform -1 0 6550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__2897_
timestamp 0
transform 1 0 7290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2898_
timestamp 0
transform 1 0 11710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2899_
timestamp 0
transform -1 0 6490 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2900_
timestamp 0
transform -1 0 6690 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2901_
timestamp 0
transform -1 0 8130 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2902_
timestamp 0
transform 1 0 9590 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2903_
timestamp 0
transform -1 0 11530 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2904_
timestamp 0
transform 1 0 8310 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2905_
timestamp 0
transform -1 0 6890 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2906_
timestamp 0
transform -1 0 7270 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2907_
timestamp 0
transform -1 0 6290 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2908_
timestamp 0
transform 1 0 8410 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2909_
timestamp 0
transform -1 0 10310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2910_
timestamp 0
transform 1 0 10710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2911_
timestamp 0
transform 1 0 10890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2912_
timestamp 0
transform -1 0 10750 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2913_
timestamp 0
transform -1 0 8630 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2914_
timestamp 0
transform -1 0 8510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2915_
timestamp 0
transform -1 0 11190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2916_
timestamp 0
transform -1 0 7930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2917_
timestamp 0
transform -1 0 6950 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2918_
timestamp 0
transform 1 0 6730 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2919_
timestamp 0
transform -1 0 7150 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2920_
timestamp 0
transform 1 0 7110 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2921_
timestamp 0
transform 1 0 6910 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2922_
timestamp 0
transform 1 0 6570 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2923_
timestamp 0
transform -1 0 5790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2924_
timestamp 0
transform 1 0 8830 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2925_
timestamp 0
transform 1 0 10190 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2926_
timestamp 0
transform 1 0 11930 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2927_
timestamp 0
transform 1 0 8650 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2928_
timestamp 0
transform 1 0 7450 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2929_
timestamp 0
transform 1 0 8170 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2930_
timestamp 0
transform -1 0 8390 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2931_
timestamp 0
transform -1 0 8030 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2932_
timestamp 0
transform 1 0 7830 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2933_
timestamp 0
transform 1 0 7870 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2934_
timestamp 0
transform -1 0 10170 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2935_
timestamp 0
transform 1 0 11290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__2936_
timestamp 0
transform -1 0 8150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2937_
timestamp 0
transform 1 0 8630 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2938_
timestamp 0
transform -1 0 11750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2939_
timestamp 0
transform -1 0 11190 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2940_
timestamp 0
transform -1 0 6530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2941_
timestamp 0
transform 1 0 8810 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2942_
timestamp 0
transform 1 0 8890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2943_
timestamp 0
transform 1 0 9650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2944_
timestamp 0
transform 1 0 9830 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__2945_
timestamp 0
transform 1 0 9010 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2946_
timestamp 0
transform -1 0 9110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2947_
timestamp 0
transform -1 0 8670 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2948_
timestamp 0
transform -1 0 8610 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2949_
timestamp 0
transform 1 0 10790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2950_
timestamp 0
transform 1 0 11610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2951_
timestamp 0
transform -1 0 6930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2952_
timestamp 0
transform -1 0 6730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2953_
timestamp 0
transform 1 0 11230 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2954_
timestamp 0
transform -1 0 8910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2955_
timestamp 0
transform -1 0 10050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__2956_
timestamp 0
transform -1 0 11310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2957_
timestamp 0
transform 1 0 9630 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2958_
timestamp 0
transform 1 0 11590 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__2959_
timestamp 0
transform 1 0 5070 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2960_
timestamp 0
transform -1 0 7330 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2961_
timestamp 0
transform -1 0 7930 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2962_
timestamp 0
transform -1 0 7530 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2963_
timestamp 0
transform -1 0 6450 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__2964_
timestamp 0
transform -1 0 7730 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2965_
timestamp 0
transform -1 0 11710 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__2966_
timestamp 0
transform 1 0 8530 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2967_
timestamp 0
transform 1 0 9230 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__2968_
timestamp 0
transform 1 0 10350 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2969_
timestamp 0
transform 1 0 10550 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__2970_
timestamp 0
transform -1 0 11230 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2971_
timestamp 0
transform 1 0 7690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2972_
timestamp 0
transform -1 0 9290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2973_
timestamp 0
transform 1 0 7330 0 1 250
box -6 -8 26 248
use FILL  FILL_0__2974_
timestamp 0
transform -1 0 7270 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2975_
timestamp 0
transform -1 0 9030 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__2976_
timestamp 0
transform 1 0 10010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2977_
timestamp 0
transform 1 0 10410 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2978_
timestamp 0
transform -1 0 11570 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__2979_
timestamp 0
transform -1 0 11810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__2980_
timestamp 0
transform 1 0 7130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2981_
timestamp 0
transform 1 0 6530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__2982_
timestamp 0
transform 1 0 7470 0 1 730
box -6 -8 26 248
use FILL  FILL_0__2983_
timestamp 0
transform 1 0 11850 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__2984_
timestamp 0
transform 1 0 11590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__2985_
timestamp 0
transform -1 0 7090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__2986_
timestamp 0
transform -1 0 7110 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__2987_
timestamp 0
transform 1 0 5770 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__3000_
timestamp 0
transform -1 0 2170 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3001_
timestamp 0
transform 1 0 2310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3002_
timestamp 0
transform 1 0 2110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__3003_
timestamp 0
transform -1 0 3590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__3004_
timestamp 0
transform 1 0 3790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__3005_
timestamp 0
transform -1 0 3430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__3006_
timestamp 0
transform -1 0 4310 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__3007_
timestamp 0
transform -1 0 4110 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__3008_
timestamp 0
transform 1 0 3830 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__3009_
timestamp 0
transform 1 0 3930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3010_
timestamp 0
transform -1 0 3950 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__3011_
timestamp 0
transform 1 0 3750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3012_
timestamp 0
transform 1 0 2690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__3013_
timestamp 0
transform -1 0 2390 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3014_
timestamp 0
transform 1 0 2530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__3015_
timestamp 0
transform -1 0 4510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3016_
timestamp 0
transform 1 0 4430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__3017_
timestamp 0
transform 1 0 4130 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3018_
timestamp 0
transform 1 0 4330 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3019_
timestamp 0
transform -1 0 3950 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3020_
timestamp 0
transform 1 0 1770 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3021_
timestamp 0
transform 1 0 1610 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3022_
timestamp 0
transform -1 0 2010 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3023_
timestamp 0
transform -1 0 2850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3024_
timestamp 0
transform 1 0 4670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3025_
timestamp 0
transform 1 0 4290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3026_
timestamp 0
transform 1 0 3550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3027_
timestamp 0
transform 1 0 3250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__3028_
timestamp 0
transform -1 0 2750 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__3029_
timestamp 0
transform 1 0 3390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3030_
timestamp 0
transform 1 0 4830 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__3031_
timestamp 0
transform 1 0 4670 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__3032_
timestamp 0
transform 1 0 5830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3033_
timestamp 0
transform -1 0 4550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3034_
timestamp 0
transform 1 0 3770 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3035_
timestamp 0
transform -1 0 4530 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__3036_
timestamp 0
transform -1 0 2330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__3037_
timestamp 0
transform -1 0 3270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__3038_
timestamp 0
transform 1 0 2150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__3039_
timestamp 0
transform -1 0 3530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3040_
timestamp 0
transform -1 0 3750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3041_
timestamp 0
transform 1 0 3350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3042_
timestamp 0
transform -1 0 2730 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3043_
timestamp 0
transform -1 0 3770 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__3044_
timestamp 0
transform -1 0 2570 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3045_
timestamp 0
transform -1 0 2870 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__3046_
timestamp 0
transform -1 0 3210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3047_
timestamp 0
transform 1 0 2810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3048_
timestamp 0
transform 1 0 3350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__3049_
timestamp 0
transform -1 0 3650 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__3050_
timestamp 0
transform -1 0 2890 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__3051_
timestamp 0
transform -1 0 2910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__3052_
timestamp 0
transform 1 0 3070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__3053_
timestamp 0
transform -1 0 2950 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3054_
timestamp 0
transform -1 0 2550 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__3055_
timestamp 0
transform -1 0 2370 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__3056_
timestamp 0
transform -1 0 2690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3057_
timestamp 0
transform -1 0 3210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3058_
timestamp 0
transform 1 0 4130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3059_
timestamp 0
transform -1 0 5050 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__3060_
timestamp 0
transform -1 0 5250 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__3061_
timestamp 0
transform -1 0 6010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3062_
timestamp 0
transform -1 0 5070 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__3063_
timestamp 0
transform -1 0 5090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__3064_
timestamp 0
transform -1 0 4930 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3076_
timestamp 0
transform 1 0 1030 0 1 250
box -6 -8 26 248
use FILL  FILL_0__3077_
timestamp 0
transform -1 0 1250 0 1 250
box -6 -8 26 248
use FILL  FILL_0__3078_
timestamp 0
transform 1 0 870 0 1 250
box -6 -8 26 248
use FILL  FILL_0__3079_
timestamp 0
transform 1 0 950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__3080_
timestamp 0
transform -1 0 830 0 1 730
box -6 -8 26 248
use FILL  FILL_0__3081_
timestamp 0
transform 1 0 770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__3082_
timestamp 0
transform 1 0 1350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__3083_
timestamp 0
transform -1 0 1510 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__3084_
timestamp 0
transform 1 0 1430 0 1 250
box -6 -8 26 248
use FILL  FILL_0__3085_
timestamp 0
transform -1 0 1710 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__3086_
timestamp 0
transform -1 0 410 0 1 730
box -6 -8 26 248
use FILL  FILL_0__3087_
timestamp 0
transform -1 0 590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__3088_
timestamp 0
transform 1 0 390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__3089_
timestamp 0
transform -1 0 1370 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__3090_
timestamp 0
transform 1 0 1170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3091_
timestamp 0
transform -1 0 1850 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__3092_
timestamp 0
transform -1 0 630 0 1 730
box -6 -8 26 248
use FILL  FILL_0__3093_
timestamp 0
transform -1 0 30 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__3094_
timestamp 0
transform -1 0 30 0 1 730
box -6 -8 26 248
use FILL  FILL_0__3095_
timestamp 0
transform -1 0 230 0 1 730
box -6 -8 26 248
use FILL  FILL_0__3096_
timestamp 0
transform -1 0 230 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__3097_
timestamp 0
transform 1 0 1990 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__3098_
timestamp 0
transform -1 0 2290 0 1 250
box -6 -8 26 248
use FILL  FILL_0__3099_
timestamp 0
transform 1 0 1850 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__3100_
timestamp 0
transform 1 0 10 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3101_
timestamp 0
transform -1 0 30 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__3102_
timestamp 0
transform -1 0 1210 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__3103_
timestamp 0
transform -1 0 1170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__3104_
timestamp 0
transform -1 0 210 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__3105_
timestamp 0
transform -1 0 1130 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__3106_
timestamp 0
transform -1 0 2290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__3107_
timestamp 0
transform -1 0 1490 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__3108_
timestamp 0
transform -1 0 370 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3109_
timestamp 0
transform -1 0 550 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3110_
timestamp 0
transform 1 0 690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__3111_
timestamp 0
transform -1 0 890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__3112_
timestamp 0
transform -1 0 30 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__3113_
timestamp 0
transform -1 0 30 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3114_
timestamp 0
transform -1 0 4530 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__3115_
timestamp 0
transform -1 0 4590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3116_
timestamp 0
transform 1 0 4450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__3117_
timestamp 0
transform 1 0 490 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__3118_
timestamp 0
transform -1 0 1650 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__3119_
timestamp 0
transform 1 0 830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3120_
timestamp 0
transform 1 0 990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3121_
timestamp 0
transform -1 0 2310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3122_
timestamp 0
transform -1 0 410 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__3123_
timestamp 0
transform 1 0 290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__3124_
timestamp 0
transform 1 0 190 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__3125_
timestamp 0
transform 1 0 2010 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__3126_
timestamp 0
transform -1 0 2230 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__3127_
timestamp 0
transform 1 0 1530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3128_
timestamp 0
transform 1 0 1370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3129_
timestamp 0
transform 1 0 4710 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__3130_
timestamp 0
transform 1 0 4890 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__3131_
timestamp 0
transform 1 0 5110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__3132_
timestamp 0
transform 1 0 4770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3133_
timestamp 0
transform -1 0 4670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__3134_
timestamp 0
transform -1 0 4310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__3135_
timestamp 0
transform 1 0 670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__3136_
timestamp 0
transform -1 0 730 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__3137_
timestamp 0
transform 1 0 330 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__3138_
timestamp 0
transform 1 0 670 0 1 250
box -6 -8 26 248
use FILL  FILL_0__3139_
timestamp 0
transform 1 0 190 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__3140_
timestamp 0
transform -1 0 1490 0 1 730
box -6 -8 26 248
use FILL  FILL_0__3141_
timestamp 0
transform 1 0 1670 0 1 730
box -6 -8 26 248
use FILL  FILL_0__3142_
timestamp 0
transform -1 0 1650 0 1 250
box -6 -8 26 248
use FILL  FILL_0__3143_
timestamp 0
transform 1 0 2350 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__3144_
timestamp 0
transform 1 0 2470 0 1 250
box -6 -8 26 248
use FILL  FILL_0__3145_
timestamp 0
transform 1 0 2190 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__3146_
timestamp 0
transform -1 0 1890 0 1 730
box -6 -8 26 248
use FILL  FILL_0__3147_
timestamp 0
transform 1 0 1990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__3148_
timestamp 0
transform 1 0 1030 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__3149_
timestamp 0
transform -1 0 870 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__3150_
timestamp 0
transform -1 0 230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__3151_
timestamp 0
transform 1 0 10 0 1 250
box -6 -8 26 248
use FILL  FILL_0__3152_
timestamp 0
transform -1 0 2090 0 1 730
box -6 -8 26 248
use FILL  FILL_0__3284_
timestamp 0
transform -1 0 4690 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__3285_
timestamp 0
transform 1 0 4330 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__3286_
timestamp 0
transform -1 0 3370 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3287_
timestamp 0
transform 1 0 3230 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3288_
timestamp 0
transform 1 0 2150 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3289_
timestamp 0
transform 1 0 2350 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3290_
timestamp 0
transform -1 0 2030 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3291_
timestamp 0
transform 1 0 2970 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3292_
timestamp 0
transform 1 0 3170 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3293_
timestamp 0
transform 1 0 5790 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3294_
timestamp 0
transform -1 0 5830 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3295_
timestamp 0
transform 1 0 5870 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3296_
timestamp 0
transform 1 0 6350 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3297_
timestamp 0
transform 1 0 6550 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3298_
timestamp 0
transform 1 0 5250 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3299_
timestamp 0
transform 1 0 5450 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3300_
timestamp 0
transform 1 0 4590 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3301_
timestamp 0
transform 1 0 4790 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3302_
timestamp 0
transform -1 0 3350 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3303_
timestamp 0
transform -1 0 3510 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3304_
timestamp 0
transform -1 0 3390 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3305_
timestamp 0
transform -1 0 3570 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3306_
timestamp 0
transform 1 0 4310 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3307_
timestamp 0
transform 1 0 4410 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3308_
timestamp 0
transform -1 0 1070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3309_
timestamp 0
transform -1 0 990 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__3310_
timestamp 0
transform 1 0 2470 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3311_
timestamp 0
transform -1 0 2690 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3312_
timestamp 0
transform 1 0 3410 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3313_
timestamp 0
transform -1 0 2330 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3314_
timestamp 0
transform -1 0 210 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__3315_
timestamp 0
transform -1 0 410 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__3316_
timestamp 0
transform -1 0 7490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__3317_
timestamp 0
transform 1 0 6110 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3318_
timestamp 0
transform 1 0 2590 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3319_
timestamp 0
transform 1 0 6610 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3320_
timestamp 0
transform 1 0 5390 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3321_
timestamp 0
transform -1 0 6410 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__3322_
timestamp 0
transform -1 0 3770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3323_
timestamp 0
transform -1 0 3610 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3324_
timestamp 0
transform 1 0 5110 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3325_
timestamp 0
transform -1 0 5330 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3326_
timestamp 0
transform -1 0 5190 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__3327_
timestamp 0
transform 1 0 4770 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__3328_
timestamp 0
transform -1 0 5230 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3329_
timestamp 0
transform -1 0 5650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__3330_
timestamp 0
transform 1 0 5510 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3331_
timestamp 0
transform 1 0 4930 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3332_
timestamp 0
transform -1 0 4610 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__3333_
timestamp 0
transform -1 0 5910 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3334_
timestamp 0
transform 1 0 5890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__3335_
timestamp 0
transform -1 0 410 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3336_
timestamp 0
transform -1 0 230 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3337_
timestamp 0
transform -1 0 850 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3338_
timestamp 0
transform -1 0 870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3339_
timestamp 0
transform -1 0 5830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__3340_
timestamp 0
transform 1 0 6010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__3341_
timestamp 0
transform -1 0 5790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3342_
timestamp 0
transform -1 0 5410 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3343_
timestamp 0
transform -1 0 4330 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3344_
timestamp 0
transform -1 0 5450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__3345_
timestamp 0
transform 1 0 5630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__3346_
timestamp 0
transform 1 0 5230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__3347_
timestamp 0
transform 1 0 5050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__3348_
timestamp 0
transform -1 0 30 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3349_
timestamp 0
transform 1 0 210 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3350_
timestamp 0
transform 1 0 7730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__3351_
timestamp 0
transform -1 0 30 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3352_
timestamp 0
transform 1 0 250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3353_
timestamp 0
transform -1 0 1770 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3354_
timestamp 0
transform 1 0 1950 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3355_
timestamp 0
transform -1 0 270 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3356_
timestamp 0
transform -1 0 470 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3357_
timestamp 0
transform -1 0 810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3358_
timestamp 0
transform -1 0 790 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3359_
timestamp 0
transform -1 0 30 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3360_
timestamp 0
transform -1 0 230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__3361_
timestamp 0
transform -1 0 4830 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3362_
timestamp 0
transform -1 0 4950 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3363_
timestamp 0
transform 1 0 5270 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3364_
timestamp 0
transform -1 0 3370 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3365_
timestamp 0
transform 1 0 3290 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3366_
timestamp 0
transform 1 0 2870 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3367_
timestamp 0
transform 1 0 2510 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3368_
timestamp 0
transform 1 0 2310 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3369_
timestamp 0
transform -1 0 4090 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3370_
timestamp 0
transform -1 0 5250 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3371_
timestamp 0
transform -1 0 7010 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3372_
timestamp 0
transform 1 0 5050 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3373_
timestamp 0
transform -1 0 7450 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3374_
timestamp 0
transform -1 0 7230 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3375_
timestamp 0
transform -1 0 4630 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3376_
timestamp 0
transform -1 0 4670 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3377_
timestamp 0
transform 1 0 4850 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3378_
timestamp 0
transform -1 0 4270 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3379_
timestamp 0
transform 1 0 5710 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3380_
timestamp 0
transform -1 0 7770 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3381_
timestamp 0
transform 1 0 6610 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3382_
timestamp 0
transform 1 0 6430 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3383_
timestamp 0
transform -1 0 7030 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3384_
timestamp 0
transform -1 0 6830 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3385_
timestamp 0
transform 1 0 7210 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3386_
timestamp 0
transform -1 0 6470 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3387_
timestamp 0
transform 1 0 6250 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3388_
timestamp 0
transform 1 0 6670 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3389_
timestamp 0
transform -1 0 7070 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3390_
timestamp 0
transform -1 0 9670 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3391_
timestamp 0
transform -1 0 10210 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3392_
timestamp 0
transform -1 0 210 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3393_
timestamp 0
transform 1 0 190 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3394_
timestamp 0
transform -1 0 190 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3395_
timestamp 0
transform -1 0 210 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3396_
timestamp 0
transform -1 0 30 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3397_
timestamp 0
transform -1 0 1190 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3398_
timestamp 0
transform 1 0 970 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3399_
timestamp 0
transform 1 0 930 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3400_
timestamp 0
transform -1 0 570 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3401_
timestamp 0
transform -1 0 30 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3402_
timestamp 0
transform -1 0 790 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3403_
timestamp 0
transform 1 0 1550 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3404_
timestamp 0
transform -1 0 850 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3405_
timestamp 0
transform 1 0 650 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3406_
timestamp 0
transform -1 0 1830 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3407_
timestamp 0
transform -1 0 430 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__3408_
timestamp 0
transform 1 0 210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__3409_
timestamp 0
transform -1 0 30 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__3410_
timestamp 0
transform -1 0 850 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3411_
timestamp 0
transform -1 0 390 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3412_
timestamp 0
transform -1 0 210 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3413_
timestamp 0
transform -1 0 30 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3414_
timestamp 0
transform -1 0 190 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3415_
timestamp 0
transform -1 0 30 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3416_
timestamp 0
transform -1 0 30 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3417_
timestamp 0
transform -1 0 370 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3418_
timestamp 0
transform -1 0 6890 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3419_
timestamp 0
transform 1 0 6190 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3420_
timestamp 0
transform 1 0 5990 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3421_
timestamp 0
transform 1 0 5230 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3422_
timestamp 0
transform 1 0 5090 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3423_
timestamp 0
transform 1 0 7070 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3424_
timestamp 0
transform -1 0 1330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3425_
timestamp 0
transform 1 0 570 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3426_
timestamp 0
transform 1 0 370 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3427_
timestamp 0
transform -1 0 390 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3428_
timestamp 0
transform -1 0 230 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3429_
timestamp 0
transform 1 0 550 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3430_
timestamp 0
transform -1 0 30 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3431_
timestamp 0
transform -1 0 210 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3432_
timestamp 0
transform 1 0 830 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3433_
timestamp 0
transform 1 0 1430 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3434_
timestamp 0
transform -1 0 930 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3435_
timestamp 0
transform -1 0 1050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3436_
timestamp 0
transform 1 0 1230 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3437_
timestamp 0
transform -1 0 1270 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__3438_
timestamp 0
transform -1 0 950 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3439_
timestamp 0
transform -1 0 750 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3440_
timestamp 0
transform -1 0 1070 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__3441_
timestamp 0
transform 1 0 670 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3442_
timestamp 0
transform 1 0 770 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3443_
timestamp 0
transform -1 0 750 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3444_
timestamp 0
transform -1 0 570 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3445_
timestamp 0
transform -1 0 690 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__3446_
timestamp 0
transform -1 0 1350 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3447_
timestamp 0
transform -1 0 1130 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3448_
timestamp 0
transform -1 0 670 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3449_
timestamp 0
transform 1 0 1290 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3450_
timestamp 0
transform 1 0 1470 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3451_
timestamp 0
transform -1 0 2590 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3452_
timestamp 0
transform -1 0 2790 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3453_
timestamp 0
transform -1 0 3010 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3454_
timestamp 0
transform -1 0 1130 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__3455_
timestamp 0
transform -1 0 230 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3456_
timestamp 0
transform -1 0 30 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3457_
timestamp 0
transform -1 0 790 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3458_
timestamp 0
transform 1 0 570 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3459_
timestamp 0
transform -1 0 510 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__3460_
timestamp 0
transform 1 0 410 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3461_
timestamp 0
transform -1 0 1850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3462_
timestamp 0
transform 1 0 1630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3463_
timestamp 0
transform -1 0 1890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__3464_
timestamp 0
transform -1 0 2010 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3465_
timestamp 0
transform -1 0 1590 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3466_
timestamp 0
transform -1 0 1970 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__3467_
timestamp 0
transform -1 0 1830 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3468_
timestamp 0
transform -1 0 2230 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3469_
timestamp 0
transform -1 0 230 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3470_
timestamp 0
transform -1 0 1170 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3471_
timestamp 0
transform -1 0 1150 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3472_
timestamp 0
transform -1 0 1530 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3473_
timestamp 0
transform 1 0 1710 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3474_
timestamp 0
transform -1 0 2010 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3475_
timestamp 0
transform -1 0 1690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3476_
timestamp 0
transform -1 0 1650 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3477_
timestamp 0
transform -1 0 1830 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3478_
timestamp 0
transform 1 0 1910 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3479_
timestamp 0
transform -1 0 1370 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3480_
timestamp 0
transform -1 0 2770 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3481_
timestamp 0
transform -1 0 6010 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3482_
timestamp 0
transform -1 0 5830 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3483_
timestamp 0
transform 1 0 6670 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3484_
timestamp 0
transform -1 0 7430 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__3485_
timestamp 0
transform -1 0 7230 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__3486_
timestamp 0
transform 1 0 5690 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__3487_
timestamp 0
transform -1 0 5710 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3488_
timestamp 0
transform 1 0 2930 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3489_
timestamp 0
transform -1 0 6070 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__3490_
timestamp 0
transform 1 0 1490 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3491_
timestamp 0
transform 1 0 1310 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3492_
timestamp 0
transform 1 0 1870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3493_
timestamp 0
transform -1 0 1710 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3494_
timestamp 0
transform 1 0 7150 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3495_
timestamp 0
transform -1 0 7530 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3496_
timestamp 0
transform -1 0 7730 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3497_
timestamp 0
transform -1 0 8150 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3498_
timestamp 0
transform -1 0 7370 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3499_
timestamp 0
transform 1 0 1110 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__3500_
timestamp 0
transform 1 0 1310 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__3501_
timestamp 0
transform -1 0 3090 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3502_
timestamp 0
transform -1 0 3690 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3503_
timestamp 0
transform -1 0 3190 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3504_
timestamp 0
transform 1 0 2890 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__3505_
timestamp 0
transform 1 0 3090 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__3506_
timestamp 0
transform -1 0 710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__3507_
timestamp 0
transform -1 0 910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__3508_
timestamp 0
transform 1 0 6310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__3509_
timestamp 0
transform -1 0 6550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__3510_
timestamp 0
transform 1 0 6770 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__3511_
timestamp 0
transform -1 0 6590 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__3512_
timestamp 0
transform 1 0 6530 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__3513_
timestamp 0
transform 1 0 6710 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__3514_
timestamp 0
transform -1 0 6450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3515_
timestamp 0
transform 1 0 7110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__3516_
timestamp 0
transform -1 0 1170 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3517_
timestamp 0
transform 1 0 950 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3518_
timestamp 0
transform -1 0 7430 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3519_
timestamp 0
transform -1 0 7250 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3520_
timestamp 0
transform 1 0 5270 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3521_
timestamp 0
transform -1 0 5470 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3522_
timestamp 0
transform -1 0 30 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__3523_
timestamp 0
transform 1 0 190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3524_
timestamp 0
transform -1 0 410 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__3525_
timestamp 0
transform 1 0 1990 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__3526_
timestamp 0
transform 1 0 2170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__3527_
timestamp 0
transform 1 0 6970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__3528_
timestamp 0
transform -1 0 6910 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__3529_
timestamp 0
transform -1 0 30 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3530_
timestamp 0
transform 1 0 10050 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3531_
timestamp 0
transform 1 0 6010 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3532_
timestamp 0
transform 1 0 5630 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3533_
timestamp 0
transform 1 0 11790 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3534_
timestamp 0
transform -1 0 9090 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3535_
timestamp 0
transform 1 0 7590 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3536_
timestamp 0
transform 1 0 5990 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__3537_
timestamp 0
transform 1 0 5530 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3538_
timestamp 0
transform 1 0 5510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3539_
timestamp 0
transform 1 0 6110 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3540_
timestamp 0
transform 1 0 6310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3541_
timestamp 0
transform -1 0 6190 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3542_
timestamp 0
transform -1 0 6010 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3543_
timestamp 0
transform 1 0 5910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3544_
timestamp 0
transform 1 0 5790 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3545_
timestamp 0
transform 1 0 5790 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3546_
timestamp 0
transform -1 0 6170 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__3547_
timestamp 0
transform 1 0 6330 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3548_
timestamp 0
transform 1 0 6430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3549_
timestamp 0
transform 1 0 6630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3550_
timestamp 0
transform 1 0 6490 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3551_
timestamp 0
transform -1 0 6690 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3552_
timestamp 0
transform 1 0 6770 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3553_
timestamp 0
transform -1 0 7210 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__3554_
timestamp 0
transform 1 0 11170 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3555_
timestamp 0
transform 1 0 10830 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3556_
timestamp 0
transform 1 0 10090 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3557_
timestamp 0
transform -1 0 9170 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3558_
timestamp 0
transform -1 0 10670 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3559_
timestamp 0
transform 1 0 11510 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3560_
timestamp 0
transform 1 0 9970 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3561_
timestamp 0
transform 1 0 9950 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3562_
timestamp 0
transform 1 0 9750 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3563_
timestamp 0
transform -1 0 9830 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3564_
timestamp 0
transform -1 0 11770 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3565_
timestamp 0
transform 1 0 11950 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3566_
timestamp 0
transform 1 0 11370 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3567_
timestamp 0
transform 1 0 11010 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3568_
timestamp 0
transform 1 0 11150 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3569_
timestamp 0
transform 1 0 9690 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3570_
timestamp 0
transform 1 0 10590 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3571_
timestamp 0
transform 1 0 9510 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3572_
timestamp 0
transform -1 0 9350 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3573_
timestamp 0
transform 1 0 10950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3574_
timestamp 0
transform -1 0 9290 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3575_
timestamp 0
transform 1 0 8490 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3576_
timestamp 0
transform -1 0 7970 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3577_
timestamp 0
transform -1 0 8950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3578_
timestamp 0
transform -1 0 9030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3579_
timestamp 0
transform -1 0 8150 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3580_
timestamp 0
transform -1 0 8610 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3581_
timestamp 0
transform 1 0 9550 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3582_
timestamp 0
transform 1 0 9350 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3583_
timestamp 0
transform 1 0 8410 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3584_
timestamp 0
transform -1 0 8350 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3585_
timestamp 0
transform 1 0 9070 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3586_
timestamp 0
transform -1 0 8910 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3587_
timestamp 0
transform -1 0 9150 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3588_
timestamp 0
transform 1 0 8150 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3589_
timestamp 0
transform -1 0 8970 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3590_
timestamp 0
transform -1 0 10550 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3591_
timestamp 0
transform -1 0 10710 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3592_
timestamp 0
transform 1 0 8170 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3593_
timestamp 0
transform -1 0 6150 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3594_
timestamp 0
transform -1 0 10310 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3595_
timestamp 0
transform -1 0 10470 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3596_
timestamp 0
transform 1 0 6910 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3597_
timestamp 0
transform 1 0 6570 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3598_
timestamp 0
transform 1 0 11790 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3599_
timestamp 0
transform -1 0 8850 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3600_
timestamp 0
transform 1 0 8630 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3601_
timestamp 0
transform 1 0 8770 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3602_
timestamp 0
transform -1 0 9890 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3603_
timestamp 0
transform -1 0 10210 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3604_
timestamp 0
transform -1 0 8370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3605_
timestamp 0
transform -1 0 7810 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3606_
timestamp 0
transform -1 0 7950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3607_
timestamp 0
transform 1 0 7750 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3608_
timestamp 0
transform 1 0 11350 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3609_
timestamp 0
transform 1 0 11570 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3610_
timestamp 0
transform 1 0 11430 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3611_
timestamp 0
transform 1 0 11230 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3612_
timestamp 0
transform 1 0 11590 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3613_
timestamp 0
transform 1 0 11330 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3614_
timestamp 0
transform 1 0 11530 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3615_
timestamp 0
transform 1 0 11270 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3616_
timestamp 0
transform -1 0 8050 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3617_
timestamp 0
transform 1 0 11970 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3618_
timestamp 0
transform 1 0 11910 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3619_
timestamp 0
transform -1 0 11490 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3620_
timestamp 0
transform 1 0 8730 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3621_
timestamp 0
transform 1 0 8110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3622_
timestamp 0
transform 1 0 8070 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3623_
timestamp 0
transform 1 0 11070 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3624_
timestamp 0
transform -1 0 11050 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3625_
timestamp 0
transform 1 0 10730 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3626_
timestamp 0
transform 1 0 10930 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3627_
timestamp 0
transform 1 0 10870 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3628_
timestamp 0
transform 1 0 7910 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3629_
timestamp 0
transform 1 0 7570 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3630_
timestamp 0
transform 1 0 7550 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3631_
timestamp 0
transform -1 0 7410 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3632_
timestamp 0
transform 1 0 6970 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3633_
timestamp 0
transform 1 0 7970 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3634_
timestamp 0
transform 1 0 8650 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3635_
timestamp 0
transform 1 0 8310 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3636_
timestamp 0
transform -1 0 6790 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3637_
timestamp 0
transform 1 0 8670 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3638_
timestamp 0
transform 1 0 10770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3639_
timestamp 0
transform 1 0 8530 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3640_
timestamp 0
transform 1 0 9390 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3641_
timestamp 0
transform 1 0 8890 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3642_
timestamp 0
transform -1 0 7250 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3643_
timestamp 0
transform 1 0 7050 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3644_
timestamp 0
transform -1 0 9270 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3645_
timestamp 0
transform -1 0 10350 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3646_
timestamp 0
transform 1 0 9050 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3647_
timestamp 0
transform 1 0 10490 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3648_
timestamp 0
transform 1 0 10810 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3649_
timestamp 0
transform 1 0 10910 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3650_
timestamp 0
transform -1 0 11330 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3651_
timestamp 0
transform 1 0 6710 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3652_
timestamp 0
transform 1 0 4770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3653_
timestamp 0
transform 1 0 4570 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3654_
timestamp 0
transform 1 0 4370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3655_
timestamp 0
transform 1 0 4170 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3656_
timestamp 0
transform 1 0 5370 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3657_
timestamp 0
transform 1 0 5330 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3658_
timestamp 0
transform 1 0 5170 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3659_
timestamp 0
transform 1 0 4590 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3660_
timestamp 0
transform 1 0 4390 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3661_
timestamp 0
transform 1 0 4770 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3662_
timestamp 0
transform 1 0 6510 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3663_
timestamp 0
transform 1 0 6310 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3664_
timestamp 0
transform 1 0 5550 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3665_
timestamp 0
transform 1 0 5150 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3666_
timestamp 0
transform 1 0 5750 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3667_
timestamp 0
transform -1 0 3630 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3668_
timestamp 0
transform 1 0 3850 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3669_
timestamp 0
transform -1 0 3350 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3670_
timestamp 0
transform -1 0 3470 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3671_
timestamp 0
transform 1 0 4110 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3672_
timestamp 0
transform 1 0 4170 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3673_
timestamp 0
transform 1 0 5930 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3674_
timestamp 0
transform -1 0 10670 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3675_
timestamp 0
transform -1 0 10490 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3676_
timestamp 0
transform 1 0 4090 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3677_
timestamp 0
transform -1 0 4150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3678_
timestamp 0
transform 1 0 4590 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3679_
timestamp 0
transform -1 0 4810 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3680_
timestamp 0
transform -1 0 5010 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3681_
timestamp 0
transform -1 0 4710 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3682_
timestamp 0
transform 1 0 1590 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__3683_
timestamp 0
transform 1 0 6210 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3684_
timestamp 0
transform 1 0 6550 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3685_
timestamp 0
transform 1 0 6830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3686_
timestamp 0
transform 1 0 6610 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3687_
timestamp 0
transform 1 0 4830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3688_
timestamp 0
transform -1 0 4850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3689_
timestamp 0
transform 1 0 5030 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3690_
timestamp 0
transform -1 0 4690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3691_
timestamp 0
transform -1 0 4630 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3692_
timestamp 0
transform 1 0 4430 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3693_
timestamp 0
transform 1 0 4810 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3694_
timestamp 0
transform -1 0 6010 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3695_
timestamp 0
transform 1 0 1650 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3696_
timestamp 0
transform 1 0 7530 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3697_
timestamp 0
transform 1 0 7730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3698_
timestamp 0
transform 1 0 6630 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3699_
timestamp 0
transform 1 0 6830 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3700_
timestamp 0
transform -1 0 7030 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3701_
timestamp 0
transform 1 0 4590 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__3702_
timestamp 0
transform 1 0 4290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3703_
timestamp 0
transform 1 0 4350 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3704_
timestamp 0
transform 1 0 4770 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3705_
timestamp 0
transform -1 0 4850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3706_
timestamp 0
transform -1 0 4630 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__3707_
timestamp 0
transform -1 0 4970 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3708_
timestamp 0
transform 1 0 4550 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3709_
timestamp 0
transform 1 0 2410 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3710_
timestamp 0
transform 1 0 9730 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3711_
timestamp 0
transform 1 0 9610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3712_
timestamp 0
transform 1 0 9590 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3713_
timestamp 0
transform 1 0 9970 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3714_
timestamp 0
transform 1 0 8670 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3715_
timestamp 0
transform -1 0 8870 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3716_
timestamp 0
transform -1 0 9470 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3717_
timestamp 0
transform -1 0 10370 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3718_
timestamp 0
transform 1 0 10530 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3719_
timestamp 0
transform -1 0 9070 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3720_
timestamp 0
transform 1 0 9250 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3721_
timestamp 0
transform -1 0 10590 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3722_
timestamp 0
transform -1 0 10410 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3723_
timestamp 0
transform 1 0 10730 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3724_
timestamp 0
transform 1 0 9410 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3725_
timestamp 0
transform 1 0 8270 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3726_
timestamp 0
transform -1 0 8150 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3727_
timestamp 0
transform 1 0 9590 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3728_
timestamp 0
transform -1 0 10150 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3729_
timestamp 0
transform 1 0 9990 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3730_
timestamp 0
transform 1 0 9950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3731_
timestamp 0
transform 1 0 8390 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3732_
timestamp 0
transform 1 0 8770 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3733_
timestamp 0
transform -1 0 3830 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3734_
timestamp 0
transform -1 0 4010 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3735_
timestamp 0
transform 1 0 7590 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3736_
timestamp 0
transform -1 0 7190 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3737_
timestamp 0
transform -1 0 5750 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3738_
timestamp 0
transform 1 0 9530 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3739_
timestamp 0
transform 1 0 9330 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3740_
timestamp 0
transform 1 0 9210 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3741_
timestamp 0
transform -1 0 10710 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3742_
timestamp 0
transform 1 0 11210 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3743_
timestamp 0
transform 1 0 11390 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3744_
timestamp 0
transform 1 0 11130 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3745_
timestamp 0
transform -1 0 10550 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3746_
timestamp 0
transform -1 0 10210 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3747_
timestamp 0
transform -1 0 10150 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3748_
timestamp 0
transform -1 0 10890 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3749_
timestamp 0
transform -1 0 11210 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3750_
timestamp 0
transform 1 0 11010 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3751_
timestamp 0
transform -1 0 8010 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3752_
timestamp 0
transform -1 0 6810 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3753_
timestamp 0
transform -1 0 6710 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3754_
timestamp 0
transform 1 0 4350 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3755_
timestamp 0
transform 1 0 2990 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3756_
timestamp 0
transform 1 0 4030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3757_
timestamp 0
transform 1 0 4510 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3758_
timestamp 0
transform -1 0 5030 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__3759_
timestamp 0
transform -1 0 4810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__3760_
timestamp 0
transform -1 0 4250 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3761_
timestamp 0
transform -1 0 4270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__3762_
timestamp 0
transform -1 0 4370 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__3763_
timestamp 0
transform -1 0 4110 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3764_
timestamp 0
transform -1 0 3390 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3765_
timestamp 0
transform -1 0 4570 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__3766_
timestamp 0
transform 1 0 2190 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3767_
timestamp 0
transform -1 0 2410 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3768_
timestamp 0
transform -1 0 2570 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3769_
timestamp 0
transform -1 0 2770 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3770_
timestamp 0
transform -1 0 3770 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3771_
timestamp 0
transform 1 0 3350 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3772_
timestamp 0
transform -1 0 990 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3773_
timestamp 0
transform 1 0 5770 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__3774_
timestamp 0
transform 1 0 4990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__3775_
timestamp 0
transform -1 0 4950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3776_
timestamp 0
transform -1 0 4790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3777_
timestamp 0
transform 1 0 4850 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3778_
timestamp 0
transform 1 0 4690 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3779_
timestamp 0
transform 1 0 4490 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3780_
timestamp 0
transform 1 0 5170 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3781_
timestamp 0
transform -1 0 5350 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3782_
timestamp 0
transform -1 0 4330 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3783_
timestamp 0
transform 1 0 3770 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3784_
timestamp 0
transform -1 0 5210 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3785_
timestamp 0
transform 1 0 7490 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__3786_
timestamp 0
transform 1 0 7350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__3787_
timestamp 0
transform -1 0 7330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3788_
timestamp 0
transform -1 0 7170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3789_
timestamp 0
transform -1 0 7190 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3790_
timestamp 0
transform -1 0 6170 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3791_
timestamp 0
transform -1 0 6550 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3792_
timestamp 0
transform 1 0 6970 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3793_
timestamp 0
transform -1 0 6770 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3794_
timestamp 0
transform 1 0 7930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__3795_
timestamp 0
transform -1 0 9550 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3796_
timestamp 0
transform 1 0 8250 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3797_
timestamp 0
transform 1 0 7630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3798_
timestamp 0
transform 1 0 6910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3799_
timestamp 0
transform -1 0 7090 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3800_
timestamp 0
transform -1 0 7270 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3801_
timestamp 0
transform 1 0 5610 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3802_
timestamp 0
transform -1 0 5870 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3803_
timestamp 0
transform 1 0 5650 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3804_
timestamp 0
transform 1 0 5270 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3805_
timestamp 0
transform 1 0 5310 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3806_
timestamp 0
transform 1 0 4990 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3807_
timestamp 0
transform -1 0 5470 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3808_
timestamp 0
transform -1 0 7850 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3809_
timestamp 0
transform -1 0 7970 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3810_
timestamp 0
transform 1 0 7770 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3811_
timestamp 0
transform -1 0 7450 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3812_
timestamp 0
transform 1 0 10390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3813_
timestamp 0
transform -1 0 9810 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3814_
timestamp 0
transform 1 0 9790 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3815_
timestamp 0
transform -1 0 9790 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3816_
timestamp 0
transform -1 0 9630 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3817_
timestamp 0
transform 1 0 9090 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3818_
timestamp 0
transform -1 0 8910 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3819_
timestamp 0
transform 1 0 10090 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3820_
timestamp 0
transform 1 0 10170 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3821_
timestamp 0
transform 1 0 6490 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3822_
timestamp 0
transform -1 0 3290 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3823_
timestamp 0
transform -1 0 8210 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3824_
timestamp 0
transform 1 0 7230 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3825_
timestamp 0
transform -1 0 9930 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3826_
timestamp 0
transform 1 0 9410 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3827_
timestamp 0
transform -1 0 9250 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3828_
timestamp 0
transform 1 0 9050 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3829_
timestamp 0
transform 1 0 8850 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3830_
timestamp 0
transform 1 0 7350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3831_
timestamp 0
transform 1 0 7630 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3832_
timestamp 0
transform 1 0 8490 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3833_
timestamp 0
transform 1 0 8670 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3834_
timestamp 0
transform -1 0 8650 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3835_
timestamp 0
transform 1 0 8850 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3836_
timestamp 0
transform 1 0 9150 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3837_
timestamp 0
transform -1 0 8410 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3838_
timestamp 0
transform 1 0 8590 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3839_
timestamp 0
transform 1 0 8830 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3840_
timestamp 0
transform -1 0 8470 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3841_
timestamp 0
transform -1 0 8270 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3842_
timestamp 0
transform 1 0 9030 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3843_
timestamp 0
transform -1 0 8290 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3844_
timestamp 0
transform 1 0 7590 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3845_
timestamp 0
transform 1 0 9250 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__3846_
timestamp 0
transform 1 0 8810 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3847_
timestamp 0
transform 1 0 8090 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3848_
timestamp 0
transform -1 0 7950 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__3849_
timestamp 0
transform 1 0 7730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__3850_
timestamp 0
transform 1 0 7910 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3851_
timestamp 0
transform 1 0 7570 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3852_
timestamp 0
transform -1 0 7770 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3853_
timestamp 0
transform -1 0 7530 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3854_
timestamp 0
transform -1 0 7390 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3855_
timestamp 0
transform 1 0 7770 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__3856_
timestamp 0
transform -1 0 7170 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3857_
timestamp 0
transform -1 0 8270 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3858_
timestamp 0
transform 1 0 8610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3859_
timestamp 0
transform 1 0 7790 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3860_
timestamp 0
transform 1 0 4730 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3861_
timestamp 0
transform 1 0 8470 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3862_
timestamp 0
transform -1 0 8710 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3863_
timestamp 0
transform -1 0 10170 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3864_
timestamp 0
transform 1 0 9410 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3865_
timestamp 0
transform 1 0 7990 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3866_
timestamp 0
transform 1 0 5590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3867_
timestamp 0
transform -1 0 7430 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3868_
timestamp 0
transform -1 0 8490 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3869_
timestamp 0
transform 1 0 7910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3870_
timestamp 0
transform -1 0 7790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3871_
timestamp 0
transform 1 0 6330 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3872_
timestamp 0
transform 1 0 5630 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3873_
timestamp 0
transform -1 0 9470 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3874_
timestamp 0
transform 1 0 9810 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__3875_
timestamp 0
transform 1 0 6850 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3876_
timestamp 0
transform 1 0 4950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3877_
timestamp 0
transform -1 0 4590 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3878_
timestamp 0
transform 1 0 4750 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3879_
timestamp 0
transform 1 0 4510 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3880_
timestamp 0
transform 1 0 5070 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3881_
timestamp 0
transform -1 0 5290 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3882_
timestamp 0
transform -1 0 4310 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3883_
timestamp 0
transform -1 0 4930 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3884_
timestamp 0
transform -1 0 4750 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3885_
timestamp 0
transform 1 0 5110 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3886_
timestamp 0
transform 1 0 9610 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__3887_
timestamp 0
transform 1 0 10330 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__3888_
timestamp 0
transform 1 0 10290 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__3889_
timestamp 0
transform -1 0 10790 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__3890_
timestamp 0
transform -1 0 10710 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3891_
timestamp 0
transform 1 0 10870 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3892_
timestamp 0
transform -1 0 8730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__3893_
timestamp 0
transform -1 0 8530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__3894_
timestamp 0
transform -1 0 11230 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3895_
timestamp 0
transform 1 0 11010 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3896_
timestamp 0
transform 1 0 11770 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3897_
timestamp 0
transform 1 0 11030 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__3898_
timestamp 0
transform 1 0 8210 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3899_
timestamp 0
transform -1 0 5570 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3900_
timestamp 0
transform 1 0 4030 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3901_
timestamp 0
transform -1 0 4990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__3902_
timestamp 0
transform 1 0 4910 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3903_
timestamp 0
transform 1 0 7390 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3904_
timestamp 0
transform -1 0 6970 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3905_
timestamp 0
transform -1 0 6410 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3906_
timestamp 0
transform 1 0 4990 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3907_
timestamp 0
transform -1 0 8150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__3908_
timestamp 0
transform -1 0 6750 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3909_
timestamp 0
transform -1 0 5930 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__3910_
timestamp 0
transform 1 0 5810 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__3911_
timestamp 0
transform -1 0 4490 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3912_
timestamp 0
transform 1 0 4290 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__3913_
timestamp 0
transform -1 0 4510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3914_
timestamp 0
transform 1 0 4170 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__3915_
timestamp 0
transform 1 0 4710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3916_
timestamp 0
transform 1 0 4910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3917_
timestamp 0
transform 1 0 5290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3918_
timestamp 0
transform -1 0 4610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3919_
timestamp 0
transform 1 0 4710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__3920_
timestamp 0
transform 1 0 4430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3921_
timestamp 0
transform 1 0 750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3922_
timestamp 0
transform 1 0 850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3923_
timestamp 0
transform 1 0 370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3924_
timestamp 0
transform 1 0 730 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__3925_
timestamp 0
transform 1 0 5030 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3926_
timestamp 0
transform 1 0 5230 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3927_
timestamp 0
transform -1 0 4650 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3928_
timestamp 0
transform 1 0 5410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3929_
timestamp 0
transform -1 0 4530 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__3930_
timestamp 0
transform 1 0 3370 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__3931_
timestamp 0
transform 1 0 3410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__3932_
timestamp 0
transform 1 0 2270 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__3933_
timestamp 0
transform 1 0 3170 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__3934_
timestamp 0
transform -1 0 4410 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__3935_
timestamp 0
transform 1 0 3770 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3936_
timestamp 0
transform 1 0 3570 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__3937_
timestamp 0
transform 1 0 4150 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__3938_
timestamp 0
transform -1 0 3430 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__3939_
timestamp 0
transform 1 0 3530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__3940_
timestamp 0
transform -1 0 4670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__3941_
timestamp 0
transform 1 0 6870 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3942_
timestamp 0
transform -1 0 9950 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3943_
timestamp 0
transform -1 0 9930 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__3944_
timestamp 0
transform -1 0 9630 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__3945_
timestamp 0
transform -1 0 10150 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3946_
timestamp 0
transform 1 0 9730 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__3947_
timestamp 0
transform 1 0 10330 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3948_
timestamp 0
transform 1 0 10510 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3949_
timestamp 0
transform 1 0 7630 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__3950_
timestamp 0
transform -1 0 6910 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3951_
timestamp 0
transform 1 0 6510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3952_
timestamp 0
transform -1 0 5730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__3953_
timestamp 0
transform 1 0 5390 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3954_
timestamp 0
transform -1 0 5790 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3955_
timestamp 0
transform 1 0 5850 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3956_
timestamp 0
transform -1 0 6070 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3957_
timestamp 0
transform 1 0 6090 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3958_
timestamp 0
transform 1 0 6290 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3959_
timestamp 0
transform 1 0 6410 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3960_
timestamp 0
transform 1 0 2330 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3961_
timestamp 0
transform -1 0 2730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3962_
timestamp 0
transform 1 0 2870 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3963_
timestamp 0
transform 1 0 3470 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3964_
timestamp 0
transform -1 0 4050 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3965_
timestamp 0
transform -1 0 3290 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3966_
timestamp 0
transform -1 0 4250 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3967_
timestamp 0
transform -1 0 5050 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3968_
timestamp 0
transform -1 0 5250 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3969_
timestamp 0
transform -1 0 4250 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3970_
timestamp 0
transform 1 0 3870 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3971_
timestamp 0
transform 1 0 5570 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__3972_
timestamp 0
transform 1 0 5390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__3973_
timestamp 0
transform 1 0 5390 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3974_
timestamp 0
transform -1 0 5610 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3975_
timestamp 0
transform -1 0 5610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3976_
timestamp 0
transform -1 0 5610 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3977_
timestamp 0
transform 1 0 5490 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__3978_
timestamp 0
transform 1 0 6310 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3979_
timestamp 0
transform -1 0 2670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3980_
timestamp 0
transform 1 0 1970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__3981_
timestamp 0
transform 1 0 1810 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__3982_
timestamp 0
transform 1 0 1750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__3983_
timestamp 0
transform -1 0 1890 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__3984_
timestamp 0
transform 1 0 8210 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__3985_
timestamp 0
transform 1 0 6790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3986_
timestamp 0
transform -1 0 7290 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__3987_
timestamp 0
transform 1 0 7570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3988_
timestamp 0
transform 1 0 7490 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3989_
timestamp 0
transform 1 0 7290 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3990_
timestamp 0
transform 1 0 7090 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3991_
timestamp 0
transform -1 0 7250 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__3992_
timestamp 0
transform -1 0 7910 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3993_
timestamp 0
transform 1 0 7670 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3994_
timestamp 0
transform -1 0 7010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__3995_
timestamp 0
transform -1 0 9370 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3996_
timestamp 0
transform -1 0 5970 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__3997_
timestamp 0
transform 1 0 5930 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__3998_
timestamp 0
transform -1 0 6010 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__3999_
timestamp 0
transform 1 0 5790 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4000_
timestamp 0
transform -1 0 5210 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4001_
timestamp 0
transform -1 0 5050 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4002_
timestamp 0
transform -1 0 6910 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4003_
timestamp 0
transform -1 0 6550 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4004_
timestamp 0
transform 1 0 2590 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4005_
timestamp 0
transform 1 0 2790 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4006_
timestamp 0
transform -1 0 2610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4007_
timestamp 0
transform 1 0 2390 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4008_
timestamp 0
transform -1 0 7070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4009_
timestamp 0
transform 1 0 6850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4010_
timestamp 0
transform -1 0 6710 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4011_
timestamp 0
transform 1 0 8590 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4012_
timestamp 0
transform 1 0 6690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4013_
timestamp 0
transform 1 0 6570 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4014_
timestamp 0
transform 1 0 6110 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4015_
timestamp 0
transform 1 0 6470 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4016_
timestamp 0
transform 1 0 9290 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4017_
timestamp 0
transform -1 0 9610 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4018_
timestamp 0
transform -1 0 9790 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4019_
timestamp 0
transform 1 0 9950 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4020_
timestamp 0
transform -1 0 7430 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4021_
timestamp 0
transform -1 0 9990 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4022_
timestamp 0
transform -1 0 6770 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4023_
timestamp 0
transform -1 0 7110 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4024_
timestamp 0
transform 1 0 8910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4025_
timestamp 0
transform -1 0 7630 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4026_
timestamp 0
transform -1 0 7790 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4027_
timestamp 0
transform 1 0 8330 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4028_
timestamp 0
transform 1 0 7870 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4029_
timestamp 0
transform 1 0 10970 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4030_
timestamp 0
transform 1 0 10790 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4031_
timestamp 0
transform 1 0 9170 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4032_
timestamp 0
transform 1 0 8610 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4033_
timestamp 0
transform -1 0 9270 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4034_
timestamp 0
transform 1 0 3930 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4035_
timestamp 0
transform 1 0 9730 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4036_
timestamp 0
transform -1 0 9590 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4037_
timestamp 0
transform -1 0 9110 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4038_
timestamp 0
transform -1 0 8070 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4039_
timestamp 0
transform -1 0 7010 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4040_
timestamp 0
transform 1 0 11950 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4041_
timestamp 0
transform 1 0 9230 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4042_
timestamp 0
transform -1 0 5950 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__4043_
timestamp 0
transform 1 0 5270 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4044_
timestamp 0
transform -1 0 5350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4045_
timestamp 0
transform -1 0 5410 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4046_
timestamp 0
transform -1 0 5770 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4047_
timestamp 0
transform -1 0 5950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4048_
timestamp 0
transform -1 0 5950 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4049_
timestamp 0
transform 1 0 5430 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4050_
timestamp 0
transform -1 0 5210 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4051_
timestamp 0
transform 1 0 5550 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4052_
timestamp 0
transform -1 0 6170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4053_
timestamp 0
transform -1 0 8150 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4054_
timestamp 0
transform 1 0 3670 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4055_
timestamp 0
transform -1 0 3510 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4056_
timestamp 0
transform 1 0 2670 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4057_
timestamp 0
transform 1 0 3290 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4058_
timestamp 0
transform -1 0 7430 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4059_
timestamp 0
transform 1 0 7290 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4060_
timestamp 0
transform -1 0 7970 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4061_
timestamp 0
transform -1 0 8910 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4062_
timestamp 0
transform -1 0 3090 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4063_
timestamp 0
transform 1 0 5010 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4064_
timestamp 0
transform -1 0 4990 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4065_
timestamp 0
transform 1 0 5210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4066_
timestamp 0
transform 1 0 4410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4067_
timestamp 0
transform -1 0 7050 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4068_
timestamp 0
transform 1 0 3070 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4069_
timestamp 0
transform -1 0 610 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__4070_
timestamp 0
transform 1 0 1090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__4071_
timestamp 0
transform 1 0 490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__4072_
timestamp 0
transform -1 0 810 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__4073_
timestamp 0
transform 1 0 4030 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4074_
timestamp 0
transform 1 0 4230 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4075_
timestamp 0
transform 1 0 4150 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4076_
timestamp 0
transform -1 0 5410 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4077_
timestamp 0
transform 1 0 5430 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4078_
timestamp 0
transform -1 0 5450 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4079_
timestamp 0
transform 1 0 3710 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4080_
timestamp 0
transform 1 0 5810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4081_
timestamp 0
transform 1 0 850 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4082_
timestamp 0
transform 1 0 4090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4083_
timestamp 0
transform -1 0 3890 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4084_
timestamp 0
transform 1 0 1590 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4085_
timestamp 0
transform 1 0 1410 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4086_
timestamp 0
transform 1 0 1550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4087_
timestamp 0
transform 1 0 1510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4088_
timestamp 0
transform -1 0 4450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4089_
timestamp 0
transform -1 0 4410 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4090_
timestamp 0
transform -1 0 3910 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4091_
timestamp 0
transform -1 0 3350 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4092_
timestamp 0
transform -1 0 5630 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4093_
timestamp 0
transform 1 0 4570 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4094_
timestamp 0
transform 1 0 4150 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4095_
timestamp 0
transform 1 0 1890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4096_
timestamp 0
transform 1 0 1710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4097_
timestamp 0
transform 1 0 1590 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4098_
timestamp 0
transform 1 0 1510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4099_
timestamp 0
transform 1 0 7090 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4100_
timestamp 0
transform 1 0 7970 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4101_
timestamp 0
transform 1 0 8130 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4102_
timestamp 0
transform -1 0 8330 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4103_
timestamp 0
transform 1 0 7950 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4104_
timestamp 0
transform -1 0 8170 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4105_
timestamp 0
transform 1 0 8610 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4106_
timestamp 0
transform 1 0 6650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4107_
timestamp 0
transform -1 0 1050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0__4108_
timestamp 0
transform -1 0 450 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__4109_
timestamp 0
transform -1 0 1790 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4110_
timestamp 0
transform -1 0 7730 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4111_
timestamp 0
transform -1 0 9470 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4112_
timestamp 0
transform 1 0 2850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__4113_
timestamp 0
transform 1 0 3050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__4114_
timestamp 0
transform 1 0 3550 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4115_
timestamp 0
transform 1 0 4430 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4116_
timestamp 0
transform -1 0 5310 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4117_
timestamp 0
transform 1 0 4850 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4118_
timestamp 0
transform 1 0 4770 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4119_
timestamp 0
transform 1 0 3930 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4120_
timestamp 0
transform -1 0 3670 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4121_
timestamp 0
transform -1 0 4510 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4122_
timestamp 0
transform 1 0 4650 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4123_
timestamp 0
transform 1 0 8010 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4124_
timestamp 0
transform 1 0 8530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4125_
timestamp 0
transform -1 0 4250 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4126_
timestamp 0
transform 1 0 4210 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4127_
timestamp 0
transform 1 0 4030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4128_
timestamp 0
transform 1 0 4450 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4129_
timestamp 0
transform -1 0 4870 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4130_
timestamp 0
transform 1 0 5990 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4131_
timestamp 0
transform 1 0 4270 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4132_
timestamp 0
transform -1 0 4490 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4133_
timestamp 0
transform -1 0 1970 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4134_
timestamp 0
transform 1 0 1750 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4135_
timestamp 0
transform -1 0 2110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4136_
timestamp 0
transform -1 0 2110 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4137_
timestamp 0
transform -1 0 1950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4138_
timestamp 0
transform -1 0 2190 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4139_
timestamp 0
transform 1 0 1970 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4140_
timestamp 0
transform -1 0 2990 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4141_
timestamp 0
transform 1 0 1770 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4142_
timestamp 0
transform 1 0 1570 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4143_
timestamp 0
transform -1 0 1410 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4144_
timestamp 0
transform 1 0 1550 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4145_
timestamp 0
transform -1 0 1030 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4146_
timestamp 0
transform 1 0 3050 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4147_
timestamp 0
transform -1 0 1990 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4148_
timestamp 0
transform -1 0 3170 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4149_
timestamp 0
transform 1 0 3150 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4150_
timestamp 0
transform 1 0 3150 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4151_
timestamp 0
transform 1 0 3690 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4152_
timestamp 0
transform -1 0 3630 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4153_
timestamp 0
transform -1 0 2010 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4154_
timestamp 0
transform -1 0 2210 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4155_
timestamp 0
transform 1 0 590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4156_
timestamp 0
transform 1 0 950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4157_
timestamp 0
transform -1 0 5890 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4158_
timestamp 0
transform 1 0 6050 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4159_
timestamp 0
transform 1 0 6250 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4160_
timestamp 0
transform 1 0 5330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4161_
timestamp 0
transform -1 0 5550 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4162_
timestamp 0
transform 1 0 5130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4163_
timestamp 0
transform -1 0 5150 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4164_
timestamp 0
transform 1 0 5690 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4165_
timestamp 0
transform -1 0 5690 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4166_
timestamp 0
transform 1 0 5710 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4167_
timestamp 0
transform 1 0 6410 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4168_
timestamp 0
transform -1 0 5850 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4169_
timestamp 0
transform 1 0 5650 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4170_
timestamp 0
transform 1 0 6050 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4171_
timestamp 0
transform 1 0 5470 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4172_
timestamp 0
transform 1 0 5090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4173_
timestamp 0
transform 1 0 3770 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4174_
timestamp 0
transform 1 0 5490 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4175_
timestamp 0
transform 1 0 5110 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4176_
timestamp 0
transform -1 0 3290 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4177_
timestamp 0
transform 1 0 2970 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4178_
timestamp 0
transform -1 0 2190 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4179_
timestamp 0
transform -1 0 2310 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4180_
timestamp 0
transform 1 0 2770 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4181_
timestamp 0
transform -1 0 2390 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4182_
timestamp 0
transform 1 0 2230 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4183_
timestamp 0
transform -1 0 3210 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4184_
timestamp 0
transform 1 0 3370 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4185_
timestamp 0
transform 1 0 2790 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4186_
timestamp 0
transform -1 0 2410 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4187_
timestamp 0
transform 1 0 4030 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4188_
timestamp 0
transform 1 0 4230 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4189_
timestamp 0
transform -1 0 4050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4190_
timestamp 0
transform -1 0 3870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4191_
timestamp 0
transform -1 0 3690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4192_
timestamp 0
transform -1 0 5150 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4193_
timestamp 0
transform -1 0 5010 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4194_
timestamp 0
transform -1 0 3870 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4195_
timestamp 0
transform 1 0 3410 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4196_
timestamp 0
transform 1 0 3710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4197_
timestamp 0
transform 1 0 1570 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4198_
timestamp 0
transform -1 0 1690 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4199_
timestamp 0
transform -1 0 1890 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4200_
timestamp 0
transform -1 0 2290 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4201_
timestamp 0
transform -1 0 1510 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4202_
timestamp 0
transform -1 0 1390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__4203_
timestamp 0
transform -1 0 1770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__4204_
timestamp 0
transform -1 0 2570 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4205_
timestamp 0
transform 1 0 2570 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4206_
timestamp 0
transform -1 0 8550 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4207_
timestamp 0
transform -1 0 7890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4208_
timestamp 0
transform -1 0 6230 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4209_
timestamp 0
transform -1 0 230 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4210_
timestamp 0
transform 1 0 10 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4211_
timestamp 0
transform -1 0 30 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4212_
timestamp 0
transform -1 0 410 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4213_
timestamp 0
transform 1 0 870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4214_
timestamp 0
transform -1 0 1390 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4215_
timestamp 0
transform 1 0 1370 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4216_
timestamp 0
transform -1 0 1970 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4217_
timestamp 0
transform -1 0 2950 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4218_
timestamp 0
transform -1 0 2170 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4219_
timestamp 0
transform 1 0 2250 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4220_
timestamp 0
transform 1 0 2450 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4221_
timestamp 0
transform -1 0 230 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4222_
timestamp 0
transform -1 0 30 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4223_
timestamp 0
transform -1 0 410 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4224_
timestamp 0
transform -1 0 410 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4225_
timestamp 0
transform -1 0 390 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4226_
timestamp 0
transform 1 0 10 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4227_
timestamp 0
transform -1 0 230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4228_
timestamp 0
transform -1 0 2370 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4229_
timestamp 0
transform 1 0 2570 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4230_
timestamp 0
transform -1 0 2790 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4231_
timestamp 0
transform 1 0 3130 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4232_
timestamp 0
transform -1 0 3590 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4233_
timestamp 0
transform -1 0 2170 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4234_
timestamp 0
transform -1 0 3030 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4235_
timestamp 0
transform -1 0 3790 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4236_
timestamp 0
transform 1 0 3870 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4237_
timestamp 0
transform -1 0 4090 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4238_
timestamp 0
transform 1 0 3410 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4239_
timestamp 0
transform 1 0 2570 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4240_
timestamp 0
transform 1 0 2210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4241_
timestamp 0
transform -1 0 2070 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4242_
timestamp 0
transform 1 0 2250 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4243_
timestamp 0
transform -1 0 4430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4244_
timestamp 0
transform -1 0 5430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4245_
timestamp 0
transform -1 0 6010 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4246_
timestamp 0
transform -1 0 4130 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4247_
timestamp 0
transform 1 0 2530 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4248_
timestamp 0
transform -1 0 5610 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4249_
timestamp 0
transform -1 0 2310 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4250_
timestamp 0
transform -1 0 4230 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4251_
timestamp 0
transform 1 0 5610 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4252_
timestamp 0
transform -1 0 5810 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4253_
timestamp 0
transform -1 0 3710 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4254_
timestamp 0
transform -1 0 2130 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4255_
timestamp 0
transform 1 0 2470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4256_
timestamp 0
transform -1 0 3830 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4257_
timestamp 0
transform 1 0 4010 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4258_
timestamp 0
transform 1 0 4210 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4259_
timestamp 0
transform 1 0 3970 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4260_
timestamp 0
transform -1 0 2930 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4261_
timestamp 0
transform -1 0 3990 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4262_
timestamp 0
transform 1 0 1510 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4263_
timestamp 0
transform -1 0 7930 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4264_
timestamp 0
transform 1 0 7550 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4265_
timestamp 0
transform 1 0 7370 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4266_
timestamp 0
transform 1 0 7050 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4267_
timestamp 0
transform 1 0 7490 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4268_
timestamp 0
transform -1 0 6730 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4269_
timestamp 0
transform -1 0 9410 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4270_
timestamp 0
transform -1 0 11110 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4271_
timestamp 0
transform 1 0 11090 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4272_
timestamp 0
transform 1 0 9190 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4273_
timestamp 0
transform 1 0 8990 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4274_
timestamp 0
transform -1 0 8910 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4275_
timestamp 0
transform 1 0 8730 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4276_
timestamp 0
transform 1 0 8810 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4277_
timestamp 0
transform 1 0 8830 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4278_
timestamp 0
transform 1 0 7710 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4279_
timestamp 0
transform 1 0 10490 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4280_
timestamp 0
transform 1 0 10690 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4281_
timestamp 0
transform -1 0 10650 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4282_
timestamp 0
transform -1 0 1190 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4283_
timestamp 0
transform -1 0 7030 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4284_
timestamp 0
transform 1 0 7610 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4285_
timestamp 0
transform 1 0 7350 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4286_
timestamp 0
transform -1 0 1030 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4287_
timestamp 0
transform -1 0 1230 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4288_
timestamp 0
transform -1 0 1630 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4289_
timestamp 0
transform -1 0 4330 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4290_
timestamp 0
transform 1 0 6810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4291_
timestamp 0
transform 1 0 6830 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4292_
timestamp 0
transform -1 0 2490 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4293_
timestamp 0
transform -1 0 1770 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4294_
timestamp 0
transform -1 0 7250 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4295_
timestamp 0
transform 1 0 1450 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4296_
timestamp 0
transform -1 0 30 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4297_
timestamp 0
transform 1 0 1110 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4298_
timestamp 0
transform -1 0 3230 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4299_
timestamp 0
transform 1 0 3310 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4300_
timestamp 0
transform -1 0 3790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4301_
timestamp 0
transform -1 0 3510 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4302_
timestamp 0
transform -1 0 3630 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4303_
timestamp 0
transform -1 0 1550 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4304_
timestamp 0
transform 1 0 1130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4305_
timestamp 0
transform -1 0 2250 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4306_
timestamp 0
transform -1 0 2810 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4307_
timestamp 0
transform 1 0 6170 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4308_
timestamp 0
transform -1 0 6250 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4309_
timestamp 0
transform 1 0 2810 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4310_
timestamp 0
transform -1 0 2390 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4311_
timestamp 0
transform 1 0 2290 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4312_
timestamp 0
transform 1 0 870 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4313_
timestamp 0
transform 1 0 1450 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4314_
timestamp 0
transform 1 0 1630 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4315_
timestamp 0
transform -1 0 2670 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4316_
timestamp 0
transform -1 0 2730 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4317_
timestamp 0
transform 1 0 4370 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4318_
timestamp 0
transform 1 0 4050 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4319_
timestamp 0
transform 1 0 3550 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4320_
timestamp 0
transform -1 0 2990 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4321_
timestamp 0
transform 1 0 2770 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4322_
timestamp 0
transform 1 0 1510 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4323_
timestamp 0
transform -1 0 2630 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4324_
timestamp 0
transform -1 0 1770 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4325_
timestamp 0
transform -1 0 4030 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4326_
timestamp 0
transform 1 0 3930 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4327_
timestamp 0
transform 1 0 4070 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4328_
timestamp 0
transform -1 0 8510 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4329_
timestamp 0
transform 1 0 1670 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4330_
timestamp 0
transform 1 0 2070 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4331_
timestamp 0
transform -1 0 1390 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4332_
timestamp 0
transform -1 0 1930 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4333_
timestamp 0
transform -1 0 2850 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4334_
timestamp 0
transform -1 0 3050 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4335_
timestamp 0
transform -1 0 3630 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4336_
timestamp 0
transform 1 0 2790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4337_
timestamp 0
transform 1 0 2590 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4338_
timestamp 0
transform 1 0 2630 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4339_
timestamp 0
transform -1 0 3250 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4340_
timestamp 0
transform -1 0 3430 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4341_
timestamp 0
transform 1 0 3370 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4342_
timestamp 0
transform -1 0 3190 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4343_
timestamp 0
transform 1 0 3430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4344_
timestamp 0
transform 1 0 1730 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4345_
timestamp 0
transform -1 0 2370 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4346_
timestamp 0
transform 1 0 6850 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4347_
timestamp 0
transform -1 0 6670 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4348_
timestamp 0
transform -1 0 570 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4349_
timestamp 0
transform -1 0 990 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4350_
timestamp 0
transform 1 0 2110 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4351_
timestamp 0
transform -1 0 2730 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4352_
timestamp 0
transform 1 0 3710 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4353_
timestamp 0
transform -1 0 6110 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4354_
timestamp 0
transform -1 0 3390 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4355_
timestamp 0
transform -1 0 810 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4356_
timestamp 0
transform -1 0 450 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4357_
timestamp 0
transform 1 0 2310 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4358_
timestamp 0
transform -1 0 5170 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4359_
timestamp 0
transform 1 0 5090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4360_
timestamp 0
transform -1 0 5050 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4361_
timestamp 0
transform 1 0 2990 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4362_
timestamp 0
transform 1 0 4830 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4363_
timestamp 0
transform -1 0 4670 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4364_
timestamp 0
transform 1 0 3630 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4365_
timestamp 0
transform -1 0 5610 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4366_
timestamp 0
transform -1 0 5810 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4367_
timestamp 0
transform -1 0 2850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4368_
timestamp 0
transform 1 0 7490 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4369_
timestamp 0
transform -1 0 7330 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4370_
timestamp 0
transform 1 0 610 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4371_
timestamp 0
transform -1 0 1750 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4372_
timestamp 0
transform 1 0 1870 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4373_
timestamp 0
transform 1 0 2070 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4374_
timestamp 0
transform 1 0 2430 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4375_
timestamp 0
transform -1 0 3750 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4376_
timestamp 0
transform 1 0 7430 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4377_
timestamp 0
transform 1 0 11490 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4378_
timestamp 0
transform -1 0 1210 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4379_
timestamp 0
transform -1 0 5170 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4380_
timestamp 0
transform 1 0 4750 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4381_
timestamp 0
transform 1 0 5850 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4382_
timestamp 0
transform 1 0 190 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4383_
timestamp 0
transform 1 0 10 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4384_
timestamp 0
transform 1 0 6190 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4385_
timestamp 0
transform 1 0 6390 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4386_
timestamp 0
transform 1 0 6790 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4387_
timestamp 0
transform 1 0 6590 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4388_
timestamp 0
transform -1 0 5390 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4389_
timestamp 0
transform -1 0 6490 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4390_
timestamp 0
transform 1 0 6990 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4391_
timestamp 0
transform 1 0 4950 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4392_
timestamp 0
transform -1 0 6290 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4393_
timestamp 0
transform 1 0 6450 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4394_
timestamp 0
transform 1 0 6630 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4395_
timestamp 0
transform 1 0 6750 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4396_
timestamp 0
transform -1 0 6230 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4397_
timestamp 0
transform 1 0 3990 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4398_
timestamp 0
transform 1 0 2970 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4399_
timestamp 0
transform 1 0 2090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4400_
timestamp 0
transform -1 0 6270 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4401_
timestamp 0
transform 1 0 6190 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4402_
timestamp 0
transform -1 0 6030 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4403_
timestamp 0
transform -1 0 5570 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4404_
timestamp 0
transform 1 0 1350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4405_
timestamp 0
transform -1 0 1790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4406_
timestamp 0
transform -1 0 2490 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4407_
timestamp 0
transform -1 0 2290 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4408_
timestamp 0
transform 1 0 1510 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4409_
timestamp 0
transform -1 0 1730 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4410_
timestamp 0
transform 1 0 3530 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4411_
timestamp 0
transform 1 0 3850 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4412_
timestamp 0
transform 1 0 1690 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4413_
timestamp 0
transform -1 0 210 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4414_
timestamp 0
transform 1 0 210 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4415_
timestamp 0
transform 1 0 390 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4416_
timestamp 0
transform 1 0 1470 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__4417_
timestamp 0
transform -1 0 1690 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__4418_
timestamp 0
transform -1 0 2510 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__4419_
timestamp 0
transform 1 0 2070 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__4420_
timestamp 0
transform 1 0 2190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4421_
timestamp 0
transform 1 0 2390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4422_
timestamp 0
transform -1 0 1930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4423_
timestamp 0
transform -1 0 570 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4424_
timestamp 0
transform 1 0 1990 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4425_
timestamp 0
transform 1 0 1030 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4426_
timestamp 0
transform 1 0 1230 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4427_
timestamp 0
transform 1 0 3490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4428_
timestamp 0
transform -1 0 3330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4429_
timestamp 0
transform 1 0 1210 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4430_
timestamp 0
transform 1 0 1410 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4431_
timestamp 0
transform -1 0 690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4432_
timestamp 0
transform -1 0 570 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4433_
timestamp 0
transform -1 0 810 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4434_
timestamp 0
transform -1 0 1270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__4435_
timestamp 0
transform 1 0 1450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__4436_
timestamp 0
transform 1 0 3050 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__4437_
timestamp 0
transform -1 0 3270 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__4438_
timestamp 0
transform -1 0 6510 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4439_
timestamp 0
transform 1 0 5910 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4440_
timestamp 0
transform -1 0 4690 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4441_
timestamp 0
transform 1 0 4090 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4442_
timestamp 0
transform 1 0 3870 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4443_
timestamp 0
transform 1 0 3750 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4444_
timestamp 0
transform 1 0 3570 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4445_
timestamp 0
transform 1 0 3910 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4446_
timestamp 0
transform 1 0 4330 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4447_
timestamp 0
transform 1 0 4510 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4448_
timestamp 0
transform 1 0 2430 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4449_
timestamp 0
transform 1 0 990 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4450_
timestamp 0
transform -1 0 1750 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4451_
timestamp 0
transform 1 0 1350 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4452_
timestamp 0
transform -1 0 2150 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4453_
timestamp 0
transform 1 0 7170 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4454_
timestamp 0
transform -1 0 990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4455_
timestamp 0
transform 1 0 6710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4456_
timestamp 0
transform 1 0 6930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4457_
timestamp 0
transform 1 0 7130 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4458_
timestamp 0
transform -1 0 7330 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4459_
timestamp 0
transform -1 0 6950 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4460_
timestamp 0
transform -1 0 8270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4461_
timestamp 0
transform 1 0 7550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4462_
timestamp 0
transform -1 0 6650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4463_
timestamp 0
transform 1 0 1170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4464_
timestamp 0
transform -1 0 2470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4465_
timestamp 0
transform -1 0 5810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4466_
timestamp 0
transform 1 0 5950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4467_
timestamp 0
transform 1 0 6370 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4468_
timestamp 0
transform 1 0 6610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4469_
timestamp 0
transform 1 0 6810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4470_
timestamp 0
transform -1 0 6570 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4471_
timestamp 0
transform 1 0 7170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4472_
timestamp 0
transform -1 0 6370 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4473_
timestamp 0
transform 1 0 8090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4474_
timestamp 0
transform -1 0 6190 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4475_
timestamp 0
transform 1 0 2650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4476_
timestamp 0
transform -1 0 1150 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4477_
timestamp 0
transform -1 0 2550 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4478_
timestamp 0
transform 1 0 2530 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4479_
timestamp 0
transform 1 0 5250 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4480_
timestamp 0
transform 1 0 1330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4481_
timestamp 0
transform 1 0 170 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4482_
timestamp 0
transform 1 0 370 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4483_
timestamp 0
transform 1 0 3130 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4484_
timestamp 0
transform -1 0 4890 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4485_
timestamp 0
transform 1 0 5270 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4486_
timestamp 0
transform -1 0 5090 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4487_
timestamp 0
transform -1 0 5470 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4488_
timestamp 0
transform 1 0 5630 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4489_
timestamp 0
transform -1 0 5750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4490_
timestamp 0
transform -1 0 5710 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4491_
timestamp 0
transform -1 0 5790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4492_
timestamp 0
transform 1 0 10 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4493_
timestamp 0
transform -1 0 5630 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4494_
timestamp 0
transform 1 0 5430 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4495_
timestamp 0
transform 1 0 4290 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4496_
timestamp 0
transform 1 0 3750 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4497_
timestamp 0
transform -1 0 3530 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4498_
timestamp 0
transform -1 0 4570 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4499_
timestamp 0
transform 1 0 1190 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4500_
timestamp 0
transform 1 0 6290 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4501_
timestamp 0
transform 1 0 6010 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4502_
timestamp 0
transform -1 0 4450 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4503_
timestamp 0
transform 1 0 6410 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4504_
timestamp 0
transform -1 0 1650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__4505_
timestamp 0
transform -1 0 4770 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__4506_
timestamp 0
transform -1 0 5210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4507_
timestamp 0
transform 1 0 5590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__4508_
timestamp 0
transform 1 0 5470 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4509_
timestamp 0
transform -1 0 5690 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4510_
timestamp 0
transform -1 0 5870 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4511_
timestamp 0
transform 1 0 6030 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4512_
timestamp 0
transform 1 0 6130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4513_
timestamp 0
transform 1 0 6150 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4514_
timestamp 0
transform -1 0 1650 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__4515_
timestamp 0
transform -1 0 2490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__4516_
timestamp 0
transform -1 0 4610 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__4517_
timestamp 0
transform -1 0 5090 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4518_
timestamp 0
transform 1 0 5050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4519_
timestamp 0
transform 1 0 5410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4520_
timestamp 0
transform -1 0 5610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4521_
timestamp 0
transform 1 0 6450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4522_
timestamp 0
transform -1 0 8870 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4523_
timestamp 0
transform 1 0 5250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4524_
timestamp 0
transform 1 0 5950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4525_
timestamp 0
transform 1 0 5810 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4526_
timestamp 0
transform -1 0 6390 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4527_
timestamp 0
transform -1 0 4890 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4528_
timestamp 0
transform 1 0 6290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4529_
timestamp 0
transform 1 0 5990 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4530_
timestamp 0
transform 1 0 5970 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4531_
timestamp 0
transform -1 0 2210 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__4532_
timestamp 0
transform -1 0 6230 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4533_
timestamp 0
transform -1 0 6170 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4534_
timestamp 0
transform 1 0 4210 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4535_
timestamp 0
transform 1 0 3610 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4536_
timestamp 0
transform -1 0 1030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4537_
timestamp 0
transform 1 0 4390 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4538_
timestamp 0
transform -1 0 7630 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4539_
timestamp 0
transform -1 0 3010 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4540_
timestamp 0
transform 1 0 7590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4541_
timestamp 0
transform 1 0 6450 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4542_
timestamp 0
transform 1 0 2990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4543_
timestamp 0
transform -1 0 2830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4544_
timestamp 0
transform -1 0 850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4545_
timestamp 0
transform 1 0 2070 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4546_
timestamp 0
transform 1 0 2850 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4547_
timestamp 0
transform -1 0 2310 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4548_
timestamp 0
transform -1 0 1690 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4549_
timestamp 0
transform 1 0 2550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4550_
timestamp 0
transform 1 0 2750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4551_
timestamp 0
transform -1 0 2950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4552_
timestamp 0
transform -1 0 2930 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4553_
timestamp 0
transform -1 0 6490 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4554_
timestamp 0
transform 1 0 930 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4555_
timestamp 0
transform -1 0 690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__4556_
timestamp 0
transform 1 0 4290 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4557_
timestamp 0
transform 1 0 4110 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4558_
timestamp 0
transform -1 0 3950 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4559_
timestamp 0
transform 1 0 4970 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4560_
timestamp 0
transform -1 0 8430 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4561_
timestamp 0
transform -1 0 8830 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4562_
timestamp 0
transform 1 0 8350 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4563_
timestamp 0
transform -1 0 6330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4564_
timestamp 0
transform -1 0 1830 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4565_
timestamp 0
transform 1 0 2650 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4566_
timestamp 0
transform 1 0 3030 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4567_
timestamp 0
transform -1 0 6730 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4568_
timestamp 0
transform 1 0 6650 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4569_
timestamp 0
transform 1 0 1870 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4570_
timestamp 0
transform -1 0 6530 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4571_
timestamp 0
transform 1 0 6230 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4572_
timestamp 0
transform -1 0 9470 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4573_
timestamp 0
transform -1 0 10330 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4574_
timestamp 0
transform -1 0 9510 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4575_
timestamp 0
transform -1 0 6930 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4576_
timestamp 0
transform -1 0 8450 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4577_
timestamp 0
transform -1 0 2970 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4578_
timestamp 0
transform -1 0 5930 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4579_
timestamp 0
transform 1 0 7950 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4580_
timestamp 0
transform 1 0 10130 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4581_
timestamp 0
transform -1 0 7470 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4582_
timestamp 0
transform 1 0 1230 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4583_
timestamp 0
transform -1 0 2310 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4584_
timestamp 0
transform -1 0 2150 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4585_
timestamp 0
transform -1 0 2050 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4586_
timestamp 0
transform -1 0 1870 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4587_
timestamp 0
transform -1 0 1530 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4588_
timestamp 0
transform 1 0 3250 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4589_
timestamp 0
transform 1 0 3790 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4590_
timestamp 0
transform 1 0 1170 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4591_
timestamp 0
transform -1 0 1590 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4592_
timestamp 0
transform 1 0 1390 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4593_
timestamp 0
transform -1 0 3950 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4594_
timestamp 0
transform -1 0 3110 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__4595_
timestamp 0
transform -1 0 2670 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4596_
timestamp 0
transform -1 0 2870 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4597_
timestamp 0
transform 1 0 2730 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__4598_
timestamp 0
transform -1 0 2650 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4599_
timestamp 0
transform -1 0 2830 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4600_
timestamp 0
transform -1 0 3990 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4601_
timestamp 0
transform -1 0 3950 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4602_
timestamp 0
transform -1 0 1370 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4603_
timestamp 0
transform -1 0 1310 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4604_
timestamp 0
transform -1 0 2910 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__4605_
timestamp 0
transform 1 0 1730 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4606_
timestamp 0
transform -1 0 630 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4607_
timestamp 0
transform -1 0 450 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4608_
timestamp 0
transform -1 0 3190 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4609_
timestamp 0
transform 1 0 1570 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__4610_
timestamp 0
transform 1 0 2450 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4611_
timestamp 0
transform -1 0 2290 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4612_
timestamp 0
transform -1 0 1950 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4613_
timestamp 0
transform 1 0 1930 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__4614_
timestamp 0
transform -1 0 590 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4615_
timestamp 0
transform -1 0 410 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4616_
timestamp 0
transform -1 0 1770 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__4617_
timestamp 0
transform -1 0 1570 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__4618_
timestamp 0
transform -1 0 2470 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4619_
timestamp 0
transform -1 0 1810 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4620_
timestamp 0
transform -1 0 1410 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4621_
timestamp 0
transform 1 0 2070 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4622_
timestamp 0
transform 1 0 2490 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4623_
timestamp 0
transform 1 0 1990 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4624_
timestamp 0
transform 1 0 1190 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4625_
timestamp 0
transform 1 0 810 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4626_
timestamp 0
transform -1 0 650 0 1 11290
box -6 -8 26 248
use FILL  FILL_0__4627_
timestamp 0
transform -1 0 2150 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__4628_
timestamp 0
transform -1 0 1210 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__4629_
timestamp 0
transform 1 0 990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0__4630_
timestamp 0
transform 1 0 950 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4631_
timestamp 0
transform 1 0 1530 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4632_
timestamp 0
transform -1 0 690 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4633_
timestamp 0
transform -1 0 510 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4634_
timestamp 0
transform -1 0 7530 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4635_
timestamp 0
transform -1 0 1470 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4636_
timestamp 0
transform 1 0 1270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4637_
timestamp 0
transform -1 0 1670 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4638_
timestamp 0
transform -1 0 830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0__4639_
timestamp 0
transform 1 0 1030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4640_
timestamp 0
transform 1 0 890 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4641_
timestamp 0
transform -1 0 1050 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4642_
timestamp 0
transform -1 0 2870 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__4643_
timestamp 0
transform 1 0 3010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0__4644_
timestamp 0
transform -1 0 3450 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__4645_
timestamp 0
transform -1 0 810 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4646_
timestamp 0
transform 1 0 590 0 1 10810
box -6 -8 26 248
use FILL  FILL_0__4647_
timestamp 0
transform -1 0 1210 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4648_
timestamp 0
transform -1 0 1150 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4649_
timestamp 0
transform -1 0 510 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4650_
timestamp 0
transform -1 0 750 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0__4651_
timestamp 0
transform 1 0 4050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__4652_
timestamp 0
transform 1 0 3770 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__4653_
timestamp 0
transform -1 0 4270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__4654_
timestamp 0
transform -1 0 6830 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4655_
timestamp 0
transform 1 0 2490 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4656_
timestamp 0
transform -1 0 2310 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4657_
timestamp 0
transform -1 0 2230 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4658_
timestamp 0
transform 1 0 3670 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4659_
timestamp 0
transform -1 0 3890 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4660_
timestamp 0
transform -1 0 4270 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4661_
timestamp 0
transform 1 0 4450 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4662_
timestamp 0
transform 1 0 3910 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4663_
timestamp 0
transform 1 0 3350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4664_
timestamp 0
transform 1 0 2490 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4665_
timestamp 0
transform -1 0 7770 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4666_
timestamp 0
transform 1 0 7670 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__4667_
timestamp 0
transform 1 0 6190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__4668_
timestamp 0
transform -1 0 6410 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0__4669_
timestamp 0
transform 1 0 390 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4670_
timestamp 0
transform 1 0 3970 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4671_
timestamp 0
transform 1 0 3790 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4672_
timestamp 0
transform 1 0 2730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4673_
timestamp 0
transform -1 0 2930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4674_
timestamp 0
transform -1 0 3090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4675_
timestamp 0
transform -1 0 2970 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4676_
timestamp 0
transform -1 0 3570 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4677_
timestamp 0
transform -1 0 3510 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4678_
timestamp 0
transform 1 0 3330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4679_
timestamp 0
transform -1 0 3170 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4680_
timestamp 0
transform -1 0 2170 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__4681_
timestamp 0
transform 1 0 1950 0 1 2650
box -6 -8 26 248
use FILL  FILL_0__4682_
timestamp 0
transform -1 0 7010 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4683_
timestamp 0
transform -1 0 1810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4684_
timestamp 0
transform 1 0 3710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4685_
timestamp 0
transform 1 0 3530 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4686_
timestamp 0
transform 1 0 11070 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4687_
timestamp 0
transform 1 0 11250 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4688_
timestamp 0
transform 1 0 11430 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4689_
timestamp 0
transform 1 0 11610 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4690_
timestamp 0
transform 1 0 10450 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4691_
timestamp 0
transform 1 0 10090 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4692_
timestamp 0
transform 1 0 10170 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4693_
timestamp 0
transform -1 0 9690 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4694_
timestamp 0
transform -1 0 9710 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4695_
timestamp 0
transform 1 0 10550 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4696_
timestamp 0
transform 1 0 10870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4697_
timestamp 0
transform 1 0 11350 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4698_
timestamp 0
transform 1 0 11190 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4699_
timestamp 0
transform 1 0 11190 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4700_
timestamp 0
transform 1 0 11030 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4701_
timestamp 0
transform -1 0 11410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4702_
timestamp 0
transform 1 0 11390 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4703_
timestamp 0
transform 1 0 11670 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4704_
timestamp 0
transform -1 0 11570 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4705_
timestamp 0
transform -1 0 11770 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4706_
timestamp 0
transform -1 0 11710 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4707_
timestamp 0
transform 1 0 10650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4708_
timestamp 0
transform 1 0 10850 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4709_
timestamp 0
transform -1 0 10850 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4710_
timestamp 0
transform -1 0 10650 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4711_
timestamp 0
transform 1 0 10110 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4712_
timestamp 0
transform -1 0 9890 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4713_
timestamp 0
transform 1 0 9690 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4714_
timestamp 0
transform 1 0 9490 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4715_
timestamp 0
transform -1 0 9810 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4716_
timestamp 0
transform 1 0 9230 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4717_
timestamp 0
transform 1 0 9570 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4718_
timestamp 0
transform -1 0 8710 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4719_
timestamp 0
transform 1 0 11250 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4720_
timestamp 0
transform 1 0 9990 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4721_
timestamp 0
transform 1 0 9810 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4722_
timestamp 0
transform -1 0 9890 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4723_
timestamp 0
transform -1 0 9890 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4724_
timestamp 0
transform 1 0 4190 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4725_
timestamp 0
transform -1 0 10090 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4726_
timestamp 0
transform -1 0 10290 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4727_
timestamp 0
transform -1 0 11050 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4728_
timestamp 0
transform 1 0 10130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4729_
timestamp 0
transform -1 0 10070 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4730_
timestamp 0
transform -1 0 9950 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4731_
timestamp 0
transform -1 0 11630 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4732_
timestamp 0
transform -1 0 9790 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4733_
timestamp 0
transform 1 0 9770 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4734_
timestamp 0
transform -1 0 7750 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4735_
timestamp 0
transform 1 0 9290 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4736_
timestamp 0
transform -1 0 9990 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4737_
timestamp 0
transform 1 0 9490 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4738_
timestamp 0
transform -1 0 9690 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4739_
timestamp 0
transform -1 0 9870 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4740_
timestamp 0
transform -1 0 10250 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4741_
timestamp 0
transform -1 0 10070 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4742_
timestamp 0
transform 1 0 10290 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4743_
timestamp 0
transform 1 0 10050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4744_
timestamp 0
transform 1 0 10550 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4745_
timestamp 0
transform 1 0 10870 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4746_
timestamp 0
transform 1 0 10350 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4747_
timestamp 0
transform 1 0 8290 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4748_
timestamp 0
transform 1 0 8490 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4749_
timestamp 0
transform -1 0 8730 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4750_
timestamp 0
transform 1 0 8490 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4751_
timestamp 0
transform 1 0 3690 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4752_
timestamp 0
transform -1 0 9090 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4753_
timestamp 0
transform -1 0 7970 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4754_
timestamp 0
transform 1 0 8090 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4755_
timestamp 0
transform 1 0 7210 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4756_
timestamp 0
transform 1 0 6870 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4757_
timestamp 0
transform 1 0 8310 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4758_
timestamp 0
transform -1 0 10370 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4759_
timestamp 0
transform 1 0 10730 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4760_
timestamp 0
transform -1 0 11010 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4761_
timestamp 0
transform 1 0 11290 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4762_
timestamp 0
transform -1 0 10450 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4763_
timestamp 0
transform 1 0 11790 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4764_
timestamp 0
transform 1 0 10830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4765_
timestamp 0
transform -1 0 11090 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4766_
timestamp 0
transform -1 0 10450 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4767_
timestamp 0
transform -1 0 10470 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4768_
timestamp 0
transform 1 0 10250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4769_
timestamp 0
transform 1 0 10630 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4770_
timestamp 0
transform 1 0 11110 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4771_
timestamp 0
transform 1 0 11970 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4772_
timestamp 0
transform 1 0 9310 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4773_
timestamp 0
transform -1 0 8770 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4774_
timestamp 0
transform 1 0 2510 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4775_
timestamp 0
transform 1 0 2670 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4776_
timestamp 0
transform 1 0 2830 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4777_
timestamp 0
transform -1 0 3050 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4778_
timestamp 0
transform -1 0 3650 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4779_
timestamp 0
transform 1 0 3830 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4780_
timestamp 0
transform -1 0 8710 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4781_
timestamp 0
transform 1 0 3550 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4782_
timestamp 0
transform 1 0 3230 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4783_
timestamp 0
transform 1 0 9050 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4784_
timestamp 0
transform 1 0 7690 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4785_
timestamp 0
transform 1 0 2050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4786_
timestamp 0
transform -1 0 3930 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__4787_
timestamp 0
transform -1 0 3610 0 1 3130
box -6 -8 26 248
use FILL  FILL_0__4788_
timestamp 0
transform -1 0 4130 0 1 3610
box -6 -8 26 248
use FILL  FILL_0__4789_
timestamp 0
transform 1 0 7170 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4790_
timestamp 0
transform 1 0 7230 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4791_
timestamp 0
transform -1 0 7770 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4792_
timestamp 0
transform -1 0 7830 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4793_
timestamp 0
transform -1 0 7770 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4794_
timestamp 0
transform -1 0 7410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4795_
timestamp 0
transform -1 0 7470 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4796_
timestamp 0
transform 1 0 11770 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4797_
timestamp 0
transform 1 0 8510 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4798_
timestamp 0
transform 1 0 9970 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4799_
timestamp 0
transform -1 0 9810 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4800_
timestamp 0
transform 1 0 8450 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4801_
timestamp 0
transform 1 0 10910 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4802_
timestamp 0
transform -1 0 10450 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4803_
timestamp 0
transform -1 0 7350 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4804_
timestamp 0
transform -1 0 7030 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4805_
timestamp 0
transform -1 0 6910 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4806_
timestamp 0
transform -1 0 9270 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4807_
timestamp 0
transform -1 0 9050 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4808_
timestamp 0
transform -1 0 8670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4809_
timestamp 0
transform -1 0 8670 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4810_
timestamp 0
transform -1 0 8910 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4811_
timestamp 0
transform 1 0 11890 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4812_
timestamp 0
transform 1 0 11970 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4813_
timestamp 0
transform 1 0 11430 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4814_
timestamp 0
transform 1 0 11310 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4815_
timestamp 0
transform -1 0 9010 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4816_
timestamp 0
transform -1 0 9450 0 1 7450
box -6 -8 26 248
use FILL  FILL_0__4817_
timestamp 0
transform -1 0 11510 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4818_
timestamp 0
transform -1 0 11450 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4819_
timestamp 0
transform -1 0 6390 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4820_
timestamp 0
transform 1 0 7950 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4821_
timestamp 0
transform 1 0 11590 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4822_
timestamp 0
transform 1 0 11790 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4823_
timestamp 0
transform 1 0 11570 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4824_
timestamp 0
transform -1 0 11430 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4825_
timestamp 0
transform 1 0 11130 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4826_
timestamp 0
transform -1 0 10970 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4827_
timestamp 0
transform -1 0 11670 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4828_
timestamp 0
transform -1 0 11750 0 1 10330
box -6 -8 26 248
use FILL  FILL_0__4829_
timestamp 0
transform 1 0 11590 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4830_
timestamp 0
transform 1 0 8950 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4831_
timestamp 0
transform -1 0 9310 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4832_
timestamp 0
transform 1 0 11850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4833_
timestamp 0
transform 1 0 8330 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4834_
timestamp 0
transform 1 0 8130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4835_
timestamp 0
transform -1 0 8330 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4836_
timestamp 0
transform 1 0 9610 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4837_
timestamp 0
transform -1 0 10750 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4838_
timestamp 0
transform 1 0 11770 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4839_
timestamp 0
transform 1 0 12030 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4840_
timestamp 0
transform 1 0 9210 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4841_
timestamp 0
transform 1 0 10250 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4842_
timestamp 0
transform 1 0 11950 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4843_
timestamp 0
transform 1 0 11110 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4844_
timestamp 0
transform -1 0 11090 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4845_
timestamp 0
transform -1 0 11870 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4846_
timestamp 0
transform 1 0 11850 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4847_
timestamp 0
transform -1 0 8330 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0__4848_
timestamp 0
transform -1 0 8350 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4849_
timestamp 0
transform 1 0 9010 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4850_
timestamp 0
transform 1 0 9250 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4851_
timestamp 0
transform 1 0 11230 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4852_
timestamp 0
transform 1 0 11610 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4853_
timestamp 0
transform 1 0 12010 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4854_
timestamp 0
transform -1 0 11150 0 1 11770
box -6 -8 26 248
use FILL  FILL_0__4855_
timestamp 0
transform -1 0 8170 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4856_
timestamp 0
transform -1 0 8190 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4857_
timestamp 0
transform -1 0 10270 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4858_
timestamp 0
transform -1 0 10410 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4859_
timestamp 0
transform -1 0 7150 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4860_
timestamp 0
transform -1 0 10330 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4861_
timestamp 0
transform -1 0 10590 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4862_
timestamp 0
transform 1 0 11390 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4863_
timestamp 0
transform -1 0 10650 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4864_
timestamp 0
transform -1 0 10490 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4865_
timestamp 0
transform 1 0 10510 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4866_
timestamp 0
transform 1 0 11590 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4867_
timestamp 0
transform 1 0 11770 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4868_
timestamp 0
transform -1 0 11270 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4869_
timestamp 0
transform -1 0 10810 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0__4870_
timestamp 0
transform 1 0 8050 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4871_
timestamp 0
transform 1 0 7890 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4872_
timestamp 0
transform 1 0 7790 0 1 7930
box -6 -8 26 248
use FILL  FILL_0__4873_
timestamp 0
transform -1 0 11310 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4874_
timestamp 0
transform 1 0 11830 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4875_
timestamp 0
transform -1 0 7530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0__4876_
timestamp 0
transform -1 0 10450 0 -1 9370
box -6 -8 26 248
use FILL  FILL_0__4877_
timestamp 0
transform 1 0 10850 0 1 8410
box -6 -8 26 248
use FILL  FILL_0__4878_
timestamp 0
transform 1 0 11290 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4879_
timestamp 0
transform 1 0 11950 0 1 9850
box -6 -8 26 248
use FILL  FILL_0__4880_
timestamp 0
transform -1 0 12010 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4881_
timestamp 0
transform -1 0 9050 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4882_
timestamp 0
transform 1 0 11970 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4883_
timestamp 0
transform 1 0 11790 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4884_
timestamp 0
transform 1 0 11610 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4885_
timestamp 0
transform -1 0 11650 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4886_
timestamp 0
transform 1 0 10910 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4887_
timestamp 0
transform 1 0 10950 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4888_
timestamp 0
transform 1 0 11610 0 1 8890
box -6 -8 26 248
use FILL  FILL_0__4889_
timestamp 0
transform 1 0 11950 0 1 9370
box -6 -8 26 248
use FILL  FILL_0__4890_
timestamp 0
transform 1 0 11470 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4891_
timestamp 0
transform 1 0 11810 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0__4892_
timestamp 0
transform -1 0 12030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0__4893_
timestamp 0
transform -1 0 2450 0 -1 7450
box -6 -8 26 248
use FILL  FILL_0__4894_
timestamp 0
transform 1 0 9650 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4895_
timestamp 0
transform 1 0 8390 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4896_
timestamp 0
transform -1 0 9430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4897_
timestamp 0
transform 1 0 9470 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4898_
timestamp 0
transform 1 0 9650 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4899_
timestamp 0
transform -1 0 9130 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4900_
timestamp 0
transform -1 0 9470 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4901_
timestamp 0
transform -1 0 9850 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4902_
timestamp 0
transform 1 0 10170 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4903_
timestamp 0
transform 1 0 9630 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4904_
timestamp 0
transform -1 0 10350 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4905_
timestamp 0
transform 1 0 9630 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4906_
timestamp 0
transform -1 0 9810 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4907_
timestamp 0
transform -1 0 9470 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4908_
timestamp 0
transform 1 0 9970 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4909_
timestamp 0
transform 1 0 10910 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4910_
timestamp 0
transform -1 0 11290 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4911_
timestamp 0
transform 1 0 11230 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4912_
timestamp 0
transform 1 0 11050 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4913_
timestamp 0
transform -1 0 10870 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4914_
timestamp 0
transform 1 0 11430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4915_
timestamp 0
transform -1 0 10730 0 1 6970
box -6 -8 26 248
use FILL  FILL_0__4916_
timestamp 0
transform 1 0 10490 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4917_
timestamp 0
transform -1 0 10550 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4918_
timestamp 0
transform -1 0 10910 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4919_
timestamp 0
transform 1 0 11070 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4920_
timestamp 0
transform 1 0 8490 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4921_
timestamp 0
transform -1 0 8710 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4922_
timestamp 0
transform -1 0 8910 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4923_
timestamp 0
transform 1 0 9290 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4924_
timestamp 0
transform 1 0 9270 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4925_
timestamp 0
transform -1 0 9090 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4926_
timestamp 0
transform 1 0 8850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4927_
timestamp 0
transform -1 0 11250 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4928_
timestamp 0
transform 1 0 11430 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4929_
timestamp 0
transform 1 0 12010 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4930_
timestamp 0
transform 1 0 11590 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4931_
timestamp 0
transform -1 0 11810 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4932_
timestamp 0
transform -1 0 11650 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4933_
timestamp 0
transform -1 0 11090 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4934_
timestamp 0
transform 1 0 10870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4935_
timestamp 0
transform -1 0 10690 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4936_
timestamp 0
transform -1 0 9590 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4937_
timestamp 0
transform -1 0 9810 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4938_
timestamp 0
transform 1 0 9970 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4939_
timestamp 0
transform 1 0 10050 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4940_
timestamp 0
transform 1 0 10150 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0__4941_
timestamp 0
transform 1 0 10250 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4942_
timestamp 0
transform -1 0 10650 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4943_
timestamp 0
transform 1 0 11630 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4944_
timestamp 0
transform -1 0 11850 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4945_
timestamp 0
transform 1 0 11790 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4946_
timestamp 0
transform -1 0 11770 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4947_
timestamp 0
transform -1 0 8590 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4948_
timestamp 0
transform 1 0 8910 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4949_
timestamp 0
transform 1 0 12030 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__4950_
timestamp 0
transform -1 0 11990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4951_
timestamp 0
transform -1 0 8530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4952_
timestamp 0
transform 1 0 8910 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4953_
timestamp 0
transform -1 0 8810 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4954_
timestamp 0
transform -1 0 9110 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4955_
timestamp 0
transform -1 0 8670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__4956_
timestamp 0
transform -1 0 8750 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4957_
timestamp 0
transform -1 0 8610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4958_
timestamp 0
transform -1 0 10990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4959_
timestamp 0
transform 1 0 11170 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4960_
timestamp 0
transform -1 0 11390 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4961_
timestamp 0
transform 1 0 11570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4962_
timestamp 0
transform 1 0 11970 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4963_
timestamp 0
transform 1 0 11930 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4964_
timestamp 0
transform 1 0 11930 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4965_
timestamp 0
transform -1 0 11770 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4966_
timestamp 0
transform -1 0 9110 0 1 4090
box -6 -8 26 248
use FILL  FILL_0__4967_
timestamp 0
transform 1 0 8030 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__4968_
timestamp 0
transform 1 0 11610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4969_
timestamp 0
transform 1 0 11970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4970_
timestamp 0
transform 1 0 9010 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4971_
timestamp 0
transform -1 0 8230 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4972_
timestamp 0
transform -1 0 8630 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4973_
timestamp 0
transform -1 0 8790 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4974_
timestamp 0
transform 1 0 8690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4975_
timestamp 0
transform 1 0 8890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4976_
timestamp 0
transform 1 0 11550 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4977_
timestamp 0
transform 1 0 11350 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4978_
timestamp 0
transform 1 0 11370 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4979_
timestamp 0
transform 1 0 11390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4980_
timestamp 0
transform 1 0 11770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4981_
timestamp 0
transform -1 0 11770 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4982_
timestamp 0
transform -1 0 11790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4983_
timestamp 0
transform 1 0 11570 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4984_
timestamp 0
transform 1 0 11190 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4985_
timestamp 0
transform -1 0 8010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4986_
timestamp 0
transform 1 0 9050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4987_
timestamp 0
transform 1 0 11570 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4988_
timestamp 0
transform -1 0 11790 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4989_
timestamp 0
transform -1 0 11390 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4990_
timestamp 0
transform -1 0 11210 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__4991_
timestamp 0
transform 1 0 11590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__4992_
timestamp 0
transform -1 0 11450 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4993_
timestamp 0
transform 1 0 11230 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__4994_
timestamp 0
transform 1 0 9250 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__4995_
timestamp 0
transform -1 0 9830 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4996_
timestamp 0
transform 1 0 9190 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4997_
timestamp 0
transform -1 0 9270 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__4998_
timestamp 0
transform 1 0 9370 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__4999_
timestamp 0
transform -1 0 9230 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5000_
timestamp 0
transform 1 0 10970 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__5001_
timestamp 0
transform -1 0 10790 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__5002_
timestamp 0
transform -1 0 10610 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5003_
timestamp 0
transform -1 0 10670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5004_
timestamp 0
transform 1 0 10850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5005_
timestamp 0
transform -1 0 10830 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5006_
timestamp 0
transform 1 0 11350 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5007_
timestamp 0
transform 1 0 11950 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5008_
timestamp 0
transform 1 0 11930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__5009_
timestamp 0
transform 1 0 11950 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5010_
timestamp 0
transform -1 0 11250 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__5011_
timestamp 0
transform 1 0 11750 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5012_
timestamp 0
transform 1 0 11550 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5013_
timestamp 0
transform -1 0 10230 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5014_
timestamp 0
transform -1 0 9450 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5015_
timestamp 0
transform 1 0 8210 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5016_
timestamp 0
transform 1 0 10610 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5017_
timestamp 0
transform 1 0 8870 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5018_
timestamp 0
transform 1 0 8410 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5019_
timestamp 0
transform 1 0 9090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5020_
timestamp 0
transform 1 0 8990 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5021_
timestamp 0
transform 1 0 9270 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5022_
timestamp 0
transform -1 0 9070 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5023_
timestamp 0
transform -1 0 10790 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__5024_
timestamp 0
transform 1 0 10790 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5025_
timestamp 0
transform -1 0 11010 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5026_
timestamp 0
transform 1 0 11030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__5027_
timestamp 0
transform -1 0 10830 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5028_
timestamp 0
transform -1 0 10650 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5029_
timestamp 0
transform 1 0 10990 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5030_
timestamp 0
transform 1 0 11010 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5031_
timestamp 0
transform 1 0 11770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__5032_
timestamp 0
transform 1 0 11610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__5033_
timestamp 0
transform -1 0 8930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__5034_
timestamp 0
transform -1 0 9130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__5035_
timestamp 0
transform 1 0 11150 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5036_
timestamp 0
transform 1 0 9830 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5037_
timestamp 0
transform 1 0 9630 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5038_
timestamp 0
transform 1 0 9470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5039_
timestamp 0
transform 1 0 9410 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5040_
timestamp 0
transform 1 0 9650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5041_
timestamp 0
transform 1 0 9850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5042_
timestamp 0
transform 1 0 10570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__5043_
timestamp 0
transform 1 0 10390 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5044_
timestamp 0
transform 1 0 10450 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5045_
timestamp 0
transform -1 0 10430 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5046_
timestamp 0
transform 1 0 10870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__5047_
timestamp 0
transform 1 0 10970 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5048_
timestamp 0
transform 1 0 11410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__5049_
timestamp 0
transform -1 0 11250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__5050_
timestamp 0
transform -1 0 9310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__5051_
timestamp 0
transform 1 0 8310 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__5052_
timestamp 0
transform -1 0 10470 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__5053_
timestamp 0
transform -1 0 10710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__5054_
timestamp 0
transform -1 0 10350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__5055_
timestamp 0
transform 1 0 8470 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__5056_
timestamp 0
transform 1 0 8090 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__5057_
timestamp 0
transform 1 0 8310 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__5058_
timestamp 0
transform -1 0 8130 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__5059_
timestamp 0
transform 1 0 7950 0 1 6490
box -6 -8 26 248
use FILL  FILL_0__5060_
timestamp 0
transform -1 0 7590 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__5061_
timestamp 0
transform -1 0 7770 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__5062_
timestamp 0
transform 1 0 7930 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0__5063_
timestamp 0
transform -1 0 7970 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__5064_
timestamp 0
transform -1 0 7490 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5065_
timestamp 0
transform -1 0 7690 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5066_
timestamp 0
transform -1 0 7630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5067_
timestamp 0
transform -1 0 8330 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5068_
timestamp 0
transform -1 0 8350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5069_
timestamp 0
transform -1 0 8190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5070_
timestamp 0
transform -1 0 7810 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5071_
timestamp 0
transform 1 0 7990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5072_
timestamp 0
transform -1 0 7450 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5073_
timestamp 0
transform 1 0 7250 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5074_
timestamp 0
transform 1 0 4810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0__5075_
timestamp 0
transform 1 0 10210 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__5076_
timestamp 0
transform 1 0 10010 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__5077_
timestamp 0
transform 1 0 9790 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__5078_
timestamp 0
transform 1 0 9570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__5079_
timestamp 0
transform 1 0 9970 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__5080_
timestamp 0
transform 1 0 10170 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__5081_
timestamp 0
transform 1 0 10390 0 1 6010
box -6 -8 26 248
use FILL  FILL_0__5082_
timestamp 0
transform 1 0 10370 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0__5083_
timestamp 0
transform -1 0 10270 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5084_
timestamp 0
transform -1 0 9650 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5085_
timestamp 0
transform 1 0 8490 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5086_
timestamp 0
transform -1 0 8690 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5087_
timestamp 0
transform -1 0 10850 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__5088_
timestamp 0
transform -1 0 10630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__5089_
timestamp 0
transform -1 0 10430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__5090_
timestamp 0
transform -1 0 10210 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5091_
timestamp 0
transform 1 0 10050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0__5092_
timestamp 0
transform 1 0 9890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__5093_
timestamp 0
transform -1 0 10070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__5094_
timestamp 0
transform 1 0 10210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__5095_
timestamp 0
transform -1 0 9730 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__5096_
timestamp 0
transform 1 0 8870 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__5097_
timestamp 0
transform 1 0 8190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0__5098_
timestamp 0
transform 1 0 9690 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5099_
timestamp 0
transform 1 0 9870 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5100_
timestamp 0
transform 1 0 9310 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5101_
timestamp 0
transform -1 0 10030 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5102_
timestamp 0
transform -1 0 9850 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5103_
timestamp 0
transform 1 0 9990 0 1 5050
box -6 -8 26 248
use FILL  FILL_0__5104_
timestamp 0
transform -1 0 10290 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5105_
timestamp 0
transform -1 0 10090 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5106_
timestamp 0
transform -1 0 10470 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5107_
timestamp 0
transform 1 0 10450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__5108_
timestamp 0
transform -1 0 11050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__5109_
timestamp 0
transform 1 0 10650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0__5110_
timestamp 0
transform -1 0 9510 0 1 4570
box -6 -8 26 248
use FILL  FILL_0__5111_
timestamp 0
transform -1 0 7870 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5112_
timestamp 0
transform -1 0 8050 0 1 5530
box -6 -8 26 248
use FILL  FILL_0__5124_
timestamp 0
transform 1 0 1730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__5125_
timestamp 0
transform -1 0 590 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__5126_
timestamp 0
transform -1 0 770 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__5127_
timestamp 0
transform 1 0 730 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__5128_
timestamp 0
transform 1 0 490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__5129_
timestamp 0
transform 1 0 930 0 1 2170
box -6 -8 26 248
use FILL  FILL_0__5130_
timestamp 0
transform 1 0 930 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__5131_
timestamp 0
transform -1 0 2250 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5132_
timestamp 0
transform -1 0 5490 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5133_
timestamp 0
transform 1 0 5230 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5134_
timestamp 0
transform 1 0 1310 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__5135_
timestamp 0
transform 1 0 2110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__5136_
timestamp 0
transform 1 0 1910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__5137_
timestamp 0
transform -1 0 1050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__5138_
timestamp 0
transform -1 0 1230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__5139_
timestamp 0
transform -1 0 3610 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5140_
timestamp 0
transform 1 0 4070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__5141_
timestamp 0
transform -1 0 4250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__5142_
timestamp 0
transform -1 0 4130 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__5143_
timestamp 0
transform -1 0 4350 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5144_
timestamp 0
transform 1 0 5510 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5145_
timestamp 0
transform -1 0 4050 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5146_
timestamp 0
transform -1 0 4570 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5147_
timestamp 0
transform 1 0 4670 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5148_
timestamp 0
transform 1 0 4870 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5149_
timestamp 0
transform 1 0 5390 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5150_
timestamp 0
transform -1 0 6010 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5151_
timestamp 0
transform 1 0 3390 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5152_
timestamp 0
transform 1 0 5650 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5153_
timestamp 0
transform 1 0 4130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__5154_
timestamp 0
transform 1 0 5330 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5155_
timestamp 0
transform 1 0 5290 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5156_
timestamp 0
transform 1 0 5450 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5157_
timestamp 0
transform 1 0 5590 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5158_
timestamp 0
transform 1 0 4470 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5159_
timestamp 0
transform -1 0 4590 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5160_
timestamp 0
transform 1 0 4910 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5161_
timestamp 0
transform 1 0 4750 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5162_
timestamp 0
transform 1 0 5790 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5163_
timestamp 0
transform -1 0 2690 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5164_
timestamp 0
transform 1 0 5810 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5165_
timestamp 0
transform -1 0 3750 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__5166_
timestamp 0
transform 1 0 4190 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5167_
timestamp 0
transform 1 0 4150 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5168_
timestamp 0
transform -1 0 3970 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5169_
timestamp 0
transform 1 0 2650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__5170_
timestamp 0
transform 1 0 3770 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5171_
timestamp 0
transform -1 0 4070 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__5172_
timestamp 0
transform -1 0 3570 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__5173_
timestamp 0
transform -1 0 4850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__5174_
timestamp 0
transform -1 0 3750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__5175_
timestamp 0
transform 1 0 3590 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5176_
timestamp 0
transform -1 0 2590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__5177_
timestamp 0
transform 1 0 3030 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5178_
timestamp 0
transform 1 0 4370 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5179_
timestamp 0
transform 1 0 4390 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5180_
timestamp 0
transform 1 0 4190 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5181_
timestamp 0
transform 1 0 3190 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5182_
timestamp 0
transform -1 0 2390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__5183_
timestamp 0
transform 1 0 2190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__5184_
timestamp 0
transform -1 0 2410 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__5185_
timestamp 0
transform -1 0 3970 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__5186_
timestamp 0
transform -1 0 3250 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__5187_
timestamp 0
transform -1 0 2990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__5188_
timestamp 0
transform 1 0 3690 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5189_
timestamp 0
transform -1 0 3630 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5190_
timestamp 0
transform 1 0 3170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__5191_
timestamp 0
transform 1 0 2850 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5192_
timestamp 0
transform -1 0 3570 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__5193_
timestamp 0
transform 1 0 6010 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5194_
timestamp 0
transform -1 0 2870 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__5195_
timestamp 0
transform -1 0 2790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__5196_
timestamp 0
transform 1 0 3530 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5197_
timestamp 0
transform -1 0 3450 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5198_
timestamp 0
transform -1 0 2850 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5199_
timestamp 0
transform 1 0 2410 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5200_
timestamp 0
transform -1 0 2630 0 -1 730
box -6 -8 26 248
use FILL  FILL_0__5201_
timestamp 0
transform -1 0 3910 0 1 1690
box -6 -8 26 248
use FILL  FILL_0__5202_
timestamp 0
transform 1 0 3870 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5203_
timestamp 0
transform -1 0 3410 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5204_
timestamp 0
transform 1 0 4030 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5205_
timestamp 0
transform -1 0 3870 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5206_
timestamp 0
transform -1 0 3210 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5207_
timestamp 0
transform 1 0 2430 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5208_
timestamp 0
transform 1 0 2970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__5209_
timestamp 0
transform -1 0 4430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0__5210_
timestamp 0
transform 1 0 2630 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5211_
timestamp 0
transform 1 0 2790 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5212_
timestamp 0
transform 1 0 3370 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5213_
timestamp 0
transform 1 0 3250 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5214_
timestamp 0
transform -1 0 3010 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5215_
timestamp 0
transform 1 0 2230 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5216_
timestamp 0
transform -1 0 3030 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__5217_
timestamp 0
transform -1 0 6190 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5218_
timestamp 0
transform 1 0 3370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__5219_
timestamp 0
transform 1 0 3530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__5220_
timestamp 0
transform 1 0 4710 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5221_
timestamp 0
transform 1 0 4530 0 -1 250
box -6 -8 26 248
use FILL  FILL_0__5222_
timestamp 0
transform -1 0 4010 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5223_
timestamp 0
transform 1 0 3050 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5224_
timestamp 0
transform -1 0 3810 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5225_
timestamp 0
transform 1 0 5310 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__5226_
timestamp 0
transform 1 0 5090 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5227_
timestamp 0
transform -1 0 5270 0 1 250
box -6 -8 26 248
use FILL  FILL_0__5228_
timestamp 0
transform -1 0 4710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0__5229_
timestamp 0
transform -1 0 4750 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5230_
timestamp 0
transform 1 0 4930 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5231_
timestamp 0
transform 1 0 5130 0 1 730
box -6 -8 26 248
use FILL  FILL_0__5232_
timestamp 0
transform 1 0 3930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0__5233_
timestamp 0
transform 1 0 4310 0 1 1210
box -6 -8 26 248
use FILL  FILL_0__5234_
timestamp 0
transform -1 0 5110 0 1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert0
timestamp 0
transform -1 0 4150 0 1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert1
timestamp 0
transform 1 0 6070 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert2
timestamp 0
transform -1 0 3250 0 1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert3
timestamp 0
transform -1 0 3630 0 1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert4
timestamp 0
transform 1 0 9410 0 1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert5
timestamp 0
transform 1 0 11210 0 1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert6
timestamp 0
transform -1 0 9410 0 1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert7
timestamp 0
transform 1 0 11950 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert8
timestamp 0
transform -1 0 7110 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert9
timestamp 0
transform 1 0 6610 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert10
timestamp 0
transform 1 0 8650 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert11
timestamp 0
transform 1 0 6810 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert12
timestamp 0
transform 1 0 8850 0 1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert13
timestamp 0
transform 1 0 7330 0 1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert14
timestamp 0
transform 1 0 590 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert15
timestamp 0
transform 1 0 10 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert16
timestamp 0
transform 1 0 1830 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert17
timestamp 0
transform -1 0 9090 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert18
timestamp 0
transform -1 0 11450 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert19
timestamp 0
transform 1 0 10610 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert20
timestamp 0
transform -1 0 9130 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert21
timestamp 0
transform 1 0 2470 0 1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert22
timestamp 0
transform -1 0 1210 0 1 11290
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert23
timestamp 0
transform -1 0 1390 0 1 11290
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert24
timestamp 0
transform -1 0 1590 0 1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert38
timestamp 0
transform -1 0 11470 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert39
timestamp 0
transform -1 0 10610 0 1 6010
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert40
timestamp 0
transform 1 0 11970 0 1 6970
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert41
timestamp 0
transform -1 0 11190 0 1 6010
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert42
timestamp 0
transform 1 0 11390 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert43
timestamp 0
transform -1 0 10950 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert44
timestamp 0
transform -1 0 10430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert45
timestamp 0
transform -1 0 11310 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert46
timestamp 0
transform -1 0 10690 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert47
timestamp 0
transform 1 0 6150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert48
timestamp 0
transform -1 0 4710 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert49
timestamp 0
transform 1 0 11510 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert50
timestamp 0
transform -1 0 10350 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert51
timestamp 0
transform 1 0 8110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert52
timestamp 0
transform 1 0 9970 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert53
timestamp 0
transform 1 0 9130 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert54
timestamp 0
transform 1 0 8950 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert55
timestamp 0
transform -1 0 9490 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert56
timestamp 0
transform -1 0 8790 0 1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert57
timestamp 0
transform 1 0 11410 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert58
timestamp 0
transform 1 0 10590 0 -1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert59
timestamp 0
transform -1 0 7670 0 -1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert60
timestamp 0
transform 1 0 11750 0 -1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert61
timestamp 0
transform 1 0 11850 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert62
timestamp 0
transform -1 0 4750 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert63
timestamp 0
transform -1 0 9270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert64
timestamp 0
transform -1 0 11610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert65
timestamp 0
transform -1 0 9270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert66
timestamp 0
transform -1 0 11450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert67
timestamp 0
transform 1 0 6870 0 1 11290
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert68
timestamp 0
transform -1 0 3110 0 -1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert69
timestamp 0
transform -1 0 5570 0 1 10810
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert70
timestamp 0
transform 1 0 5050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert71
timestamp 0
transform -1 0 3510 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert72
timestamp 0
transform 1 0 7050 0 1 11290
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert73
timestamp 0
transform 1 0 7070 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert74
timestamp 0
transform -1 0 6410 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert75
timestamp 0
transform 1 0 7030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert76
timestamp 0
transform 1 0 6490 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert77
timestamp 0
transform 1 0 10210 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert78
timestamp 0
transform 1 0 9070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert79
timestamp 0
transform 1 0 10230 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert80
timestamp 0
transform -1 0 4890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert81
timestamp 0
transform -1 0 2750 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert82
timestamp 0
transform -1 0 3970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert83
timestamp 0
transform -1 0 6230 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert84
timestamp 0
transform 1 0 7290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert85
timestamp 0
transform -1 0 3210 0 1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert86
timestamp 0
transform 1 0 3910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert87
timestamp 0
transform -1 0 3170 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert88
timestamp 0
transform 1 0 7830 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert89
timestamp 0
transform -1 0 4670 0 1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert90
timestamp 0
transform 1 0 5510 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert91
timestamp 0
transform 1 0 8970 0 1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert92
timestamp 0
transform -1 0 8470 0 1 10810
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert93
timestamp 0
transform -1 0 10870 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert94
timestamp 0
transform 1 0 7210 0 1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert95
timestamp 0
transform 1 0 11470 0 1 10810
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert96
timestamp 0
transform -1 0 4930 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert97
timestamp 0
transform 1 0 550 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert98
timestamp 0
transform -1 0 3950 0 1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert99
timestamp 0
transform 1 0 490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert100
timestamp 0
transform 1 0 2970 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert101
timestamp 0
transform -1 0 430 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert102
timestamp 0
transform 1 0 3670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert103
timestamp 0
transform -1 0 3590 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert104
timestamp 0
transform 1 0 4570 0 1 10330
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert105
timestamp 0
transform 1 0 230 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert106
timestamp 0
transform 1 0 6450 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert107
timestamp 0
transform -1 0 6150 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert108
timestamp 0
transform 1 0 5630 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert109
timestamp 0
transform 1 0 7770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert110
timestamp 0
transform -1 0 5270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert111
timestamp 0
transform 1 0 7230 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert112
timestamp 0
transform 1 0 10610 0 1 11770
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert113
timestamp 0
transform -1 0 12050 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert114
timestamp 0
transform -1 0 10250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert115
timestamp 0
transform 1 0 7310 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert116
timestamp 0
transform -1 0 5450 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert117
timestamp 0
transform -1 0 5430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert118
timestamp 0
transform -1 0 11130 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert119
timestamp 0
transform 1 0 10310 0 1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert120
timestamp 0
transform -1 0 11050 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert121
timestamp 0
transform -1 0 8110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert122
timestamp 0
transform 1 0 11130 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert123
timestamp 0
transform -1 0 9970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert124
timestamp 0
transform -1 0 7950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert125
timestamp 0
transform -1 0 5270 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert126
timestamp 0
transform 1 0 11950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert127
timestamp 0
transform 1 0 10710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert128
timestamp 0
transform -1 0 11990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert129
timestamp 0
transform 1 0 10390 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert130
timestamp 0
transform 1 0 11950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert131
timestamp 0
transform -1 0 9310 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert132
timestamp 0
transform -1 0 8650 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert133
timestamp 0
transform 1 0 11950 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert134
timestamp 0
transform -1 0 11330 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert135
timestamp 0
transform -1 0 9050 0 -1 250
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert136
timestamp 0
transform 1 0 9410 0 -1 250
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert137
timestamp 0
transform -1 0 6330 0 1 730
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert138
timestamp 0
transform 1 0 8310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert139
timestamp 0
transform -1 0 6350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert140
timestamp 0
transform 1 0 9370 0 1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert141
timestamp 0
transform -1 0 6990 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert142
timestamp 0
transform -1 0 6970 0 1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert143
timestamp 0
transform -1 0 6390 0 -1 6970
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert144
timestamp 0
transform -1 0 6210 0 1 6970
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert145
timestamp 0
transform 1 0 9490 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert146
timestamp 0
transform 1 0 9590 0 1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert147
timestamp 0
transform -1 0 7670 0 1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert148
timestamp 0
transform -1 0 7590 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert149
timestamp 0
transform -1 0 9170 0 -1 7930
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert150
timestamp 0
transform -1 0 7170 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert151
timestamp 0
transform 1 0 7270 0 -1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert152
timestamp 0
transform -1 0 8170 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert153
timestamp 0
transform 1 0 10010 0 -1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert154
timestamp 0
transform 1 0 10690 0 -1 8410
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert155
timestamp 0
transform 1 0 6330 0 1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert156
timestamp 0
transform 1 0 9070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert157
timestamp 0
transform -1 0 5810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert158
timestamp 0
transform 1 0 9810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert159
timestamp 0
transform 1 0 8670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert160
timestamp 0
transform 1 0 10310 0 1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert161
timestamp 0
transform 1 0 9210 0 1 9850
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert162
timestamp 0
transform 1 0 10170 0 1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert163
timestamp 0
transform -1 0 8270 0 1 8890
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert164
timestamp 0
transform 1 0 11670 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert165
timestamp 0
transform -1 0 8730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert166
timestamp 0
transform -1 0 11510 0 1 4090
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert167
timestamp 0
transform 1 0 11670 0 1 11770
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert168
timestamp 0
transform -1 0 11250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_BUFX2_insert169
timestamp 0
transform 1 0 4870 0 1 1690
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert25
timestamp 0
transform 1 0 1310 0 1 2170
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert26
timestamp 0
transform 1 0 3970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert27
timestamp 0
transform -1 0 30 0 -1 2650
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert28
timestamp 0
transform -1 0 2670 0 1 9370
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert29
timestamp 0
transform 1 0 10 0 -1 2170
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert30
timestamp 0
transform 1 0 6130 0 -1 5050
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert31
timestamp 0
transform 1 0 730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert32
timestamp 0
transform -1 0 4770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert33
timestamp 0
transform -1 0 910 0 -1 10810
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert34
timestamp 0
transform 1 0 1350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert35
timestamp 0
transform -1 0 270 0 -1 11770
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert36
timestamp 0
transform 1 0 10 0 1 5530
box -6 -8 26 248
use FILL  FILL_0_CLKBUF1_insert37
timestamp 0
transform 1 0 6090 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__2478_
timestamp 0
transform -1 0 50 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2479_
timestamp 0
transform -1 0 50 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2480_
timestamp 0
transform 1 0 1890 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2481_
timestamp 0
transform 1 0 2710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2482_
timestamp 0
transform -1 0 50 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__2483_
timestamp 0
transform -1 0 530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__2484_
timestamp 0
transform -1 0 2090 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2485_
timestamp 0
transform 1 0 3910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2486_
timestamp 0
transform 1 0 12030 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2487_
timestamp 0
transform -1 0 6610 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2488_
timestamp 0
transform -1 0 6790 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2489_
timestamp 0
transform 1 0 11990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2490_
timestamp 0
transform 1 0 11990 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2491_
timestamp 0
transform 1 0 6410 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2492_
timestamp 0
transform 1 0 11810 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2493_
timestamp 0
transform -1 0 11910 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2494_
timestamp 0
transform -1 0 1010 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__2495_
timestamp 0
transform -1 0 1170 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2496_
timestamp 0
transform -1 0 50 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__2497_
timestamp 0
transform -1 0 4390 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2498_
timestamp 0
transform 1 0 4430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2499_
timestamp 0
transform -1 0 3250 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2500_
timestamp 0
transform -1 0 430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2501_
timestamp 0
transform -1 0 3630 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2502_
timestamp 0
transform -1 0 50 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__2503_
timestamp 0
transform -1 0 50 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2504_
timestamp 0
transform 1 0 4530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2505_
timestamp 0
transform 1 0 5070 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2506_
timestamp 0
transform -1 0 2510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2507_
timestamp 0
transform 1 0 3790 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2508_
timestamp 0
transform 1 0 3410 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2509_
timestamp 0
transform 1 0 4190 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2510_
timestamp 0
transform 1 0 3050 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2511_
timestamp 0
transform -1 0 4910 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2519_
timestamp 0
transform -1 0 5650 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2520_
timestamp 0
transform -1 0 7510 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2521_
timestamp 0
transform -1 0 7710 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2522_
timestamp 0
transform 1 0 7710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2523_
timestamp 0
transform 1 0 9450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2524_
timestamp 0
transform -1 0 7770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2525_
timestamp 0
transform 1 0 7510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2526_
timestamp 0
transform 1 0 8250 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2527_
timestamp 0
transform 1 0 8450 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2528_
timestamp 0
transform -1 0 9590 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2529_
timestamp 0
transform 1 0 8530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2530_
timestamp 0
transform -1 0 8170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2531_
timestamp 0
transform -1 0 8310 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2532_
timestamp 0
transform -1 0 8730 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2533_
timestamp 0
transform 1 0 9470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2534_
timestamp 0
transform 1 0 10030 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__2535_
timestamp 0
transform -1 0 10230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2536_
timestamp 0
transform -1 0 8730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2537_
timestamp 0
transform -1 0 8530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2538_
timestamp 0
transform -1 0 8330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2539_
timestamp 0
transform 1 0 7930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2540_
timestamp 0
transform -1 0 10630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2541_
timestamp 0
transform -1 0 10830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2542_
timestamp 0
transform 1 0 10870 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2543_
timestamp 0
transform -1 0 10570 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2544_
timestamp 0
transform -1 0 5670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2545_
timestamp 0
transform -1 0 5870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2546_
timestamp 0
transform -1 0 6090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2547_
timestamp 0
transform -1 0 5970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2548_
timestamp 0
transform -1 0 6170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2549_
timestamp 0
transform 1 0 5550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2550_
timestamp 0
transform 1 0 5750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2551_
timestamp 0
transform -1 0 6870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2552_
timestamp 0
transform -1 0 7230 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2553_
timestamp 0
transform -1 0 5690 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2554_
timestamp 0
transform -1 0 6330 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2555_
timestamp 0
transform 1 0 6370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2556_
timestamp 0
transform -1 0 6710 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2557_
timestamp 0
transform -1 0 6190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2558_
timestamp 0
transform 1 0 6470 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2559_
timestamp 0
transform 1 0 6850 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2560_
timestamp 0
transform -1 0 5890 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2561_
timestamp 0
transform -1 0 6530 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2562_
timestamp 0
transform 1 0 6710 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2563_
timestamp 0
transform -1 0 6090 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2564_
timestamp 0
transform 1 0 7750 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2565_
timestamp 0
transform 1 0 7970 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2566_
timestamp 0
transform 1 0 7550 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2567_
timestamp 0
transform 1 0 6950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2568_
timestamp 0
transform -1 0 6590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2569_
timestamp 0
transform 1 0 7170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2570_
timestamp 0
transform -1 0 9350 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2571_
timestamp 0
transform -1 0 9250 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2572_
timestamp 0
transform 1 0 9270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2573_
timestamp 0
transform 1 0 9150 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2574_
timestamp 0
transform -1 0 9230 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2575_
timestamp 0
transform -1 0 9050 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2576_
timestamp 0
transform -1 0 8770 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2577_
timestamp 0
transform -1 0 8970 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2578_
timestamp 0
transform 1 0 9530 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2579_
timestamp 0
transform -1 0 9470 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2580_
timestamp 0
transform -1 0 8270 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2581_
timestamp 0
transform 1 0 8230 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2582_
timestamp 0
transform 1 0 8350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2583_
timestamp 0
transform -1 0 9750 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2584_
timestamp 0
transform 1 0 9410 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2585_
timestamp 0
transform -1 0 11150 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2586_
timestamp 0
transform 1 0 8830 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2587_
timestamp 0
transform 1 0 8630 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2588_
timestamp 0
transform -1 0 8450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2589_
timestamp 0
transform 1 0 8490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2590_
timestamp 0
transform 1 0 8230 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2591_
timestamp 0
transform -1 0 8570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2592_
timestamp 0
transform 1 0 7830 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2593_
timestamp 0
transform -1 0 9070 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2594_
timestamp 0
transform -1 0 8970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2595_
timestamp 0
transform -1 0 9230 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2596_
timestamp 0
transform 1 0 10410 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2597_
timestamp 0
transform 1 0 10590 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2598_
timestamp 0
transform -1 0 10430 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2599_
timestamp 0
transform 1 0 10790 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2600_
timestamp 0
transform -1 0 11390 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2601_
timestamp 0
transform 1 0 8250 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2602_
timestamp 0
transform -1 0 8050 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2603_
timestamp 0
transform 1 0 7050 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2604_
timestamp 0
transform 1 0 8210 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2605_
timestamp 0
transform -1 0 8090 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2606_
timestamp 0
transform -1 0 7690 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2607_
timestamp 0
transform -1 0 6550 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2608_
timestamp 0
transform 1 0 6730 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2609_
timestamp 0
transform 1 0 6930 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2610_
timestamp 0
transform -1 0 7870 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2611_
timestamp 0
transform -1 0 10090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2612_
timestamp 0
transform 1 0 9870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2613_
timestamp 0
transform 1 0 10270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2614_
timestamp 0
transform -1 0 10970 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__2615_
timestamp 0
transform -1 0 7150 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2616_
timestamp 0
transform 1 0 8290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2617_
timestamp 0
transform -1 0 7150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2618_
timestamp 0
transform -1 0 6490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2619_
timestamp 0
transform 1 0 6270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2620_
timestamp 0
transform -1 0 7970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2621_
timestamp 0
transform -1 0 8070 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2622_
timestamp 0
transform 1 0 8330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2623_
timestamp 0
transform -1 0 8930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2624_
timestamp 0
transform 1 0 8070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2625_
timestamp 0
transform 1 0 6830 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2626_
timestamp 0
transform -1 0 8290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2627_
timestamp 0
transform 1 0 9890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2628_
timestamp 0
transform 1 0 11510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2629_
timestamp 0
transform 1 0 11410 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2630_
timestamp 0
transform 1 0 11690 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2631_
timestamp 0
transform -1 0 11510 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2632_
timestamp 0
transform 1 0 9410 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2633_
timestamp 0
transform -1 0 8510 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2634_
timestamp 0
transform 1 0 8910 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2635_
timestamp 0
transform -1 0 9150 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2636_
timestamp 0
transform -1 0 9930 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2637_
timestamp 0
transform -1 0 8630 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2638_
timestamp 0
transform 1 0 9710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2639_
timestamp 0
transform 1 0 9970 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2640_
timestamp 0
transform 1 0 8090 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2641_
timestamp 0
transform 1 0 7890 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2642_
timestamp 0
transform 1 0 9370 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2643_
timestamp 0
transform 1 0 9370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2644_
timestamp 0
transform 1 0 8390 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2645_
timestamp 0
transform 1 0 7610 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2646_
timestamp 0
transform 1 0 7410 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2647_
timestamp 0
transform 1 0 8190 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2648_
timestamp 0
transform -1 0 8030 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2649_
timestamp 0
transform -1 0 9030 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2650_
timestamp 0
transform 1 0 11090 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2651_
timestamp 0
transform -1 0 9230 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2652_
timestamp 0
transform -1 0 8530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2653_
timestamp 0
transform 1 0 8710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2654_
timestamp 0
transform 1 0 5830 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2655_
timestamp 0
transform -1 0 6050 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2656_
timestamp 0
transform -1 0 6230 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2657_
timestamp 0
transform -1 0 7630 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2658_
timestamp 0
transform 1 0 7390 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2659_
timestamp 0
transform -1 0 7150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2660_
timestamp 0
transform -1 0 7330 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2661_
timestamp 0
transform -1 0 10770 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2662_
timestamp 0
transform 1 0 10950 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2663_
timestamp 0
transform 1 0 10010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2664_
timestamp 0
transform 1 0 10190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2665_
timestamp 0
transform -1 0 6610 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2666_
timestamp 0
transform 1 0 7190 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2667_
timestamp 0
transform -1 0 6990 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2668_
timestamp 0
transform -1 0 6810 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2669_
timestamp 0
transform 1 0 6730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2670_
timestamp 0
transform -1 0 10590 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2671_
timestamp 0
transform 1 0 11650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2672_
timestamp 0
transform 1 0 11690 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2673_
timestamp 0
transform -1 0 11490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2674_
timestamp 0
transform 1 0 11430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2675_
timestamp 0
transform -1 0 10790 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2676_
timestamp 0
transform 1 0 11410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2677_
timestamp 0
transform -1 0 11490 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2678_
timestamp 0
transform -1 0 10110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2679_
timestamp 0
transform 1 0 9710 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2680_
timestamp 0
transform 1 0 9630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2681_
timestamp 0
transform 1 0 9310 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2682_
timestamp 0
transform -1 0 9530 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2683_
timestamp 0
transform -1 0 10190 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2684_
timestamp 0
transform -1 0 10490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2685_
timestamp 0
transform -1 0 10770 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__2686_
timestamp 0
transform 1 0 10670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2687_
timestamp 0
transform -1 0 9790 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2688_
timestamp 0
transform 1 0 9190 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2689_
timestamp 0
transform 1 0 10510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2690_
timestamp 0
transform -1 0 10870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2691_
timestamp 0
transform -1 0 11070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2692_
timestamp 0
transform 1 0 11250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2693_
timestamp 0
transform -1 0 10410 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2694_
timestamp 0
transform 1 0 9610 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2695_
timestamp 0
transform -1 0 10530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2696_
timestamp 0
transform 1 0 10290 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2697_
timestamp 0
transform 1 0 9950 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2698_
timestamp 0
transform 1 0 9930 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2699_
timestamp 0
transform 1 0 9050 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2700_
timestamp 0
transform 1 0 8830 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2701_
timestamp 0
transform -1 0 8470 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2702_
timestamp 0
transform 1 0 8830 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2703_
timestamp 0
transform 1 0 10850 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2704_
timestamp 0
transform -1 0 9110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2705_
timestamp 0
transform -1 0 9670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2706_
timestamp 0
transform -1 0 10070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2707_
timestamp 0
transform -1 0 9590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2708_
timestamp 0
transform 1 0 8890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2709_
timestamp 0
transform 1 0 9010 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2710_
timestamp 0
transform -1 0 8710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2711_
timestamp 0
transform -1 0 10770 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2712_
timestamp 0
transform -1 0 10750 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2713_
timestamp 0
transform 1 0 10790 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2714_
timestamp 0
transform 1 0 10790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2715_
timestamp 0
transform -1 0 11430 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2716_
timestamp 0
transform 1 0 11590 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2717_
timestamp 0
transform -1 0 10710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2718_
timestamp 0
transform 1 0 11050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2719_
timestamp 0
transform 1 0 11770 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2720_
timestamp 0
transform -1 0 10970 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2721_
timestamp 0
transform -1 0 10870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2722_
timestamp 0
transform -1 0 10910 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2723_
timestamp 0
transform 1 0 11350 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2724_
timestamp 0
transform 1 0 11330 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2725_
timestamp 0
transform 1 0 10310 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2726_
timestamp 0
transform -1 0 9690 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2727_
timestamp 0
transform 1 0 9890 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2728_
timestamp 0
transform -1 0 9870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2729_
timestamp 0
transform -1 0 9470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2730_
timestamp 0
transform 1 0 11210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2731_
timestamp 0
transform 1 0 9450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2732_
timestamp 0
transform 1 0 6670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2733_
timestamp 0
transform -1 0 9090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2734_
timestamp 0
transform 1 0 9450 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2735_
timestamp 0
transform 1 0 9470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2736_
timestamp 0
transform -1 0 8890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2737_
timestamp 0
transform -1 0 9270 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2738_
timestamp 0
transform -1 0 10350 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2739_
timestamp 0
transform 1 0 10530 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2740_
timestamp 0
transform 1 0 11150 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2741_
timestamp 0
transform 1 0 11550 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2742_
timestamp 0
transform -1 0 10550 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2743_
timestamp 0
transform -1 0 10390 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2744_
timestamp 0
transform 1 0 10470 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2745_
timestamp 0
transform -1 0 11130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2746_
timestamp 0
transform -1 0 10130 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2747_
timestamp 0
transform 1 0 10930 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2748_
timestamp 0
transform 1 0 9790 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2749_
timestamp 0
transform 1 0 10650 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2750_
timestamp 0
transform 1 0 10990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2751_
timestamp 0
transform -1 0 10110 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2752_
timestamp 0
transform 1 0 5730 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2753_
timestamp 0
transform -1 0 5950 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2754_
timestamp 0
transform -1 0 6010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2755_
timestamp 0
transform -1 0 7370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2756_
timestamp 0
transform -1 0 7490 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2757_
timestamp 0
transform 1 0 8090 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2758_
timestamp 0
transform -1 0 7550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2759_
timestamp 0
transform -1 0 9690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2760_
timestamp 0
transform -1 0 6210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2761_
timestamp 0
transform -1 0 8850 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2762_
timestamp 0
transform -1 0 8830 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2763_
timestamp 0
transform -1 0 6290 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2764_
timestamp 0
transform -1 0 6370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2765_
timestamp 0
transform -1 0 9330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2766_
timestamp 0
transform -1 0 6670 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2767_
timestamp 0
transform 1 0 8890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2768_
timestamp 0
transform -1 0 5970 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2769_
timestamp 0
transform -1 0 6910 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2770_
timestamp 0
transform 1 0 7090 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2771_
timestamp 0
transform 1 0 10010 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2772_
timestamp 0
transform -1 0 7370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2773_
timestamp 0
transform -1 0 7570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2774_
timestamp 0
transform -1 0 6010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2775_
timestamp 0
transform -1 0 7310 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2776_
timestamp 0
transform 1 0 6130 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2777_
timestamp 0
transform -1 0 9850 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2778_
timestamp 0
transform 1 0 7670 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2779_
timestamp 0
transform 1 0 7890 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2780_
timestamp 0
transform 1 0 7950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2781_
timestamp 0
transform -1 0 7770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2782_
timestamp 0
transform 1 0 7630 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2783_
timestamp 0
transform -1 0 8430 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2784_
timestamp 0
transform -1 0 10970 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2785_
timestamp 0
transform 1 0 9490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2786_
timestamp 0
transform -1 0 7750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2787_
timestamp 0
transform -1 0 9190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2788_
timestamp 0
transform -1 0 10170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2789_
timestamp 0
transform 1 0 10350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2790_
timestamp 0
transform 1 0 7950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2791_
timestamp 0
transform 1 0 8150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2792_
timestamp 0
transform -1 0 7610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2793_
timestamp 0
transform -1 0 7830 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2794_
timestamp 0
transform -1 0 7830 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2795_
timestamp 0
transform -1 0 7550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2796_
timestamp 0
transform -1 0 6950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2797_
timestamp 0
transform -1 0 8370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2798_
timestamp 0
transform 1 0 11910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2799_
timestamp 0
transform -1 0 7330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2800_
timestamp 0
transform -1 0 7450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2801_
timestamp 0
transform 1 0 7090 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2802_
timestamp 0
transform 1 0 6750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2803_
timestamp 0
transform -1 0 6970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2804_
timestamp 0
transform -1 0 8470 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2805_
timestamp 0
transform 1 0 6890 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2806_
timestamp 0
transform -1 0 6790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2807_
timestamp 0
transform -1 0 7050 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2808_
timestamp 0
transform 1 0 10130 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2809_
timestamp 0
transform -1 0 10550 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2810_
timestamp 0
transform 1 0 10530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2811_
timestamp 0
transform 1 0 10350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2812_
timestamp 0
transform 1 0 10210 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2813_
timestamp 0
transform -1 0 10050 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2814_
timestamp 0
transform -1 0 10450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2815_
timestamp 0
transform -1 0 10650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2816_
timestamp 0
transform 1 0 10170 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2817_
timestamp 0
transform -1 0 10270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2818_
timestamp 0
transform -1 0 10930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2819_
timestamp 0
transform -1 0 11030 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2820_
timestamp 0
transform -1 0 11230 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2821_
timestamp 0
transform 1 0 10990 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2822_
timestamp 0
transform -1 0 11930 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2823_
timestamp 0
transform 1 0 11110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2824_
timestamp 0
transform 1 0 10610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2825_
timestamp 0
transform 1 0 11130 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2826_
timestamp 0
transform 1 0 11330 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2827_
timestamp 0
transform -1 0 11790 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2828_
timestamp 0
transform -1 0 11910 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2829_
timestamp 0
transform -1 0 11350 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2830_
timestamp 0
transform 1 0 10990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2831_
timestamp 0
transform 1 0 11050 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2832_
timestamp 0
transform -1 0 11290 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2833_
timestamp 0
transform 1 0 11350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2834_
timestamp 0
transform 1 0 11850 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2835_
timestamp 0
transform 1 0 12030 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__2836_
timestamp 0
transform 1 0 11650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2837_
timestamp 0
transform 1 0 11850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2838_
timestamp 0
transform 1 0 11970 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2839_
timestamp 0
transform 1 0 11550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2840_
timestamp 0
transform -1 0 11750 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2841_
timestamp 0
transform -1 0 11610 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2842_
timestamp 0
transform -1 0 9790 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2843_
timestamp 0
transform -1 0 9990 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2844_
timestamp 0
transform -1 0 11770 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2845_
timestamp 0
transform 1 0 11950 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2846_
timestamp 0
transform 1 0 11510 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__2847_
timestamp 0
transform 1 0 11930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2848_
timestamp 0
transform -1 0 11570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2849_
timestamp 0
transform -1 0 11670 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2850_
timestamp 0
transform 1 0 11850 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2851_
timestamp 0
transform -1 0 9850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2852_
timestamp 0
transform -1 0 11030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2853_
timestamp 0
transform 1 0 11210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2854_
timestamp 0
transform 1 0 11790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2855_
timestamp 0
transform 1 0 11790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2856_
timestamp 0
transform -1 0 9810 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2857_
timestamp 0
transform -1 0 9870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2858_
timestamp 0
transform -1 0 8030 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2859_
timestamp 0
transform 1 0 9650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2860_
timestamp 0
transform -1 0 9110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2861_
timestamp 0
transform 1 0 9930 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2862_
timestamp 0
transform 1 0 9530 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2863_
timestamp 0
transform 1 0 8750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2864_
timestamp 0
transform -1 0 7750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2865_
timestamp 0
transform -1 0 6410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2866_
timestamp 0
transform -1 0 8830 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2867_
timestamp 0
transform -1 0 9370 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2868_
timestamp 0
transform 1 0 9170 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2869_
timestamp 0
transform -1 0 10530 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2870_
timestamp 0
transform -1 0 9290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2871_
timestamp 0
transform -1 0 8530 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2872_
timestamp 0
transform 1 0 9730 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2873_
timestamp 0
transform 1 0 9770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2874_
timestamp 0
transform 1 0 9570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2875_
timestamp 0
transform -1 0 11170 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__2876_
timestamp 0
transform 1 0 10170 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2877_
timestamp 0
transform -1 0 10710 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2878_
timestamp 0
transform 1 0 9610 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2879_
timestamp 0
transform -1 0 9830 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2880_
timestamp 0
transform -1 0 10150 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2881_
timestamp 0
transform -1 0 5930 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2882_
timestamp 0
transform -1 0 6110 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2883_
timestamp 0
transform -1 0 5470 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2884_
timestamp 0
transform -1 0 5470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2885_
timestamp 0
transform 1 0 5450 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2886_
timestamp 0
transform -1 0 5270 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__2887_
timestamp 0
transform 1 0 5610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2888_
timestamp 0
transform 1 0 6030 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2889_
timestamp 0
transform -1 0 6270 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2890_
timestamp 0
transform -1 0 6650 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2891_
timestamp 0
transform 1 0 8130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2892_
timestamp 0
transform -1 0 7250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2893_
timestamp 0
transform -1 0 5850 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2894_
timestamp 0
transform 1 0 5350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2895_
timestamp 0
transform -1 0 7450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2896_
timestamp 0
transform -1 0 6570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__2897_
timestamp 0
transform 1 0 7310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2898_
timestamp 0
transform 1 0 11730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2899_
timestamp 0
transform -1 0 6510 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2900_
timestamp 0
transform -1 0 6710 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2901_
timestamp 0
transform -1 0 8150 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2902_
timestamp 0
transform 1 0 9610 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2903_
timestamp 0
transform -1 0 11550 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2904_
timestamp 0
transform 1 0 8330 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2905_
timestamp 0
transform -1 0 6910 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2906_
timestamp 0
transform -1 0 7290 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2907_
timestamp 0
transform -1 0 6310 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2908_
timestamp 0
transform 1 0 8430 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2909_
timestamp 0
transform -1 0 10330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2910_
timestamp 0
transform 1 0 10730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2911_
timestamp 0
transform 1 0 10910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2912_
timestamp 0
transform -1 0 10770 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2913_
timestamp 0
transform -1 0 8650 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2914_
timestamp 0
transform -1 0 8530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2915_
timestamp 0
transform -1 0 11210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2916_
timestamp 0
transform -1 0 7950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2917_
timestamp 0
transform -1 0 6970 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2918_
timestamp 0
transform 1 0 6750 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2919_
timestamp 0
transform -1 0 7170 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2920_
timestamp 0
transform 1 0 7130 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2921_
timestamp 0
transform 1 0 6930 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2922_
timestamp 0
transform 1 0 6590 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2923_
timestamp 0
transform -1 0 5810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2924_
timestamp 0
transform 1 0 8850 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2925_
timestamp 0
transform 1 0 10210 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2926_
timestamp 0
transform 1 0 11950 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2927_
timestamp 0
transform 1 0 8670 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2928_
timestamp 0
transform 1 0 7470 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2929_
timestamp 0
transform 1 0 8190 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2930_
timestamp 0
transform -1 0 8410 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2931_
timestamp 0
transform -1 0 8050 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2932_
timestamp 0
transform 1 0 7850 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2933_
timestamp 0
transform 1 0 7890 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2934_
timestamp 0
transform -1 0 10190 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2935_
timestamp 0
transform 1 0 11310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__2936_
timestamp 0
transform -1 0 8170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2937_
timestamp 0
transform 1 0 8650 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2938_
timestamp 0
transform -1 0 11770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2939_
timestamp 0
transform -1 0 11210 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2940_
timestamp 0
transform -1 0 6550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2941_
timestamp 0
transform 1 0 8830 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2942_
timestamp 0
transform 1 0 8910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2943_
timestamp 0
transform 1 0 9670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2944_
timestamp 0
transform 1 0 9850 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__2945_
timestamp 0
transform 1 0 9030 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2946_
timestamp 0
transform -1 0 9130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2947_
timestamp 0
transform -1 0 8690 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2948_
timestamp 0
transform -1 0 8630 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2949_
timestamp 0
transform 1 0 10810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2950_
timestamp 0
transform 1 0 11630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2951_
timestamp 0
transform -1 0 6950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2952_
timestamp 0
transform -1 0 6750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2953_
timestamp 0
transform 1 0 11250 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2954_
timestamp 0
transform -1 0 8930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2955_
timestamp 0
transform -1 0 10070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__2956_
timestamp 0
transform -1 0 11330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2957_
timestamp 0
transform 1 0 9650 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2958_
timestamp 0
transform 1 0 11610 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__2959_
timestamp 0
transform 1 0 5090 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2960_
timestamp 0
transform -1 0 7350 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2961_
timestamp 0
transform -1 0 7950 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2962_
timestamp 0
transform -1 0 7550 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2963_
timestamp 0
transform -1 0 6470 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__2964_
timestamp 0
transform -1 0 7750 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2965_
timestamp 0
transform -1 0 11730 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__2966_
timestamp 0
transform 1 0 8550 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2967_
timestamp 0
transform 1 0 9250 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__2968_
timestamp 0
transform 1 0 10370 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2969_
timestamp 0
transform 1 0 10570 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__2970_
timestamp 0
transform -1 0 11250 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2971_
timestamp 0
transform 1 0 7710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2972_
timestamp 0
transform -1 0 9310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2973_
timestamp 0
transform 1 0 7350 0 1 250
box -6 -8 26 248
use FILL  FILL_1__2974_
timestamp 0
transform -1 0 7290 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2975_
timestamp 0
transform -1 0 9050 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__2976_
timestamp 0
transform 1 0 10030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2977_
timestamp 0
transform 1 0 10430 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2978_
timestamp 0
transform -1 0 11590 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__2979_
timestamp 0
transform -1 0 11830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__2980_
timestamp 0
transform 1 0 7150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2981_
timestamp 0
transform 1 0 6550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__2982_
timestamp 0
transform 1 0 7490 0 1 730
box -6 -8 26 248
use FILL  FILL_1__2983_
timestamp 0
transform 1 0 11870 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__2984_
timestamp 0
transform 1 0 11610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__2985_
timestamp 0
transform -1 0 7110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__2986_
timestamp 0
transform -1 0 7130 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__2987_
timestamp 0
transform 1 0 5790 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__3000_
timestamp 0
transform -1 0 2190 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3001_
timestamp 0
transform 1 0 2330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3002_
timestamp 0
transform 1 0 2130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__3003_
timestamp 0
transform -1 0 3610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__3004_
timestamp 0
transform 1 0 3810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__3005_
timestamp 0
transform -1 0 3450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__3006_
timestamp 0
transform -1 0 4330 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__3007_
timestamp 0
transform -1 0 4130 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__3008_
timestamp 0
transform 1 0 3850 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__3009_
timestamp 0
transform 1 0 3950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3010_
timestamp 0
transform -1 0 3970 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__3011_
timestamp 0
transform 1 0 3770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3012_
timestamp 0
transform 1 0 2710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__3013_
timestamp 0
transform -1 0 2410 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3014_
timestamp 0
transform 1 0 2550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__3015_
timestamp 0
transform -1 0 4530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3016_
timestamp 0
transform 1 0 4450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__3017_
timestamp 0
transform 1 0 4150 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3018_
timestamp 0
transform 1 0 4350 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3019_
timestamp 0
transform -1 0 3970 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3020_
timestamp 0
transform 1 0 1790 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3021_
timestamp 0
transform 1 0 1630 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3022_
timestamp 0
transform -1 0 2030 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3023_
timestamp 0
transform -1 0 2870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3024_
timestamp 0
transform 1 0 4690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3025_
timestamp 0
transform 1 0 4310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3026_
timestamp 0
transform 1 0 3570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3027_
timestamp 0
transform 1 0 3270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__3028_
timestamp 0
transform -1 0 2770 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__3029_
timestamp 0
transform 1 0 3410 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3030_
timestamp 0
transform 1 0 4850 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__3031_
timestamp 0
transform 1 0 4690 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__3032_
timestamp 0
transform 1 0 5850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3033_
timestamp 0
transform -1 0 4570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3034_
timestamp 0
transform 1 0 3790 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3035_
timestamp 0
transform -1 0 4550 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__3036_
timestamp 0
transform -1 0 2350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__3037_
timestamp 0
transform -1 0 3290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__3038_
timestamp 0
transform 1 0 2170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__3039_
timestamp 0
transform -1 0 3550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3040_
timestamp 0
transform -1 0 3770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3041_
timestamp 0
transform 1 0 3370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3042_
timestamp 0
transform -1 0 2750 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3043_
timestamp 0
transform -1 0 3790 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__3044_
timestamp 0
transform -1 0 2590 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3045_
timestamp 0
transform -1 0 2890 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__3046_
timestamp 0
transform -1 0 3230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3047_
timestamp 0
transform 1 0 2830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3048_
timestamp 0
transform 1 0 3370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__3049_
timestamp 0
transform -1 0 3670 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__3050_
timestamp 0
transform -1 0 2910 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__3051_
timestamp 0
transform -1 0 2930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__3052_
timestamp 0
transform 1 0 3090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__3053_
timestamp 0
transform -1 0 2970 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3054_
timestamp 0
transform -1 0 2570 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__3055_
timestamp 0
transform -1 0 2390 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__3056_
timestamp 0
transform -1 0 2710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3057_
timestamp 0
transform -1 0 3230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3058_
timestamp 0
transform 1 0 4150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3059_
timestamp 0
transform -1 0 5070 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__3060_
timestamp 0
transform -1 0 5270 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__3061_
timestamp 0
transform -1 0 6030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3062_
timestamp 0
transform -1 0 5090 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__3063_
timestamp 0
transform -1 0 5110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__3064_
timestamp 0
transform -1 0 4950 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3076_
timestamp 0
transform 1 0 1050 0 1 250
box -6 -8 26 248
use FILL  FILL_1__3077_
timestamp 0
transform -1 0 1270 0 1 250
box -6 -8 26 248
use FILL  FILL_1__3078_
timestamp 0
transform 1 0 890 0 1 250
box -6 -8 26 248
use FILL  FILL_1__3079_
timestamp 0
transform 1 0 970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__3080_
timestamp 0
transform -1 0 850 0 1 730
box -6 -8 26 248
use FILL  FILL_1__3081_
timestamp 0
transform 1 0 790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__3082_
timestamp 0
transform 1 0 1370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__3083_
timestamp 0
transform -1 0 1530 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__3084_
timestamp 0
transform 1 0 1450 0 1 250
box -6 -8 26 248
use FILL  FILL_1__3085_
timestamp 0
transform -1 0 1730 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__3086_
timestamp 0
transform -1 0 430 0 1 730
box -6 -8 26 248
use FILL  FILL_1__3087_
timestamp 0
transform -1 0 610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__3088_
timestamp 0
transform 1 0 410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__3089_
timestamp 0
transform -1 0 1390 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__3090_
timestamp 0
transform 1 0 1190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3091_
timestamp 0
transform -1 0 1870 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__3092_
timestamp 0
transform -1 0 650 0 1 730
box -6 -8 26 248
use FILL  FILL_1__3093_
timestamp 0
transform -1 0 50 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__3094_
timestamp 0
transform -1 0 50 0 1 730
box -6 -8 26 248
use FILL  FILL_1__3095_
timestamp 0
transform -1 0 250 0 1 730
box -6 -8 26 248
use FILL  FILL_1__3096_
timestamp 0
transform -1 0 250 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__3097_
timestamp 0
transform 1 0 2010 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__3098_
timestamp 0
transform -1 0 2310 0 1 250
box -6 -8 26 248
use FILL  FILL_1__3099_
timestamp 0
transform 1 0 1870 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__3100_
timestamp 0
transform 1 0 30 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3101_
timestamp 0
transform -1 0 50 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__3102_
timestamp 0
transform -1 0 1230 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__3103_
timestamp 0
transform -1 0 1190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__3104_
timestamp 0
transform -1 0 230 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__3105_
timestamp 0
transform -1 0 1150 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__3106_
timestamp 0
transform -1 0 2310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__3107_
timestamp 0
transform -1 0 1510 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__3108_
timestamp 0
transform -1 0 390 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3109_
timestamp 0
transform -1 0 570 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3110_
timestamp 0
transform 1 0 710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__3111_
timestamp 0
transform -1 0 910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__3112_
timestamp 0
transform -1 0 50 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__3113_
timestamp 0
transform -1 0 50 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3114_
timestamp 0
transform -1 0 4550 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__3115_
timestamp 0
transform -1 0 4610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3116_
timestamp 0
transform 1 0 4470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__3117_
timestamp 0
transform 1 0 510 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__3118_
timestamp 0
transform -1 0 1670 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__3119_
timestamp 0
transform 1 0 850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3120_
timestamp 0
transform 1 0 1010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3121_
timestamp 0
transform -1 0 2330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3122_
timestamp 0
transform -1 0 430 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__3123_
timestamp 0
transform 1 0 310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__3124_
timestamp 0
transform 1 0 210 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__3125_
timestamp 0
transform 1 0 2030 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__3126_
timestamp 0
transform -1 0 2250 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__3127_
timestamp 0
transform 1 0 1550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3128_
timestamp 0
transform 1 0 1390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3129_
timestamp 0
transform 1 0 4730 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__3130_
timestamp 0
transform 1 0 4910 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__3131_
timestamp 0
transform 1 0 5130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__3132_
timestamp 0
transform 1 0 4790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3133_
timestamp 0
transform -1 0 4690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__3134_
timestamp 0
transform -1 0 4330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__3135_
timestamp 0
transform 1 0 690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__3136_
timestamp 0
transform -1 0 750 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__3137_
timestamp 0
transform 1 0 350 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__3138_
timestamp 0
transform 1 0 690 0 1 250
box -6 -8 26 248
use FILL  FILL_1__3139_
timestamp 0
transform 1 0 210 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__3140_
timestamp 0
transform -1 0 1510 0 1 730
box -6 -8 26 248
use FILL  FILL_1__3141_
timestamp 0
transform 1 0 1690 0 1 730
box -6 -8 26 248
use FILL  FILL_1__3142_
timestamp 0
transform -1 0 1670 0 1 250
box -6 -8 26 248
use FILL  FILL_1__3143_
timestamp 0
transform 1 0 2370 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__3144_
timestamp 0
transform 1 0 2490 0 1 250
box -6 -8 26 248
use FILL  FILL_1__3145_
timestamp 0
transform 1 0 2210 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__3146_
timestamp 0
transform -1 0 1910 0 1 730
box -6 -8 26 248
use FILL  FILL_1__3147_
timestamp 0
transform 1 0 2010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__3148_
timestamp 0
transform 1 0 1050 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__3149_
timestamp 0
transform -1 0 890 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__3150_
timestamp 0
transform -1 0 250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__3151_
timestamp 0
transform 1 0 30 0 1 250
box -6 -8 26 248
use FILL  FILL_1__3152_
timestamp 0
transform -1 0 2110 0 1 730
box -6 -8 26 248
use FILL  FILL_1__3284_
timestamp 0
transform -1 0 4710 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__3285_
timestamp 0
transform 1 0 4350 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__3286_
timestamp 0
transform -1 0 3390 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3287_
timestamp 0
transform 1 0 3250 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3288_
timestamp 0
transform 1 0 2170 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3289_
timestamp 0
transform 1 0 2370 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3290_
timestamp 0
transform -1 0 2050 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3291_
timestamp 0
transform 1 0 2990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3292_
timestamp 0
transform 1 0 3190 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3293_
timestamp 0
transform 1 0 5810 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3294_
timestamp 0
transform -1 0 5850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3295_
timestamp 0
transform 1 0 5890 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3296_
timestamp 0
transform 1 0 6370 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3297_
timestamp 0
transform 1 0 6570 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3298_
timestamp 0
transform 1 0 5270 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3299_
timestamp 0
transform 1 0 5470 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3300_
timestamp 0
transform 1 0 4610 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3301_
timestamp 0
transform 1 0 4810 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3302_
timestamp 0
transform -1 0 3370 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3303_
timestamp 0
transform -1 0 3530 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3304_
timestamp 0
transform -1 0 3410 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3305_
timestamp 0
transform -1 0 3590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3306_
timestamp 0
transform 1 0 4330 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3307_
timestamp 0
transform 1 0 4430 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3308_
timestamp 0
transform -1 0 1090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3309_
timestamp 0
transform -1 0 1010 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__3310_
timestamp 0
transform 1 0 2490 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3311_
timestamp 0
transform -1 0 2710 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3312_
timestamp 0
transform 1 0 3430 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3313_
timestamp 0
transform -1 0 2350 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3314_
timestamp 0
transform -1 0 230 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__3315_
timestamp 0
transform -1 0 430 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__3316_
timestamp 0
transform -1 0 7510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__3317_
timestamp 0
transform 1 0 6130 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3318_
timestamp 0
transform 1 0 2610 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3319_
timestamp 0
transform 1 0 6630 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3320_
timestamp 0
transform 1 0 5410 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3321_
timestamp 0
transform -1 0 6430 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__3322_
timestamp 0
transform -1 0 3790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3323_
timestamp 0
transform -1 0 3630 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3324_
timestamp 0
transform 1 0 5130 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3325_
timestamp 0
transform -1 0 5350 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3326_
timestamp 0
transform -1 0 5210 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__3327_
timestamp 0
transform 1 0 4790 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__3328_
timestamp 0
transform -1 0 5250 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3329_
timestamp 0
transform -1 0 5670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__3330_
timestamp 0
transform 1 0 5530 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3331_
timestamp 0
transform 1 0 4950 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3332_
timestamp 0
transform -1 0 4630 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__3333_
timestamp 0
transform -1 0 5930 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3334_
timestamp 0
transform 1 0 5910 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__3335_
timestamp 0
transform -1 0 430 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3336_
timestamp 0
transform -1 0 250 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3337_
timestamp 0
transform -1 0 870 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3338_
timestamp 0
transform -1 0 890 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3339_
timestamp 0
transform -1 0 5850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__3340_
timestamp 0
transform 1 0 6030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__3341_
timestamp 0
transform -1 0 5810 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3342_
timestamp 0
transform -1 0 5430 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3343_
timestamp 0
transform -1 0 4350 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3344_
timestamp 0
transform -1 0 5470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__3345_
timestamp 0
transform 1 0 5650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__3346_
timestamp 0
transform 1 0 5250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__3347_
timestamp 0
transform 1 0 5070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__3348_
timestamp 0
transform -1 0 50 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3349_
timestamp 0
transform 1 0 230 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3350_
timestamp 0
transform 1 0 7750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__3351_
timestamp 0
transform -1 0 50 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3352_
timestamp 0
transform 1 0 270 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3353_
timestamp 0
transform -1 0 1790 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3354_
timestamp 0
transform 1 0 1970 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3355_
timestamp 0
transform -1 0 290 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3356_
timestamp 0
transform -1 0 490 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3357_
timestamp 0
transform -1 0 830 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3358_
timestamp 0
transform -1 0 810 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3359_
timestamp 0
transform -1 0 50 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3360_
timestamp 0
transform -1 0 250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__3361_
timestamp 0
transform -1 0 4850 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3362_
timestamp 0
transform -1 0 4970 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3363_
timestamp 0
transform 1 0 5290 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3364_
timestamp 0
transform -1 0 3390 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3365_
timestamp 0
transform 1 0 3310 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3366_
timestamp 0
transform 1 0 2890 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3367_
timestamp 0
transform 1 0 2530 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3368_
timestamp 0
transform 1 0 2330 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3369_
timestamp 0
transform -1 0 4110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3370_
timestamp 0
transform -1 0 5270 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3371_
timestamp 0
transform -1 0 7030 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3372_
timestamp 0
transform 1 0 5070 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3373_
timestamp 0
transform -1 0 7470 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3374_
timestamp 0
transform -1 0 7250 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3375_
timestamp 0
transform -1 0 4650 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3376_
timestamp 0
transform -1 0 4690 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3377_
timestamp 0
transform 1 0 4870 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3378_
timestamp 0
transform -1 0 4290 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3379_
timestamp 0
transform 1 0 5730 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3380_
timestamp 0
transform -1 0 7790 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3381_
timestamp 0
transform 1 0 6630 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3382_
timestamp 0
transform 1 0 6450 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3383_
timestamp 0
transform -1 0 7050 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3384_
timestamp 0
transform -1 0 6850 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3385_
timestamp 0
transform 1 0 7230 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3386_
timestamp 0
transform -1 0 6490 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3387_
timestamp 0
transform 1 0 6270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3388_
timestamp 0
transform 1 0 6690 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3389_
timestamp 0
transform -1 0 7090 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3390_
timestamp 0
transform -1 0 9690 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3391_
timestamp 0
transform -1 0 10230 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3392_
timestamp 0
transform -1 0 230 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3393_
timestamp 0
transform 1 0 210 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3394_
timestamp 0
transform -1 0 210 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3395_
timestamp 0
transform -1 0 230 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3396_
timestamp 0
transform -1 0 50 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3397_
timestamp 0
transform -1 0 1210 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3398_
timestamp 0
transform 1 0 990 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3399_
timestamp 0
transform 1 0 950 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3400_
timestamp 0
transform -1 0 590 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3401_
timestamp 0
transform -1 0 50 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3402_
timestamp 0
transform -1 0 810 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3403_
timestamp 0
transform 1 0 1570 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3404_
timestamp 0
transform -1 0 870 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3405_
timestamp 0
transform 1 0 670 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3406_
timestamp 0
transform -1 0 1850 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3407_
timestamp 0
transform -1 0 450 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__3408_
timestamp 0
transform 1 0 230 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__3409_
timestamp 0
transform -1 0 50 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__3410_
timestamp 0
transform -1 0 870 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3411_
timestamp 0
transform -1 0 410 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3412_
timestamp 0
transform -1 0 230 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3413_
timestamp 0
transform -1 0 50 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3414_
timestamp 0
transform -1 0 210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3415_
timestamp 0
transform -1 0 50 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3416_
timestamp 0
transform -1 0 50 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3417_
timestamp 0
transform -1 0 390 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3418_
timestamp 0
transform -1 0 6910 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3419_
timestamp 0
transform 1 0 6210 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3420_
timestamp 0
transform 1 0 6010 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3421_
timestamp 0
transform 1 0 5250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3422_
timestamp 0
transform 1 0 5110 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3423_
timestamp 0
transform 1 0 7090 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3424_
timestamp 0
transform -1 0 1350 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3425_
timestamp 0
transform 1 0 590 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3426_
timestamp 0
transform 1 0 390 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3427_
timestamp 0
transform -1 0 410 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3428_
timestamp 0
transform -1 0 250 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3429_
timestamp 0
transform 1 0 570 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3430_
timestamp 0
transform -1 0 50 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3431_
timestamp 0
transform -1 0 230 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3432_
timestamp 0
transform 1 0 850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3433_
timestamp 0
transform 1 0 1450 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3434_
timestamp 0
transform -1 0 950 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3435_
timestamp 0
transform -1 0 1070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3436_
timestamp 0
transform 1 0 1250 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3437_
timestamp 0
transform -1 0 1290 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__3438_
timestamp 0
transform -1 0 970 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3439_
timestamp 0
transform -1 0 770 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3440_
timestamp 0
transform -1 0 1090 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__3441_
timestamp 0
transform 1 0 690 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3442_
timestamp 0
transform 1 0 790 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3443_
timestamp 0
transform -1 0 770 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3444_
timestamp 0
transform -1 0 590 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3445_
timestamp 0
transform -1 0 710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__3446_
timestamp 0
transform -1 0 1370 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3447_
timestamp 0
transform -1 0 1150 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3448_
timestamp 0
transform -1 0 690 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3449_
timestamp 0
transform 1 0 1310 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3450_
timestamp 0
transform 1 0 1490 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3451_
timestamp 0
transform -1 0 2610 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3452_
timestamp 0
transform -1 0 2810 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3453_
timestamp 0
transform -1 0 3030 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3454_
timestamp 0
transform -1 0 1150 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__3455_
timestamp 0
transform -1 0 250 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3456_
timestamp 0
transform -1 0 50 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3457_
timestamp 0
transform -1 0 810 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3458_
timestamp 0
transform 1 0 590 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3459_
timestamp 0
transform -1 0 530 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__3460_
timestamp 0
transform 1 0 430 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3461_
timestamp 0
transform -1 0 1870 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3462_
timestamp 0
transform 1 0 1650 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3463_
timestamp 0
transform -1 0 1910 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__3464_
timestamp 0
transform -1 0 2030 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3465_
timestamp 0
transform -1 0 1610 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3466_
timestamp 0
transform -1 0 1990 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__3467_
timestamp 0
transform -1 0 1850 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3468_
timestamp 0
transform -1 0 2250 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3469_
timestamp 0
transform -1 0 250 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3470_
timestamp 0
transform -1 0 1190 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3471_
timestamp 0
transform -1 0 1170 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3472_
timestamp 0
transform -1 0 1550 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3473_
timestamp 0
transform 1 0 1730 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3474_
timestamp 0
transform -1 0 2030 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3475_
timestamp 0
transform -1 0 1710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3476_
timestamp 0
transform -1 0 1670 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3477_
timestamp 0
transform -1 0 1850 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3478_
timestamp 0
transform 1 0 1930 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3479_
timestamp 0
transform -1 0 1390 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3480_
timestamp 0
transform -1 0 2790 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3481_
timestamp 0
transform -1 0 6030 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3482_
timestamp 0
transform -1 0 5850 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3483_
timestamp 0
transform 1 0 6690 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3484_
timestamp 0
transform -1 0 7450 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__3485_
timestamp 0
transform -1 0 7250 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__3486_
timestamp 0
transform 1 0 5710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__3487_
timestamp 0
transform -1 0 5730 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3488_
timestamp 0
transform 1 0 2950 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3489_
timestamp 0
transform -1 0 6090 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__3490_
timestamp 0
transform 1 0 1510 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3491_
timestamp 0
transform 1 0 1330 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3492_
timestamp 0
transform 1 0 1890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3493_
timestamp 0
transform -1 0 1730 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3494_
timestamp 0
transform 1 0 7170 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3495_
timestamp 0
transform -1 0 7550 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3496_
timestamp 0
transform -1 0 7750 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3497_
timestamp 0
transform -1 0 8170 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3498_
timestamp 0
transform -1 0 7390 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3499_
timestamp 0
transform 1 0 1130 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__3500_
timestamp 0
transform 1 0 1330 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__3501_
timestamp 0
transform -1 0 3110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3502_
timestamp 0
transform -1 0 3710 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3503_
timestamp 0
transform -1 0 3210 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3504_
timestamp 0
transform 1 0 2910 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__3505_
timestamp 0
transform 1 0 3110 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__3506_
timestamp 0
transform -1 0 730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__3507_
timestamp 0
transform -1 0 930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__3508_
timestamp 0
transform 1 0 6330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__3509_
timestamp 0
transform -1 0 6570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__3510_
timestamp 0
transform 1 0 6790 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__3511_
timestamp 0
transform -1 0 6610 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__3512_
timestamp 0
transform 1 0 6550 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__3513_
timestamp 0
transform 1 0 6730 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__3514_
timestamp 0
transform -1 0 6470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3515_
timestamp 0
transform 1 0 7130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__3516_
timestamp 0
transform -1 0 1190 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3517_
timestamp 0
transform 1 0 970 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3518_
timestamp 0
transform -1 0 7450 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3519_
timestamp 0
transform -1 0 7270 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3520_
timestamp 0
transform 1 0 5290 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3521_
timestamp 0
transform -1 0 5490 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3522_
timestamp 0
transform -1 0 50 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__3523_
timestamp 0
transform 1 0 210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3524_
timestamp 0
transform -1 0 430 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__3525_
timestamp 0
transform 1 0 2010 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__3526_
timestamp 0
transform 1 0 2190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__3527_
timestamp 0
transform 1 0 6990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__3528_
timestamp 0
transform -1 0 6930 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__3529_
timestamp 0
transform -1 0 50 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3530_
timestamp 0
transform 1 0 10070 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3531_
timestamp 0
transform 1 0 6030 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3532_
timestamp 0
transform 1 0 5650 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3533_
timestamp 0
transform 1 0 11810 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3534_
timestamp 0
transform -1 0 9110 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3535_
timestamp 0
transform 1 0 7610 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3536_
timestamp 0
transform 1 0 6010 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__3537_
timestamp 0
transform 1 0 5550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3538_
timestamp 0
transform 1 0 5530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3539_
timestamp 0
transform 1 0 6130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3540_
timestamp 0
transform 1 0 6330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3541_
timestamp 0
transform -1 0 6210 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3542_
timestamp 0
transform -1 0 6030 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3543_
timestamp 0
transform 1 0 5930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3544_
timestamp 0
transform 1 0 5810 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3545_
timestamp 0
transform 1 0 5810 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3546_
timestamp 0
transform -1 0 6190 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__3547_
timestamp 0
transform 1 0 6350 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3548_
timestamp 0
transform 1 0 6450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3549_
timestamp 0
transform 1 0 6650 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3550_
timestamp 0
transform 1 0 6510 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3551_
timestamp 0
transform -1 0 6710 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3552_
timestamp 0
transform 1 0 6790 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3553_
timestamp 0
transform -1 0 7230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__3554_
timestamp 0
transform 1 0 11190 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3555_
timestamp 0
transform 1 0 10850 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3556_
timestamp 0
transform 1 0 10110 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3557_
timestamp 0
transform -1 0 9190 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3558_
timestamp 0
transform -1 0 10690 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3559_
timestamp 0
transform 1 0 11530 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3560_
timestamp 0
transform 1 0 9990 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3561_
timestamp 0
transform 1 0 9970 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3562_
timestamp 0
transform 1 0 9770 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3563_
timestamp 0
transform -1 0 9850 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3564_
timestamp 0
transform -1 0 11790 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3565_
timestamp 0
transform 1 0 11970 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3566_
timestamp 0
transform 1 0 11390 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3567_
timestamp 0
transform 1 0 11030 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3568_
timestamp 0
transform 1 0 11170 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3569_
timestamp 0
transform 1 0 9710 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3570_
timestamp 0
transform 1 0 10610 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3571_
timestamp 0
transform 1 0 9530 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3572_
timestamp 0
transform -1 0 9370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3573_
timestamp 0
transform 1 0 10970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3574_
timestamp 0
transform -1 0 9310 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3575_
timestamp 0
transform 1 0 8510 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3576_
timestamp 0
transform -1 0 7990 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3577_
timestamp 0
transform -1 0 8970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3578_
timestamp 0
transform -1 0 9050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3579_
timestamp 0
transform -1 0 8170 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3580_
timestamp 0
transform -1 0 8630 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3581_
timestamp 0
transform 1 0 9570 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3582_
timestamp 0
transform 1 0 9370 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3583_
timestamp 0
transform 1 0 8430 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3584_
timestamp 0
transform -1 0 8370 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3585_
timestamp 0
transform 1 0 9090 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3586_
timestamp 0
transform -1 0 8930 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3587_
timestamp 0
transform -1 0 9170 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3588_
timestamp 0
transform 1 0 8170 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3589_
timestamp 0
transform -1 0 8990 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3590_
timestamp 0
transform -1 0 10570 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3591_
timestamp 0
transform -1 0 10730 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3592_
timestamp 0
transform 1 0 8190 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3593_
timestamp 0
transform -1 0 6170 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3594_
timestamp 0
transform -1 0 10330 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3595_
timestamp 0
transform -1 0 10490 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3596_
timestamp 0
transform 1 0 6930 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3597_
timestamp 0
transform 1 0 6590 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3598_
timestamp 0
transform 1 0 11810 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3599_
timestamp 0
transform -1 0 8870 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3600_
timestamp 0
transform 1 0 8650 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3601_
timestamp 0
transform 1 0 8790 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3602_
timestamp 0
transform -1 0 9910 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3603_
timestamp 0
transform -1 0 10230 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3604_
timestamp 0
transform -1 0 8390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3605_
timestamp 0
transform -1 0 7830 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3606_
timestamp 0
transform -1 0 7970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3607_
timestamp 0
transform 1 0 7770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3608_
timestamp 0
transform 1 0 11370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3609_
timestamp 0
transform 1 0 11590 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3610_
timestamp 0
transform 1 0 11450 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3611_
timestamp 0
transform 1 0 11250 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3612_
timestamp 0
transform 1 0 11610 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3613_
timestamp 0
transform 1 0 11350 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3614_
timestamp 0
transform 1 0 11550 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3615_
timestamp 0
transform 1 0 11290 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3616_
timestamp 0
transform -1 0 8070 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3617_
timestamp 0
transform 1 0 11990 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3618_
timestamp 0
transform 1 0 11930 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3619_
timestamp 0
transform -1 0 11510 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3620_
timestamp 0
transform 1 0 8750 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3621_
timestamp 0
transform 1 0 8130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3622_
timestamp 0
transform 1 0 8090 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3623_
timestamp 0
transform 1 0 11090 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3624_
timestamp 0
transform -1 0 11070 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3625_
timestamp 0
transform 1 0 10750 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3626_
timestamp 0
transform 1 0 10950 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3627_
timestamp 0
transform 1 0 10890 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3628_
timestamp 0
transform 1 0 7930 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3629_
timestamp 0
transform 1 0 7590 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3630_
timestamp 0
transform 1 0 7570 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3631_
timestamp 0
transform -1 0 7430 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3632_
timestamp 0
transform 1 0 6990 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3633_
timestamp 0
transform 1 0 7990 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3634_
timestamp 0
transform 1 0 8670 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3635_
timestamp 0
transform 1 0 8330 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3636_
timestamp 0
transform -1 0 6810 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3637_
timestamp 0
transform 1 0 8690 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3638_
timestamp 0
transform 1 0 10790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3639_
timestamp 0
transform 1 0 8550 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3640_
timestamp 0
transform 1 0 9410 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3641_
timestamp 0
transform 1 0 8910 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3642_
timestamp 0
transform -1 0 7270 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3643_
timestamp 0
transform 1 0 7070 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3644_
timestamp 0
transform -1 0 9290 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3645_
timestamp 0
transform -1 0 10370 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3646_
timestamp 0
transform 1 0 9070 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3647_
timestamp 0
transform 1 0 10510 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3648_
timestamp 0
transform 1 0 10830 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3649_
timestamp 0
transform 1 0 10930 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3650_
timestamp 0
transform -1 0 11350 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3651_
timestamp 0
transform 1 0 6730 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3652_
timestamp 0
transform 1 0 4790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3653_
timestamp 0
transform 1 0 4590 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3654_
timestamp 0
transform 1 0 4390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3655_
timestamp 0
transform 1 0 4190 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3656_
timestamp 0
transform 1 0 5390 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3657_
timestamp 0
transform 1 0 5350 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3658_
timestamp 0
transform 1 0 5190 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3659_
timestamp 0
transform 1 0 4610 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3660_
timestamp 0
transform 1 0 4410 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3661_
timestamp 0
transform 1 0 4790 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3662_
timestamp 0
transform 1 0 6530 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3663_
timestamp 0
transform 1 0 6330 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3664_
timestamp 0
transform 1 0 5570 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3665_
timestamp 0
transform 1 0 5170 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3666_
timestamp 0
transform 1 0 5770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3667_
timestamp 0
transform -1 0 3650 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3668_
timestamp 0
transform 1 0 3870 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3669_
timestamp 0
transform -1 0 3370 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3670_
timestamp 0
transform -1 0 3490 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3671_
timestamp 0
transform 1 0 4130 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3672_
timestamp 0
transform 1 0 4190 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3673_
timestamp 0
transform 1 0 5950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3674_
timestamp 0
transform -1 0 10690 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3675_
timestamp 0
transform -1 0 10510 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3676_
timestamp 0
transform 1 0 4110 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3677_
timestamp 0
transform -1 0 4170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3678_
timestamp 0
transform 1 0 4610 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3679_
timestamp 0
transform -1 0 4830 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3680_
timestamp 0
transform -1 0 5030 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3681_
timestamp 0
transform -1 0 4730 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3682_
timestamp 0
transform 1 0 1610 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__3683_
timestamp 0
transform 1 0 6230 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3684_
timestamp 0
transform 1 0 6570 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3685_
timestamp 0
transform 1 0 6850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3686_
timestamp 0
transform 1 0 6630 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3687_
timestamp 0
transform 1 0 4850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3688_
timestamp 0
transform -1 0 4870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3689_
timestamp 0
transform 1 0 5050 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3690_
timestamp 0
transform -1 0 4710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3691_
timestamp 0
transform -1 0 4650 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3692_
timestamp 0
transform 1 0 4450 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3693_
timestamp 0
transform 1 0 4830 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3694_
timestamp 0
transform -1 0 6030 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3695_
timestamp 0
transform 1 0 1670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3696_
timestamp 0
transform 1 0 7550 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3697_
timestamp 0
transform 1 0 7750 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3698_
timestamp 0
transform 1 0 6650 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3699_
timestamp 0
transform 1 0 6850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3700_
timestamp 0
transform -1 0 7050 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3701_
timestamp 0
transform 1 0 4610 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__3702_
timestamp 0
transform 1 0 4310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3703_
timestamp 0
transform 1 0 4370 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3704_
timestamp 0
transform 1 0 4790 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3705_
timestamp 0
transform -1 0 4870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3706_
timestamp 0
transform -1 0 4650 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__3707_
timestamp 0
transform -1 0 4990 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3708_
timestamp 0
transform 1 0 4570 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3709_
timestamp 0
transform 1 0 2430 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3710_
timestamp 0
transform 1 0 9750 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3711_
timestamp 0
transform 1 0 9630 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3712_
timestamp 0
transform 1 0 9610 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3713_
timestamp 0
transform 1 0 9990 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3714_
timestamp 0
transform 1 0 8690 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3715_
timestamp 0
transform -1 0 8890 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3716_
timestamp 0
transform -1 0 9490 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3717_
timestamp 0
transform -1 0 10390 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3718_
timestamp 0
transform 1 0 10550 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3719_
timestamp 0
transform -1 0 9090 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3720_
timestamp 0
transform 1 0 9270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3721_
timestamp 0
transform -1 0 10610 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3722_
timestamp 0
transform -1 0 10430 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3723_
timestamp 0
transform 1 0 10750 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3724_
timestamp 0
transform 1 0 9430 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3725_
timestamp 0
transform 1 0 8290 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3726_
timestamp 0
transform -1 0 8170 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3727_
timestamp 0
transform 1 0 9610 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3728_
timestamp 0
transform -1 0 10170 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3729_
timestamp 0
transform 1 0 10010 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3730_
timestamp 0
transform 1 0 9970 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3731_
timestamp 0
transform 1 0 8410 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3732_
timestamp 0
transform 1 0 8790 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3733_
timestamp 0
transform -1 0 3850 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3734_
timestamp 0
transform -1 0 4030 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3735_
timestamp 0
transform 1 0 7610 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3736_
timestamp 0
transform -1 0 7210 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3737_
timestamp 0
transform -1 0 5770 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3738_
timestamp 0
transform 1 0 9550 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3739_
timestamp 0
transform 1 0 9350 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3740_
timestamp 0
transform 1 0 9230 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3741_
timestamp 0
transform -1 0 10730 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3742_
timestamp 0
transform 1 0 11230 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3743_
timestamp 0
transform 1 0 11410 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3744_
timestamp 0
transform 1 0 11150 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3745_
timestamp 0
transform -1 0 10570 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3746_
timestamp 0
transform -1 0 10230 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3747_
timestamp 0
transform -1 0 10170 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3748_
timestamp 0
transform -1 0 10910 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3749_
timestamp 0
transform -1 0 11230 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3750_
timestamp 0
transform 1 0 11030 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3751_
timestamp 0
transform -1 0 8030 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3752_
timestamp 0
transform -1 0 6830 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3753_
timestamp 0
transform -1 0 6730 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3754_
timestamp 0
transform 1 0 4370 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3755_
timestamp 0
transform 1 0 3010 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3756_
timestamp 0
transform 1 0 4050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3757_
timestamp 0
transform 1 0 4530 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3758_
timestamp 0
transform -1 0 5050 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__3759_
timestamp 0
transform -1 0 4830 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__3760_
timestamp 0
transform -1 0 4270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3761_
timestamp 0
transform -1 0 4290 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__3762_
timestamp 0
transform -1 0 4390 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__3763_
timestamp 0
transform -1 0 4130 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3764_
timestamp 0
transform -1 0 3410 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3765_
timestamp 0
transform -1 0 4590 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__3766_
timestamp 0
transform 1 0 2210 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3767_
timestamp 0
transform -1 0 2430 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3768_
timestamp 0
transform -1 0 2590 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3769_
timestamp 0
transform -1 0 2790 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3770_
timestamp 0
transform -1 0 3790 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3771_
timestamp 0
transform 1 0 3370 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3772_
timestamp 0
transform -1 0 1010 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3773_
timestamp 0
transform 1 0 5790 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__3774_
timestamp 0
transform 1 0 5010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__3775_
timestamp 0
transform -1 0 4970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3776_
timestamp 0
transform -1 0 4810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3777_
timestamp 0
transform 1 0 4870 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3778_
timestamp 0
transform 1 0 4710 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3779_
timestamp 0
transform 1 0 4510 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3780_
timestamp 0
transform 1 0 5190 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3781_
timestamp 0
transform -1 0 5370 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3782_
timestamp 0
transform -1 0 4350 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3783_
timestamp 0
transform 1 0 3790 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3784_
timestamp 0
transform -1 0 5230 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3785_
timestamp 0
transform 1 0 7510 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__3786_
timestamp 0
transform 1 0 7370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__3787_
timestamp 0
transform -1 0 7350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3788_
timestamp 0
transform -1 0 7190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3789_
timestamp 0
transform -1 0 7210 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3790_
timestamp 0
transform -1 0 6190 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3791_
timestamp 0
transform -1 0 6570 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3792_
timestamp 0
transform 1 0 6990 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3793_
timestamp 0
transform -1 0 6790 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3794_
timestamp 0
transform 1 0 7950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__3795_
timestamp 0
transform -1 0 9570 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3796_
timestamp 0
transform 1 0 8270 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3797_
timestamp 0
transform 1 0 7650 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3798_
timestamp 0
transform 1 0 6930 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3799_
timestamp 0
transform -1 0 7110 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3800_
timestamp 0
transform -1 0 7290 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3801_
timestamp 0
transform 1 0 5630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3802_
timestamp 0
transform -1 0 5890 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3803_
timestamp 0
transform 1 0 5670 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3804_
timestamp 0
transform 1 0 5290 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3805_
timestamp 0
transform 1 0 5330 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3806_
timestamp 0
transform 1 0 5010 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3807_
timestamp 0
transform -1 0 5490 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3808_
timestamp 0
transform -1 0 7870 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3809_
timestamp 0
transform -1 0 7990 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3810_
timestamp 0
transform 1 0 7790 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3811_
timestamp 0
transform -1 0 7470 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3812_
timestamp 0
transform 1 0 10410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3813_
timestamp 0
transform -1 0 9830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3814_
timestamp 0
transform 1 0 9810 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3815_
timestamp 0
transform -1 0 9810 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3816_
timestamp 0
transform -1 0 9650 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3817_
timestamp 0
transform 1 0 9110 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3818_
timestamp 0
transform -1 0 8930 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3819_
timestamp 0
transform 1 0 10110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3820_
timestamp 0
transform 1 0 10190 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3821_
timestamp 0
transform 1 0 6510 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3822_
timestamp 0
transform -1 0 3310 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3823_
timestamp 0
transform -1 0 8230 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3824_
timestamp 0
transform 1 0 7250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3825_
timestamp 0
transform -1 0 9950 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3826_
timestamp 0
transform 1 0 9430 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3827_
timestamp 0
transform -1 0 9270 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3828_
timestamp 0
transform 1 0 9070 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3829_
timestamp 0
transform 1 0 8870 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3830_
timestamp 0
transform 1 0 7370 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3831_
timestamp 0
transform 1 0 7650 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3832_
timestamp 0
transform 1 0 8510 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3833_
timestamp 0
transform 1 0 8690 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3834_
timestamp 0
transform -1 0 8670 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3835_
timestamp 0
transform 1 0 8870 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3836_
timestamp 0
transform 1 0 9170 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3837_
timestamp 0
transform -1 0 8430 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3838_
timestamp 0
transform 1 0 8610 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3839_
timestamp 0
transform 1 0 8850 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3840_
timestamp 0
transform -1 0 8490 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3841_
timestamp 0
transform -1 0 8290 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3842_
timestamp 0
transform 1 0 9050 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3843_
timestamp 0
transform -1 0 8310 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3844_
timestamp 0
transform 1 0 7610 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3845_
timestamp 0
transform 1 0 9270 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__3846_
timestamp 0
transform 1 0 8830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3847_
timestamp 0
transform 1 0 8110 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3848_
timestamp 0
transform -1 0 7970 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__3849_
timestamp 0
transform 1 0 7750 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__3850_
timestamp 0
transform 1 0 7930 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3851_
timestamp 0
transform 1 0 7590 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3852_
timestamp 0
transform -1 0 7790 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3853_
timestamp 0
transform -1 0 7550 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3854_
timestamp 0
transform -1 0 7410 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3855_
timestamp 0
transform 1 0 7790 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__3856_
timestamp 0
transform -1 0 7190 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3857_
timestamp 0
transform -1 0 8290 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3858_
timestamp 0
transform 1 0 8630 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3859_
timestamp 0
transform 1 0 7810 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3860_
timestamp 0
transform 1 0 4750 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3861_
timestamp 0
transform 1 0 8490 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3862_
timestamp 0
transform -1 0 8730 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3863_
timestamp 0
transform -1 0 10190 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3864_
timestamp 0
transform 1 0 9430 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3865_
timestamp 0
transform 1 0 8010 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3866_
timestamp 0
transform 1 0 5610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3867_
timestamp 0
transform -1 0 7450 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3868_
timestamp 0
transform -1 0 8510 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3869_
timestamp 0
transform 1 0 7930 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3870_
timestamp 0
transform -1 0 7810 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3871_
timestamp 0
transform 1 0 6350 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3872_
timestamp 0
transform 1 0 5650 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3873_
timestamp 0
transform -1 0 9490 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3874_
timestamp 0
transform 1 0 9830 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__3875_
timestamp 0
transform 1 0 6870 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3876_
timestamp 0
transform 1 0 4970 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3877_
timestamp 0
transform -1 0 4610 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3878_
timestamp 0
transform 1 0 4770 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3879_
timestamp 0
transform 1 0 4530 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3880_
timestamp 0
transform 1 0 5090 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3881_
timestamp 0
transform -1 0 5310 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3882_
timestamp 0
transform -1 0 4330 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3883_
timestamp 0
transform -1 0 4950 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3884_
timestamp 0
transform -1 0 4770 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3885_
timestamp 0
transform 1 0 5130 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3886_
timestamp 0
transform 1 0 9630 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__3887_
timestamp 0
transform 1 0 10350 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__3888_
timestamp 0
transform 1 0 10310 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__3889_
timestamp 0
transform -1 0 10810 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__3890_
timestamp 0
transform -1 0 10730 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3891_
timestamp 0
transform 1 0 10890 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3892_
timestamp 0
transform -1 0 8750 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__3893_
timestamp 0
transform -1 0 8550 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__3894_
timestamp 0
transform -1 0 11250 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3895_
timestamp 0
transform 1 0 11030 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3896_
timestamp 0
transform 1 0 11790 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3897_
timestamp 0
transform 1 0 11050 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__3898_
timestamp 0
transform 1 0 8230 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3899_
timestamp 0
transform -1 0 5590 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3900_
timestamp 0
transform 1 0 4050 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3901_
timestamp 0
transform -1 0 5010 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__3902_
timestamp 0
transform 1 0 4930 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3903_
timestamp 0
transform 1 0 7410 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3904_
timestamp 0
transform -1 0 6990 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3905_
timestamp 0
transform -1 0 6430 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3906_
timestamp 0
transform 1 0 5010 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3907_
timestamp 0
transform -1 0 8170 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__3908_
timestamp 0
transform -1 0 6770 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3909_
timestamp 0
transform -1 0 5950 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__3910_
timestamp 0
transform 1 0 5830 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__3911_
timestamp 0
transform -1 0 4510 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3912_
timestamp 0
transform 1 0 4310 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__3913_
timestamp 0
transform -1 0 4530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3914_
timestamp 0
transform 1 0 4190 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__3915_
timestamp 0
transform 1 0 4730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3916_
timestamp 0
transform 1 0 4930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3917_
timestamp 0
transform 1 0 5310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3918_
timestamp 0
transform -1 0 4630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3919_
timestamp 0
transform 1 0 4730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__3920_
timestamp 0
transform 1 0 4450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3921_
timestamp 0
transform 1 0 770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3922_
timestamp 0
transform 1 0 870 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3923_
timestamp 0
transform 1 0 390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3924_
timestamp 0
transform 1 0 750 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__3925_
timestamp 0
transform 1 0 5050 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3926_
timestamp 0
transform 1 0 5250 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3927_
timestamp 0
transform -1 0 4670 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3928_
timestamp 0
transform 1 0 5430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3929_
timestamp 0
transform -1 0 4550 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__3930_
timestamp 0
transform 1 0 3390 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__3931_
timestamp 0
transform 1 0 3430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__3932_
timestamp 0
transform 1 0 2290 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__3933_
timestamp 0
transform 1 0 3190 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__3934_
timestamp 0
transform -1 0 4430 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__3935_
timestamp 0
transform 1 0 3790 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3936_
timestamp 0
transform 1 0 3590 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__3937_
timestamp 0
transform 1 0 4170 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__3938_
timestamp 0
transform -1 0 3450 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__3939_
timestamp 0
transform 1 0 3550 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__3940_
timestamp 0
transform -1 0 4690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__3941_
timestamp 0
transform 1 0 6890 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3942_
timestamp 0
transform -1 0 9970 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3943_
timestamp 0
transform -1 0 9950 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__3944_
timestamp 0
transform -1 0 9650 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__3945_
timestamp 0
transform -1 0 10170 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3946_
timestamp 0
transform 1 0 9750 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__3947_
timestamp 0
transform 1 0 10350 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3948_
timestamp 0
transform 1 0 10530 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3949_
timestamp 0
transform 1 0 7650 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__3950_
timestamp 0
transform -1 0 6930 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3951_
timestamp 0
transform 1 0 6530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3952_
timestamp 0
transform -1 0 5750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__3953_
timestamp 0
transform 1 0 5410 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3954_
timestamp 0
transform -1 0 5810 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3955_
timestamp 0
transform 1 0 5870 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3956_
timestamp 0
transform -1 0 6090 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3957_
timestamp 0
transform 1 0 6110 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3958_
timestamp 0
transform 1 0 6310 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3959_
timestamp 0
transform 1 0 6430 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3960_
timestamp 0
transform 1 0 2350 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3961_
timestamp 0
transform -1 0 2750 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3962_
timestamp 0
transform 1 0 2890 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3963_
timestamp 0
transform 1 0 3490 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3964_
timestamp 0
transform -1 0 4070 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3965_
timestamp 0
transform -1 0 3310 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3966_
timestamp 0
transform -1 0 4270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3967_
timestamp 0
transform -1 0 5070 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3968_
timestamp 0
transform -1 0 5270 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3969_
timestamp 0
transform -1 0 4270 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3970_
timestamp 0
transform 1 0 3890 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3971_
timestamp 0
transform 1 0 5590 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__3972_
timestamp 0
transform 1 0 5410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__3973_
timestamp 0
transform 1 0 5410 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3974_
timestamp 0
transform -1 0 5630 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3975_
timestamp 0
transform -1 0 5630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3976_
timestamp 0
transform -1 0 5630 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3977_
timestamp 0
transform 1 0 5510 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__3978_
timestamp 0
transform 1 0 6330 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3979_
timestamp 0
transform -1 0 2690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3980_
timestamp 0
transform 1 0 1990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__3981_
timestamp 0
transform 1 0 1830 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__3982_
timestamp 0
transform 1 0 1770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__3983_
timestamp 0
transform -1 0 1910 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__3984_
timestamp 0
transform 1 0 8230 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__3985_
timestamp 0
transform 1 0 6810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3986_
timestamp 0
transform -1 0 7310 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__3987_
timestamp 0
transform 1 0 7590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3988_
timestamp 0
transform 1 0 7510 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3989_
timestamp 0
transform 1 0 7310 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3990_
timestamp 0
transform 1 0 7110 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3991_
timestamp 0
transform -1 0 7270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__3992_
timestamp 0
transform -1 0 7930 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3993_
timestamp 0
transform 1 0 7690 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3994_
timestamp 0
transform -1 0 7030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__3995_
timestamp 0
transform -1 0 9390 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3996_
timestamp 0
transform -1 0 5990 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__3997_
timestamp 0
transform 1 0 5950 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__3998_
timestamp 0
transform -1 0 6030 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__3999_
timestamp 0
transform 1 0 5810 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4000_
timestamp 0
transform -1 0 5230 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4001_
timestamp 0
transform -1 0 5070 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4002_
timestamp 0
transform -1 0 6930 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4003_
timestamp 0
transform -1 0 6570 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4004_
timestamp 0
transform 1 0 2610 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4005_
timestamp 0
transform 1 0 2810 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4006_
timestamp 0
transform -1 0 2630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4007_
timestamp 0
transform 1 0 2410 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4008_
timestamp 0
transform -1 0 7090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4009_
timestamp 0
transform 1 0 6870 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4010_
timestamp 0
transform -1 0 6730 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4011_
timestamp 0
transform 1 0 8610 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4012_
timestamp 0
transform 1 0 6710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4013_
timestamp 0
transform 1 0 6590 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4014_
timestamp 0
transform 1 0 6130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4015_
timestamp 0
transform 1 0 6490 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4016_
timestamp 0
transform 1 0 9310 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4017_
timestamp 0
transform -1 0 9630 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4018_
timestamp 0
transform -1 0 9810 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4019_
timestamp 0
transform 1 0 9970 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4020_
timestamp 0
transform -1 0 7450 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4021_
timestamp 0
transform -1 0 10010 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4022_
timestamp 0
transform -1 0 6790 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4023_
timestamp 0
transform -1 0 7130 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4024_
timestamp 0
transform 1 0 8930 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4025_
timestamp 0
transform -1 0 7650 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4026_
timestamp 0
transform -1 0 7810 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4027_
timestamp 0
transform 1 0 8350 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4028_
timestamp 0
transform 1 0 7890 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4029_
timestamp 0
transform 1 0 10990 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4030_
timestamp 0
transform 1 0 10810 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4031_
timestamp 0
transform 1 0 9190 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4032_
timestamp 0
transform 1 0 8630 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4033_
timestamp 0
transform -1 0 9290 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4034_
timestamp 0
transform 1 0 3950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4035_
timestamp 0
transform 1 0 9750 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4036_
timestamp 0
transform -1 0 9610 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4037_
timestamp 0
transform -1 0 9130 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4038_
timestamp 0
transform -1 0 8090 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4039_
timestamp 0
transform -1 0 7030 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4040_
timestamp 0
transform 1 0 11970 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4041_
timestamp 0
transform 1 0 9250 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4042_
timestamp 0
transform -1 0 5970 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__4043_
timestamp 0
transform 1 0 5290 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4044_
timestamp 0
transform -1 0 5370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4045_
timestamp 0
transform -1 0 5430 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4046_
timestamp 0
transform -1 0 5790 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4047_
timestamp 0
transform -1 0 5970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4048_
timestamp 0
transform -1 0 5970 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4049_
timestamp 0
transform 1 0 5450 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4050_
timestamp 0
transform -1 0 5230 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4051_
timestamp 0
transform 1 0 5570 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4052_
timestamp 0
transform -1 0 6190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4053_
timestamp 0
transform -1 0 8170 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4054_
timestamp 0
transform 1 0 3690 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4055_
timestamp 0
transform -1 0 3530 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4056_
timestamp 0
transform 1 0 2690 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4057_
timestamp 0
transform 1 0 3310 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4058_
timestamp 0
transform -1 0 7450 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4059_
timestamp 0
transform 1 0 7310 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4060_
timestamp 0
transform -1 0 7990 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4061_
timestamp 0
transform -1 0 8930 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4062_
timestamp 0
transform -1 0 3110 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4063_
timestamp 0
transform 1 0 5030 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4064_
timestamp 0
transform -1 0 5010 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4065_
timestamp 0
transform 1 0 5230 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4066_
timestamp 0
transform 1 0 4430 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4067_
timestamp 0
transform -1 0 7070 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4068_
timestamp 0
transform 1 0 3090 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4069_
timestamp 0
transform -1 0 630 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__4070_
timestamp 0
transform 1 0 1110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__4071_
timestamp 0
transform 1 0 510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__4072_
timestamp 0
transform -1 0 830 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__4073_
timestamp 0
transform 1 0 4050 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4074_
timestamp 0
transform 1 0 4250 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4075_
timestamp 0
transform 1 0 4170 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4076_
timestamp 0
transform -1 0 5430 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4077_
timestamp 0
transform 1 0 5450 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4078_
timestamp 0
transform -1 0 5470 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4079_
timestamp 0
transform 1 0 3730 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4080_
timestamp 0
transform 1 0 5830 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4081_
timestamp 0
transform 1 0 870 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4082_
timestamp 0
transform 1 0 4110 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4083_
timestamp 0
transform -1 0 3910 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4084_
timestamp 0
transform 1 0 1610 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4085_
timestamp 0
transform 1 0 1430 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4086_
timestamp 0
transform 1 0 1570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4087_
timestamp 0
transform 1 0 1530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4088_
timestamp 0
transform -1 0 4470 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4089_
timestamp 0
transform -1 0 4430 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4090_
timestamp 0
transform -1 0 3930 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4091_
timestamp 0
transform -1 0 3370 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4092_
timestamp 0
transform -1 0 5650 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4093_
timestamp 0
transform 1 0 4590 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4094_
timestamp 0
transform 1 0 4170 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4095_
timestamp 0
transform 1 0 1910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4096_
timestamp 0
transform 1 0 1730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4097_
timestamp 0
transform 1 0 1610 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4098_
timestamp 0
transform 1 0 1530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4099_
timestamp 0
transform 1 0 7110 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4100_
timestamp 0
transform 1 0 7990 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4101_
timestamp 0
transform 1 0 8150 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4102_
timestamp 0
transform -1 0 8350 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4103_
timestamp 0
transform 1 0 7970 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4104_
timestamp 0
transform -1 0 8190 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4105_
timestamp 0
transform 1 0 8630 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4106_
timestamp 0
transform 1 0 6670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4107_
timestamp 0
transform -1 0 1070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1__4108_
timestamp 0
transform -1 0 470 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__4109_
timestamp 0
transform -1 0 1810 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4110_
timestamp 0
transform -1 0 7750 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4111_
timestamp 0
transform -1 0 9490 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4112_
timestamp 0
transform 1 0 2870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__4113_
timestamp 0
transform 1 0 3070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__4114_
timestamp 0
transform 1 0 3570 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4115_
timestamp 0
transform 1 0 4450 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4116_
timestamp 0
transform -1 0 5330 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4117_
timestamp 0
transform 1 0 4870 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4118_
timestamp 0
transform 1 0 4790 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4119_
timestamp 0
transform 1 0 3950 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4120_
timestamp 0
transform -1 0 3690 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4121_
timestamp 0
transform -1 0 4530 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4122_
timestamp 0
transform 1 0 4670 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4123_
timestamp 0
transform 1 0 8030 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4124_
timestamp 0
transform 1 0 8550 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4125_
timestamp 0
transform -1 0 4270 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4126_
timestamp 0
transform 1 0 4230 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4127_
timestamp 0
transform 1 0 4050 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4128_
timestamp 0
transform 1 0 4470 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4129_
timestamp 0
transform -1 0 4890 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4130_
timestamp 0
transform 1 0 6010 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4131_
timestamp 0
transform 1 0 4290 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4132_
timestamp 0
transform -1 0 4510 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4133_
timestamp 0
transform -1 0 1990 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4134_
timestamp 0
transform 1 0 1770 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4135_
timestamp 0
transform -1 0 2130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4136_
timestamp 0
transform -1 0 2130 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4137_
timestamp 0
transform -1 0 1970 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4138_
timestamp 0
transform -1 0 2210 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4139_
timestamp 0
transform 1 0 1990 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4140_
timestamp 0
transform -1 0 3010 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4141_
timestamp 0
transform 1 0 1790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4142_
timestamp 0
transform 1 0 1590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4143_
timestamp 0
transform -1 0 1430 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4144_
timestamp 0
transform 1 0 1570 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4145_
timestamp 0
transform -1 0 1050 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4146_
timestamp 0
transform 1 0 3070 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4147_
timestamp 0
transform -1 0 2010 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4148_
timestamp 0
transform -1 0 3190 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4149_
timestamp 0
transform 1 0 3170 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4150_
timestamp 0
transform 1 0 3170 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4151_
timestamp 0
transform 1 0 3710 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4152_
timestamp 0
transform -1 0 3650 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4153_
timestamp 0
transform -1 0 2030 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4154_
timestamp 0
transform -1 0 2230 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4155_
timestamp 0
transform 1 0 610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4156_
timestamp 0
transform 1 0 970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4157_
timestamp 0
transform -1 0 5910 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4158_
timestamp 0
transform 1 0 6070 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4159_
timestamp 0
transform 1 0 6270 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4160_
timestamp 0
transform 1 0 5350 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4161_
timestamp 0
transform -1 0 5570 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4162_
timestamp 0
transform 1 0 5150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4163_
timestamp 0
transform -1 0 5170 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4164_
timestamp 0
transform 1 0 5710 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4165_
timestamp 0
transform -1 0 5710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4166_
timestamp 0
transform 1 0 5730 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4167_
timestamp 0
transform 1 0 6430 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4168_
timestamp 0
transform -1 0 5870 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4169_
timestamp 0
transform 1 0 5670 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4170_
timestamp 0
transform 1 0 6070 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4171_
timestamp 0
transform 1 0 5490 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4172_
timestamp 0
transform 1 0 5110 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4173_
timestamp 0
transform 1 0 3790 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4174_
timestamp 0
transform 1 0 5510 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4175_
timestamp 0
transform 1 0 5130 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4176_
timestamp 0
transform -1 0 3310 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4177_
timestamp 0
transform 1 0 2990 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4178_
timestamp 0
transform -1 0 2210 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4179_
timestamp 0
transform -1 0 2330 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4180_
timestamp 0
transform 1 0 2790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4181_
timestamp 0
transform -1 0 2410 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4182_
timestamp 0
transform 1 0 2250 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4183_
timestamp 0
transform -1 0 3230 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4184_
timestamp 0
transform 1 0 3390 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4185_
timestamp 0
transform 1 0 2810 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4186_
timestamp 0
transform -1 0 2430 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4187_
timestamp 0
transform 1 0 4050 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4188_
timestamp 0
transform 1 0 4250 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4189_
timestamp 0
transform -1 0 4070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4190_
timestamp 0
transform -1 0 3890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4191_
timestamp 0
transform -1 0 3710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4192_
timestamp 0
transform -1 0 5170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4193_
timestamp 0
transform -1 0 5030 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4194_
timestamp 0
transform -1 0 3890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4195_
timestamp 0
transform 1 0 3430 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4196_
timestamp 0
transform 1 0 3730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4197_
timestamp 0
transform 1 0 1590 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4198_
timestamp 0
transform -1 0 1710 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4199_
timestamp 0
transform -1 0 1910 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4200_
timestamp 0
transform -1 0 2310 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4201_
timestamp 0
transform -1 0 1530 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4202_
timestamp 0
transform -1 0 1410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__4203_
timestamp 0
transform -1 0 1790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__4204_
timestamp 0
transform -1 0 2590 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4205_
timestamp 0
transform 1 0 2590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4206_
timestamp 0
transform -1 0 8570 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4207_
timestamp 0
transform -1 0 7910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4208_
timestamp 0
transform -1 0 6250 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4209_
timestamp 0
transform -1 0 250 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4210_
timestamp 0
transform 1 0 30 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4211_
timestamp 0
transform -1 0 50 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4212_
timestamp 0
transform -1 0 430 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4213_
timestamp 0
transform 1 0 890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4214_
timestamp 0
transform -1 0 1410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4215_
timestamp 0
transform 1 0 1390 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4216_
timestamp 0
transform -1 0 1990 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4217_
timestamp 0
transform -1 0 2970 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4218_
timestamp 0
transform -1 0 2190 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4219_
timestamp 0
transform 1 0 2270 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4220_
timestamp 0
transform 1 0 2470 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4221_
timestamp 0
transform -1 0 250 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4222_
timestamp 0
transform -1 0 50 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4223_
timestamp 0
transform -1 0 430 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4224_
timestamp 0
transform -1 0 430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4225_
timestamp 0
transform -1 0 410 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4226_
timestamp 0
transform 1 0 30 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4227_
timestamp 0
transform -1 0 250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4228_
timestamp 0
transform -1 0 2390 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4229_
timestamp 0
transform 1 0 2590 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4230_
timestamp 0
transform -1 0 2810 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4231_
timestamp 0
transform 1 0 3150 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4232_
timestamp 0
transform -1 0 3610 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4233_
timestamp 0
transform -1 0 2190 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4234_
timestamp 0
transform -1 0 3050 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4235_
timestamp 0
transform -1 0 3810 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4236_
timestamp 0
transform 1 0 3890 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4237_
timestamp 0
transform -1 0 4110 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4238_
timestamp 0
transform 1 0 3430 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4239_
timestamp 0
transform 1 0 2590 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4240_
timestamp 0
transform 1 0 2230 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4241_
timestamp 0
transform -1 0 2090 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4242_
timestamp 0
transform 1 0 2270 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4243_
timestamp 0
transform -1 0 4450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4244_
timestamp 0
transform -1 0 5450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4245_
timestamp 0
transform -1 0 6030 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4246_
timestamp 0
transform -1 0 4150 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4247_
timestamp 0
transform 1 0 2550 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4248_
timestamp 0
transform -1 0 5630 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4249_
timestamp 0
transform -1 0 2330 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4250_
timestamp 0
transform -1 0 4250 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4251_
timestamp 0
transform 1 0 5630 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4252_
timestamp 0
transform -1 0 5830 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4253_
timestamp 0
transform -1 0 3730 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4254_
timestamp 0
transform -1 0 2150 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4255_
timestamp 0
transform 1 0 2490 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4256_
timestamp 0
transform -1 0 3850 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4257_
timestamp 0
transform 1 0 4030 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4258_
timestamp 0
transform 1 0 4230 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4259_
timestamp 0
transform 1 0 3990 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4260_
timestamp 0
transform -1 0 2950 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4261_
timestamp 0
transform -1 0 4010 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4262_
timestamp 0
transform 1 0 1530 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4263_
timestamp 0
transform -1 0 7950 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4264_
timestamp 0
transform 1 0 7570 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4265_
timestamp 0
transform 1 0 7390 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4266_
timestamp 0
transform 1 0 7070 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4267_
timestamp 0
transform 1 0 7510 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4268_
timestamp 0
transform -1 0 6750 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4269_
timestamp 0
transform -1 0 9430 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4270_
timestamp 0
transform -1 0 11130 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4271_
timestamp 0
transform 1 0 11110 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4272_
timestamp 0
transform 1 0 9210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4273_
timestamp 0
transform 1 0 9010 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4274_
timestamp 0
transform -1 0 8930 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4275_
timestamp 0
transform 1 0 8750 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4276_
timestamp 0
transform 1 0 8830 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4277_
timestamp 0
transform 1 0 8850 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4278_
timestamp 0
transform 1 0 7730 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4279_
timestamp 0
transform 1 0 10510 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4280_
timestamp 0
transform 1 0 10710 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4281_
timestamp 0
transform -1 0 10670 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4282_
timestamp 0
transform -1 0 1210 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4283_
timestamp 0
transform -1 0 7050 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4284_
timestamp 0
transform 1 0 7630 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4285_
timestamp 0
transform 1 0 7370 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4286_
timestamp 0
transform -1 0 1050 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4287_
timestamp 0
transform -1 0 1250 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4288_
timestamp 0
transform -1 0 1650 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4289_
timestamp 0
transform -1 0 4350 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4290_
timestamp 0
transform 1 0 6830 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4291_
timestamp 0
transform 1 0 6850 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4292_
timestamp 0
transform -1 0 2510 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4293_
timestamp 0
transform -1 0 1790 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4294_
timestamp 0
transform -1 0 7270 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4295_
timestamp 0
transform 1 0 1470 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4296_
timestamp 0
transform -1 0 50 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4297_
timestamp 0
transform 1 0 1130 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4298_
timestamp 0
transform -1 0 3250 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4299_
timestamp 0
transform 1 0 3330 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4300_
timestamp 0
transform -1 0 3810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4301_
timestamp 0
transform -1 0 3530 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4302_
timestamp 0
transform -1 0 3650 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4303_
timestamp 0
transform -1 0 1570 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4304_
timestamp 0
transform 1 0 1150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4305_
timestamp 0
transform -1 0 2270 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4306_
timestamp 0
transform -1 0 2830 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4307_
timestamp 0
transform 1 0 6190 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4308_
timestamp 0
transform -1 0 6270 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4309_
timestamp 0
transform 1 0 2830 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4310_
timestamp 0
transform -1 0 2410 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4311_
timestamp 0
transform 1 0 2310 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4312_
timestamp 0
transform 1 0 890 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4313_
timestamp 0
transform 1 0 1470 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4314_
timestamp 0
transform 1 0 1650 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4315_
timestamp 0
transform -1 0 2690 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4316_
timestamp 0
transform -1 0 2750 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4317_
timestamp 0
transform 1 0 4390 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4318_
timestamp 0
transform 1 0 4070 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4319_
timestamp 0
transform 1 0 3570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4320_
timestamp 0
transform -1 0 3010 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4321_
timestamp 0
transform 1 0 2790 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4322_
timestamp 0
transform 1 0 1530 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4323_
timestamp 0
transform -1 0 2650 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4324_
timestamp 0
transform -1 0 1790 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4325_
timestamp 0
transform -1 0 4050 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4326_
timestamp 0
transform 1 0 3950 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4327_
timestamp 0
transform 1 0 4090 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4328_
timestamp 0
transform -1 0 8530 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4329_
timestamp 0
transform 1 0 1690 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4330_
timestamp 0
transform 1 0 2090 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4331_
timestamp 0
transform -1 0 1410 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4332_
timestamp 0
transform -1 0 1950 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4333_
timestamp 0
transform -1 0 2870 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4334_
timestamp 0
transform -1 0 3070 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4335_
timestamp 0
transform -1 0 3650 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4336_
timestamp 0
transform 1 0 2810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4337_
timestamp 0
transform 1 0 2610 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4338_
timestamp 0
transform 1 0 2650 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4339_
timestamp 0
transform -1 0 3270 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4340_
timestamp 0
transform -1 0 3450 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4341_
timestamp 0
transform 1 0 3390 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4342_
timestamp 0
transform -1 0 3210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4343_
timestamp 0
transform 1 0 3450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4344_
timestamp 0
transform 1 0 1750 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4345_
timestamp 0
transform -1 0 2390 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4346_
timestamp 0
transform 1 0 6870 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4347_
timestamp 0
transform -1 0 6690 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4348_
timestamp 0
transform -1 0 590 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4349_
timestamp 0
transform -1 0 1010 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4350_
timestamp 0
transform 1 0 2130 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4351_
timestamp 0
transform -1 0 2750 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4352_
timestamp 0
transform 1 0 3730 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4353_
timestamp 0
transform -1 0 6130 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4354_
timestamp 0
transform -1 0 3410 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4355_
timestamp 0
transform -1 0 830 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4356_
timestamp 0
transform -1 0 470 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4357_
timestamp 0
transform 1 0 2330 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4358_
timestamp 0
transform -1 0 5190 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4359_
timestamp 0
transform 1 0 5110 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4360_
timestamp 0
transform -1 0 5070 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4361_
timestamp 0
transform 1 0 3010 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4362_
timestamp 0
transform 1 0 4850 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4363_
timestamp 0
transform -1 0 4690 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4364_
timestamp 0
transform 1 0 3650 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4365_
timestamp 0
transform -1 0 5630 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4366_
timestamp 0
transform -1 0 5830 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4367_
timestamp 0
transform -1 0 2870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4368_
timestamp 0
transform 1 0 7510 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4369_
timestamp 0
transform -1 0 7350 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4370_
timestamp 0
transform 1 0 630 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4371_
timestamp 0
transform -1 0 1770 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4372_
timestamp 0
transform 1 0 1890 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4373_
timestamp 0
transform 1 0 2090 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4374_
timestamp 0
transform 1 0 2450 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4375_
timestamp 0
transform -1 0 3770 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4376_
timestamp 0
transform 1 0 7450 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4377_
timestamp 0
transform 1 0 11510 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4378_
timestamp 0
transform -1 0 1230 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4379_
timestamp 0
transform -1 0 5190 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4380_
timestamp 0
transform 1 0 4770 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4381_
timestamp 0
transform 1 0 5870 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4382_
timestamp 0
transform 1 0 210 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4383_
timestamp 0
transform 1 0 30 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4384_
timestamp 0
transform 1 0 6210 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4385_
timestamp 0
transform 1 0 6410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4386_
timestamp 0
transform 1 0 6810 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4387_
timestamp 0
transform 1 0 6610 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4388_
timestamp 0
transform -1 0 5410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4389_
timestamp 0
transform -1 0 6510 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4390_
timestamp 0
transform 1 0 7010 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4391_
timestamp 0
transform 1 0 4970 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4392_
timestamp 0
transform -1 0 6310 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4393_
timestamp 0
transform 1 0 6470 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4394_
timestamp 0
transform 1 0 6650 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4395_
timestamp 0
transform 1 0 6770 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4396_
timestamp 0
transform -1 0 6250 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4397_
timestamp 0
transform 1 0 4010 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4398_
timestamp 0
transform 1 0 2990 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4399_
timestamp 0
transform 1 0 2110 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4400_
timestamp 0
transform -1 0 6290 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4401_
timestamp 0
transform 1 0 6210 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4402_
timestamp 0
transform -1 0 6050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4403_
timestamp 0
transform -1 0 5590 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4404_
timestamp 0
transform 1 0 1370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4405_
timestamp 0
transform -1 0 1810 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4406_
timestamp 0
transform -1 0 2510 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4407_
timestamp 0
transform -1 0 2310 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4408_
timestamp 0
transform 1 0 1530 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4409_
timestamp 0
transform -1 0 1750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4410_
timestamp 0
transform 1 0 3550 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4411_
timestamp 0
transform 1 0 3870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4412_
timestamp 0
transform 1 0 1710 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4413_
timestamp 0
transform -1 0 230 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4414_
timestamp 0
transform 1 0 230 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4415_
timestamp 0
transform 1 0 410 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4416_
timestamp 0
transform 1 0 1490 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__4417_
timestamp 0
transform -1 0 1710 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__4418_
timestamp 0
transform -1 0 2530 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__4419_
timestamp 0
transform 1 0 2090 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__4420_
timestamp 0
transform 1 0 2210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4421_
timestamp 0
transform 1 0 2410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4422_
timestamp 0
transform -1 0 1950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4423_
timestamp 0
transform -1 0 590 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4424_
timestamp 0
transform 1 0 2010 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4425_
timestamp 0
transform 1 0 1050 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4426_
timestamp 0
transform 1 0 1250 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4427_
timestamp 0
transform 1 0 3510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4428_
timestamp 0
transform -1 0 3350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4429_
timestamp 0
transform 1 0 1230 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4430_
timestamp 0
transform 1 0 1430 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4431_
timestamp 0
transform -1 0 710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4432_
timestamp 0
transform -1 0 590 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4433_
timestamp 0
transform -1 0 830 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4434_
timestamp 0
transform -1 0 1290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__4435_
timestamp 0
transform 1 0 1470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__4436_
timestamp 0
transform 1 0 3070 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__4437_
timestamp 0
transform -1 0 3290 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__4438_
timestamp 0
transform -1 0 6530 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4439_
timestamp 0
transform 1 0 5930 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4440_
timestamp 0
transform -1 0 4710 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4441_
timestamp 0
transform 1 0 4110 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4442_
timestamp 0
transform 1 0 3890 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4443_
timestamp 0
transform 1 0 3770 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4444_
timestamp 0
transform 1 0 3590 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4445_
timestamp 0
transform 1 0 3930 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4446_
timestamp 0
transform 1 0 4350 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4447_
timestamp 0
transform 1 0 4530 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4448_
timestamp 0
transform 1 0 2450 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4449_
timestamp 0
transform 1 0 1010 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4450_
timestamp 0
transform -1 0 1770 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4451_
timestamp 0
transform 1 0 1370 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4452_
timestamp 0
transform -1 0 2170 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4453_
timestamp 0
transform 1 0 7190 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4454_
timestamp 0
transform -1 0 1010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4455_
timestamp 0
transform 1 0 6730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4456_
timestamp 0
transform 1 0 6950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4457_
timestamp 0
transform 1 0 7150 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4458_
timestamp 0
transform -1 0 7350 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4459_
timestamp 0
transform -1 0 6970 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4460_
timestamp 0
transform -1 0 8290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4461_
timestamp 0
transform 1 0 7570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4462_
timestamp 0
transform -1 0 6670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4463_
timestamp 0
transform 1 0 1190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4464_
timestamp 0
transform -1 0 2490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4465_
timestamp 0
transform -1 0 5830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4466_
timestamp 0
transform 1 0 5970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4467_
timestamp 0
transform 1 0 6390 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4468_
timestamp 0
transform 1 0 6630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4469_
timestamp 0
transform 1 0 6830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4470_
timestamp 0
transform -1 0 6590 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4471_
timestamp 0
transform 1 0 7190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4472_
timestamp 0
transform -1 0 6390 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4473_
timestamp 0
transform 1 0 8110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4474_
timestamp 0
transform -1 0 6210 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4475_
timestamp 0
transform 1 0 2670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4476_
timestamp 0
transform -1 0 1170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4477_
timestamp 0
transform -1 0 2570 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4478_
timestamp 0
transform 1 0 2550 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4479_
timestamp 0
transform 1 0 5270 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4480_
timestamp 0
transform 1 0 1350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4481_
timestamp 0
transform 1 0 190 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4482_
timestamp 0
transform 1 0 390 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4483_
timestamp 0
transform 1 0 3150 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4484_
timestamp 0
transform -1 0 4910 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4485_
timestamp 0
transform 1 0 5290 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4486_
timestamp 0
transform -1 0 5110 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4487_
timestamp 0
transform -1 0 5490 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4488_
timestamp 0
transform 1 0 5650 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4489_
timestamp 0
transform -1 0 5770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4490_
timestamp 0
transform -1 0 5730 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4491_
timestamp 0
transform -1 0 5810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4492_
timestamp 0
transform 1 0 30 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4493_
timestamp 0
transform -1 0 5650 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4494_
timestamp 0
transform 1 0 5450 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4495_
timestamp 0
transform 1 0 4310 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4496_
timestamp 0
transform 1 0 3770 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4497_
timestamp 0
transform -1 0 3550 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4498_
timestamp 0
transform -1 0 4590 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4499_
timestamp 0
transform 1 0 1210 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4500_
timestamp 0
transform 1 0 6310 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4501_
timestamp 0
transform 1 0 6030 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4502_
timestamp 0
transform -1 0 4470 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4503_
timestamp 0
transform 1 0 6430 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4504_
timestamp 0
transform -1 0 1670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__4505_
timestamp 0
transform -1 0 4790 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__4506_
timestamp 0
transform -1 0 5230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4507_
timestamp 0
transform 1 0 5610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__4508_
timestamp 0
transform 1 0 5490 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4509_
timestamp 0
transform -1 0 5710 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4510_
timestamp 0
transform -1 0 5890 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4511_
timestamp 0
transform 1 0 6050 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4512_
timestamp 0
transform 1 0 6150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4513_
timestamp 0
transform 1 0 6170 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4514_
timestamp 0
transform -1 0 1670 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__4515_
timestamp 0
transform -1 0 2510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__4516_
timestamp 0
transform -1 0 4630 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__4517_
timestamp 0
transform -1 0 5110 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4518_
timestamp 0
transform 1 0 5070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4519_
timestamp 0
transform 1 0 5430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4520_
timestamp 0
transform -1 0 5630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4521_
timestamp 0
transform 1 0 6470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4522_
timestamp 0
transform -1 0 8890 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4523_
timestamp 0
transform 1 0 5270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4524_
timestamp 0
transform 1 0 5970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4525_
timestamp 0
transform 1 0 5830 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4526_
timestamp 0
transform -1 0 6410 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4527_
timestamp 0
transform -1 0 4910 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4528_
timestamp 0
transform 1 0 6310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4529_
timestamp 0
transform 1 0 6010 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4530_
timestamp 0
transform 1 0 5990 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4531_
timestamp 0
transform -1 0 2230 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__4532_
timestamp 0
transform -1 0 6250 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4533_
timestamp 0
transform -1 0 6190 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4534_
timestamp 0
transform 1 0 4230 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4535_
timestamp 0
transform 1 0 3630 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4536_
timestamp 0
transform -1 0 1050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4537_
timestamp 0
transform 1 0 4410 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4538_
timestamp 0
transform -1 0 7650 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4539_
timestamp 0
transform -1 0 3030 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4540_
timestamp 0
transform 1 0 7610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4541_
timestamp 0
transform 1 0 6470 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4542_
timestamp 0
transform 1 0 3010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4543_
timestamp 0
transform -1 0 2850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4544_
timestamp 0
transform -1 0 870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4545_
timestamp 0
transform 1 0 2090 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4546_
timestamp 0
transform 1 0 2870 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4547_
timestamp 0
transform -1 0 2330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4548_
timestamp 0
transform -1 0 1710 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4549_
timestamp 0
transform 1 0 2570 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4550_
timestamp 0
transform 1 0 2770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4551_
timestamp 0
transform -1 0 2970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4552_
timestamp 0
transform -1 0 2950 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4553_
timestamp 0
transform -1 0 6510 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4554_
timestamp 0
transform 1 0 950 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4555_
timestamp 0
transform -1 0 710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__4556_
timestamp 0
transform 1 0 4310 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4557_
timestamp 0
transform 1 0 4130 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4558_
timestamp 0
transform -1 0 3970 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4559_
timestamp 0
transform 1 0 4990 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4560_
timestamp 0
transform -1 0 8450 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4561_
timestamp 0
transform -1 0 8850 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4562_
timestamp 0
transform 1 0 8370 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4563_
timestamp 0
transform -1 0 6350 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4564_
timestamp 0
transform -1 0 1850 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4565_
timestamp 0
transform 1 0 2670 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4566_
timestamp 0
transform 1 0 3050 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4567_
timestamp 0
transform -1 0 6750 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4568_
timestamp 0
transform 1 0 6670 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4569_
timestamp 0
transform 1 0 1890 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4570_
timestamp 0
transform -1 0 6550 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4571_
timestamp 0
transform 1 0 6250 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4572_
timestamp 0
transform -1 0 9490 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4573_
timestamp 0
transform -1 0 10350 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4574_
timestamp 0
transform -1 0 9530 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4575_
timestamp 0
transform -1 0 6950 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4576_
timestamp 0
transform -1 0 8470 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4577_
timestamp 0
transform -1 0 2990 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4578_
timestamp 0
transform -1 0 5950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4579_
timestamp 0
transform 1 0 7970 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4580_
timestamp 0
transform 1 0 10150 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4581_
timestamp 0
transform -1 0 7490 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4582_
timestamp 0
transform 1 0 1250 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4583_
timestamp 0
transform -1 0 2330 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4584_
timestamp 0
transform -1 0 2170 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4585_
timestamp 0
transform -1 0 2070 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4586_
timestamp 0
transform -1 0 1890 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4587_
timestamp 0
transform -1 0 1550 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4588_
timestamp 0
transform 1 0 3270 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4589_
timestamp 0
transform 1 0 3810 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4590_
timestamp 0
transform 1 0 1190 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4591_
timestamp 0
transform -1 0 1610 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4592_
timestamp 0
transform 1 0 1410 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4593_
timestamp 0
transform -1 0 3970 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4594_
timestamp 0
transform -1 0 3130 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__4595_
timestamp 0
transform -1 0 2690 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4596_
timestamp 0
transform -1 0 2890 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4597_
timestamp 0
transform 1 0 2750 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__4598_
timestamp 0
transform -1 0 2670 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4599_
timestamp 0
transform -1 0 2850 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4600_
timestamp 0
transform -1 0 4010 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4601_
timestamp 0
transform -1 0 3970 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4602_
timestamp 0
transform -1 0 1390 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4603_
timestamp 0
transform -1 0 1330 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4604_
timestamp 0
transform -1 0 2930 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__4605_
timestamp 0
transform 1 0 1750 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4606_
timestamp 0
transform -1 0 650 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4607_
timestamp 0
transform -1 0 470 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4608_
timestamp 0
transform -1 0 3210 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4609_
timestamp 0
transform 1 0 1590 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__4610_
timestamp 0
transform 1 0 2470 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4611_
timestamp 0
transform -1 0 2310 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4612_
timestamp 0
transform -1 0 1970 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4613_
timestamp 0
transform 1 0 1950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__4614_
timestamp 0
transform -1 0 610 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4615_
timestamp 0
transform -1 0 430 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4616_
timestamp 0
transform -1 0 1790 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__4617_
timestamp 0
transform -1 0 1590 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__4618_
timestamp 0
transform -1 0 2490 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4619_
timestamp 0
transform -1 0 1830 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4620_
timestamp 0
transform -1 0 1430 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4621_
timestamp 0
transform 1 0 2090 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4622_
timestamp 0
transform 1 0 2510 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4623_
timestamp 0
transform 1 0 2010 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4624_
timestamp 0
transform 1 0 1210 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4625_
timestamp 0
transform 1 0 830 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4626_
timestamp 0
transform -1 0 670 0 1 11290
box -6 -8 26 248
use FILL  FILL_1__4627_
timestamp 0
transform -1 0 2170 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__4628_
timestamp 0
transform -1 0 1230 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__4629_
timestamp 0
transform 1 0 1010 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1__4630_
timestamp 0
transform 1 0 970 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4631_
timestamp 0
transform 1 0 1550 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4632_
timestamp 0
transform -1 0 710 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4633_
timestamp 0
transform -1 0 530 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4634_
timestamp 0
transform -1 0 7550 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4635_
timestamp 0
transform -1 0 1490 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4636_
timestamp 0
transform 1 0 1290 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4637_
timestamp 0
transform -1 0 1690 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4638_
timestamp 0
transform -1 0 850 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1__4639_
timestamp 0
transform 1 0 1050 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4640_
timestamp 0
transform 1 0 910 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4641_
timestamp 0
transform -1 0 1070 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4642_
timestamp 0
transform -1 0 2890 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__4643_
timestamp 0
transform 1 0 3030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1__4644_
timestamp 0
transform -1 0 3470 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__4645_
timestamp 0
transform -1 0 830 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4646_
timestamp 0
transform 1 0 610 0 1 10810
box -6 -8 26 248
use FILL  FILL_1__4647_
timestamp 0
transform -1 0 1230 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4648_
timestamp 0
transform -1 0 1170 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4649_
timestamp 0
transform -1 0 530 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4650_
timestamp 0
transform -1 0 770 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1__4651_
timestamp 0
transform 1 0 4070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__4652_
timestamp 0
transform 1 0 3790 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__4653_
timestamp 0
transform -1 0 4290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__4654_
timestamp 0
transform -1 0 6850 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4655_
timestamp 0
transform 1 0 2510 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4656_
timestamp 0
transform -1 0 2330 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4657_
timestamp 0
transform -1 0 2250 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4658_
timestamp 0
transform 1 0 3690 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4659_
timestamp 0
transform -1 0 3910 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4660_
timestamp 0
transform -1 0 4290 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4661_
timestamp 0
transform 1 0 4470 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4662_
timestamp 0
transform 1 0 3930 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4663_
timestamp 0
transform 1 0 3370 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4664_
timestamp 0
transform 1 0 2510 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4665_
timestamp 0
transform -1 0 7790 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4666_
timestamp 0
transform 1 0 7690 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__4667_
timestamp 0
transform 1 0 6210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__4668_
timestamp 0
transform -1 0 6430 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1__4669_
timestamp 0
transform 1 0 410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4670_
timestamp 0
transform 1 0 3990 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4671_
timestamp 0
transform 1 0 3810 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4672_
timestamp 0
transform 1 0 2750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4673_
timestamp 0
transform -1 0 2950 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4674_
timestamp 0
transform -1 0 3110 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4675_
timestamp 0
transform -1 0 2990 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4676_
timestamp 0
transform -1 0 3590 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4677_
timestamp 0
transform -1 0 3530 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4678_
timestamp 0
transform 1 0 3350 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4679_
timestamp 0
transform -1 0 3190 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4680_
timestamp 0
transform -1 0 2190 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__4681_
timestamp 0
transform 1 0 1970 0 1 2650
box -6 -8 26 248
use FILL  FILL_1__4682_
timestamp 0
transform -1 0 7030 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4683_
timestamp 0
transform -1 0 1830 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4684_
timestamp 0
transform 1 0 3730 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4685_
timestamp 0
transform 1 0 3550 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4686_
timestamp 0
transform 1 0 11090 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4687_
timestamp 0
transform 1 0 11270 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4688_
timestamp 0
transform 1 0 11450 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4689_
timestamp 0
transform 1 0 11630 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4690_
timestamp 0
transform 1 0 10470 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4691_
timestamp 0
transform 1 0 10110 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4692_
timestamp 0
transform 1 0 10190 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4693_
timestamp 0
transform -1 0 9710 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4694_
timestamp 0
transform -1 0 9730 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4695_
timestamp 0
transform 1 0 10570 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4696_
timestamp 0
transform 1 0 10890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4697_
timestamp 0
transform 1 0 11370 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4698_
timestamp 0
transform 1 0 11210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4699_
timestamp 0
transform 1 0 11210 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4700_
timestamp 0
transform 1 0 11050 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4701_
timestamp 0
transform -1 0 11430 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4702_
timestamp 0
transform 1 0 11410 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4703_
timestamp 0
transform 1 0 11690 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4704_
timestamp 0
transform -1 0 11590 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4705_
timestamp 0
transform -1 0 11790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4706_
timestamp 0
transform -1 0 11730 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4707_
timestamp 0
transform 1 0 10670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4708_
timestamp 0
transform 1 0 10870 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4709_
timestamp 0
transform -1 0 10870 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4710_
timestamp 0
transform -1 0 10670 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4711_
timestamp 0
transform 1 0 10130 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4712_
timestamp 0
transform -1 0 9910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4713_
timestamp 0
transform 1 0 9710 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4714_
timestamp 0
transform 1 0 9510 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4715_
timestamp 0
transform -1 0 9830 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4716_
timestamp 0
transform 1 0 9250 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4717_
timestamp 0
transform 1 0 9590 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4718_
timestamp 0
transform -1 0 8730 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4719_
timestamp 0
transform 1 0 11270 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4720_
timestamp 0
transform 1 0 10010 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4721_
timestamp 0
transform 1 0 9830 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4722_
timestamp 0
transform -1 0 9910 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4723_
timestamp 0
transform -1 0 9910 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4724_
timestamp 0
transform 1 0 4210 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4725_
timestamp 0
transform -1 0 10110 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4726_
timestamp 0
transform -1 0 10310 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4727_
timestamp 0
transform -1 0 11070 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4728_
timestamp 0
transform 1 0 10150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4729_
timestamp 0
transform -1 0 10090 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4730_
timestamp 0
transform -1 0 9970 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4731_
timestamp 0
transform -1 0 11650 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4732_
timestamp 0
transform -1 0 9810 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4733_
timestamp 0
transform 1 0 9790 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4734_
timestamp 0
transform -1 0 7770 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4735_
timestamp 0
transform 1 0 9310 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4736_
timestamp 0
transform -1 0 10010 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4737_
timestamp 0
transform 1 0 9510 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4738_
timestamp 0
transform -1 0 9710 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4739_
timestamp 0
transform -1 0 9890 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4740_
timestamp 0
transform -1 0 10270 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4741_
timestamp 0
transform -1 0 10090 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4742_
timestamp 0
transform 1 0 10310 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4743_
timestamp 0
transform 1 0 10070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4744_
timestamp 0
transform 1 0 10570 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4745_
timestamp 0
transform 1 0 10890 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4746_
timestamp 0
transform 1 0 10370 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4747_
timestamp 0
transform 1 0 8310 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4748_
timestamp 0
transform 1 0 8510 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4749_
timestamp 0
transform -1 0 8750 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4750_
timestamp 0
transform 1 0 8510 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4751_
timestamp 0
transform 1 0 3710 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4752_
timestamp 0
transform -1 0 9110 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4753_
timestamp 0
transform -1 0 7990 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4754_
timestamp 0
transform 1 0 8110 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4755_
timestamp 0
transform 1 0 7230 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4756_
timestamp 0
transform 1 0 6890 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4757_
timestamp 0
transform 1 0 8330 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4758_
timestamp 0
transform -1 0 10390 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4759_
timestamp 0
transform 1 0 10750 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4760_
timestamp 0
transform -1 0 11030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4761_
timestamp 0
transform 1 0 11310 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4762_
timestamp 0
transform -1 0 10470 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4763_
timestamp 0
transform 1 0 11810 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4764_
timestamp 0
transform 1 0 10850 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4765_
timestamp 0
transform -1 0 11110 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4766_
timestamp 0
transform -1 0 10470 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4767_
timestamp 0
transform -1 0 10490 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4768_
timestamp 0
transform 1 0 10270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4769_
timestamp 0
transform 1 0 10650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4770_
timestamp 0
transform 1 0 11130 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4771_
timestamp 0
transform 1 0 11990 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4772_
timestamp 0
transform 1 0 9330 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4773_
timestamp 0
transform -1 0 8790 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4774_
timestamp 0
transform 1 0 2530 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4775_
timestamp 0
transform 1 0 2690 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4776_
timestamp 0
transform 1 0 2850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4777_
timestamp 0
transform -1 0 3070 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4778_
timestamp 0
transform -1 0 3670 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4779_
timestamp 0
transform 1 0 3850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4780_
timestamp 0
transform -1 0 8730 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4781_
timestamp 0
transform 1 0 3570 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4782_
timestamp 0
transform 1 0 3250 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4783_
timestamp 0
transform 1 0 9070 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4784_
timestamp 0
transform 1 0 7710 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4785_
timestamp 0
transform 1 0 2070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4786_
timestamp 0
transform -1 0 3950 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__4787_
timestamp 0
transform -1 0 3630 0 1 3130
box -6 -8 26 248
use FILL  FILL_1__4788_
timestamp 0
transform -1 0 4150 0 1 3610
box -6 -8 26 248
use FILL  FILL_1__4789_
timestamp 0
transform 1 0 7190 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4790_
timestamp 0
transform 1 0 7250 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4791_
timestamp 0
transform -1 0 7790 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4792_
timestamp 0
transform -1 0 7850 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4793_
timestamp 0
transform -1 0 7790 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4794_
timestamp 0
transform -1 0 7430 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4795_
timestamp 0
transform -1 0 7490 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4796_
timestamp 0
transform 1 0 11790 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4797_
timestamp 0
transform 1 0 8530 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4798_
timestamp 0
transform 1 0 9990 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4799_
timestamp 0
transform -1 0 9830 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4800_
timestamp 0
transform 1 0 8470 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4801_
timestamp 0
transform 1 0 10930 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4802_
timestamp 0
transform -1 0 10470 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4803_
timestamp 0
transform -1 0 7370 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4804_
timestamp 0
transform -1 0 7050 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4805_
timestamp 0
transform -1 0 6930 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4806_
timestamp 0
transform -1 0 9290 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4807_
timestamp 0
transform -1 0 9070 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4808_
timestamp 0
transform -1 0 8690 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4809_
timestamp 0
transform -1 0 8690 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4810_
timestamp 0
transform -1 0 8930 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4811_
timestamp 0
transform 1 0 11910 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4812_
timestamp 0
transform 1 0 11990 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4813_
timestamp 0
transform 1 0 11450 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4814_
timestamp 0
transform 1 0 11330 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4815_
timestamp 0
transform -1 0 9030 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4816_
timestamp 0
transform -1 0 9470 0 1 7450
box -6 -8 26 248
use FILL  FILL_1__4817_
timestamp 0
transform -1 0 11530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4818_
timestamp 0
transform -1 0 11470 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4819_
timestamp 0
transform -1 0 6410 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4820_
timestamp 0
transform 1 0 7970 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4821_
timestamp 0
transform 1 0 11610 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4822_
timestamp 0
transform 1 0 11810 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4823_
timestamp 0
transform 1 0 11590 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4824_
timestamp 0
transform -1 0 11450 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4825_
timestamp 0
transform 1 0 11150 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4826_
timestamp 0
transform -1 0 10990 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4827_
timestamp 0
transform -1 0 11690 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4828_
timestamp 0
transform -1 0 11770 0 1 10330
box -6 -8 26 248
use FILL  FILL_1__4829_
timestamp 0
transform 1 0 11610 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4830_
timestamp 0
transform 1 0 8970 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4831_
timestamp 0
transform -1 0 9330 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4832_
timestamp 0
transform 1 0 11870 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4833_
timestamp 0
transform 1 0 8350 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4834_
timestamp 0
transform 1 0 8150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4835_
timestamp 0
transform -1 0 8350 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4836_
timestamp 0
transform 1 0 9630 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4837_
timestamp 0
transform -1 0 10770 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4838_
timestamp 0
transform 1 0 11790 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4839_
timestamp 0
transform 1 0 12050 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4840_
timestamp 0
transform 1 0 9230 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4841_
timestamp 0
transform 1 0 10270 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4842_
timestamp 0
transform 1 0 11970 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4843_
timestamp 0
transform 1 0 11130 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4844_
timestamp 0
transform -1 0 11110 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4845_
timestamp 0
transform -1 0 11890 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4846_
timestamp 0
transform 1 0 11870 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4847_
timestamp 0
transform -1 0 8350 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1__4848_
timestamp 0
transform -1 0 8370 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4849_
timestamp 0
transform 1 0 9030 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4850_
timestamp 0
transform 1 0 9270 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4851_
timestamp 0
transform 1 0 11250 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4852_
timestamp 0
transform 1 0 11630 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4853_
timestamp 0
transform 1 0 12030 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4854_
timestamp 0
transform -1 0 11170 0 1 11770
box -6 -8 26 248
use FILL  FILL_1__4855_
timestamp 0
transform -1 0 8190 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4856_
timestamp 0
transform -1 0 8210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4857_
timestamp 0
transform -1 0 10290 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4858_
timestamp 0
transform -1 0 10430 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4859_
timestamp 0
transform -1 0 7170 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4860_
timestamp 0
transform -1 0 10350 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4861_
timestamp 0
transform -1 0 10610 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4862_
timestamp 0
transform 1 0 11410 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4863_
timestamp 0
transform -1 0 10670 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4864_
timestamp 0
transform -1 0 10510 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4865_
timestamp 0
transform 1 0 10530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4866_
timestamp 0
transform 1 0 11610 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4867_
timestamp 0
transform 1 0 11790 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4868_
timestamp 0
transform -1 0 11290 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4869_
timestamp 0
transform -1 0 10830 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1__4870_
timestamp 0
transform 1 0 8070 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4871_
timestamp 0
transform 1 0 7910 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4872_
timestamp 0
transform 1 0 7810 0 1 7930
box -6 -8 26 248
use FILL  FILL_1__4873_
timestamp 0
transform -1 0 11330 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4874_
timestamp 0
transform 1 0 11850 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4875_
timestamp 0
transform -1 0 7550 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1__4876_
timestamp 0
transform -1 0 10470 0 -1 9370
box -6 -8 26 248
use FILL  FILL_1__4877_
timestamp 0
transform 1 0 10870 0 1 8410
box -6 -8 26 248
use FILL  FILL_1__4878_
timestamp 0
transform 1 0 11310 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4879_
timestamp 0
transform 1 0 11970 0 1 9850
box -6 -8 26 248
use FILL  FILL_1__4880_
timestamp 0
transform -1 0 12030 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4881_
timestamp 0
transform -1 0 9070 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4882_
timestamp 0
transform 1 0 11990 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4883_
timestamp 0
transform 1 0 11810 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4884_
timestamp 0
transform 1 0 11630 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4885_
timestamp 0
transform -1 0 11670 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4886_
timestamp 0
transform 1 0 10930 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4887_
timestamp 0
transform 1 0 10970 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4888_
timestamp 0
transform 1 0 11630 0 1 8890
box -6 -8 26 248
use FILL  FILL_1__4889_
timestamp 0
transform 1 0 11970 0 1 9370
box -6 -8 26 248
use FILL  FILL_1__4890_
timestamp 0
transform 1 0 11490 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4891_
timestamp 0
transform 1 0 11830 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1__4892_
timestamp 0
transform -1 0 12050 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1__4893_
timestamp 0
transform -1 0 2470 0 -1 7450
box -6 -8 26 248
use FILL  FILL_1__4894_
timestamp 0
transform 1 0 9670 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4895_
timestamp 0
transform 1 0 8410 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4896_
timestamp 0
transform -1 0 9450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4897_
timestamp 0
transform 1 0 9490 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4898_
timestamp 0
transform 1 0 9670 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4899_
timestamp 0
transform -1 0 9150 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4900_
timestamp 0
transform -1 0 9490 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4901_
timestamp 0
transform -1 0 9870 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4902_
timestamp 0
transform 1 0 10190 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4903_
timestamp 0
transform 1 0 9650 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4904_
timestamp 0
transform -1 0 10370 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4905_
timestamp 0
transform 1 0 9650 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4906_
timestamp 0
transform -1 0 9830 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4907_
timestamp 0
transform -1 0 9490 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4908_
timestamp 0
transform 1 0 9990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4909_
timestamp 0
transform 1 0 10930 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4910_
timestamp 0
transform -1 0 11310 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4911_
timestamp 0
transform 1 0 11250 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4912_
timestamp 0
transform 1 0 11070 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4913_
timestamp 0
transform -1 0 10890 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4914_
timestamp 0
transform 1 0 11450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4915_
timestamp 0
transform -1 0 10750 0 1 6970
box -6 -8 26 248
use FILL  FILL_1__4916_
timestamp 0
transform 1 0 10510 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4917_
timestamp 0
transform -1 0 10570 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4918_
timestamp 0
transform -1 0 10930 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4919_
timestamp 0
transform 1 0 11090 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4920_
timestamp 0
transform 1 0 8510 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4921_
timestamp 0
transform -1 0 8730 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4922_
timestamp 0
transform -1 0 8930 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4923_
timestamp 0
transform 1 0 9310 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4924_
timestamp 0
transform 1 0 9290 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4925_
timestamp 0
transform -1 0 9110 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4926_
timestamp 0
transform 1 0 8870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4927_
timestamp 0
transform -1 0 11270 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4928_
timestamp 0
transform 1 0 11450 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4929_
timestamp 0
transform 1 0 12030 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4930_
timestamp 0
transform 1 0 11610 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4931_
timestamp 0
transform -1 0 11830 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4932_
timestamp 0
transform -1 0 11670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4933_
timestamp 0
transform -1 0 11110 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4934_
timestamp 0
transform 1 0 10890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4935_
timestamp 0
transform -1 0 10710 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4936_
timestamp 0
transform -1 0 9610 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4937_
timestamp 0
transform -1 0 9830 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4938_
timestamp 0
transform 1 0 9990 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4939_
timestamp 0
transform 1 0 10070 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4940_
timestamp 0
transform 1 0 10170 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1__4941_
timestamp 0
transform 1 0 10270 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4942_
timestamp 0
transform -1 0 10670 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4943_
timestamp 0
transform 1 0 11650 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4944_
timestamp 0
transform -1 0 11870 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4945_
timestamp 0
transform 1 0 11810 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4946_
timestamp 0
transform -1 0 11790 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4947_
timestamp 0
transform -1 0 8610 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4948_
timestamp 0
transform 1 0 8930 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4949_
timestamp 0
transform 1 0 12050 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__4950_
timestamp 0
transform -1 0 12010 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4951_
timestamp 0
transform -1 0 8550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4952_
timestamp 0
transform 1 0 8930 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4953_
timestamp 0
transform -1 0 8830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4954_
timestamp 0
transform -1 0 9130 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4955_
timestamp 0
transform -1 0 8690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__4956_
timestamp 0
transform -1 0 8770 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4957_
timestamp 0
transform -1 0 8630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4958_
timestamp 0
transform -1 0 11010 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4959_
timestamp 0
transform 1 0 11190 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4960_
timestamp 0
transform -1 0 11410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4961_
timestamp 0
transform 1 0 11590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4962_
timestamp 0
transform 1 0 11990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4963_
timestamp 0
transform 1 0 11950 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4964_
timestamp 0
transform 1 0 11950 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4965_
timestamp 0
transform -1 0 11790 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4966_
timestamp 0
transform -1 0 9130 0 1 4090
box -6 -8 26 248
use FILL  FILL_1__4967_
timestamp 0
transform 1 0 8050 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__4968_
timestamp 0
transform 1 0 11630 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4969_
timestamp 0
transform 1 0 11990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4970_
timestamp 0
transform 1 0 9030 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4971_
timestamp 0
transform -1 0 8250 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4972_
timestamp 0
transform -1 0 8650 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4973_
timestamp 0
transform -1 0 8810 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4974_
timestamp 0
transform 1 0 8710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4975_
timestamp 0
transform 1 0 8910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4976_
timestamp 0
transform 1 0 11570 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4977_
timestamp 0
transform 1 0 11370 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4978_
timestamp 0
transform 1 0 11390 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4979_
timestamp 0
transform 1 0 11410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4980_
timestamp 0
transform 1 0 11790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4981_
timestamp 0
transform -1 0 11790 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4982_
timestamp 0
transform -1 0 11810 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4983_
timestamp 0
transform 1 0 11590 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4984_
timestamp 0
transform 1 0 11210 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4985_
timestamp 0
transform -1 0 8030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4986_
timestamp 0
transform 1 0 9070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4987_
timestamp 0
transform 1 0 11590 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4988_
timestamp 0
transform -1 0 11810 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4989_
timestamp 0
transform -1 0 11410 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4990_
timestamp 0
transform -1 0 11230 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__4991_
timestamp 0
transform 1 0 11610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__4992_
timestamp 0
transform -1 0 11470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4993_
timestamp 0
transform 1 0 11250 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__4994_
timestamp 0
transform 1 0 9270 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__4995_
timestamp 0
transform -1 0 9850 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4996_
timestamp 0
transform 1 0 9210 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4997_
timestamp 0
transform -1 0 9290 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__4998_
timestamp 0
transform 1 0 9390 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__4999_
timestamp 0
transform -1 0 9250 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5000_
timestamp 0
transform 1 0 10990 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__5001_
timestamp 0
transform -1 0 10810 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__5002_
timestamp 0
transform -1 0 10630 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5003_
timestamp 0
transform -1 0 10690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5004_
timestamp 0
transform 1 0 10870 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5005_
timestamp 0
transform -1 0 10850 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5006_
timestamp 0
transform 1 0 11370 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5007_
timestamp 0
transform 1 0 11970 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5008_
timestamp 0
transform 1 0 11950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__5009_
timestamp 0
transform 1 0 11970 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5010_
timestamp 0
transform -1 0 11270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__5011_
timestamp 0
transform 1 0 11770 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5012_
timestamp 0
transform 1 0 11570 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5013_
timestamp 0
transform -1 0 10250 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5014_
timestamp 0
transform -1 0 9470 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5015_
timestamp 0
transform 1 0 8230 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5016_
timestamp 0
transform 1 0 10630 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5017_
timestamp 0
transform 1 0 8890 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5018_
timestamp 0
transform 1 0 8430 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5019_
timestamp 0
transform 1 0 9110 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5020_
timestamp 0
transform 1 0 9010 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5021_
timestamp 0
transform 1 0 9290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5022_
timestamp 0
transform -1 0 9090 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5023_
timestamp 0
transform -1 0 10810 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__5024_
timestamp 0
transform 1 0 10810 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5025_
timestamp 0
transform -1 0 11030 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5026_
timestamp 0
transform 1 0 11050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__5027_
timestamp 0
transform -1 0 10850 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5028_
timestamp 0
transform -1 0 10670 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5029_
timestamp 0
transform 1 0 11010 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5030_
timestamp 0
transform 1 0 11030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5031_
timestamp 0
transform 1 0 11790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__5032_
timestamp 0
transform 1 0 11630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__5033_
timestamp 0
transform -1 0 8950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__5034_
timestamp 0
transform -1 0 9150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__5035_
timestamp 0
transform 1 0 11170 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5036_
timestamp 0
transform 1 0 9850 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5037_
timestamp 0
transform 1 0 9650 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5038_
timestamp 0
transform 1 0 9490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5039_
timestamp 0
transform 1 0 9430 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5040_
timestamp 0
transform 1 0 9670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5041_
timestamp 0
transform 1 0 9870 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5042_
timestamp 0
transform 1 0 10590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__5043_
timestamp 0
transform 1 0 10410 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5044_
timestamp 0
transform 1 0 10470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5045_
timestamp 0
transform -1 0 10450 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5046_
timestamp 0
transform 1 0 10890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__5047_
timestamp 0
transform 1 0 10990 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5048_
timestamp 0
transform 1 0 11430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__5049_
timestamp 0
transform -1 0 11270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__5050_
timestamp 0
transform -1 0 9330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__5051_
timestamp 0
transform 1 0 8330 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__5052_
timestamp 0
transform -1 0 10490 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__5053_
timestamp 0
transform -1 0 10730 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__5054_
timestamp 0
transform -1 0 10370 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__5055_
timestamp 0
transform 1 0 8490 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__5056_
timestamp 0
transform 1 0 8110 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__5057_
timestamp 0
transform 1 0 8330 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__5058_
timestamp 0
transform -1 0 8150 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__5059_
timestamp 0
transform 1 0 7970 0 1 6490
box -6 -8 26 248
use FILL  FILL_1__5060_
timestamp 0
transform -1 0 7610 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__5061_
timestamp 0
transform -1 0 7790 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__5062_
timestamp 0
transform 1 0 7950 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1__5063_
timestamp 0
transform -1 0 7990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__5064_
timestamp 0
transform -1 0 7510 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5065_
timestamp 0
transform -1 0 7710 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5066_
timestamp 0
transform -1 0 7650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5067_
timestamp 0
transform -1 0 8350 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5068_
timestamp 0
transform -1 0 8370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5069_
timestamp 0
transform -1 0 8210 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5070_
timestamp 0
transform -1 0 7830 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5071_
timestamp 0
transform 1 0 8010 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5072_
timestamp 0
transform -1 0 7470 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5073_
timestamp 0
transform 1 0 7270 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5074_
timestamp 0
transform 1 0 4830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1__5075_
timestamp 0
transform 1 0 10230 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__5076_
timestamp 0
transform 1 0 10030 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__5077_
timestamp 0
transform 1 0 9810 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__5078_
timestamp 0
transform 1 0 9590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__5079_
timestamp 0
transform 1 0 9990 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__5080_
timestamp 0
transform 1 0 10190 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__5081_
timestamp 0
transform 1 0 10410 0 1 6010
box -6 -8 26 248
use FILL  FILL_1__5082_
timestamp 0
transform 1 0 10390 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1__5083_
timestamp 0
transform -1 0 10290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5084_
timestamp 0
transform -1 0 9670 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5085_
timestamp 0
transform 1 0 8510 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5086_
timestamp 0
transform -1 0 8710 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5087_
timestamp 0
transform -1 0 10870 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__5088_
timestamp 0
transform -1 0 10650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__5089_
timestamp 0
transform -1 0 10450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__5090_
timestamp 0
transform -1 0 10230 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5091_
timestamp 0
transform 1 0 10070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1__5092_
timestamp 0
transform 1 0 9910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__5093_
timestamp 0
transform -1 0 10090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__5094_
timestamp 0
transform 1 0 10230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__5095_
timestamp 0
transform -1 0 9750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__5096_
timestamp 0
transform 1 0 8890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__5097_
timestamp 0
transform 1 0 8210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1__5098_
timestamp 0
transform 1 0 9710 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5099_
timestamp 0
transform 1 0 9890 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5100_
timestamp 0
transform 1 0 9330 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5101_
timestamp 0
transform -1 0 10050 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5102_
timestamp 0
transform -1 0 9870 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5103_
timestamp 0
transform 1 0 10010 0 1 5050
box -6 -8 26 248
use FILL  FILL_1__5104_
timestamp 0
transform -1 0 10310 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5105_
timestamp 0
transform -1 0 10110 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5106_
timestamp 0
transform -1 0 10490 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5107_
timestamp 0
transform 1 0 10470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__5108_
timestamp 0
transform -1 0 11070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__5109_
timestamp 0
transform 1 0 10670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1__5110_
timestamp 0
transform -1 0 9530 0 1 4570
box -6 -8 26 248
use FILL  FILL_1__5111_
timestamp 0
transform -1 0 7890 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5112_
timestamp 0
transform -1 0 8070 0 1 5530
box -6 -8 26 248
use FILL  FILL_1__5124_
timestamp 0
transform 1 0 1750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__5125_
timestamp 0
transform -1 0 610 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__5126_
timestamp 0
transform -1 0 790 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__5127_
timestamp 0
transform 1 0 750 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__5128_
timestamp 0
transform 1 0 510 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__5129_
timestamp 0
transform 1 0 950 0 1 2170
box -6 -8 26 248
use FILL  FILL_1__5130_
timestamp 0
transform 1 0 950 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__5131_
timestamp 0
transform -1 0 2270 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5132_
timestamp 0
transform -1 0 5510 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5133_
timestamp 0
transform 1 0 5250 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5134_
timestamp 0
transform 1 0 1330 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__5135_
timestamp 0
transform 1 0 2130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__5136_
timestamp 0
transform 1 0 1930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__5137_
timestamp 0
transform -1 0 1070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__5138_
timestamp 0
transform -1 0 1250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__5139_
timestamp 0
transform -1 0 3630 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5140_
timestamp 0
transform 1 0 4090 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__5141_
timestamp 0
transform -1 0 4270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__5142_
timestamp 0
transform -1 0 4150 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__5143_
timestamp 0
transform -1 0 4370 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5144_
timestamp 0
transform 1 0 5530 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5145_
timestamp 0
transform -1 0 4070 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5146_
timestamp 0
transform -1 0 4590 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5147_
timestamp 0
transform 1 0 4690 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5148_
timestamp 0
transform 1 0 4890 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5149_
timestamp 0
transform 1 0 5410 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5150_
timestamp 0
transform -1 0 6030 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5151_
timestamp 0
transform 1 0 3410 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5152_
timestamp 0
transform 1 0 5670 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5153_
timestamp 0
transform 1 0 4150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__5154_
timestamp 0
transform 1 0 5350 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5155_
timestamp 0
transform 1 0 5310 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5156_
timestamp 0
transform 1 0 5470 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5157_
timestamp 0
transform 1 0 5610 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5158_
timestamp 0
transform 1 0 4490 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5159_
timestamp 0
transform -1 0 4610 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5160_
timestamp 0
transform 1 0 4930 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5161_
timestamp 0
transform 1 0 4770 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5162_
timestamp 0
transform 1 0 5810 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5163_
timestamp 0
transform -1 0 2710 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5164_
timestamp 0
transform 1 0 5830 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5165_
timestamp 0
transform -1 0 3770 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__5166_
timestamp 0
transform 1 0 4210 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5167_
timestamp 0
transform 1 0 4170 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5168_
timestamp 0
transform -1 0 3990 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5169_
timestamp 0
transform 1 0 2670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__5170_
timestamp 0
transform 1 0 3790 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5171_
timestamp 0
transform -1 0 4090 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__5172_
timestamp 0
transform -1 0 3590 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__5173_
timestamp 0
transform -1 0 4870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__5174_
timestamp 0
transform -1 0 3770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__5175_
timestamp 0
transform 1 0 3610 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5176_
timestamp 0
transform -1 0 2610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__5177_
timestamp 0
transform 1 0 3050 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5178_
timestamp 0
transform 1 0 4390 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5179_
timestamp 0
transform 1 0 4410 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5180_
timestamp 0
transform 1 0 4210 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5181_
timestamp 0
transform 1 0 3210 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5182_
timestamp 0
transform -1 0 2410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__5183_
timestamp 0
transform 1 0 2210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__5184_
timestamp 0
transform -1 0 2430 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__5185_
timestamp 0
transform -1 0 3990 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__5186_
timestamp 0
transform -1 0 3270 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__5187_
timestamp 0
transform -1 0 3010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__5188_
timestamp 0
transform 1 0 3710 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5189_
timestamp 0
transform -1 0 3650 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5190_
timestamp 0
transform 1 0 3190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__5191_
timestamp 0
transform 1 0 2870 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5192_
timestamp 0
transform -1 0 3590 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__5193_
timestamp 0
transform 1 0 6030 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5194_
timestamp 0
transform -1 0 2890 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__5195_
timestamp 0
transform -1 0 2810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__5196_
timestamp 0
transform 1 0 3550 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5197_
timestamp 0
transform -1 0 3470 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5198_
timestamp 0
transform -1 0 2870 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5199_
timestamp 0
transform 1 0 2430 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5200_
timestamp 0
transform -1 0 2650 0 -1 730
box -6 -8 26 248
use FILL  FILL_1__5201_
timestamp 0
transform -1 0 3930 0 1 1690
box -6 -8 26 248
use FILL  FILL_1__5202_
timestamp 0
transform 1 0 3890 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5203_
timestamp 0
transform -1 0 3430 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5204_
timestamp 0
transform 1 0 4050 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5205_
timestamp 0
transform -1 0 3890 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5206_
timestamp 0
transform -1 0 3230 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5207_
timestamp 0
transform 1 0 2450 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5208_
timestamp 0
transform 1 0 2990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__5209_
timestamp 0
transform -1 0 4450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1__5210_
timestamp 0
transform 1 0 2650 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5211_
timestamp 0
transform 1 0 2810 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5212_
timestamp 0
transform 1 0 3390 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5213_
timestamp 0
transform 1 0 3270 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5214_
timestamp 0
transform -1 0 3030 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5215_
timestamp 0
transform 1 0 2250 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5216_
timestamp 0
transform -1 0 3050 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__5217_
timestamp 0
transform -1 0 6210 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5218_
timestamp 0
transform 1 0 3390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__5219_
timestamp 0
transform 1 0 3550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__5220_
timestamp 0
transform 1 0 4730 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5221_
timestamp 0
transform 1 0 4550 0 -1 250
box -6 -8 26 248
use FILL  FILL_1__5222_
timestamp 0
transform -1 0 4030 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5223_
timestamp 0
transform 1 0 3070 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5224_
timestamp 0
transform -1 0 3830 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5225_
timestamp 0
transform 1 0 5330 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__5226_
timestamp 0
transform 1 0 5110 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5227_
timestamp 0
transform -1 0 5290 0 1 250
box -6 -8 26 248
use FILL  FILL_1__5228_
timestamp 0
transform -1 0 4730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1__5229_
timestamp 0
transform -1 0 4770 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5230_
timestamp 0
transform 1 0 4950 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5231_
timestamp 0
transform 1 0 5150 0 1 730
box -6 -8 26 248
use FILL  FILL_1__5232_
timestamp 0
transform 1 0 3950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1__5233_
timestamp 0
transform 1 0 4330 0 1 1210
box -6 -8 26 248
use FILL  FILL_1__5234_
timestamp 0
transform -1 0 5130 0 1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert0
timestamp 0
transform -1 0 4170 0 1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert1
timestamp 0
transform 1 0 6090 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert2
timestamp 0
transform -1 0 3270 0 1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert3
timestamp 0
transform -1 0 3650 0 1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert4
timestamp 0
transform 1 0 9430 0 1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert5
timestamp 0
transform 1 0 11230 0 1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert6
timestamp 0
transform -1 0 9430 0 1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert7
timestamp 0
transform 1 0 11970 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert8
timestamp 0
transform -1 0 7130 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert9
timestamp 0
transform 1 0 6630 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert10
timestamp 0
transform 1 0 8670 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert11
timestamp 0
transform 1 0 6830 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert12
timestamp 0
transform 1 0 8870 0 1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert13
timestamp 0
transform 1 0 7350 0 1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert14
timestamp 0
transform 1 0 610 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert15
timestamp 0
transform 1 0 30 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert16
timestamp 0
transform 1 0 1850 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert17
timestamp 0
transform -1 0 9110 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert18
timestamp 0
transform -1 0 11470 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert19
timestamp 0
transform 1 0 10630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert20
timestamp 0
transform -1 0 9150 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert21
timestamp 0
transform 1 0 2490 0 1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert22
timestamp 0
transform -1 0 1230 0 1 11290
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert23
timestamp 0
transform -1 0 1410 0 1 11290
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert24
timestamp 0
transform -1 0 1610 0 1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert38
timestamp 0
transform -1 0 11490 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert39
timestamp 0
transform -1 0 10630 0 1 6010
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert40
timestamp 0
transform 1 0 11990 0 1 6970
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert41
timestamp 0
transform -1 0 11210 0 1 6010
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert42
timestamp 0
transform 1 0 11410 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert43
timestamp 0
transform -1 0 10970 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert44
timestamp 0
transform -1 0 10450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert45
timestamp 0
transform -1 0 11330 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert46
timestamp 0
transform -1 0 10710 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert47
timestamp 0
transform 1 0 6170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert48
timestamp 0
transform -1 0 4730 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert49
timestamp 0
transform 1 0 11530 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert50
timestamp 0
transform -1 0 10370 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert51
timestamp 0
transform 1 0 8130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert52
timestamp 0
transform 1 0 9990 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert53
timestamp 0
transform 1 0 9150 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert54
timestamp 0
transform 1 0 8970 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert55
timestamp 0
transform -1 0 9510 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert56
timestamp 0
transform -1 0 8810 0 1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert57
timestamp 0
transform 1 0 11430 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert58
timestamp 0
transform 1 0 10610 0 -1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert59
timestamp 0
transform -1 0 7690 0 -1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert60
timestamp 0
transform 1 0 11770 0 -1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert61
timestamp 0
transform 1 0 11870 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert62
timestamp 0
transform -1 0 4770 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert63
timestamp 0
transform -1 0 9290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert64
timestamp 0
transform -1 0 11630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert65
timestamp 0
transform -1 0 9290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert66
timestamp 0
transform -1 0 11470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert67
timestamp 0
transform 1 0 6890 0 1 11290
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert68
timestamp 0
transform -1 0 3130 0 -1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert69
timestamp 0
transform -1 0 5590 0 1 10810
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert70
timestamp 0
transform 1 0 5070 0 -1 11290
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert71
timestamp 0
transform -1 0 3530 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert72
timestamp 0
transform 1 0 7070 0 1 11290
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert73
timestamp 0
transform 1 0 7090 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert74
timestamp 0
transform -1 0 6430 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert75
timestamp 0
transform 1 0 7050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert76
timestamp 0
transform 1 0 6510 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert77
timestamp 0
transform 1 0 10230 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert78
timestamp 0
transform 1 0 9090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert79
timestamp 0
transform 1 0 10250 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert80
timestamp 0
transform -1 0 4910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert81
timestamp 0
transform -1 0 2770 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert82
timestamp 0
transform -1 0 3990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert83
timestamp 0
transform -1 0 6250 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert84
timestamp 0
transform 1 0 7310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert85
timestamp 0
transform -1 0 3230 0 1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert86
timestamp 0
transform 1 0 3930 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert87
timestamp 0
transform -1 0 3190 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert88
timestamp 0
transform 1 0 7850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert89
timestamp 0
transform -1 0 4690 0 1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert90
timestamp 0
transform 1 0 5530 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert91
timestamp 0
transform 1 0 8990 0 1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert92
timestamp 0
transform -1 0 8490 0 1 10810
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert93
timestamp 0
transform -1 0 10890 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert94
timestamp 0
transform 1 0 7230 0 1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert95
timestamp 0
transform 1 0 11490 0 1 10810
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert96
timestamp 0
transform -1 0 4950 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert97
timestamp 0
transform 1 0 570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert98
timestamp 0
transform -1 0 3970 0 1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert99
timestamp 0
transform 1 0 510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert100
timestamp 0
transform 1 0 2990 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert101
timestamp 0
transform -1 0 450 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert102
timestamp 0
transform 1 0 3690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert103
timestamp 0
transform -1 0 3610 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert104
timestamp 0
transform 1 0 4590 0 1 10330
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert105
timestamp 0
transform 1 0 250 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert106
timestamp 0
transform 1 0 6470 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert107
timestamp 0
transform -1 0 6170 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert108
timestamp 0
transform 1 0 5650 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert109
timestamp 0
transform 1 0 7790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert110
timestamp 0
transform -1 0 5290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert111
timestamp 0
transform 1 0 7250 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert112
timestamp 0
transform 1 0 10630 0 1 11770
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert113
timestamp 0
transform -1 0 12070 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert114
timestamp 0
transform -1 0 10270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert115
timestamp 0
transform 1 0 7330 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert116
timestamp 0
transform -1 0 5470 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert117
timestamp 0
transform -1 0 5450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert118
timestamp 0
transform -1 0 11150 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert119
timestamp 0
transform 1 0 10330 0 1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert120
timestamp 0
transform -1 0 11070 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert121
timestamp 0
transform -1 0 8130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert122
timestamp 0
transform 1 0 11150 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert123
timestamp 0
transform -1 0 9990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert124
timestamp 0
transform -1 0 7970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert125
timestamp 0
transform -1 0 5290 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert126
timestamp 0
transform 1 0 11970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert127
timestamp 0
transform 1 0 10730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert128
timestamp 0
transform -1 0 12010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert129
timestamp 0
transform 1 0 10410 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert130
timestamp 0
transform 1 0 11970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert131
timestamp 0
transform -1 0 9330 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert132
timestamp 0
transform -1 0 8670 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert133
timestamp 0
transform 1 0 11970 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert134
timestamp 0
transform -1 0 11350 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert135
timestamp 0
transform -1 0 9070 0 -1 250
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert136
timestamp 0
transform 1 0 9430 0 -1 250
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert137
timestamp 0
transform -1 0 6350 0 1 730
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert138
timestamp 0
transform 1 0 8330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert139
timestamp 0
transform -1 0 6370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert140
timestamp 0
transform 1 0 9390 0 1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert141
timestamp 0
transform -1 0 7010 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert142
timestamp 0
transform -1 0 6990 0 1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert143
timestamp 0
transform -1 0 6410 0 -1 6970
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert144
timestamp 0
transform -1 0 6230 0 1 6970
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert145
timestamp 0
transform 1 0 9510 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert146
timestamp 0
transform 1 0 9610 0 1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert147
timestamp 0
transform -1 0 7690 0 1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert148
timestamp 0
transform -1 0 7610 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert149
timestamp 0
transform -1 0 9190 0 -1 7930
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert150
timestamp 0
transform -1 0 7190 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert151
timestamp 0
transform 1 0 7290 0 -1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert152
timestamp 0
transform -1 0 8190 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert153
timestamp 0
transform 1 0 10030 0 -1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert154
timestamp 0
transform 1 0 10710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert155
timestamp 0
transform 1 0 6350 0 1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert156
timestamp 0
transform 1 0 9090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert157
timestamp 0
transform -1 0 5830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert158
timestamp 0
transform 1 0 9830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert159
timestamp 0
transform 1 0 8690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert160
timestamp 0
transform 1 0 10330 0 1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert161
timestamp 0
transform 1 0 9230 0 1 9850
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert162
timestamp 0
transform 1 0 10190 0 1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert163
timestamp 0
transform -1 0 8290 0 1 8890
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert164
timestamp 0
transform 1 0 11690 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert165
timestamp 0
transform -1 0 8750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert166
timestamp 0
transform -1 0 11530 0 1 4090
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert167
timestamp 0
transform 1 0 11690 0 1 11770
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert168
timestamp 0
transform -1 0 11270 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_BUFX2_insert169
timestamp 0
transform 1 0 4890 0 1 1690
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert25
timestamp 0
transform 1 0 1330 0 1 2170
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert26
timestamp 0
transform 1 0 3990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert27
timestamp 0
transform -1 0 50 0 -1 2650
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert28
timestamp 0
transform -1 0 2690 0 1 9370
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert29
timestamp 0
transform 1 0 30 0 -1 2170
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert30
timestamp 0
transform 1 0 6150 0 -1 5050
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert31
timestamp 0
transform 1 0 750 0 -1 6010
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert32
timestamp 0
transform -1 0 4790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert33
timestamp 0
transform -1 0 930 0 -1 10810
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert34
timestamp 0
transform 1 0 1370 0 -1 6490
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert35
timestamp 0
transform -1 0 290 0 -1 11770
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert36
timestamp 0
transform 1 0 30 0 1 5530
box -6 -8 26 248
use FILL  FILL_1_CLKBUF1_insert37
timestamp 0
transform 1 0 6110 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__2478_
timestamp 0
transform -1 0 70 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2479_
timestamp 0
transform -1 0 70 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2480_
timestamp 0
transform 1 0 1910 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2481_
timestamp 0
transform 1 0 2730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2482_
timestamp 0
transform -1 0 70 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__2483_
timestamp 0
transform -1 0 550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__2484_
timestamp 0
transform -1 0 2110 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2485_
timestamp 0
transform 1 0 3930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2486_
timestamp 0
transform 1 0 12050 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2487_
timestamp 0
transform -1 0 6630 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2488_
timestamp 0
transform -1 0 6810 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2489_
timestamp 0
transform 1 0 12010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2490_
timestamp 0
transform 1 0 12010 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2491_
timestamp 0
transform 1 0 6430 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2492_
timestamp 0
transform 1 0 11830 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2493_
timestamp 0
transform -1 0 11930 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2494_
timestamp 0
transform -1 0 1030 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__2495_
timestamp 0
transform -1 0 1190 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2496_
timestamp 0
transform -1 0 70 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__2497_
timestamp 0
transform -1 0 4410 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2498_
timestamp 0
transform 1 0 4450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2499_
timestamp 0
transform -1 0 3270 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2500_
timestamp 0
transform -1 0 450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2501_
timestamp 0
transform -1 0 3650 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2502_
timestamp 0
transform -1 0 70 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__2503_
timestamp 0
transform -1 0 70 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2504_
timestamp 0
transform 1 0 4550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2505_
timestamp 0
transform 1 0 5090 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2506_
timestamp 0
transform -1 0 2530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2507_
timestamp 0
transform 1 0 3810 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2508_
timestamp 0
transform 1 0 3430 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2509_
timestamp 0
transform 1 0 4210 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2510_
timestamp 0
transform 1 0 3070 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2511_
timestamp 0
transform -1 0 4930 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2519_
timestamp 0
transform -1 0 5670 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2520_
timestamp 0
transform -1 0 7530 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2521_
timestamp 0
transform -1 0 7730 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2522_
timestamp 0
transform 1 0 7730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2523_
timestamp 0
transform 1 0 9470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2524_
timestamp 0
transform -1 0 7790 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2525_
timestamp 0
transform 1 0 7530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2526_
timestamp 0
transform 1 0 8270 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2527_
timestamp 0
transform 1 0 8470 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2528_
timestamp 0
transform -1 0 9610 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2529_
timestamp 0
transform 1 0 8550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2530_
timestamp 0
transform -1 0 8190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2531_
timestamp 0
transform -1 0 8330 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2532_
timestamp 0
transform -1 0 8750 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2533_
timestamp 0
transform 1 0 9490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2534_
timestamp 0
transform 1 0 10050 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__2535_
timestamp 0
transform -1 0 10250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2536_
timestamp 0
transform -1 0 8750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2537_
timestamp 0
transform -1 0 8550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2538_
timestamp 0
transform -1 0 8350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2539_
timestamp 0
transform 1 0 7950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2540_
timestamp 0
transform -1 0 10650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2541_
timestamp 0
transform -1 0 10850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2542_
timestamp 0
transform 1 0 10890 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2543_
timestamp 0
transform -1 0 10590 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2544_
timestamp 0
transform -1 0 5690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2545_
timestamp 0
transform -1 0 5890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2546_
timestamp 0
transform -1 0 6110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2547_
timestamp 0
transform -1 0 5990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2548_
timestamp 0
transform -1 0 6190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2549_
timestamp 0
transform 1 0 5570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2550_
timestamp 0
transform 1 0 5770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2551_
timestamp 0
transform -1 0 6890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2552_
timestamp 0
transform -1 0 7250 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2553_
timestamp 0
transform -1 0 5710 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2554_
timestamp 0
transform -1 0 6350 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2555_
timestamp 0
transform 1 0 6390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2556_
timestamp 0
transform -1 0 6730 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2557_
timestamp 0
transform -1 0 6210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2558_
timestamp 0
transform 1 0 6490 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2559_
timestamp 0
transform 1 0 6870 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2560_
timestamp 0
transform -1 0 5910 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2561_
timestamp 0
transform -1 0 6550 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2562_
timestamp 0
transform 1 0 6730 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2563_
timestamp 0
transform -1 0 6110 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2564_
timestamp 0
transform 1 0 7770 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2565_
timestamp 0
transform 1 0 7990 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2566_
timestamp 0
transform 1 0 7570 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2567_
timestamp 0
transform 1 0 6970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2568_
timestamp 0
transform -1 0 6610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2569_
timestamp 0
transform 1 0 7190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2570_
timestamp 0
transform -1 0 9370 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2571_
timestamp 0
transform -1 0 9270 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2572_
timestamp 0
transform 1 0 9290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2573_
timestamp 0
transform 1 0 9170 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2574_
timestamp 0
transform -1 0 9250 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2575_
timestamp 0
transform -1 0 9070 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2576_
timestamp 0
transform -1 0 8790 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2577_
timestamp 0
transform -1 0 8990 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2578_
timestamp 0
transform 1 0 9550 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2579_
timestamp 0
transform -1 0 9490 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2580_
timestamp 0
transform -1 0 8290 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2581_
timestamp 0
transform 1 0 8250 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2582_
timestamp 0
transform 1 0 8370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2583_
timestamp 0
transform -1 0 9770 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2584_
timestamp 0
transform 1 0 9430 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2585_
timestamp 0
transform -1 0 11170 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2586_
timestamp 0
transform 1 0 8850 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2587_
timestamp 0
transform 1 0 8650 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2588_
timestamp 0
transform -1 0 8470 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2589_
timestamp 0
transform 1 0 8510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2590_
timestamp 0
transform 1 0 8250 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2591_
timestamp 0
transform -1 0 8590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2592_
timestamp 0
transform 1 0 7850 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2593_
timestamp 0
transform -1 0 9090 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2594_
timestamp 0
transform -1 0 8990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2595_
timestamp 0
transform -1 0 9250 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2596_
timestamp 0
transform 1 0 10430 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2597_
timestamp 0
transform 1 0 10610 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2598_
timestamp 0
transform -1 0 10450 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2599_
timestamp 0
transform 1 0 10810 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2600_
timestamp 0
transform -1 0 11410 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2601_
timestamp 0
transform 1 0 8270 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2602_
timestamp 0
transform -1 0 8070 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2603_
timestamp 0
transform 1 0 7070 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2604_
timestamp 0
transform 1 0 8230 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2605_
timestamp 0
transform -1 0 8110 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2606_
timestamp 0
transform -1 0 7710 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2607_
timestamp 0
transform -1 0 6570 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2608_
timestamp 0
transform 1 0 6750 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2609_
timestamp 0
transform 1 0 6950 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2610_
timestamp 0
transform -1 0 7890 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2611_
timestamp 0
transform -1 0 10110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2612_
timestamp 0
transform 1 0 9890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2613_
timestamp 0
transform 1 0 10290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2614_
timestamp 0
transform -1 0 10990 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__2615_
timestamp 0
transform -1 0 7170 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2616_
timestamp 0
transform 1 0 8310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2617_
timestamp 0
transform -1 0 7170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2618_
timestamp 0
transform -1 0 6510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2619_
timestamp 0
transform 1 0 6290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2620_
timestamp 0
transform -1 0 7990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2621_
timestamp 0
transform -1 0 8090 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2622_
timestamp 0
transform 1 0 8350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2623_
timestamp 0
transform -1 0 8950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2624_
timestamp 0
transform 1 0 8090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2625_
timestamp 0
transform 1 0 6850 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2626_
timestamp 0
transform -1 0 8310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2627_
timestamp 0
transform 1 0 9910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2628_
timestamp 0
transform 1 0 11530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2629_
timestamp 0
transform 1 0 11430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2630_
timestamp 0
transform 1 0 11710 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2631_
timestamp 0
transform -1 0 11530 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2632_
timestamp 0
transform 1 0 9430 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2633_
timestamp 0
transform -1 0 8530 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2634_
timestamp 0
transform 1 0 8930 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2635_
timestamp 0
transform -1 0 9170 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2636_
timestamp 0
transform -1 0 9950 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2637_
timestamp 0
transform -1 0 8650 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2638_
timestamp 0
transform 1 0 9730 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2639_
timestamp 0
transform 1 0 9990 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2640_
timestamp 0
transform 1 0 8110 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2641_
timestamp 0
transform 1 0 7910 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2642_
timestamp 0
transform 1 0 9390 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2643_
timestamp 0
transform 1 0 9390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2644_
timestamp 0
transform 1 0 8410 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2645_
timestamp 0
transform 1 0 7630 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2646_
timestamp 0
transform 1 0 7430 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2647_
timestamp 0
transform 1 0 8210 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2648_
timestamp 0
transform -1 0 8050 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2649_
timestamp 0
transform -1 0 9050 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2650_
timestamp 0
transform 1 0 11110 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2651_
timestamp 0
transform -1 0 9250 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2652_
timestamp 0
transform -1 0 8550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2653_
timestamp 0
transform 1 0 8730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2654_
timestamp 0
transform 1 0 5850 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2655_
timestamp 0
transform -1 0 6070 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2656_
timestamp 0
transform -1 0 6250 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2657_
timestamp 0
transform -1 0 7650 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2658_
timestamp 0
transform 1 0 7410 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2659_
timestamp 0
transform -1 0 7170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2660_
timestamp 0
transform -1 0 7350 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2661_
timestamp 0
transform -1 0 10790 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2662_
timestamp 0
transform 1 0 10970 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2663_
timestamp 0
transform 1 0 10030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2664_
timestamp 0
transform 1 0 10210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2665_
timestamp 0
transform -1 0 6630 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2666_
timestamp 0
transform 1 0 7210 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2667_
timestamp 0
transform -1 0 7010 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2668_
timestamp 0
transform -1 0 6830 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2669_
timestamp 0
transform 1 0 6750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2670_
timestamp 0
transform -1 0 10610 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2671_
timestamp 0
transform 1 0 11670 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2672_
timestamp 0
transform 1 0 11710 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2673_
timestamp 0
transform -1 0 11510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2674_
timestamp 0
transform 1 0 11450 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2675_
timestamp 0
transform -1 0 10810 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2676_
timestamp 0
transform 1 0 11430 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2677_
timestamp 0
transform -1 0 11510 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2678_
timestamp 0
transform -1 0 10130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2679_
timestamp 0
transform 1 0 9730 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2680_
timestamp 0
transform 1 0 9650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2681_
timestamp 0
transform 1 0 9330 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2682_
timestamp 0
transform -1 0 9550 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2683_
timestamp 0
transform -1 0 10210 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2684_
timestamp 0
transform -1 0 10510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2685_
timestamp 0
transform -1 0 10790 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__2686_
timestamp 0
transform 1 0 10690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2687_
timestamp 0
transform -1 0 9810 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2688_
timestamp 0
transform 1 0 9210 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2689_
timestamp 0
transform 1 0 10530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2690_
timestamp 0
transform -1 0 10890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2691_
timestamp 0
transform -1 0 11090 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2692_
timestamp 0
transform 1 0 11270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2693_
timestamp 0
transform -1 0 10430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2694_
timestamp 0
transform 1 0 9630 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2695_
timestamp 0
transform -1 0 10550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2696_
timestamp 0
transform 1 0 10310 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2697_
timestamp 0
transform 1 0 9970 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2698_
timestamp 0
transform 1 0 9950 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2699_
timestamp 0
transform 1 0 9070 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2700_
timestamp 0
transform 1 0 8850 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2701_
timestamp 0
transform -1 0 8490 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2702_
timestamp 0
transform 1 0 8850 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2703_
timestamp 0
transform 1 0 10870 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2704_
timestamp 0
transform -1 0 9130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2705_
timestamp 0
transform -1 0 9690 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2706_
timestamp 0
transform -1 0 10090 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2707_
timestamp 0
transform -1 0 9610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2708_
timestamp 0
transform 1 0 8910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2709_
timestamp 0
transform 1 0 9030 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2710_
timestamp 0
transform -1 0 8730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2711_
timestamp 0
transform -1 0 10790 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2712_
timestamp 0
transform -1 0 10770 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2713_
timestamp 0
transform 1 0 10810 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2714_
timestamp 0
transform 1 0 10810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2715_
timestamp 0
transform -1 0 11450 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2716_
timestamp 0
transform 1 0 11610 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2717_
timestamp 0
transform -1 0 10730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2718_
timestamp 0
transform 1 0 11070 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2719_
timestamp 0
transform 1 0 11790 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2720_
timestamp 0
transform -1 0 10990 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2721_
timestamp 0
transform -1 0 10890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2722_
timestamp 0
transform -1 0 10930 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2723_
timestamp 0
transform 1 0 11370 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2724_
timestamp 0
transform 1 0 11350 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2725_
timestamp 0
transform 1 0 10330 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2726_
timestamp 0
transform -1 0 9710 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2727_
timestamp 0
transform 1 0 9910 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2728_
timestamp 0
transform -1 0 9890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2729_
timestamp 0
transform -1 0 9490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2730_
timestamp 0
transform 1 0 11230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2731_
timestamp 0
transform 1 0 9470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2732_
timestamp 0
transform 1 0 6690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2733_
timestamp 0
transform -1 0 9110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2734_
timestamp 0
transform 1 0 9470 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2735_
timestamp 0
transform 1 0 9490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2736_
timestamp 0
transform -1 0 8910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2737_
timestamp 0
transform -1 0 9290 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2738_
timestamp 0
transform -1 0 10370 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2739_
timestamp 0
transform 1 0 10550 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2740_
timestamp 0
transform 1 0 11170 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2741_
timestamp 0
transform 1 0 11570 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2742_
timestamp 0
transform -1 0 10570 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2743_
timestamp 0
transform -1 0 10410 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2744_
timestamp 0
transform 1 0 10490 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2745_
timestamp 0
transform -1 0 11150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2746_
timestamp 0
transform -1 0 10150 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2747_
timestamp 0
transform 1 0 10950 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2748_
timestamp 0
transform 1 0 9810 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2749_
timestamp 0
transform 1 0 10670 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2750_
timestamp 0
transform 1 0 11010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2751_
timestamp 0
transform -1 0 10130 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2752_
timestamp 0
transform 1 0 5750 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2753_
timestamp 0
transform -1 0 5970 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2754_
timestamp 0
transform -1 0 6030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2755_
timestamp 0
transform -1 0 7390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2756_
timestamp 0
transform -1 0 7510 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2757_
timestamp 0
transform 1 0 8110 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2758_
timestamp 0
transform -1 0 7570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2759_
timestamp 0
transform -1 0 9710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2760_
timestamp 0
transform -1 0 6230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2761_
timestamp 0
transform -1 0 8870 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2762_
timestamp 0
transform -1 0 8850 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2763_
timestamp 0
transform -1 0 6310 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2764_
timestamp 0
transform -1 0 6390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2765_
timestamp 0
transform -1 0 9350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2766_
timestamp 0
transform -1 0 6690 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2767_
timestamp 0
transform 1 0 8910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2768_
timestamp 0
transform -1 0 5990 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2769_
timestamp 0
transform -1 0 6930 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2770_
timestamp 0
transform 1 0 7110 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2771_
timestamp 0
transform 1 0 10030 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2772_
timestamp 0
transform -1 0 7390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2773_
timestamp 0
transform -1 0 7590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2774_
timestamp 0
transform -1 0 6030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2775_
timestamp 0
transform -1 0 7330 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2776_
timestamp 0
transform 1 0 6150 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2777_
timestamp 0
transform -1 0 9870 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2778_
timestamp 0
transform 1 0 7690 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2779_
timestamp 0
transform 1 0 7910 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2780_
timestamp 0
transform 1 0 7970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2781_
timestamp 0
transform -1 0 7790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2782_
timestamp 0
transform 1 0 7650 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2783_
timestamp 0
transform -1 0 8450 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2784_
timestamp 0
transform -1 0 10990 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2785_
timestamp 0
transform 1 0 9510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2786_
timestamp 0
transform -1 0 7770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2787_
timestamp 0
transform -1 0 9210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2788_
timestamp 0
transform -1 0 10190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2789_
timestamp 0
transform 1 0 10370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2790_
timestamp 0
transform 1 0 7970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2791_
timestamp 0
transform 1 0 8170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2792_
timestamp 0
transform -1 0 7630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2793_
timestamp 0
transform -1 0 7850 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2794_
timestamp 0
transform -1 0 7850 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2795_
timestamp 0
transform -1 0 7570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2796_
timestamp 0
transform -1 0 6970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2797_
timestamp 0
transform -1 0 8390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2798_
timestamp 0
transform 1 0 11930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2799_
timestamp 0
transform -1 0 7350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2800_
timestamp 0
transform -1 0 7470 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2801_
timestamp 0
transform 1 0 7110 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2802_
timestamp 0
transform 1 0 6770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2803_
timestamp 0
transform -1 0 6990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2804_
timestamp 0
transform -1 0 8490 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2805_
timestamp 0
transform 1 0 6910 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2806_
timestamp 0
transform -1 0 6810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2807_
timestamp 0
transform -1 0 7070 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2808_
timestamp 0
transform 1 0 10150 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2809_
timestamp 0
transform -1 0 10570 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2810_
timestamp 0
transform 1 0 10550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2811_
timestamp 0
transform 1 0 10370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2812_
timestamp 0
transform 1 0 10230 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2813_
timestamp 0
transform -1 0 10070 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2814_
timestamp 0
transform -1 0 10470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2815_
timestamp 0
transform -1 0 10670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2816_
timestamp 0
transform 1 0 10190 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2817_
timestamp 0
transform -1 0 10290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2818_
timestamp 0
transform -1 0 10950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2819_
timestamp 0
transform -1 0 11050 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2820_
timestamp 0
transform -1 0 11250 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2821_
timestamp 0
transform 1 0 11010 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2822_
timestamp 0
transform -1 0 11950 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2823_
timestamp 0
transform 1 0 11130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2824_
timestamp 0
transform 1 0 10630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2825_
timestamp 0
transform 1 0 11150 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2826_
timestamp 0
transform 1 0 11350 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2827_
timestamp 0
transform -1 0 11810 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2828_
timestamp 0
transform -1 0 11930 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2829_
timestamp 0
transform -1 0 11370 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2830_
timestamp 0
transform 1 0 11010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2831_
timestamp 0
transform 1 0 11070 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2832_
timestamp 0
transform -1 0 11310 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2833_
timestamp 0
transform 1 0 11370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2834_
timestamp 0
transform 1 0 11870 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2835_
timestamp 0
transform 1 0 12050 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__2836_
timestamp 0
transform 1 0 11670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2837_
timestamp 0
transform 1 0 11870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2838_
timestamp 0
transform 1 0 11990 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2839_
timestamp 0
transform 1 0 11570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2840_
timestamp 0
transform -1 0 11770 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2841_
timestamp 0
transform -1 0 11630 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2842_
timestamp 0
transform -1 0 9810 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2843_
timestamp 0
transform -1 0 10010 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2844_
timestamp 0
transform -1 0 11790 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2845_
timestamp 0
transform 1 0 11970 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2846_
timestamp 0
transform 1 0 11530 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__2847_
timestamp 0
transform 1 0 11950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2848_
timestamp 0
transform -1 0 11590 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2849_
timestamp 0
transform -1 0 11690 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2850_
timestamp 0
transform 1 0 11870 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2851_
timestamp 0
transform -1 0 9870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2852_
timestamp 0
transform -1 0 11050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2853_
timestamp 0
transform 1 0 11230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2854_
timestamp 0
transform 1 0 11810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2855_
timestamp 0
transform 1 0 11810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2856_
timestamp 0
transform -1 0 9830 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2857_
timestamp 0
transform -1 0 9890 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2858_
timestamp 0
transform -1 0 8050 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2859_
timestamp 0
transform 1 0 9670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2860_
timestamp 0
transform -1 0 9130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2861_
timestamp 0
transform 1 0 9950 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2862_
timestamp 0
transform 1 0 9550 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2863_
timestamp 0
transform 1 0 8770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2864_
timestamp 0
transform -1 0 7770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2865_
timestamp 0
transform -1 0 6430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2866_
timestamp 0
transform -1 0 8850 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2867_
timestamp 0
transform -1 0 9390 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2868_
timestamp 0
transform 1 0 9190 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2869_
timestamp 0
transform -1 0 10550 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2870_
timestamp 0
transform -1 0 9310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2871_
timestamp 0
transform -1 0 8550 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2872_
timestamp 0
transform 1 0 9750 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2873_
timestamp 0
transform 1 0 9790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2874_
timestamp 0
transform 1 0 9590 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2875_
timestamp 0
transform -1 0 11190 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__2876_
timestamp 0
transform 1 0 10190 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2877_
timestamp 0
transform -1 0 10730 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2878_
timestamp 0
transform 1 0 9630 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2879_
timestamp 0
transform -1 0 9850 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2880_
timestamp 0
transform -1 0 10170 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2881_
timestamp 0
transform -1 0 5950 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2882_
timestamp 0
transform -1 0 6130 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2883_
timestamp 0
transform -1 0 5490 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2884_
timestamp 0
transform -1 0 5490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2885_
timestamp 0
transform 1 0 5470 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2886_
timestamp 0
transform -1 0 5290 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__2887_
timestamp 0
transform 1 0 5630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2888_
timestamp 0
transform 1 0 6050 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2889_
timestamp 0
transform -1 0 6290 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2890_
timestamp 0
transform -1 0 6670 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2891_
timestamp 0
transform 1 0 8150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2892_
timestamp 0
transform -1 0 7270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2893_
timestamp 0
transform -1 0 5870 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2894_
timestamp 0
transform 1 0 5370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2895_
timestamp 0
transform -1 0 7470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2896_
timestamp 0
transform -1 0 6590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__2897_
timestamp 0
transform 1 0 7330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2898_
timestamp 0
transform 1 0 11750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2899_
timestamp 0
transform -1 0 6530 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2900_
timestamp 0
transform -1 0 6730 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2901_
timestamp 0
transform -1 0 8170 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2902_
timestamp 0
transform 1 0 9630 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2903_
timestamp 0
transform -1 0 11570 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2904_
timestamp 0
transform 1 0 8350 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2905_
timestamp 0
transform -1 0 6930 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2906_
timestamp 0
transform -1 0 7310 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2907_
timestamp 0
transform -1 0 6330 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2908_
timestamp 0
transform 1 0 8450 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2909_
timestamp 0
transform -1 0 10350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2910_
timestamp 0
transform 1 0 10750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2911_
timestamp 0
transform 1 0 10930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2912_
timestamp 0
transform -1 0 10790 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2913_
timestamp 0
transform -1 0 8670 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2914_
timestamp 0
transform -1 0 8550 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2915_
timestamp 0
transform -1 0 11230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2916_
timestamp 0
transform -1 0 7970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2917_
timestamp 0
transform -1 0 6990 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2918_
timestamp 0
transform 1 0 6770 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2919_
timestamp 0
transform -1 0 7190 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2920_
timestamp 0
transform 1 0 7150 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2921_
timestamp 0
transform 1 0 6950 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2922_
timestamp 0
transform 1 0 6610 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2923_
timestamp 0
transform -1 0 5830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2924_
timestamp 0
transform 1 0 8870 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2925_
timestamp 0
transform 1 0 10230 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2926_
timestamp 0
transform 1 0 11970 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2927_
timestamp 0
transform 1 0 8690 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2928_
timestamp 0
transform 1 0 7490 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2929_
timestamp 0
transform 1 0 8210 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2930_
timestamp 0
transform -1 0 8430 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2931_
timestamp 0
transform -1 0 8070 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2932_
timestamp 0
transform 1 0 7870 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2933_
timestamp 0
transform 1 0 7910 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2934_
timestamp 0
transform -1 0 10210 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2935_
timestamp 0
transform 1 0 11330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__2936_
timestamp 0
transform -1 0 8190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2937_
timestamp 0
transform 1 0 8670 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2938_
timestamp 0
transform -1 0 11790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2939_
timestamp 0
transform -1 0 11230 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2940_
timestamp 0
transform -1 0 6570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2941_
timestamp 0
transform 1 0 8850 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2942_
timestamp 0
transform 1 0 8930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2943_
timestamp 0
transform 1 0 9690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2944_
timestamp 0
transform 1 0 9870 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__2945_
timestamp 0
transform 1 0 9050 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2946_
timestamp 0
transform -1 0 9150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2947_
timestamp 0
transform -1 0 8710 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2948_
timestamp 0
transform -1 0 8650 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2949_
timestamp 0
transform 1 0 10830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2950_
timestamp 0
transform 1 0 11650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2951_
timestamp 0
transform -1 0 6970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2952_
timestamp 0
transform -1 0 6770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2953_
timestamp 0
transform 1 0 11270 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2954_
timestamp 0
transform -1 0 8950 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2955_
timestamp 0
transform -1 0 10090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__2956_
timestamp 0
transform -1 0 11350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2957_
timestamp 0
transform 1 0 9670 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2958_
timestamp 0
transform 1 0 11630 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__2959_
timestamp 0
transform 1 0 5110 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2960_
timestamp 0
transform -1 0 7370 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2961_
timestamp 0
transform -1 0 7970 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2962_
timestamp 0
transform -1 0 7570 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2963_
timestamp 0
transform -1 0 6490 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__2964_
timestamp 0
transform -1 0 7770 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2965_
timestamp 0
transform -1 0 11750 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__2966_
timestamp 0
transform 1 0 8570 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2967_
timestamp 0
transform 1 0 9270 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__2968_
timestamp 0
transform 1 0 10390 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2969_
timestamp 0
transform 1 0 10590 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__2970_
timestamp 0
transform -1 0 11270 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2971_
timestamp 0
transform 1 0 7730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2972_
timestamp 0
transform -1 0 9330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2973_
timestamp 0
transform 1 0 7370 0 1 250
box -6 -8 26 248
use FILL  FILL_2__2974_
timestamp 0
transform -1 0 7310 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2975_
timestamp 0
transform -1 0 9070 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__2976_
timestamp 0
transform 1 0 10050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2977_
timestamp 0
transform 1 0 10450 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2978_
timestamp 0
transform -1 0 11610 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__2979_
timestamp 0
transform -1 0 11850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__2980_
timestamp 0
transform 1 0 7170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2981_
timestamp 0
transform 1 0 6570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__2982_
timestamp 0
transform 1 0 7510 0 1 730
box -6 -8 26 248
use FILL  FILL_2__2983_
timestamp 0
transform 1 0 11890 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__2984_
timestamp 0
transform 1 0 11630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__2985_
timestamp 0
transform -1 0 7130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__2986_
timestamp 0
transform -1 0 7150 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__2987_
timestamp 0
transform 1 0 5810 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__3000_
timestamp 0
transform -1 0 2210 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3001_
timestamp 0
transform 1 0 2350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3002_
timestamp 0
transform 1 0 2150 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__3003_
timestamp 0
transform -1 0 3630 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__3004_
timestamp 0
transform 1 0 3830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__3005_
timestamp 0
transform -1 0 3470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__3006_
timestamp 0
transform -1 0 4350 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__3007_
timestamp 0
transform -1 0 4150 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__3008_
timestamp 0
transform 1 0 3870 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__3009_
timestamp 0
transform 1 0 3970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3010_
timestamp 0
transform -1 0 3990 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__3011_
timestamp 0
transform 1 0 3790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3012_
timestamp 0
transform 1 0 2730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__3013_
timestamp 0
transform -1 0 2430 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3014_
timestamp 0
transform 1 0 2570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__3015_
timestamp 0
transform -1 0 4550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3016_
timestamp 0
transform 1 0 4470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__3017_
timestamp 0
transform 1 0 4170 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3018_
timestamp 0
transform 1 0 4370 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3019_
timestamp 0
transform -1 0 3990 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3020_
timestamp 0
transform 1 0 1810 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3021_
timestamp 0
transform 1 0 1650 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3022_
timestamp 0
transform -1 0 2050 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3023_
timestamp 0
transform -1 0 2890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3024_
timestamp 0
transform 1 0 4710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3025_
timestamp 0
transform 1 0 4330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3026_
timestamp 0
transform 1 0 3590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3027_
timestamp 0
transform 1 0 3290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__3028_
timestamp 0
transform -1 0 2790 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__3029_
timestamp 0
transform 1 0 3430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3030_
timestamp 0
transform 1 0 4870 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__3031_
timestamp 0
transform 1 0 4710 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__3032_
timestamp 0
transform 1 0 5870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3033_
timestamp 0
transform -1 0 4590 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3034_
timestamp 0
transform 1 0 3810 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3035_
timestamp 0
transform -1 0 4570 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__3036_
timestamp 0
transform -1 0 2370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__3037_
timestamp 0
transform -1 0 3310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__3038_
timestamp 0
transform 1 0 2190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__3039_
timestamp 0
transform -1 0 3570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3040_
timestamp 0
transform -1 0 3790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3041_
timestamp 0
transform 1 0 3390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3042_
timestamp 0
transform -1 0 2770 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3043_
timestamp 0
transform -1 0 3810 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__3044_
timestamp 0
transform -1 0 2610 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3045_
timestamp 0
transform -1 0 2910 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__3046_
timestamp 0
transform -1 0 3250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3047_
timestamp 0
transform 1 0 2850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3048_
timestamp 0
transform 1 0 3390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__3049_
timestamp 0
transform -1 0 3690 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__3050_
timestamp 0
transform -1 0 2930 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__3051_
timestamp 0
transform -1 0 2950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__3052_
timestamp 0
transform 1 0 3110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__3053_
timestamp 0
transform -1 0 2990 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3054_
timestamp 0
transform -1 0 2590 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__3055_
timestamp 0
transform -1 0 2410 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__3056_
timestamp 0
transform -1 0 2730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3057_
timestamp 0
transform -1 0 3250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3058_
timestamp 0
transform 1 0 4170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3059_
timestamp 0
transform -1 0 5090 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__3060_
timestamp 0
transform -1 0 5290 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__3061_
timestamp 0
transform -1 0 6050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3062_
timestamp 0
transform -1 0 5110 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__3063_
timestamp 0
transform -1 0 5130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__3064_
timestamp 0
transform -1 0 4970 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3076_
timestamp 0
transform 1 0 1070 0 1 250
box -6 -8 26 248
use FILL  FILL_2__3077_
timestamp 0
transform -1 0 1290 0 1 250
box -6 -8 26 248
use FILL  FILL_2__3078_
timestamp 0
transform 1 0 910 0 1 250
box -6 -8 26 248
use FILL  FILL_2__3079_
timestamp 0
transform 1 0 990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__3080_
timestamp 0
transform -1 0 870 0 1 730
box -6 -8 26 248
use FILL  FILL_2__3081_
timestamp 0
transform 1 0 810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__3082_
timestamp 0
transform 1 0 1390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__3083_
timestamp 0
transform -1 0 1550 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__3084_
timestamp 0
transform 1 0 1470 0 1 250
box -6 -8 26 248
use FILL  FILL_2__3085_
timestamp 0
transform -1 0 1750 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__3086_
timestamp 0
transform -1 0 450 0 1 730
box -6 -8 26 248
use FILL  FILL_2__3087_
timestamp 0
transform -1 0 630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__3088_
timestamp 0
transform 1 0 430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__3089_
timestamp 0
transform -1 0 1410 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__3090_
timestamp 0
transform 1 0 1210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3091_
timestamp 0
transform -1 0 1890 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__3092_
timestamp 0
transform -1 0 670 0 1 730
box -6 -8 26 248
use FILL  FILL_2__3093_
timestamp 0
transform -1 0 70 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__3094_
timestamp 0
transform -1 0 70 0 1 730
box -6 -8 26 248
use FILL  FILL_2__3095_
timestamp 0
transform -1 0 270 0 1 730
box -6 -8 26 248
use FILL  FILL_2__3096_
timestamp 0
transform -1 0 270 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__3097_
timestamp 0
transform 1 0 2030 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__3098_
timestamp 0
transform -1 0 2330 0 1 250
box -6 -8 26 248
use FILL  FILL_2__3099_
timestamp 0
transform 1 0 1890 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__3100_
timestamp 0
transform 1 0 50 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3101_
timestamp 0
transform -1 0 70 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__3102_
timestamp 0
transform -1 0 1250 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__3103_
timestamp 0
transform -1 0 1210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__3104_
timestamp 0
transform -1 0 250 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__3105_
timestamp 0
transform -1 0 1170 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__3106_
timestamp 0
transform -1 0 2330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__3107_
timestamp 0
transform -1 0 1530 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__3108_
timestamp 0
transform -1 0 410 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3109_
timestamp 0
transform -1 0 590 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3110_
timestamp 0
transform 1 0 730 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__3111_
timestamp 0
transform -1 0 930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__3112_
timestamp 0
transform -1 0 70 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__3113_
timestamp 0
transform -1 0 70 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3114_
timestamp 0
transform -1 0 4570 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__3115_
timestamp 0
transform -1 0 4630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3116_
timestamp 0
transform 1 0 4490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__3117_
timestamp 0
transform 1 0 530 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__3118_
timestamp 0
transform -1 0 1690 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__3119_
timestamp 0
transform 1 0 870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3120_
timestamp 0
transform 1 0 1030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3121_
timestamp 0
transform -1 0 2350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3122_
timestamp 0
transform -1 0 450 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__3123_
timestamp 0
transform 1 0 330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__3124_
timestamp 0
transform 1 0 230 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__3125_
timestamp 0
transform 1 0 2050 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__3126_
timestamp 0
transform -1 0 2270 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__3127_
timestamp 0
transform 1 0 1570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3128_
timestamp 0
transform 1 0 1410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3129_
timestamp 0
transform 1 0 4750 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__3130_
timestamp 0
transform 1 0 4930 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__3131_
timestamp 0
transform 1 0 5150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__3132_
timestamp 0
transform 1 0 4810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3133_
timestamp 0
transform -1 0 4710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__3134_
timestamp 0
transform -1 0 4350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__3135_
timestamp 0
transform 1 0 710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__3136_
timestamp 0
transform -1 0 770 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__3137_
timestamp 0
transform 1 0 370 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__3138_
timestamp 0
transform 1 0 710 0 1 250
box -6 -8 26 248
use FILL  FILL_2__3139_
timestamp 0
transform 1 0 230 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__3140_
timestamp 0
transform -1 0 1530 0 1 730
box -6 -8 26 248
use FILL  FILL_2__3141_
timestamp 0
transform 1 0 1710 0 1 730
box -6 -8 26 248
use FILL  FILL_2__3142_
timestamp 0
transform -1 0 1690 0 1 250
box -6 -8 26 248
use FILL  FILL_2__3143_
timestamp 0
transform 1 0 2390 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__3144_
timestamp 0
transform 1 0 2510 0 1 250
box -6 -8 26 248
use FILL  FILL_2__3145_
timestamp 0
transform 1 0 2230 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__3146_
timestamp 0
transform -1 0 1930 0 1 730
box -6 -8 26 248
use FILL  FILL_2__3147_
timestamp 0
transform 1 0 2030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__3148_
timestamp 0
transform 1 0 1070 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__3149_
timestamp 0
transform -1 0 910 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__3150_
timestamp 0
transform -1 0 270 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__3151_
timestamp 0
transform 1 0 50 0 1 250
box -6 -8 26 248
use FILL  FILL_2__3152_
timestamp 0
transform -1 0 2130 0 1 730
box -6 -8 26 248
use FILL  FILL_2__3284_
timestamp 0
transform -1 0 4730 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__3285_
timestamp 0
transform 1 0 4370 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__3286_
timestamp 0
transform -1 0 3410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3287_
timestamp 0
transform 1 0 3270 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3288_
timestamp 0
transform 1 0 2190 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3289_
timestamp 0
transform 1 0 2390 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3290_
timestamp 0
transform -1 0 2070 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3291_
timestamp 0
transform 1 0 3010 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3292_
timestamp 0
transform 1 0 3210 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3293_
timestamp 0
transform 1 0 5830 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3294_
timestamp 0
transform -1 0 5870 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3295_
timestamp 0
transform 1 0 5910 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3296_
timestamp 0
transform 1 0 6390 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3297_
timestamp 0
transform 1 0 6590 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3298_
timestamp 0
transform 1 0 5290 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3299_
timestamp 0
transform 1 0 5490 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3300_
timestamp 0
transform 1 0 4630 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3301_
timestamp 0
transform 1 0 4830 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3302_
timestamp 0
transform -1 0 3390 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3303_
timestamp 0
transform -1 0 3550 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3304_
timestamp 0
transform -1 0 3430 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3305_
timestamp 0
transform -1 0 3610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3306_
timestamp 0
transform 1 0 4350 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3307_
timestamp 0
transform 1 0 4450 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3308_
timestamp 0
transform -1 0 1110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3309_
timestamp 0
transform -1 0 1030 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__3310_
timestamp 0
transform 1 0 2510 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3311_
timestamp 0
transform -1 0 2730 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3312_
timestamp 0
transform 1 0 3450 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3313_
timestamp 0
transform -1 0 2370 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3314_
timestamp 0
transform -1 0 250 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__3315_
timestamp 0
transform -1 0 450 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__3316_
timestamp 0
transform -1 0 7530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__3317_
timestamp 0
transform 1 0 6150 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3318_
timestamp 0
transform 1 0 2630 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3319_
timestamp 0
transform 1 0 6650 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3320_
timestamp 0
transform 1 0 5430 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3321_
timestamp 0
transform -1 0 6450 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__3322_
timestamp 0
transform -1 0 3810 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3323_
timestamp 0
transform -1 0 3650 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3324_
timestamp 0
transform 1 0 5150 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3325_
timestamp 0
transform -1 0 5370 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3326_
timestamp 0
transform -1 0 5230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__3327_
timestamp 0
transform 1 0 4810 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__3328_
timestamp 0
transform -1 0 5270 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3329_
timestamp 0
transform -1 0 5690 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__3330_
timestamp 0
transform 1 0 5550 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3331_
timestamp 0
transform 1 0 4970 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3332_
timestamp 0
transform -1 0 4650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__3333_
timestamp 0
transform -1 0 5950 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3334_
timestamp 0
transform 1 0 5930 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__3335_
timestamp 0
transform -1 0 450 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3336_
timestamp 0
transform -1 0 270 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3337_
timestamp 0
transform -1 0 890 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3338_
timestamp 0
transform -1 0 910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3339_
timestamp 0
transform -1 0 5870 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__3340_
timestamp 0
transform 1 0 6050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__3341_
timestamp 0
transform -1 0 5830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3342_
timestamp 0
transform -1 0 5450 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3343_
timestamp 0
transform -1 0 4370 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3344_
timestamp 0
transform -1 0 5490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__3345_
timestamp 0
transform 1 0 5670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__3346_
timestamp 0
transform 1 0 5270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__3347_
timestamp 0
transform 1 0 5090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__3348_
timestamp 0
transform -1 0 70 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3349_
timestamp 0
transform 1 0 250 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3350_
timestamp 0
transform 1 0 7770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__3351_
timestamp 0
transform -1 0 70 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3352_
timestamp 0
transform 1 0 290 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3353_
timestamp 0
transform -1 0 1810 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3354_
timestamp 0
transform 1 0 1990 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3355_
timestamp 0
transform -1 0 310 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3356_
timestamp 0
transform -1 0 510 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3357_
timestamp 0
transform -1 0 850 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3358_
timestamp 0
transform -1 0 830 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3359_
timestamp 0
transform -1 0 70 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3360_
timestamp 0
transform -1 0 270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__3361_
timestamp 0
transform -1 0 4870 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3362_
timestamp 0
transform -1 0 4990 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3363_
timestamp 0
transform 1 0 5310 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3364_
timestamp 0
transform -1 0 3410 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3365_
timestamp 0
transform 1 0 3330 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3366_
timestamp 0
transform 1 0 2910 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3367_
timestamp 0
transform 1 0 2550 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3368_
timestamp 0
transform 1 0 2350 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3369_
timestamp 0
transform -1 0 4130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3370_
timestamp 0
transform -1 0 5290 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3371_
timestamp 0
transform -1 0 7050 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3372_
timestamp 0
transform 1 0 5090 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3373_
timestamp 0
transform -1 0 7490 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3374_
timestamp 0
transform -1 0 7270 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3375_
timestamp 0
transform -1 0 4670 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3376_
timestamp 0
transform -1 0 4710 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3377_
timestamp 0
transform 1 0 4890 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3378_
timestamp 0
transform -1 0 4310 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3379_
timestamp 0
transform 1 0 5750 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3380_
timestamp 0
transform -1 0 7810 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3381_
timestamp 0
transform 1 0 6650 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3382_
timestamp 0
transform 1 0 6470 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3383_
timestamp 0
transform -1 0 7070 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3384_
timestamp 0
transform -1 0 6870 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3385_
timestamp 0
transform 1 0 7250 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3386_
timestamp 0
transform -1 0 6510 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3387_
timestamp 0
transform 1 0 6290 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3388_
timestamp 0
transform 1 0 6710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3389_
timestamp 0
transform -1 0 7110 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3390_
timestamp 0
transform -1 0 9710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3391_
timestamp 0
transform -1 0 10250 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3392_
timestamp 0
transform -1 0 250 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3393_
timestamp 0
transform 1 0 230 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3394_
timestamp 0
transform -1 0 230 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3395_
timestamp 0
transform -1 0 250 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3396_
timestamp 0
transform -1 0 70 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3397_
timestamp 0
transform -1 0 1230 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3398_
timestamp 0
transform 1 0 1010 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3399_
timestamp 0
transform 1 0 970 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3400_
timestamp 0
transform -1 0 610 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3401_
timestamp 0
transform -1 0 70 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3402_
timestamp 0
transform -1 0 830 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3403_
timestamp 0
transform 1 0 1590 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3404_
timestamp 0
transform -1 0 890 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3405_
timestamp 0
transform 1 0 690 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3406_
timestamp 0
transform -1 0 1870 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3407_
timestamp 0
transform -1 0 470 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__3408_
timestamp 0
transform 1 0 250 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__3409_
timestamp 0
transform -1 0 70 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__3410_
timestamp 0
transform -1 0 890 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3411_
timestamp 0
transform -1 0 430 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3412_
timestamp 0
transform -1 0 250 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3413_
timestamp 0
transform -1 0 70 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3414_
timestamp 0
transform -1 0 230 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3415_
timestamp 0
transform -1 0 70 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3416_
timestamp 0
transform -1 0 70 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3417_
timestamp 0
transform -1 0 410 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3418_
timestamp 0
transform -1 0 6930 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3419_
timestamp 0
transform 1 0 6230 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3420_
timestamp 0
transform 1 0 6030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3421_
timestamp 0
transform 1 0 5270 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3422_
timestamp 0
transform 1 0 5130 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3423_
timestamp 0
transform 1 0 7110 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3424_
timestamp 0
transform -1 0 1370 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3425_
timestamp 0
transform 1 0 610 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3426_
timestamp 0
transform 1 0 410 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3427_
timestamp 0
transform -1 0 430 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3428_
timestamp 0
transform -1 0 270 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3429_
timestamp 0
transform 1 0 590 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3430_
timestamp 0
transform -1 0 70 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3431_
timestamp 0
transform -1 0 250 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3432_
timestamp 0
transform 1 0 870 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3433_
timestamp 0
transform 1 0 1470 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3434_
timestamp 0
transform -1 0 970 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3435_
timestamp 0
transform -1 0 1090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3436_
timestamp 0
transform 1 0 1270 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3437_
timestamp 0
transform -1 0 1310 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__3438_
timestamp 0
transform -1 0 990 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3439_
timestamp 0
transform -1 0 790 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3440_
timestamp 0
transform -1 0 1110 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__3441_
timestamp 0
transform 1 0 710 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3442_
timestamp 0
transform 1 0 810 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3443_
timestamp 0
transform -1 0 790 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3444_
timestamp 0
transform -1 0 610 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3445_
timestamp 0
transform -1 0 730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__3446_
timestamp 0
transform -1 0 1390 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3447_
timestamp 0
transform -1 0 1170 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3448_
timestamp 0
transform -1 0 710 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3449_
timestamp 0
transform 1 0 1330 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3450_
timestamp 0
transform 1 0 1510 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3451_
timestamp 0
transform -1 0 2630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3452_
timestamp 0
transform -1 0 2830 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3453_
timestamp 0
transform -1 0 3050 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3454_
timestamp 0
transform -1 0 1170 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__3455_
timestamp 0
transform -1 0 270 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3456_
timestamp 0
transform -1 0 70 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3457_
timestamp 0
transform -1 0 830 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3458_
timestamp 0
transform 1 0 610 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3459_
timestamp 0
transform -1 0 550 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__3460_
timestamp 0
transform 1 0 450 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3461_
timestamp 0
transform -1 0 1890 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3462_
timestamp 0
transform 1 0 1670 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3463_
timestamp 0
transform -1 0 1930 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__3464_
timestamp 0
transform -1 0 2050 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3465_
timestamp 0
transform -1 0 1630 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3466_
timestamp 0
transform -1 0 2010 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__3467_
timestamp 0
transform -1 0 1870 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3468_
timestamp 0
transform -1 0 2270 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3469_
timestamp 0
transform -1 0 270 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3470_
timestamp 0
transform -1 0 1210 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3471_
timestamp 0
transform -1 0 1190 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3472_
timestamp 0
transform -1 0 1570 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3473_
timestamp 0
transform 1 0 1750 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3474_
timestamp 0
transform -1 0 2050 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3475_
timestamp 0
transform -1 0 1730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3476_
timestamp 0
transform -1 0 1690 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3477_
timestamp 0
transform -1 0 1870 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3478_
timestamp 0
transform 1 0 1950 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3479_
timestamp 0
transform -1 0 1410 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3480_
timestamp 0
transform -1 0 2810 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3481_
timestamp 0
transform -1 0 6050 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3482_
timestamp 0
transform -1 0 5870 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3483_
timestamp 0
transform 1 0 6710 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3484_
timestamp 0
transform -1 0 7470 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__3485_
timestamp 0
transform -1 0 7270 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__3486_
timestamp 0
transform 1 0 5730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__3487_
timestamp 0
transform -1 0 5750 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3488_
timestamp 0
transform 1 0 2970 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3489_
timestamp 0
transform -1 0 6110 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__3490_
timestamp 0
transform 1 0 1530 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3491_
timestamp 0
transform 1 0 1350 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3492_
timestamp 0
transform 1 0 1910 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3493_
timestamp 0
transform -1 0 1750 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3494_
timestamp 0
transform 1 0 7190 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3495_
timestamp 0
transform -1 0 7570 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3496_
timestamp 0
transform -1 0 7770 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3497_
timestamp 0
transform -1 0 8190 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3498_
timestamp 0
transform -1 0 7410 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3499_
timestamp 0
transform 1 0 1150 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__3500_
timestamp 0
transform 1 0 1350 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__3501_
timestamp 0
transform -1 0 3130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3502_
timestamp 0
transform -1 0 3730 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3503_
timestamp 0
transform -1 0 3230 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3504_
timestamp 0
transform 1 0 2930 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__3505_
timestamp 0
transform 1 0 3130 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__3506_
timestamp 0
transform -1 0 750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__3507_
timestamp 0
transform -1 0 950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__3508_
timestamp 0
transform 1 0 6350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__3509_
timestamp 0
transform -1 0 6590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__3510_
timestamp 0
transform 1 0 6810 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__3511_
timestamp 0
transform -1 0 6630 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__3512_
timestamp 0
transform 1 0 6570 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__3513_
timestamp 0
transform 1 0 6750 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__3514_
timestamp 0
transform -1 0 6490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3515_
timestamp 0
transform 1 0 7150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__3516_
timestamp 0
transform -1 0 1210 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3517_
timestamp 0
transform 1 0 990 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3518_
timestamp 0
transform -1 0 7470 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3519_
timestamp 0
transform -1 0 7290 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3520_
timestamp 0
transform 1 0 5310 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3521_
timestamp 0
transform -1 0 5510 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3522_
timestamp 0
transform -1 0 70 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__3523_
timestamp 0
transform 1 0 230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3524_
timestamp 0
transform -1 0 450 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__3525_
timestamp 0
transform 1 0 2030 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__3526_
timestamp 0
transform 1 0 2210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__3527_
timestamp 0
transform 1 0 7010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__3528_
timestamp 0
transform -1 0 6950 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__3529_
timestamp 0
transform -1 0 70 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3530_
timestamp 0
transform 1 0 10090 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3531_
timestamp 0
transform 1 0 6050 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3532_
timestamp 0
transform 1 0 5670 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3533_
timestamp 0
transform 1 0 11830 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3534_
timestamp 0
transform -1 0 9130 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3535_
timestamp 0
transform 1 0 7630 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3536_
timestamp 0
transform 1 0 6030 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__3537_
timestamp 0
transform 1 0 5570 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3538_
timestamp 0
transform 1 0 5550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3539_
timestamp 0
transform 1 0 6150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3540_
timestamp 0
transform 1 0 6350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3541_
timestamp 0
transform -1 0 6230 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3542_
timestamp 0
transform -1 0 6050 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3543_
timestamp 0
transform 1 0 5950 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3544_
timestamp 0
transform 1 0 5830 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3545_
timestamp 0
transform 1 0 5830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3546_
timestamp 0
transform -1 0 6210 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__3547_
timestamp 0
transform 1 0 6370 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3548_
timestamp 0
transform 1 0 6470 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3549_
timestamp 0
transform 1 0 6670 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3550_
timestamp 0
transform 1 0 6530 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3551_
timestamp 0
transform -1 0 6730 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3552_
timestamp 0
transform 1 0 6810 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3553_
timestamp 0
transform -1 0 7250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__3554_
timestamp 0
transform 1 0 11210 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3555_
timestamp 0
transform 1 0 10870 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3556_
timestamp 0
transform 1 0 10130 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3557_
timestamp 0
transform -1 0 9210 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3558_
timestamp 0
transform -1 0 10710 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3559_
timestamp 0
transform 1 0 11550 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3560_
timestamp 0
transform 1 0 10010 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3561_
timestamp 0
transform 1 0 9990 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3562_
timestamp 0
transform 1 0 9790 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3563_
timestamp 0
transform -1 0 9870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3564_
timestamp 0
transform -1 0 11810 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3565_
timestamp 0
transform 1 0 11990 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3566_
timestamp 0
transform 1 0 11410 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3567_
timestamp 0
transform 1 0 11050 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3568_
timestamp 0
transform 1 0 11190 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3569_
timestamp 0
transform 1 0 9730 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3570_
timestamp 0
transform 1 0 10630 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3571_
timestamp 0
transform 1 0 9550 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3572_
timestamp 0
transform -1 0 9390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3573_
timestamp 0
transform 1 0 10990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3574_
timestamp 0
transform -1 0 9330 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3575_
timestamp 0
transform 1 0 8530 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3576_
timestamp 0
transform -1 0 8010 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3577_
timestamp 0
transform -1 0 8990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3578_
timestamp 0
transform -1 0 9070 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3579_
timestamp 0
transform -1 0 8190 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3580_
timestamp 0
transform -1 0 8650 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3581_
timestamp 0
transform 1 0 9590 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3582_
timestamp 0
transform 1 0 9390 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3583_
timestamp 0
transform 1 0 8450 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3584_
timestamp 0
transform -1 0 8390 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3585_
timestamp 0
transform 1 0 9110 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3586_
timestamp 0
transform -1 0 8950 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3587_
timestamp 0
transform -1 0 9190 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3588_
timestamp 0
transform 1 0 8190 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3589_
timestamp 0
transform -1 0 9010 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3590_
timestamp 0
transform -1 0 10590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3591_
timestamp 0
transform -1 0 10750 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3592_
timestamp 0
transform 1 0 8210 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3593_
timestamp 0
transform -1 0 6190 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3594_
timestamp 0
transform -1 0 10350 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3595_
timestamp 0
transform -1 0 10510 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3596_
timestamp 0
transform 1 0 6950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3597_
timestamp 0
transform 1 0 6610 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3598_
timestamp 0
transform 1 0 11830 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3599_
timestamp 0
transform -1 0 8890 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3600_
timestamp 0
transform 1 0 8670 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3601_
timestamp 0
transform 1 0 8810 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3602_
timestamp 0
transform -1 0 9930 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3603_
timestamp 0
transform -1 0 10250 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3604_
timestamp 0
transform -1 0 8410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3605_
timestamp 0
transform -1 0 7850 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3606_
timestamp 0
transform -1 0 7990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3607_
timestamp 0
transform 1 0 7790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3608_
timestamp 0
transform 1 0 11390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3609_
timestamp 0
transform 1 0 11610 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3610_
timestamp 0
transform 1 0 11470 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3611_
timestamp 0
transform 1 0 11270 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3612_
timestamp 0
transform 1 0 11630 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3613_
timestamp 0
transform 1 0 11370 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3614_
timestamp 0
transform 1 0 11570 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3615_
timestamp 0
transform 1 0 11310 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3616_
timestamp 0
transform -1 0 8090 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3617_
timestamp 0
transform 1 0 12010 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3618_
timestamp 0
transform 1 0 11950 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3619_
timestamp 0
transform -1 0 11530 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3620_
timestamp 0
transform 1 0 8770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3621_
timestamp 0
transform 1 0 8150 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3622_
timestamp 0
transform 1 0 8110 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3623_
timestamp 0
transform 1 0 11110 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3624_
timestamp 0
transform -1 0 11090 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3625_
timestamp 0
transform 1 0 10770 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3626_
timestamp 0
transform 1 0 10970 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3627_
timestamp 0
transform 1 0 10910 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3628_
timestamp 0
transform 1 0 7950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3629_
timestamp 0
transform 1 0 7610 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3630_
timestamp 0
transform 1 0 7590 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3631_
timestamp 0
transform -1 0 7450 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3632_
timestamp 0
transform 1 0 7010 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3633_
timestamp 0
transform 1 0 8010 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3634_
timestamp 0
transform 1 0 8690 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3635_
timestamp 0
transform 1 0 8350 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3636_
timestamp 0
transform -1 0 6830 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3637_
timestamp 0
transform 1 0 8710 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3638_
timestamp 0
transform 1 0 10810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3639_
timestamp 0
transform 1 0 8570 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3640_
timestamp 0
transform 1 0 9430 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3641_
timestamp 0
transform 1 0 8930 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3642_
timestamp 0
transform -1 0 7290 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3643_
timestamp 0
transform 1 0 7090 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3644_
timestamp 0
transform -1 0 9310 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3645_
timestamp 0
transform -1 0 10390 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3646_
timestamp 0
transform 1 0 9090 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3647_
timestamp 0
transform 1 0 10530 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3648_
timestamp 0
transform 1 0 10850 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3649_
timestamp 0
transform 1 0 10950 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3650_
timestamp 0
transform -1 0 11370 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3651_
timestamp 0
transform 1 0 6750 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3652_
timestamp 0
transform 1 0 4810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3653_
timestamp 0
transform 1 0 4610 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3654_
timestamp 0
transform 1 0 4410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3655_
timestamp 0
transform 1 0 4210 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3656_
timestamp 0
transform 1 0 5410 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3657_
timestamp 0
transform 1 0 5370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3658_
timestamp 0
transform 1 0 5210 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3659_
timestamp 0
transform 1 0 4630 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3660_
timestamp 0
transform 1 0 4430 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3661_
timestamp 0
transform 1 0 4810 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3662_
timestamp 0
transform 1 0 6550 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3663_
timestamp 0
transform 1 0 6350 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3664_
timestamp 0
transform 1 0 5590 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3665_
timestamp 0
transform 1 0 5190 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3666_
timestamp 0
transform 1 0 5790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3667_
timestamp 0
transform -1 0 3670 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3668_
timestamp 0
transform 1 0 3890 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3669_
timestamp 0
transform -1 0 3390 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3670_
timestamp 0
transform -1 0 3510 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3671_
timestamp 0
transform 1 0 4150 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3672_
timestamp 0
transform 1 0 4210 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3673_
timestamp 0
transform 1 0 5970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3674_
timestamp 0
transform -1 0 10710 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3675_
timestamp 0
transform -1 0 10530 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3676_
timestamp 0
transform 1 0 4130 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3677_
timestamp 0
transform -1 0 4190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3678_
timestamp 0
transform 1 0 4630 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3679_
timestamp 0
transform -1 0 4850 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3680_
timestamp 0
transform -1 0 5050 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3681_
timestamp 0
transform -1 0 4750 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3682_
timestamp 0
transform 1 0 1630 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__3683_
timestamp 0
transform 1 0 6250 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3684_
timestamp 0
transform 1 0 6590 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3685_
timestamp 0
transform 1 0 6870 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3686_
timestamp 0
transform 1 0 6650 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3687_
timestamp 0
transform 1 0 4870 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3688_
timestamp 0
transform -1 0 4890 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3689_
timestamp 0
transform 1 0 5070 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3690_
timestamp 0
transform -1 0 4730 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3691_
timestamp 0
transform -1 0 4670 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3692_
timestamp 0
transform 1 0 4470 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3693_
timestamp 0
transform 1 0 4850 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3694_
timestamp 0
transform -1 0 6050 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3695_
timestamp 0
transform 1 0 1690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3696_
timestamp 0
transform 1 0 7570 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3697_
timestamp 0
transform 1 0 7770 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3698_
timestamp 0
transform 1 0 6670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3699_
timestamp 0
transform 1 0 6870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3700_
timestamp 0
transform -1 0 7070 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3701_
timestamp 0
transform 1 0 4630 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__3702_
timestamp 0
transform 1 0 4330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3703_
timestamp 0
transform 1 0 4390 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3704_
timestamp 0
transform 1 0 4810 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3705_
timestamp 0
transform -1 0 4890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3706_
timestamp 0
transform -1 0 4670 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__3707_
timestamp 0
transform -1 0 5010 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3708_
timestamp 0
transform 1 0 4590 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3709_
timestamp 0
transform 1 0 2450 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3710_
timestamp 0
transform 1 0 9770 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3711_
timestamp 0
transform 1 0 9650 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3712_
timestamp 0
transform 1 0 9630 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3713_
timestamp 0
transform 1 0 10010 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3714_
timestamp 0
transform 1 0 8710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3715_
timestamp 0
transform -1 0 8910 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3716_
timestamp 0
transform -1 0 9510 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3717_
timestamp 0
transform -1 0 10410 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3718_
timestamp 0
transform 1 0 10570 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3719_
timestamp 0
transform -1 0 9110 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3720_
timestamp 0
transform 1 0 9290 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3721_
timestamp 0
transform -1 0 10630 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3722_
timestamp 0
transform -1 0 10450 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3723_
timestamp 0
transform 1 0 10770 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3724_
timestamp 0
transform 1 0 9450 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3725_
timestamp 0
transform 1 0 8310 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3726_
timestamp 0
transform -1 0 8190 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3727_
timestamp 0
transform 1 0 9630 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3728_
timestamp 0
transform -1 0 10190 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3729_
timestamp 0
transform 1 0 10030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3730_
timestamp 0
transform 1 0 9990 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3731_
timestamp 0
transform 1 0 8430 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3732_
timestamp 0
transform 1 0 8810 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3733_
timestamp 0
transform -1 0 3870 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3734_
timestamp 0
transform -1 0 4050 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3735_
timestamp 0
transform 1 0 7630 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3736_
timestamp 0
transform -1 0 7230 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3737_
timestamp 0
transform -1 0 5790 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3738_
timestamp 0
transform 1 0 9570 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3739_
timestamp 0
transform 1 0 9370 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3740_
timestamp 0
transform 1 0 9250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3741_
timestamp 0
transform -1 0 10750 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3742_
timestamp 0
transform 1 0 11250 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3743_
timestamp 0
transform 1 0 11430 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3744_
timestamp 0
transform 1 0 11170 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3745_
timestamp 0
transform -1 0 10590 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3746_
timestamp 0
transform -1 0 10250 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3747_
timestamp 0
transform -1 0 10190 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3748_
timestamp 0
transform -1 0 10930 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3749_
timestamp 0
transform -1 0 11250 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3750_
timestamp 0
transform 1 0 11050 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3751_
timestamp 0
transform -1 0 8050 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3752_
timestamp 0
transform -1 0 6850 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3753_
timestamp 0
transform -1 0 6750 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3754_
timestamp 0
transform 1 0 4390 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3755_
timestamp 0
transform 1 0 3030 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3756_
timestamp 0
transform 1 0 4070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3757_
timestamp 0
transform 1 0 4550 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3758_
timestamp 0
transform -1 0 5070 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__3759_
timestamp 0
transform -1 0 4850 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__3760_
timestamp 0
transform -1 0 4290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3761_
timestamp 0
transform -1 0 4310 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__3762_
timestamp 0
transform -1 0 4410 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__3763_
timestamp 0
transform -1 0 4150 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3764_
timestamp 0
transform -1 0 3430 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3765_
timestamp 0
transform -1 0 4610 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__3766_
timestamp 0
transform 1 0 2230 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3767_
timestamp 0
transform -1 0 2450 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3768_
timestamp 0
transform -1 0 2610 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3769_
timestamp 0
transform -1 0 2810 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3770_
timestamp 0
transform -1 0 3810 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3771_
timestamp 0
transform 1 0 3390 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3772_
timestamp 0
transform -1 0 1030 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3773_
timestamp 0
transform 1 0 5810 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__3774_
timestamp 0
transform 1 0 5030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__3775_
timestamp 0
transform -1 0 4990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3776_
timestamp 0
transform -1 0 4830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3777_
timestamp 0
transform 1 0 4890 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3778_
timestamp 0
transform 1 0 4730 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3779_
timestamp 0
transform 1 0 4530 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3780_
timestamp 0
transform 1 0 5210 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3781_
timestamp 0
transform -1 0 5390 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3782_
timestamp 0
transform -1 0 4370 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3783_
timestamp 0
transform 1 0 3810 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3784_
timestamp 0
transform -1 0 5250 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3785_
timestamp 0
transform 1 0 7530 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__3786_
timestamp 0
transform 1 0 7390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__3787_
timestamp 0
transform -1 0 7370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3788_
timestamp 0
transform -1 0 7210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3789_
timestamp 0
transform -1 0 7230 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3790_
timestamp 0
transform -1 0 6210 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3791_
timestamp 0
transform -1 0 6590 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3792_
timestamp 0
transform 1 0 7010 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3793_
timestamp 0
transform -1 0 6810 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3794_
timestamp 0
transform 1 0 7970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__3795_
timestamp 0
transform -1 0 9590 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3796_
timestamp 0
transform 1 0 8290 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3797_
timestamp 0
transform 1 0 7670 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3798_
timestamp 0
transform 1 0 6950 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3799_
timestamp 0
transform -1 0 7130 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3800_
timestamp 0
transform -1 0 7310 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3801_
timestamp 0
transform 1 0 5650 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3802_
timestamp 0
transform -1 0 5910 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3803_
timestamp 0
transform 1 0 5690 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3804_
timestamp 0
transform 1 0 5310 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3805_
timestamp 0
transform 1 0 5350 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3806_
timestamp 0
transform 1 0 5030 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3807_
timestamp 0
transform -1 0 5510 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3808_
timestamp 0
transform -1 0 7890 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3809_
timestamp 0
transform -1 0 8010 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3810_
timestamp 0
transform 1 0 7810 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3811_
timestamp 0
transform -1 0 7490 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3812_
timestamp 0
transform 1 0 10430 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3813_
timestamp 0
transform -1 0 9850 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3814_
timestamp 0
transform 1 0 9830 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3815_
timestamp 0
transform -1 0 9830 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3816_
timestamp 0
transform -1 0 9670 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3817_
timestamp 0
transform 1 0 9130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3818_
timestamp 0
transform -1 0 8950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3819_
timestamp 0
transform 1 0 10130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3820_
timestamp 0
transform 1 0 10210 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3821_
timestamp 0
transform 1 0 6530 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3822_
timestamp 0
transform -1 0 3330 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3823_
timestamp 0
transform -1 0 8250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3824_
timestamp 0
transform 1 0 7270 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3825_
timestamp 0
transform -1 0 9970 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3826_
timestamp 0
transform 1 0 9450 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3827_
timestamp 0
transform -1 0 9290 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3828_
timestamp 0
transform 1 0 9090 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3829_
timestamp 0
transform 1 0 8890 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3830_
timestamp 0
transform 1 0 7390 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3831_
timestamp 0
transform 1 0 7670 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3832_
timestamp 0
transform 1 0 8530 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3833_
timestamp 0
transform 1 0 8710 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3834_
timestamp 0
transform -1 0 8690 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3835_
timestamp 0
transform 1 0 8890 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3836_
timestamp 0
transform 1 0 9190 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3837_
timestamp 0
transform -1 0 8450 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3838_
timestamp 0
transform 1 0 8630 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3839_
timestamp 0
transform 1 0 8870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3840_
timestamp 0
transform -1 0 8510 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3841_
timestamp 0
transform -1 0 8310 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3842_
timestamp 0
transform 1 0 9070 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3843_
timestamp 0
transform -1 0 8330 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3844_
timestamp 0
transform 1 0 7630 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3845_
timestamp 0
transform 1 0 9290 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__3846_
timestamp 0
transform 1 0 8850 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3847_
timestamp 0
transform 1 0 8130 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3848_
timestamp 0
transform -1 0 7990 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__3849_
timestamp 0
transform 1 0 7770 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__3850_
timestamp 0
transform 1 0 7950 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3851_
timestamp 0
transform 1 0 7610 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3852_
timestamp 0
transform -1 0 7810 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3853_
timestamp 0
transform -1 0 7570 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3854_
timestamp 0
transform -1 0 7430 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3855_
timestamp 0
transform 1 0 7810 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__3856_
timestamp 0
transform -1 0 7210 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3857_
timestamp 0
transform -1 0 8310 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3858_
timestamp 0
transform 1 0 8650 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3859_
timestamp 0
transform 1 0 7830 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3860_
timestamp 0
transform 1 0 4770 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3861_
timestamp 0
transform 1 0 8510 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3862_
timestamp 0
transform -1 0 8750 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3863_
timestamp 0
transform -1 0 10210 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3864_
timestamp 0
transform 1 0 9450 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3865_
timestamp 0
transform 1 0 8030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3866_
timestamp 0
transform 1 0 5630 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3867_
timestamp 0
transform -1 0 7470 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3868_
timestamp 0
transform -1 0 8530 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3869_
timestamp 0
transform 1 0 7950 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3870_
timestamp 0
transform -1 0 7830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3871_
timestamp 0
transform 1 0 6370 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3872_
timestamp 0
transform 1 0 5670 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3873_
timestamp 0
transform -1 0 9510 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3874_
timestamp 0
transform 1 0 9850 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__3875_
timestamp 0
transform 1 0 6890 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3876_
timestamp 0
transform 1 0 4990 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3877_
timestamp 0
transform -1 0 4630 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3878_
timestamp 0
transform 1 0 4790 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3879_
timestamp 0
transform 1 0 4550 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3880_
timestamp 0
transform 1 0 5110 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3881_
timestamp 0
transform -1 0 5330 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3882_
timestamp 0
transform -1 0 4350 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3883_
timestamp 0
transform -1 0 4970 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3884_
timestamp 0
transform -1 0 4790 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3885_
timestamp 0
transform 1 0 5150 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3886_
timestamp 0
transform 1 0 9650 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__3887_
timestamp 0
transform 1 0 10370 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__3888_
timestamp 0
transform 1 0 10330 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__3889_
timestamp 0
transform -1 0 10830 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__3890_
timestamp 0
transform -1 0 10750 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3891_
timestamp 0
transform 1 0 10910 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3892_
timestamp 0
transform -1 0 8770 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__3893_
timestamp 0
transform -1 0 8570 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__3894_
timestamp 0
transform -1 0 11270 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3895_
timestamp 0
transform 1 0 11050 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3896_
timestamp 0
transform 1 0 11810 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3897_
timestamp 0
transform 1 0 11070 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__3898_
timestamp 0
transform 1 0 8250 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3899_
timestamp 0
transform -1 0 5610 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3900_
timestamp 0
transform 1 0 4070 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3901_
timestamp 0
transform -1 0 5030 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__3902_
timestamp 0
transform 1 0 4950 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3903_
timestamp 0
transform 1 0 7430 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3904_
timestamp 0
transform -1 0 7010 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3905_
timestamp 0
transform -1 0 6450 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3906_
timestamp 0
transform 1 0 5030 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3907_
timestamp 0
transform -1 0 8190 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__3908_
timestamp 0
transform -1 0 6790 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3909_
timestamp 0
transform -1 0 5970 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__3910_
timestamp 0
transform 1 0 5850 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__3911_
timestamp 0
transform -1 0 4530 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3912_
timestamp 0
transform 1 0 4330 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__3913_
timestamp 0
transform -1 0 4550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3914_
timestamp 0
transform 1 0 4210 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__3915_
timestamp 0
transform 1 0 4750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3916_
timestamp 0
transform 1 0 4950 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3917_
timestamp 0
transform 1 0 5330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3918_
timestamp 0
transform -1 0 4650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3919_
timestamp 0
transform 1 0 4750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__3920_
timestamp 0
transform 1 0 4470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3921_
timestamp 0
transform 1 0 790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3922_
timestamp 0
transform 1 0 890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3923_
timestamp 0
transform 1 0 410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3924_
timestamp 0
transform 1 0 770 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__3925_
timestamp 0
transform 1 0 5070 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3926_
timestamp 0
transform 1 0 5270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3927_
timestamp 0
transform -1 0 4690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3928_
timestamp 0
transform 1 0 5450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3929_
timestamp 0
transform -1 0 4570 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__3930_
timestamp 0
transform 1 0 3410 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__3931_
timestamp 0
transform 1 0 3450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__3932_
timestamp 0
transform 1 0 2310 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__3933_
timestamp 0
transform 1 0 3210 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__3934_
timestamp 0
transform -1 0 4450 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__3935_
timestamp 0
transform 1 0 3810 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3936_
timestamp 0
transform 1 0 3610 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__3937_
timestamp 0
transform 1 0 4190 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__3938_
timestamp 0
transform -1 0 3470 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__3939_
timestamp 0
transform 1 0 3570 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__3940_
timestamp 0
transform -1 0 4710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__3941_
timestamp 0
transform 1 0 6910 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3942_
timestamp 0
transform -1 0 9990 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3943_
timestamp 0
transform -1 0 9970 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__3944_
timestamp 0
transform -1 0 9670 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__3945_
timestamp 0
transform -1 0 10190 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3946_
timestamp 0
transform 1 0 9770 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__3947_
timestamp 0
transform 1 0 10370 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3948_
timestamp 0
transform 1 0 10550 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3949_
timestamp 0
transform 1 0 7670 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__3950_
timestamp 0
transform -1 0 6950 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3951_
timestamp 0
transform 1 0 6550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3952_
timestamp 0
transform -1 0 5770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__3953_
timestamp 0
transform 1 0 5430 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3954_
timestamp 0
transform -1 0 5830 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3955_
timestamp 0
transform 1 0 5890 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3956_
timestamp 0
transform -1 0 6110 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3957_
timestamp 0
transform 1 0 6130 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3958_
timestamp 0
transform 1 0 6330 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3959_
timestamp 0
transform 1 0 6450 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3960_
timestamp 0
transform 1 0 2370 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3961_
timestamp 0
transform -1 0 2770 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3962_
timestamp 0
transform 1 0 2910 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3963_
timestamp 0
transform 1 0 3510 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3964_
timestamp 0
transform -1 0 4090 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3965_
timestamp 0
transform -1 0 3330 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3966_
timestamp 0
transform -1 0 4290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3967_
timestamp 0
transform -1 0 5090 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3968_
timestamp 0
transform -1 0 5290 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3969_
timestamp 0
transform -1 0 4290 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3970_
timestamp 0
transform 1 0 3910 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3971_
timestamp 0
transform 1 0 5610 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__3972_
timestamp 0
transform 1 0 5430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__3973_
timestamp 0
transform 1 0 5430 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3974_
timestamp 0
transform -1 0 5650 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3975_
timestamp 0
transform -1 0 5650 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3976_
timestamp 0
transform -1 0 5650 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3977_
timestamp 0
transform 1 0 5530 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__3978_
timestamp 0
transform 1 0 6350 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3979_
timestamp 0
transform -1 0 2710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3980_
timestamp 0
transform 1 0 2010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__3981_
timestamp 0
transform 1 0 1850 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__3982_
timestamp 0
transform 1 0 1790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__3983_
timestamp 0
transform -1 0 1930 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__3984_
timestamp 0
transform 1 0 8250 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__3985_
timestamp 0
transform 1 0 6830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3986_
timestamp 0
transform -1 0 7330 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__3987_
timestamp 0
transform 1 0 7610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3988_
timestamp 0
transform 1 0 7530 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3989_
timestamp 0
transform 1 0 7330 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3990_
timestamp 0
transform 1 0 7130 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3991_
timestamp 0
transform -1 0 7290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__3992_
timestamp 0
transform -1 0 7950 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3993_
timestamp 0
transform 1 0 7710 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3994_
timestamp 0
transform -1 0 7050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__3995_
timestamp 0
transform -1 0 9410 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3996_
timestamp 0
transform -1 0 6010 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__3997_
timestamp 0
transform 1 0 5970 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__3998_
timestamp 0
transform -1 0 6050 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__3999_
timestamp 0
transform 1 0 5830 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4000_
timestamp 0
transform -1 0 5250 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4001_
timestamp 0
transform -1 0 5090 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4002_
timestamp 0
transform -1 0 6950 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4003_
timestamp 0
transform -1 0 6590 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4004_
timestamp 0
transform 1 0 2630 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4005_
timestamp 0
transform 1 0 2830 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4006_
timestamp 0
transform -1 0 2650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4007_
timestamp 0
transform 1 0 2430 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4008_
timestamp 0
transform -1 0 7110 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4009_
timestamp 0
transform 1 0 6890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4010_
timestamp 0
transform -1 0 6750 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4011_
timestamp 0
transform 1 0 8630 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4012_
timestamp 0
transform 1 0 6730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4013_
timestamp 0
transform 1 0 6610 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4014_
timestamp 0
transform 1 0 6150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4015_
timestamp 0
transform 1 0 6510 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4016_
timestamp 0
transform 1 0 9330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4017_
timestamp 0
transform -1 0 9650 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4018_
timestamp 0
transform -1 0 9830 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4019_
timestamp 0
transform 1 0 9990 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4020_
timestamp 0
transform -1 0 7470 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4021_
timestamp 0
transform -1 0 10030 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4022_
timestamp 0
transform -1 0 6810 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4023_
timestamp 0
transform -1 0 7150 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4024_
timestamp 0
transform 1 0 8950 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4025_
timestamp 0
transform -1 0 7670 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4026_
timestamp 0
transform -1 0 7830 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4027_
timestamp 0
transform 1 0 8370 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4028_
timestamp 0
transform 1 0 7910 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4029_
timestamp 0
transform 1 0 11010 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4030_
timestamp 0
transform 1 0 10830 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4031_
timestamp 0
transform 1 0 9210 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4032_
timestamp 0
transform 1 0 8650 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4033_
timestamp 0
transform -1 0 9310 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4034_
timestamp 0
transform 1 0 3970 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4035_
timestamp 0
transform 1 0 9770 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4036_
timestamp 0
transform -1 0 9630 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4037_
timestamp 0
transform -1 0 9150 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4038_
timestamp 0
transform -1 0 8110 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4039_
timestamp 0
transform -1 0 7050 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4040_
timestamp 0
transform 1 0 11990 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4041_
timestamp 0
transform 1 0 9270 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4042_
timestamp 0
transform -1 0 5990 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__4043_
timestamp 0
transform 1 0 5310 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4044_
timestamp 0
transform -1 0 5390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4045_
timestamp 0
transform -1 0 5450 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4046_
timestamp 0
transform -1 0 5810 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4047_
timestamp 0
transform -1 0 5990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4048_
timestamp 0
transform -1 0 5990 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4049_
timestamp 0
transform 1 0 5470 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4050_
timestamp 0
transform -1 0 5250 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4051_
timestamp 0
transform 1 0 5590 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4052_
timestamp 0
transform -1 0 6210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4053_
timestamp 0
transform -1 0 8190 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4054_
timestamp 0
transform 1 0 3710 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4055_
timestamp 0
transform -1 0 3550 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4056_
timestamp 0
transform 1 0 2710 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4057_
timestamp 0
transform 1 0 3330 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4058_
timestamp 0
transform -1 0 7470 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4059_
timestamp 0
transform 1 0 7330 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4060_
timestamp 0
transform -1 0 8010 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4061_
timestamp 0
transform -1 0 8950 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4062_
timestamp 0
transform -1 0 3130 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4063_
timestamp 0
transform 1 0 5050 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4064_
timestamp 0
transform -1 0 5030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4065_
timestamp 0
transform 1 0 5250 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4066_
timestamp 0
transform 1 0 4450 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4067_
timestamp 0
transform -1 0 7090 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4068_
timestamp 0
transform 1 0 3110 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4069_
timestamp 0
transform -1 0 650 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__4070_
timestamp 0
transform 1 0 1130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__4071_
timestamp 0
transform 1 0 530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__4072_
timestamp 0
transform -1 0 850 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__4073_
timestamp 0
transform 1 0 4070 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4074_
timestamp 0
transform 1 0 4270 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4075_
timestamp 0
transform 1 0 4190 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4076_
timestamp 0
transform -1 0 5450 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4077_
timestamp 0
transform 1 0 5470 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4078_
timestamp 0
transform -1 0 5490 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4079_
timestamp 0
transform 1 0 3750 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4080_
timestamp 0
transform 1 0 5850 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4081_
timestamp 0
transform 1 0 890 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4082_
timestamp 0
transform 1 0 4130 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4083_
timestamp 0
transform -1 0 3930 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4084_
timestamp 0
transform 1 0 1630 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4085_
timestamp 0
transform 1 0 1450 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4086_
timestamp 0
transform 1 0 1590 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4087_
timestamp 0
transform 1 0 1550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4088_
timestamp 0
transform -1 0 4490 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4089_
timestamp 0
transform -1 0 4450 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4090_
timestamp 0
transform -1 0 3950 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4091_
timestamp 0
transform -1 0 3390 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4092_
timestamp 0
transform -1 0 5670 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4093_
timestamp 0
transform 1 0 4610 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4094_
timestamp 0
transform 1 0 4190 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4095_
timestamp 0
transform 1 0 1930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4096_
timestamp 0
transform 1 0 1750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4097_
timestamp 0
transform 1 0 1630 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4098_
timestamp 0
transform 1 0 1550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4099_
timestamp 0
transform 1 0 7130 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4100_
timestamp 0
transform 1 0 8010 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4101_
timestamp 0
transform 1 0 8170 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4102_
timestamp 0
transform -1 0 8370 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4103_
timestamp 0
transform 1 0 7990 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4104_
timestamp 0
transform -1 0 8210 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4105_
timestamp 0
transform 1 0 8650 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4106_
timestamp 0
transform 1 0 6690 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4107_
timestamp 0
transform -1 0 1090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2__4108_
timestamp 0
transform -1 0 490 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__4109_
timestamp 0
transform -1 0 1830 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4110_
timestamp 0
transform -1 0 7770 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4111_
timestamp 0
transform -1 0 9510 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4112_
timestamp 0
transform 1 0 2890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__4113_
timestamp 0
transform 1 0 3090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__4114_
timestamp 0
transform 1 0 3590 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4115_
timestamp 0
transform 1 0 4470 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4116_
timestamp 0
transform -1 0 5350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4117_
timestamp 0
transform 1 0 4890 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4118_
timestamp 0
transform 1 0 4810 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4119_
timestamp 0
transform 1 0 3970 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4120_
timestamp 0
transform -1 0 3710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4121_
timestamp 0
transform -1 0 4550 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4122_
timestamp 0
transform 1 0 4690 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4123_
timestamp 0
transform 1 0 8050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4124_
timestamp 0
transform 1 0 8570 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4125_
timestamp 0
transform -1 0 4290 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4126_
timestamp 0
transform 1 0 4250 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4127_
timestamp 0
transform 1 0 4070 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4128_
timestamp 0
transform 1 0 4490 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4129_
timestamp 0
transform -1 0 4910 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4130_
timestamp 0
transform 1 0 6030 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4131_
timestamp 0
transform 1 0 4310 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4132_
timestamp 0
transform -1 0 4530 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4133_
timestamp 0
transform -1 0 2010 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4134_
timestamp 0
transform 1 0 1790 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4135_
timestamp 0
transform -1 0 2150 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4136_
timestamp 0
transform -1 0 2150 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4137_
timestamp 0
transform -1 0 1990 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4138_
timestamp 0
transform -1 0 2230 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4139_
timestamp 0
transform 1 0 2010 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4140_
timestamp 0
transform -1 0 3030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4141_
timestamp 0
transform 1 0 1810 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4142_
timestamp 0
transform 1 0 1610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4143_
timestamp 0
transform -1 0 1450 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4144_
timestamp 0
transform 1 0 1590 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4145_
timestamp 0
transform -1 0 1070 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4146_
timestamp 0
transform 1 0 3090 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4147_
timestamp 0
transform -1 0 2030 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4148_
timestamp 0
transform -1 0 3210 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4149_
timestamp 0
transform 1 0 3190 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4150_
timestamp 0
transform 1 0 3190 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4151_
timestamp 0
transform 1 0 3730 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4152_
timestamp 0
transform -1 0 3670 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4153_
timestamp 0
transform -1 0 2050 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4154_
timestamp 0
transform -1 0 2250 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4155_
timestamp 0
transform 1 0 630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4156_
timestamp 0
transform 1 0 990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4157_
timestamp 0
transform -1 0 5930 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4158_
timestamp 0
transform 1 0 6090 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4159_
timestamp 0
transform 1 0 6290 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4160_
timestamp 0
transform 1 0 5370 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4161_
timestamp 0
transform -1 0 5590 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4162_
timestamp 0
transform 1 0 5170 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4163_
timestamp 0
transform -1 0 5190 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4164_
timestamp 0
transform 1 0 5730 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4165_
timestamp 0
transform -1 0 5730 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4166_
timestamp 0
transform 1 0 5750 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4167_
timestamp 0
transform 1 0 6450 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4168_
timestamp 0
transform -1 0 5890 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4169_
timestamp 0
transform 1 0 5690 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4170_
timestamp 0
transform 1 0 6090 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4171_
timestamp 0
transform 1 0 5510 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4172_
timestamp 0
transform 1 0 5130 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4173_
timestamp 0
transform 1 0 3810 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4174_
timestamp 0
transform 1 0 5530 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4175_
timestamp 0
transform 1 0 5150 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4176_
timestamp 0
transform -1 0 3330 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4177_
timestamp 0
transform 1 0 3010 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4178_
timestamp 0
transform -1 0 2230 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4179_
timestamp 0
transform -1 0 2350 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4180_
timestamp 0
transform 1 0 2810 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4181_
timestamp 0
transform -1 0 2430 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4182_
timestamp 0
transform 1 0 2270 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4183_
timestamp 0
transform -1 0 3250 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4184_
timestamp 0
transform 1 0 3410 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4185_
timestamp 0
transform 1 0 2830 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4186_
timestamp 0
transform -1 0 2450 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4187_
timestamp 0
transform 1 0 4070 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4188_
timestamp 0
transform 1 0 4270 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4189_
timestamp 0
transform -1 0 4090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4190_
timestamp 0
transform -1 0 3910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4191_
timestamp 0
transform -1 0 3730 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4192_
timestamp 0
transform -1 0 5190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4193_
timestamp 0
transform -1 0 5050 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4194_
timestamp 0
transform -1 0 3910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4195_
timestamp 0
transform 1 0 3450 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4196_
timestamp 0
transform 1 0 3750 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4197_
timestamp 0
transform 1 0 1610 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4198_
timestamp 0
transform -1 0 1730 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4199_
timestamp 0
transform -1 0 1930 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4200_
timestamp 0
transform -1 0 2330 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4201_
timestamp 0
transform -1 0 1550 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4202_
timestamp 0
transform -1 0 1430 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__4203_
timestamp 0
transform -1 0 1810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__4204_
timestamp 0
transform -1 0 2610 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4205_
timestamp 0
transform 1 0 2610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4206_
timestamp 0
transform -1 0 8590 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4207_
timestamp 0
transform -1 0 7930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4208_
timestamp 0
transform -1 0 6270 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4209_
timestamp 0
transform -1 0 270 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4210_
timestamp 0
transform 1 0 50 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4211_
timestamp 0
transform -1 0 70 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4212_
timestamp 0
transform -1 0 450 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4213_
timestamp 0
transform 1 0 910 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4214_
timestamp 0
transform -1 0 1430 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4215_
timestamp 0
transform 1 0 1410 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4216_
timestamp 0
transform -1 0 2010 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4217_
timestamp 0
transform -1 0 2990 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4218_
timestamp 0
transform -1 0 2210 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4219_
timestamp 0
transform 1 0 2290 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4220_
timestamp 0
transform 1 0 2490 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4221_
timestamp 0
transform -1 0 270 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4222_
timestamp 0
transform -1 0 70 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4223_
timestamp 0
transform -1 0 450 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4224_
timestamp 0
transform -1 0 450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4225_
timestamp 0
transform -1 0 430 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4226_
timestamp 0
transform 1 0 50 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4227_
timestamp 0
transform -1 0 270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4228_
timestamp 0
transform -1 0 2410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4229_
timestamp 0
transform 1 0 2610 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4230_
timestamp 0
transform -1 0 2830 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4231_
timestamp 0
transform 1 0 3170 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4232_
timestamp 0
transform -1 0 3630 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4233_
timestamp 0
transform -1 0 2210 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4234_
timestamp 0
transform -1 0 3070 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4235_
timestamp 0
transform -1 0 3830 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4236_
timestamp 0
transform 1 0 3910 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4237_
timestamp 0
transform -1 0 4130 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4238_
timestamp 0
transform 1 0 3450 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4239_
timestamp 0
transform 1 0 2610 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4240_
timestamp 0
transform 1 0 2250 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4241_
timestamp 0
transform -1 0 2110 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4242_
timestamp 0
transform 1 0 2290 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4243_
timestamp 0
transform -1 0 4470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4244_
timestamp 0
transform -1 0 5470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4245_
timestamp 0
transform -1 0 6050 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4246_
timestamp 0
transform -1 0 4170 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4247_
timestamp 0
transform 1 0 2570 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4248_
timestamp 0
transform -1 0 5650 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4249_
timestamp 0
transform -1 0 2350 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4250_
timestamp 0
transform -1 0 4270 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4251_
timestamp 0
transform 1 0 5650 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4252_
timestamp 0
transform -1 0 5850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4253_
timestamp 0
transform -1 0 3750 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4254_
timestamp 0
transform -1 0 2170 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4255_
timestamp 0
transform 1 0 2510 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4256_
timestamp 0
transform -1 0 3870 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4257_
timestamp 0
transform 1 0 4050 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4258_
timestamp 0
transform 1 0 4250 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4259_
timestamp 0
transform 1 0 4010 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4260_
timestamp 0
transform -1 0 2970 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4261_
timestamp 0
transform -1 0 4030 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4262_
timestamp 0
transform 1 0 1550 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4263_
timestamp 0
transform -1 0 7970 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4264_
timestamp 0
transform 1 0 7590 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4265_
timestamp 0
transform 1 0 7410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4266_
timestamp 0
transform 1 0 7090 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4267_
timestamp 0
transform 1 0 7530 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4268_
timestamp 0
transform -1 0 6770 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4269_
timestamp 0
transform -1 0 9450 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4270_
timestamp 0
transform -1 0 11150 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4271_
timestamp 0
transform 1 0 11130 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4272_
timestamp 0
transform 1 0 9230 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4273_
timestamp 0
transform 1 0 9030 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4274_
timestamp 0
transform -1 0 8950 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4275_
timestamp 0
transform 1 0 8770 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4276_
timestamp 0
transform 1 0 8850 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4277_
timestamp 0
transform 1 0 8870 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4278_
timestamp 0
transform 1 0 7750 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4279_
timestamp 0
transform 1 0 10530 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4280_
timestamp 0
transform 1 0 10730 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4281_
timestamp 0
transform -1 0 10690 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4282_
timestamp 0
transform -1 0 1230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4283_
timestamp 0
transform -1 0 7070 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4284_
timestamp 0
transform 1 0 7650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4285_
timestamp 0
transform 1 0 7390 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4286_
timestamp 0
transform -1 0 1070 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4287_
timestamp 0
transform -1 0 1270 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4288_
timestamp 0
transform -1 0 1670 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4289_
timestamp 0
transform -1 0 4370 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4290_
timestamp 0
transform 1 0 6850 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4291_
timestamp 0
transform 1 0 6870 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4292_
timestamp 0
transform -1 0 2530 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4293_
timestamp 0
transform -1 0 1810 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4294_
timestamp 0
transform -1 0 7290 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4295_
timestamp 0
transform 1 0 1490 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4296_
timestamp 0
transform -1 0 70 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4297_
timestamp 0
transform 1 0 1150 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4298_
timestamp 0
transform -1 0 3270 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4299_
timestamp 0
transform 1 0 3350 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4300_
timestamp 0
transform -1 0 3830 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4301_
timestamp 0
transform -1 0 3550 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4302_
timestamp 0
transform -1 0 3670 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4303_
timestamp 0
transform -1 0 1590 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4304_
timestamp 0
transform 1 0 1170 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4305_
timestamp 0
transform -1 0 2290 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4306_
timestamp 0
transform -1 0 2850 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4307_
timestamp 0
transform 1 0 6210 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4308_
timestamp 0
transform -1 0 6290 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4309_
timestamp 0
transform 1 0 2850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4310_
timestamp 0
transform -1 0 2430 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4311_
timestamp 0
transform 1 0 2330 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4312_
timestamp 0
transform 1 0 910 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4313_
timestamp 0
transform 1 0 1490 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4314_
timestamp 0
transform 1 0 1670 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4315_
timestamp 0
transform -1 0 2710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4316_
timestamp 0
transform -1 0 2770 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4317_
timestamp 0
transform 1 0 4410 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4318_
timestamp 0
transform 1 0 4090 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4319_
timestamp 0
transform 1 0 3590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4320_
timestamp 0
transform -1 0 3030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4321_
timestamp 0
transform 1 0 2810 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4322_
timestamp 0
transform 1 0 1550 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4323_
timestamp 0
transform -1 0 2670 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4324_
timestamp 0
transform -1 0 1810 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4325_
timestamp 0
transform -1 0 4070 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4326_
timestamp 0
transform 1 0 3970 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4327_
timestamp 0
transform 1 0 4110 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4328_
timestamp 0
transform -1 0 8550 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4329_
timestamp 0
transform 1 0 1710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4330_
timestamp 0
transform 1 0 2110 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4331_
timestamp 0
transform -1 0 1430 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4332_
timestamp 0
transform -1 0 1970 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4333_
timestamp 0
transform -1 0 2890 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4334_
timestamp 0
transform -1 0 3090 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4335_
timestamp 0
transform -1 0 3670 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4336_
timestamp 0
transform 1 0 2830 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4337_
timestamp 0
transform 1 0 2630 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4338_
timestamp 0
transform 1 0 2670 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4339_
timestamp 0
transform -1 0 3290 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4340_
timestamp 0
transform -1 0 3470 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4341_
timestamp 0
transform 1 0 3410 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4342_
timestamp 0
transform -1 0 3230 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4343_
timestamp 0
transform 1 0 3470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4344_
timestamp 0
transform 1 0 1770 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4345_
timestamp 0
transform -1 0 2410 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4346_
timestamp 0
transform 1 0 6890 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4347_
timestamp 0
transform -1 0 6710 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4348_
timestamp 0
transform -1 0 610 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4349_
timestamp 0
transform -1 0 1030 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4350_
timestamp 0
transform 1 0 2150 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4351_
timestamp 0
transform -1 0 2770 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4352_
timestamp 0
transform 1 0 3750 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4353_
timestamp 0
transform -1 0 6150 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4354_
timestamp 0
transform -1 0 3430 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4355_
timestamp 0
transform -1 0 850 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4356_
timestamp 0
transform -1 0 490 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4357_
timestamp 0
transform 1 0 2350 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4358_
timestamp 0
transform -1 0 5210 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4359_
timestamp 0
transform 1 0 5130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4360_
timestamp 0
transform -1 0 5090 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4361_
timestamp 0
transform 1 0 3030 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4362_
timestamp 0
transform 1 0 4870 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4363_
timestamp 0
transform -1 0 4710 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4364_
timestamp 0
transform 1 0 3670 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4365_
timestamp 0
transform -1 0 5650 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4366_
timestamp 0
transform -1 0 5850 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4367_
timestamp 0
transform -1 0 2890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4368_
timestamp 0
transform 1 0 7530 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4369_
timestamp 0
transform -1 0 7370 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4370_
timestamp 0
transform 1 0 650 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4371_
timestamp 0
transform -1 0 1790 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4372_
timestamp 0
transform 1 0 1910 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4373_
timestamp 0
transform 1 0 2110 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4374_
timestamp 0
transform 1 0 2470 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4375_
timestamp 0
transform -1 0 3790 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4376_
timestamp 0
transform 1 0 7470 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4377_
timestamp 0
transform 1 0 11530 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4378_
timestamp 0
transform -1 0 1250 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4379_
timestamp 0
transform -1 0 5210 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4380_
timestamp 0
transform 1 0 4790 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4381_
timestamp 0
transform 1 0 5890 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4382_
timestamp 0
transform 1 0 230 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4383_
timestamp 0
transform 1 0 50 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4384_
timestamp 0
transform 1 0 6230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4385_
timestamp 0
transform 1 0 6430 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4386_
timestamp 0
transform 1 0 6830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4387_
timestamp 0
transform 1 0 6630 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4388_
timestamp 0
transform -1 0 5430 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4389_
timestamp 0
transform -1 0 6530 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4390_
timestamp 0
transform 1 0 7030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4391_
timestamp 0
transform 1 0 4990 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4392_
timestamp 0
transform -1 0 6330 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4393_
timestamp 0
transform 1 0 6490 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4394_
timestamp 0
transform 1 0 6670 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4395_
timestamp 0
transform 1 0 6790 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4396_
timestamp 0
transform -1 0 6270 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4397_
timestamp 0
transform 1 0 4030 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4398_
timestamp 0
transform 1 0 3010 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4399_
timestamp 0
transform 1 0 2130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4400_
timestamp 0
transform -1 0 6310 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4401_
timestamp 0
transform 1 0 6230 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4402_
timestamp 0
transform -1 0 6070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4403_
timestamp 0
transform -1 0 5610 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4404_
timestamp 0
transform 1 0 1390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4405_
timestamp 0
transform -1 0 1830 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4406_
timestamp 0
transform -1 0 2530 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4407_
timestamp 0
transform -1 0 2330 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4408_
timestamp 0
transform 1 0 1550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4409_
timestamp 0
transform -1 0 1770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4410_
timestamp 0
transform 1 0 3570 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4411_
timestamp 0
transform 1 0 3890 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4412_
timestamp 0
transform 1 0 1730 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4413_
timestamp 0
transform -1 0 250 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4414_
timestamp 0
transform 1 0 250 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4415_
timestamp 0
transform 1 0 430 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4416_
timestamp 0
transform 1 0 1510 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__4417_
timestamp 0
transform -1 0 1730 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__4418_
timestamp 0
transform -1 0 2550 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__4419_
timestamp 0
transform 1 0 2110 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__4420_
timestamp 0
transform 1 0 2230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4421_
timestamp 0
transform 1 0 2430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4422_
timestamp 0
transform -1 0 1970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4423_
timestamp 0
transform -1 0 610 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4424_
timestamp 0
transform 1 0 2030 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4425_
timestamp 0
transform 1 0 1070 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4426_
timestamp 0
transform 1 0 1270 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4427_
timestamp 0
transform 1 0 3530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4428_
timestamp 0
transform -1 0 3370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4429_
timestamp 0
transform 1 0 1250 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4430_
timestamp 0
transform 1 0 1450 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4431_
timestamp 0
transform -1 0 730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4432_
timestamp 0
transform -1 0 610 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4433_
timestamp 0
transform -1 0 850 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4434_
timestamp 0
transform -1 0 1310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__4435_
timestamp 0
transform 1 0 1490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__4436_
timestamp 0
transform 1 0 3090 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__4437_
timestamp 0
transform -1 0 3310 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__4438_
timestamp 0
transform -1 0 6550 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4439_
timestamp 0
transform 1 0 5950 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4440_
timestamp 0
transform -1 0 4730 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4441_
timestamp 0
transform 1 0 4130 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4442_
timestamp 0
transform 1 0 3910 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4443_
timestamp 0
transform 1 0 3790 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4444_
timestamp 0
transform 1 0 3610 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4445_
timestamp 0
transform 1 0 3950 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4446_
timestamp 0
transform 1 0 4370 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4447_
timestamp 0
transform 1 0 4550 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4448_
timestamp 0
transform 1 0 2470 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4449_
timestamp 0
transform 1 0 1030 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4450_
timestamp 0
transform -1 0 1790 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4451_
timestamp 0
transform 1 0 1390 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4452_
timestamp 0
transform -1 0 2190 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4453_
timestamp 0
transform 1 0 7210 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4454_
timestamp 0
transform -1 0 1030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4455_
timestamp 0
transform 1 0 6750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4456_
timestamp 0
transform 1 0 6970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4457_
timestamp 0
transform 1 0 7170 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4458_
timestamp 0
transform -1 0 7370 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4459_
timestamp 0
transform -1 0 6990 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4460_
timestamp 0
transform -1 0 8310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4461_
timestamp 0
transform 1 0 7590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4462_
timestamp 0
transform -1 0 6690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4463_
timestamp 0
transform 1 0 1210 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4464_
timestamp 0
transform -1 0 2510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4465_
timestamp 0
transform -1 0 5850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4466_
timestamp 0
transform 1 0 5990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4467_
timestamp 0
transform 1 0 6410 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4468_
timestamp 0
transform 1 0 6650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4469_
timestamp 0
transform 1 0 6850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4470_
timestamp 0
transform -1 0 6610 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4471_
timestamp 0
transform 1 0 7210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4472_
timestamp 0
transform -1 0 6410 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4473_
timestamp 0
transform 1 0 8130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4474_
timestamp 0
transform -1 0 6230 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4475_
timestamp 0
transform 1 0 2690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4476_
timestamp 0
transform -1 0 1190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4477_
timestamp 0
transform -1 0 2590 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4478_
timestamp 0
transform 1 0 2570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4479_
timestamp 0
transform 1 0 5290 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4480_
timestamp 0
transform 1 0 1370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4481_
timestamp 0
transform 1 0 210 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4482_
timestamp 0
transform 1 0 410 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4483_
timestamp 0
transform 1 0 3170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4484_
timestamp 0
transform -1 0 4930 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4485_
timestamp 0
transform 1 0 5310 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4486_
timestamp 0
transform -1 0 5130 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4487_
timestamp 0
transform -1 0 5510 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4488_
timestamp 0
transform 1 0 5670 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4489_
timestamp 0
transform -1 0 5790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4490_
timestamp 0
transform -1 0 5750 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4491_
timestamp 0
transform -1 0 5830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4492_
timestamp 0
transform 1 0 50 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4493_
timestamp 0
transform -1 0 5670 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4494_
timestamp 0
transform 1 0 5470 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4495_
timestamp 0
transform 1 0 4330 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4496_
timestamp 0
transform 1 0 3790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4497_
timestamp 0
transform -1 0 3570 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4498_
timestamp 0
transform -1 0 4610 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4499_
timestamp 0
transform 1 0 1230 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4500_
timestamp 0
transform 1 0 6330 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4501_
timestamp 0
transform 1 0 6050 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4502_
timestamp 0
transform -1 0 4490 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4503_
timestamp 0
transform 1 0 6450 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4504_
timestamp 0
transform -1 0 1690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__4505_
timestamp 0
transform -1 0 4810 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__4506_
timestamp 0
transform -1 0 5250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4507_
timestamp 0
transform 1 0 5630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__4508_
timestamp 0
transform 1 0 5510 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4509_
timestamp 0
transform -1 0 5730 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4510_
timestamp 0
transform -1 0 5910 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4511_
timestamp 0
transform 1 0 6070 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4512_
timestamp 0
transform 1 0 6170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4513_
timestamp 0
transform 1 0 6190 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4514_
timestamp 0
transform -1 0 1690 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__4515_
timestamp 0
transform -1 0 2530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__4516_
timestamp 0
transform -1 0 4650 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__4517_
timestamp 0
transform -1 0 5130 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4518_
timestamp 0
transform 1 0 5090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4519_
timestamp 0
transform 1 0 5450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4520_
timestamp 0
transform -1 0 5650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4521_
timestamp 0
transform 1 0 6490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4522_
timestamp 0
transform -1 0 8910 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4523_
timestamp 0
transform 1 0 5290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4524_
timestamp 0
transform 1 0 5990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4525_
timestamp 0
transform 1 0 5850 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4526_
timestamp 0
transform -1 0 6430 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4527_
timestamp 0
transform -1 0 4930 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4528_
timestamp 0
transform 1 0 6330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4529_
timestamp 0
transform 1 0 6030 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4530_
timestamp 0
transform 1 0 6010 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4531_
timestamp 0
transform -1 0 2250 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__4532_
timestamp 0
transform -1 0 6270 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4533_
timestamp 0
transform -1 0 6210 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4534_
timestamp 0
transform 1 0 4250 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4535_
timestamp 0
transform 1 0 3650 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4536_
timestamp 0
transform -1 0 1070 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4537_
timestamp 0
transform 1 0 4430 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4538_
timestamp 0
transform -1 0 7670 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4539_
timestamp 0
transform -1 0 3050 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4540_
timestamp 0
transform 1 0 7630 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4541_
timestamp 0
transform 1 0 6490 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4542_
timestamp 0
transform 1 0 3030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4543_
timestamp 0
transform -1 0 2870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4544_
timestamp 0
transform -1 0 890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4545_
timestamp 0
transform 1 0 2110 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4546_
timestamp 0
transform 1 0 2890 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4547_
timestamp 0
transform -1 0 2350 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4548_
timestamp 0
transform -1 0 1730 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4549_
timestamp 0
transform 1 0 2590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4550_
timestamp 0
transform 1 0 2790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4551_
timestamp 0
transform -1 0 2990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4552_
timestamp 0
transform -1 0 2970 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4553_
timestamp 0
transform -1 0 6530 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4554_
timestamp 0
transform 1 0 970 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4555_
timestamp 0
transform -1 0 730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__4556_
timestamp 0
transform 1 0 4330 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4557_
timestamp 0
transform 1 0 4150 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4558_
timestamp 0
transform -1 0 3990 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4559_
timestamp 0
transform 1 0 5010 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4560_
timestamp 0
transform -1 0 8470 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4561_
timestamp 0
transform -1 0 8870 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4562_
timestamp 0
transform 1 0 8390 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4563_
timestamp 0
transform -1 0 6370 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4564_
timestamp 0
transform -1 0 1870 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4565_
timestamp 0
transform 1 0 2690 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4566_
timestamp 0
transform 1 0 3070 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4567_
timestamp 0
transform -1 0 6770 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4568_
timestamp 0
transform 1 0 6690 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4569_
timestamp 0
transform 1 0 1910 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4570_
timestamp 0
transform -1 0 6570 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4571_
timestamp 0
transform 1 0 6270 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4572_
timestamp 0
transform -1 0 9510 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4573_
timestamp 0
transform -1 0 10370 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4574_
timestamp 0
transform -1 0 9550 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4575_
timestamp 0
transform -1 0 6970 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4576_
timestamp 0
transform -1 0 8490 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4577_
timestamp 0
transform -1 0 3010 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4578_
timestamp 0
transform -1 0 5970 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4579_
timestamp 0
transform 1 0 7990 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4580_
timestamp 0
transform 1 0 10170 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4581_
timestamp 0
transform -1 0 7510 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4582_
timestamp 0
transform 1 0 1270 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4583_
timestamp 0
transform -1 0 2350 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4584_
timestamp 0
transform -1 0 2190 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4585_
timestamp 0
transform -1 0 2090 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4586_
timestamp 0
transform -1 0 1910 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4587_
timestamp 0
transform -1 0 1570 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4588_
timestamp 0
transform 1 0 3290 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4589_
timestamp 0
transform 1 0 3830 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4590_
timestamp 0
transform 1 0 1210 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4591_
timestamp 0
transform -1 0 1630 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4592_
timestamp 0
transform 1 0 1430 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4593_
timestamp 0
transform -1 0 3990 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4594_
timestamp 0
transform -1 0 3150 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__4595_
timestamp 0
transform -1 0 2710 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4596_
timestamp 0
transform -1 0 2910 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4597_
timestamp 0
transform 1 0 2770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__4598_
timestamp 0
transform -1 0 2690 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4599_
timestamp 0
transform -1 0 2870 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4600_
timestamp 0
transform -1 0 4030 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4601_
timestamp 0
transform -1 0 3990 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4602_
timestamp 0
transform -1 0 1410 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4603_
timestamp 0
transform -1 0 1350 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4604_
timestamp 0
transform -1 0 2950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__4605_
timestamp 0
transform 1 0 1770 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4606_
timestamp 0
transform -1 0 670 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4607_
timestamp 0
transform -1 0 490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4608_
timestamp 0
transform -1 0 3230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4609_
timestamp 0
transform 1 0 1610 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__4610_
timestamp 0
transform 1 0 2490 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4611_
timestamp 0
transform -1 0 2330 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4612_
timestamp 0
transform -1 0 1990 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4613_
timestamp 0
transform 1 0 1970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__4614_
timestamp 0
transform -1 0 630 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4615_
timestamp 0
transform -1 0 450 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4616_
timestamp 0
transform -1 0 1810 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__4617_
timestamp 0
transform -1 0 1610 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__4618_
timestamp 0
transform -1 0 2510 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4619_
timestamp 0
transform -1 0 1850 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4620_
timestamp 0
transform -1 0 1450 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4621_
timestamp 0
transform 1 0 2110 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4622_
timestamp 0
transform 1 0 2530 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4623_
timestamp 0
transform 1 0 2030 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4624_
timestamp 0
transform 1 0 1230 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4625_
timestamp 0
transform 1 0 850 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4626_
timestamp 0
transform -1 0 690 0 1 11290
box -6 -8 26 248
use FILL  FILL_2__4627_
timestamp 0
transform -1 0 2190 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__4628_
timestamp 0
transform -1 0 1250 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__4629_
timestamp 0
transform 1 0 1030 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2__4630_
timestamp 0
transform 1 0 990 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4631_
timestamp 0
transform 1 0 1570 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4632_
timestamp 0
transform -1 0 730 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4633_
timestamp 0
transform -1 0 550 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4634_
timestamp 0
transform -1 0 7570 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4635_
timestamp 0
transform -1 0 1510 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4636_
timestamp 0
transform 1 0 1310 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4637_
timestamp 0
transform -1 0 1710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4638_
timestamp 0
transform -1 0 870 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2__4639_
timestamp 0
transform 1 0 1070 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4640_
timestamp 0
transform 1 0 930 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4641_
timestamp 0
transform -1 0 1090 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4642_
timestamp 0
transform -1 0 2910 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__4643_
timestamp 0
transform 1 0 3050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2__4644_
timestamp 0
transform -1 0 3490 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__4645_
timestamp 0
transform -1 0 850 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4646_
timestamp 0
transform 1 0 630 0 1 10810
box -6 -8 26 248
use FILL  FILL_2__4647_
timestamp 0
transform -1 0 1250 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4648_
timestamp 0
transform -1 0 1190 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4649_
timestamp 0
transform -1 0 550 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4650_
timestamp 0
transform -1 0 790 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2__4651_
timestamp 0
transform 1 0 4090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__4652_
timestamp 0
transform 1 0 3810 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__4653_
timestamp 0
transform -1 0 4310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__4654_
timestamp 0
transform -1 0 6870 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4655_
timestamp 0
transform 1 0 2530 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4656_
timestamp 0
transform -1 0 2350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4657_
timestamp 0
transform -1 0 2270 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4658_
timestamp 0
transform 1 0 3710 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4659_
timestamp 0
transform -1 0 3930 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4660_
timestamp 0
transform -1 0 4310 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4661_
timestamp 0
transform 1 0 4490 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4662_
timestamp 0
transform 1 0 3950 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4663_
timestamp 0
transform 1 0 3390 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4664_
timestamp 0
transform 1 0 2530 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4665_
timestamp 0
transform -1 0 7810 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4666_
timestamp 0
transform 1 0 7710 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__4667_
timestamp 0
transform 1 0 6230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__4668_
timestamp 0
transform -1 0 6450 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2__4669_
timestamp 0
transform 1 0 430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4670_
timestamp 0
transform 1 0 4010 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4671_
timestamp 0
transform 1 0 3830 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4672_
timestamp 0
transform 1 0 2770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4673_
timestamp 0
transform -1 0 2970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4674_
timestamp 0
transform -1 0 3130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4675_
timestamp 0
transform -1 0 3010 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4676_
timestamp 0
transform -1 0 3610 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4677_
timestamp 0
transform -1 0 3550 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4678_
timestamp 0
transform 1 0 3370 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4679_
timestamp 0
transform -1 0 3210 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4680_
timestamp 0
transform -1 0 2210 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__4681_
timestamp 0
transform 1 0 1990 0 1 2650
box -6 -8 26 248
use FILL  FILL_2__4682_
timestamp 0
transform -1 0 7050 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4683_
timestamp 0
transform -1 0 1850 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4684_
timestamp 0
transform 1 0 3750 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4685_
timestamp 0
transform 1 0 3570 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4686_
timestamp 0
transform 1 0 11110 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4687_
timestamp 0
transform 1 0 11290 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4688_
timestamp 0
transform 1 0 11470 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4689_
timestamp 0
transform 1 0 11650 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4690_
timestamp 0
transform 1 0 10490 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4691_
timestamp 0
transform 1 0 10130 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4692_
timestamp 0
transform 1 0 10210 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4693_
timestamp 0
transform -1 0 9730 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4694_
timestamp 0
transform -1 0 9750 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4695_
timestamp 0
transform 1 0 10590 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4696_
timestamp 0
transform 1 0 10910 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4697_
timestamp 0
transform 1 0 11390 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4698_
timestamp 0
transform 1 0 11230 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4699_
timestamp 0
transform 1 0 11230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4700_
timestamp 0
transform 1 0 11070 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4701_
timestamp 0
transform -1 0 11450 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4702_
timestamp 0
transform 1 0 11430 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4703_
timestamp 0
transform 1 0 11710 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4704_
timestamp 0
transform -1 0 11610 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4705_
timestamp 0
transform -1 0 11810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4706_
timestamp 0
transform -1 0 11750 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4707_
timestamp 0
transform 1 0 10690 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4708_
timestamp 0
transform 1 0 10890 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4709_
timestamp 0
transform -1 0 10890 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4710_
timestamp 0
transform -1 0 10690 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4711_
timestamp 0
transform 1 0 10150 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4712_
timestamp 0
transform -1 0 9930 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4713_
timestamp 0
transform 1 0 9730 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4714_
timestamp 0
transform 1 0 9530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4715_
timestamp 0
transform -1 0 9850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4716_
timestamp 0
transform 1 0 9270 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4717_
timestamp 0
transform 1 0 9610 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4718_
timestamp 0
transform -1 0 8750 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4719_
timestamp 0
transform 1 0 11290 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4720_
timestamp 0
transform 1 0 10030 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4721_
timestamp 0
transform 1 0 9850 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4722_
timestamp 0
transform -1 0 9930 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4723_
timestamp 0
transform -1 0 9930 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4724_
timestamp 0
transform 1 0 4230 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4725_
timestamp 0
transform -1 0 10130 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4726_
timestamp 0
transform -1 0 10330 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4727_
timestamp 0
transform -1 0 11090 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4728_
timestamp 0
transform 1 0 10170 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4729_
timestamp 0
transform -1 0 10110 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4730_
timestamp 0
transform -1 0 9990 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4731_
timestamp 0
transform -1 0 11670 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4732_
timestamp 0
transform -1 0 9830 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4733_
timestamp 0
transform 1 0 9810 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4734_
timestamp 0
transform -1 0 7790 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4735_
timestamp 0
transform 1 0 9330 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4736_
timestamp 0
transform -1 0 10030 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4737_
timestamp 0
transform 1 0 9530 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4738_
timestamp 0
transform -1 0 9730 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4739_
timestamp 0
transform -1 0 9910 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4740_
timestamp 0
transform -1 0 10290 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4741_
timestamp 0
transform -1 0 10110 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4742_
timestamp 0
transform 1 0 10330 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4743_
timestamp 0
transform 1 0 10090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4744_
timestamp 0
transform 1 0 10590 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4745_
timestamp 0
transform 1 0 10910 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4746_
timestamp 0
transform 1 0 10390 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4747_
timestamp 0
transform 1 0 8330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4748_
timestamp 0
transform 1 0 8530 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4749_
timestamp 0
transform -1 0 8770 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4750_
timestamp 0
transform 1 0 8530 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4751_
timestamp 0
transform 1 0 3730 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4752_
timestamp 0
transform -1 0 9130 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4753_
timestamp 0
transform -1 0 8010 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4754_
timestamp 0
transform 1 0 8130 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4755_
timestamp 0
transform 1 0 7250 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4756_
timestamp 0
transform 1 0 6910 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4757_
timestamp 0
transform 1 0 8350 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4758_
timestamp 0
transform -1 0 10410 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4759_
timestamp 0
transform 1 0 10770 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4760_
timestamp 0
transform -1 0 11050 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4761_
timestamp 0
transform 1 0 11330 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4762_
timestamp 0
transform -1 0 10490 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4763_
timestamp 0
transform 1 0 11830 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4764_
timestamp 0
transform 1 0 10870 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4765_
timestamp 0
transform -1 0 11130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4766_
timestamp 0
transform -1 0 10490 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4767_
timestamp 0
transform -1 0 10510 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4768_
timestamp 0
transform 1 0 10290 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4769_
timestamp 0
transform 1 0 10670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4770_
timestamp 0
transform 1 0 11150 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4771_
timestamp 0
transform 1 0 12010 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4772_
timestamp 0
transform 1 0 9350 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4773_
timestamp 0
transform -1 0 8810 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4774_
timestamp 0
transform 1 0 2550 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4775_
timestamp 0
transform 1 0 2710 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4776_
timestamp 0
transform 1 0 2870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4777_
timestamp 0
transform -1 0 3090 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4778_
timestamp 0
transform -1 0 3690 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4779_
timestamp 0
transform 1 0 3870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4780_
timestamp 0
transform -1 0 8750 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4781_
timestamp 0
transform 1 0 3590 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4782_
timestamp 0
transform 1 0 3270 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4783_
timestamp 0
transform 1 0 9090 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4784_
timestamp 0
transform 1 0 7730 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4785_
timestamp 0
transform 1 0 2090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4786_
timestamp 0
transform -1 0 3970 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__4787_
timestamp 0
transform -1 0 3650 0 1 3130
box -6 -8 26 248
use FILL  FILL_2__4788_
timestamp 0
transform -1 0 4170 0 1 3610
box -6 -8 26 248
use FILL  FILL_2__4789_
timestamp 0
transform 1 0 7210 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4790_
timestamp 0
transform 1 0 7270 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4791_
timestamp 0
transform -1 0 7810 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4792_
timestamp 0
transform -1 0 7870 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4793_
timestamp 0
transform -1 0 7810 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4794_
timestamp 0
transform -1 0 7450 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4795_
timestamp 0
transform -1 0 7510 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4796_
timestamp 0
transform 1 0 11810 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4797_
timestamp 0
transform 1 0 8550 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4798_
timestamp 0
transform 1 0 10010 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4799_
timestamp 0
transform -1 0 9850 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4800_
timestamp 0
transform 1 0 8490 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4801_
timestamp 0
transform 1 0 10950 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4802_
timestamp 0
transform -1 0 10490 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4803_
timestamp 0
transform -1 0 7390 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4804_
timestamp 0
transform -1 0 7070 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4805_
timestamp 0
transform -1 0 6950 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4806_
timestamp 0
transform -1 0 9310 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4807_
timestamp 0
transform -1 0 9090 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4808_
timestamp 0
transform -1 0 8710 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4809_
timestamp 0
transform -1 0 8710 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4810_
timestamp 0
transform -1 0 8950 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4811_
timestamp 0
transform 1 0 11930 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4812_
timestamp 0
transform 1 0 12010 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4813_
timestamp 0
transform 1 0 11470 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4814_
timestamp 0
transform 1 0 11350 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4815_
timestamp 0
transform -1 0 9050 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4816_
timestamp 0
transform -1 0 9490 0 1 7450
box -6 -8 26 248
use FILL  FILL_2__4817_
timestamp 0
transform -1 0 11550 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4818_
timestamp 0
transform -1 0 11490 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4819_
timestamp 0
transform -1 0 6430 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4820_
timestamp 0
transform 1 0 7990 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4821_
timestamp 0
transform 1 0 11630 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4822_
timestamp 0
transform 1 0 11830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4823_
timestamp 0
transform 1 0 11610 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4824_
timestamp 0
transform -1 0 11470 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4825_
timestamp 0
transform 1 0 11170 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4826_
timestamp 0
transform -1 0 11010 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4827_
timestamp 0
transform -1 0 11710 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4828_
timestamp 0
transform -1 0 11790 0 1 10330
box -6 -8 26 248
use FILL  FILL_2__4829_
timestamp 0
transform 1 0 11630 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4830_
timestamp 0
transform 1 0 8990 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4831_
timestamp 0
transform -1 0 9350 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4832_
timestamp 0
transform 1 0 11890 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4833_
timestamp 0
transform 1 0 8370 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4834_
timestamp 0
transform 1 0 8170 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4835_
timestamp 0
transform -1 0 8370 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4836_
timestamp 0
transform 1 0 9650 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4837_
timestamp 0
transform -1 0 10790 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4838_
timestamp 0
transform 1 0 11810 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4839_
timestamp 0
transform 1 0 12070 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4840_
timestamp 0
transform 1 0 9250 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4841_
timestamp 0
transform 1 0 10290 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4842_
timestamp 0
transform 1 0 11990 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4843_
timestamp 0
transform 1 0 11150 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4844_
timestamp 0
transform -1 0 11130 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4845_
timestamp 0
transform -1 0 11910 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4846_
timestamp 0
transform 1 0 11890 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4847_
timestamp 0
transform -1 0 8370 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2__4848_
timestamp 0
transform -1 0 8390 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4849_
timestamp 0
transform 1 0 9050 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4850_
timestamp 0
transform 1 0 9290 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4851_
timestamp 0
transform 1 0 11270 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4852_
timestamp 0
transform 1 0 11650 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4853_
timestamp 0
transform 1 0 12050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4854_
timestamp 0
transform -1 0 11190 0 1 11770
box -6 -8 26 248
use FILL  FILL_2__4855_
timestamp 0
transform -1 0 8210 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4856_
timestamp 0
transform -1 0 8230 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4857_
timestamp 0
transform -1 0 10310 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4858_
timestamp 0
transform -1 0 10450 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4859_
timestamp 0
transform -1 0 7190 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4860_
timestamp 0
transform -1 0 10370 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4861_
timestamp 0
transform -1 0 10630 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4862_
timestamp 0
transform 1 0 11430 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4863_
timestamp 0
transform -1 0 10690 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4864_
timestamp 0
transform -1 0 10530 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4865_
timestamp 0
transform 1 0 10550 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4866_
timestamp 0
transform 1 0 11630 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4867_
timestamp 0
transform 1 0 11810 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4868_
timestamp 0
transform -1 0 11310 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4869_
timestamp 0
transform -1 0 10850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2__4870_
timestamp 0
transform 1 0 8090 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4871_
timestamp 0
transform 1 0 7930 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4872_
timestamp 0
transform 1 0 7830 0 1 7930
box -6 -8 26 248
use FILL  FILL_2__4873_
timestamp 0
transform -1 0 11350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4874_
timestamp 0
transform 1 0 11870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4875_
timestamp 0
transform -1 0 7570 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2__4876_
timestamp 0
transform -1 0 10490 0 -1 9370
box -6 -8 26 248
use FILL  FILL_2__4877_
timestamp 0
transform 1 0 10890 0 1 8410
box -6 -8 26 248
use FILL  FILL_2__4878_
timestamp 0
transform 1 0 11330 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4879_
timestamp 0
transform 1 0 11990 0 1 9850
box -6 -8 26 248
use FILL  FILL_2__4880_
timestamp 0
transform -1 0 12050 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4881_
timestamp 0
transform -1 0 9090 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4882_
timestamp 0
transform 1 0 12010 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4883_
timestamp 0
transform 1 0 11830 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4884_
timestamp 0
transform 1 0 11650 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4885_
timestamp 0
transform -1 0 11690 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4886_
timestamp 0
transform 1 0 10950 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4887_
timestamp 0
transform 1 0 10990 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4888_
timestamp 0
transform 1 0 11650 0 1 8890
box -6 -8 26 248
use FILL  FILL_2__4889_
timestamp 0
transform 1 0 11990 0 1 9370
box -6 -8 26 248
use FILL  FILL_2__4890_
timestamp 0
transform 1 0 11510 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4891_
timestamp 0
transform 1 0 11850 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2__4892_
timestamp 0
transform -1 0 12070 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2__4893_
timestamp 0
transform -1 0 2490 0 -1 7450
box -6 -8 26 248
use FILL  FILL_2__4894_
timestamp 0
transform 1 0 9690 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4895_
timestamp 0
transform 1 0 8430 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4896_
timestamp 0
transform -1 0 9470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4897_
timestamp 0
transform 1 0 9510 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4898_
timestamp 0
transform 1 0 9690 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4899_
timestamp 0
transform -1 0 9170 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4900_
timestamp 0
transform -1 0 9510 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4901_
timestamp 0
transform -1 0 9890 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4902_
timestamp 0
transform 1 0 10210 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4903_
timestamp 0
transform 1 0 9670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4904_
timestamp 0
transform -1 0 10390 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4905_
timestamp 0
transform 1 0 9670 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4906_
timestamp 0
transform -1 0 9850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4907_
timestamp 0
transform -1 0 9510 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4908_
timestamp 0
transform 1 0 10010 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4909_
timestamp 0
transform 1 0 10950 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4910_
timestamp 0
transform -1 0 11330 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4911_
timestamp 0
transform 1 0 11270 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4912_
timestamp 0
transform 1 0 11090 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4913_
timestamp 0
transform -1 0 10910 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4914_
timestamp 0
transform 1 0 11470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4915_
timestamp 0
transform -1 0 10770 0 1 6970
box -6 -8 26 248
use FILL  FILL_2__4916_
timestamp 0
transform 1 0 10530 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4917_
timestamp 0
transform -1 0 10590 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4918_
timestamp 0
transform -1 0 10950 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4919_
timestamp 0
transform 1 0 11110 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4920_
timestamp 0
transform 1 0 8530 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4921_
timestamp 0
transform -1 0 8750 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4922_
timestamp 0
transform -1 0 8950 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4923_
timestamp 0
transform 1 0 9330 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4924_
timestamp 0
transform 1 0 9310 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4925_
timestamp 0
transform -1 0 9130 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4926_
timestamp 0
transform 1 0 8890 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4927_
timestamp 0
transform -1 0 11290 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4928_
timestamp 0
transform 1 0 11470 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4929_
timestamp 0
transform 1 0 12050 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4930_
timestamp 0
transform 1 0 11630 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4931_
timestamp 0
transform -1 0 11850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4932_
timestamp 0
transform -1 0 11690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4933_
timestamp 0
transform -1 0 11130 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4934_
timestamp 0
transform 1 0 10910 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4935_
timestamp 0
transform -1 0 10730 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4936_
timestamp 0
transform -1 0 9630 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4937_
timestamp 0
transform -1 0 9850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4938_
timestamp 0
transform 1 0 10010 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4939_
timestamp 0
transform 1 0 10090 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4940_
timestamp 0
transform 1 0 10190 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2__4941_
timestamp 0
transform 1 0 10290 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4942_
timestamp 0
transform -1 0 10690 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4943_
timestamp 0
transform 1 0 11670 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4944_
timestamp 0
transform -1 0 11890 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4945_
timestamp 0
transform 1 0 11830 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4946_
timestamp 0
transform -1 0 11810 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4947_
timestamp 0
transform -1 0 8630 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4948_
timestamp 0
transform 1 0 8950 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4949_
timestamp 0
transform 1 0 12070 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__4950_
timestamp 0
transform -1 0 12030 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4951_
timestamp 0
transform -1 0 8570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4952_
timestamp 0
transform 1 0 8950 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4953_
timestamp 0
transform -1 0 8850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4954_
timestamp 0
transform -1 0 9150 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4955_
timestamp 0
transform -1 0 8710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__4956_
timestamp 0
transform -1 0 8790 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4957_
timestamp 0
transform -1 0 8650 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4958_
timestamp 0
transform -1 0 11030 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4959_
timestamp 0
transform 1 0 11210 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4960_
timestamp 0
transform -1 0 11430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4961_
timestamp 0
transform 1 0 11610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4962_
timestamp 0
transform 1 0 12010 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4963_
timestamp 0
transform 1 0 11970 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4964_
timestamp 0
transform 1 0 11970 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4965_
timestamp 0
transform -1 0 11810 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4966_
timestamp 0
transform -1 0 9150 0 1 4090
box -6 -8 26 248
use FILL  FILL_2__4967_
timestamp 0
transform 1 0 8070 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__4968_
timestamp 0
transform 1 0 11650 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4969_
timestamp 0
transform 1 0 12010 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4970_
timestamp 0
transform 1 0 9050 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4971_
timestamp 0
transform -1 0 8270 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4972_
timestamp 0
transform -1 0 8670 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4973_
timestamp 0
transform -1 0 8830 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4974_
timestamp 0
transform 1 0 8730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4975_
timestamp 0
transform 1 0 8930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4976_
timestamp 0
transform 1 0 11590 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4977_
timestamp 0
transform 1 0 11390 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4978_
timestamp 0
transform 1 0 11410 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4979_
timestamp 0
transform 1 0 11430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4980_
timestamp 0
transform 1 0 11810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4981_
timestamp 0
transform -1 0 11810 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4982_
timestamp 0
transform -1 0 11830 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4983_
timestamp 0
transform 1 0 11610 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4984_
timestamp 0
transform 1 0 11230 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4985_
timestamp 0
transform -1 0 8050 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4986_
timestamp 0
transform 1 0 9090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4987_
timestamp 0
transform 1 0 11610 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4988_
timestamp 0
transform -1 0 11830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4989_
timestamp 0
transform -1 0 11430 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4990_
timestamp 0
transform -1 0 11250 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__4991_
timestamp 0
transform 1 0 11630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__4992_
timestamp 0
transform -1 0 11490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4993_
timestamp 0
transform 1 0 11270 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__4994_
timestamp 0
transform 1 0 9290 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__4995_
timestamp 0
transform -1 0 9870 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4996_
timestamp 0
transform 1 0 9230 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4997_
timestamp 0
transform -1 0 9310 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__4998_
timestamp 0
transform 1 0 9410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__4999_
timestamp 0
transform -1 0 9270 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5000_
timestamp 0
transform 1 0 11010 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__5001_
timestamp 0
transform -1 0 10830 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__5002_
timestamp 0
transform -1 0 10650 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5003_
timestamp 0
transform -1 0 10710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5004_
timestamp 0
transform 1 0 10890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5005_
timestamp 0
transform -1 0 10870 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5006_
timestamp 0
transform 1 0 11390 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5007_
timestamp 0
transform 1 0 11990 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5008_
timestamp 0
transform 1 0 11970 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__5009_
timestamp 0
transform 1 0 11990 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5010_
timestamp 0
transform -1 0 11290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__5011_
timestamp 0
transform 1 0 11790 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5012_
timestamp 0
transform 1 0 11590 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5013_
timestamp 0
transform -1 0 10270 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5014_
timestamp 0
transform -1 0 9490 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5015_
timestamp 0
transform 1 0 8250 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5016_
timestamp 0
transform 1 0 10650 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5017_
timestamp 0
transform 1 0 8910 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5018_
timestamp 0
transform 1 0 8450 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5019_
timestamp 0
transform 1 0 9130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5020_
timestamp 0
transform 1 0 9030 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5021_
timestamp 0
transform 1 0 9310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5022_
timestamp 0
transform -1 0 9110 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5023_
timestamp 0
transform -1 0 10830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__5024_
timestamp 0
transform 1 0 10830 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5025_
timestamp 0
transform -1 0 11050 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5026_
timestamp 0
transform 1 0 11070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__5027_
timestamp 0
transform -1 0 10870 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5028_
timestamp 0
transform -1 0 10690 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5029_
timestamp 0
transform 1 0 11030 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5030_
timestamp 0
transform 1 0 11050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5031_
timestamp 0
transform 1 0 11810 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__5032_
timestamp 0
transform 1 0 11650 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__5033_
timestamp 0
transform -1 0 8970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__5034_
timestamp 0
transform -1 0 9170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__5035_
timestamp 0
transform 1 0 11190 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5036_
timestamp 0
transform 1 0 9870 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5037_
timestamp 0
transform 1 0 9670 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5038_
timestamp 0
transform 1 0 9510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5039_
timestamp 0
transform 1 0 9450 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5040_
timestamp 0
transform 1 0 9690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5041_
timestamp 0
transform 1 0 9890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5042_
timestamp 0
transform 1 0 10610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__5043_
timestamp 0
transform 1 0 10430 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5044_
timestamp 0
transform 1 0 10490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5045_
timestamp 0
transform -1 0 10470 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5046_
timestamp 0
transform 1 0 10910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__5047_
timestamp 0
transform 1 0 11010 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5048_
timestamp 0
transform 1 0 11450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__5049_
timestamp 0
transform -1 0 11290 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__5050_
timestamp 0
transform -1 0 9350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__5051_
timestamp 0
transform 1 0 8350 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__5052_
timestamp 0
transform -1 0 10510 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__5053_
timestamp 0
transform -1 0 10750 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__5054_
timestamp 0
transform -1 0 10390 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__5055_
timestamp 0
transform 1 0 8510 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__5056_
timestamp 0
transform 1 0 8130 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__5057_
timestamp 0
transform 1 0 8350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__5058_
timestamp 0
transform -1 0 8170 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__5059_
timestamp 0
transform 1 0 7990 0 1 6490
box -6 -8 26 248
use FILL  FILL_2__5060_
timestamp 0
transform -1 0 7630 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__5061_
timestamp 0
transform -1 0 7810 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__5062_
timestamp 0
transform 1 0 7970 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2__5063_
timestamp 0
transform -1 0 8010 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__5064_
timestamp 0
transform -1 0 7530 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5065_
timestamp 0
transform -1 0 7730 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5066_
timestamp 0
transform -1 0 7670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5067_
timestamp 0
transform -1 0 8370 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5068_
timestamp 0
transform -1 0 8390 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5069_
timestamp 0
transform -1 0 8230 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5070_
timestamp 0
transform -1 0 7850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5071_
timestamp 0
transform 1 0 8030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5072_
timestamp 0
transform -1 0 7490 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5073_
timestamp 0
transform 1 0 7290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5074_
timestamp 0
transform 1 0 4850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2__5075_
timestamp 0
transform 1 0 10250 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__5076_
timestamp 0
transform 1 0 10050 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__5077_
timestamp 0
transform 1 0 9830 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__5078_
timestamp 0
transform 1 0 9610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__5079_
timestamp 0
transform 1 0 10010 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__5080_
timestamp 0
transform 1 0 10210 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__5081_
timestamp 0
transform 1 0 10430 0 1 6010
box -6 -8 26 248
use FILL  FILL_2__5082_
timestamp 0
transform 1 0 10410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2__5083_
timestamp 0
transform -1 0 10310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5084_
timestamp 0
transform -1 0 9690 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5085_
timestamp 0
transform 1 0 8530 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5086_
timestamp 0
transform -1 0 8730 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5087_
timestamp 0
transform -1 0 10890 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__5088_
timestamp 0
transform -1 0 10670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__5089_
timestamp 0
transform -1 0 10470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__5090_
timestamp 0
transform -1 0 10250 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5091_
timestamp 0
transform 1 0 10090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2__5092_
timestamp 0
transform 1 0 9930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__5093_
timestamp 0
transform -1 0 10110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__5094_
timestamp 0
transform 1 0 10250 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__5095_
timestamp 0
transform -1 0 9770 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__5096_
timestamp 0
transform 1 0 8910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__5097_
timestamp 0
transform 1 0 8230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2__5098_
timestamp 0
transform 1 0 9730 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5099_
timestamp 0
transform 1 0 9910 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5100_
timestamp 0
transform 1 0 9350 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5101_
timestamp 0
transform -1 0 10070 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5102_
timestamp 0
transform -1 0 9890 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5103_
timestamp 0
transform 1 0 10030 0 1 5050
box -6 -8 26 248
use FILL  FILL_2__5104_
timestamp 0
transform -1 0 10330 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5105_
timestamp 0
transform -1 0 10130 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5106_
timestamp 0
transform -1 0 10510 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5107_
timestamp 0
transform 1 0 10490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__5108_
timestamp 0
transform -1 0 11090 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__5109_
timestamp 0
transform 1 0 10690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2__5110_
timestamp 0
transform -1 0 9550 0 1 4570
box -6 -8 26 248
use FILL  FILL_2__5111_
timestamp 0
transform -1 0 7910 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5112_
timestamp 0
transform -1 0 8090 0 1 5530
box -6 -8 26 248
use FILL  FILL_2__5124_
timestamp 0
transform 1 0 1770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__5125_
timestamp 0
transform -1 0 630 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__5126_
timestamp 0
transform -1 0 810 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__5127_
timestamp 0
transform 1 0 770 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__5128_
timestamp 0
transform 1 0 530 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__5129_
timestamp 0
transform 1 0 970 0 1 2170
box -6 -8 26 248
use FILL  FILL_2__5130_
timestamp 0
transform 1 0 970 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__5131_
timestamp 0
transform -1 0 2290 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5132_
timestamp 0
transform -1 0 5530 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5133_
timestamp 0
transform 1 0 5270 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5134_
timestamp 0
transform 1 0 1350 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__5135_
timestamp 0
transform 1 0 2150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__5136_
timestamp 0
transform 1 0 1950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__5137_
timestamp 0
transform -1 0 1090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__5138_
timestamp 0
transform -1 0 1270 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__5139_
timestamp 0
transform -1 0 3650 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5140_
timestamp 0
transform 1 0 4110 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__5141_
timestamp 0
transform -1 0 4290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__5142_
timestamp 0
transform -1 0 4170 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__5143_
timestamp 0
transform -1 0 4390 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5144_
timestamp 0
transform 1 0 5550 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5145_
timestamp 0
transform -1 0 4090 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5146_
timestamp 0
transform -1 0 4610 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5147_
timestamp 0
transform 1 0 4710 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5148_
timestamp 0
transform 1 0 4910 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5149_
timestamp 0
transform 1 0 5430 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5150_
timestamp 0
transform -1 0 6050 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5151_
timestamp 0
transform 1 0 3430 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5152_
timestamp 0
transform 1 0 5690 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5153_
timestamp 0
transform 1 0 4170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__5154_
timestamp 0
transform 1 0 5370 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5155_
timestamp 0
transform 1 0 5330 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5156_
timestamp 0
transform 1 0 5490 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5157_
timestamp 0
transform 1 0 5630 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5158_
timestamp 0
transform 1 0 4510 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5159_
timestamp 0
transform -1 0 4630 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5160_
timestamp 0
transform 1 0 4950 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5161_
timestamp 0
transform 1 0 4790 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5162_
timestamp 0
transform 1 0 5830 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5163_
timestamp 0
transform -1 0 2730 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5164_
timestamp 0
transform 1 0 5850 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5165_
timestamp 0
transform -1 0 3790 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__5166_
timestamp 0
transform 1 0 4230 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5167_
timestamp 0
transform 1 0 4190 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5168_
timestamp 0
transform -1 0 4010 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5169_
timestamp 0
transform 1 0 2690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__5170_
timestamp 0
transform 1 0 3810 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5171_
timestamp 0
transform -1 0 4110 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__5172_
timestamp 0
transform -1 0 3610 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__5173_
timestamp 0
transform -1 0 4890 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__5174_
timestamp 0
transform -1 0 3790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__5175_
timestamp 0
transform 1 0 3630 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5176_
timestamp 0
transform -1 0 2630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__5177_
timestamp 0
transform 1 0 3070 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5178_
timestamp 0
transform 1 0 4410 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5179_
timestamp 0
transform 1 0 4430 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5180_
timestamp 0
transform 1 0 4230 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5181_
timestamp 0
transform 1 0 3230 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5182_
timestamp 0
transform -1 0 2430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__5183_
timestamp 0
transform 1 0 2230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__5184_
timestamp 0
transform -1 0 2450 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__5185_
timestamp 0
transform -1 0 4010 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__5186_
timestamp 0
transform -1 0 3290 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__5187_
timestamp 0
transform -1 0 3030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__5188_
timestamp 0
transform 1 0 3730 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5189_
timestamp 0
transform -1 0 3670 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5190_
timestamp 0
transform 1 0 3210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__5191_
timestamp 0
transform 1 0 2890 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5192_
timestamp 0
transform -1 0 3610 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__5193_
timestamp 0
transform 1 0 6050 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5194_
timestamp 0
transform -1 0 2910 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__5195_
timestamp 0
transform -1 0 2830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__5196_
timestamp 0
transform 1 0 3570 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5197_
timestamp 0
transform -1 0 3490 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5198_
timestamp 0
transform -1 0 2890 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5199_
timestamp 0
transform 1 0 2450 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5200_
timestamp 0
transform -1 0 2670 0 -1 730
box -6 -8 26 248
use FILL  FILL_2__5201_
timestamp 0
transform -1 0 3950 0 1 1690
box -6 -8 26 248
use FILL  FILL_2__5202_
timestamp 0
transform 1 0 3910 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5203_
timestamp 0
transform -1 0 3450 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5204_
timestamp 0
transform 1 0 4070 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5205_
timestamp 0
transform -1 0 3910 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5206_
timestamp 0
transform -1 0 3250 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5207_
timestamp 0
transform 1 0 2470 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5208_
timestamp 0
transform 1 0 3010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__5209_
timestamp 0
transform -1 0 4470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2__5210_
timestamp 0
transform 1 0 2670 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5211_
timestamp 0
transform 1 0 2830 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5212_
timestamp 0
transform 1 0 3410 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5213_
timestamp 0
transform 1 0 3290 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5214_
timestamp 0
transform -1 0 3050 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5215_
timestamp 0
transform 1 0 2270 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5216_
timestamp 0
transform -1 0 3070 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__5217_
timestamp 0
transform -1 0 6230 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5218_
timestamp 0
transform 1 0 3410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__5219_
timestamp 0
transform 1 0 3570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__5220_
timestamp 0
transform 1 0 4750 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5221_
timestamp 0
transform 1 0 4570 0 -1 250
box -6 -8 26 248
use FILL  FILL_2__5222_
timestamp 0
transform -1 0 4050 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5223_
timestamp 0
transform 1 0 3090 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5224_
timestamp 0
transform -1 0 3850 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5225_
timestamp 0
transform 1 0 5350 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__5226_
timestamp 0
transform 1 0 5130 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5227_
timestamp 0
transform -1 0 5310 0 1 250
box -6 -8 26 248
use FILL  FILL_2__5228_
timestamp 0
transform -1 0 4750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2__5229_
timestamp 0
transform -1 0 4790 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5230_
timestamp 0
transform 1 0 4970 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5231_
timestamp 0
transform 1 0 5170 0 1 730
box -6 -8 26 248
use FILL  FILL_2__5232_
timestamp 0
transform 1 0 3970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2__5233_
timestamp 0
transform 1 0 4350 0 1 1210
box -6 -8 26 248
use FILL  FILL_2__5234_
timestamp 0
transform -1 0 5150 0 1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert0
timestamp 0
transform -1 0 4190 0 1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert1
timestamp 0
transform 1 0 6110 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert2
timestamp 0
transform -1 0 3290 0 1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert3
timestamp 0
transform -1 0 3670 0 1 9850
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert4
timestamp 0
transform 1 0 9450 0 1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert5
timestamp 0
transform 1 0 11250 0 1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert6
timestamp 0
transform -1 0 9450 0 1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert7
timestamp 0
transform 1 0 11990 0 1 7930
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert8
timestamp 0
transform -1 0 7150 0 1 5530
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert9
timestamp 0
transform 1 0 6650 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert10
timestamp 0
transform 1 0 8690 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert11
timestamp 0
transform 1 0 6850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert12
timestamp 0
transform 1 0 8890 0 1 9850
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert13
timestamp 0
transform 1 0 7370 0 1 9850
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert14
timestamp 0
transform 1 0 630 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert15
timestamp 0
transform 1 0 50 0 1 9370
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert16
timestamp 0
transform 1 0 1870 0 1 5530
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert17
timestamp 0
transform -1 0 9130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert18
timestamp 0
transform -1 0 11490 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert19
timestamp 0
transform 1 0 10650 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert20
timestamp 0
transform -1 0 9170 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert21
timestamp 0
transform 1 0 2510 0 1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert22
timestamp 0
transform -1 0 1250 0 1 11290
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert23
timestamp 0
transform -1 0 1430 0 1 11290
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert24
timestamp 0
transform -1 0 1630 0 1 10330
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert38
timestamp 0
transform -1 0 11510 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert39
timestamp 0
transform -1 0 10650 0 1 6010
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert40
timestamp 0
transform 1 0 12010 0 1 6970
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert41
timestamp 0
transform -1 0 11230 0 1 6010
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert42
timestamp 0
transform 1 0 11430 0 1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert43
timestamp 0
transform -1 0 10990 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert44
timestamp 0
transform -1 0 10470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert45
timestamp 0
transform -1 0 11350 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert46
timestamp 0
transform -1 0 10730 0 1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert47
timestamp 0
transform 1 0 6190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert48
timestamp 0
transform -1 0 4750 0 1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert49
timestamp 0
transform 1 0 11550 0 1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert50
timestamp 0
transform -1 0 10390 0 1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert51
timestamp 0
transform 1 0 8150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert52
timestamp 0
transform 1 0 10010 0 1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert53
timestamp 0
transform 1 0 9170 0 1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert54
timestamp 0
transform 1 0 8990 0 1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert55
timestamp 0
transform -1 0 9530 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert56
timestamp 0
transform -1 0 8830 0 1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert57
timestamp 0
transform 1 0 11450 0 1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert58
timestamp 0
transform 1 0 10630 0 -1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert59
timestamp 0
transform -1 0 7710 0 -1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert60
timestamp 0
transform 1 0 11790 0 -1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert61
timestamp 0
transform 1 0 11890 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert62
timestamp 0
transform -1 0 4790 0 1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert63
timestamp 0
transform -1 0 9310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert64
timestamp 0
transform -1 0 11650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert65
timestamp 0
transform -1 0 9310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert66
timestamp 0
transform -1 0 11490 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert67
timestamp 0
transform 1 0 6910 0 1 11290
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert68
timestamp 0
transform -1 0 3150 0 -1 10330
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert69
timestamp 0
transform -1 0 5610 0 1 10810
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert70
timestamp 0
transform 1 0 5090 0 -1 11290
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert71
timestamp 0
transform -1 0 3550 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert72
timestamp 0
transform 1 0 7090 0 1 11290
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert73
timestamp 0
transform 1 0 7110 0 1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert74
timestamp 0
transform -1 0 6450 0 1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert75
timestamp 0
transform 1 0 7070 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert76
timestamp 0
transform 1 0 6530 0 1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert77
timestamp 0
transform 1 0 10250 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert78
timestamp 0
transform 1 0 9110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert79
timestamp 0
transform 1 0 10270 0 1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert80
timestamp 0
transform -1 0 4930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert81
timestamp 0
transform -1 0 2790 0 1 5530
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert82
timestamp 0
transform -1 0 4010 0 -1 5530
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert83
timestamp 0
transform -1 0 6270 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert84
timestamp 0
transform 1 0 7330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert85
timestamp 0
transform -1 0 3250 0 1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert86
timestamp 0
transform 1 0 3950 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert87
timestamp 0
transform -1 0 3210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert88
timestamp 0
transform 1 0 7870 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert89
timestamp 0
transform -1 0 4710 0 1 9850
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert90
timestamp 0
transform 1 0 5550 0 1 9370
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert91
timestamp 0
transform 1 0 9010 0 1 10330
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert92
timestamp 0
transform -1 0 8510 0 1 10810
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert93
timestamp 0
transform -1 0 10910 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert94
timestamp 0
transform 1 0 7250 0 1 10330
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert95
timestamp 0
transform 1 0 11510 0 1 10810
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert96
timestamp 0
transform -1 0 4970 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert97
timestamp 0
transform 1 0 590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert98
timestamp 0
transform -1 0 3990 0 1 7930
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert99
timestamp 0
transform 1 0 530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert100
timestamp 0
transform 1 0 3010 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert101
timestamp 0
transform -1 0 470 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert102
timestamp 0
transform 1 0 3710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert103
timestamp 0
transform -1 0 3630 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert104
timestamp 0
transform 1 0 4610 0 1 10330
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert105
timestamp 0
transform 1 0 270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert106
timestamp 0
transform 1 0 6490 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert107
timestamp 0
transform -1 0 6190 0 1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert108
timestamp 0
transform 1 0 5670 0 1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert109
timestamp 0
transform 1 0 7810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert110
timestamp 0
transform -1 0 5310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert111
timestamp 0
transform 1 0 7270 0 1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert112
timestamp 0
transform 1 0 10650 0 1 11770
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert113
timestamp 0
transform -1 0 12090 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert114
timestamp 0
transform -1 0 10290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert115
timestamp 0
transform 1 0 7350 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert116
timestamp 0
transform -1 0 5490 0 1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert117
timestamp 0
transform -1 0 5470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert118
timestamp 0
transform -1 0 11170 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert119
timestamp 0
transform 1 0 10350 0 1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert120
timestamp 0
transform -1 0 11090 0 1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert121
timestamp 0
transform -1 0 8150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert122
timestamp 0
transform 1 0 11170 0 1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert123
timestamp 0
transform -1 0 10010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert124
timestamp 0
transform -1 0 7990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert125
timestamp 0
transform -1 0 5310 0 1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert126
timestamp 0
transform 1 0 11990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert127
timestamp 0
transform 1 0 10750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert128
timestamp 0
transform -1 0 12030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert129
timestamp 0
transform 1 0 10430 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert130
timestamp 0
transform 1 0 11990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert131
timestamp 0
transform -1 0 9350 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert132
timestamp 0
transform -1 0 8690 0 1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert133
timestamp 0
transform 1 0 11990 0 1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert134
timestamp 0
transform -1 0 11370 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert135
timestamp 0
transform -1 0 9090 0 -1 250
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert136
timestamp 0
transform 1 0 9450 0 -1 250
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert137
timestamp 0
transform -1 0 6370 0 1 730
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert138
timestamp 0
transform 1 0 8350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert139
timestamp 0
transform -1 0 6390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert140
timestamp 0
transform 1 0 9410 0 1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert141
timestamp 0
transform -1 0 7030 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert142
timestamp 0
transform -1 0 7010 0 1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert143
timestamp 0
transform -1 0 6430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert144
timestamp 0
transform -1 0 6250 0 1 6970
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert145
timestamp 0
transform 1 0 9530 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert146
timestamp 0
transform 1 0 9630 0 1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert147
timestamp 0
transform -1 0 7710 0 1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert148
timestamp 0
transform -1 0 7630 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert149
timestamp 0
transform -1 0 9210 0 -1 7930
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert150
timestamp 0
transform -1 0 7210 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert151
timestamp 0
transform 1 0 7310 0 -1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert152
timestamp 0
transform -1 0 8210 0 1 9370
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert153
timestamp 0
transform 1 0 10050 0 -1 9850
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert154
timestamp 0
transform 1 0 10730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert155
timestamp 0
transform 1 0 6370 0 1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert156
timestamp 0
transform 1 0 9110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert157
timestamp 0
transform -1 0 5850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert158
timestamp 0
transform 1 0 9850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert159
timestamp 0
transform 1 0 8710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert160
timestamp 0
transform 1 0 10350 0 1 9850
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert161
timestamp 0
transform 1 0 9250 0 1 9850
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert162
timestamp 0
transform 1 0 10210 0 1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert163
timestamp 0
transform -1 0 8310 0 1 8890
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert164
timestamp 0
transform 1 0 11710 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert165
timestamp 0
transform -1 0 8770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert166
timestamp 0
transform -1 0 11550 0 1 4090
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert167
timestamp 0
transform 1 0 11710 0 1 11770
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert168
timestamp 0
transform -1 0 11290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_BUFX2_insert169
timestamp 0
transform 1 0 4910 0 1 1690
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert25
timestamp 0
transform 1 0 1350 0 1 2170
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert26
timestamp 0
transform 1 0 4010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert27
timestamp 0
transform -1 0 70 0 -1 2650
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert28
timestamp 0
transform -1 0 2710 0 1 9370
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert29
timestamp 0
transform 1 0 50 0 -1 2170
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert30
timestamp 0
transform 1 0 6170 0 -1 5050
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert31
timestamp 0
transform 1 0 770 0 -1 6010
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert32
timestamp 0
transform -1 0 4810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert33
timestamp 0
transform -1 0 950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert34
timestamp 0
transform 1 0 1390 0 -1 6490
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert35
timestamp 0
transform -1 0 310 0 -1 11770
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert36
timestamp 0
transform 1 0 50 0 1 5530
box -6 -8 26 248
use FILL  FILL_2_CLKBUF1_insert37
timestamp 0
transform 1 0 6130 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__2478_
timestamp 0
transform -1 0 90 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2479_
timestamp 0
transform -1 0 90 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2480_
timestamp 0
transform 1 0 1930 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2481_
timestamp 0
transform 1 0 2750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2482_
timestamp 0
transform -1 0 90 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__2483_
timestamp 0
transform -1 0 570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__2484_
timestamp 0
transform -1 0 2130 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2485_
timestamp 0
transform 1 0 3950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2486_
timestamp 0
transform 1 0 12070 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2487_
timestamp 0
transform -1 0 6650 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2488_
timestamp 0
transform -1 0 6830 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2489_
timestamp 0
transform 1 0 12030 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2490_
timestamp 0
transform 1 0 12030 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2491_
timestamp 0
transform 1 0 6450 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2492_
timestamp 0
transform 1 0 11850 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2493_
timestamp 0
transform -1 0 11950 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2494_
timestamp 0
transform -1 0 1050 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__2495_
timestamp 0
transform -1 0 1210 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2496_
timestamp 0
transform -1 0 90 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__2497_
timestamp 0
transform -1 0 4430 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2498_
timestamp 0
transform 1 0 4470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2499_
timestamp 0
transform -1 0 3290 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2500_
timestamp 0
transform -1 0 470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2501_
timestamp 0
transform -1 0 3670 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2502_
timestamp 0
transform -1 0 90 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__2503_
timestamp 0
transform -1 0 90 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2504_
timestamp 0
transform 1 0 4570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2505_
timestamp 0
transform 1 0 5110 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2506_
timestamp 0
transform -1 0 2550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2507_
timestamp 0
transform 1 0 3830 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2508_
timestamp 0
transform 1 0 3450 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2509_
timestamp 0
transform 1 0 4230 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2510_
timestamp 0
transform 1 0 3090 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2511_
timestamp 0
transform -1 0 4950 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2519_
timestamp 0
transform -1 0 5690 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2520_
timestamp 0
transform -1 0 7550 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2521_
timestamp 0
transform -1 0 7750 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2522_
timestamp 0
transform 1 0 7750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2523_
timestamp 0
transform 1 0 9490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2524_
timestamp 0
transform -1 0 7810 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2525_
timestamp 0
transform 1 0 7550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2526_
timestamp 0
transform 1 0 8290 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2527_
timestamp 0
transform 1 0 8490 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2528_
timestamp 0
transform -1 0 9630 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2529_
timestamp 0
transform 1 0 8570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2530_
timestamp 0
transform -1 0 8210 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2531_
timestamp 0
transform -1 0 8350 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2532_
timestamp 0
transform -1 0 8770 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2533_
timestamp 0
transform 1 0 9510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2534_
timestamp 0
transform 1 0 10070 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__2535_
timestamp 0
transform -1 0 10270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2536_
timestamp 0
transform -1 0 8770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2537_
timestamp 0
transform -1 0 8570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2538_
timestamp 0
transform -1 0 8370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2539_
timestamp 0
transform 1 0 7970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2540_
timestamp 0
transform -1 0 10670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2541_
timestamp 0
transform -1 0 10870 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2542_
timestamp 0
transform 1 0 10910 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2543_
timestamp 0
transform -1 0 10610 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2544_
timestamp 0
transform -1 0 5710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2545_
timestamp 0
transform -1 0 5910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2546_
timestamp 0
transform -1 0 6130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2547_
timestamp 0
transform -1 0 6010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2548_
timestamp 0
transform -1 0 6210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2549_
timestamp 0
transform 1 0 5590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2550_
timestamp 0
transform 1 0 5790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2551_
timestamp 0
transform -1 0 6910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2552_
timestamp 0
transform -1 0 7270 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2553_
timestamp 0
transform -1 0 5730 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2554_
timestamp 0
transform -1 0 6370 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2555_
timestamp 0
transform 1 0 6410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2556_
timestamp 0
transform -1 0 6750 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2557_
timestamp 0
transform -1 0 6230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2558_
timestamp 0
transform 1 0 6510 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2559_
timestamp 0
transform 1 0 6890 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2560_
timestamp 0
transform -1 0 5930 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2561_
timestamp 0
transform -1 0 6570 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2562_
timestamp 0
transform 1 0 6750 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2563_
timestamp 0
transform -1 0 6130 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2564_
timestamp 0
transform 1 0 7790 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2565_
timestamp 0
transform 1 0 8010 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2566_
timestamp 0
transform 1 0 7590 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2567_
timestamp 0
transform 1 0 6990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2568_
timestamp 0
transform -1 0 6630 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2569_
timestamp 0
transform 1 0 7210 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2570_
timestamp 0
transform -1 0 9390 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2571_
timestamp 0
transform -1 0 9290 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2572_
timestamp 0
transform 1 0 9310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2573_
timestamp 0
transform 1 0 9190 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2574_
timestamp 0
transform -1 0 9270 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2575_
timestamp 0
transform -1 0 9090 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2576_
timestamp 0
transform -1 0 8810 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2577_
timestamp 0
transform -1 0 9010 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2578_
timestamp 0
transform 1 0 9570 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2579_
timestamp 0
transform -1 0 9510 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2580_
timestamp 0
transform -1 0 8310 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2581_
timestamp 0
transform 1 0 8270 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2582_
timestamp 0
transform 1 0 8390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2583_
timestamp 0
transform -1 0 9790 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2584_
timestamp 0
transform 1 0 9450 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2585_
timestamp 0
transform -1 0 11190 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2586_
timestamp 0
transform 1 0 8870 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2587_
timestamp 0
transform 1 0 8670 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2588_
timestamp 0
transform -1 0 8490 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2589_
timestamp 0
transform 1 0 8530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2590_
timestamp 0
transform 1 0 8270 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2591_
timestamp 0
transform -1 0 8610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2592_
timestamp 0
transform 1 0 7870 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2593_
timestamp 0
transform -1 0 9110 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2594_
timestamp 0
transform -1 0 9010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2595_
timestamp 0
transform -1 0 9270 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2596_
timestamp 0
transform 1 0 10450 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2597_
timestamp 0
transform 1 0 10630 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2598_
timestamp 0
transform -1 0 10470 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2599_
timestamp 0
transform 1 0 10830 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2600_
timestamp 0
transform -1 0 11430 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2601_
timestamp 0
transform 1 0 8290 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2602_
timestamp 0
transform -1 0 8090 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2603_
timestamp 0
transform 1 0 7090 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2604_
timestamp 0
transform 1 0 8250 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2605_
timestamp 0
transform -1 0 8130 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2606_
timestamp 0
transform -1 0 7730 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2607_
timestamp 0
transform -1 0 6590 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2608_
timestamp 0
transform 1 0 6770 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2609_
timestamp 0
transform 1 0 6970 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2610_
timestamp 0
transform -1 0 7910 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2611_
timestamp 0
transform -1 0 10130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2612_
timestamp 0
transform 1 0 9910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2613_
timestamp 0
transform 1 0 10310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2614_
timestamp 0
transform -1 0 11010 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__2615_
timestamp 0
transform -1 0 7190 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2616_
timestamp 0
transform 1 0 8330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2617_
timestamp 0
transform -1 0 7190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2618_
timestamp 0
transform -1 0 6530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2619_
timestamp 0
transform 1 0 6310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2620_
timestamp 0
transform -1 0 8010 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2621_
timestamp 0
transform -1 0 8110 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2622_
timestamp 0
transform 1 0 8370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2623_
timestamp 0
transform -1 0 8970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2624_
timestamp 0
transform 1 0 8110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2625_
timestamp 0
transform 1 0 6870 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2626_
timestamp 0
transform -1 0 8330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2627_
timestamp 0
transform 1 0 9930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2628_
timestamp 0
transform 1 0 11550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2629_
timestamp 0
transform 1 0 11450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2630_
timestamp 0
transform 1 0 11730 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2631_
timestamp 0
transform -1 0 11550 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2632_
timestamp 0
transform 1 0 9450 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2633_
timestamp 0
transform -1 0 8550 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2634_
timestamp 0
transform 1 0 8950 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2635_
timestamp 0
transform -1 0 9190 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2636_
timestamp 0
transform -1 0 9970 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2637_
timestamp 0
transform -1 0 8670 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2638_
timestamp 0
transform 1 0 9750 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2639_
timestamp 0
transform 1 0 10010 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2640_
timestamp 0
transform 1 0 8130 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2641_
timestamp 0
transform 1 0 7930 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2642_
timestamp 0
transform 1 0 9410 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2643_
timestamp 0
transform 1 0 9410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2644_
timestamp 0
transform 1 0 8430 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2645_
timestamp 0
transform 1 0 7650 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2646_
timestamp 0
transform 1 0 7450 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2647_
timestamp 0
transform 1 0 8230 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2648_
timestamp 0
transform -1 0 8070 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2649_
timestamp 0
transform -1 0 9070 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2650_
timestamp 0
transform 1 0 11130 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2651_
timestamp 0
transform -1 0 9270 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2652_
timestamp 0
transform -1 0 8570 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2653_
timestamp 0
transform 1 0 8750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2654_
timestamp 0
transform 1 0 5870 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2655_
timestamp 0
transform -1 0 6090 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2656_
timestamp 0
transform -1 0 6270 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2657_
timestamp 0
transform -1 0 7670 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2658_
timestamp 0
transform 1 0 7430 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2659_
timestamp 0
transform -1 0 7190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2660_
timestamp 0
transform -1 0 7370 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2661_
timestamp 0
transform -1 0 10810 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2662_
timestamp 0
transform 1 0 10990 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2663_
timestamp 0
transform 1 0 10050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2664_
timestamp 0
transform 1 0 10230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2665_
timestamp 0
transform -1 0 6650 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2666_
timestamp 0
transform 1 0 7230 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2667_
timestamp 0
transform -1 0 7030 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2668_
timestamp 0
transform -1 0 6850 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2669_
timestamp 0
transform 1 0 6770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2670_
timestamp 0
transform -1 0 10630 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2671_
timestamp 0
transform 1 0 11690 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2672_
timestamp 0
transform 1 0 11730 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2673_
timestamp 0
transform -1 0 11530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2674_
timestamp 0
transform 1 0 11470 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2675_
timestamp 0
transform -1 0 10830 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2676_
timestamp 0
transform 1 0 11450 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2677_
timestamp 0
transform -1 0 11530 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2678_
timestamp 0
transform -1 0 10150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2679_
timestamp 0
transform 1 0 9750 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2680_
timestamp 0
transform 1 0 9670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2681_
timestamp 0
transform 1 0 9350 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2682_
timestamp 0
transform -1 0 9570 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2683_
timestamp 0
transform -1 0 10230 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2684_
timestamp 0
transform -1 0 10530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2685_
timestamp 0
transform -1 0 10810 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__2686_
timestamp 0
transform 1 0 10710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2687_
timestamp 0
transform -1 0 9830 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2688_
timestamp 0
transform 1 0 9230 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2689_
timestamp 0
transform 1 0 10550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2690_
timestamp 0
transform -1 0 10910 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2691_
timestamp 0
transform -1 0 11110 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2692_
timestamp 0
transform 1 0 11290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2693_
timestamp 0
transform -1 0 10450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2694_
timestamp 0
transform 1 0 9650 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2695_
timestamp 0
transform -1 0 10570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2696_
timestamp 0
transform 1 0 10330 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2697_
timestamp 0
transform 1 0 9990 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2698_
timestamp 0
transform 1 0 9970 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2699_
timestamp 0
transform 1 0 9090 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2700_
timestamp 0
transform 1 0 8870 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2701_
timestamp 0
transform -1 0 8510 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2702_
timestamp 0
transform 1 0 8870 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2703_
timestamp 0
transform 1 0 10890 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2704_
timestamp 0
transform -1 0 9150 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2705_
timestamp 0
transform -1 0 9710 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2706_
timestamp 0
transform -1 0 10110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2707_
timestamp 0
transform -1 0 9630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2708_
timestamp 0
transform 1 0 8930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2709_
timestamp 0
transform 1 0 9050 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2710_
timestamp 0
transform -1 0 8750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2711_
timestamp 0
transform -1 0 10810 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2712_
timestamp 0
transform -1 0 10790 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2713_
timestamp 0
transform 1 0 10830 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2714_
timestamp 0
transform 1 0 10830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2715_
timestamp 0
transform -1 0 11470 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2716_
timestamp 0
transform 1 0 11630 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2717_
timestamp 0
transform -1 0 10750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2718_
timestamp 0
transform 1 0 11090 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2719_
timestamp 0
transform 1 0 11810 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2720_
timestamp 0
transform -1 0 11010 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2721_
timestamp 0
transform -1 0 10910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2722_
timestamp 0
transform -1 0 10950 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2723_
timestamp 0
transform 1 0 11390 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2724_
timestamp 0
transform 1 0 11370 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2725_
timestamp 0
transform 1 0 10350 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2726_
timestamp 0
transform -1 0 9730 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2727_
timestamp 0
transform 1 0 9930 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2728_
timestamp 0
transform -1 0 9910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2729_
timestamp 0
transform -1 0 9510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2730_
timestamp 0
transform 1 0 11250 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2731_
timestamp 0
transform 1 0 9490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2732_
timestamp 0
transform 1 0 6710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2733_
timestamp 0
transform -1 0 9130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2734_
timestamp 0
transform 1 0 9490 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2735_
timestamp 0
transform 1 0 9510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2736_
timestamp 0
transform -1 0 8930 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2737_
timestamp 0
transform -1 0 9310 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2738_
timestamp 0
transform -1 0 10390 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2739_
timestamp 0
transform 1 0 10570 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2740_
timestamp 0
transform 1 0 11190 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2741_
timestamp 0
transform 1 0 11590 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2742_
timestamp 0
transform -1 0 10590 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2743_
timestamp 0
transform -1 0 10430 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2744_
timestamp 0
transform 1 0 10510 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2745_
timestamp 0
transform -1 0 11170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2746_
timestamp 0
transform -1 0 10170 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2747_
timestamp 0
transform 1 0 10970 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2748_
timestamp 0
transform 1 0 9830 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2749_
timestamp 0
transform 1 0 10690 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2750_
timestamp 0
transform 1 0 11030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2751_
timestamp 0
transform -1 0 10150 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2752_
timestamp 0
transform 1 0 5770 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2753_
timestamp 0
transform -1 0 5990 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2754_
timestamp 0
transform -1 0 6050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2755_
timestamp 0
transform -1 0 7410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2756_
timestamp 0
transform -1 0 7530 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2757_
timestamp 0
transform 1 0 8130 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2758_
timestamp 0
transform -1 0 7590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2759_
timestamp 0
transform -1 0 9730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2760_
timestamp 0
transform -1 0 6250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2761_
timestamp 0
transform -1 0 8890 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2762_
timestamp 0
transform -1 0 8870 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2763_
timestamp 0
transform -1 0 6330 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2764_
timestamp 0
transform -1 0 6410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2765_
timestamp 0
transform -1 0 9370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2766_
timestamp 0
transform -1 0 6710 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2767_
timestamp 0
transform 1 0 8930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2768_
timestamp 0
transform -1 0 6010 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2769_
timestamp 0
transform -1 0 6950 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2770_
timestamp 0
transform 1 0 7130 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2771_
timestamp 0
transform 1 0 10050 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2772_
timestamp 0
transform -1 0 7410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2773_
timestamp 0
transform -1 0 7610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2774_
timestamp 0
transform -1 0 6050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2775_
timestamp 0
transform -1 0 7350 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2776_
timestamp 0
transform 1 0 6170 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2777_
timestamp 0
transform -1 0 9890 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2778_
timestamp 0
transform 1 0 7710 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2779_
timestamp 0
transform 1 0 7930 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2780_
timestamp 0
transform 1 0 7990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2781_
timestamp 0
transform -1 0 7810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2782_
timestamp 0
transform 1 0 7670 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2783_
timestamp 0
transform -1 0 8470 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2784_
timestamp 0
transform -1 0 11010 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2785_
timestamp 0
transform 1 0 9530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2786_
timestamp 0
transform -1 0 7790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2787_
timestamp 0
transform -1 0 9230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2788_
timestamp 0
transform -1 0 10210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2789_
timestamp 0
transform 1 0 10390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2790_
timestamp 0
transform 1 0 7990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2791_
timestamp 0
transform 1 0 8190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2792_
timestamp 0
transform -1 0 7650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2793_
timestamp 0
transform -1 0 7870 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2794_
timestamp 0
transform -1 0 7870 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2795_
timestamp 0
transform -1 0 7590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2796_
timestamp 0
transform -1 0 6990 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2797_
timestamp 0
transform -1 0 8410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2798_
timestamp 0
transform 1 0 11950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2799_
timestamp 0
transform -1 0 7370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2800_
timestamp 0
transform -1 0 7490 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2801_
timestamp 0
transform 1 0 7130 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2802_
timestamp 0
transform 1 0 6790 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2803_
timestamp 0
transform -1 0 7010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2804_
timestamp 0
transform -1 0 8510 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2805_
timestamp 0
transform 1 0 6930 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2806_
timestamp 0
transform -1 0 6830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2807_
timestamp 0
transform -1 0 7090 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2808_
timestamp 0
transform 1 0 10170 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2809_
timestamp 0
transform -1 0 10590 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2810_
timestamp 0
transform 1 0 10570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2811_
timestamp 0
transform 1 0 10390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2812_
timestamp 0
transform 1 0 10250 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2813_
timestamp 0
transform -1 0 10090 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2814_
timestamp 0
transform -1 0 10490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2815_
timestamp 0
transform -1 0 10690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2816_
timestamp 0
transform 1 0 10210 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2817_
timestamp 0
transform -1 0 10310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2818_
timestamp 0
transform -1 0 10970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2819_
timestamp 0
transform -1 0 11070 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2820_
timestamp 0
transform -1 0 11270 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2821_
timestamp 0
transform 1 0 11030 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2822_
timestamp 0
transform -1 0 11970 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2823_
timestamp 0
transform 1 0 11150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2824_
timestamp 0
transform 1 0 10650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2825_
timestamp 0
transform 1 0 11170 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2826_
timestamp 0
transform 1 0 11370 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2827_
timestamp 0
transform -1 0 11830 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2828_
timestamp 0
transform -1 0 11950 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2829_
timestamp 0
transform -1 0 11390 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2830_
timestamp 0
transform 1 0 11030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2831_
timestamp 0
transform 1 0 11090 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2832_
timestamp 0
transform -1 0 11330 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2833_
timestamp 0
transform 1 0 11390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2834_
timestamp 0
transform 1 0 11890 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2835_
timestamp 0
transform 1 0 12070 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__2836_
timestamp 0
transform 1 0 11690 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2837_
timestamp 0
transform 1 0 11890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2838_
timestamp 0
transform 1 0 12010 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2839_
timestamp 0
transform 1 0 11590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2840_
timestamp 0
transform -1 0 11790 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2841_
timestamp 0
transform -1 0 11650 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2842_
timestamp 0
transform -1 0 9830 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2843_
timestamp 0
transform -1 0 10030 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2844_
timestamp 0
transform -1 0 11810 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2845_
timestamp 0
transform 1 0 11990 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2846_
timestamp 0
transform 1 0 11550 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__2847_
timestamp 0
transform 1 0 11970 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2848_
timestamp 0
transform -1 0 11610 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2849_
timestamp 0
transform -1 0 11710 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2850_
timestamp 0
transform 1 0 11890 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2851_
timestamp 0
transform -1 0 9890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2852_
timestamp 0
transform -1 0 11070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2853_
timestamp 0
transform 1 0 11250 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2854_
timestamp 0
transform 1 0 11830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2855_
timestamp 0
transform 1 0 11830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2856_
timestamp 0
transform -1 0 9850 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2857_
timestamp 0
transform -1 0 9910 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2858_
timestamp 0
transform -1 0 8070 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2859_
timestamp 0
transform 1 0 9690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2860_
timestamp 0
transform -1 0 9150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2861_
timestamp 0
transform 1 0 9970 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2862_
timestamp 0
transform 1 0 9570 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2863_
timestamp 0
transform 1 0 8790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2864_
timestamp 0
transform -1 0 7790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2865_
timestamp 0
transform -1 0 6450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2866_
timestamp 0
transform -1 0 8870 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2867_
timestamp 0
transform -1 0 9410 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2868_
timestamp 0
transform 1 0 9210 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2869_
timestamp 0
transform -1 0 10570 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2870_
timestamp 0
transform -1 0 9330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2871_
timestamp 0
transform -1 0 8570 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2872_
timestamp 0
transform 1 0 9770 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2873_
timestamp 0
transform 1 0 9810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2874_
timestamp 0
transform 1 0 9610 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2875_
timestamp 0
transform -1 0 11210 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__2876_
timestamp 0
transform 1 0 10210 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2877_
timestamp 0
transform -1 0 10750 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2878_
timestamp 0
transform 1 0 9650 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2879_
timestamp 0
transform -1 0 9870 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2880_
timestamp 0
transform -1 0 10190 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2881_
timestamp 0
transform -1 0 5970 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2882_
timestamp 0
transform -1 0 6150 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2883_
timestamp 0
transform -1 0 5510 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2884_
timestamp 0
transform -1 0 5510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2885_
timestamp 0
transform 1 0 5490 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2886_
timestamp 0
transform -1 0 5310 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__2887_
timestamp 0
transform 1 0 5650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2888_
timestamp 0
transform 1 0 6070 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2889_
timestamp 0
transform -1 0 6310 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2890_
timestamp 0
transform -1 0 6690 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2891_
timestamp 0
transform 1 0 8170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2892_
timestamp 0
transform -1 0 7290 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2893_
timestamp 0
transform -1 0 5890 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2894_
timestamp 0
transform 1 0 5390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2895_
timestamp 0
transform -1 0 7490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2896_
timestamp 0
transform -1 0 6610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__2897_
timestamp 0
transform 1 0 7350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2898_
timestamp 0
transform 1 0 11770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2899_
timestamp 0
transform -1 0 6550 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2900_
timestamp 0
transform -1 0 6750 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2901_
timestamp 0
transform -1 0 8190 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2902_
timestamp 0
transform 1 0 9650 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2903_
timestamp 0
transform -1 0 11590 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2904_
timestamp 0
transform 1 0 8370 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2905_
timestamp 0
transform -1 0 6950 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2906_
timestamp 0
transform -1 0 7330 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2907_
timestamp 0
transform -1 0 6350 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2908_
timestamp 0
transform 1 0 8470 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2909_
timestamp 0
transform -1 0 10370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2910_
timestamp 0
transform 1 0 10770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2911_
timestamp 0
transform 1 0 10950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2912_
timestamp 0
transform -1 0 10810 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2913_
timestamp 0
transform -1 0 8690 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2914_
timestamp 0
transform -1 0 8570 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2915_
timestamp 0
transform -1 0 11250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2916_
timestamp 0
transform -1 0 7990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2917_
timestamp 0
transform -1 0 7010 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2918_
timestamp 0
transform 1 0 6790 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2919_
timestamp 0
transform -1 0 7210 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2920_
timestamp 0
transform 1 0 7170 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2921_
timestamp 0
transform 1 0 6970 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2922_
timestamp 0
transform 1 0 6630 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2923_
timestamp 0
transform -1 0 5850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2924_
timestamp 0
transform 1 0 8890 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2925_
timestamp 0
transform 1 0 10250 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2926_
timestamp 0
transform 1 0 11990 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2927_
timestamp 0
transform 1 0 8710 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2928_
timestamp 0
transform 1 0 7510 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2929_
timestamp 0
transform 1 0 8230 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2930_
timestamp 0
transform -1 0 8450 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2931_
timestamp 0
transform -1 0 8090 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2932_
timestamp 0
transform 1 0 7890 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2933_
timestamp 0
transform 1 0 7930 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2934_
timestamp 0
transform -1 0 10230 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2935_
timestamp 0
transform 1 0 11350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__2936_
timestamp 0
transform -1 0 8210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2937_
timestamp 0
transform 1 0 8690 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2938_
timestamp 0
transform -1 0 11810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2939_
timestamp 0
transform -1 0 11250 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2940_
timestamp 0
transform -1 0 6590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2941_
timestamp 0
transform 1 0 8870 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2942_
timestamp 0
transform 1 0 8950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2943_
timestamp 0
transform 1 0 9710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2944_
timestamp 0
transform 1 0 9890 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__2945_
timestamp 0
transform 1 0 9070 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2946_
timestamp 0
transform -1 0 9170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2947_
timestamp 0
transform -1 0 8730 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2948_
timestamp 0
transform -1 0 8670 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2949_
timestamp 0
transform 1 0 10850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2950_
timestamp 0
transform 1 0 11670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2951_
timestamp 0
transform -1 0 6990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2952_
timestamp 0
transform -1 0 6790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2953_
timestamp 0
transform 1 0 11290 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2954_
timestamp 0
transform -1 0 8970 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2955_
timestamp 0
transform -1 0 10110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__2956_
timestamp 0
transform -1 0 11370 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2957_
timestamp 0
transform 1 0 9690 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2958_
timestamp 0
transform 1 0 11650 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__2959_
timestamp 0
transform 1 0 5130 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2960_
timestamp 0
transform -1 0 7390 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2961_
timestamp 0
transform -1 0 7990 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2962_
timestamp 0
transform -1 0 7590 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2963_
timestamp 0
transform -1 0 6510 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__2964_
timestamp 0
transform -1 0 7790 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2965_
timestamp 0
transform -1 0 11770 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__2966_
timestamp 0
transform 1 0 8590 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2967_
timestamp 0
transform 1 0 9290 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__2968_
timestamp 0
transform 1 0 10410 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2969_
timestamp 0
transform 1 0 10610 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__2970_
timestamp 0
transform -1 0 11290 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2971_
timestamp 0
transform 1 0 7750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2972_
timestamp 0
transform -1 0 9350 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2973_
timestamp 0
transform 1 0 7390 0 1 250
box -6 -8 26 248
use FILL  FILL_3__2974_
timestamp 0
transform -1 0 7330 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2975_
timestamp 0
transform -1 0 9090 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__2976_
timestamp 0
transform 1 0 10070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2977_
timestamp 0
transform 1 0 10470 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2978_
timestamp 0
transform -1 0 11630 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__2979_
timestamp 0
transform -1 0 11870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__2980_
timestamp 0
transform 1 0 7190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2981_
timestamp 0
transform 1 0 6590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__2982_
timestamp 0
transform 1 0 7530 0 1 730
box -6 -8 26 248
use FILL  FILL_3__2983_
timestamp 0
transform 1 0 11910 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__2984_
timestamp 0
transform 1 0 11650 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__2985_
timestamp 0
transform -1 0 7150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__2986_
timestamp 0
transform -1 0 7170 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__2987_
timestamp 0
transform 1 0 5830 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__3000_
timestamp 0
transform -1 0 2230 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3001_
timestamp 0
transform 1 0 2370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3002_
timestamp 0
transform 1 0 2170 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__3003_
timestamp 0
transform -1 0 3650 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__3004_
timestamp 0
transform 1 0 3850 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__3005_
timestamp 0
transform -1 0 3490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__3006_
timestamp 0
transform -1 0 4370 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__3007_
timestamp 0
transform -1 0 4170 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__3008_
timestamp 0
transform 1 0 3890 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__3009_
timestamp 0
transform 1 0 3990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3010_
timestamp 0
transform -1 0 4010 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__3011_
timestamp 0
transform 1 0 3810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3012_
timestamp 0
transform 1 0 2750 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__3013_
timestamp 0
transform -1 0 2450 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3014_
timestamp 0
transform 1 0 2590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__3015_
timestamp 0
transform -1 0 4570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3016_
timestamp 0
transform 1 0 4490 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__3017_
timestamp 0
transform 1 0 4190 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3018_
timestamp 0
transform 1 0 4390 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3019_
timestamp 0
transform -1 0 4010 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3020_
timestamp 0
transform 1 0 1830 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3021_
timestamp 0
transform 1 0 1670 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3022_
timestamp 0
transform -1 0 2070 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3023_
timestamp 0
transform -1 0 2910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3024_
timestamp 0
transform 1 0 4730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3025_
timestamp 0
transform 1 0 4350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3026_
timestamp 0
transform 1 0 3610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3027_
timestamp 0
transform 1 0 3310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__3028_
timestamp 0
transform -1 0 2810 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__3029_
timestamp 0
transform 1 0 3450 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3030_
timestamp 0
transform 1 0 4890 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__3031_
timestamp 0
transform 1 0 4730 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__3032_
timestamp 0
transform 1 0 5890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3033_
timestamp 0
transform -1 0 4610 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3034_
timestamp 0
transform 1 0 3830 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3035_
timestamp 0
transform -1 0 4590 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__3036_
timestamp 0
transform -1 0 2390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__3037_
timestamp 0
transform -1 0 3330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__3038_
timestamp 0
transform 1 0 2210 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__3039_
timestamp 0
transform -1 0 3590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3040_
timestamp 0
transform -1 0 3810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3041_
timestamp 0
transform 1 0 3410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3042_
timestamp 0
transform -1 0 2790 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3043_
timestamp 0
transform -1 0 3830 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__3044_
timestamp 0
transform -1 0 2630 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3045_
timestamp 0
transform -1 0 2930 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__3046_
timestamp 0
transform -1 0 3270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3047_
timestamp 0
transform 1 0 2870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3048_
timestamp 0
transform 1 0 3410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__3049_
timestamp 0
transform -1 0 3710 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__3050_
timestamp 0
transform -1 0 2950 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__3051_
timestamp 0
transform -1 0 2970 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__3052_
timestamp 0
transform 1 0 3130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__3053_
timestamp 0
transform -1 0 3010 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3054_
timestamp 0
transform -1 0 2610 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__3055_
timestamp 0
transform -1 0 2430 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__3056_
timestamp 0
transform -1 0 2750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3057_
timestamp 0
transform -1 0 3270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3058_
timestamp 0
transform 1 0 4190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3059_
timestamp 0
transform -1 0 5110 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__3060_
timestamp 0
transform -1 0 5310 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__3061_
timestamp 0
transform -1 0 6070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3062_
timestamp 0
transform -1 0 5130 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__3063_
timestamp 0
transform -1 0 5150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__3064_
timestamp 0
transform -1 0 4990 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3076_
timestamp 0
transform 1 0 1090 0 1 250
box -6 -8 26 248
use FILL  FILL_3__3077_
timestamp 0
transform -1 0 1310 0 1 250
box -6 -8 26 248
use FILL  FILL_3__3078_
timestamp 0
transform 1 0 930 0 1 250
box -6 -8 26 248
use FILL  FILL_3__3079_
timestamp 0
transform 1 0 1010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__3080_
timestamp 0
transform -1 0 890 0 1 730
box -6 -8 26 248
use FILL  FILL_3__3081_
timestamp 0
transform 1 0 830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__3082_
timestamp 0
transform 1 0 1410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__3083_
timestamp 0
transform -1 0 1570 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__3084_
timestamp 0
transform 1 0 1490 0 1 250
box -6 -8 26 248
use FILL  FILL_3__3085_
timestamp 0
transform -1 0 1770 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__3086_
timestamp 0
transform -1 0 470 0 1 730
box -6 -8 26 248
use FILL  FILL_3__3087_
timestamp 0
transform -1 0 650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__3088_
timestamp 0
transform 1 0 450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__3089_
timestamp 0
transform -1 0 1430 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__3090_
timestamp 0
transform 1 0 1230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3091_
timestamp 0
transform -1 0 1910 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__3092_
timestamp 0
transform -1 0 690 0 1 730
box -6 -8 26 248
use FILL  FILL_3__3093_
timestamp 0
transform -1 0 90 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__3094_
timestamp 0
transform -1 0 90 0 1 730
box -6 -8 26 248
use FILL  FILL_3__3095_
timestamp 0
transform -1 0 290 0 1 730
box -6 -8 26 248
use FILL  FILL_3__3096_
timestamp 0
transform -1 0 290 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__3097_
timestamp 0
transform 1 0 2050 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__3098_
timestamp 0
transform -1 0 2350 0 1 250
box -6 -8 26 248
use FILL  FILL_3__3099_
timestamp 0
transform 1 0 1910 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__3100_
timestamp 0
transform 1 0 70 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3101_
timestamp 0
transform -1 0 90 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__3102_
timestamp 0
transform -1 0 1270 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__3103_
timestamp 0
transform -1 0 1230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__3104_
timestamp 0
transform -1 0 270 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__3105_
timestamp 0
transform -1 0 1190 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__3106_
timestamp 0
transform -1 0 2350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__3107_
timestamp 0
transform -1 0 1550 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__3108_
timestamp 0
transform -1 0 430 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3109_
timestamp 0
transform -1 0 610 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3110_
timestamp 0
transform 1 0 750 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__3111_
timestamp 0
transform -1 0 950 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__3112_
timestamp 0
transform -1 0 90 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__3113_
timestamp 0
transform -1 0 90 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3114_
timestamp 0
transform -1 0 4590 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__3115_
timestamp 0
transform -1 0 4650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3116_
timestamp 0
transform 1 0 4510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__3117_
timestamp 0
transform 1 0 550 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__3118_
timestamp 0
transform -1 0 1710 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__3119_
timestamp 0
transform 1 0 890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3120_
timestamp 0
transform 1 0 1050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3121_
timestamp 0
transform -1 0 2370 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3122_
timestamp 0
transform -1 0 470 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__3123_
timestamp 0
transform 1 0 350 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__3124_
timestamp 0
transform 1 0 250 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__3125_
timestamp 0
transform 1 0 2070 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__3126_
timestamp 0
transform -1 0 2290 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__3127_
timestamp 0
transform 1 0 1590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3128_
timestamp 0
transform 1 0 1430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3129_
timestamp 0
transform 1 0 4770 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__3130_
timestamp 0
transform 1 0 4950 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__3131_
timestamp 0
transform 1 0 5170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__3132_
timestamp 0
transform 1 0 4830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3133_
timestamp 0
transform -1 0 4730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__3134_
timestamp 0
transform -1 0 4370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__3135_
timestamp 0
transform 1 0 730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__3136_
timestamp 0
transform -1 0 790 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__3137_
timestamp 0
transform 1 0 390 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__3138_
timestamp 0
transform 1 0 730 0 1 250
box -6 -8 26 248
use FILL  FILL_3__3139_
timestamp 0
transform 1 0 250 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__3140_
timestamp 0
transform -1 0 1550 0 1 730
box -6 -8 26 248
use FILL  FILL_3__3141_
timestamp 0
transform 1 0 1730 0 1 730
box -6 -8 26 248
use FILL  FILL_3__3142_
timestamp 0
transform -1 0 1710 0 1 250
box -6 -8 26 248
use FILL  FILL_3__3143_
timestamp 0
transform 1 0 2410 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__3144_
timestamp 0
transform 1 0 2530 0 1 250
box -6 -8 26 248
use FILL  FILL_3__3145_
timestamp 0
transform 1 0 2250 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__3146_
timestamp 0
transform -1 0 1950 0 1 730
box -6 -8 26 248
use FILL  FILL_3__3147_
timestamp 0
transform 1 0 2050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__3148_
timestamp 0
transform 1 0 1090 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__3149_
timestamp 0
transform -1 0 930 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__3150_
timestamp 0
transform -1 0 290 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__3151_
timestamp 0
transform 1 0 70 0 1 250
box -6 -8 26 248
use FILL  FILL_3__3152_
timestamp 0
transform -1 0 2150 0 1 730
box -6 -8 26 248
use FILL  FILL_3__3284_
timestamp 0
transform -1 0 4750 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__3285_
timestamp 0
transform 1 0 4390 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__3286_
timestamp 0
transform -1 0 3430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3287_
timestamp 0
transform 1 0 3290 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3288_
timestamp 0
transform 1 0 2210 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3289_
timestamp 0
transform 1 0 2410 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3290_
timestamp 0
transform -1 0 2090 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3291_
timestamp 0
transform 1 0 3030 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3292_
timestamp 0
transform 1 0 3230 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3293_
timestamp 0
transform 1 0 5850 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3294_
timestamp 0
transform -1 0 5890 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3295_
timestamp 0
transform 1 0 5930 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3296_
timestamp 0
transform 1 0 6410 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3297_
timestamp 0
transform 1 0 6610 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3298_
timestamp 0
transform 1 0 5310 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3299_
timestamp 0
transform 1 0 5510 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3300_
timestamp 0
transform 1 0 4650 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3301_
timestamp 0
transform 1 0 4850 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3302_
timestamp 0
transform -1 0 3410 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3303_
timestamp 0
transform -1 0 3570 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3304_
timestamp 0
transform -1 0 3450 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3305_
timestamp 0
transform -1 0 3630 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3306_
timestamp 0
transform 1 0 4370 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3307_
timestamp 0
transform 1 0 4470 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3308_
timestamp 0
transform -1 0 1130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3309_
timestamp 0
transform -1 0 1050 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__3310_
timestamp 0
transform 1 0 2530 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3311_
timestamp 0
transform -1 0 2750 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3312_
timestamp 0
transform 1 0 3470 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3313_
timestamp 0
transform -1 0 2390 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3314_
timestamp 0
transform -1 0 270 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__3315_
timestamp 0
transform -1 0 470 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__3316_
timestamp 0
transform -1 0 7550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__3317_
timestamp 0
transform 1 0 6170 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3318_
timestamp 0
transform 1 0 2650 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3319_
timestamp 0
transform 1 0 6670 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3320_
timestamp 0
transform 1 0 5450 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3321_
timestamp 0
transform -1 0 6470 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__3322_
timestamp 0
transform -1 0 3830 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3323_
timestamp 0
transform -1 0 3670 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3324_
timestamp 0
transform 1 0 5170 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3325_
timestamp 0
transform -1 0 5390 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3326_
timestamp 0
transform -1 0 5250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__3327_
timestamp 0
transform 1 0 4830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__3328_
timestamp 0
transform -1 0 5290 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3329_
timestamp 0
transform -1 0 5710 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__3330_
timestamp 0
transform 1 0 5570 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3331_
timestamp 0
transform 1 0 4990 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3332_
timestamp 0
transform -1 0 4670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__3333_
timestamp 0
transform -1 0 5970 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3334_
timestamp 0
transform 1 0 5950 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__3335_
timestamp 0
transform -1 0 470 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3336_
timestamp 0
transform -1 0 290 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3337_
timestamp 0
transform -1 0 910 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3338_
timestamp 0
transform -1 0 930 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3339_
timestamp 0
transform -1 0 5890 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__3340_
timestamp 0
transform 1 0 6070 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__3341_
timestamp 0
transform -1 0 5850 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3342_
timestamp 0
transform -1 0 5470 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3343_
timestamp 0
transform -1 0 4390 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3344_
timestamp 0
transform -1 0 5510 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__3345_
timestamp 0
transform 1 0 5690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__3346_
timestamp 0
transform 1 0 5290 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__3347_
timestamp 0
transform 1 0 5110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__3348_
timestamp 0
transform -1 0 90 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3349_
timestamp 0
transform 1 0 270 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3350_
timestamp 0
transform 1 0 7790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__3351_
timestamp 0
transform -1 0 90 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3352_
timestamp 0
transform 1 0 310 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3353_
timestamp 0
transform -1 0 1830 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3354_
timestamp 0
transform 1 0 2010 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3355_
timestamp 0
transform -1 0 330 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3356_
timestamp 0
transform -1 0 530 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3357_
timestamp 0
transform -1 0 870 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3358_
timestamp 0
transform -1 0 850 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3359_
timestamp 0
transform -1 0 90 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3360_
timestamp 0
transform -1 0 290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__3361_
timestamp 0
transform -1 0 4890 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3362_
timestamp 0
transform -1 0 5010 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3363_
timestamp 0
transform 1 0 5330 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3364_
timestamp 0
transform -1 0 3430 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3365_
timestamp 0
transform 1 0 3350 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3366_
timestamp 0
transform 1 0 2930 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3367_
timestamp 0
transform 1 0 2570 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3368_
timestamp 0
transform 1 0 2370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3369_
timestamp 0
transform -1 0 4150 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3370_
timestamp 0
transform -1 0 5310 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3371_
timestamp 0
transform -1 0 7070 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3372_
timestamp 0
transform 1 0 5110 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3373_
timestamp 0
transform -1 0 7510 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3374_
timestamp 0
transform -1 0 7290 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3375_
timestamp 0
transform -1 0 4690 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3376_
timestamp 0
transform -1 0 4730 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3377_
timestamp 0
transform 1 0 4910 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3378_
timestamp 0
transform -1 0 4330 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3379_
timestamp 0
transform 1 0 5770 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3380_
timestamp 0
transform -1 0 7830 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3381_
timestamp 0
transform 1 0 6670 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3382_
timestamp 0
transform 1 0 6490 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3383_
timestamp 0
transform -1 0 7090 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3384_
timestamp 0
transform -1 0 6890 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3385_
timestamp 0
transform 1 0 7270 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3386_
timestamp 0
transform -1 0 6530 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3387_
timestamp 0
transform 1 0 6310 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3388_
timestamp 0
transform 1 0 6730 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3389_
timestamp 0
transform -1 0 7130 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3390_
timestamp 0
transform -1 0 9730 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3391_
timestamp 0
transform -1 0 10270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3392_
timestamp 0
transform -1 0 270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3393_
timestamp 0
transform 1 0 250 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3394_
timestamp 0
transform -1 0 250 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3395_
timestamp 0
transform -1 0 270 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3396_
timestamp 0
transform -1 0 90 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3397_
timestamp 0
transform -1 0 1250 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3398_
timestamp 0
transform 1 0 1030 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3399_
timestamp 0
transform 1 0 990 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3400_
timestamp 0
transform -1 0 630 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3401_
timestamp 0
transform -1 0 90 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3402_
timestamp 0
transform -1 0 850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3403_
timestamp 0
transform 1 0 1610 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3404_
timestamp 0
transform -1 0 910 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3405_
timestamp 0
transform 1 0 710 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3406_
timestamp 0
transform -1 0 1890 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3407_
timestamp 0
transform -1 0 490 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__3408_
timestamp 0
transform 1 0 270 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__3409_
timestamp 0
transform -1 0 90 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__3410_
timestamp 0
transform -1 0 910 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3411_
timestamp 0
transform -1 0 450 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3412_
timestamp 0
transform -1 0 270 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3413_
timestamp 0
transform -1 0 90 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3414_
timestamp 0
transform -1 0 250 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3415_
timestamp 0
transform -1 0 90 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3416_
timestamp 0
transform -1 0 90 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3417_
timestamp 0
transform -1 0 430 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3418_
timestamp 0
transform -1 0 6950 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3419_
timestamp 0
transform 1 0 6250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3420_
timestamp 0
transform 1 0 6050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3421_
timestamp 0
transform 1 0 5290 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3422_
timestamp 0
transform 1 0 5150 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3423_
timestamp 0
transform 1 0 7130 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3424_
timestamp 0
transform -1 0 1390 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3425_
timestamp 0
transform 1 0 630 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3426_
timestamp 0
transform 1 0 430 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3427_
timestamp 0
transform -1 0 450 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3428_
timestamp 0
transform -1 0 290 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3429_
timestamp 0
transform 1 0 610 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3430_
timestamp 0
transform -1 0 90 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3431_
timestamp 0
transform -1 0 270 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3432_
timestamp 0
transform 1 0 890 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3433_
timestamp 0
transform 1 0 1490 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3434_
timestamp 0
transform -1 0 990 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3435_
timestamp 0
transform -1 0 1110 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3436_
timestamp 0
transform 1 0 1290 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3437_
timestamp 0
transform -1 0 1330 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__3438_
timestamp 0
transform -1 0 1010 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3439_
timestamp 0
transform -1 0 810 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3440_
timestamp 0
transform -1 0 1130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__3441_
timestamp 0
transform 1 0 730 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3442_
timestamp 0
transform 1 0 830 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3443_
timestamp 0
transform -1 0 810 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3444_
timestamp 0
transform -1 0 630 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3445_
timestamp 0
transform -1 0 750 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__3446_
timestamp 0
transform -1 0 1410 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3447_
timestamp 0
transform -1 0 1190 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3448_
timestamp 0
transform -1 0 730 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3449_
timestamp 0
transform 1 0 1350 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3450_
timestamp 0
transform 1 0 1530 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3451_
timestamp 0
transform -1 0 2650 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3452_
timestamp 0
transform -1 0 2850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3453_
timestamp 0
transform -1 0 3070 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3454_
timestamp 0
transform -1 0 1190 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__3455_
timestamp 0
transform -1 0 290 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3456_
timestamp 0
transform -1 0 90 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3457_
timestamp 0
transform -1 0 850 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3458_
timestamp 0
transform 1 0 630 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3459_
timestamp 0
transform -1 0 570 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__3460_
timestamp 0
transform 1 0 470 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3461_
timestamp 0
transform -1 0 1910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3462_
timestamp 0
transform 1 0 1690 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3463_
timestamp 0
transform -1 0 1950 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__3464_
timestamp 0
transform -1 0 2070 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3465_
timestamp 0
transform -1 0 1650 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3466_
timestamp 0
transform -1 0 2030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__3467_
timestamp 0
transform -1 0 1890 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3468_
timestamp 0
transform -1 0 2290 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3469_
timestamp 0
transform -1 0 290 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3470_
timestamp 0
transform -1 0 1230 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3471_
timestamp 0
transform -1 0 1210 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3472_
timestamp 0
transform -1 0 1590 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3473_
timestamp 0
transform 1 0 1770 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3474_
timestamp 0
transform -1 0 2070 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3475_
timestamp 0
transform -1 0 1750 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3476_
timestamp 0
transform -1 0 1710 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3477_
timestamp 0
transform -1 0 1890 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3478_
timestamp 0
transform 1 0 1970 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3479_
timestamp 0
transform -1 0 1430 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3480_
timestamp 0
transform -1 0 2830 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3481_
timestamp 0
transform -1 0 6070 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3482_
timestamp 0
transform -1 0 5890 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3483_
timestamp 0
transform 1 0 6730 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3484_
timestamp 0
transform -1 0 7490 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__3485_
timestamp 0
transform -1 0 7290 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__3486_
timestamp 0
transform 1 0 5750 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__3487_
timestamp 0
transform -1 0 5770 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3488_
timestamp 0
transform 1 0 2990 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3489_
timestamp 0
transform -1 0 6130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__3490_
timestamp 0
transform 1 0 1550 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3491_
timestamp 0
transform 1 0 1370 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3492_
timestamp 0
transform 1 0 1930 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3493_
timestamp 0
transform -1 0 1770 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3494_
timestamp 0
transform 1 0 7210 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3495_
timestamp 0
transform -1 0 7590 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3496_
timestamp 0
transform -1 0 7790 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3497_
timestamp 0
transform -1 0 8210 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3498_
timestamp 0
transform -1 0 7430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3499_
timestamp 0
transform 1 0 1170 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__3500_
timestamp 0
transform 1 0 1370 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__3501_
timestamp 0
transform -1 0 3150 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3502_
timestamp 0
transform -1 0 3750 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3503_
timestamp 0
transform -1 0 3250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3504_
timestamp 0
transform 1 0 2950 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__3505_
timestamp 0
transform 1 0 3150 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__3506_
timestamp 0
transform -1 0 770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__3507_
timestamp 0
transform -1 0 970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__3508_
timestamp 0
transform 1 0 6370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__3509_
timestamp 0
transform -1 0 6610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__3510_
timestamp 0
transform 1 0 6830 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__3511_
timestamp 0
transform -1 0 6650 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__3512_
timestamp 0
transform 1 0 6590 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__3513_
timestamp 0
transform 1 0 6770 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__3514_
timestamp 0
transform -1 0 6510 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3515_
timestamp 0
transform 1 0 7170 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__3516_
timestamp 0
transform -1 0 1230 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3517_
timestamp 0
transform 1 0 1010 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3518_
timestamp 0
transform -1 0 7490 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3519_
timestamp 0
transform -1 0 7310 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3520_
timestamp 0
transform 1 0 5330 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3521_
timestamp 0
transform -1 0 5530 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3522_
timestamp 0
transform -1 0 90 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__3523_
timestamp 0
transform 1 0 250 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3524_
timestamp 0
transform -1 0 470 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__3525_
timestamp 0
transform 1 0 2050 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__3526_
timestamp 0
transform 1 0 2230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__3527_
timestamp 0
transform 1 0 7030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__3528_
timestamp 0
transform -1 0 6970 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__3529_
timestamp 0
transform -1 0 90 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3530_
timestamp 0
transform 1 0 10110 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3531_
timestamp 0
transform 1 0 6070 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3532_
timestamp 0
transform 1 0 5690 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3533_
timestamp 0
transform 1 0 11850 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3534_
timestamp 0
transform -1 0 9150 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3535_
timestamp 0
transform 1 0 7650 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3536_
timestamp 0
transform 1 0 6050 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__3537_
timestamp 0
transform 1 0 5590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3538_
timestamp 0
transform 1 0 5570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3539_
timestamp 0
transform 1 0 6170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3540_
timestamp 0
transform 1 0 6370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3541_
timestamp 0
transform -1 0 6250 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3542_
timestamp 0
transform -1 0 6070 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3543_
timestamp 0
transform 1 0 5970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3544_
timestamp 0
transform 1 0 5850 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3545_
timestamp 0
transform 1 0 5850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3546_
timestamp 0
transform -1 0 6230 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__3547_
timestamp 0
transform 1 0 6390 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3548_
timestamp 0
transform 1 0 6490 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3549_
timestamp 0
transform 1 0 6690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3550_
timestamp 0
transform 1 0 6550 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3551_
timestamp 0
transform -1 0 6750 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3552_
timestamp 0
transform 1 0 6830 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3553_
timestamp 0
transform -1 0 7270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__3554_
timestamp 0
transform 1 0 11230 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3555_
timestamp 0
transform 1 0 10890 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3556_
timestamp 0
transform 1 0 10150 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3557_
timestamp 0
transform -1 0 9230 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3558_
timestamp 0
transform -1 0 10730 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3559_
timestamp 0
transform 1 0 11570 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3560_
timestamp 0
transform 1 0 10030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3561_
timestamp 0
transform 1 0 10010 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3562_
timestamp 0
transform 1 0 9810 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3563_
timestamp 0
transform -1 0 9890 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3564_
timestamp 0
transform -1 0 11830 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3565_
timestamp 0
transform 1 0 12010 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3566_
timestamp 0
transform 1 0 11430 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3567_
timestamp 0
transform 1 0 11070 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3568_
timestamp 0
transform 1 0 11210 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3569_
timestamp 0
transform 1 0 9750 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3570_
timestamp 0
transform 1 0 10650 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3571_
timestamp 0
transform 1 0 9570 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3572_
timestamp 0
transform -1 0 9410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3573_
timestamp 0
transform 1 0 11010 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3574_
timestamp 0
transform -1 0 9350 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3575_
timestamp 0
transform 1 0 8550 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3576_
timestamp 0
transform -1 0 8030 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3577_
timestamp 0
transform -1 0 9010 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3578_
timestamp 0
transform -1 0 9090 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3579_
timestamp 0
transform -1 0 8210 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3580_
timestamp 0
transform -1 0 8670 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3581_
timestamp 0
transform 1 0 9610 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3582_
timestamp 0
transform 1 0 9410 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3583_
timestamp 0
transform 1 0 8470 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3584_
timestamp 0
transform -1 0 8410 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3585_
timestamp 0
transform 1 0 9130 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3586_
timestamp 0
transform -1 0 8970 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3587_
timestamp 0
transform -1 0 9210 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3588_
timestamp 0
transform 1 0 8210 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3589_
timestamp 0
transform -1 0 9030 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3590_
timestamp 0
transform -1 0 10610 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3591_
timestamp 0
transform -1 0 10770 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3592_
timestamp 0
transform 1 0 8230 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3593_
timestamp 0
transform -1 0 6210 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3594_
timestamp 0
transform -1 0 10370 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3595_
timestamp 0
transform -1 0 10530 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3596_
timestamp 0
transform 1 0 6970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3597_
timestamp 0
transform 1 0 6630 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3598_
timestamp 0
transform 1 0 11850 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3599_
timestamp 0
transform -1 0 8910 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3600_
timestamp 0
transform 1 0 8690 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3601_
timestamp 0
transform 1 0 8830 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3602_
timestamp 0
transform -1 0 9950 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3603_
timestamp 0
transform -1 0 10270 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3604_
timestamp 0
transform -1 0 8430 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3605_
timestamp 0
transform -1 0 7870 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3606_
timestamp 0
transform -1 0 8010 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3607_
timestamp 0
transform 1 0 7810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3608_
timestamp 0
transform 1 0 11410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3609_
timestamp 0
transform 1 0 11630 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3610_
timestamp 0
transform 1 0 11490 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3611_
timestamp 0
transform 1 0 11290 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3612_
timestamp 0
transform 1 0 11650 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3613_
timestamp 0
transform 1 0 11390 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3614_
timestamp 0
transform 1 0 11590 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3615_
timestamp 0
transform 1 0 11330 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3616_
timestamp 0
transform -1 0 8110 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3617_
timestamp 0
transform 1 0 12030 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3618_
timestamp 0
transform 1 0 11970 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3619_
timestamp 0
transform -1 0 11550 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3620_
timestamp 0
transform 1 0 8790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3621_
timestamp 0
transform 1 0 8170 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3622_
timestamp 0
transform 1 0 8130 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3623_
timestamp 0
transform 1 0 11130 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3624_
timestamp 0
transform -1 0 11110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3625_
timestamp 0
transform 1 0 10790 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3626_
timestamp 0
transform 1 0 10990 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3627_
timestamp 0
transform 1 0 10930 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3628_
timestamp 0
transform 1 0 7970 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3629_
timestamp 0
transform 1 0 7630 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3630_
timestamp 0
transform 1 0 7610 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3631_
timestamp 0
transform -1 0 7470 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3632_
timestamp 0
transform 1 0 7030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3633_
timestamp 0
transform 1 0 8030 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3634_
timestamp 0
transform 1 0 8710 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3635_
timestamp 0
transform 1 0 8370 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3636_
timestamp 0
transform -1 0 6850 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3637_
timestamp 0
transform 1 0 8730 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3638_
timestamp 0
transform 1 0 10830 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3639_
timestamp 0
transform 1 0 8590 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3640_
timestamp 0
transform 1 0 9450 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3641_
timestamp 0
transform 1 0 8950 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3642_
timestamp 0
transform -1 0 7310 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3643_
timestamp 0
transform 1 0 7110 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3644_
timestamp 0
transform -1 0 9330 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3645_
timestamp 0
transform -1 0 10410 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3646_
timestamp 0
transform 1 0 9110 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3647_
timestamp 0
transform 1 0 10550 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3648_
timestamp 0
transform 1 0 10870 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3649_
timestamp 0
transform 1 0 10970 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3650_
timestamp 0
transform -1 0 11390 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3651_
timestamp 0
transform 1 0 6770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3652_
timestamp 0
transform 1 0 4830 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3653_
timestamp 0
transform 1 0 4630 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3654_
timestamp 0
transform 1 0 4430 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3655_
timestamp 0
transform 1 0 4230 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3656_
timestamp 0
transform 1 0 5430 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3657_
timestamp 0
transform 1 0 5390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3658_
timestamp 0
transform 1 0 5230 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3659_
timestamp 0
transform 1 0 4650 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3660_
timestamp 0
transform 1 0 4450 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3661_
timestamp 0
transform 1 0 4830 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3662_
timestamp 0
transform 1 0 6570 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3663_
timestamp 0
transform 1 0 6370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3664_
timestamp 0
transform 1 0 5610 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3665_
timestamp 0
transform 1 0 5210 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3666_
timestamp 0
transform 1 0 5810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3667_
timestamp 0
transform -1 0 3690 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3668_
timestamp 0
transform 1 0 3910 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3669_
timestamp 0
transform -1 0 3410 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3670_
timestamp 0
transform -1 0 3530 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3671_
timestamp 0
transform 1 0 4170 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3672_
timestamp 0
transform 1 0 4230 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3673_
timestamp 0
transform 1 0 5990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3674_
timestamp 0
transform -1 0 10730 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3675_
timestamp 0
transform -1 0 10550 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3676_
timestamp 0
transform 1 0 4150 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3677_
timestamp 0
transform -1 0 4210 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3678_
timestamp 0
transform 1 0 4650 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3679_
timestamp 0
transform -1 0 4870 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3680_
timestamp 0
transform -1 0 5070 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3681_
timestamp 0
transform -1 0 4770 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3682_
timestamp 0
transform 1 0 1650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__3683_
timestamp 0
transform 1 0 6270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3684_
timestamp 0
transform 1 0 6610 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3685_
timestamp 0
transform 1 0 6890 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3686_
timestamp 0
transform 1 0 6670 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3687_
timestamp 0
transform 1 0 4890 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3688_
timestamp 0
transform -1 0 4910 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3689_
timestamp 0
transform 1 0 5090 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3690_
timestamp 0
transform -1 0 4750 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3691_
timestamp 0
transform -1 0 4690 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3692_
timestamp 0
transform 1 0 4490 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3693_
timestamp 0
transform 1 0 4870 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3694_
timestamp 0
transform -1 0 6070 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3695_
timestamp 0
transform 1 0 1710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3696_
timestamp 0
transform 1 0 7590 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3697_
timestamp 0
transform 1 0 7790 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3698_
timestamp 0
transform 1 0 6690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3699_
timestamp 0
transform 1 0 6890 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3700_
timestamp 0
transform -1 0 7090 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3701_
timestamp 0
transform 1 0 4650 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__3702_
timestamp 0
transform 1 0 4350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3703_
timestamp 0
transform 1 0 4410 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3704_
timestamp 0
transform 1 0 4830 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3705_
timestamp 0
transform -1 0 4910 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3706_
timestamp 0
transform -1 0 4690 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__3707_
timestamp 0
transform -1 0 5030 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3708_
timestamp 0
transform 1 0 4610 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3709_
timestamp 0
transform 1 0 2470 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3710_
timestamp 0
transform 1 0 9790 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3711_
timestamp 0
transform 1 0 9670 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3712_
timestamp 0
transform 1 0 9650 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3713_
timestamp 0
transform 1 0 10030 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3714_
timestamp 0
transform 1 0 8730 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3715_
timestamp 0
transform -1 0 8930 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3716_
timestamp 0
transform -1 0 9530 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3717_
timestamp 0
transform -1 0 10430 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3718_
timestamp 0
transform 1 0 10590 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3719_
timestamp 0
transform -1 0 9130 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3720_
timestamp 0
transform 1 0 9310 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3721_
timestamp 0
transform -1 0 10650 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3722_
timestamp 0
transform -1 0 10470 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3723_
timestamp 0
transform 1 0 10790 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3724_
timestamp 0
transform 1 0 9470 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3725_
timestamp 0
transform 1 0 8330 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3726_
timestamp 0
transform -1 0 8210 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3727_
timestamp 0
transform 1 0 9650 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3728_
timestamp 0
transform -1 0 10210 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3729_
timestamp 0
transform 1 0 10050 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3730_
timestamp 0
transform 1 0 10010 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3731_
timestamp 0
transform 1 0 8450 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3732_
timestamp 0
transform 1 0 8830 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3733_
timestamp 0
transform -1 0 3890 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3734_
timestamp 0
transform -1 0 4070 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3735_
timestamp 0
transform 1 0 7650 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3736_
timestamp 0
transform -1 0 7250 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3737_
timestamp 0
transform -1 0 5810 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3738_
timestamp 0
transform 1 0 9590 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3739_
timestamp 0
transform 1 0 9390 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3740_
timestamp 0
transform 1 0 9270 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3741_
timestamp 0
transform -1 0 10770 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3742_
timestamp 0
transform 1 0 11270 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3743_
timestamp 0
transform 1 0 11450 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3744_
timestamp 0
transform 1 0 11190 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3745_
timestamp 0
transform -1 0 10610 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3746_
timestamp 0
transform -1 0 10270 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3747_
timestamp 0
transform -1 0 10210 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3748_
timestamp 0
transform -1 0 10950 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3749_
timestamp 0
transform -1 0 11270 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3750_
timestamp 0
transform 1 0 11070 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3751_
timestamp 0
transform -1 0 8070 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3752_
timestamp 0
transform -1 0 6870 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3753_
timestamp 0
transform -1 0 6770 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3754_
timestamp 0
transform 1 0 4410 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3755_
timestamp 0
transform 1 0 3050 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3756_
timestamp 0
transform 1 0 4090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3757_
timestamp 0
transform 1 0 4570 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3758_
timestamp 0
transform -1 0 5090 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__3759_
timestamp 0
transform -1 0 4870 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__3760_
timestamp 0
transform -1 0 4310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3761_
timestamp 0
transform -1 0 4330 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__3762_
timestamp 0
transform -1 0 4430 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__3763_
timestamp 0
transform -1 0 4170 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3764_
timestamp 0
transform -1 0 3450 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3765_
timestamp 0
transform -1 0 4630 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__3766_
timestamp 0
transform 1 0 2250 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3767_
timestamp 0
transform -1 0 2470 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3768_
timestamp 0
transform -1 0 2630 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3769_
timestamp 0
transform -1 0 2830 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3770_
timestamp 0
transform -1 0 3830 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3771_
timestamp 0
transform 1 0 3410 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3772_
timestamp 0
transform -1 0 1050 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3773_
timestamp 0
transform 1 0 5830 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__3774_
timestamp 0
transform 1 0 5050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__3775_
timestamp 0
transform -1 0 5010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3776_
timestamp 0
transform -1 0 4850 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3777_
timestamp 0
transform 1 0 4910 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3778_
timestamp 0
transform 1 0 4750 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3779_
timestamp 0
transform 1 0 4550 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3780_
timestamp 0
transform 1 0 5230 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3781_
timestamp 0
transform -1 0 5410 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3782_
timestamp 0
transform -1 0 4390 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3783_
timestamp 0
transform 1 0 3830 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3784_
timestamp 0
transform -1 0 5270 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3785_
timestamp 0
transform 1 0 7550 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__3786_
timestamp 0
transform 1 0 7410 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__3787_
timestamp 0
transform -1 0 7390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3788_
timestamp 0
transform -1 0 7230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3789_
timestamp 0
transform -1 0 7250 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3790_
timestamp 0
transform -1 0 6230 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3791_
timestamp 0
transform -1 0 6610 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3792_
timestamp 0
transform 1 0 7030 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3793_
timestamp 0
transform -1 0 6830 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3794_
timestamp 0
transform 1 0 7990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__3795_
timestamp 0
transform -1 0 9610 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3796_
timestamp 0
transform 1 0 8310 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3797_
timestamp 0
transform 1 0 7690 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3798_
timestamp 0
transform 1 0 6970 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3799_
timestamp 0
transform -1 0 7150 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3800_
timestamp 0
transform -1 0 7330 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3801_
timestamp 0
transform 1 0 5670 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3802_
timestamp 0
transform -1 0 5930 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3803_
timestamp 0
transform 1 0 5710 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3804_
timestamp 0
transform 1 0 5330 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3805_
timestamp 0
transform 1 0 5370 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3806_
timestamp 0
transform 1 0 5050 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3807_
timestamp 0
transform -1 0 5530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3808_
timestamp 0
transform -1 0 7910 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3809_
timestamp 0
transform -1 0 8030 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3810_
timestamp 0
transform 1 0 7830 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3811_
timestamp 0
transform -1 0 7510 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3812_
timestamp 0
transform 1 0 10450 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3813_
timestamp 0
transform -1 0 9870 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3814_
timestamp 0
transform 1 0 9850 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3815_
timestamp 0
transform -1 0 9850 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3816_
timestamp 0
transform -1 0 9690 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3817_
timestamp 0
transform 1 0 9150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3818_
timestamp 0
transform -1 0 8970 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3819_
timestamp 0
transform 1 0 10150 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3820_
timestamp 0
transform 1 0 10230 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3821_
timestamp 0
transform 1 0 6550 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3822_
timestamp 0
transform -1 0 3350 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3823_
timestamp 0
transform -1 0 8270 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3824_
timestamp 0
transform 1 0 7290 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3825_
timestamp 0
transform -1 0 9990 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3826_
timestamp 0
transform 1 0 9470 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3827_
timestamp 0
transform -1 0 9310 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3828_
timestamp 0
transform 1 0 9110 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3829_
timestamp 0
transform 1 0 8910 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3830_
timestamp 0
transform 1 0 7410 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3831_
timestamp 0
transform 1 0 7690 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3832_
timestamp 0
transform 1 0 8550 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3833_
timestamp 0
transform 1 0 8730 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3834_
timestamp 0
transform -1 0 8710 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3835_
timestamp 0
transform 1 0 8910 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3836_
timestamp 0
transform 1 0 9210 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3837_
timestamp 0
transform -1 0 8470 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3838_
timestamp 0
transform 1 0 8650 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3839_
timestamp 0
transform 1 0 8890 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3840_
timestamp 0
transform -1 0 8530 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3841_
timestamp 0
transform -1 0 8330 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3842_
timestamp 0
transform 1 0 9090 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3843_
timestamp 0
transform -1 0 8350 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3844_
timestamp 0
transform 1 0 7650 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3845_
timestamp 0
transform 1 0 9310 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__3846_
timestamp 0
transform 1 0 8870 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3847_
timestamp 0
transform 1 0 8150 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3848_
timestamp 0
transform -1 0 8010 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__3849_
timestamp 0
transform 1 0 7790 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__3850_
timestamp 0
transform 1 0 7970 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3851_
timestamp 0
transform 1 0 7630 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3852_
timestamp 0
transform -1 0 7830 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3853_
timestamp 0
transform -1 0 7590 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3854_
timestamp 0
transform -1 0 7450 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3855_
timestamp 0
transform 1 0 7830 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__3856_
timestamp 0
transform -1 0 7230 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3857_
timestamp 0
transform -1 0 8330 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3858_
timestamp 0
transform 1 0 8670 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3859_
timestamp 0
transform 1 0 7850 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3860_
timestamp 0
transform 1 0 4790 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3861_
timestamp 0
transform 1 0 8530 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3862_
timestamp 0
transform -1 0 8770 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3863_
timestamp 0
transform -1 0 10230 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3864_
timestamp 0
transform 1 0 9470 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3865_
timestamp 0
transform 1 0 8050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3866_
timestamp 0
transform 1 0 5650 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3867_
timestamp 0
transform -1 0 7490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3868_
timestamp 0
transform -1 0 8550 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3869_
timestamp 0
transform 1 0 7970 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3870_
timestamp 0
transform -1 0 7850 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3871_
timestamp 0
transform 1 0 6390 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3872_
timestamp 0
transform 1 0 5690 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3873_
timestamp 0
transform -1 0 9530 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3874_
timestamp 0
transform 1 0 9870 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__3875_
timestamp 0
transform 1 0 6910 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3876_
timestamp 0
transform 1 0 5010 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3877_
timestamp 0
transform -1 0 4650 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3878_
timestamp 0
transform 1 0 4810 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3879_
timestamp 0
transform 1 0 4570 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3880_
timestamp 0
transform 1 0 5130 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3881_
timestamp 0
transform -1 0 5350 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3882_
timestamp 0
transform -1 0 4370 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3883_
timestamp 0
transform -1 0 4990 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3884_
timestamp 0
transform -1 0 4810 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3885_
timestamp 0
transform 1 0 5170 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3886_
timestamp 0
transform 1 0 9670 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__3887_
timestamp 0
transform 1 0 10390 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__3888_
timestamp 0
transform 1 0 10350 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__3889_
timestamp 0
transform -1 0 10850 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__3890_
timestamp 0
transform -1 0 10770 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3891_
timestamp 0
transform 1 0 10930 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3892_
timestamp 0
transform -1 0 8790 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__3893_
timestamp 0
transform -1 0 8590 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__3894_
timestamp 0
transform -1 0 11290 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3895_
timestamp 0
transform 1 0 11070 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3896_
timestamp 0
transform 1 0 11830 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3897_
timestamp 0
transform 1 0 11090 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__3898_
timestamp 0
transform 1 0 8270 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3899_
timestamp 0
transform -1 0 5630 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3900_
timestamp 0
transform 1 0 4090 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3901_
timestamp 0
transform -1 0 5050 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__3902_
timestamp 0
transform 1 0 4970 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3903_
timestamp 0
transform 1 0 7450 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3904_
timestamp 0
transform -1 0 7030 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3905_
timestamp 0
transform -1 0 6470 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3906_
timestamp 0
transform 1 0 5050 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3907_
timestamp 0
transform -1 0 8210 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__3908_
timestamp 0
transform -1 0 6810 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3909_
timestamp 0
transform -1 0 5990 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__3910_
timestamp 0
transform 1 0 5870 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__3911_
timestamp 0
transform -1 0 4550 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3912_
timestamp 0
transform 1 0 4350 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__3913_
timestamp 0
transform -1 0 4570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3914_
timestamp 0
transform 1 0 4230 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__3915_
timestamp 0
transform 1 0 4770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3916_
timestamp 0
transform 1 0 4970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3917_
timestamp 0
transform 1 0 5350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3918_
timestamp 0
transform -1 0 4670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3919_
timestamp 0
transform 1 0 4770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__3920_
timestamp 0
transform 1 0 4490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3921_
timestamp 0
transform 1 0 810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3922_
timestamp 0
transform 1 0 910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3923_
timestamp 0
transform 1 0 430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3924_
timestamp 0
transform 1 0 790 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__3925_
timestamp 0
transform 1 0 5090 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3926_
timestamp 0
transform 1 0 5290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3927_
timestamp 0
transform -1 0 4710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3928_
timestamp 0
transform 1 0 5470 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3929_
timestamp 0
transform -1 0 4590 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__3930_
timestamp 0
transform 1 0 3430 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__3931_
timestamp 0
transform 1 0 3470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__3932_
timestamp 0
transform 1 0 2330 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__3933_
timestamp 0
transform 1 0 3230 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__3934_
timestamp 0
transform -1 0 4470 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__3935_
timestamp 0
transform 1 0 3830 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3936_
timestamp 0
transform 1 0 3630 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__3937_
timestamp 0
transform 1 0 4210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__3938_
timestamp 0
transform -1 0 3490 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__3939_
timestamp 0
transform 1 0 3590 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__3940_
timestamp 0
transform -1 0 4730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__3941_
timestamp 0
transform 1 0 6930 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3942_
timestamp 0
transform -1 0 10010 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3943_
timestamp 0
transform -1 0 9990 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__3944_
timestamp 0
transform -1 0 9690 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__3945_
timestamp 0
transform -1 0 10210 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3946_
timestamp 0
transform 1 0 9790 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__3947_
timestamp 0
transform 1 0 10390 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3948_
timestamp 0
transform 1 0 10570 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3949_
timestamp 0
transform 1 0 7690 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__3950_
timestamp 0
transform -1 0 6970 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3951_
timestamp 0
transform 1 0 6570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3952_
timestamp 0
transform -1 0 5790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__3953_
timestamp 0
transform 1 0 5450 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3954_
timestamp 0
transform -1 0 5850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3955_
timestamp 0
transform 1 0 5910 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3956_
timestamp 0
transform -1 0 6130 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3957_
timestamp 0
transform 1 0 6150 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3958_
timestamp 0
transform 1 0 6350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3959_
timestamp 0
transform 1 0 6470 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3960_
timestamp 0
transform 1 0 2390 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3961_
timestamp 0
transform -1 0 2790 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3962_
timestamp 0
transform 1 0 2930 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3963_
timestamp 0
transform 1 0 3530 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3964_
timestamp 0
transform -1 0 4110 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3965_
timestamp 0
transform -1 0 3350 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3966_
timestamp 0
transform -1 0 4310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3967_
timestamp 0
transform -1 0 5110 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3968_
timestamp 0
transform -1 0 5310 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3969_
timestamp 0
transform -1 0 4310 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3970_
timestamp 0
transform 1 0 3930 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3971_
timestamp 0
transform 1 0 5630 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__3972_
timestamp 0
transform 1 0 5450 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__3973_
timestamp 0
transform 1 0 5450 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3974_
timestamp 0
transform -1 0 5670 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3975_
timestamp 0
transform -1 0 5670 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3976_
timestamp 0
transform -1 0 5670 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3977_
timestamp 0
transform 1 0 5550 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__3978_
timestamp 0
transform 1 0 6370 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3979_
timestamp 0
transform -1 0 2730 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3980_
timestamp 0
transform 1 0 2030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__3981_
timestamp 0
transform 1 0 1870 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__3982_
timestamp 0
transform 1 0 1810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__3983_
timestamp 0
transform -1 0 1950 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__3984_
timestamp 0
transform 1 0 8270 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__3985_
timestamp 0
transform 1 0 6850 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3986_
timestamp 0
transform -1 0 7350 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__3987_
timestamp 0
transform 1 0 7630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3988_
timestamp 0
transform 1 0 7550 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3989_
timestamp 0
transform 1 0 7350 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3990_
timestamp 0
transform 1 0 7150 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3991_
timestamp 0
transform -1 0 7310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__3992_
timestamp 0
transform -1 0 7970 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3993_
timestamp 0
transform 1 0 7730 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3994_
timestamp 0
transform -1 0 7070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__3995_
timestamp 0
transform -1 0 9430 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3996_
timestamp 0
transform -1 0 6030 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__3997_
timestamp 0
transform 1 0 5990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__3998_
timestamp 0
transform -1 0 6070 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__3999_
timestamp 0
transform 1 0 5850 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4000_
timestamp 0
transform -1 0 5270 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4001_
timestamp 0
transform -1 0 5110 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4002_
timestamp 0
transform -1 0 6970 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4003_
timestamp 0
transform -1 0 6610 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4004_
timestamp 0
transform 1 0 2650 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4005_
timestamp 0
transform 1 0 2850 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4006_
timestamp 0
transform -1 0 2670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4007_
timestamp 0
transform 1 0 2450 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4008_
timestamp 0
transform -1 0 7130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4009_
timestamp 0
transform 1 0 6910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4010_
timestamp 0
transform -1 0 6770 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4011_
timestamp 0
transform 1 0 8650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4012_
timestamp 0
transform 1 0 6750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4013_
timestamp 0
transform 1 0 6630 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4014_
timestamp 0
transform 1 0 6170 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4015_
timestamp 0
transform 1 0 6530 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4016_
timestamp 0
transform 1 0 9350 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4017_
timestamp 0
transform -1 0 9670 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4018_
timestamp 0
transform -1 0 9850 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4019_
timestamp 0
transform 1 0 10010 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4020_
timestamp 0
transform -1 0 7490 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4021_
timestamp 0
transform -1 0 10050 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4022_
timestamp 0
transform -1 0 6830 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4023_
timestamp 0
transform -1 0 7170 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4024_
timestamp 0
transform 1 0 8970 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4025_
timestamp 0
transform -1 0 7690 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4026_
timestamp 0
transform -1 0 7850 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4027_
timestamp 0
transform 1 0 8390 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4028_
timestamp 0
transform 1 0 7930 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4029_
timestamp 0
transform 1 0 11030 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4030_
timestamp 0
transform 1 0 10850 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4031_
timestamp 0
transform 1 0 9230 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4032_
timestamp 0
transform 1 0 8670 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4033_
timestamp 0
transform -1 0 9330 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4034_
timestamp 0
transform 1 0 3990 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4035_
timestamp 0
transform 1 0 9790 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4036_
timestamp 0
transform -1 0 9650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4037_
timestamp 0
transform -1 0 9170 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4038_
timestamp 0
transform -1 0 8130 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4039_
timestamp 0
transform -1 0 7070 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4040_
timestamp 0
transform 1 0 12010 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4041_
timestamp 0
transform 1 0 9290 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4042_
timestamp 0
transform -1 0 6010 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__4043_
timestamp 0
transform 1 0 5330 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4044_
timestamp 0
transform -1 0 5410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4045_
timestamp 0
transform -1 0 5470 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4046_
timestamp 0
transform -1 0 5830 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4047_
timestamp 0
transform -1 0 6010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4048_
timestamp 0
transform -1 0 6010 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4049_
timestamp 0
transform 1 0 5490 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4050_
timestamp 0
transform -1 0 5270 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4051_
timestamp 0
transform 1 0 5610 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4052_
timestamp 0
transform -1 0 6230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4053_
timestamp 0
transform -1 0 8210 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4054_
timestamp 0
transform 1 0 3730 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4055_
timestamp 0
transform -1 0 3570 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4056_
timestamp 0
transform 1 0 2730 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4057_
timestamp 0
transform 1 0 3350 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4058_
timestamp 0
transform -1 0 7490 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4059_
timestamp 0
transform 1 0 7350 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4060_
timestamp 0
transform -1 0 8030 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4061_
timestamp 0
transform -1 0 8970 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4062_
timestamp 0
transform -1 0 3150 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4063_
timestamp 0
transform 1 0 5070 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4064_
timestamp 0
transform -1 0 5050 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4065_
timestamp 0
transform 1 0 5270 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4066_
timestamp 0
transform 1 0 4470 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4067_
timestamp 0
transform -1 0 7110 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4068_
timestamp 0
transform 1 0 3130 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4069_
timestamp 0
transform -1 0 670 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__4070_
timestamp 0
transform 1 0 1150 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__4071_
timestamp 0
transform 1 0 550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__4072_
timestamp 0
transform -1 0 870 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__4073_
timestamp 0
transform 1 0 4090 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4074_
timestamp 0
transform 1 0 4290 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4075_
timestamp 0
transform 1 0 4210 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4076_
timestamp 0
transform -1 0 5470 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4077_
timestamp 0
transform 1 0 5490 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4078_
timestamp 0
transform -1 0 5510 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4079_
timestamp 0
transform 1 0 3770 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4080_
timestamp 0
transform 1 0 5870 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4081_
timestamp 0
transform 1 0 910 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4082_
timestamp 0
transform 1 0 4150 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4083_
timestamp 0
transform -1 0 3950 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4084_
timestamp 0
transform 1 0 1650 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4085_
timestamp 0
transform 1 0 1470 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4086_
timestamp 0
transform 1 0 1610 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4087_
timestamp 0
transform 1 0 1570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4088_
timestamp 0
transform -1 0 4510 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4089_
timestamp 0
transform -1 0 4470 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4090_
timestamp 0
transform -1 0 3970 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4091_
timestamp 0
transform -1 0 3410 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4092_
timestamp 0
transform -1 0 5690 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4093_
timestamp 0
transform 1 0 4630 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4094_
timestamp 0
transform 1 0 4210 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4095_
timestamp 0
transform 1 0 1950 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4096_
timestamp 0
transform 1 0 1770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4097_
timestamp 0
transform 1 0 1650 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4098_
timestamp 0
transform 1 0 1570 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4099_
timestamp 0
transform 1 0 7150 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4100_
timestamp 0
transform 1 0 8030 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4101_
timestamp 0
transform 1 0 8190 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4102_
timestamp 0
transform -1 0 8390 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4103_
timestamp 0
transform 1 0 8010 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4104_
timestamp 0
transform -1 0 8230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4105_
timestamp 0
transform 1 0 8670 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4106_
timestamp 0
transform 1 0 6710 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4107_
timestamp 0
transform -1 0 1110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3__4108_
timestamp 0
transform -1 0 510 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__4109_
timestamp 0
transform -1 0 1850 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4110_
timestamp 0
transform -1 0 7790 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4111_
timestamp 0
transform -1 0 9530 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4112_
timestamp 0
transform 1 0 2910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__4113_
timestamp 0
transform 1 0 3110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__4114_
timestamp 0
transform 1 0 3610 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4115_
timestamp 0
transform 1 0 4490 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4116_
timestamp 0
transform -1 0 5370 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4117_
timestamp 0
transform 1 0 4910 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4118_
timestamp 0
transform 1 0 4830 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4119_
timestamp 0
transform 1 0 3990 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4120_
timestamp 0
transform -1 0 3730 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4121_
timestamp 0
transform -1 0 4570 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4122_
timestamp 0
transform 1 0 4710 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4123_
timestamp 0
transform 1 0 8070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4124_
timestamp 0
transform 1 0 8590 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4125_
timestamp 0
transform -1 0 4310 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4126_
timestamp 0
transform 1 0 4270 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4127_
timestamp 0
transform 1 0 4090 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4128_
timestamp 0
transform 1 0 4510 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4129_
timestamp 0
transform -1 0 4930 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4130_
timestamp 0
transform 1 0 6050 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4131_
timestamp 0
transform 1 0 4330 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4132_
timestamp 0
transform -1 0 4550 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4133_
timestamp 0
transform -1 0 2030 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4134_
timestamp 0
transform 1 0 1810 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4135_
timestamp 0
transform -1 0 2170 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4136_
timestamp 0
transform -1 0 2170 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4137_
timestamp 0
transform -1 0 2010 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4138_
timestamp 0
transform -1 0 2250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4139_
timestamp 0
transform 1 0 2030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4140_
timestamp 0
transform -1 0 3050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4141_
timestamp 0
transform 1 0 1830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4142_
timestamp 0
transform 1 0 1630 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4143_
timestamp 0
transform -1 0 1470 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4144_
timestamp 0
transform 1 0 1610 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4145_
timestamp 0
transform -1 0 1090 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4146_
timestamp 0
transform 1 0 3110 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4147_
timestamp 0
transform -1 0 2050 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4148_
timestamp 0
transform -1 0 3230 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4149_
timestamp 0
transform 1 0 3210 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4150_
timestamp 0
transform 1 0 3210 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4151_
timestamp 0
transform 1 0 3750 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4152_
timestamp 0
transform -1 0 3690 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4153_
timestamp 0
transform -1 0 2070 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4154_
timestamp 0
transform -1 0 2270 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4155_
timestamp 0
transform 1 0 650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4156_
timestamp 0
transform 1 0 1010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4157_
timestamp 0
transform -1 0 5950 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4158_
timestamp 0
transform 1 0 6110 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4159_
timestamp 0
transform 1 0 6310 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4160_
timestamp 0
transform 1 0 5390 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4161_
timestamp 0
transform -1 0 5610 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4162_
timestamp 0
transform 1 0 5190 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4163_
timestamp 0
transform -1 0 5210 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4164_
timestamp 0
transform 1 0 5750 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4165_
timestamp 0
transform -1 0 5750 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4166_
timestamp 0
transform 1 0 5770 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4167_
timestamp 0
transform 1 0 6470 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4168_
timestamp 0
transform -1 0 5910 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4169_
timestamp 0
transform 1 0 5710 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4170_
timestamp 0
transform 1 0 6110 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4171_
timestamp 0
transform 1 0 5530 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4172_
timestamp 0
transform 1 0 5150 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4173_
timestamp 0
transform 1 0 3830 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4174_
timestamp 0
transform 1 0 5550 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4175_
timestamp 0
transform 1 0 5170 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4176_
timestamp 0
transform -1 0 3350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4177_
timestamp 0
transform 1 0 3030 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4178_
timestamp 0
transform -1 0 2250 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4179_
timestamp 0
transform -1 0 2370 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4180_
timestamp 0
transform 1 0 2830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4181_
timestamp 0
transform -1 0 2450 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4182_
timestamp 0
transform 1 0 2290 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4183_
timestamp 0
transform -1 0 3270 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4184_
timestamp 0
transform 1 0 3430 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4185_
timestamp 0
transform 1 0 2850 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4186_
timestamp 0
transform -1 0 2470 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4187_
timestamp 0
transform 1 0 4090 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4188_
timestamp 0
transform 1 0 4290 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4189_
timestamp 0
transform -1 0 4110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4190_
timestamp 0
transform -1 0 3930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4191_
timestamp 0
transform -1 0 3750 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4192_
timestamp 0
transform -1 0 5210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4193_
timestamp 0
transform -1 0 5070 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4194_
timestamp 0
transform -1 0 3930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4195_
timestamp 0
transform 1 0 3470 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4196_
timestamp 0
transform 1 0 3770 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4197_
timestamp 0
transform 1 0 1630 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4198_
timestamp 0
transform -1 0 1750 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4199_
timestamp 0
transform -1 0 1950 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4200_
timestamp 0
transform -1 0 2350 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4201_
timestamp 0
transform -1 0 1570 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4202_
timestamp 0
transform -1 0 1450 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__4203_
timestamp 0
transform -1 0 1830 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__4204_
timestamp 0
transform -1 0 2630 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4205_
timestamp 0
transform 1 0 2630 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4206_
timestamp 0
transform -1 0 8610 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4207_
timestamp 0
transform -1 0 7950 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4208_
timestamp 0
transform -1 0 6290 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4209_
timestamp 0
transform -1 0 290 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4210_
timestamp 0
transform 1 0 70 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4211_
timestamp 0
transform -1 0 90 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4212_
timestamp 0
transform -1 0 470 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4213_
timestamp 0
transform 1 0 930 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4214_
timestamp 0
transform -1 0 1450 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4215_
timestamp 0
transform 1 0 1430 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4216_
timestamp 0
transform -1 0 2030 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4217_
timestamp 0
transform -1 0 3010 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4218_
timestamp 0
transform -1 0 2230 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4219_
timestamp 0
transform 1 0 2310 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4220_
timestamp 0
transform 1 0 2510 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4221_
timestamp 0
transform -1 0 290 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4222_
timestamp 0
transform -1 0 90 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4223_
timestamp 0
transform -1 0 470 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4224_
timestamp 0
transform -1 0 470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4225_
timestamp 0
transform -1 0 450 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4226_
timestamp 0
transform 1 0 70 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4227_
timestamp 0
transform -1 0 290 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4228_
timestamp 0
transform -1 0 2430 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4229_
timestamp 0
transform 1 0 2630 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4230_
timestamp 0
transform -1 0 2850 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4231_
timestamp 0
transform 1 0 3190 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4232_
timestamp 0
transform -1 0 3650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4233_
timestamp 0
transform -1 0 2230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4234_
timestamp 0
transform -1 0 3090 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4235_
timestamp 0
transform -1 0 3850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4236_
timestamp 0
transform 1 0 3930 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4237_
timestamp 0
transform -1 0 4150 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4238_
timestamp 0
transform 1 0 3470 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4239_
timestamp 0
transform 1 0 2630 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4240_
timestamp 0
transform 1 0 2270 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4241_
timestamp 0
transform -1 0 2130 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4242_
timestamp 0
transform 1 0 2310 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4243_
timestamp 0
transform -1 0 4490 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4244_
timestamp 0
transform -1 0 5490 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4245_
timestamp 0
transform -1 0 6070 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4246_
timestamp 0
transform -1 0 4190 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4247_
timestamp 0
transform 1 0 2590 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4248_
timestamp 0
transform -1 0 5670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4249_
timestamp 0
transform -1 0 2370 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4250_
timestamp 0
transform -1 0 4290 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4251_
timestamp 0
transform 1 0 5670 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4252_
timestamp 0
transform -1 0 5870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4253_
timestamp 0
transform -1 0 3770 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4254_
timestamp 0
transform -1 0 2190 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4255_
timestamp 0
transform 1 0 2530 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4256_
timestamp 0
transform -1 0 3890 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4257_
timestamp 0
transform 1 0 4070 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4258_
timestamp 0
transform 1 0 4270 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4259_
timestamp 0
transform 1 0 4030 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4260_
timestamp 0
transform -1 0 2990 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4261_
timestamp 0
transform -1 0 4050 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4262_
timestamp 0
transform 1 0 1570 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4263_
timestamp 0
transform -1 0 7990 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4264_
timestamp 0
transform 1 0 7610 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4265_
timestamp 0
transform 1 0 7430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4266_
timestamp 0
transform 1 0 7110 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4267_
timestamp 0
transform 1 0 7550 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4268_
timestamp 0
transform -1 0 6790 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4269_
timestamp 0
transform -1 0 9470 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4270_
timestamp 0
transform -1 0 11170 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4271_
timestamp 0
transform 1 0 11150 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4272_
timestamp 0
transform 1 0 9250 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4273_
timestamp 0
transform 1 0 9050 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4274_
timestamp 0
transform -1 0 8970 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4275_
timestamp 0
transform 1 0 8790 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4276_
timestamp 0
transform 1 0 8870 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4277_
timestamp 0
transform 1 0 8890 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4278_
timestamp 0
transform 1 0 7770 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4279_
timestamp 0
transform 1 0 10550 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4280_
timestamp 0
transform 1 0 10750 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4281_
timestamp 0
transform -1 0 10710 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4282_
timestamp 0
transform -1 0 1250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4283_
timestamp 0
transform -1 0 7090 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4284_
timestamp 0
transform 1 0 7670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4285_
timestamp 0
transform 1 0 7410 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4286_
timestamp 0
transform -1 0 1090 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4287_
timestamp 0
transform -1 0 1290 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4288_
timestamp 0
transform -1 0 1690 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4289_
timestamp 0
transform -1 0 4390 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4290_
timestamp 0
transform 1 0 6870 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4291_
timestamp 0
transform 1 0 6890 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4292_
timestamp 0
transform -1 0 2550 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4293_
timestamp 0
transform -1 0 1830 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4294_
timestamp 0
transform -1 0 7310 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4295_
timestamp 0
transform 1 0 1510 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4296_
timestamp 0
transform -1 0 90 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4297_
timestamp 0
transform 1 0 1170 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4298_
timestamp 0
transform -1 0 3290 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4299_
timestamp 0
transform 1 0 3370 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4300_
timestamp 0
transform -1 0 3850 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4301_
timestamp 0
transform -1 0 3570 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4302_
timestamp 0
transform -1 0 3690 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4303_
timestamp 0
transform -1 0 1610 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4304_
timestamp 0
transform 1 0 1190 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4305_
timestamp 0
transform -1 0 2310 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4306_
timestamp 0
transform -1 0 2870 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4307_
timestamp 0
transform 1 0 6230 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4308_
timestamp 0
transform -1 0 6310 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4309_
timestamp 0
transform 1 0 2870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4310_
timestamp 0
transform -1 0 2450 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4311_
timestamp 0
transform 1 0 2350 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4312_
timestamp 0
transform 1 0 930 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4313_
timestamp 0
transform 1 0 1510 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4314_
timestamp 0
transform 1 0 1690 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4315_
timestamp 0
transform -1 0 2730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4316_
timestamp 0
transform -1 0 2790 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4317_
timestamp 0
transform 1 0 4430 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4318_
timestamp 0
transform 1 0 4110 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4319_
timestamp 0
transform 1 0 3610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4320_
timestamp 0
transform -1 0 3050 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4321_
timestamp 0
transform 1 0 2830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4322_
timestamp 0
transform 1 0 1570 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4323_
timestamp 0
transform -1 0 2690 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4324_
timestamp 0
transform -1 0 1830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4325_
timestamp 0
transform -1 0 4090 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4326_
timestamp 0
transform 1 0 3990 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4327_
timestamp 0
transform 1 0 4130 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4328_
timestamp 0
transform -1 0 8570 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4329_
timestamp 0
transform 1 0 1730 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4330_
timestamp 0
transform 1 0 2130 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4331_
timestamp 0
transform -1 0 1450 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4332_
timestamp 0
transform -1 0 1990 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4333_
timestamp 0
transform -1 0 2910 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4334_
timestamp 0
transform -1 0 3110 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4335_
timestamp 0
transform -1 0 3690 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4336_
timestamp 0
transform 1 0 2850 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4337_
timestamp 0
transform 1 0 2650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4338_
timestamp 0
transform 1 0 2690 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4339_
timestamp 0
transform -1 0 3310 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4340_
timestamp 0
transform -1 0 3490 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4341_
timestamp 0
transform 1 0 3430 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4342_
timestamp 0
transform -1 0 3250 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4343_
timestamp 0
transform 1 0 3490 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4344_
timestamp 0
transform 1 0 1790 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4345_
timestamp 0
transform -1 0 2430 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4346_
timestamp 0
transform 1 0 6910 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4347_
timestamp 0
transform -1 0 6730 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4348_
timestamp 0
transform -1 0 630 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4349_
timestamp 0
transform -1 0 1050 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4350_
timestamp 0
transform 1 0 2170 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4351_
timestamp 0
transform -1 0 2790 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4352_
timestamp 0
transform 1 0 3770 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4353_
timestamp 0
transform -1 0 6170 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4354_
timestamp 0
transform -1 0 3450 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4355_
timestamp 0
transform -1 0 870 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4356_
timestamp 0
transform -1 0 510 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4357_
timestamp 0
transform 1 0 2370 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4358_
timestamp 0
transform -1 0 5230 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4359_
timestamp 0
transform 1 0 5150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4360_
timestamp 0
transform -1 0 5110 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4361_
timestamp 0
transform 1 0 3050 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4362_
timestamp 0
transform 1 0 4890 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4363_
timestamp 0
transform -1 0 4730 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4364_
timestamp 0
transform 1 0 3690 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4365_
timestamp 0
transform -1 0 5670 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4366_
timestamp 0
transform -1 0 5870 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4367_
timestamp 0
transform -1 0 2910 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4368_
timestamp 0
transform 1 0 7550 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4369_
timestamp 0
transform -1 0 7390 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4370_
timestamp 0
transform 1 0 670 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4371_
timestamp 0
transform -1 0 1810 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4372_
timestamp 0
transform 1 0 1930 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4373_
timestamp 0
transform 1 0 2130 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4374_
timestamp 0
transform 1 0 2490 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4375_
timestamp 0
transform -1 0 3810 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4376_
timestamp 0
transform 1 0 7490 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4377_
timestamp 0
transform 1 0 11550 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4378_
timestamp 0
transform -1 0 1270 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4379_
timestamp 0
transform -1 0 5230 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4380_
timestamp 0
transform 1 0 4810 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4381_
timestamp 0
transform 1 0 5910 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4382_
timestamp 0
transform 1 0 250 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4383_
timestamp 0
transform 1 0 70 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4384_
timestamp 0
transform 1 0 6250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4385_
timestamp 0
transform 1 0 6450 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4386_
timestamp 0
transform 1 0 6850 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4387_
timestamp 0
transform 1 0 6650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4388_
timestamp 0
transform -1 0 5450 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4389_
timestamp 0
transform -1 0 6550 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4390_
timestamp 0
transform 1 0 7050 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4391_
timestamp 0
transform 1 0 5010 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4392_
timestamp 0
transform -1 0 6350 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4393_
timestamp 0
transform 1 0 6510 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4394_
timestamp 0
transform 1 0 6690 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4395_
timestamp 0
transform 1 0 6810 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4396_
timestamp 0
transform -1 0 6290 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4397_
timestamp 0
transform 1 0 4050 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4398_
timestamp 0
transform 1 0 3030 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4399_
timestamp 0
transform 1 0 2150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4400_
timestamp 0
transform -1 0 6330 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4401_
timestamp 0
transform 1 0 6250 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4402_
timestamp 0
transform -1 0 6090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4403_
timestamp 0
transform -1 0 5630 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4404_
timestamp 0
transform 1 0 1410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4405_
timestamp 0
transform -1 0 1850 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4406_
timestamp 0
transform -1 0 2550 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4407_
timestamp 0
transform -1 0 2350 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4408_
timestamp 0
transform 1 0 1570 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4409_
timestamp 0
transform -1 0 1790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4410_
timestamp 0
transform 1 0 3590 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4411_
timestamp 0
transform 1 0 3910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4412_
timestamp 0
transform 1 0 1750 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4413_
timestamp 0
transform -1 0 270 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4414_
timestamp 0
transform 1 0 270 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4415_
timestamp 0
transform 1 0 450 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4416_
timestamp 0
transform 1 0 1530 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__4417_
timestamp 0
transform -1 0 1750 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__4418_
timestamp 0
transform -1 0 2570 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__4419_
timestamp 0
transform 1 0 2130 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__4420_
timestamp 0
transform 1 0 2250 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4421_
timestamp 0
transform 1 0 2450 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4422_
timestamp 0
transform -1 0 1990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4423_
timestamp 0
transform -1 0 630 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4424_
timestamp 0
transform 1 0 2050 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4425_
timestamp 0
transform 1 0 1090 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4426_
timestamp 0
transform 1 0 1290 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4427_
timestamp 0
transform 1 0 3550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4428_
timestamp 0
transform -1 0 3390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4429_
timestamp 0
transform 1 0 1270 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4430_
timestamp 0
transform 1 0 1470 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4431_
timestamp 0
transform -1 0 750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4432_
timestamp 0
transform -1 0 630 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4433_
timestamp 0
transform -1 0 870 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4434_
timestamp 0
transform -1 0 1330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__4435_
timestamp 0
transform 1 0 1510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__4436_
timestamp 0
transform 1 0 3110 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__4437_
timestamp 0
transform -1 0 3330 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__4438_
timestamp 0
transform -1 0 6570 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4439_
timestamp 0
transform 1 0 5970 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4440_
timestamp 0
transform -1 0 4750 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4441_
timestamp 0
transform 1 0 4150 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4442_
timestamp 0
transform 1 0 3930 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4443_
timestamp 0
transform 1 0 3810 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4444_
timestamp 0
transform 1 0 3630 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4445_
timestamp 0
transform 1 0 3970 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4446_
timestamp 0
transform 1 0 4390 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4447_
timestamp 0
transform 1 0 4570 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4448_
timestamp 0
transform 1 0 2490 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4449_
timestamp 0
transform 1 0 1050 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4450_
timestamp 0
transform -1 0 1810 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4451_
timestamp 0
transform 1 0 1410 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4452_
timestamp 0
transform -1 0 2210 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4453_
timestamp 0
transform 1 0 7230 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4454_
timestamp 0
transform -1 0 1050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4455_
timestamp 0
transform 1 0 6770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4456_
timestamp 0
transform 1 0 6990 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4457_
timestamp 0
transform 1 0 7190 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4458_
timestamp 0
transform -1 0 7390 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4459_
timestamp 0
transform -1 0 7010 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4460_
timestamp 0
transform -1 0 8330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4461_
timestamp 0
transform 1 0 7610 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4462_
timestamp 0
transform -1 0 6710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4463_
timestamp 0
transform 1 0 1230 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4464_
timestamp 0
transform -1 0 2530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4465_
timestamp 0
transform -1 0 5870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4466_
timestamp 0
transform 1 0 6010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4467_
timestamp 0
transform 1 0 6430 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4468_
timestamp 0
transform 1 0 6670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4469_
timestamp 0
transform 1 0 6870 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4470_
timestamp 0
transform -1 0 6630 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4471_
timestamp 0
transform 1 0 7230 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4472_
timestamp 0
transform -1 0 6430 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4473_
timestamp 0
transform 1 0 8150 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4474_
timestamp 0
transform -1 0 6250 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4475_
timestamp 0
transform 1 0 2710 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4476_
timestamp 0
transform -1 0 1210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4477_
timestamp 0
transform -1 0 2610 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4478_
timestamp 0
transform 1 0 2590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4479_
timestamp 0
transform 1 0 5310 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4480_
timestamp 0
transform 1 0 1390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4481_
timestamp 0
transform 1 0 230 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4482_
timestamp 0
transform 1 0 430 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4483_
timestamp 0
transform 1 0 3190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4484_
timestamp 0
transform -1 0 4950 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4485_
timestamp 0
transform 1 0 5330 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4486_
timestamp 0
transform -1 0 5150 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4487_
timestamp 0
transform -1 0 5530 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4488_
timestamp 0
transform 1 0 5690 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4489_
timestamp 0
transform -1 0 5810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4490_
timestamp 0
transform -1 0 5770 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4491_
timestamp 0
transform -1 0 5850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4492_
timestamp 0
transform 1 0 70 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4493_
timestamp 0
transform -1 0 5690 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4494_
timestamp 0
transform 1 0 5490 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4495_
timestamp 0
transform 1 0 4350 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4496_
timestamp 0
transform 1 0 3810 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4497_
timestamp 0
transform -1 0 3590 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4498_
timestamp 0
transform -1 0 4630 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4499_
timestamp 0
transform 1 0 1250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4500_
timestamp 0
transform 1 0 6350 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4501_
timestamp 0
transform 1 0 6070 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4502_
timestamp 0
transform -1 0 4510 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4503_
timestamp 0
transform 1 0 6470 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4504_
timestamp 0
transform -1 0 1710 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__4505_
timestamp 0
transform -1 0 4830 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__4506_
timestamp 0
transform -1 0 5270 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4507_
timestamp 0
transform 1 0 5650 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__4508_
timestamp 0
transform 1 0 5530 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4509_
timestamp 0
transform -1 0 5750 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4510_
timestamp 0
transform -1 0 5930 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4511_
timestamp 0
transform 1 0 6090 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4512_
timestamp 0
transform 1 0 6190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4513_
timestamp 0
transform 1 0 6210 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4514_
timestamp 0
transform -1 0 1710 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__4515_
timestamp 0
transform -1 0 2550 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__4516_
timestamp 0
transform -1 0 4670 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__4517_
timestamp 0
transform -1 0 5150 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4518_
timestamp 0
transform 1 0 5110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4519_
timestamp 0
transform 1 0 5470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4520_
timestamp 0
transform -1 0 5670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4521_
timestamp 0
transform 1 0 6510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4522_
timestamp 0
transform -1 0 8930 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4523_
timestamp 0
transform 1 0 5310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4524_
timestamp 0
transform 1 0 6010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4525_
timestamp 0
transform 1 0 5870 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4526_
timestamp 0
transform -1 0 6450 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4527_
timestamp 0
transform -1 0 4950 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4528_
timestamp 0
transform 1 0 6350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4529_
timestamp 0
transform 1 0 6050 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4530_
timestamp 0
transform 1 0 6030 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4531_
timestamp 0
transform -1 0 2270 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__4532_
timestamp 0
transform -1 0 6290 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4533_
timestamp 0
transform -1 0 6230 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4534_
timestamp 0
transform 1 0 4270 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4535_
timestamp 0
transform 1 0 3670 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4536_
timestamp 0
transform -1 0 1090 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4537_
timestamp 0
transform 1 0 4450 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4538_
timestamp 0
transform -1 0 7690 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4539_
timestamp 0
transform -1 0 3070 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4540_
timestamp 0
transform 1 0 7650 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4541_
timestamp 0
transform 1 0 6510 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4542_
timestamp 0
transform 1 0 3050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4543_
timestamp 0
transform -1 0 2890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4544_
timestamp 0
transform -1 0 910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4545_
timestamp 0
transform 1 0 2130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4546_
timestamp 0
transform 1 0 2910 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4547_
timestamp 0
transform -1 0 2370 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4548_
timestamp 0
transform -1 0 1750 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4549_
timestamp 0
transform 1 0 2610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4550_
timestamp 0
transform 1 0 2810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4551_
timestamp 0
transform -1 0 3010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4552_
timestamp 0
transform -1 0 2990 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4553_
timestamp 0
transform -1 0 6550 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4554_
timestamp 0
transform 1 0 990 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4555_
timestamp 0
transform -1 0 750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__4556_
timestamp 0
transform 1 0 4350 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4557_
timestamp 0
transform 1 0 4170 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4558_
timestamp 0
transform -1 0 4010 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4559_
timestamp 0
transform 1 0 5030 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4560_
timestamp 0
transform -1 0 8490 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4561_
timestamp 0
transform -1 0 8890 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4562_
timestamp 0
transform 1 0 8410 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4563_
timestamp 0
transform -1 0 6390 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4564_
timestamp 0
transform -1 0 1890 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4565_
timestamp 0
transform 1 0 2710 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4566_
timestamp 0
transform 1 0 3090 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4567_
timestamp 0
transform -1 0 6790 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4568_
timestamp 0
transform 1 0 6710 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4569_
timestamp 0
transform 1 0 1930 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4570_
timestamp 0
transform -1 0 6590 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4571_
timestamp 0
transform 1 0 6290 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4572_
timestamp 0
transform -1 0 9530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4573_
timestamp 0
transform -1 0 10390 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4574_
timestamp 0
transform -1 0 9570 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4575_
timestamp 0
transform -1 0 6990 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4576_
timestamp 0
transform -1 0 8510 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4577_
timestamp 0
transform -1 0 3030 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4578_
timestamp 0
transform -1 0 5990 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4579_
timestamp 0
transform 1 0 8010 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4580_
timestamp 0
transform 1 0 10190 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4581_
timestamp 0
transform -1 0 7530 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4582_
timestamp 0
transform 1 0 1290 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4583_
timestamp 0
transform -1 0 2370 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4584_
timestamp 0
transform -1 0 2210 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4585_
timestamp 0
transform -1 0 2110 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4586_
timestamp 0
transform -1 0 1930 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4587_
timestamp 0
transform -1 0 1590 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4588_
timestamp 0
transform 1 0 3310 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4589_
timestamp 0
transform 1 0 3850 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4590_
timestamp 0
transform 1 0 1230 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4591_
timestamp 0
transform -1 0 1650 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4592_
timestamp 0
transform 1 0 1450 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4593_
timestamp 0
transform -1 0 4010 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4594_
timestamp 0
transform -1 0 3170 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__4595_
timestamp 0
transform -1 0 2730 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4596_
timestamp 0
transform -1 0 2930 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4597_
timestamp 0
transform 1 0 2790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__4598_
timestamp 0
transform -1 0 2710 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4599_
timestamp 0
transform -1 0 2890 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4600_
timestamp 0
transform -1 0 4050 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4601_
timestamp 0
transform -1 0 4010 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4602_
timestamp 0
transform -1 0 1430 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4603_
timestamp 0
transform -1 0 1370 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4604_
timestamp 0
transform -1 0 2970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__4605_
timestamp 0
transform 1 0 1790 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4606_
timestamp 0
transform -1 0 690 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4607_
timestamp 0
transform -1 0 510 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4608_
timestamp 0
transform -1 0 3250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4609_
timestamp 0
transform 1 0 1630 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__4610_
timestamp 0
transform 1 0 2510 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4611_
timestamp 0
transform -1 0 2350 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4612_
timestamp 0
transform -1 0 2010 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4613_
timestamp 0
transform 1 0 1990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__4614_
timestamp 0
transform -1 0 650 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4615_
timestamp 0
transform -1 0 470 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4616_
timestamp 0
transform -1 0 1830 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__4617_
timestamp 0
transform -1 0 1630 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__4618_
timestamp 0
transform -1 0 2530 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4619_
timestamp 0
transform -1 0 1870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4620_
timestamp 0
transform -1 0 1470 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4621_
timestamp 0
transform 1 0 2130 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4622_
timestamp 0
transform 1 0 2550 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4623_
timestamp 0
transform 1 0 2050 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4624_
timestamp 0
transform 1 0 1250 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4625_
timestamp 0
transform 1 0 870 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4626_
timestamp 0
transform -1 0 710 0 1 11290
box -6 -8 26 248
use FILL  FILL_3__4627_
timestamp 0
transform -1 0 2210 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__4628_
timestamp 0
transform -1 0 1270 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__4629_
timestamp 0
transform 1 0 1050 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3__4630_
timestamp 0
transform 1 0 1010 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4631_
timestamp 0
transform 1 0 1590 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4632_
timestamp 0
transform -1 0 750 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4633_
timestamp 0
transform -1 0 570 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4634_
timestamp 0
transform -1 0 7590 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4635_
timestamp 0
transform -1 0 1530 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4636_
timestamp 0
transform 1 0 1330 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4637_
timestamp 0
transform -1 0 1730 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4638_
timestamp 0
transform -1 0 890 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3__4639_
timestamp 0
transform 1 0 1090 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4640_
timestamp 0
transform 1 0 950 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4641_
timestamp 0
transform -1 0 1110 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4642_
timestamp 0
transform -1 0 2930 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__4643_
timestamp 0
transform 1 0 3070 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3__4644_
timestamp 0
transform -1 0 3510 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__4645_
timestamp 0
transform -1 0 870 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4646_
timestamp 0
transform 1 0 650 0 1 10810
box -6 -8 26 248
use FILL  FILL_3__4647_
timestamp 0
transform -1 0 1270 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4648_
timestamp 0
transform -1 0 1210 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4649_
timestamp 0
transform -1 0 570 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4650_
timestamp 0
transform -1 0 810 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3__4651_
timestamp 0
transform 1 0 4110 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__4652_
timestamp 0
transform 1 0 3830 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__4653_
timestamp 0
transform -1 0 4330 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__4654_
timestamp 0
transform -1 0 6890 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4655_
timestamp 0
transform 1 0 2550 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4656_
timestamp 0
transform -1 0 2370 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4657_
timestamp 0
transform -1 0 2290 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4658_
timestamp 0
transform 1 0 3730 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4659_
timestamp 0
transform -1 0 3950 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4660_
timestamp 0
transform -1 0 4330 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4661_
timestamp 0
transform 1 0 4510 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4662_
timestamp 0
transform 1 0 3970 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4663_
timestamp 0
transform 1 0 3410 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4664_
timestamp 0
transform 1 0 2550 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4665_
timestamp 0
transform -1 0 7830 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4666_
timestamp 0
transform 1 0 7730 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__4667_
timestamp 0
transform 1 0 6250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__4668_
timestamp 0
transform -1 0 6470 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3__4669_
timestamp 0
transform 1 0 450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4670_
timestamp 0
transform 1 0 4030 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4671_
timestamp 0
transform 1 0 3850 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4672_
timestamp 0
transform 1 0 2790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4673_
timestamp 0
transform -1 0 2990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4674_
timestamp 0
transform -1 0 3150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4675_
timestamp 0
transform -1 0 3030 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4676_
timestamp 0
transform -1 0 3630 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4677_
timestamp 0
transform -1 0 3570 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4678_
timestamp 0
transform 1 0 3390 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4679_
timestamp 0
transform -1 0 3230 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4680_
timestamp 0
transform -1 0 2230 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__4681_
timestamp 0
transform 1 0 2010 0 1 2650
box -6 -8 26 248
use FILL  FILL_3__4682_
timestamp 0
transform -1 0 7070 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4683_
timestamp 0
transform -1 0 1870 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4684_
timestamp 0
transform 1 0 3770 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4685_
timestamp 0
transform 1 0 3590 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4686_
timestamp 0
transform 1 0 11130 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4687_
timestamp 0
transform 1 0 11310 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4688_
timestamp 0
transform 1 0 11490 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4689_
timestamp 0
transform 1 0 11670 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4690_
timestamp 0
transform 1 0 10510 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4691_
timestamp 0
transform 1 0 10150 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4692_
timestamp 0
transform 1 0 10230 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4693_
timestamp 0
transform -1 0 9750 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4694_
timestamp 0
transform -1 0 9770 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4695_
timestamp 0
transform 1 0 10610 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4696_
timestamp 0
transform 1 0 10930 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4697_
timestamp 0
transform 1 0 11410 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4698_
timestamp 0
transform 1 0 11250 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4699_
timestamp 0
transform 1 0 11250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4700_
timestamp 0
transform 1 0 11090 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4701_
timestamp 0
transform -1 0 11470 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4702_
timestamp 0
transform 1 0 11450 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4703_
timestamp 0
transform 1 0 11730 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4704_
timestamp 0
transform -1 0 11630 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4705_
timestamp 0
transform -1 0 11830 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4706_
timestamp 0
transform -1 0 11770 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4707_
timestamp 0
transform 1 0 10710 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4708_
timestamp 0
transform 1 0 10910 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4709_
timestamp 0
transform -1 0 10910 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4710_
timestamp 0
transform -1 0 10710 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4711_
timestamp 0
transform 1 0 10170 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4712_
timestamp 0
transform -1 0 9950 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4713_
timestamp 0
transform 1 0 9750 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4714_
timestamp 0
transform 1 0 9550 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4715_
timestamp 0
transform -1 0 9870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4716_
timestamp 0
transform 1 0 9290 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4717_
timestamp 0
transform 1 0 9630 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4718_
timestamp 0
transform -1 0 8770 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4719_
timestamp 0
transform 1 0 11310 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4720_
timestamp 0
transform 1 0 10050 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4721_
timestamp 0
transform 1 0 9870 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4722_
timestamp 0
transform -1 0 9950 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4723_
timestamp 0
transform -1 0 9950 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4724_
timestamp 0
transform 1 0 4250 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4725_
timestamp 0
transform -1 0 10150 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4726_
timestamp 0
transform -1 0 10350 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4727_
timestamp 0
transform -1 0 11110 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4728_
timestamp 0
transform 1 0 10190 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4729_
timestamp 0
transform -1 0 10130 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4730_
timestamp 0
transform -1 0 10010 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4731_
timestamp 0
transform -1 0 11690 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4732_
timestamp 0
transform -1 0 9850 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4733_
timestamp 0
transform 1 0 9830 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4734_
timestamp 0
transform -1 0 7810 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4735_
timestamp 0
transform 1 0 9350 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4736_
timestamp 0
transform -1 0 10050 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4737_
timestamp 0
transform 1 0 9550 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4738_
timestamp 0
transform -1 0 9750 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4739_
timestamp 0
transform -1 0 9930 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4740_
timestamp 0
transform -1 0 10310 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4741_
timestamp 0
transform -1 0 10130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4742_
timestamp 0
transform 1 0 10350 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4743_
timestamp 0
transform 1 0 10110 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4744_
timestamp 0
transform 1 0 10610 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4745_
timestamp 0
transform 1 0 10930 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4746_
timestamp 0
transform 1 0 10410 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4747_
timestamp 0
transform 1 0 8350 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4748_
timestamp 0
transform 1 0 8550 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4749_
timestamp 0
transform -1 0 8790 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4750_
timestamp 0
transform 1 0 8550 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4751_
timestamp 0
transform 1 0 3750 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4752_
timestamp 0
transform -1 0 9150 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4753_
timestamp 0
transform -1 0 8030 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4754_
timestamp 0
transform 1 0 8150 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4755_
timestamp 0
transform 1 0 7270 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4756_
timestamp 0
transform 1 0 6930 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4757_
timestamp 0
transform 1 0 8370 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4758_
timestamp 0
transform -1 0 10430 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4759_
timestamp 0
transform 1 0 10790 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4760_
timestamp 0
transform -1 0 11070 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4761_
timestamp 0
transform 1 0 11350 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4762_
timestamp 0
transform -1 0 10510 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4763_
timestamp 0
transform 1 0 11850 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4764_
timestamp 0
transform 1 0 10890 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4765_
timestamp 0
transform -1 0 11150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4766_
timestamp 0
transform -1 0 10510 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4767_
timestamp 0
transform -1 0 10530 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4768_
timestamp 0
transform 1 0 10310 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4769_
timestamp 0
transform 1 0 10690 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4770_
timestamp 0
transform 1 0 11170 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4771_
timestamp 0
transform 1 0 12030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4772_
timestamp 0
transform 1 0 9370 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4773_
timestamp 0
transform -1 0 8830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4774_
timestamp 0
transform 1 0 2570 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4775_
timestamp 0
transform 1 0 2730 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4776_
timestamp 0
transform 1 0 2890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4777_
timestamp 0
transform -1 0 3110 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4778_
timestamp 0
transform -1 0 3710 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4779_
timestamp 0
transform 1 0 3890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4780_
timestamp 0
transform -1 0 8770 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4781_
timestamp 0
transform 1 0 3610 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4782_
timestamp 0
transform 1 0 3290 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4783_
timestamp 0
transform 1 0 9110 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4784_
timestamp 0
transform 1 0 7750 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4785_
timestamp 0
transform 1 0 2110 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4786_
timestamp 0
transform -1 0 3990 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__4787_
timestamp 0
transform -1 0 3670 0 1 3130
box -6 -8 26 248
use FILL  FILL_3__4788_
timestamp 0
transform -1 0 4190 0 1 3610
box -6 -8 26 248
use FILL  FILL_3__4789_
timestamp 0
transform 1 0 7230 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4790_
timestamp 0
transform 1 0 7290 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4791_
timestamp 0
transform -1 0 7830 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4792_
timestamp 0
transform -1 0 7890 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4793_
timestamp 0
transform -1 0 7830 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4794_
timestamp 0
transform -1 0 7470 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4795_
timestamp 0
transform -1 0 7530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4796_
timestamp 0
transform 1 0 11830 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4797_
timestamp 0
transform 1 0 8570 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4798_
timestamp 0
transform 1 0 10030 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4799_
timestamp 0
transform -1 0 9870 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4800_
timestamp 0
transform 1 0 8510 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4801_
timestamp 0
transform 1 0 10970 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4802_
timestamp 0
transform -1 0 10510 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4803_
timestamp 0
transform -1 0 7410 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4804_
timestamp 0
transform -1 0 7090 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4805_
timestamp 0
transform -1 0 6970 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4806_
timestamp 0
transform -1 0 9330 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4807_
timestamp 0
transform -1 0 9110 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4808_
timestamp 0
transform -1 0 8730 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4809_
timestamp 0
transform -1 0 8730 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4810_
timestamp 0
transform -1 0 8970 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4811_
timestamp 0
transform 1 0 11950 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4812_
timestamp 0
transform 1 0 12030 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4813_
timestamp 0
transform 1 0 11490 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4814_
timestamp 0
transform 1 0 11370 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4815_
timestamp 0
transform -1 0 9070 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4816_
timestamp 0
transform -1 0 9510 0 1 7450
box -6 -8 26 248
use FILL  FILL_3__4817_
timestamp 0
transform -1 0 11570 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4818_
timestamp 0
transform -1 0 11510 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4819_
timestamp 0
transform -1 0 6450 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4820_
timestamp 0
transform 1 0 8010 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4821_
timestamp 0
transform 1 0 11650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4822_
timestamp 0
transform 1 0 11850 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4823_
timestamp 0
transform 1 0 11630 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4824_
timestamp 0
transform -1 0 11490 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4825_
timestamp 0
transform 1 0 11190 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4826_
timestamp 0
transform -1 0 11030 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4827_
timestamp 0
transform -1 0 11730 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4828_
timestamp 0
transform -1 0 11810 0 1 10330
box -6 -8 26 248
use FILL  FILL_3__4829_
timestamp 0
transform 1 0 11650 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4830_
timestamp 0
transform 1 0 9010 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4831_
timestamp 0
transform -1 0 9370 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4832_
timestamp 0
transform 1 0 11910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4833_
timestamp 0
transform 1 0 8390 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4834_
timestamp 0
transform 1 0 8190 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4835_
timestamp 0
transform -1 0 8390 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4836_
timestamp 0
transform 1 0 9670 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4837_
timestamp 0
transform -1 0 10810 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4838_
timestamp 0
transform 1 0 11830 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4839_
timestamp 0
transform 1 0 12090 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4840_
timestamp 0
transform 1 0 9270 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4841_
timestamp 0
transform 1 0 10310 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4842_
timestamp 0
transform 1 0 12010 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4843_
timestamp 0
transform 1 0 11170 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4844_
timestamp 0
transform -1 0 11150 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4845_
timestamp 0
transform -1 0 11930 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4846_
timestamp 0
transform 1 0 11910 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4847_
timestamp 0
transform -1 0 8390 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3__4848_
timestamp 0
transform -1 0 8410 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4849_
timestamp 0
transform 1 0 9070 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4850_
timestamp 0
transform 1 0 9310 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4851_
timestamp 0
transform 1 0 11290 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4852_
timestamp 0
transform 1 0 11670 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4853_
timestamp 0
transform 1 0 12070 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4854_
timestamp 0
transform -1 0 11210 0 1 11770
box -6 -8 26 248
use FILL  FILL_3__4855_
timestamp 0
transform -1 0 8230 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4856_
timestamp 0
transform -1 0 8250 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4857_
timestamp 0
transform -1 0 10330 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4858_
timestamp 0
transform -1 0 10470 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4859_
timestamp 0
transform -1 0 7210 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4860_
timestamp 0
transform -1 0 10390 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4861_
timestamp 0
transform -1 0 10650 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4862_
timestamp 0
transform 1 0 11450 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4863_
timestamp 0
transform -1 0 10710 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4864_
timestamp 0
transform -1 0 10550 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4865_
timestamp 0
transform 1 0 10570 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4866_
timestamp 0
transform 1 0 11650 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4867_
timestamp 0
transform 1 0 11830 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4868_
timestamp 0
transform -1 0 11330 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4869_
timestamp 0
transform -1 0 10870 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3__4870_
timestamp 0
transform 1 0 8110 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4871_
timestamp 0
transform 1 0 7950 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4872_
timestamp 0
transform 1 0 7850 0 1 7930
box -6 -8 26 248
use FILL  FILL_3__4873_
timestamp 0
transform -1 0 11370 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4874_
timestamp 0
transform 1 0 11890 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4875_
timestamp 0
transform -1 0 7590 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3__4876_
timestamp 0
transform -1 0 10510 0 -1 9370
box -6 -8 26 248
use FILL  FILL_3__4877_
timestamp 0
transform 1 0 10910 0 1 8410
box -6 -8 26 248
use FILL  FILL_3__4878_
timestamp 0
transform 1 0 11350 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4879_
timestamp 0
transform 1 0 12010 0 1 9850
box -6 -8 26 248
use FILL  FILL_3__4880_
timestamp 0
transform -1 0 12070 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4881_
timestamp 0
transform -1 0 9110 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4882_
timestamp 0
transform 1 0 12030 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4883_
timestamp 0
transform 1 0 11850 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4884_
timestamp 0
transform 1 0 11670 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4885_
timestamp 0
transform -1 0 11710 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4886_
timestamp 0
transform 1 0 10970 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4887_
timestamp 0
transform 1 0 11010 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4888_
timestamp 0
transform 1 0 11670 0 1 8890
box -6 -8 26 248
use FILL  FILL_3__4889_
timestamp 0
transform 1 0 12010 0 1 9370
box -6 -8 26 248
use FILL  FILL_3__4890_
timestamp 0
transform 1 0 11530 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4891_
timestamp 0
transform 1 0 11870 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3__4892_
timestamp 0
transform -1 0 12090 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3__4893_
timestamp 0
transform -1 0 2510 0 -1 7450
box -6 -8 26 248
use FILL  FILL_3__4894_
timestamp 0
transform 1 0 9710 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4895_
timestamp 0
transform 1 0 8450 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4896_
timestamp 0
transform -1 0 9490 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4897_
timestamp 0
transform 1 0 9530 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4898_
timestamp 0
transform 1 0 9710 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4899_
timestamp 0
transform -1 0 9190 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4900_
timestamp 0
transform -1 0 9530 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4901_
timestamp 0
transform -1 0 9910 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4902_
timestamp 0
transform 1 0 10230 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4903_
timestamp 0
transform 1 0 9690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4904_
timestamp 0
transform -1 0 10410 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4905_
timestamp 0
transform 1 0 9690 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4906_
timestamp 0
transform -1 0 9870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4907_
timestamp 0
transform -1 0 9530 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4908_
timestamp 0
transform 1 0 10030 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4909_
timestamp 0
transform 1 0 10970 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4910_
timestamp 0
transform -1 0 11350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4911_
timestamp 0
transform 1 0 11290 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4912_
timestamp 0
transform 1 0 11110 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4913_
timestamp 0
transform -1 0 10930 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4914_
timestamp 0
transform 1 0 11490 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4915_
timestamp 0
transform -1 0 10790 0 1 6970
box -6 -8 26 248
use FILL  FILL_3__4916_
timestamp 0
transform 1 0 10550 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4917_
timestamp 0
transform -1 0 10610 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4918_
timestamp 0
transform -1 0 10970 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4919_
timestamp 0
transform 1 0 11130 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4920_
timestamp 0
transform 1 0 8550 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4921_
timestamp 0
transform -1 0 8770 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4922_
timestamp 0
transform -1 0 8970 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4923_
timestamp 0
transform 1 0 9350 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4924_
timestamp 0
transform 1 0 9330 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4925_
timestamp 0
transform -1 0 9150 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4926_
timestamp 0
transform 1 0 8910 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4927_
timestamp 0
transform -1 0 11310 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4928_
timestamp 0
transform 1 0 11490 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4929_
timestamp 0
transform 1 0 12070 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4930_
timestamp 0
transform 1 0 11650 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4931_
timestamp 0
transform -1 0 11870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4932_
timestamp 0
transform -1 0 11710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4933_
timestamp 0
transform -1 0 11150 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4934_
timestamp 0
transform 1 0 10930 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4935_
timestamp 0
transform -1 0 10750 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4936_
timestamp 0
transform -1 0 9650 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4937_
timestamp 0
transform -1 0 9870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4938_
timestamp 0
transform 1 0 10030 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4939_
timestamp 0
transform 1 0 10110 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4940_
timestamp 0
transform 1 0 10210 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3__4941_
timestamp 0
transform 1 0 10310 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4942_
timestamp 0
transform -1 0 10710 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4943_
timestamp 0
transform 1 0 11690 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4944_
timestamp 0
transform -1 0 11910 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4945_
timestamp 0
transform 1 0 11850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4946_
timestamp 0
transform -1 0 11830 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4947_
timestamp 0
transform -1 0 8650 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4948_
timestamp 0
transform 1 0 8970 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4949_
timestamp 0
transform 1 0 12090 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__4950_
timestamp 0
transform -1 0 12050 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4951_
timestamp 0
transform -1 0 8590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4952_
timestamp 0
transform 1 0 8970 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4953_
timestamp 0
transform -1 0 8870 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4954_
timestamp 0
transform -1 0 9170 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4955_
timestamp 0
transform -1 0 8730 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__4956_
timestamp 0
transform -1 0 8810 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4957_
timestamp 0
transform -1 0 8670 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4958_
timestamp 0
transform -1 0 11050 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4959_
timestamp 0
transform 1 0 11230 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4960_
timestamp 0
transform -1 0 11450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4961_
timestamp 0
transform 1 0 11630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4962_
timestamp 0
transform 1 0 12030 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4963_
timestamp 0
transform 1 0 11990 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4964_
timestamp 0
transform 1 0 11990 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4965_
timestamp 0
transform -1 0 11830 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4966_
timestamp 0
transform -1 0 9170 0 1 4090
box -6 -8 26 248
use FILL  FILL_3__4967_
timestamp 0
transform 1 0 8090 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__4968_
timestamp 0
transform 1 0 11670 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4969_
timestamp 0
transform 1 0 12030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4970_
timestamp 0
transform 1 0 9070 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4971_
timestamp 0
transform -1 0 8290 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4972_
timestamp 0
transform -1 0 8690 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4973_
timestamp 0
transform -1 0 8850 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4974_
timestamp 0
transform 1 0 8750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4975_
timestamp 0
transform 1 0 8950 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4976_
timestamp 0
transform 1 0 11610 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4977_
timestamp 0
transform 1 0 11410 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4978_
timestamp 0
transform 1 0 11430 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4979_
timestamp 0
transform 1 0 11450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4980_
timestamp 0
transform 1 0 11830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4981_
timestamp 0
transform -1 0 11830 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4982_
timestamp 0
transform -1 0 11850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4983_
timestamp 0
transform 1 0 11630 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4984_
timestamp 0
transform 1 0 11250 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4985_
timestamp 0
transform -1 0 8070 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4986_
timestamp 0
transform 1 0 9110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4987_
timestamp 0
transform 1 0 11630 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4988_
timestamp 0
transform -1 0 11850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4989_
timestamp 0
transform -1 0 11450 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4990_
timestamp 0
transform -1 0 11270 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__4991_
timestamp 0
transform 1 0 11650 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__4992_
timestamp 0
transform -1 0 11510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4993_
timestamp 0
transform 1 0 11290 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__4994_
timestamp 0
transform 1 0 9310 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__4995_
timestamp 0
transform -1 0 9890 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4996_
timestamp 0
transform 1 0 9250 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4997_
timestamp 0
transform -1 0 9330 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__4998_
timestamp 0
transform 1 0 9430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__4999_
timestamp 0
transform -1 0 9290 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5000_
timestamp 0
transform 1 0 11030 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__5001_
timestamp 0
transform -1 0 10850 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__5002_
timestamp 0
transform -1 0 10670 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5003_
timestamp 0
transform -1 0 10730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5004_
timestamp 0
transform 1 0 10910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5005_
timestamp 0
transform -1 0 10890 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5006_
timestamp 0
transform 1 0 11410 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5007_
timestamp 0
transform 1 0 12010 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5008_
timestamp 0
transform 1 0 11990 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__5009_
timestamp 0
transform 1 0 12010 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5010_
timestamp 0
transform -1 0 11310 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__5011_
timestamp 0
transform 1 0 11810 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5012_
timestamp 0
transform 1 0 11610 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5013_
timestamp 0
transform -1 0 10290 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5014_
timestamp 0
transform -1 0 9510 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5015_
timestamp 0
transform 1 0 8270 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5016_
timestamp 0
transform 1 0 10670 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5017_
timestamp 0
transform 1 0 8930 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5018_
timestamp 0
transform 1 0 8470 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5019_
timestamp 0
transform 1 0 9150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5020_
timestamp 0
transform 1 0 9050 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5021_
timestamp 0
transform 1 0 9330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5022_
timestamp 0
transform -1 0 9130 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5023_
timestamp 0
transform -1 0 10850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__5024_
timestamp 0
transform 1 0 10850 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5025_
timestamp 0
transform -1 0 11070 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5026_
timestamp 0
transform 1 0 11090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__5027_
timestamp 0
transform -1 0 10890 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5028_
timestamp 0
transform -1 0 10710 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5029_
timestamp 0
transform 1 0 11050 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5030_
timestamp 0
transform 1 0 11070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5031_
timestamp 0
transform 1 0 11830 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__5032_
timestamp 0
transform 1 0 11670 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__5033_
timestamp 0
transform -1 0 8990 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__5034_
timestamp 0
transform -1 0 9190 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__5035_
timestamp 0
transform 1 0 11210 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5036_
timestamp 0
transform 1 0 9890 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5037_
timestamp 0
transform 1 0 9690 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5038_
timestamp 0
transform 1 0 9530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5039_
timestamp 0
transform 1 0 9470 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5040_
timestamp 0
transform 1 0 9710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5041_
timestamp 0
transform 1 0 9910 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5042_
timestamp 0
transform 1 0 10630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__5043_
timestamp 0
transform 1 0 10450 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5044_
timestamp 0
transform 1 0 10510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5045_
timestamp 0
transform -1 0 10490 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5046_
timestamp 0
transform 1 0 10930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__5047_
timestamp 0
transform 1 0 11030 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5048_
timestamp 0
transform 1 0 11470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__5049_
timestamp 0
transform -1 0 11310 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__5050_
timestamp 0
transform -1 0 9370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__5051_
timestamp 0
transform 1 0 8370 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__5052_
timestamp 0
transform -1 0 10530 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__5053_
timestamp 0
transform -1 0 10770 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__5054_
timestamp 0
transform -1 0 10410 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__5055_
timestamp 0
transform 1 0 8530 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__5056_
timestamp 0
transform 1 0 8150 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__5057_
timestamp 0
transform 1 0 8370 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__5058_
timestamp 0
transform -1 0 8190 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__5059_
timestamp 0
transform 1 0 8010 0 1 6490
box -6 -8 26 248
use FILL  FILL_3__5060_
timestamp 0
transform -1 0 7650 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__5061_
timestamp 0
transform -1 0 7830 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__5062_
timestamp 0
transform 1 0 7990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3__5063_
timestamp 0
transform -1 0 8030 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__5064_
timestamp 0
transform -1 0 7550 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5065_
timestamp 0
transform -1 0 7750 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5066_
timestamp 0
transform -1 0 7690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5067_
timestamp 0
transform -1 0 8390 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5068_
timestamp 0
transform -1 0 8410 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5069_
timestamp 0
transform -1 0 8250 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5070_
timestamp 0
transform -1 0 7870 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5071_
timestamp 0
transform 1 0 8050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5072_
timestamp 0
transform -1 0 7510 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5073_
timestamp 0
transform 1 0 7310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5074_
timestamp 0
transform 1 0 4870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3__5075_
timestamp 0
transform 1 0 10270 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__5076_
timestamp 0
transform 1 0 10070 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__5077_
timestamp 0
transform 1 0 9850 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__5078_
timestamp 0
transform 1 0 9630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__5079_
timestamp 0
transform 1 0 10030 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__5080_
timestamp 0
transform 1 0 10230 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__5081_
timestamp 0
transform 1 0 10450 0 1 6010
box -6 -8 26 248
use FILL  FILL_3__5082_
timestamp 0
transform 1 0 10430 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3__5083_
timestamp 0
transform -1 0 10330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5084_
timestamp 0
transform -1 0 9710 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5085_
timestamp 0
transform 1 0 8550 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5086_
timestamp 0
transform -1 0 8750 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5087_
timestamp 0
transform -1 0 10910 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__5088_
timestamp 0
transform -1 0 10690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__5089_
timestamp 0
transform -1 0 10490 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__5090_
timestamp 0
transform -1 0 10270 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5091_
timestamp 0
transform 1 0 10110 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3__5092_
timestamp 0
transform 1 0 9950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__5093_
timestamp 0
transform -1 0 10130 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__5094_
timestamp 0
transform 1 0 10270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__5095_
timestamp 0
transform -1 0 9790 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__5096_
timestamp 0
transform 1 0 8930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__5097_
timestamp 0
transform 1 0 8250 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3__5098_
timestamp 0
transform 1 0 9750 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5099_
timestamp 0
transform 1 0 9930 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5100_
timestamp 0
transform 1 0 9370 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5101_
timestamp 0
transform -1 0 10090 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5102_
timestamp 0
transform -1 0 9910 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5103_
timestamp 0
transform 1 0 10050 0 1 5050
box -6 -8 26 248
use FILL  FILL_3__5104_
timestamp 0
transform -1 0 10350 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5105_
timestamp 0
transform -1 0 10150 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5106_
timestamp 0
transform -1 0 10530 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5107_
timestamp 0
transform 1 0 10510 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__5108_
timestamp 0
transform -1 0 11110 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__5109_
timestamp 0
transform 1 0 10710 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3__5110_
timestamp 0
transform -1 0 9570 0 1 4570
box -6 -8 26 248
use FILL  FILL_3__5111_
timestamp 0
transform -1 0 7930 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5112_
timestamp 0
transform -1 0 8110 0 1 5530
box -6 -8 26 248
use FILL  FILL_3__5124_
timestamp 0
transform 1 0 1790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__5125_
timestamp 0
transform -1 0 650 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__5126_
timestamp 0
transform -1 0 830 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__5127_
timestamp 0
transform 1 0 790 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__5128_
timestamp 0
transform 1 0 550 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__5129_
timestamp 0
transform 1 0 990 0 1 2170
box -6 -8 26 248
use FILL  FILL_3__5130_
timestamp 0
transform 1 0 990 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__5131_
timestamp 0
transform -1 0 2310 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5132_
timestamp 0
transform -1 0 5550 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5133_
timestamp 0
transform 1 0 5290 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5134_
timestamp 0
transform 1 0 1370 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__5135_
timestamp 0
transform 1 0 2170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__5136_
timestamp 0
transform 1 0 1970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__5137_
timestamp 0
transform -1 0 1110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__5138_
timestamp 0
transform -1 0 1290 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__5139_
timestamp 0
transform -1 0 3670 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5140_
timestamp 0
transform 1 0 4130 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__5141_
timestamp 0
transform -1 0 4310 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__5142_
timestamp 0
transform -1 0 4190 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__5143_
timestamp 0
transform -1 0 4410 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5144_
timestamp 0
transform 1 0 5570 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5145_
timestamp 0
transform -1 0 4110 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5146_
timestamp 0
transform -1 0 4630 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5147_
timestamp 0
transform 1 0 4730 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5148_
timestamp 0
transform 1 0 4930 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5149_
timestamp 0
transform 1 0 5450 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5150_
timestamp 0
transform -1 0 6070 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5151_
timestamp 0
transform 1 0 3450 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5152_
timestamp 0
transform 1 0 5710 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5153_
timestamp 0
transform 1 0 4190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__5154_
timestamp 0
transform 1 0 5390 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5155_
timestamp 0
transform 1 0 5350 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5156_
timestamp 0
transform 1 0 5510 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5157_
timestamp 0
transform 1 0 5650 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5158_
timestamp 0
transform 1 0 4530 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5159_
timestamp 0
transform -1 0 4650 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5160_
timestamp 0
transform 1 0 4970 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5161_
timestamp 0
transform 1 0 4810 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5162_
timestamp 0
transform 1 0 5850 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5163_
timestamp 0
transform -1 0 2750 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5164_
timestamp 0
transform 1 0 5870 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5165_
timestamp 0
transform -1 0 3810 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__5166_
timestamp 0
transform 1 0 4250 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5167_
timestamp 0
transform 1 0 4210 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5168_
timestamp 0
transform -1 0 4030 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5169_
timestamp 0
transform 1 0 2710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__5170_
timestamp 0
transform 1 0 3830 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5171_
timestamp 0
transform -1 0 4130 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__5172_
timestamp 0
transform -1 0 3630 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__5173_
timestamp 0
transform -1 0 4910 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__5174_
timestamp 0
transform -1 0 3810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__5175_
timestamp 0
transform 1 0 3650 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5176_
timestamp 0
transform -1 0 2650 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__5177_
timestamp 0
transform 1 0 3090 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5178_
timestamp 0
transform 1 0 4430 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5179_
timestamp 0
transform 1 0 4450 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5180_
timestamp 0
transform 1 0 4250 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5181_
timestamp 0
transform 1 0 3250 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5182_
timestamp 0
transform -1 0 2450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__5183_
timestamp 0
transform 1 0 2250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__5184_
timestamp 0
transform -1 0 2470 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__5185_
timestamp 0
transform -1 0 4030 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__5186_
timestamp 0
transform -1 0 3310 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__5187_
timestamp 0
transform -1 0 3050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__5188_
timestamp 0
transform 1 0 3750 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5189_
timestamp 0
transform -1 0 3690 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5190_
timestamp 0
transform 1 0 3230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__5191_
timestamp 0
transform 1 0 2910 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5192_
timestamp 0
transform -1 0 3630 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__5193_
timestamp 0
transform 1 0 6070 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5194_
timestamp 0
transform -1 0 2930 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__5195_
timestamp 0
transform -1 0 2850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__5196_
timestamp 0
transform 1 0 3590 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5197_
timestamp 0
transform -1 0 3510 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5198_
timestamp 0
transform -1 0 2910 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5199_
timestamp 0
transform 1 0 2470 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5200_
timestamp 0
transform -1 0 2690 0 -1 730
box -6 -8 26 248
use FILL  FILL_3__5201_
timestamp 0
transform -1 0 3970 0 1 1690
box -6 -8 26 248
use FILL  FILL_3__5202_
timestamp 0
transform 1 0 3930 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5203_
timestamp 0
transform -1 0 3470 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5204_
timestamp 0
transform 1 0 4090 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5205_
timestamp 0
transform -1 0 3930 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5206_
timestamp 0
transform -1 0 3270 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5207_
timestamp 0
transform 1 0 2490 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5208_
timestamp 0
transform 1 0 3030 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__5209_
timestamp 0
transform -1 0 4490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3__5210_
timestamp 0
transform 1 0 2690 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5211_
timestamp 0
transform 1 0 2850 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5212_
timestamp 0
transform 1 0 3430 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5213_
timestamp 0
transform 1 0 3310 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5214_
timestamp 0
transform -1 0 3070 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5215_
timestamp 0
transform 1 0 2290 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5216_
timestamp 0
transform -1 0 3090 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__5217_
timestamp 0
transform -1 0 6250 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5218_
timestamp 0
transform 1 0 3430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__5219_
timestamp 0
transform 1 0 3590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__5220_
timestamp 0
transform 1 0 4770 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5221_
timestamp 0
transform 1 0 4590 0 -1 250
box -6 -8 26 248
use FILL  FILL_3__5222_
timestamp 0
transform -1 0 4070 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5223_
timestamp 0
transform 1 0 3110 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5224_
timestamp 0
transform -1 0 3870 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5225_
timestamp 0
transform 1 0 5370 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__5226_
timestamp 0
transform 1 0 5150 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5227_
timestamp 0
transform -1 0 5330 0 1 250
box -6 -8 26 248
use FILL  FILL_3__5228_
timestamp 0
transform -1 0 4770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3__5229_
timestamp 0
transform -1 0 4810 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5230_
timestamp 0
transform 1 0 4990 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5231_
timestamp 0
transform 1 0 5190 0 1 730
box -6 -8 26 248
use FILL  FILL_3__5232_
timestamp 0
transform 1 0 3990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3__5233_
timestamp 0
transform 1 0 4370 0 1 1210
box -6 -8 26 248
use FILL  FILL_3__5234_
timestamp 0
transform -1 0 5170 0 1 1210
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert0
timestamp 0
transform -1 0 4210 0 1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert1
timestamp 0
transform 1 0 6130 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert2
timestamp 0
transform -1 0 3310 0 1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert3
timestamp 0
transform -1 0 3690 0 1 9850
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert4
timestamp 0
transform 1 0 9470 0 1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert5
timestamp 0
transform 1 0 11270 0 1 8410
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert6
timestamp 0
transform -1 0 9470 0 1 8410
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert7
timestamp 0
transform 1 0 12010 0 1 7930
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert8
timestamp 0
transform -1 0 7170 0 1 5530
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert9
timestamp 0
transform 1 0 6670 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert10
timestamp 0
transform 1 0 8710 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert11
timestamp 0
transform 1 0 6870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert12
timestamp 0
transform 1 0 8910 0 1 9850
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert13
timestamp 0
transform 1 0 7390 0 1 9850
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert14
timestamp 0
transform 1 0 650 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert15
timestamp 0
transform 1 0 70 0 1 9370
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert16
timestamp 0
transform 1 0 1890 0 1 5530
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert17
timestamp 0
transform -1 0 9150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert18
timestamp 0
transform -1 0 11510 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert19
timestamp 0
transform 1 0 10670 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert20
timestamp 0
transform -1 0 9190 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert21
timestamp 0
transform 1 0 2530 0 1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert22
timestamp 0
transform -1 0 1270 0 1 11290
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert23
timestamp 0
transform -1 0 1450 0 1 11290
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert24
timestamp 0
transform -1 0 1650 0 1 10330
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert38
timestamp 0
transform -1 0 11530 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert39
timestamp 0
transform -1 0 10670 0 1 6010
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert40
timestamp 0
transform 1 0 12030 0 1 6970
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert41
timestamp 0
transform -1 0 11250 0 1 6010
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert42
timestamp 0
transform 1 0 11450 0 1 730
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert43
timestamp 0
transform -1 0 11010 0 1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert44
timestamp 0
transform -1 0 10490 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert45
timestamp 0
transform -1 0 11370 0 1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert46
timestamp 0
transform -1 0 10750 0 1 3130
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert47
timestamp 0
transform 1 0 6210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert48
timestamp 0
transform -1 0 4770 0 1 1690
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert49
timestamp 0
transform 1 0 11570 0 1 1690
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert50
timestamp 0
transform -1 0 10410 0 1 1690
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert51
timestamp 0
transform 1 0 8170 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert52
timestamp 0
transform 1 0 10030 0 1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert53
timestamp 0
transform 1 0 9190 0 1 4570
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert54
timestamp 0
transform 1 0 9010 0 1 4570
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert55
timestamp 0
transform -1 0 9550 0 1 4090
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert56
timestamp 0
transform -1 0 8850 0 1 4570
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert57
timestamp 0
transform 1 0 11470 0 1 3130
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert58
timestamp 0
transform 1 0 10650 0 -1 730
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert59
timestamp 0
transform -1 0 7730 0 -1 730
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert60
timestamp 0
transform 1 0 11810 0 -1 730
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert61
timestamp 0
transform 1 0 11910 0 1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert62
timestamp 0
transform -1 0 4810 0 1 2170
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert63
timestamp 0
transform -1 0 9330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert64
timestamp 0
transform -1 0 11670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert65
timestamp 0
transform -1 0 9330 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert66
timestamp 0
transform -1 0 11510 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert67
timestamp 0
transform 1 0 6930 0 1 11290
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert68
timestamp 0
transform -1 0 3170 0 -1 10330
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert69
timestamp 0
transform -1 0 5630 0 1 10810
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert70
timestamp 0
transform 1 0 5110 0 -1 11290
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert71
timestamp 0
transform -1 0 3570 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert72
timestamp 0
transform 1 0 7110 0 1 11290
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert73
timestamp 0
transform 1 0 7130 0 1 730
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert74
timestamp 0
transform -1 0 6470 0 1 2170
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert75
timestamp 0
transform 1 0 7090 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert76
timestamp 0
transform 1 0 6550 0 1 730
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert77
timestamp 0
transform 1 0 10270 0 1 4090
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert78
timestamp 0
transform 1 0 9130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert79
timestamp 0
transform 1 0 10290 0 1 730
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert80
timestamp 0
transform -1 0 4950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert81
timestamp 0
transform -1 0 2810 0 1 5530
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert82
timestamp 0
transform -1 0 4030 0 -1 5530
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert83
timestamp 0
transform -1 0 6290 0 1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert84
timestamp 0
transform 1 0 7350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert85
timestamp 0
transform -1 0 3270 0 1 8410
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert86
timestamp 0
transform 1 0 3970 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert87
timestamp 0
transform -1 0 3230 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert88
timestamp 0
transform 1 0 7890 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert89
timestamp 0
transform -1 0 4730 0 1 9850
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert90
timestamp 0
transform 1 0 5570 0 1 9370
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert91
timestamp 0
transform 1 0 9030 0 1 10330
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert92
timestamp 0
transform -1 0 8530 0 1 10810
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert93
timestamp 0
transform -1 0 10930 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert94
timestamp 0
transform 1 0 7270 0 1 10330
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert95
timestamp 0
transform 1 0 11530 0 1 10810
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert96
timestamp 0
transform -1 0 4990 0 1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert97
timestamp 0
transform 1 0 610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert98
timestamp 0
transform -1 0 4010 0 1 7930
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert99
timestamp 0
transform 1 0 550 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert100
timestamp 0
transform 1 0 3030 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert101
timestamp 0
transform -1 0 490 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert102
timestamp 0
transform 1 0 3730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert103
timestamp 0
transform -1 0 3650 0 1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert104
timestamp 0
transform 1 0 4630 0 1 10330
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert105
timestamp 0
transform 1 0 290 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert106
timestamp 0
transform 1 0 6510 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert107
timestamp 0
transform -1 0 6210 0 1 730
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert108
timestamp 0
transform 1 0 5690 0 1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert109
timestamp 0
transform 1 0 7830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert110
timestamp 0
transform -1 0 5330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert111
timestamp 0
transform 1 0 7290 0 1 1690
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert112
timestamp 0
transform 1 0 10670 0 1 11770
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert113
timestamp 0
transform -1 0 12110 0 1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert114
timestamp 0
transform -1 0 10310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert115
timestamp 0
transform 1 0 7370 0 1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert116
timestamp 0
transform -1 0 5510 0 1 2170
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert117
timestamp 0
transform -1 0 5490 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert118
timestamp 0
transform -1 0 11190 0 1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert119
timestamp 0
transform 1 0 10370 0 1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert120
timestamp 0
transform -1 0 11110 0 1 730
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert121
timestamp 0
transform -1 0 8170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert122
timestamp 0
transform 1 0 11190 0 1 2170
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert123
timestamp 0
transform -1 0 10030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert124
timestamp 0
transform -1 0 8010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert125
timestamp 0
transform -1 0 5330 0 1 2170
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert126
timestamp 0
transform 1 0 12010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert127
timestamp 0
transform 1 0 10770 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert128
timestamp 0
transform -1 0 12050 0 -1 4090
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert129
timestamp 0
transform 1 0 10450 0 1 4090
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert130
timestamp 0
transform 1 0 12010 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert131
timestamp 0
transform -1 0 9370 0 1 4090
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert132
timestamp 0
transform -1 0 8710 0 1 730
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert133
timestamp 0
transform 1 0 12010 0 1 730
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert134
timestamp 0
transform -1 0 11390 0 1 4090
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert135
timestamp 0
transform -1 0 9110 0 -1 250
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert136
timestamp 0
transform 1 0 9470 0 -1 250
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert137
timestamp 0
transform -1 0 6390 0 1 730
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert138
timestamp 0
transform 1 0 8370 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert139
timestamp 0
transform -1 0 6410 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert140
timestamp 0
transform 1 0 9430 0 1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert141
timestamp 0
transform -1 0 7050 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert142
timestamp 0
transform -1 0 7030 0 1 8410
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert143
timestamp 0
transform -1 0 6450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert144
timestamp 0
transform -1 0 6270 0 1 6970
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert145
timestamp 0
transform 1 0 9550 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert146
timestamp 0
transform 1 0 9650 0 1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert147
timestamp 0
transform -1 0 7730 0 1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert148
timestamp 0
transform -1 0 7650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert149
timestamp 0
transform -1 0 9230 0 -1 7930
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert150
timestamp 0
transform -1 0 7230 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert151
timestamp 0
transform 1 0 7330 0 -1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert152
timestamp 0
transform -1 0 8230 0 1 9370
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert153
timestamp 0
transform 1 0 10070 0 -1 9850
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert154
timestamp 0
transform 1 0 10750 0 -1 8410
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert155
timestamp 0
transform 1 0 6390 0 1 3130
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert156
timestamp 0
transform 1 0 9130 0 -1 3130
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert157
timestamp 0
transform -1 0 5870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert158
timestamp 0
transform 1 0 9870 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert159
timestamp 0
transform 1 0 8730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert160
timestamp 0
transform 1 0 10370 0 1 9850
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert161
timestamp 0
transform 1 0 9270 0 1 9850
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert162
timestamp 0
transform 1 0 10230 0 1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert163
timestamp 0
transform -1 0 8330 0 1 8890
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert164
timestamp 0
transform 1 0 11730 0 1 4090
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert165
timestamp 0
transform -1 0 8790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert166
timestamp 0
transform -1 0 11570 0 1 4090
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert167
timestamp 0
transform 1 0 11730 0 1 11770
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert168
timestamp 0
transform -1 0 11310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3_BUFX2_insert169
timestamp 0
transform 1 0 4930 0 1 1690
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert25
timestamp 0
transform 1 0 1370 0 1 2170
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert26
timestamp 0
transform 1 0 4030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert27
timestamp 0
transform -1 0 90 0 -1 2650
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert28
timestamp 0
transform -1 0 2730 0 1 9370
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert29
timestamp 0
transform 1 0 70 0 -1 2170
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert30
timestamp 0
transform 1 0 6190 0 -1 5050
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert31
timestamp 0
transform 1 0 790 0 -1 6010
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert32
timestamp 0
transform -1 0 4830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert33
timestamp 0
transform -1 0 970 0 -1 10810
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert34
timestamp 0
transform 1 0 1410 0 -1 6490
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert35
timestamp 0
transform -1 0 330 0 -1 11770
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert36
timestamp 0
transform 1 0 70 0 1 5530
box -6 -8 26 248
use FILL  FILL_3_CLKBUF1_insert37
timestamp 0
transform 1 0 6150 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__2478_
timestamp 0
transform -1 0 110 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2479_
timestamp 0
transform -1 0 110 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2480_
timestamp 0
transform 1 0 1950 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2481_
timestamp 0
transform 1 0 2770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2482_
timestamp 0
transform -1 0 110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__2483_
timestamp 0
transform -1 0 590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__2484_
timestamp 0
transform -1 0 2150 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2485_
timestamp 0
transform 1 0 3970 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2486_
timestamp 0
transform 1 0 12090 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2487_
timestamp 0
transform -1 0 6670 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2489_
timestamp 0
transform 1 0 12050 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2490_
timestamp 0
transform 1 0 12050 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2491_
timestamp 0
transform 1 0 6470 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2492_
timestamp 0
transform 1 0 11870 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2493_
timestamp 0
transform -1 0 11970 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2494_
timestamp 0
transform -1 0 1070 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__2495_
timestamp 0
transform -1 0 1230 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2496_
timestamp 0
transform -1 0 110 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__2497_
timestamp 0
transform -1 0 4450 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2498_
timestamp 0
transform 1 0 4490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2499_
timestamp 0
transform -1 0 3310 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2500_
timestamp 0
transform -1 0 490 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2501_
timestamp 0
transform -1 0 3690 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2502_
timestamp 0
transform -1 0 110 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__2503_
timestamp 0
transform -1 0 110 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2504_
timestamp 0
transform 1 0 4590 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2505_
timestamp 0
transform 1 0 5130 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2506_
timestamp 0
transform -1 0 2570 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2507_
timestamp 0
transform 1 0 3850 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2509_
timestamp 0
transform 1 0 4250 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2510_
timestamp 0
transform 1 0 3110 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2511_
timestamp 0
transform -1 0 4970 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2519_
timestamp 0
transform -1 0 5710 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2520_
timestamp 0
transform -1 0 7570 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2521_
timestamp 0
transform -1 0 7770 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2522_
timestamp 0
transform 1 0 7770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2523_
timestamp 0
transform 1 0 9510 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2524_
timestamp 0
transform -1 0 7830 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2525_
timestamp 0
transform 1 0 7570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2526_
timestamp 0
transform 1 0 8310 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2527_
timestamp 0
transform 1 0 8510 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2528_
timestamp 0
transform -1 0 9650 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2529_
timestamp 0
transform 1 0 8590 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2530_
timestamp 0
transform -1 0 8230 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2531_
timestamp 0
transform -1 0 8370 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2532_
timestamp 0
transform -1 0 8790 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2533_
timestamp 0
transform 1 0 9530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2534_
timestamp 0
transform 1 0 10090 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__2536_
timestamp 0
transform -1 0 8790 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2537_
timestamp 0
transform -1 0 8590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2538_
timestamp 0
transform -1 0 8390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2539_
timestamp 0
transform 1 0 7990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2540_
timestamp 0
transform -1 0 10690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2541_
timestamp 0
transform -1 0 10890 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2542_
timestamp 0
transform 1 0 10930 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2543_
timestamp 0
transform -1 0 10630 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2544_
timestamp 0
transform -1 0 5730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2545_
timestamp 0
transform -1 0 5930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2546_
timestamp 0
transform -1 0 6150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2547_
timestamp 0
transform -1 0 6030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2548_
timestamp 0
transform -1 0 6230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2549_
timestamp 0
transform 1 0 5610 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2550_
timestamp 0
transform 1 0 5810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2551_
timestamp 0
transform -1 0 6930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2552_
timestamp 0
transform -1 0 7290 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2553_
timestamp 0
transform -1 0 5750 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2554_
timestamp 0
transform -1 0 6390 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2556_
timestamp 0
transform -1 0 6770 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2557_
timestamp 0
transform -1 0 6250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2558_
timestamp 0
transform 1 0 6530 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2559_
timestamp 0
transform 1 0 6910 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2560_
timestamp 0
transform -1 0 5950 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2561_
timestamp 0
transform -1 0 6590 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2562_
timestamp 0
transform 1 0 6770 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2563_
timestamp 0
transform -1 0 6150 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2564_
timestamp 0
transform 1 0 7810 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2565_
timestamp 0
transform 1 0 8030 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2566_
timestamp 0
transform 1 0 7610 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2567_
timestamp 0
transform 1 0 7010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2568_
timestamp 0
transform -1 0 6650 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2569_
timestamp 0
transform 1 0 7230 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2570_
timestamp 0
transform -1 0 9410 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2571_
timestamp 0
transform -1 0 9310 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2572_
timestamp 0
transform 1 0 9330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2573_
timestamp 0
transform 1 0 9210 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2574_
timestamp 0
transform -1 0 9290 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2576_
timestamp 0
transform -1 0 8830 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2577_
timestamp 0
transform -1 0 9030 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2578_
timestamp 0
transform 1 0 9590 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2579_
timestamp 0
transform -1 0 9530 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2580_
timestamp 0
transform -1 0 8330 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2581_
timestamp 0
transform 1 0 8290 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2582_
timestamp 0
transform 1 0 8410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2583_
timestamp 0
transform -1 0 9810 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2584_
timestamp 0
transform 1 0 9470 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2585_
timestamp 0
transform -1 0 11210 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2586_
timestamp 0
transform 1 0 8890 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2587_
timestamp 0
transform 1 0 8690 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2588_
timestamp 0
transform -1 0 8510 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2589_
timestamp 0
transform 1 0 8550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2590_
timestamp 0
transform 1 0 8290 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2591_
timestamp 0
transform -1 0 8630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2592_
timestamp 0
transform 1 0 7890 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2593_
timestamp 0
transform -1 0 9130 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2594_
timestamp 0
transform -1 0 9030 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2596_
timestamp 0
transform 1 0 10470 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2597_
timestamp 0
transform 1 0 10650 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2598_
timestamp 0
transform -1 0 10490 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2599_
timestamp 0
transform 1 0 10850 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2600_
timestamp 0
transform -1 0 11450 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2601_
timestamp 0
transform 1 0 8310 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2602_
timestamp 0
transform -1 0 8110 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2603_
timestamp 0
transform 1 0 7110 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2604_
timestamp 0
transform 1 0 8270 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2605_
timestamp 0
transform -1 0 8150 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2606_
timestamp 0
transform -1 0 7750 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2607_
timestamp 0
transform -1 0 6610 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2608_
timestamp 0
transform 1 0 6790 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2609_
timestamp 0
transform 1 0 6990 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2610_
timestamp 0
transform -1 0 7930 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2611_
timestamp 0
transform -1 0 10150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2612_
timestamp 0
transform 1 0 9930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2613_
timestamp 0
transform 1 0 10330 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2614_
timestamp 0
transform -1 0 11030 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__2616_
timestamp 0
transform 1 0 8350 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2617_
timestamp 0
transform -1 0 7210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2618_
timestamp 0
transform -1 0 6550 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2619_
timestamp 0
transform 1 0 6330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2620_
timestamp 0
transform -1 0 8030 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2621_
timestamp 0
transform -1 0 8130 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2622_
timestamp 0
transform 1 0 8390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2623_
timestamp 0
transform -1 0 8990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2624_
timestamp 0
transform 1 0 8130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2625_
timestamp 0
transform 1 0 6890 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2626_
timestamp 0
transform -1 0 8350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2627_
timestamp 0
transform 1 0 9950 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2628_
timestamp 0
transform 1 0 11570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2629_
timestamp 0
transform 1 0 11470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2630_
timestamp 0
transform 1 0 11750 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2631_
timestamp 0
transform -1 0 11570 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2632_
timestamp 0
transform 1 0 9470 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2633_
timestamp 0
transform -1 0 8570 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2634_
timestamp 0
transform 1 0 8970 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2636_
timestamp 0
transform -1 0 9990 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2637_
timestamp 0
transform -1 0 8690 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2638_
timestamp 0
transform 1 0 9770 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2639_
timestamp 0
transform 1 0 10030 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2640_
timestamp 0
transform 1 0 8150 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2641_
timestamp 0
transform 1 0 7950 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2642_
timestamp 0
transform 1 0 9430 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2643_
timestamp 0
transform 1 0 9430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2644_
timestamp 0
transform 1 0 8450 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2645_
timestamp 0
transform 1 0 7670 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2646_
timestamp 0
transform 1 0 7470 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2647_
timestamp 0
transform 1 0 8250 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2648_
timestamp 0
transform -1 0 8090 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2649_
timestamp 0
transform -1 0 9090 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2650_
timestamp 0
transform 1 0 11150 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2651_
timestamp 0
transform -1 0 9290 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2652_
timestamp 0
transform -1 0 8590 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2653_
timestamp 0
transform 1 0 8770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2654_
timestamp 0
transform 1 0 5890 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2656_
timestamp 0
transform -1 0 6290 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2657_
timestamp 0
transform -1 0 7690 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2658_
timestamp 0
transform 1 0 7450 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2659_
timestamp 0
transform -1 0 7210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2660_
timestamp 0
transform -1 0 7390 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2661_
timestamp 0
transform -1 0 10830 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2662_
timestamp 0
transform 1 0 11010 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2663_
timestamp 0
transform 1 0 10070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2664_
timestamp 0
transform 1 0 10250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2665_
timestamp 0
transform -1 0 6670 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2666_
timestamp 0
transform 1 0 7250 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2667_
timestamp 0
transform -1 0 7050 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2668_
timestamp 0
transform -1 0 6870 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2669_
timestamp 0
transform 1 0 6790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2670_
timestamp 0
transform -1 0 10650 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2671_
timestamp 0
transform 1 0 11710 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2672_
timestamp 0
transform 1 0 11750 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2673_
timestamp 0
transform -1 0 11550 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2674_
timestamp 0
transform 1 0 11490 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2676_
timestamp 0
transform 1 0 11470 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2677_
timestamp 0
transform -1 0 11550 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2678_
timestamp 0
transform -1 0 10170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2679_
timestamp 0
transform 1 0 9770 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2680_
timestamp 0
transform 1 0 9690 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2681_
timestamp 0
transform 1 0 9370 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2682_
timestamp 0
transform -1 0 9590 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2683_
timestamp 0
transform -1 0 10250 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2684_
timestamp 0
transform -1 0 10550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2685_
timestamp 0
transform -1 0 10830 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__2686_
timestamp 0
transform 1 0 10730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2687_
timestamp 0
transform -1 0 9850 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2688_
timestamp 0
transform 1 0 9250 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2689_
timestamp 0
transform 1 0 10570 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2690_
timestamp 0
transform -1 0 10930 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2691_
timestamp 0
transform -1 0 11130 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2692_
timestamp 0
transform 1 0 11310 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2693_
timestamp 0
transform -1 0 10470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2694_
timestamp 0
transform 1 0 9670 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2696_
timestamp 0
transform 1 0 10350 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2697_
timestamp 0
transform 1 0 10010 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2698_
timestamp 0
transform 1 0 9990 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2699_
timestamp 0
transform 1 0 9110 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2700_
timestamp 0
transform 1 0 8890 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2701_
timestamp 0
transform -1 0 8530 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2702_
timestamp 0
transform 1 0 8890 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2703_
timestamp 0
transform 1 0 10910 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2704_
timestamp 0
transform -1 0 9170 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2705_
timestamp 0
transform -1 0 9730 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2706_
timestamp 0
transform -1 0 10130 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2707_
timestamp 0
transform -1 0 9650 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2708_
timestamp 0
transform 1 0 8950 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2709_
timestamp 0
transform 1 0 9070 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2710_
timestamp 0
transform -1 0 8770 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2711_
timestamp 0
transform -1 0 10830 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2712_
timestamp 0
transform -1 0 10810 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2713_
timestamp 0
transform 1 0 10850 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2714_
timestamp 0
transform 1 0 10850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2716_
timestamp 0
transform 1 0 11650 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2717_
timestamp 0
transform -1 0 10770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2718_
timestamp 0
transform 1 0 11110 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2719_
timestamp 0
transform 1 0 11830 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2720_
timestamp 0
transform -1 0 11030 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2721_
timestamp 0
transform -1 0 10930 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2722_
timestamp 0
transform -1 0 10970 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2723_
timestamp 0
transform 1 0 11410 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2724_
timestamp 0
transform 1 0 11390 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2725_
timestamp 0
transform 1 0 10370 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2726_
timestamp 0
transform -1 0 9750 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2727_
timestamp 0
transform 1 0 9950 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2728_
timestamp 0
transform -1 0 9930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2729_
timestamp 0
transform -1 0 9530 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2730_
timestamp 0
transform 1 0 11270 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2731_
timestamp 0
transform 1 0 9510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2732_
timestamp 0
transform 1 0 6730 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2733_
timestamp 0
transform -1 0 9150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2734_
timestamp 0
transform 1 0 9510 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2736_
timestamp 0
transform -1 0 8950 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2737_
timestamp 0
transform -1 0 9330 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2738_
timestamp 0
transform -1 0 10410 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2739_
timestamp 0
transform 1 0 10590 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2740_
timestamp 0
transform 1 0 11210 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2741_
timestamp 0
transform 1 0 11610 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2742_
timestamp 0
transform -1 0 10610 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2743_
timestamp 0
transform -1 0 10450 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2744_
timestamp 0
transform 1 0 10530 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2745_
timestamp 0
transform -1 0 11190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2746_
timestamp 0
transform -1 0 10190 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2747_
timestamp 0
transform 1 0 10990 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2748_
timestamp 0
transform 1 0 9850 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2749_
timestamp 0
transform 1 0 10710 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2750_
timestamp 0
transform 1 0 11050 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2751_
timestamp 0
transform -1 0 10170 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2752_
timestamp 0
transform 1 0 5790 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2753_
timestamp 0
transform -1 0 6010 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2754_
timestamp 0
transform -1 0 6070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2756_
timestamp 0
transform -1 0 7550 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2757_
timestamp 0
transform 1 0 8150 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2758_
timestamp 0
transform -1 0 7610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2759_
timestamp 0
transform -1 0 9750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2760_
timestamp 0
transform -1 0 6270 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2761_
timestamp 0
transform -1 0 8910 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2762_
timestamp 0
transform -1 0 8890 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2763_
timestamp 0
transform -1 0 6350 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2764_
timestamp 0
transform -1 0 6430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2765_
timestamp 0
transform -1 0 9390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2766_
timestamp 0
transform -1 0 6730 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2767_
timestamp 0
transform 1 0 8950 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2768_
timestamp 0
transform -1 0 6030 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2769_
timestamp 0
transform -1 0 6970 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2770_
timestamp 0
transform 1 0 7150 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2771_
timestamp 0
transform 1 0 10070 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2772_
timestamp 0
transform -1 0 7430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2773_
timestamp 0
transform -1 0 7630 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2774_
timestamp 0
transform -1 0 6070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2776_
timestamp 0
transform 1 0 6190 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2777_
timestamp 0
transform -1 0 9910 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2778_
timestamp 0
transform 1 0 7730 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2779_
timestamp 0
transform 1 0 7950 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2780_
timestamp 0
transform 1 0 8010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2781_
timestamp 0
transform -1 0 7830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2782_
timestamp 0
transform 1 0 7690 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2783_
timestamp 0
transform -1 0 8490 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2784_
timestamp 0
transform -1 0 11030 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2785_
timestamp 0
transform 1 0 9550 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2786_
timestamp 0
transform -1 0 7810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2787_
timestamp 0
transform -1 0 9250 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2788_
timestamp 0
transform -1 0 10230 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2789_
timestamp 0
transform 1 0 10410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2790_
timestamp 0
transform 1 0 8010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2791_
timestamp 0
transform 1 0 8210 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2792_
timestamp 0
transform -1 0 7670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2793_
timestamp 0
transform -1 0 7890 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2794_
timestamp 0
transform -1 0 7890 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2796_
timestamp 0
transform -1 0 7010 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2797_
timestamp 0
transform -1 0 8430 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2798_
timestamp 0
transform 1 0 11970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2799_
timestamp 0
transform -1 0 7390 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2800_
timestamp 0
transform -1 0 7510 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2801_
timestamp 0
transform 1 0 7150 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2802_
timestamp 0
transform 1 0 6810 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2803_
timestamp 0
transform -1 0 7030 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2804_
timestamp 0
transform -1 0 8530 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2805_
timestamp 0
transform 1 0 6950 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2806_
timestamp 0
transform -1 0 6850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2807_
timestamp 0
transform -1 0 7110 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2808_
timestamp 0
transform 1 0 10190 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2809_
timestamp 0
transform -1 0 10610 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2810_
timestamp 0
transform 1 0 10590 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2811_
timestamp 0
transform 1 0 10410 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2812_
timestamp 0
transform 1 0 10270 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2813_
timestamp 0
transform -1 0 10110 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2814_
timestamp 0
transform -1 0 10510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2816_
timestamp 0
transform 1 0 10230 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2817_
timestamp 0
transform -1 0 10330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2818_
timestamp 0
transform -1 0 10990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2819_
timestamp 0
transform -1 0 11090 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2820_
timestamp 0
transform -1 0 11290 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2821_
timestamp 0
transform 1 0 11050 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2822_
timestamp 0
transform -1 0 11990 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2823_
timestamp 0
transform 1 0 11170 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2824_
timestamp 0
transform 1 0 10670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2825_
timestamp 0
transform 1 0 11190 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2826_
timestamp 0
transform 1 0 11390 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2827_
timestamp 0
transform -1 0 11850 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2828_
timestamp 0
transform -1 0 11970 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2829_
timestamp 0
transform -1 0 11410 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2830_
timestamp 0
transform 1 0 11050 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2831_
timestamp 0
transform 1 0 11110 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2832_
timestamp 0
transform -1 0 11350 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2833_
timestamp 0
transform 1 0 11410 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2834_
timestamp 0
transform 1 0 11910 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2836_
timestamp 0
transform 1 0 11710 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2837_
timestamp 0
transform 1 0 11910 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2838_
timestamp 0
transform 1 0 12030 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2839_
timestamp 0
transform 1 0 11610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2840_
timestamp 0
transform -1 0 11810 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2841_
timestamp 0
transform -1 0 11670 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2842_
timestamp 0
transform -1 0 9850 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2843_
timestamp 0
transform -1 0 10050 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2844_
timestamp 0
transform -1 0 11830 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2845_
timestamp 0
transform 1 0 12010 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2846_
timestamp 0
transform 1 0 11570 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__2847_
timestamp 0
transform 1 0 11990 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2848_
timestamp 0
transform -1 0 11630 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2849_
timestamp 0
transform -1 0 11730 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2850_
timestamp 0
transform 1 0 11910 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2851_
timestamp 0
transform -1 0 9910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2852_
timestamp 0
transform -1 0 11090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2853_
timestamp 0
transform 1 0 11270 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2854_
timestamp 0
transform 1 0 11850 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2856_
timestamp 0
transform -1 0 9870 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2857_
timestamp 0
transform -1 0 9930 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2858_
timestamp 0
transform -1 0 8090 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2859_
timestamp 0
transform 1 0 9710 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2860_
timestamp 0
transform -1 0 9170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2861_
timestamp 0
transform 1 0 9990 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2862_
timestamp 0
transform 1 0 9590 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2863_
timestamp 0
transform 1 0 8810 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2864_
timestamp 0
transform -1 0 7810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2865_
timestamp 0
transform -1 0 6470 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2866_
timestamp 0
transform -1 0 8890 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2867_
timestamp 0
transform -1 0 9430 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2868_
timestamp 0
transform 1 0 9230 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2869_
timestamp 0
transform -1 0 10590 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2870_
timestamp 0
transform -1 0 9350 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2871_
timestamp 0
transform -1 0 8590 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2872_
timestamp 0
transform 1 0 9790 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2873_
timestamp 0
transform 1 0 9830 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2874_
timestamp 0
transform 1 0 9630 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2876_
timestamp 0
transform 1 0 10230 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2877_
timestamp 0
transform -1 0 10770 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2878_
timestamp 0
transform 1 0 9670 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2879_
timestamp 0
transform -1 0 9890 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2880_
timestamp 0
transform -1 0 10210 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2881_
timestamp 0
transform -1 0 5990 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2882_
timestamp 0
transform -1 0 6170 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2883_
timestamp 0
transform -1 0 5530 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2884_
timestamp 0
transform -1 0 5530 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2885_
timestamp 0
transform 1 0 5510 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2886_
timestamp 0
transform -1 0 5330 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__2887_
timestamp 0
transform 1 0 5670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2888_
timestamp 0
transform 1 0 6090 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2889_
timestamp 0
transform -1 0 6330 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2890_
timestamp 0
transform -1 0 6710 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2891_
timestamp 0
transform 1 0 8190 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2892_
timestamp 0
transform -1 0 7310 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2893_
timestamp 0
transform -1 0 5910 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2894_
timestamp 0
transform 1 0 5410 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2896_
timestamp 0
transform -1 0 6630 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__2897_
timestamp 0
transform 1 0 7370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2898_
timestamp 0
transform 1 0 11790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2899_
timestamp 0
transform -1 0 6570 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2900_
timestamp 0
transform -1 0 6770 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2901_
timestamp 0
transform -1 0 8210 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2902_
timestamp 0
transform 1 0 9670 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2903_
timestamp 0
transform -1 0 11610 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2904_
timestamp 0
transform 1 0 8390 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2905_
timestamp 0
transform -1 0 6970 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2906_
timestamp 0
transform -1 0 7350 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2907_
timestamp 0
transform -1 0 6370 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2908_
timestamp 0
transform 1 0 8490 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2909_
timestamp 0
transform -1 0 10390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2910_
timestamp 0
transform 1 0 10790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2911_
timestamp 0
transform 1 0 10970 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2912_
timestamp 0
transform -1 0 10830 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2913_
timestamp 0
transform -1 0 8710 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2914_
timestamp 0
transform -1 0 8590 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2916_
timestamp 0
transform -1 0 8010 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__2917_
timestamp 0
transform -1 0 7030 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2918_
timestamp 0
transform 1 0 6810 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2919_
timestamp 0
transform -1 0 7230 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2920_
timestamp 0
transform 1 0 7190 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2921_
timestamp 0
transform 1 0 6990 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2922_
timestamp 0
transform 1 0 6650 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2923_
timestamp 0
transform -1 0 5870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2924_
timestamp 0
transform 1 0 8910 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2925_
timestamp 0
transform 1 0 10270 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2926_
timestamp 0
transform 1 0 12010 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2927_
timestamp 0
transform 1 0 8730 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2928_
timestamp 0
transform 1 0 7530 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2929_
timestamp 0
transform 1 0 8250 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2930_
timestamp 0
transform -1 0 8470 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2931_
timestamp 0
transform -1 0 8110 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2932_
timestamp 0
transform 1 0 7910 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2933_
timestamp 0
transform 1 0 7950 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2934_
timestamp 0
transform -1 0 10250 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2936_
timestamp 0
transform -1 0 8230 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2937_
timestamp 0
transform 1 0 8710 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2938_
timestamp 0
transform -1 0 11830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2939_
timestamp 0
transform -1 0 11270 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2940_
timestamp 0
transform -1 0 6610 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2941_
timestamp 0
transform 1 0 8890 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2942_
timestamp 0
transform 1 0 8970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2943_
timestamp 0
transform 1 0 9730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2944_
timestamp 0
transform 1 0 9910 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__2945_
timestamp 0
transform 1 0 9090 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2946_
timestamp 0
transform -1 0 9190 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2947_
timestamp 0
transform -1 0 8750 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2948_
timestamp 0
transform -1 0 8690 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2949_
timestamp 0
transform 1 0 10870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__2950_
timestamp 0
transform 1 0 11690 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2951_
timestamp 0
transform -1 0 7010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2952_
timestamp 0
transform -1 0 6810 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2953_
timestamp 0
transform 1 0 11310 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2954_
timestamp 0
transform -1 0 8990 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2956_
timestamp 0
transform -1 0 11390 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2957_
timestamp 0
transform 1 0 9710 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2958_
timestamp 0
transform 1 0 11670 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__2959_
timestamp 0
transform 1 0 5150 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__2960_
timestamp 0
transform -1 0 7410 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2961_
timestamp 0
transform -1 0 8010 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2962_
timestamp 0
transform -1 0 7610 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2963_
timestamp 0
transform -1 0 6530 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__2964_
timestamp 0
transform -1 0 7810 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2965_
timestamp 0
transform -1 0 11790 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__2966_
timestamp 0
transform 1 0 8610 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2967_
timestamp 0
transform 1 0 9310 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__2968_
timestamp 0
transform 1 0 10430 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2969_
timestamp 0
transform 1 0 10630 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__2970_
timestamp 0
transform -1 0 11310 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2971_
timestamp 0
transform 1 0 7770 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2972_
timestamp 0
transform -1 0 9370 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2973_
timestamp 0
transform 1 0 7410 0 1 250
box -6 -8 26 248
use FILL  FILL_4__2974_
timestamp 0
transform -1 0 7350 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2976_
timestamp 0
transform 1 0 10090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2977_
timestamp 0
transform 1 0 10490 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2978_
timestamp 0
transform -1 0 11650 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__2979_
timestamp 0
transform -1 0 11890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__2980_
timestamp 0
transform 1 0 7210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2981_
timestamp 0
transform 1 0 6610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__2982_
timestamp 0
transform 1 0 7550 0 1 730
box -6 -8 26 248
use FILL  FILL_4__2983_
timestamp 0
transform 1 0 11930 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__2984_
timestamp 0
transform 1 0 11670 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__2985_
timestamp 0
transform -1 0 7170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__2986_
timestamp 0
transform -1 0 7190 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__2987_
timestamp 0
transform 1 0 5850 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__3000_
timestamp 0
transform -1 0 2250 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3001_
timestamp 0
transform 1 0 2390 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3002_
timestamp 0
transform 1 0 2190 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__3003_
timestamp 0
transform -1 0 3670 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__3004_
timestamp 0
transform 1 0 3870 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__3005_
timestamp 0
transform -1 0 3510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__3006_
timestamp 0
transform -1 0 4390 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__3007_
timestamp 0
transform -1 0 4190 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__3009_
timestamp 0
transform 1 0 4010 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3010_
timestamp 0
transform -1 0 4030 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__3011_
timestamp 0
transform 1 0 3830 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3012_
timestamp 0
transform 1 0 2770 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__3013_
timestamp 0
transform -1 0 2470 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3014_
timestamp 0
transform 1 0 2610 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__3015_
timestamp 0
transform -1 0 4590 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3016_
timestamp 0
transform 1 0 4510 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__3017_
timestamp 0
transform 1 0 4210 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3018_
timestamp 0
transform 1 0 4410 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3019_
timestamp 0
transform -1 0 4030 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3020_
timestamp 0
transform 1 0 1850 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3021_
timestamp 0
transform 1 0 1690 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3022_
timestamp 0
transform -1 0 2090 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3023_
timestamp 0
transform -1 0 2930 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3024_
timestamp 0
transform 1 0 4750 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3025_
timestamp 0
transform 1 0 4370 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3026_
timestamp 0
transform 1 0 3630 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3027_
timestamp 0
transform 1 0 3330 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__3029_
timestamp 0
transform 1 0 3470 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3030_
timestamp 0
transform 1 0 4910 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__3031_
timestamp 0
transform 1 0 4750 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__3032_
timestamp 0
transform 1 0 5910 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3033_
timestamp 0
transform -1 0 4630 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3034_
timestamp 0
transform 1 0 3850 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3035_
timestamp 0
transform -1 0 4610 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__3036_
timestamp 0
transform -1 0 2410 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__3037_
timestamp 0
transform -1 0 3350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__3038_
timestamp 0
transform 1 0 2230 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__3039_
timestamp 0
transform -1 0 3610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3040_
timestamp 0
transform -1 0 3830 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3041_
timestamp 0
transform 1 0 3430 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3042_
timestamp 0
transform -1 0 2810 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3043_
timestamp 0
transform -1 0 3850 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__3044_
timestamp 0
transform -1 0 2650 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3045_
timestamp 0
transform -1 0 2950 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__3046_
timestamp 0
transform -1 0 3290 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3047_
timestamp 0
transform 1 0 2890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3049_
timestamp 0
transform -1 0 3730 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__3050_
timestamp 0
transform -1 0 2970 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__3051_
timestamp 0
transform -1 0 2990 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__3052_
timestamp 0
transform 1 0 3150 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__3053_
timestamp 0
transform -1 0 3030 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3054_
timestamp 0
transform -1 0 2630 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__3055_
timestamp 0
transform -1 0 2450 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__3056_
timestamp 0
transform -1 0 2770 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3057_
timestamp 0
transform -1 0 3290 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3058_
timestamp 0
transform 1 0 4210 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3059_
timestamp 0
transform -1 0 5130 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__3060_
timestamp 0
transform -1 0 5330 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__3061_
timestamp 0
transform -1 0 6090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3062_
timestamp 0
transform -1 0 5150 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__3063_
timestamp 0
transform -1 0 5170 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__3064_
timestamp 0
transform -1 0 5010 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3076_
timestamp 0
transform 1 0 1110 0 1 250
box -6 -8 26 248
use FILL  FILL_4__3077_
timestamp 0
transform -1 0 1330 0 1 250
box -6 -8 26 248
use FILL  FILL_4__3078_
timestamp 0
transform 1 0 950 0 1 250
box -6 -8 26 248
use FILL  FILL_4__3080_
timestamp 0
transform -1 0 910 0 1 730
box -6 -8 26 248
use FILL  FILL_4__3081_
timestamp 0
transform 1 0 850 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__3082_
timestamp 0
transform 1 0 1430 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__3083_
timestamp 0
transform -1 0 1590 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__3084_
timestamp 0
transform 1 0 1510 0 1 250
box -6 -8 26 248
use FILL  FILL_4__3085_
timestamp 0
transform -1 0 1790 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__3086_
timestamp 0
transform -1 0 490 0 1 730
box -6 -8 26 248
use FILL  FILL_4__3087_
timestamp 0
transform -1 0 670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__3088_
timestamp 0
transform 1 0 470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__3089_
timestamp 0
transform -1 0 1450 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__3090_
timestamp 0
transform 1 0 1250 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3091_
timestamp 0
transform -1 0 1930 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__3092_
timestamp 0
transform -1 0 710 0 1 730
box -6 -8 26 248
use FILL  FILL_4__3093_
timestamp 0
transform -1 0 110 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__3094_
timestamp 0
transform -1 0 110 0 1 730
box -6 -8 26 248
use FILL  FILL_4__3095_
timestamp 0
transform -1 0 310 0 1 730
box -6 -8 26 248
use FILL  FILL_4__3096_
timestamp 0
transform -1 0 310 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__3097_
timestamp 0
transform 1 0 2070 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__3098_
timestamp 0
transform -1 0 2370 0 1 250
box -6 -8 26 248
use FILL  FILL_4__3100_
timestamp 0
transform 1 0 90 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3101_
timestamp 0
transform -1 0 110 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__3102_
timestamp 0
transform -1 0 1290 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__3103_
timestamp 0
transform -1 0 1250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__3104_
timestamp 0
transform -1 0 290 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__3105_
timestamp 0
transform -1 0 1210 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__3106_
timestamp 0
transform -1 0 2370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__3107_
timestamp 0
transform -1 0 1570 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__3108_
timestamp 0
transform -1 0 450 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3109_
timestamp 0
transform -1 0 630 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3110_
timestamp 0
transform 1 0 770 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__3111_
timestamp 0
transform -1 0 970 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__3112_
timestamp 0
transform -1 0 110 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__3113_
timestamp 0
transform -1 0 110 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3114_
timestamp 0
transform -1 0 4610 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__3115_
timestamp 0
transform -1 0 4670 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3116_
timestamp 0
transform 1 0 4530 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__3117_
timestamp 0
transform 1 0 570 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__3118_
timestamp 0
transform -1 0 1730 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__3120_
timestamp 0
transform 1 0 1070 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3121_
timestamp 0
transform -1 0 2390 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3122_
timestamp 0
transform -1 0 490 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__3123_
timestamp 0
transform 1 0 370 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__3124_
timestamp 0
transform 1 0 270 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__3125_
timestamp 0
transform 1 0 2090 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__3126_
timestamp 0
transform -1 0 2310 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__3127_
timestamp 0
transform 1 0 1610 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3128_
timestamp 0
transform 1 0 1450 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3129_
timestamp 0
transform 1 0 4790 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__3130_
timestamp 0
transform 1 0 4970 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__3131_
timestamp 0
transform 1 0 5190 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__3132_
timestamp 0
transform 1 0 4850 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3133_
timestamp 0
transform -1 0 4750 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__3134_
timestamp 0
transform -1 0 4390 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__3135_
timestamp 0
transform 1 0 750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__3136_
timestamp 0
transform -1 0 810 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__3137_
timestamp 0
transform 1 0 410 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__3138_
timestamp 0
transform 1 0 750 0 1 250
box -6 -8 26 248
use FILL  FILL_4__3140_
timestamp 0
transform -1 0 1570 0 1 730
box -6 -8 26 248
use FILL  FILL_4__3141_
timestamp 0
transform 1 0 1750 0 1 730
box -6 -8 26 248
use FILL  FILL_4__3142_
timestamp 0
transform -1 0 1730 0 1 250
box -6 -8 26 248
use FILL  FILL_4__3143_
timestamp 0
transform 1 0 2430 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__3144_
timestamp 0
transform 1 0 2550 0 1 250
box -6 -8 26 248
use FILL  FILL_4__3145_
timestamp 0
transform 1 0 2270 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__3146_
timestamp 0
transform -1 0 1970 0 1 730
box -6 -8 26 248
use FILL  FILL_4__3147_
timestamp 0
transform 1 0 2070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__3148_
timestamp 0
transform 1 0 1110 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__3149_
timestamp 0
transform -1 0 950 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__3150_
timestamp 0
transform -1 0 310 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__3151_
timestamp 0
transform 1 0 90 0 1 250
box -6 -8 26 248
use FILL  FILL_4__3152_
timestamp 0
transform -1 0 2170 0 1 730
box -6 -8 26 248
use FILL  FILL_4__3284_
timestamp 0
transform -1 0 4770 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__3285_
timestamp 0
transform 1 0 4410 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__3286_
timestamp 0
transform -1 0 3450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3287_
timestamp 0
transform 1 0 3310 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3288_
timestamp 0
transform 1 0 2230 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3289_
timestamp 0
transform 1 0 2430 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3291_
timestamp 0
transform 1 0 3050 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3292_
timestamp 0
transform 1 0 3250 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3293_
timestamp 0
transform 1 0 5870 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3294_
timestamp 0
transform -1 0 5910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3295_
timestamp 0
transform 1 0 5950 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3296_
timestamp 0
transform 1 0 6430 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3297_
timestamp 0
transform 1 0 6630 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3298_
timestamp 0
transform 1 0 5330 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3299_
timestamp 0
transform 1 0 5530 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3300_
timestamp 0
transform 1 0 4670 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3301_
timestamp 0
transform 1 0 4870 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3302_
timestamp 0
transform -1 0 3430 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3303_
timestamp 0
transform -1 0 3590 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3304_
timestamp 0
transform -1 0 3470 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3305_
timestamp 0
transform -1 0 3650 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3306_
timestamp 0
transform 1 0 4390 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3307_
timestamp 0
transform 1 0 4490 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3308_
timestamp 0
transform -1 0 1150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3309_
timestamp 0
transform -1 0 1070 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__3311_
timestamp 0
transform -1 0 2770 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3312_
timestamp 0
transform 1 0 3490 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3313_
timestamp 0
transform -1 0 2410 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3314_
timestamp 0
transform -1 0 290 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__3315_
timestamp 0
transform -1 0 490 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__3316_
timestamp 0
transform -1 0 7570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__3317_
timestamp 0
transform 1 0 6190 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3318_
timestamp 0
transform 1 0 2670 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3319_
timestamp 0
transform 1 0 6690 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3320_
timestamp 0
transform 1 0 5470 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3321_
timestamp 0
transform -1 0 6490 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__3322_
timestamp 0
transform -1 0 3850 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__3323_
timestamp 0
transform -1 0 3690 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3324_
timestamp 0
transform 1 0 5190 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__3325_
timestamp 0
transform -1 0 5410 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__3326_
timestamp 0
transform -1 0 5270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__3327_
timestamp 0
transform 1 0 4850 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__3328_
timestamp 0
transform -1 0 5310 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3329_
timestamp 0
transform -1 0 5730 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__3331_
timestamp 0
transform 1 0 5010 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__3332_
timestamp 0
transform -1 0 4690 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__3333_
timestamp 0
transform -1 0 5990 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__3334_
timestamp 0
transform 1 0 5970 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__3335_
timestamp 0
transform -1 0 490 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3336_
timestamp 0
transform -1 0 310 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3337_
timestamp 0
transform -1 0 930 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3338_
timestamp 0
transform -1 0 950 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3339_
timestamp 0
transform -1 0 5910 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__3340_
timestamp 0
transform 1 0 6090 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__3341_
timestamp 0
transform -1 0 5870 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3342_
timestamp 0
transform -1 0 5490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3343_
timestamp 0
transform -1 0 4410 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3344_
timestamp 0
transform -1 0 5530 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__3345_
timestamp 0
transform 1 0 5710 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__3346_
timestamp 0
transform 1 0 5310 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__3347_
timestamp 0
transform 1 0 5130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__3348_
timestamp 0
transform -1 0 110 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3349_
timestamp 0
transform 1 0 290 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3351_
timestamp 0
transform -1 0 110 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3352_
timestamp 0
transform 1 0 330 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3353_
timestamp 0
transform -1 0 1850 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3354_
timestamp 0
transform 1 0 2030 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3355_
timestamp 0
transform -1 0 350 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3356_
timestamp 0
transform -1 0 550 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3357_
timestamp 0
transform -1 0 890 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3358_
timestamp 0
transform -1 0 870 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3359_
timestamp 0
transform -1 0 110 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3360_
timestamp 0
transform -1 0 310 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__3361_
timestamp 0
transform -1 0 4910 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3362_
timestamp 0
transform -1 0 5030 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3363_
timestamp 0
transform 1 0 5350 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3364_
timestamp 0
transform -1 0 3450 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3365_
timestamp 0
transform 1 0 3370 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3366_
timestamp 0
transform 1 0 2950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3367_
timestamp 0
transform 1 0 2590 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3368_
timestamp 0
transform 1 0 2390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3369_
timestamp 0
transform -1 0 4170 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3371_
timestamp 0
transform -1 0 7090 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3372_
timestamp 0
transform 1 0 5130 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3373_
timestamp 0
transform -1 0 7530 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3374_
timestamp 0
transform -1 0 7310 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3375_
timestamp 0
transform -1 0 4710 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3376_
timestamp 0
transform -1 0 4750 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3377_
timestamp 0
transform 1 0 4930 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3378_
timestamp 0
transform -1 0 4350 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3379_
timestamp 0
transform 1 0 5790 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3380_
timestamp 0
transform -1 0 7850 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3381_
timestamp 0
transform 1 0 6690 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3382_
timestamp 0
transform 1 0 6510 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3383_
timestamp 0
transform -1 0 7110 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3384_
timestamp 0
transform -1 0 6910 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3385_
timestamp 0
transform 1 0 7290 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3386_
timestamp 0
transform -1 0 6550 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3387_
timestamp 0
transform 1 0 6330 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3388_
timestamp 0
transform 1 0 6750 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3389_
timestamp 0
transform -1 0 7150 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3391_
timestamp 0
transform -1 0 10290 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3392_
timestamp 0
transform -1 0 290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3393_
timestamp 0
transform 1 0 270 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3394_
timestamp 0
transform -1 0 270 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3395_
timestamp 0
transform -1 0 290 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3396_
timestamp 0
transform -1 0 110 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3397_
timestamp 0
transform -1 0 1270 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3398_
timestamp 0
transform 1 0 1050 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3399_
timestamp 0
transform 1 0 1010 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3400_
timestamp 0
transform -1 0 650 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3401_
timestamp 0
transform -1 0 110 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__3402_
timestamp 0
transform -1 0 870 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3403_
timestamp 0
transform 1 0 1630 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3404_
timestamp 0
transform -1 0 930 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3405_
timestamp 0
transform 1 0 730 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3406_
timestamp 0
transform -1 0 1910 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3407_
timestamp 0
transform -1 0 510 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__3408_
timestamp 0
transform 1 0 290 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__3409_
timestamp 0
transform -1 0 110 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__3411_
timestamp 0
transform -1 0 470 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3412_
timestamp 0
transform -1 0 290 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3413_
timestamp 0
transform -1 0 110 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3414_
timestamp 0
transform -1 0 270 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3415_
timestamp 0
transform -1 0 110 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3416_
timestamp 0
transform -1 0 110 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3417_
timestamp 0
transform -1 0 450 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3418_
timestamp 0
transform -1 0 6970 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3419_
timestamp 0
transform 1 0 6270 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3420_
timestamp 0
transform 1 0 6070 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3421_
timestamp 0
transform 1 0 5310 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3422_
timestamp 0
transform 1 0 5170 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3423_
timestamp 0
transform 1 0 7150 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3424_
timestamp 0
transform -1 0 1410 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3425_
timestamp 0
transform 1 0 650 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3426_
timestamp 0
transform 1 0 450 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3427_
timestamp 0
transform -1 0 470 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3428_
timestamp 0
transform -1 0 310 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3429_
timestamp 0
transform 1 0 630 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3431_
timestamp 0
transform -1 0 290 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3432_
timestamp 0
transform 1 0 910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3433_
timestamp 0
transform 1 0 1510 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3434_
timestamp 0
transform -1 0 1010 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3435_
timestamp 0
transform -1 0 1130 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3436_
timestamp 0
transform 1 0 1310 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3437_
timestamp 0
transform -1 0 1350 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__3438_
timestamp 0
transform -1 0 1030 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3439_
timestamp 0
transform -1 0 830 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3440_
timestamp 0
transform -1 0 1150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__3441_
timestamp 0
transform 1 0 750 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3442_
timestamp 0
transform 1 0 850 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3443_
timestamp 0
transform -1 0 830 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3444_
timestamp 0
transform -1 0 650 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3445_
timestamp 0
transform -1 0 770 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__3446_
timestamp 0
transform -1 0 1430 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3447_
timestamp 0
transform -1 0 1210 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3448_
timestamp 0
transform -1 0 750 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3449_
timestamp 0
transform 1 0 1370 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3451_
timestamp 0
transform -1 0 2670 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3452_
timestamp 0
transform -1 0 2870 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3453_
timestamp 0
transform -1 0 3090 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3454_
timestamp 0
transform -1 0 1210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__3455_
timestamp 0
transform -1 0 310 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3456_
timestamp 0
transform -1 0 110 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3457_
timestamp 0
transform -1 0 870 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3458_
timestamp 0
transform 1 0 650 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3459_
timestamp 0
transform -1 0 590 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__3460_
timestamp 0
transform 1 0 490 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3461_
timestamp 0
transform -1 0 1930 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3462_
timestamp 0
transform 1 0 1710 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3463_
timestamp 0
transform -1 0 1970 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__3464_
timestamp 0
transform -1 0 2090 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3465_
timestamp 0
transform -1 0 1670 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__3466_
timestamp 0
transform -1 0 2050 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__3467_
timestamp 0
transform -1 0 1910 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3468_
timestamp 0
transform -1 0 2310 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3469_
timestamp 0
transform -1 0 310 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__3471_
timestamp 0
transform -1 0 1230 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3472_
timestamp 0
transform -1 0 1610 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3473_
timestamp 0
transform 1 0 1790 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3474_
timestamp 0
transform -1 0 2090 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3475_
timestamp 0
transform -1 0 1770 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3476_
timestamp 0
transform -1 0 1730 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3477_
timestamp 0
transform -1 0 1910 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3478_
timestamp 0
transform 1 0 1990 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3479_
timestamp 0
transform -1 0 1450 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3480_
timestamp 0
transform -1 0 2850 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3481_
timestamp 0
transform -1 0 6090 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3482_
timestamp 0
transform -1 0 5910 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3483_
timestamp 0
transform 1 0 6750 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3484_
timestamp 0
transform -1 0 7510 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__3485_
timestamp 0
transform -1 0 7310 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__3486_
timestamp 0
transform 1 0 5770 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__3487_
timestamp 0
transform -1 0 5790 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__3488_
timestamp 0
transform 1 0 3010 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3489_
timestamp 0
transform -1 0 6150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__3491_
timestamp 0
transform 1 0 1390 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3492_
timestamp 0
transform 1 0 1950 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3493_
timestamp 0
transform -1 0 1790 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3494_
timestamp 0
transform 1 0 7230 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3495_
timestamp 0
transform -1 0 7610 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3496_
timestamp 0
transform -1 0 7810 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3497_
timestamp 0
transform -1 0 8230 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3498_
timestamp 0
transform -1 0 7450 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3499_
timestamp 0
transform 1 0 1190 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__3500_
timestamp 0
transform 1 0 1390 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__3501_
timestamp 0
transform -1 0 3170 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3502_
timestamp 0
transform -1 0 3770 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3503_
timestamp 0
transform -1 0 3270 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3504_
timestamp 0
transform 1 0 2970 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__3505_
timestamp 0
transform 1 0 3170 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__3506_
timestamp 0
transform -1 0 790 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__3507_
timestamp 0
transform -1 0 990 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__3508_
timestamp 0
transform 1 0 6390 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__3509_
timestamp 0
transform -1 0 6630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__3511_
timestamp 0
transform -1 0 6670 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__3512_
timestamp 0
transform 1 0 6610 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__3513_
timestamp 0
transform 1 0 6790 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__3514_
timestamp 0
transform -1 0 6530 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3515_
timestamp 0
transform 1 0 7190 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__3516_
timestamp 0
transform -1 0 1250 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3517_
timestamp 0
transform 1 0 1030 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3518_
timestamp 0
transform -1 0 7510 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3519_
timestamp 0
transform -1 0 7330 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3520_
timestamp 0
transform 1 0 5350 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3521_
timestamp 0
transform -1 0 5550 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3522_
timestamp 0
transform -1 0 110 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__3523_
timestamp 0
transform 1 0 270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3524_
timestamp 0
transform -1 0 490 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__3525_
timestamp 0
transform 1 0 2070 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__3526_
timestamp 0
transform 1 0 2250 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__3527_
timestamp 0
transform 1 0 7050 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__3528_
timestamp 0
transform -1 0 6990 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__3529_
timestamp 0
transform -1 0 110 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3531_
timestamp 0
transform 1 0 6090 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3532_
timestamp 0
transform 1 0 5710 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3533_
timestamp 0
transform 1 0 11870 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3534_
timestamp 0
transform -1 0 9170 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3535_
timestamp 0
transform 1 0 7670 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3536_
timestamp 0
transform 1 0 6070 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__3537_
timestamp 0
transform 1 0 5610 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3538_
timestamp 0
transform 1 0 5590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__3539_
timestamp 0
transform 1 0 6190 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__3540_
timestamp 0
transform 1 0 6390 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__3541_
timestamp 0
transform -1 0 6270 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3542_
timestamp 0
transform -1 0 6090 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3543_
timestamp 0
transform 1 0 5990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__3544_
timestamp 0
transform 1 0 5870 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3545_
timestamp 0
transform 1 0 5870 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3546_
timestamp 0
transform -1 0 6250 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__3547_
timestamp 0
transform 1 0 6410 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__3548_
timestamp 0
transform 1 0 6510 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3549_
timestamp 0
transform 1 0 6710 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3551_
timestamp 0
transform -1 0 6770 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3552_
timestamp 0
transform 1 0 6850 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3553_
timestamp 0
transform -1 0 7290 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__3554_
timestamp 0
transform 1 0 11250 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3555_
timestamp 0
transform 1 0 10910 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3556_
timestamp 0
transform 1 0 10170 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3557_
timestamp 0
transform -1 0 9250 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3558_
timestamp 0
transform -1 0 10750 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3559_
timestamp 0
transform 1 0 11590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3560_
timestamp 0
transform 1 0 10050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3561_
timestamp 0
transform 1 0 10030 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3562_
timestamp 0
transform 1 0 9830 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3563_
timestamp 0
transform -1 0 9910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3564_
timestamp 0
transform -1 0 11850 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3565_
timestamp 0
transform 1 0 12030 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3566_
timestamp 0
transform 1 0 11450 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3567_
timestamp 0
transform 1 0 11090 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3568_
timestamp 0
transform 1 0 11230 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3569_
timestamp 0
transform 1 0 9770 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3571_
timestamp 0
transform 1 0 9590 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3572_
timestamp 0
transform -1 0 9430 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3573_
timestamp 0
transform 1 0 11030 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3574_
timestamp 0
transform -1 0 9370 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3575_
timestamp 0
transform 1 0 8570 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3576_
timestamp 0
transform -1 0 8050 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3577_
timestamp 0
transform -1 0 9030 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3578_
timestamp 0
transform -1 0 9110 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3579_
timestamp 0
transform -1 0 8230 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3580_
timestamp 0
transform -1 0 8690 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3581_
timestamp 0
transform 1 0 9630 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3582_
timestamp 0
transform 1 0 9430 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3583_
timestamp 0
transform 1 0 8490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3584_
timestamp 0
transform -1 0 8430 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3585_
timestamp 0
transform 1 0 9150 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3586_
timestamp 0
transform -1 0 8990 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3587_
timestamp 0
transform -1 0 9230 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3588_
timestamp 0
transform 1 0 8230 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3589_
timestamp 0
transform -1 0 9050 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3591_
timestamp 0
transform -1 0 10790 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3592_
timestamp 0
transform 1 0 8250 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3593_
timestamp 0
transform -1 0 6230 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3594_
timestamp 0
transform -1 0 10390 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3595_
timestamp 0
transform -1 0 10550 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3596_
timestamp 0
transform 1 0 6990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3597_
timestamp 0
transform 1 0 6650 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3598_
timestamp 0
transform 1 0 11870 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3599_
timestamp 0
transform -1 0 8930 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3600_
timestamp 0
transform 1 0 8710 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3601_
timestamp 0
transform 1 0 8850 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3602_
timestamp 0
transform -1 0 9970 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3603_
timestamp 0
transform -1 0 10290 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3604_
timestamp 0
transform -1 0 8450 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3605_
timestamp 0
transform -1 0 7890 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3606_
timestamp 0
transform -1 0 8030 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3607_
timestamp 0
transform 1 0 7830 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3608_
timestamp 0
transform 1 0 11430 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3609_
timestamp 0
transform 1 0 11650 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3611_
timestamp 0
transform 1 0 11310 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3612_
timestamp 0
transform 1 0 11670 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3613_
timestamp 0
transform 1 0 11410 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3614_
timestamp 0
transform 1 0 11610 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3615_
timestamp 0
transform 1 0 11350 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3616_
timestamp 0
transform -1 0 8130 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3617_
timestamp 0
transform 1 0 12050 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3618_
timestamp 0
transform 1 0 11990 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3619_
timestamp 0
transform -1 0 11570 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3620_
timestamp 0
transform 1 0 8810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3621_
timestamp 0
transform 1 0 8190 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3622_
timestamp 0
transform 1 0 8150 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3623_
timestamp 0
transform 1 0 11150 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3624_
timestamp 0
transform -1 0 11130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3625_
timestamp 0
transform 1 0 10810 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3626_
timestamp 0
transform 1 0 11010 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3627_
timestamp 0
transform 1 0 10950 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3628_
timestamp 0
transform 1 0 7990 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3629_
timestamp 0
transform 1 0 7650 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3631_
timestamp 0
transform -1 0 7490 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3632_
timestamp 0
transform 1 0 7050 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3633_
timestamp 0
transform 1 0 8050 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3634_
timestamp 0
transform 1 0 8730 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3635_
timestamp 0
transform 1 0 8390 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3636_
timestamp 0
transform -1 0 6870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3637_
timestamp 0
transform 1 0 8750 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3638_
timestamp 0
transform 1 0 10850 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3639_
timestamp 0
transform 1 0 8610 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3640_
timestamp 0
transform 1 0 9470 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3641_
timestamp 0
transform 1 0 8970 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3642_
timestamp 0
transform -1 0 7330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3643_
timestamp 0
transform 1 0 7130 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3644_
timestamp 0
transform -1 0 9350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3645_
timestamp 0
transform -1 0 10430 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3646_
timestamp 0
transform 1 0 9130 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3647_
timestamp 0
transform 1 0 10570 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3648_
timestamp 0
transform 1 0 10890 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3649_
timestamp 0
transform 1 0 10990 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3651_
timestamp 0
transform 1 0 6790 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3652_
timestamp 0
transform 1 0 4850 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3653_
timestamp 0
transform 1 0 4650 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3654_
timestamp 0
transform 1 0 4450 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3655_
timestamp 0
transform 1 0 4250 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3656_
timestamp 0
transform 1 0 5450 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3657_
timestamp 0
transform 1 0 5410 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3658_
timestamp 0
transform 1 0 5250 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3659_
timestamp 0
transform 1 0 4670 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3660_
timestamp 0
transform 1 0 4470 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3661_
timestamp 0
transform 1 0 4850 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3662_
timestamp 0
transform 1 0 6590 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3663_
timestamp 0
transform 1 0 6390 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3664_
timestamp 0
transform 1 0 5630 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3665_
timestamp 0
transform 1 0 5230 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3666_
timestamp 0
transform 1 0 5830 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3667_
timestamp 0
transform -1 0 3710 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3668_
timestamp 0
transform 1 0 3930 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3669_
timestamp 0
transform -1 0 3430 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3671_
timestamp 0
transform 1 0 4190 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3672_
timestamp 0
transform 1 0 4250 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3673_
timestamp 0
transform 1 0 6010 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3674_
timestamp 0
transform -1 0 10750 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3675_
timestamp 0
transform -1 0 10570 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3676_
timestamp 0
transform 1 0 4170 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__3677_
timestamp 0
transform -1 0 4230 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__3678_
timestamp 0
transform 1 0 4670 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3679_
timestamp 0
transform -1 0 4890 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3680_
timestamp 0
transform -1 0 5090 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3681_
timestamp 0
transform -1 0 4790 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3682_
timestamp 0
transform 1 0 1670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__3683_
timestamp 0
transform 1 0 6290 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3684_
timestamp 0
transform 1 0 6630 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3685_
timestamp 0
transform 1 0 6910 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3686_
timestamp 0
transform 1 0 6690 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3687_
timestamp 0
transform 1 0 4910 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3688_
timestamp 0
transform -1 0 4930 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3689_
timestamp 0
transform 1 0 5110 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3691_
timestamp 0
transform -1 0 4710 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3692_
timestamp 0
transform 1 0 4510 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3693_
timestamp 0
transform 1 0 4890 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3694_
timestamp 0
transform -1 0 6090 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3695_
timestamp 0
transform 1 0 1730 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3696_
timestamp 0
transform 1 0 7610 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3697_
timestamp 0
transform 1 0 7810 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3698_
timestamp 0
transform 1 0 6710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3699_
timestamp 0
transform 1 0 6910 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3700_
timestamp 0
transform -1 0 7110 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3701_
timestamp 0
transform 1 0 4670 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__3702_
timestamp 0
transform 1 0 4370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__3703_
timestamp 0
transform 1 0 4430 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3704_
timestamp 0
transform 1 0 4850 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3705_
timestamp 0
transform -1 0 4930 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3706_
timestamp 0
transform -1 0 4710 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__3707_
timestamp 0
transform -1 0 5050 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3708_
timestamp 0
transform 1 0 4630 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3709_
timestamp 0
transform 1 0 2490 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3711_
timestamp 0
transform 1 0 9690 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3712_
timestamp 0
transform 1 0 9670 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3713_
timestamp 0
transform 1 0 10050 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3714_
timestamp 0
transform 1 0 8750 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3715_
timestamp 0
transform -1 0 8950 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3716_
timestamp 0
transform -1 0 9550 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3717_
timestamp 0
transform -1 0 10450 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3718_
timestamp 0
transform 1 0 10610 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3719_
timestamp 0
transform -1 0 9150 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3720_
timestamp 0
transform 1 0 9330 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3721_
timestamp 0
transform -1 0 10670 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3722_
timestamp 0
transform -1 0 10490 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3723_
timestamp 0
transform 1 0 10810 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3724_
timestamp 0
transform 1 0 9490 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3725_
timestamp 0
transform 1 0 8350 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3726_
timestamp 0
transform -1 0 8230 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3727_
timestamp 0
transform 1 0 9670 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3728_
timestamp 0
transform -1 0 10230 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3729_
timestamp 0
transform 1 0 10070 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3731_
timestamp 0
transform 1 0 8470 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3732_
timestamp 0
transform 1 0 8850 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3733_
timestamp 0
transform -1 0 3910 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3734_
timestamp 0
transform -1 0 4090 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3735_
timestamp 0
transform 1 0 7670 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3736_
timestamp 0
transform -1 0 7270 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3737_
timestamp 0
transform -1 0 5830 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3738_
timestamp 0
transform 1 0 9610 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3739_
timestamp 0
transform 1 0 9410 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3740_
timestamp 0
transform 1 0 9290 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3741_
timestamp 0
transform -1 0 10790 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3742_
timestamp 0
transform 1 0 11290 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3743_
timestamp 0
transform 1 0 11470 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3744_
timestamp 0
transform 1 0 11210 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3745_
timestamp 0
transform -1 0 10630 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3746_
timestamp 0
transform -1 0 10290 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3747_
timestamp 0
transform -1 0 10230 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3748_
timestamp 0
transform -1 0 10970 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3749_
timestamp 0
transform -1 0 11290 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3751_
timestamp 0
transform -1 0 8090 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3752_
timestamp 0
transform -1 0 6890 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3753_
timestamp 0
transform -1 0 6790 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3754_
timestamp 0
transform 1 0 4430 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3755_
timestamp 0
transform 1 0 3070 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3756_
timestamp 0
transform 1 0 4110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3757_
timestamp 0
transform 1 0 4590 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3758_
timestamp 0
transform -1 0 5110 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__3759_
timestamp 0
transform -1 0 4890 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__3760_
timestamp 0
transform -1 0 4330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3761_
timestamp 0
transform -1 0 4350 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__3762_
timestamp 0
transform -1 0 4450 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__3763_
timestamp 0
transform -1 0 4190 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3764_
timestamp 0
transform -1 0 3470 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3765_
timestamp 0
transform -1 0 4650 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__3766_
timestamp 0
transform 1 0 2270 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__3767_
timestamp 0
transform -1 0 2490 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__3768_
timestamp 0
transform -1 0 2650 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__3769_
timestamp 0
transform -1 0 2850 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__3771_
timestamp 0
transform 1 0 3430 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__3772_
timestamp 0
transform -1 0 1070 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3773_
timestamp 0
transform 1 0 5850 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__3774_
timestamp 0
transform 1 0 5070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__3775_
timestamp 0
transform -1 0 5030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3776_
timestamp 0
transform -1 0 4870 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3777_
timestamp 0
transform 1 0 4930 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3778_
timestamp 0
transform 1 0 4770 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3779_
timestamp 0
transform 1 0 4570 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3780_
timestamp 0
transform 1 0 5250 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3781_
timestamp 0
transform -1 0 5430 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3782_
timestamp 0
transform -1 0 4410 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3783_
timestamp 0
transform 1 0 3850 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3784_
timestamp 0
transform -1 0 5290 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3785_
timestamp 0
transform 1 0 7570 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__3786_
timestamp 0
transform 1 0 7430 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__3787_
timestamp 0
transform -1 0 7410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3788_
timestamp 0
transform -1 0 7250 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3789_
timestamp 0
transform -1 0 7270 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__3791_
timestamp 0
transform -1 0 6630 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__3792_
timestamp 0
transform 1 0 7050 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__3793_
timestamp 0
transform -1 0 6850 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__3794_
timestamp 0
transform 1 0 8010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__3795_
timestamp 0
transform -1 0 9630 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3796_
timestamp 0
transform 1 0 8330 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3797_
timestamp 0
transform 1 0 7710 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3798_
timestamp 0
transform 1 0 6990 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3799_
timestamp 0
transform -1 0 7170 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3800_
timestamp 0
transform -1 0 7350 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3801_
timestamp 0
transform 1 0 5690 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3802_
timestamp 0
transform -1 0 5950 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3803_
timestamp 0
transform 1 0 5730 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3804_
timestamp 0
transform 1 0 5350 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3805_
timestamp 0
transform 1 0 5390 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3806_
timestamp 0
transform 1 0 5070 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3807_
timestamp 0
transform -1 0 5550 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3808_
timestamp 0
transform -1 0 7930 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3809_
timestamp 0
transform -1 0 8050 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3811_
timestamp 0
transform -1 0 7530 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3812_
timestamp 0
transform 1 0 10470 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3813_
timestamp 0
transform -1 0 9890 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3814_
timestamp 0
transform 1 0 9870 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3815_
timestamp 0
transform -1 0 9870 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3816_
timestamp 0
transform -1 0 9710 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3817_
timestamp 0
transform 1 0 9170 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3818_
timestamp 0
transform -1 0 8990 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3819_
timestamp 0
transform 1 0 10170 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3820_
timestamp 0
transform 1 0 10250 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3821_
timestamp 0
transform 1 0 6570 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3822_
timestamp 0
transform -1 0 3370 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3823_
timestamp 0
transform -1 0 8290 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3824_
timestamp 0
transform 1 0 7310 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3825_
timestamp 0
transform -1 0 10010 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3826_
timestamp 0
transform 1 0 9490 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3827_
timestamp 0
transform -1 0 9330 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3828_
timestamp 0
transform 1 0 9130 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3829_
timestamp 0
transform 1 0 8930 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3830_
timestamp 0
transform 1 0 7430 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3832_
timestamp 0
transform 1 0 8570 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3833_
timestamp 0
transform 1 0 8750 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3834_
timestamp 0
transform -1 0 8730 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3835_
timestamp 0
transform 1 0 8930 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3836_
timestamp 0
transform 1 0 9230 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3837_
timestamp 0
transform -1 0 8490 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3838_
timestamp 0
transform 1 0 8670 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3839_
timestamp 0
transform 1 0 8910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3840_
timestamp 0
transform -1 0 8550 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3841_
timestamp 0
transform -1 0 8350 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3842_
timestamp 0
transform 1 0 9110 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3843_
timestamp 0
transform -1 0 8370 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3844_
timestamp 0
transform 1 0 7670 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3845_
timestamp 0
transform 1 0 9330 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__3846_
timestamp 0
transform 1 0 8890 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3847_
timestamp 0
transform 1 0 8170 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3848_
timestamp 0
transform -1 0 8030 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__3849_
timestamp 0
transform 1 0 7810 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__3850_
timestamp 0
transform 1 0 7990 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3852_
timestamp 0
transform -1 0 7850 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3853_
timestamp 0
transform -1 0 7610 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3854_
timestamp 0
transform -1 0 7470 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3855_
timestamp 0
transform 1 0 7850 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__3856_
timestamp 0
transform -1 0 7250 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3857_
timestamp 0
transform -1 0 8350 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3858_
timestamp 0
transform 1 0 8690 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3859_
timestamp 0
transform 1 0 7870 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3860_
timestamp 0
transform 1 0 4810 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3861_
timestamp 0
transform 1 0 8550 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3862_
timestamp 0
transform -1 0 8790 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3863_
timestamp 0
transform -1 0 10250 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3864_
timestamp 0
transform 1 0 9490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3865_
timestamp 0
transform 1 0 8070 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3866_
timestamp 0
transform 1 0 5670 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3867_
timestamp 0
transform -1 0 7510 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3868_
timestamp 0
transform -1 0 8570 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3869_
timestamp 0
transform 1 0 7990 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3870_
timestamp 0
transform -1 0 7870 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3872_
timestamp 0
transform 1 0 5710 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3873_
timestamp 0
transform -1 0 9550 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3874_
timestamp 0
transform 1 0 9890 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__3875_
timestamp 0
transform 1 0 6930 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3876_
timestamp 0
transform 1 0 5030 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3877_
timestamp 0
transform -1 0 4670 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3878_
timestamp 0
transform 1 0 4830 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3879_
timestamp 0
transform 1 0 4590 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3880_
timestamp 0
transform 1 0 5150 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3881_
timestamp 0
transform -1 0 5370 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3882_
timestamp 0
transform -1 0 4390 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__3883_
timestamp 0
transform -1 0 5010 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3884_
timestamp 0
transform -1 0 4830 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3885_
timestamp 0
transform 1 0 5190 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3886_
timestamp 0
transform 1 0 9690 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__3887_
timestamp 0
transform 1 0 10410 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__3888_
timestamp 0
transform 1 0 10370 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__3889_
timestamp 0
transform -1 0 10870 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__3890_
timestamp 0
transform -1 0 10790 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3892_
timestamp 0
transform -1 0 8810 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__3893_
timestamp 0
transform -1 0 8610 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__3894_
timestamp 0
transform -1 0 11310 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__3895_
timestamp 0
transform 1 0 11090 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__3896_
timestamp 0
transform 1 0 11850 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__3897_
timestamp 0
transform 1 0 11110 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__3898_
timestamp 0
transform 1 0 8290 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3899_
timestamp 0
transform -1 0 5650 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3900_
timestamp 0
transform 1 0 4110 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3901_
timestamp 0
transform -1 0 5070 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__3902_
timestamp 0
transform 1 0 4990 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3903_
timestamp 0
transform 1 0 7470 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3904_
timestamp 0
transform -1 0 7050 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3905_
timestamp 0
transform -1 0 6490 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3906_
timestamp 0
transform 1 0 5070 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3907_
timestamp 0
transform -1 0 8230 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__3908_
timestamp 0
transform -1 0 6830 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3909_
timestamp 0
transform -1 0 6010 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__3910_
timestamp 0
transform 1 0 5890 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__3912_
timestamp 0
transform 1 0 4370 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__3913_
timestamp 0
transform -1 0 4590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__3914_
timestamp 0
transform 1 0 4250 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__3915_
timestamp 0
transform 1 0 4790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__3916_
timestamp 0
transform 1 0 4990 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__3917_
timestamp 0
transform 1 0 5370 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__3918_
timestamp 0
transform -1 0 4690 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3919_
timestamp 0
transform 1 0 4790 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__3920_
timestamp 0
transform 1 0 4510 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3921_
timestamp 0
transform 1 0 830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3922_
timestamp 0
transform 1 0 930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__3923_
timestamp 0
transform 1 0 450 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3924_
timestamp 0
transform 1 0 810 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__3925_
timestamp 0
transform 1 0 5110 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3926_
timestamp 0
transform 1 0 5310 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3927_
timestamp 0
transform -1 0 4730 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3928_
timestamp 0
transform 1 0 5490 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3929_
timestamp 0
transform -1 0 4610 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__3930_
timestamp 0
transform 1 0 3450 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__3932_
timestamp 0
transform 1 0 2350 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__3933_
timestamp 0
transform 1 0 3250 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__3934_
timestamp 0
transform -1 0 4490 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__3935_
timestamp 0
transform 1 0 3850 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3936_
timestamp 0
transform 1 0 3650 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__3937_
timestamp 0
transform 1 0 4230 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__3938_
timestamp 0
transform -1 0 3510 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__3939_
timestamp 0
transform 1 0 3610 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__3940_
timestamp 0
transform -1 0 4750 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__3941_
timestamp 0
transform 1 0 6950 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3942_
timestamp 0
transform -1 0 10030 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3943_
timestamp 0
transform -1 0 10010 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__3944_
timestamp 0
transform -1 0 9710 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__3945_
timestamp 0
transform -1 0 10230 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3946_
timestamp 0
transform 1 0 9810 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__3947_
timestamp 0
transform 1 0 10410 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3948_
timestamp 0
transform 1 0 10590 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3949_
timestamp 0
transform 1 0 7710 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__3950_
timestamp 0
transform -1 0 6990 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3952_
timestamp 0
transform -1 0 5810 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__3953_
timestamp 0
transform 1 0 5470 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3954_
timestamp 0
transform -1 0 5870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3955_
timestamp 0
transform 1 0 5930 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3956_
timestamp 0
transform -1 0 6150 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3957_
timestamp 0
transform 1 0 6170 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3958_
timestamp 0
transform 1 0 6370 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3959_
timestamp 0
transform 1 0 6490 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3960_
timestamp 0
transform 1 0 2410 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3961_
timestamp 0
transform -1 0 2810 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3962_
timestamp 0
transform 1 0 2950 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3963_
timestamp 0
transform 1 0 3550 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3964_
timestamp 0
transform -1 0 4130 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3965_
timestamp 0
transform -1 0 3370 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3966_
timestamp 0
transform -1 0 4330 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3967_
timestamp 0
transform -1 0 5130 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3968_
timestamp 0
transform -1 0 5330 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3969_
timestamp 0
transform -1 0 4330 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3970_
timestamp 0
transform 1 0 3950 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3972_
timestamp 0
transform 1 0 5470 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__3973_
timestamp 0
transform 1 0 5470 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3974_
timestamp 0
transform -1 0 5690 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3975_
timestamp 0
transform -1 0 5690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3976_
timestamp 0
transform -1 0 5690 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3977_
timestamp 0
transform 1 0 5570 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__3978_
timestamp 0
transform 1 0 6390 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3979_
timestamp 0
transform -1 0 2750 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3980_
timestamp 0
transform 1 0 2050 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__3981_
timestamp 0
transform 1 0 1890 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__3982_
timestamp 0
transform 1 0 1830 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__3983_
timestamp 0
transform -1 0 1970 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__3984_
timestamp 0
transform 1 0 8290 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__3985_
timestamp 0
transform 1 0 6870 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3986_
timestamp 0
transform -1 0 7370 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__3987_
timestamp 0
transform 1 0 7650 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__3988_
timestamp 0
transform 1 0 7570 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3989_
timestamp 0
transform 1 0 7370 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3990_
timestamp 0
transform 1 0 7170 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3992_
timestamp 0
transform -1 0 7990 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3993_
timestamp 0
transform 1 0 7750 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3994_
timestamp 0
transform -1 0 7090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__3995_
timestamp 0
transform -1 0 9450 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3996_
timestamp 0
transform -1 0 6050 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__3997_
timestamp 0
transform 1 0 6010 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__3998_
timestamp 0
transform -1 0 6090 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__3999_
timestamp 0
transform 1 0 5870 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4000_
timestamp 0
transform -1 0 5290 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4001_
timestamp 0
transform -1 0 5130 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4002_
timestamp 0
transform -1 0 6990 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4003_
timestamp 0
transform -1 0 6630 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4004_
timestamp 0
transform 1 0 2670 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4005_
timestamp 0
transform 1 0 2870 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4006_
timestamp 0
transform -1 0 2690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4007_
timestamp 0
transform 1 0 2470 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4008_
timestamp 0
transform -1 0 7150 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4009_
timestamp 0
transform 1 0 6930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4010_
timestamp 0
transform -1 0 6790 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4012_
timestamp 0
transform 1 0 6770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4013_
timestamp 0
transform 1 0 6650 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4014_
timestamp 0
transform 1 0 6190 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4015_
timestamp 0
transform 1 0 6550 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4016_
timestamp 0
transform 1 0 9370 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4017_
timestamp 0
transform -1 0 9690 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4018_
timestamp 0
transform -1 0 9870 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4019_
timestamp 0
transform 1 0 10030 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4020_
timestamp 0
transform -1 0 7510 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4021_
timestamp 0
transform -1 0 10070 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4022_
timestamp 0
transform -1 0 6850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4023_
timestamp 0
transform -1 0 7190 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4024_
timestamp 0
transform 1 0 8990 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4025_
timestamp 0
transform -1 0 7710 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4026_
timestamp 0
transform -1 0 7870 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4027_
timestamp 0
transform 1 0 8410 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4028_
timestamp 0
transform 1 0 7950 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4029_
timestamp 0
transform 1 0 11050 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4030_
timestamp 0
transform 1 0 10870 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4032_
timestamp 0
transform 1 0 8690 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4033_
timestamp 0
transform -1 0 9350 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4034_
timestamp 0
transform 1 0 4010 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4035_
timestamp 0
transform 1 0 9810 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4036_
timestamp 0
transform -1 0 9670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4037_
timestamp 0
transform -1 0 9190 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4038_
timestamp 0
transform -1 0 8150 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4039_
timestamp 0
transform -1 0 7090 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4040_
timestamp 0
transform 1 0 12030 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4041_
timestamp 0
transform 1 0 9310 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4042_
timestamp 0
transform -1 0 6030 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__4043_
timestamp 0
transform 1 0 5350 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4044_
timestamp 0
transform -1 0 5430 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4045_
timestamp 0
transform -1 0 5490 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4046_
timestamp 0
transform -1 0 5850 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4047_
timestamp 0
transform -1 0 6030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4048_
timestamp 0
transform -1 0 6030 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4049_
timestamp 0
transform 1 0 5510 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4050_
timestamp 0
transform -1 0 5290 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4052_
timestamp 0
transform -1 0 6250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4053_
timestamp 0
transform -1 0 8230 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4054_
timestamp 0
transform 1 0 3750 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4055_
timestamp 0
transform -1 0 3590 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4056_
timestamp 0
transform 1 0 2750 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4057_
timestamp 0
transform 1 0 3370 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4058_
timestamp 0
transform -1 0 7510 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4059_
timestamp 0
transform 1 0 7370 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4060_
timestamp 0
transform -1 0 8050 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4061_
timestamp 0
transform -1 0 8990 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4062_
timestamp 0
transform -1 0 3170 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4063_
timestamp 0
transform 1 0 5090 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4064_
timestamp 0
transform -1 0 5070 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4065_
timestamp 0
transform 1 0 5290 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4066_
timestamp 0
transform 1 0 4490 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4067_
timestamp 0
transform -1 0 7130 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4068_
timestamp 0
transform 1 0 3150 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4069_
timestamp 0
transform -1 0 690 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__4070_
timestamp 0
transform 1 0 1170 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__4072_
timestamp 0
transform -1 0 890 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__4073_
timestamp 0
transform 1 0 4110 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4074_
timestamp 0
transform 1 0 4310 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4075_
timestamp 0
transform 1 0 4230 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4076_
timestamp 0
transform -1 0 5490 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4077_
timestamp 0
transform 1 0 5510 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4078_
timestamp 0
transform -1 0 5530 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4079_
timestamp 0
transform 1 0 3790 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4080_
timestamp 0
transform 1 0 5890 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4081_
timestamp 0
transform 1 0 930 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4082_
timestamp 0
transform 1 0 4170 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4083_
timestamp 0
transform -1 0 3970 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4084_
timestamp 0
transform 1 0 1670 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4085_
timestamp 0
transform 1 0 1490 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4086_
timestamp 0
transform 1 0 1630 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4087_
timestamp 0
transform 1 0 1590 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4088_
timestamp 0
transform -1 0 4530 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4089_
timestamp 0
transform -1 0 4490 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4090_
timestamp 0
transform -1 0 3990 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4092_
timestamp 0
transform -1 0 5710 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4093_
timestamp 0
transform 1 0 4650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4094_
timestamp 0
transform 1 0 4230 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4095_
timestamp 0
transform 1 0 1970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4096_
timestamp 0
transform 1 0 1790 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4097_
timestamp 0
transform 1 0 1670 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4098_
timestamp 0
transform 1 0 1590 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4099_
timestamp 0
transform 1 0 7170 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4100_
timestamp 0
transform 1 0 8050 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4101_
timestamp 0
transform 1 0 8210 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4102_
timestamp 0
transform -1 0 8410 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4103_
timestamp 0
transform 1 0 8030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4104_
timestamp 0
transform -1 0 8250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4105_
timestamp 0
transform 1 0 8690 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4106_
timestamp 0
transform 1 0 6730 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4107_
timestamp 0
transform -1 0 1130 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4__4108_
timestamp 0
transform -1 0 530 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__4109_
timestamp 0
transform -1 0 1870 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4110_
timestamp 0
transform -1 0 7810 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4112_
timestamp 0
transform 1 0 2930 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__4113_
timestamp 0
transform 1 0 3130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__4114_
timestamp 0
transform 1 0 3630 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4115_
timestamp 0
transform 1 0 4510 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4116_
timestamp 0
transform -1 0 5390 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4117_
timestamp 0
transform 1 0 4930 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4118_
timestamp 0
transform 1 0 4850 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4119_
timestamp 0
transform 1 0 4010 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4120_
timestamp 0
transform -1 0 3750 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4121_
timestamp 0
transform -1 0 4590 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4122_
timestamp 0
transform 1 0 4730 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4123_
timestamp 0
transform 1 0 8090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4124_
timestamp 0
transform 1 0 8610 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4125_
timestamp 0
transform -1 0 4330 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4126_
timestamp 0
transform 1 0 4290 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4127_
timestamp 0
transform 1 0 4110 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4128_
timestamp 0
transform 1 0 4530 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4129_
timestamp 0
transform -1 0 4950 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4130_
timestamp 0
transform 1 0 6070 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4132_
timestamp 0
transform -1 0 4570 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4133_
timestamp 0
transform -1 0 2050 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4134_
timestamp 0
transform 1 0 1830 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4135_
timestamp 0
transform -1 0 2190 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__4136_
timestamp 0
transform -1 0 2190 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4137_
timestamp 0
transform -1 0 2030 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__4138_
timestamp 0
transform -1 0 2270 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4139_
timestamp 0
transform 1 0 2050 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4140_
timestamp 0
transform -1 0 3070 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4141_
timestamp 0
transform 1 0 1850 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4142_
timestamp 0
transform 1 0 1650 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4143_
timestamp 0
transform -1 0 1490 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4144_
timestamp 0
transform 1 0 1630 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4145_
timestamp 0
transform -1 0 1110 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4146_
timestamp 0
transform 1 0 3130 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4147_
timestamp 0
transform -1 0 2070 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4148_
timestamp 0
transform -1 0 3250 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4149_
timestamp 0
transform 1 0 3230 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4150_
timestamp 0
transform 1 0 3230 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4152_
timestamp 0
transform -1 0 3710 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4153_
timestamp 0
transform -1 0 2090 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4154_
timestamp 0
transform -1 0 2290 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4155_
timestamp 0
transform 1 0 670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4156_
timestamp 0
transform 1 0 1030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4157_
timestamp 0
transform -1 0 5970 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4158_
timestamp 0
transform 1 0 6130 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4159_
timestamp 0
transform 1 0 6330 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4160_
timestamp 0
transform 1 0 5410 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4161_
timestamp 0
transform -1 0 5630 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4162_
timestamp 0
transform 1 0 5210 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4163_
timestamp 0
transform -1 0 5230 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4164_
timestamp 0
transform 1 0 5770 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4165_
timestamp 0
transform -1 0 5770 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4166_
timestamp 0
transform 1 0 5790 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4167_
timestamp 0
transform 1 0 6490 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4168_
timestamp 0
transform -1 0 5930 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4169_
timestamp 0
transform 1 0 5730 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4170_
timestamp 0
transform 1 0 6130 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4172_
timestamp 0
transform 1 0 5170 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4173_
timestamp 0
transform 1 0 3850 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4174_
timestamp 0
transform 1 0 5570 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4175_
timestamp 0
transform 1 0 5190 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4176_
timestamp 0
transform -1 0 3370 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4177_
timestamp 0
transform 1 0 3050 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4178_
timestamp 0
transform -1 0 2270 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4179_
timestamp 0
transform -1 0 2390 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__4180_
timestamp 0
transform 1 0 2850 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4181_
timestamp 0
transform -1 0 2470 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4182_
timestamp 0
transform 1 0 2310 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4183_
timestamp 0
transform -1 0 3290 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4184_
timestamp 0
transform 1 0 3450 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4185_
timestamp 0
transform 1 0 2870 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4186_
timestamp 0
transform -1 0 2490 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4187_
timestamp 0
transform 1 0 4110 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4188_
timestamp 0
transform 1 0 4310 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4189_
timestamp 0
transform -1 0 4130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4190_
timestamp 0
transform -1 0 3950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4192_
timestamp 0
transform -1 0 5230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4193_
timestamp 0
transform -1 0 5090 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4194_
timestamp 0
transform -1 0 3950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4195_
timestamp 0
transform 1 0 3490 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4196_
timestamp 0
transform 1 0 3790 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4197_
timestamp 0
transform 1 0 1650 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4198_
timestamp 0
transform -1 0 1770 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4199_
timestamp 0
transform -1 0 1970 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4200_
timestamp 0
transform -1 0 2370 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4201_
timestamp 0
transform -1 0 1590 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4202_
timestamp 0
transform -1 0 1470 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__4203_
timestamp 0
transform -1 0 1850 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__4204_
timestamp 0
transform -1 0 2650 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4205_
timestamp 0
transform 1 0 2650 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4206_
timestamp 0
transform -1 0 8630 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4207_
timestamp 0
transform -1 0 7970 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4208_
timestamp 0
transform -1 0 6310 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4209_
timestamp 0
transform -1 0 310 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4210_
timestamp 0
transform 1 0 90 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4212_
timestamp 0
transform -1 0 490 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4213_
timestamp 0
transform 1 0 950 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4214_
timestamp 0
transform -1 0 1470 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4215_
timestamp 0
transform 1 0 1450 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4216_
timestamp 0
transform -1 0 2050 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4217_
timestamp 0
transform -1 0 3030 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4218_
timestamp 0
transform -1 0 2250 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4219_
timestamp 0
transform 1 0 2330 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4220_
timestamp 0
transform 1 0 2530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4221_
timestamp 0
transform -1 0 310 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4222_
timestamp 0
transform -1 0 110 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4223_
timestamp 0
transform -1 0 490 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4224_
timestamp 0
transform -1 0 490 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4225_
timestamp 0
transform -1 0 470 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4226_
timestamp 0
transform 1 0 90 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4227_
timestamp 0
transform -1 0 310 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4228_
timestamp 0
transform -1 0 2450 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4229_
timestamp 0
transform 1 0 2650 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4230_
timestamp 0
transform -1 0 2870 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4232_
timestamp 0
transform -1 0 3670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4233_
timestamp 0
transform -1 0 2250 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4234_
timestamp 0
transform -1 0 3110 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4235_
timestamp 0
transform -1 0 3870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4236_
timestamp 0
transform 1 0 3950 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4237_
timestamp 0
transform -1 0 4170 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4238_
timestamp 0
transform 1 0 3490 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4239_
timestamp 0
transform 1 0 2650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4240_
timestamp 0
transform 1 0 2290 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4241_
timestamp 0
transform -1 0 2150 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4242_
timestamp 0
transform 1 0 2330 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4243_
timestamp 0
transform -1 0 4510 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4244_
timestamp 0
transform -1 0 5510 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4245_
timestamp 0
transform -1 0 6090 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4246_
timestamp 0
transform -1 0 4210 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4247_
timestamp 0
transform 1 0 2610 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4248_
timestamp 0
transform -1 0 5690 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4249_
timestamp 0
transform -1 0 2390 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4250_
timestamp 0
transform -1 0 4310 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4252_
timestamp 0
transform -1 0 5890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4253_
timestamp 0
transform -1 0 3790 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4254_
timestamp 0
transform -1 0 2210 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4255_
timestamp 0
transform 1 0 2550 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4256_
timestamp 0
transform -1 0 3910 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4257_
timestamp 0
transform 1 0 4090 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4258_
timestamp 0
transform 1 0 4290 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4259_
timestamp 0
transform 1 0 4050 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4260_
timestamp 0
transform -1 0 3010 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4261_
timestamp 0
transform -1 0 4070 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4262_
timestamp 0
transform 1 0 1590 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4263_
timestamp 0
transform -1 0 8010 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4264_
timestamp 0
transform 1 0 7630 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4265_
timestamp 0
transform 1 0 7450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4266_
timestamp 0
transform 1 0 7130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4267_
timestamp 0
transform 1 0 7570 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4268_
timestamp 0
transform -1 0 6810 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4269_
timestamp 0
transform -1 0 9490 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4270_
timestamp 0
transform -1 0 11190 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4272_
timestamp 0
transform 1 0 9270 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4273_
timestamp 0
transform 1 0 9070 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4274_
timestamp 0
transform -1 0 8990 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4275_
timestamp 0
transform 1 0 8810 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4276_
timestamp 0
transform 1 0 8890 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4277_
timestamp 0
transform 1 0 8910 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4278_
timestamp 0
transform 1 0 7790 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4279_
timestamp 0
transform 1 0 10570 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4280_
timestamp 0
transform 1 0 10770 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4281_
timestamp 0
transform -1 0 10730 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4282_
timestamp 0
transform -1 0 1270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4283_
timestamp 0
transform -1 0 7110 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4284_
timestamp 0
transform 1 0 7690 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4285_
timestamp 0
transform 1 0 7430 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4286_
timestamp 0
transform -1 0 1110 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4287_
timestamp 0
transform -1 0 1310 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4288_
timestamp 0
transform -1 0 1710 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4289_
timestamp 0
transform -1 0 4410 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4290_
timestamp 0
transform 1 0 6890 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4292_
timestamp 0
transform -1 0 2570 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4293_
timestamp 0
transform -1 0 1850 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4294_
timestamp 0
transform -1 0 7330 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4295_
timestamp 0
transform 1 0 1530 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4296_
timestamp 0
transform -1 0 110 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4297_
timestamp 0
transform 1 0 1190 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4298_
timestamp 0
transform -1 0 3310 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4299_
timestamp 0
transform 1 0 3390 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4300_
timestamp 0
transform -1 0 3870 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4301_
timestamp 0
transform -1 0 3590 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4302_
timestamp 0
transform -1 0 3710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4303_
timestamp 0
transform -1 0 1630 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4304_
timestamp 0
transform 1 0 1210 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4305_
timestamp 0
transform -1 0 2330 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4306_
timestamp 0
transform -1 0 2890 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4307_
timestamp 0
transform 1 0 6250 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4308_
timestamp 0
transform -1 0 6330 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4309_
timestamp 0
transform 1 0 2890 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4310_
timestamp 0
transform -1 0 2470 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4312_
timestamp 0
transform 1 0 950 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4313_
timestamp 0
transform 1 0 1530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4314_
timestamp 0
transform 1 0 1710 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4315_
timestamp 0
transform -1 0 2750 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4316_
timestamp 0
transform -1 0 2810 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4317_
timestamp 0
transform 1 0 4450 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4318_
timestamp 0
transform 1 0 4130 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4319_
timestamp 0
transform 1 0 3630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4320_
timestamp 0
transform -1 0 3070 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4321_
timestamp 0
transform 1 0 2850 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4322_
timestamp 0
transform 1 0 1590 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4323_
timestamp 0
transform -1 0 2710 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4324_
timestamp 0
transform -1 0 1850 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4325_
timestamp 0
transform -1 0 4110 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4326_
timestamp 0
transform 1 0 4010 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4327_
timestamp 0
transform 1 0 4150 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4328_
timestamp 0
transform -1 0 8590 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4329_
timestamp 0
transform 1 0 1750 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4330_
timestamp 0
transform 1 0 2150 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4332_
timestamp 0
transform -1 0 2010 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4333_
timestamp 0
transform -1 0 2930 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4334_
timestamp 0
transform -1 0 3130 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4335_
timestamp 0
transform -1 0 3710 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4336_
timestamp 0
transform 1 0 2870 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4337_
timestamp 0
transform 1 0 2670 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4338_
timestamp 0
transform 1 0 2710 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4339_
timestamp 0
transform -1 0 3330 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4340_
timestamp 0
transform -1 0 3510 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4341_
timestamp 0
transform 1 0 3450 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4342_
timestamp 0
transform -1 0 3270 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4343_
timestamp 0
transform 1 0 3510 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4344_
timestamp 0
transform 1 0 1810 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4345_
timestamp 0
transform -1 0 2450 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4346_
timestamp 0
transform 1 0 6930 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4347_
timestamp 0
transform -1 0 6750 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4348_
timestamp 0
transform -1 0 650 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4349_
timestamp 0
transform -1 0 1070 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4350_
timestamp 0
transform 1 0 2190 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4352_
timestamp 0
transform 1 0 3790 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4353_
timestamp 0
transform -1 0 6190 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4354_
timestamp 0
transform -1 0 3470 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4355_
timestamp 0
transform -1 0 890 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4356_
timestamp 0
transform -1 0 530 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4357_
timestamp 0
transform 1 0 2390 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4358_
timestamp 0
transform -1 0 5250 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4359_
timestamp 0
transform 1 0 5170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4360_
timestamp 0
transform -1 0 5130 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4361_
timestamp 0
transform 1 0 3070 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4362_
timestamp 0
transform 1 0 4910 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4363_
timestamp 0
transform -1 0 4750 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4364_
timestamp 0
transform 1 0 3710 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4365_
timestamp 0
transform -1 0 5690 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4366_
timestamp 0
transform -1 0 5890 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4367_
timestamp 0
transform -1 0 2930 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4368_
timestamp 0
transform 1 0 7570 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4369_
timestamp 0
transform -1 0 7410 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4370_
timestamp 0
transform 1 0 690 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4372_
timestamp 0
transform 1 0 1950 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4373_
timestamp 0
transform 1 0 2150 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4374_
timestamp 0
transform 1 0 2510 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4375_
timestamp 0
transform -1 0 3830 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4376_
timestamp 0
transform 1 0 7510 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4377_
timestamp 0
transform 1 0 11570 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4378_
timestamp 0
transform -1 0 1290 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4379_
timestamp 0
transform -1 0 5250 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4380_
timestamp 0
transform 1 0 4830 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4381_
timestamp 0
transform 1 0 5930 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4382_
timestamp 0
transform 1 0 270 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4383_
timestamp 0
transform 1 0 90 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4384_
timestamp 0
transform 1 0 6270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4385_
timestamp 0
transform 1 0 6470 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4386_
timestamp 0
transform 1 0 6870 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4387_
timestamp 0
transform 1 0 6670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4388_
timestamp 0
transform -1 0 5470 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4389_
timestamp 0
transform -1 0 6570 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4390_
timestamp 0
transform 1 0 7070 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4392_
timestamp 0
transform -1 0 6370 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4393_
timestamp 0
transform 1 0 6530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4394_
timestamp 0
transform 1 0 6710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4395_
timestamp 0
transform 1 0 6830 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4396_
timestamp 0
transform -1 0 6310 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4397_
timestamp 0
transform 1 0 4070 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4398_
timestamp 0
transform 1 0 3050 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4399_
timestamp 0
transform 1 0 2170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4400_
timestamp 0
transform -1 0 6350 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4401_
timestamp 0
transform 1 0 6270 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4402_
timestamp 0
transform -1 0 6110 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4403_
timestamp 0
transform -1 0 5650 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4404_
timestamp 0
transform 1 0 1430 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4405_
timestamp 0
transform -1 0 1870 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4406_
timestamp 0
transform -1 0 2570 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4407_
timestamp 0
transform -1 0 2370 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4408_
timestamp 0
transform 1 0 1590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4409_
timestamp 0
transform -1 0 1810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4410_
timestamp 0
transform 1 0 3610 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4412_
timestamp 0
transform 1 0 1770 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4413_
timestamp 0
transform -1 0 290 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4414_
timestamp 0
transform 1 0 290 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4415_
timestamp 0
transform 1 0 470 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4416_
timestamp 0
transform 1 0 1550 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__4417_
timestamp 0
transform -1 0 1770 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__4418_
timestamp 0
transform -1 0 2590 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__4419_
timestamp 0
transform 1 0 2150 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__4420_
timestamp 0
transform 1 0 2270 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4421_
timestamp 0
transform 1 0 2470 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4422_
timestamp 0
transform -1 0 2010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4423_
timestamp 0
transform -1 0 650 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4424_
timestamp 0
transform 1 0 2070 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4425_
timestamp 0
transform 1 0 1110 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4426_
timestamp 0
transform 1 0 1310 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4427_
timestamp 0
transform 1 0 3570 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4428_
timestamp 0
transform -1 0 3410 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4429_
timestamp 0
transform 1 0 1290 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4430_
timestamp 0
transform 1 0 1490 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4432_
timestamp 0
transform -1 0 650 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4433_
timestamp 0
transform -1 0 890 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4434_
timestamp 0
transform -1 0 1350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__4435_
timestamp 0
transform 1 0 1530 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__4436_
timestamp 0
transform 1 0 3130 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__4437_
timestamp 0
transform -1 0 3350 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__4438_
timestamp 0
transform -1 0 6590 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4439_
timestamp 0
transform 1 0 5990 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4440_
timestamp 0
transform -1 0 4770 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4441_
timestamp 0
transform 1 0 4170 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4442_
timestamp 0
transform 1 0 3950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__4443_
timestamp 0
transform 1 0 3830 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4444_
timestamp 0
transform 1 0 3650 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4445_
timestamp 0
transform 1 0 3990 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4446_
timestamp 0
transform 1 0 4410 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4447_
timestamp 0
transform 1 0 4590 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4448_
timestamp 0
transform 1 0 2510 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4449_
timestamp 0
transform 1 0 1070 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4450_
timestamp 0
transform -1 0 1830 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__4452_
timestamp 0
transform -1 0 2230 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4453_
timestamp 0
transform 1 0 7250 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4454_
timestamp 0
transform -1 0 1070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4455_
timestamp 0
transform 1 0 6790 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4456_
timestamp 0
transform 1 0 7010 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4457_
timestamp 0
transform 1 0 7210 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4458_
timestamp 0
transform -1 0 7410 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4459_
timestamp 0
transform -1 0 7030 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4460_
timestamp 0
transform -1 0 8350 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4461_
timestamp 0
transform 1 0 7630 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4462_
timestamp 0
transform -1 0 6730 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4463_
timestamp 0
transform 1 0 1250 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4464_
timestamp 0
transform -1 0 2550 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4465_
timestamp 0
transform -1 0 5890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4466_
timestamp 0
transform 1 0 6030 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4467_
timestamp 0
transform 1 0 6450 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4468_
timestamp 0
transform 1 0 6690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4469_
timestamp 0
transform 1 0 6890 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4470_
timestamp 0
transform -1 0 6650 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4472_
timestamp 0
transform -1 0 6450 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4473_
timestamp 0
transform 1 0 8170 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4474_
timestamp 0
transform -1 0 6270 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4475_
timestamp 0
transform 1 0 2730 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4476_
timestamp 0
transform -1 0 1230 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4477_
timestamp 0
transform -1 0 2630 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4478_
timestamp 0
transform 1 0 2610 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4479_
timestamp 0
transform 1 0 5330 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4480_
timestamp 0
transform 1 0 1410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4481_
timestamp 0
transform 1 0 250 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4482_
timestamp 0
transform 1 0 450 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4483_
timestamp 0
transform 1 0 3210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4484_
timestamp 0
transform -1 0 4970 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4485_
timestamp 0
transform 1 0 5350 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4486_
timestamp 0
transform -1 0 5170 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4487_
timestamp 0
transform -1 0 5550 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4488_
timestamp 0
transform 1 0 5710 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4489_
timestamp 0
transform -1 0 5830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4490_
timestamp 0
transform -1 0 5790 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4492_
timestamp 0
transform 1 0 90 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4493_
timestamp 0
transform -1 0 5710 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__4494_
timestamp 0
transform 1 0 5510 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__4495_
timestamp 0
transform 1 0 4370 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4496_
timestamp 0
transform 1 0 3830 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4497_
timestamp 0
transform -1 0 3610 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4498_
timestamp 0
transform -1 0 4650 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4499_
timestamp 0
transform 1 0 1270 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4500_
timestamp 0
transform 1 0 6370 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__4501_
timestamp 0
transform 1 0 6090 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4502_
timestamp 0
transform -1 0 4530 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__4503_
timestamp 0
transform 1 0 6490 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4504_
timestamp 0
transform -1 0 1730 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__4505_
timestamp 0
transform -1 0 4850 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__4506_
timestamp 0
transform -1 0 5290 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4507_
timestamp 0
transform 1 0 5670 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__4508_
timestamp 0
transform 1 0 5550 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4509_
timestamp 0
transform -1 0 5770 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4510_
timestamp 0
transform -1 0 5950 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4511_
timestamp 0
transform 1 0 6110 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4513_
timestamp 0
transform 1 0 6230 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4514_
timestamp 0
transform -1 0 1730 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__4515_
timestamp 0
transform -1 0 2570 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__4516_
timestamp 0
transform -1 0 4690 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__4517_
timestamp 0
transform -1 0 5170 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4518_
timestamp 0
transform 1 0 5130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4519_
timestamp 0
transform 1 0 5490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4520_
timestamp 0
transform -1 0 5690 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4521_
timestamp 0
transform 1 0 6530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4522_
timestamp 0
transform -1 0 8950 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4523_
timestamp 0
transform 1 0 5330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4524_
timestamp 0
transform 1 0 6030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4525_
timestamp 0
transform 1 0 5890 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4526_
timestamp 0
transform -1 0 6470 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4527_
timestamp 0
transform -1 0 4970 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4528_
timestamp 0
transform 1 0 6370 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4529_
timestamp 0
transform 1 0 6070 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4530_
timestamp 0
transform 1 0 6050 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4531_
timestamp 0
transform -1 0 2290 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__4533_
timestamp 0
transform -1 0 6250 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4534_
timestamp 0
transform 1 0 4290 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4535_
timestamp 0
transform 1 0 3690 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4536_
timestamp 0
transform -1 0 1110 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4537_
timestamp 0
transform 1 0 4470 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4538_
timestamp 0
transform -1 0 7710 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4539_
timestamp 0
transform -1 0 3090 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4540_
timestamp 0
transform 1 0 7670 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4541_
timestamp 0
transform 1 0 6530 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4542_
timestamp 0
transform 1 0 3070 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4543_
timestamp 0
transform -1 0 2910 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4544_
timestamp 0
transform -1 0 930 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4545_
timestamp 0
transform 1 0 2150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4546_
timestamp 0
transform 1 0 2930 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4547_
timestamp 0
transform -1 0 2390 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4548_
timestamp 0
transform -1 0 1770 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4549_
timestamp 0
transform 1 0 2630 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4550_
timestamp 0
transform 1 0 2830 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4551_
timestamp 0
transform -1 0 3030 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4553_
timestamp 0
transform -1 0 6570 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4554_
timestamp 0
transform 1 0 1010 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4555_
timestamp 0
transform -1 0 770 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__4556_
timestamp 0
transform 1 0 4370 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4557_
timestamp 0
transform 1 0 4190 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4558_
timestamp 0
transform -1 0 4030 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4559_
timestamp 0
transform 1 0 5050 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4560_
timestamp 0
transform -1 0 8510 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4561_
timestamp 0
transform -1 0 8910 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4562_
timestamp 0
transform 1 0 8430 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4563_
timestamp 0
transform -1 0 6410 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4564_
timestamp 0
transform -1 0 1910 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4565_
timestamp 0
transform 1 0 2730 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4566_
timestamp 0
transform 1 0 3110 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4567_
timestamp 0
transform -1 0 6810 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4568_
timestamp 0
transform 1 0 6730 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4569_
timestamp 0
transform 1 0 1950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4570_
timestamp 0
transform -1 0 6610 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4571_
timestamp 0
transform 1 0 6310 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4573_
timestamp 0
transform -1 0 10410 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4574_
timestamp 0
transform -1 0 9590 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4575_
timestamp 0
transform -1 0 7010 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4576_
timestamp 0
transform -1 0 8530 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4577_
timestamp 0
transform -1 0 3050 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4578_
timestamp 0
transform -1 0 6010 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4579_
timestamp 0
transform 1 0 8030 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4580_
timestamp 0
transform 1 0 10210 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4581_
timestamp 0
transform -1 0 7550 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4582_
timestamp 0
transform 1 0 1310 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4583_
timestamp 0
transform -1 0 2390 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4584_
timestamp 0
transform -1 0 2230 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4585_
timestamp 0
transform -1 0 2130 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4586_
timestamp 0
transform -1 0 1950 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4587_
timestamp 0
transform -1 0 1610 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4588_
timestamp 0
transform 1 0 3330 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4589_
timestamp 0
transform 1 0 3870 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4590_
timestamp 0
transform 1 0 1250 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4591_
timestamp 0
transform -1 0 1670 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4593_
timestamp 0
transform -1 0 4030 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4594_
timestamp 0
transform -1 0 3190 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__4595_
timestamp 0
transform -1 0 2750 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4596_
timestamp 0
transform -1 0 2950 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4597_
timestamp 0
transform 1 0 2810 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__4598_
timestamp 0
transform -1 0 2730 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4599_
timestamp 0
transform -1 0 2910 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4600_
timestamp 0
transform -1 0 4070 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4601_
timestamp 0
transform -1 0 4030 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4602_
timestamp 0
transform -1 0 1450 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4603_
timestamp 0
transform -1 0 1390 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4604_
timestamp 0
transform -1 0 2990 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__4605_
timestamp 0
transform 1 0 1810 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4606_
timestamp 0
transform -1 0 710 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4607_
timestamp 0
transform -1 0 530 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4608_
timestamp 0
transform -1 0 3270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4609_
timestamp 0
transform 1 0 1650 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__4610_
timestamp 0
transform 1 0 2530 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4611_
timestamp 0
transform -1 0 2370 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4613_
timestamp 0
transform 1 0 2010 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__4614_
timestamp 0
transform -1 0 670 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4615_
timestamp 0
transform -1 0 490 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4616_
timestamp 0
transform -1 0 1850 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__4617_
timestamp 0
transform -1 0 1650 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__4618_
timestamp 0
transform -1 0 2550 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4619_
timestamp 0
transform -1 0 1890 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4620_
timestamp 0
transform -1 0 1490 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4621_
timestamp 0
transform 1 0 2150 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4622_
timestamp 0
transform 1 0 2570 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__4623_
timestamp 0
transform 1 0 2070 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4624_
timestamp 0
transform 1 0 1270 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__4625_
timestamp 0
transform 1 0 890 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4626_
timestamp 0
transform -1 0 730 0 1 11290
box -6 -8 26 248
use FILL  FILL_4__4627_
timestamp 0
transform -1 0 2230 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__4628_
timestamp 0
transform -1 0 1290 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__4629_
timestamp 0
transform 1 0 1070 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4__4630_
timestamp 0
transform 1 0 1030 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4631_
timestamp 0
transform 1 0 1610 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__4633_
timestamp 0
transform -1 0 590 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4634_
timestamp 0
transform -1 0 7610 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4635_
timestamp 0
transform -1 0 1550 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4636_
timestamp 0
transform 1 0 1350 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4637_
timestamp 0
transform -1 0 1750 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4638_
timestamp 0
transform -1 0 910 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4__4639_
timestamp 0
transform 1 0 1110 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4640_
timestamp 0
transform 1 0 970 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4641_
timestamp 0
transform -1 0 1130 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4642_
timestamp 0
transform -1 0 2950 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__4643_
timestamp 0
transform 1 0 3090 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4__4644_
timestamp 0
transform -1 0 3530 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__4645_
timestamp 0
transform -1 0 890 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4646_
timestamp 0
transform 1 0 670 0 1 10810
box -6 -8 26 248
use FILL  FILL_4__4647_
timestamp 0
transform -1 0 1290 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4648_
timestamp 0
transform -1 0 1230 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4649_
timestamp 0
transform -1 0 590 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4650_
timestamp 0
transform -1 0 830 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4__4651_
timestamp 0
transform 1 0 4130 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__4653_
timestamp 0
transform -1 0 4350 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__4654_
timestamp 0
transform -1 0 6910 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4655_
timestamp 0
transform 1 0 2570 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4656_
timestamp 0
transform -1 0 2390 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4657_
timestamp 0
transform -1 0 2310 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4658_
timestamp 0
transform 1 0 3750 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4659_
timestamp 0
transform -1 0 3970 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4660_
timestamp 0
transform -1 0 4350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4661_
timestamp 0
transform 1 0 4530 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4662_
timestamp 0
transform 1 0 3990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4663_
timestamp 0
transform 1 0 3430 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4664_
timestamp 0
transform 1 0 2570 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4665_
timestamp 0
transform -1 0 7850 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4666_
timestamp 0
transform 1 0 7750 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__4667_
timestamp 0
transform 1 0 6270 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__4668_
timestamp 0
transform -1 0 6490 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4__4669_
timestamp 0
transform 1 0 470 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4670_
timestamp 0
transform 1 0 4050 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4671_
timestamp 0
transform 1 0 3870 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4673_
timestamp 0
transform -1 0 3010 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4674_
timestamp 0
transform -1 0 3170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4675_
timestamp 0
transform -1 0 3050 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4676_
timestamp 0
transform -1 0 3650 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4677_
timestamp 0
transform -1 0 3590 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4678_
timestamp 0
transform 1 0 3410 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4679_
timestamp 0
transform -1 0 3250 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4680_
timestamp 0
transform -1 0 2250 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__4681_
timestamp 0
transform 1 0 2030 0 1 2650
box -6 -8 26 248
use FILL  FILL_4__4682_
timestamp 0
transform -1 0 7090 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4683_
timestamp 0
transform -1 0 1890 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4684_
timestamp 0
transform 1 0 3790 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4685_
timestamp 0
transform 1 0 3610 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4686_
timestamp 0
transform 1 0 11150 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4687_
timestamp 0
transform 1 0 11330 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4688_
timestamp 0
transform 1 0 11510 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4689_
timestamp 0
transform 1 0 11690 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4690_
timestamp 0
transform 1 0 10530 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4691_
timestamp 0
transform 1 0 10170 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4693_
timestamp 0
transform -1 0 9770 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4694_
timestamp 0
transform -1 0 9790 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4695_
timestamp 0
transform 1 0 10630 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4696_
timestamp 0
transform 1 0 10950 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4697_
timestamp 0
transform 1 0 11430 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4698_
timestamp 0
transform 1 0 11270 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4699_
timestamp 0
transform 1 0 11270 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4700_
timestamp 0
transform 1 0 11110 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4701_
timestamp 0
transform -1 0 11490 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4702_
timestamp 0
transform 1 0 11470 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4703_
timestamp 0
transform 1 0 11750 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4704_
timestamp 0
transform -1 0 11650 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4705_
timestamp 0
transform -1 0 11850 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4706_
timestamp 0
transform -1 0 11790 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4707_
timestamp 0
transform 1 0 10730 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4708_
timestamp 0
transform 1 0 10930 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4709_
timestamp 0
transform -1 0 10930 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4710_
timestamp 0
transform -1 0 10730 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4711_
timestamp 0
transform 1 0 10190 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4713_
timestamp 0
transform 1 0 9770 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4714_
timestamp 0
transform 1 0 9570 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4715_
timestamp 0
transform -1 0 9890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4716_
timestamp 0
transform 1 0 9310 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4717_
timestamp 0
transform 1 0 9650 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4718_
timestamp 0
transform -1 0 8790 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4719_
timestamp 0
transform 1 0 11330 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4720_
timestamp 0
transform 1 0 10070 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4721_
timestamp 0
transform 1 0 9890 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4722_
timestamp 0
transform -1 0 9970 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4723_
timestamp 0
transform -1 0 9970 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4724_
timestamp 0
transform 1 0 4270 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4725_
timestamp 0
transform -1 0 10170 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4726_
timestamp 0
transform -1 0 10370 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4727_
timestamp 0
transform -1 0 11130 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4728_
timestamp 0
transform 1 0 10210 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4729_
timestamp 0
transform -1 0 10150 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4730_
timestamp 0
transform -1 0 10030 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4731_
timestamp 0
transform -1 0 11710 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4733_
timestamp 0
transform 1 0 9850 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4734_
timestamp 0
transform -1 0 7830 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4735_
timestamp 0
transform 1 0 9370 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4736_
timestamp 0
transform -1 0 10070 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4737_
timestamp 0
transform 1 0 9570 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4738_
timestamp 0
transform -1 0 9770 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4739_
timestamp 0
transform -1 0 9950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4740_
timestamp 0
transform -1 0 10330 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4741_
timestamp 0
transform -1 0 10150 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4742_
timestamp 0
transform 1 0 10370 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4743_
timestamp 0
transform 1 0 10130 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4744_
timestamp 0
transform 1 0 10630 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4745_
timestamp 0
transform 1 0 10950 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4746_
timestamp 0
transform 1 0 10430 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4747_
timestamp 0
transform 1 0 8370 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4748_
timestamp 0
transform 1 0 8570 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4749_
timestamp 0
transform -1 0 8810 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4750_
timestamp 0
transform 1 0 8570 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4751_
timestamp 0
transform 1 0 3770 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4753_
timestamp 0
transform -1 0 8050 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4754_
timestamp 0
transform 1 0 8170 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4755_
timestamp 0
transform 1 0 7290 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4756_
timestamp 0
transform 1 0 6950 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4757_
timestamp 0
transform 1 0 8390 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4758_
timestamp 0
transform -1 0 10450 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4759_
timestamp 0
transform 1 0 10810 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4760_
timestamp 0
transform -1 0 11090 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4761_
timestamp 0
transform 1 0 11370 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4762_
timestamp 0
transform -1 0 10530 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4763_
timestamp 0
transform 1 0 11870 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4764_
timestamp 0
transform 1 0 10910 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4765_
timestamp 0
transform -1 0 11170 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4766_
timestamp 0
transform -1 0 10530 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4767_
timestamp 0
transform -1 0 10550 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4768_
timestamp 0
transform 1 0 10330 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4769_
timestamp 0
transform 1 0 10710 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4770_
timestamp 0
transform 1 0 11190 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4771_
timestamp 0
transform 1 0 12050 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4773_
timestamp 0
transform -1 0 8850 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4774_
timestamp 0
transform 1 0 2590 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4775_
timestamp 0
transform 1 0 2750 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4776_
timestamp 0
transform 1 0 2910 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4777_
timestamp 0
transform -1 0 3130 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4778_
timestamp 0
transform -1 0 3730 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4779_
timestamp 0
transform 1 0 3910 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4780_
timestamp 0
transform -1 0 8790 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4781_
timestamp 0
transform 1 0 3630 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4782_
timestamp 0
transform 1 0 3310 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4783_
timestamp 0
transform 1 0 9130 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4784_
timestamp 0
transform 1 0 7770 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4785_
timestamp 0
transform 1 0 2130 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4786_
timestamp 0
transform -1 0 4010 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__4787_
timestamp 0
transform -1 0 3690 0 1 3130
box -6 -8 26 248
use FILL  FILL_4__4788_
timestamp 0
transform -1 0 4210 0 1 3610
box -6 -8 26 248
use FILL  FILL_4__4789_
timestamp 0
transform 1 0 7250 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4790_
timestamp 0
transform 1 0 7310 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4791_
timestamp 0
transform -1 0 7850 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4793_
timestamp 0
transform -1 0 7850 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4794_
timestamp 0
transform -1 0 7490 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4795_
timestamp 0
transform -1 0 7550 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4796_
timestamp 0
transform 1 0 11850 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4797_
timestamp 0
transform 1 0 8590 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4798_
timestamp 0
transform 1 0 10050 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4799_
timestamp 0
transform -1 0 9890 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4800_
timestamp 0
transform 1 0 8530 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4801_
timestamp 0
transform 1 0 10990 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4802_
timestamp 0
transform -1 0 10530 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4803_
timestamp 0
transform -1 0 7430 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4804_
timestamp 0
transform -1 0 7110 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4805_
timestamp 0
transform -1 0 6990 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4806_
timestamp 0
transform -1 0 9350 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4807_
timestamp 0
transform -1 0 9130 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4808_
timestamp 0
transform -1 0 8750 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4809_
timestamp 0
transform -1 0 8750 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4810_
timestamp 0
transform -1 0 8990 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4811_
timestamp 0
transform 1 0 11970 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4813_
timestamp 0
transform 1 0 11510 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4814_
timestamp 0
transform 1 0 11390 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4815_
timestamp 0
transform -1 0 9090 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4816_
timestamp 0
transform -1 0 9530 0 1 7450
box -6 -8 26 248
use FILL  FILL_4__4817_
timestamp 0
transform -1 0 11590 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4818_
timestamp 0
transform -1 0 11530 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4819_
timestamp 0
transform -1 0 6470 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4820_
timestamp 0
transform 1 0 8030 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4821_
timestamp 0
transform 1 0 11670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4822_
timestamp 0
transform 1 0 11870 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4823_
timestamp 0
transform 1 0 11650 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4824_
timestamp 0
transform -1 0 11510 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4825_
timestamp 0
transform 1 0 11210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4826_
timestamp 0
transform -1 0 11050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4827_
timestamp 0
transform -1 0 11750 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4828_
timestamp 0
transform -1 0 11830 0 1 10330
box -6 -8 26 248
use FILL  FILL_4__4829_
timestamp 0
transform 1 0 11670 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4830_
timestamp 0
transform 1 0 9030 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4831_
timestamp 0
transform -1 0 9390 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4833_
timestamp 0
transform 1 0 8410 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4834_
timestamp 0
transform 1 0 8210 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4835_
timestamp 0
transform -1 0 8410 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4836_
timestamp 0
transform 1 0 9690 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4837_
timestamp 0
transform -1 0 10830 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4838_
timestamp 0
transform 1 0 11850 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4839_
timestamp 0
transform 1 0 12110 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4840_
timestamp 0
transform 1 0 9290 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4841_
timestamp 0
transform 1 0 10330 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4842_
timestamp 0
transform 1 0 12030 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4843_
timestamp 0
transform 1 0 11190 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4844_
timestamp 0
transform -1 0 11170 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4845_
timestamp 0
transform -1 0 11950 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4846_
timestamp 0
transform 1 0 11930 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4847_
timestamp 0
transform -1 0 8410 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4__4848_
timestamp 0
transform -1 0 8430 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4849_
timestamp 0
transform 1 0 9090 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4850_
timestamp 0
transform 1 0 9330 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4851_
timestamp 0
transform 1 0 11310 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4853_
timestamp 0
transform 1 0 12090 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4854_
timestamp 0
transform -1 0 11230 0 1 11770
box -6 -8 26 248
use FILL  FILL_4__4855_
timestamp 0
transform -1 0 8250 0 1 7930
box -6 -8 26 248
use FILL  FILL_4__4856_
timestamp 0
transform -1 0 8270 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4857_
timestamp 0
transform -1 0 10350 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4858_
timestamp 0
transform -1 0 10490 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4859_
timestamp 0
transform -1 0 7230 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4860_
timestamp 0
transform -1 0 10410 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4861_
timestamp 0
transform -1 0 10670 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4862_
timestamp 0
transform 1 0 11470 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4863_
timestamp 0
transform -1 0 10730 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4864_
timestamp 0
transform -1 0 10570 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4865_
timestamp 0
transform 1 0 10590 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4866_
timestamp 0
transform 1 0 11670 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4867_
timestamp 0
transform 1 0 11850 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4868_
timestamp 0
transform -1 0 11350 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4869_
timestamp 0
transform -1 0 10890 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4__4870_
timestamp 0
transform 1 0 8130 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4871_
timestamp 0
transform 1 0 7970 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4873_
timestamp 0
transform -1 0 11390 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4874_
timestamp 0
transform 1 0 11910 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4875_
timestamp 0
transform -1 0 7610 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4__4876_
timestamp 0
transform -1 0 10530 0 -1 9370
box -6 -8 26 248
use FILL  FILL_4__4877_
timestamp 0
transform 1 0 10930 0 1 8410
box -6 -8 26 248
use FILL  FILL_4__4878_
timestamp 0
transform 1 0 11370 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4879_
timestamp 0
transform 1 0 12030 0 1 9850
box -6 -8 26 248
use FILL  FILL_4__4880_
timestamp 0
transform -1 0 12090 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4881_
timestamp 0
transform -1 0 9130 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4882_
timestamp 0
transform 1 0 12050 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4883_
timestamp 0
transform 1 0 11870 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4884_
timestamp 0
transform 1 0 11690 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4885_
timestamp 0
transform -1 0 11730 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4886_
timestamp 0
transform 1 0 10990 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4887_
timestamp 0
transform 1 0 11030 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4__4888_
timestamp 0
transform 1 0 11690 0 1 8890
box -6 -8 26 248
use FILL  FILL_4__4889_
timestamp 0
transform 1 0 12030 0 1 9370
box -6 -8 26 248
use FILL  FILL_4__4890_
timestamp 0
transform 1 0 11550 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4891_
timestamp 0
transform 1 0 11890 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4__4893_
timestamp 0
transform -1 0 2530 0 -1 7450
box -6 -8 26 248
use FILL  FILL_4__4894_
timestamp 0
transform 1 0 9730 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4895_
timestamp 0
transform 1 0 8470 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4896_
timestamp 0
transform -1 0 9510 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4897_
timestamp 0
transform 1 0 9550 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4898_
timestamp 0
transform 1 0 9730 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4899_
timestamp 0
transform -1 0 9210 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4900_
timestamp 0
transform -1 0 9550 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4901_
timestamp 0
transform -1 0 9930 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4902_
timestamp 0
transform 1 0 10250 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4903_
timestamp 0
transform 1 0 9710 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4904_
timestamp 0
transform -1 0 10430 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4905_
timestamp 0
transform 1 0 9710 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4906_
timestamp 0
transform -1 0 9890 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4907_
timestamp 0
transform -1 0 9550 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4908_
timestamp 0
transform 1 0 10050 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4909_
timestamp 0
transform 1 0 10990 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4910_
timestamp 0
transform -1 0 11370 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4911_
timestamp 0
transform 1 0 11310 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4913_
timestamp 0
transform -1 0 10950 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4914_
timestamp 0
transform 1 0 11510 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4915_
timestamp 0
transform -1 0 10810 0 1 6970
box -6 -8 26 248
use FILL  FILL_4__4916_
timestamp 0
transform 1 0 10570 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4917_
timestamp 0
transform -1 0 10630 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4918_
timestamp 0
transform -1 0 10990 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4919_
timestamp 0
transform 1 0 11150 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4920_
timestamp 0
transform 1 0 8570 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4921_
timestamp 0
transform -1 0 8790 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4922_
timestamp 0
transform -1 0 8990 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4923_
timestamp 0
transform 1 0 9370 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4924_
timestamp 0
transform 1 0 9350 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4925_
timestamp 0
transform -1 0 9170 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4926_
timestamp 0
transform 1 0 8930 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4927_
timestamp 0
transform -1 0 11330 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4928_
timestamp 0
transform 1 0 11510 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4929_
timestamp 0
transform 1 0 12090 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4930_
timestamp 0
transform 1 0 11670 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4931_
timestamp 0
transform -1 0 11890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4933_
timestamp 0
transform -1 0 11170 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4934_
timestamp 0
transform 1 0 10950 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4935_
timestamp 0
transform -1 0 10770 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4936_
timestamp 0
transform -1 0 9670 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4937_
timestamp 0
transform -1 0 9890 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4938_
timestamp 0
transform 1 0 10050 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4939_
timestamp 0
transform 1 0 10130 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4940_
timestamp 0
transform 1 0 10230 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4__4941_
timestamp 0
transform 1 0 10330 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4942_
timestamp 0
transform -1 0 10730 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4943_
timestamp 0
transform 1 0 11710 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4944_
timestamp 0
transform -1 0 11930 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4945_
timestamp 0
transform 1 0 11870 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4946_
timestamp 0
transform -1 0 11850 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4947_
timestamp 0
transform -1 0 8670 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4948_
timestamp 0
transform 1 0 8990 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4949_
timestamp 0
transform 1 0 12110 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__4950_
timestamp 0
transform -1 0 12070 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4951_
timestamp 0
transform -1 0 8610 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4953_
timestamp 0
transform -1 0 8890 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4954_
timestamp 0
transform -1 0 9190 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4955_
timestamp 0
transform -1 0 8750 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__4956_
timestamp 0
transform -1 0 8830 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4957_
timestamp 0
transform -1 0 8690 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4958_
timestamp 0
transform -1 0 11070 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4959_
timestamp 0
transform 1 0 11250 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4960_
timestamp 0
transform -1 0 11470 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4961_
timestamp 0
transform 1 0 11650 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4962_
timestamp 0
transform 1 0 12050 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4963_
timestamp 0
transform 1 0 12010 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4964_
timestamp 0
transform 1 0 12010 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4965_
timestamp 0
transform -1 0 11850 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4966_
timestamp 0
transform -1 0 9190 0 1 4090
box -6 -8 26 248
use FILL  FILL_4__4967_
timestamp 0
transform 1 0 8110 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__4968_
timestamp 0
transform 1 0 11690 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4969_
timestamp 0
transform 1 0 12050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4970_
timestamp 0
transform 1 0 9090 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4971_
timestamp 0
transform -1 0 8310 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4973_
timestamp 0
transform -1 0 8870 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4974_
timestamp 0
transform 1 0 8770 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4975_
timestamp 0
transform 1 0 8970 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4976_
timestamp 0
transform 1 0 11630 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4977_
timestamp 0
transform 1 0 11430 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4978_
timestamp 0
transform 1 0 11450 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4979_
timestamp 0
transform 1 0 11470 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4980_
timestamp 0
transform 1 0 11850 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4981_
timestamp 0
transform -1 0 11850 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4982_
timestamp 0
transform -1 0 11870 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4983_
timestamp 0
transform 1 0 11650 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4984_
timestamp 0
transform 1 0 11270 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4985_
timestamp 0
transform -1 0 8090 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4986_
timestamp 0
transform 1 0 9130 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4987_
timestamp 0
transform 1 0 11650 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4988_
timestamp 0
transform -1 0 11870 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4989_
timestamp 0
transform -1 0 11470 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4990_
timestamp 0
transform -1 0 11290 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__4991_
timestamp 0
transform 1 0 11670 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__4993_
timestamp 0
transform 1 0 11310 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__4994_
timestamp 0
transform 1 0 9330 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__4995_
timestamp 0
transform -1 0 9910 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4996_
timestamp 0
transform 1 0 9270 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4997_
timestamp 0
transform -1 0 9350 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__4998_
timestamp 0
transform 1 0 9450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__4999_
timestamp 0
transform -1 0 9310 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5000_
timestamp 0
transform 1 0 11050 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__5001_
timestamp 0
transform -1 0 10870 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__5002_
timestamp 0
transform -1 0 10690 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5003_
timestamp 0
transform -1 0 10750 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5004_
timestamp 0
transform 1 0 10930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5005_
timestamp 0
transform -1 0 10910 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5006_
timestamp 0
transform 1 0 11430 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5007_
timestamp 0
transform 1 0 12030 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5008_
timestamp 0
transform 1 0 12010 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__5009_
timestamp 0
transform 1 0 12030 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5010_
timestamp 0
transform -1 0 11330 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__5011_
timestamp 0
transform 1 0 11830 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5013_
timestamp 0
transform -1 0 10310 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5014_
timestamp 0
transform -1 0 9530 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5015_
timestamp 0
transform 1 0 8290 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5016_
timestamp 0
transform 1 0 10690 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5017_
timestamp 0
transform 1 0 8950 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5018_
timestamp 0
transform 1 0 8490 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5019_
timestamp 0
transform 1 0 9170 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5020_
timestamp 0
transform 1 0 9070 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5021_
timestamp 0
transform 1 0 9350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5022_
timestamp 0
transform -1 0 9150 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5023_
timestamp 0
transform -1 0 10870 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__5024_
timestamp 0
transform 1 0 10870 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5025_
timestamp 0
transform -1 0 11090 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5026_
timestamp 0
transform 1 0 11110 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__5027_
timestamp 0
transform -1 0 10910 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5028_
timestamp 0
transform -1 0 10730 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5029_
timestamp 0
transform 1 0 11070 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5030_
timestamp 0
transform 1 0 11090 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5031_
timestamp 0
transform 1 0 11850 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__5033_
timestamp 0
transform -1 0 9010 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__5034_
timestamp 0
transform -1 0 9210 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__5035_
timestamp 0
transform 1 0 11230 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5036_
timestamp 0
transform 1 0 9910 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5037_
timestamp 0
transform 1 0 9710 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5038_
timestamp 0
transform 1 0 9550 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5039_
timestamp 0
transform 1 0 9490 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5040_
timestamp 0
transform 1 0 9730 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5041_
timestamp 0
transform 1 0 9930 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5042_
timestamp 0
transform 1 0 10650 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__5043_
timestamp 0
transform 1 0 10470 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5044_
timestamp 0
transform 1 0 10530 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5045_
timestamp 0
transform -1 0 10510 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5046_
timestamp 0
transform 1 0 10950 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__5047_
timestamp 0
transform 1 0 11050 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5048_
timestamp 0
transform 1 0 11490 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__5049_
timestamp 0
transform -1 0 11330 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__5050_
timestamp 0
transform -1 0 9390 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__5051_
timestamp 0
transform 1 0 8390 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__5053_
timestamp 0
transform -1 0 10790 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__5054_
timestamp 0
transform -1 0 10430 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__5055_
timestamp 0
transform 1 0 8550 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__5056_
timestamp 0
transform 1 0 8170 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__5057_
timestamp 0
transform 1 0 8390 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__5058_
timestamp 0
transform -1 0 8210 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__5059_
timestamp 0
transform 1 0 8030 0 1 6490
box -6 -8 26 248
use FILL  FILL_4__5060_
timestamp 0
transform -1 0 7670 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__5061_
timestamp 0
transform -1 0 7850 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__5062_
timestamp 0
transform 1 0 8010 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4__5063_
timestamp 0
transform -1 0 8050 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__5064_
timestamp 0
transform -1 0 7570 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5065_
timestamp 0
transform -1 0 7770 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5066_
timestamp 0
transform -1 0 7710 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5067_
timestamp 0
transform -1 0 8410 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5068_
timestamp 0
transform -1 0 8430 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5069_
timestamp 0
transform -1 0 8270 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5070_
timestamp 0
transform -1 0 7890 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5071_
timestamp 0
transform 1 0 8070 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5073_
timestamp 0
transform 1 0 7330 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5074_
timestamp 0
transform 1 0 4890 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4__5075_
timestamp 0
transform 1 0 10290 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__5076_
timestamp 0
transform 1 0 10090 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__5077_
timestamp 0
transform 1 0 9870 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__5078_
timestamp 0
transform 1 0 9650 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__5079_
timestamp 0
transform 1 0 10050 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__5080_
timestamp 0
transform 1 0 10250 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__5081_
timestamp 0
transform 1 0 10470 0 1 6010
box -6 -8 26 248
use FILL  FILL_4__5082_
timestamp 0
transform 1 0 10450 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4__5083_
timestamp 0
transform -1 0 10350 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5084_
timestamp 0
transform -1 0 9730 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5085_
timestamp 0
transform 1 0 8570 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5086_
timestamp 0
transform -1 0 8770 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5087_
timestamp 0
transform -1 0 10930 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__5088_
timestamp 0
transform -1 0 10710 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__5089_
timestamp 0
transform -1 0 10510 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__5090_
timestamp 0
transform -1 0 10290 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5091_
timestamp 0
transform 1 0 10130 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4__5093_
timestamp 0
transform -1 0 10150 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__5094_
timestamp 0
transform 1 0 10290 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__5095_
timestamp 0
transform -1 0 9810 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__5096_
timestamp 0
transform 1 0 8950 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__5097_
timestamp 0
transform 1 0 8270 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4__5098_
timestamp 0
transform 1 0 9770 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5099_
timestamp 0
transform 1 0 9950 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5100_
timestamp 0
transform 1 0 9390 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5101_
timestamp 0
transform -1 0 10110 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5102_
timestamp 0
transform -1 0 9930 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5103_
timestamp 0
transform 1 0 10070 0 1 5050
box -6 -8 26 248
use FILL  FILL_4__5104_
timestamp 0
transform -1 0 10370 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5105_
timestamp 0
transform -1 0 10170 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5106_
timestamp 0
transform -1 0 10550 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5107_
timestamp 0
transform 1 0 10530 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__5108_
timestamp 0
transform -1 0 11130 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__5109_
timestamp 0
transform 1 0 10730 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4__5110_
timestamp 0
transform -1 0 9590 0 1 4570
box -6 -8 26 248
use FILL  FILL_4__5111_
timestamp 0
transform -1 0 7950 0 1 5530
box -6 -8 26 248
use FILL  FILL_4__5124_
timestamp 0
transform 1 0 1810 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__5125_
timestamp 0
transform -1 0 670 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__5126_
timestamp 0
transform -1 0 850 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__5127_
timestamp 0
transform 1 0 810 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__5128_
timestamp 0
transform 1 0 570 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__5129_
timestamp 0
transform 1 0 1010 0 1 2170
box -6 -8 26 248
use FILL  FILL_4__5130_
timestamp 0
transform 1 0 1010 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__5131_
timestamp 0
transform -1 0 2330 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5132_
timestamp 0
transform -1 0 5570 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5133_
timestamp 0
transform 1 0 5310 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__5134_
timestamp 0
transform 1 0 1390 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__5135_
timestamp 0
transform 1 0 2190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__5136_
timestamp 0
transform 1 0 1990 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__5137_
timestamp 0
transform -1 0 1130 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__5138_
timestamp 0
transform -1 0 1310 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__5139_
timestamp 0
transform -1 0 3690 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5140_
timestamp 0
transform 1 0 4150 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__5141_
timestamp 0
transform -1 0 4330 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__5142_
timestamp 0
transform -1 0 4210 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__5144_
timestamp 0
transform 1 0 5590 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5145_
timestamp 0
transform -1 0 4130 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5146_
timestamp 0
transform -1 0 4650 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5147_
timestamp 0
transform 1 0 4750 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5148_
timestamp 0
transform 1 0 4950 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5149_
timestamp 0
transform 1 0 5470 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__5150_
timestamp 0
transform -1 0 6090 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__5151_
timestamp 0
transform 1 0 3470 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5152_
timestamp 0
transform 1 0 5730 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5153_
timestamp 0
transform 1 0 4210 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__5154_
timestamp 0
transform 1 0 5410 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5155_
timestamp 0
transform 1 0 5370 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5156_
timestamp 0
transform 1 0 5530 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5157_
timestamp 0
transform 1 0 5670 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__5158_
timestamp 0
transform 1 0 4550 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5159_
timestamp 0
transform -1 0 4670 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5160_
timestamp 0
transform 1 0 4990 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5161_
timestamp 0
transform 1 0 4830 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5162_
timestamp 0
transform 1 0 5870 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__5164_
timestamp 0
transform 1 0 5890 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5165_
timestamp 0
transform -1 0 3830 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__5166_
timestamp 0
transform 1 0 4270 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5167_
timestamp 0
transform 1 0 4230 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5168_
timestamp 0
transform -1 0 4050 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5169_
timestamp 0
transform 1 0 2730 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__5170_
timestamp 0
transform 1 0 3850 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5171_
timestamp 0
transform -1 0 4150 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__5172_
timestamp 0
transform -1 0 3650 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__5173_
timestamp 0
transform -1 0 4930 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__5174_
timestamp 0
transform -1 0 3830 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__5175_
timestamp 0
transform 1 0 3670 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5176_
timestamp 0
transform -1 0 2670 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__5177_
timestamp 0
transform 1 0 3110 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__5178_
timestamp 0
transform 1 0 4450 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5179_
timestamp 0
transform 1 0 4470 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5180_
timestamp 0
transform 1 0 4270 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5181_
timestamp 0
transform 1 0 3270 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__5182_
timestamp 0
transform -1 0 2470 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__5184_
timestamp 0
transform -1 0 2490 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__5185_
timestamp 0
transform -1 0 4050 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__5186_
timestamp 0
transform -1 0 3330 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__5187_
timestamp 0
transform -1 0 3070 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__5188_
timestamp 0
transform 1 0 3770 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__5189_
timestamp 0
transform -1 0 3710 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5190_
timestamp 0
transform 1 0 3250 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__5191_
timestamp 0
transform 1 0 2930 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5192_
timestamp 0
transform -1 0 3650 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__5193_
timestamp 0
transform 1 0 6090 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5194_
timestamp 0
transform -1 0 2950 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__5195_
timestamp 0
transform -1 0 2870 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__5196_
timestamp 0
transform 1 0 3610 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__5197_
timestamp 0
transform -1 0 3530 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5198_
timestamp 0
transform -1 0 2930 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5199_
timestamp 0
transform 1 0 2490 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5200_
timestamp 0
transform -1 0 2710 0 -1 730
box -6 -8 26 248
use FILL  FILL_4__5201_
timestamp 0
transform -1 0 3990 0 1 1690
box -6 -8 26 248
use FILL  FILL_4__5202_
timestamp 0
transform 1 0 3950 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5203_
timestamp 0
transform -1 0 3490 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5205_
timestamp 0
transform -1 0 3950 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__5206_
timestamp 0
transform -1 0 3290 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5207_
timestamp 0
transform 1 0 2510 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5208_
timestamp 0
transform 1 0 3050 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__5209_
timestamp 0
transform -1 0 4510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4__5210_
timestamp 0
transform 1 0 2710 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5211_
timestamp 0
transform 1 0 2870 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5212_
timestamp 0
transform 1 0 3450 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__5213_
timestamp 0
transform 1 0 3330 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5214_
timestamp 0
transform -1 0 3090 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5215_
timestamp 0
transform 1 0 2310 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5216_
timestamp 0
transform -1 0 3110 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__5217_
timestamp 0
transform -1 0 6270 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5218_
timestamp 0
transform 1 0 3450 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__5219_
timestamp 0
transform 1 0 3610 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__5220_
timestamp 0
transform 1 0 4790 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__5221_
timestamp 0
transform 1 0 4610 0 -1 250
box -6 -8 26 248
use FILL  FILL_4__5222_
timestamp 0
transform -1 0 4090 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5223_
timestamp 0
transform 1 0 3130 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5225_
timestamp 0
transform 1 0 5390 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__5226_
timestamp 0
transform 1 0 5170 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5227_
timestamp 0
transform -1 0 5350 0 1 250
box -6 -8 26 248
use FILL  FILL_4__5228_
timestamp 0
transform -1 0 4790 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4__5229_
timestamp 0
transform -1 0 4830 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5230_
timestamp 0
transform 1 0 5010 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5231_
timestamp 0
transform 1 0 5210 0 1 730
box -6 -8 26 248
use FILL  FILL_4__5232_
timestamp 0
transform 1 0 4010 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4__5233_
timestamp 0
transform 1 0 4390 0 1 1210
box -6 -8 26 248
use FILL  FILL_4__5234_
timestamp 0
transform -1 0 5190 0 1 1210
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert0
timestamp 0
transform -1 0 4230 0 1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert1
timestamp 0
transform 1 0 6150 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert2
timestamp 0
transform -1 0 3330 0 1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert3
timestamp 0
transform -1 0 3710 0 1 9850
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert4
timestamp 0
transform 1 0 9490 0 1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert5
timestamp 0
transform 1 0 11290 0 1 8410
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert6
timestamp 0
transform -1 0 9490 0 1 8410
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert7
timestamp 0
transform 1 0 12030 0 1 7930
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert8
timestamp 0
transform -1 0 7190 0 1 5530
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert10
timestamp 0
transform 1 0 8730 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert11
timestamp 0
transform 1 0 6890 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert12
timestamp 0
transform 1 0 8930 0 1 9850
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert13
timestamp 0
transform 1 0 7410 0 1 9850
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert14
timestamp 0
transform 1 0 670 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert15
timestamp 0
transform 1 0 90 0 1 9370
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert16
timestamp 0
transform 1 0 1910 0 1 5530
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert17
timestamp 0
transform -1 0 9170 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert18
timestamp 0
transform -1 0 11530 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert19
timestamp 0
transform 1 0 10690 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert20
timestamp 0
transform -1 0 9210 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert21
timestamp 0
transform 1 0 2550 0 1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert22
timestamp 0
transform -1 0 1290 0 1 11290
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert23
timestamp 0
transform -1 0 1470 0 1 11290
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert24
timestamp 0
transform -1 0 1670 0 1 10330
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert38
timestamp 0
transform -1 0 11550 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert39
timestamp 0
transform -1 0 10690 0 1 6010
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert40
timestamp 0
transform 1 0 12050 0 1 6970
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert41
timestamp 0
transform -1 0 11270 0 1 6010
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert42
timestamp 0
transform 1 0 11470 0 1 730
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert43
timestamp 0
transform -1 0 11030 0 1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert44
timestamp 0
transform -1 0 10510 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert45
timestamp 0
transform -1 0 11390 0 1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert46
timestamp 0
transform -1 0 10770 0 1 3130
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert47
timestamp 0
transform 1 0 6230 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert48
timestamp 0
transform -1 0 4790 0 1 1690
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert50
timestamp 0
transform -1 0 10430 0 1 1690
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert51
timestamp 0
transform 1 0 8190 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert52
timestamp 0
transform 1 0 10050 0 1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert53
timestamp 0
transform 1 0 9210 0 1 4570
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert54
timestamp 0
transform 1 0 9030 0 1 4570
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert55
timestamp 0
transform -1 0 9570 0 1 4090
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert56
timestamp 0
transform -1 0 8870 0 1 4570
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert57
timestamp 0
transform 1 0 11490 0 1 3130
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert58
timestamp 0
transform 1 0 10670 0 -1 730
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert59
timestamp 0
transform -1 0 7750 0 -1 730
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert60
timestamp 0
transform 1 0 11830 0 -1 730
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert61
timestamp 0
transform 1 0 11930 0 1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert62
timestamp 0
transform -1 0 4830 0 1 2170
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert63
timestamp 0
transform -1 0 9350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert64
timestamp 0
transform -1 0 11690 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert65
timestamp 0
transform -1 0 9350 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert66
timestamp 0
transform -1 0 11530 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert67
timestamp 0
transform 1 0 6950 0 1 11290
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert68
timestamp 0
transform -1 0 3190 0 -1 10330
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert70
timestamp 0
transform 1 0 5130 0 -1 11290
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert71
timestamp 0
transform -1 0 3590 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert72
timestamp 0
transform 1 0 7130 0 1 11290
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert73
timestamp 0
transform 1 0 7150 0 1 730
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert74
timestamp 0
transform -1 0 6490 0 1 2170
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert75
timestamp 0
transform 1 0 7110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert76
timestamp 0
transform 1 0 6570 0 1 730
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert77
timestamp 0
transform 1 0 10290 0 1 4090
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert78
timestamp 0
transform 1 0 9150 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert79
timestamp 0
transform 1 0 10310 0 1 730
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert80
timestamp 0
transform -1 0 4970 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert81
timestamp 0
transform -1 0 2830 0 1 5530
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert82
timestamp 0
transform -1 0 4050 0 -1 5530
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert83
timestamp 0
transform -1 0 6310 0 1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert84
timestamp 0
transform 1 0 7370 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert85
timestamp 0
transform -1 0 3290 0 1 8410
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert86
timestamp 0
transform 1 0 3990 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert87
timestamp 0
transform -1 0 3250 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert88
timestamp 0
transform 1 0 7910 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert90
timestamp 0
transform 1 0 5590 0 1 9370
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert91
timestamp 0
transform 1 0 9050 0 1 10330
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert92
timestamp 0
transform -1 0 8550 0 1 10810
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert93
timestamp 0
transform -1 0 10950 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert94
timestamp 0
transform 1 0 7290 0 1 10330
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert95
timestamp 0
transform 1 0 11550 0 1 10810
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert96
timestamp 0
transform -1 0 5010 0 1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert97
timestamp 0
transform 1 0 630 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert98
timestamp 0
transform -1 0 4030 0 1 7930
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert99
timestamp 0
transform 1 0 570 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert100
timestamp 0
transform 1 0 3050 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert101
timestamp 0
transform -1 0 510 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert102
timestamp 0
transform 1 0 3750 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert103
timestamp 0
transform -1 0 3670 0 1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert104
timestamp 0
transform 1 0 4650 0 1 10330
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert105
timestamp 0
transform 1 0 310 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert106
timestamp 0
transform 1 0 6530 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert107
timestamp 0
transform -1 0 6230 0 1 730
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert108
timestamp 0
transform 1 0 5710 0 1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert110
timestamp 0
transform -1 0 5350 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert111
timestamp 0
transform 1 0 7310 0 1 1690
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert112
timestamp 0
transform 1 0 10690 0 1 11770
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert113
timestamp 0
transform -1 0 12130 0 1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert114
timestamp 0
transform -1 0 10330 0 -1 1210
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert115
timestamp 0
transform 1 0 7390 0 1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert116
timestamp 0
transform -1 0 5530 0 1 2170
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert117
timestamp 0
transform -1 0 5510 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert118
timestamp 0
transform -1 0 11210 0 1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert119
timestamp 0
transform 1 0 10390 0 1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert120
timestamp 0
transform -1 0 11130 0 1 730
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert121
timestamp 0
transform -1 0 8190 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert122
timestamp 0
transform 1 0 11210 0 1 2170
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert123
timestamp 0
transform -1 0 10050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert124
timestamp 0
transform -1 0 8030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert125
timestamp 0
transform -1 0 5350 0 1 2170
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert126
timestamp 0
transform 1 0 12030 0 -1 4570
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert127
timestamp 0
transform 1 0 10790 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert128
timestamp 0
transform -1 0 12070 0 -1 4090
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert130
timestamp 0
transform 1 0 12030 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert131
timestamp 0
transform -1 0 9390 0 1 4090
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert132
timestamp 0
transform -1 0 8730 0 1 730
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert133
timestamp 0
transform 1 0 12030 0 1 730
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert134
timestamp 0
transform -1 0 11410 0 1 4090
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert135
timestamp 0
transform -1 0 9130 0 -1 250
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert136
timestamp 0
transform 1 0 9490 0 -1 250
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert137
timestamp 0
transform -1 0 6410 0 1 730
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert138
timestamp 0
transform 1 0 8390 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert139
timestamp 0
transform -1 0 6430 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert140
timestamp 0
transform 1 0 9450 0 1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert141
timestamp 0
transform -1 0 7070 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert142
timestamp 0
transform -1 0 7050 0 1 8410
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert143
timestamp 0
transform -1 0 6470 0 -1 6970
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert144
timestamp 0
transform -1 0 6290 0 1 6970
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert145
timestamp 0
transform 1 0 9570 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert146
timestamp 0
transform 1 0 9670 0 1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert147
timestamp 0
transform -1 0 7750 0 1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert148
timestamp 0
transform -1 0 7670 0 -1 7930
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert150
timestamp 0
transform -1 0 7250 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert151
timestamp 0
transform 1 0 7350 0 -1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert152
timestamp 0
transform -1 0 8250 0 1 9370
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert153
timestamp 0
transform 1 0 10090 0 -1 9850
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert154
timestamp 0
transform 1 0 10770 0 -1 8410
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert155
timestamp 0
transform 1 0 6410 0 1 3130
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert156
timestamp 0
transform 1 0 9150 0 -1 3130
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert157
timestamp 0
transform -1 0 5890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert158
timestamp 0
transform 1 0 9890 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert159
timestamp 0
transform 1 0 8750 0 -1 1690
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert160
timestamp 0
transform 1 0 10390 0 1 9850
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert161
timestamp 0
transform 1 0 9290 0 1 9850
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert162
timestamp 0
transform 1 0 10250 0 1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert163
timestamp 0
transform -1 0 8350 0 1 8890
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert164
timestamp 0
transform 1 0 11750 0 1 4090
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert165
timestamp 0
transform -1 0 8810 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert166
timestamp 0
transform -1 0 11590 0 1 4090
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert167
timestamp 0
transform 1 0 11750 0 1 11770
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert168
timestamp 0
transform -1 0 11330 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4_BUFX2_insert169
timestamp 0
transform 1 0 4950 0 1 1690
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert25
timestamp 0
transform 1 0 1390 0 1 2170
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert26
timestamp 0
transform 1 0 4050 0 -1 2170
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert27
timestamp 0
transform -1 0 110 0 -1 2650
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert28
timestamp 0
transform -1 0 2750 0 1 9370
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert30
timestamp 0
transform 1 0 6210 0 -1 5050
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert31
timestamp 0
transform 1 0 810 0 -1 6010
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert32
timestamp 0
transform -1 0 4850 0 -1 3610
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert33
timestamp 0
transform -1 0 990 0 -1 10810
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert34
timestamp 0
transform 1 0 1430 0 -1 6490
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert35
timestamp 0
transform -1 0 350 0 -1 11770
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert36
timestamp 0
transform 1 0 90 0 1 5530
box -6 -8 26 248
use FILL  FILL_4_CLKBUF1_insert37
timestamp 0
transform 1 0 6170 0 1 11770
box -6 -8 26 248
<< labels >>
flabel metal1 s 12222 2 12282 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 5997 12057 6003 12063 3 FreeSans 16 90 0 0 clk
port 2 nsew
flabel metal3 s -24 2336 -16 2344 7 FreeSans 16 0 0 0 reset
port 3 nsew
flabel metal3 s -24 3716 -16 3724 7 FreeSans 16 0 0 0 AB[15]
port 4 nsew
flabel metal3 s -24 2756 -16 2764 7 FreeSans 16 0 0 0 AB[14]
port 5 nsew
flabel metal2 s 1997 -23 2003 -17 7 FreeSans 16 270 0 0 AB[13]
port 6 nsew
flabel metal2 s 2817 -23 2823 -17 7 FreeSans 16 270 0 0 AB[12]
port 7 nsew
flabel metal3 s -24 4916 -16 4924 7 FreeSans 16 0 0 0 AB[11]
port 8 nsew
flabel metal3 s -24 5396 -16 5404 7 FreeSans 16 0 0 0 AB[10]
port 9 nsew
flabel metal2 s 2177 -23 2183 -17 7 FreeSans 16 270 0 0 AB[9]
port 10 nsew
flabel metal2 s 4017 -23 4023 -17 7 FreeSans 16 270 0 0 AB[8]
port 11 nsew
flabel metal3 s 12256 2756 12264 2764 3 FreeSans 16 0 0 0 AB[7]
port 12 nsew
flabel metal2 s 6697 -23 6703 -17 7 FreeSans 16 270 0 0 AB[6]
port 13 nsew
flabel metal2 s 6857 -23 6863 -17 7 FreeSans 16 270 0 0 AB[5]
port 14 nsew
flabel metal3 s 12256 2996 12264 3004 3 FreeSans 16 0 0 0 AB[4]
port 15 nsew
flabel metal3 s 12256 3216 12264 3224 3 FreeSans 16 0 0 0 AB[3]
port 16 nsew
flabel metal2 s 6517 -23 6523 -17 7 FreeSans 16 270 0 0 AB[2]
port 17 nsew
flabel metal3 s 12256 3256 12264 3264 3 FreeSans 16 0 0 0 AB[1]
port 18 nsew
flabel metal2 s 11997 -23 12003 -17 7 FreeSans 16 270 0 0 AB[0]
port 19 nsew
flabel metal2 s 5157 -23 5163 -17 7 FreeSans 16 270 0 0 DI[7]
port 20 nsew
flabel metal2 s 6117 -23 6123 -17 7 FreeSans 16 270 0 0 DI[6]
port 21 nsew
flabel metal2 s 3117 -23 3123 -17 7 FreeSans 16 270 0 0 DI[5]
port 22 nsew
flabel metal2 s 3817 -23 3823 -17 7 FreeSans 16 270 0 0 DI[4]
port 23 nsew
flabel metal2 s 3617 -23 3623 -17 7 FreeSans 16 270 0 0 DI[3]
port 24 nsew
flabel metal2 s 4137 -23 4143 -17 7 FreeSans 16 270 0 0 DI[2]
port 25 nsew
flabel metal2 s 3457 -23 3463 -17 7 FreeSans 16 270 0 0 DI[1]
port 26 nsew
flabel metal2 s 4837 -23 4843 -17 7 FreeSans 16 270 0 0 DI[0]
port 27 nsew
flabel metal3 s -24 6116 -16 6124 7 FreeSans 16 0 0 0 DO[7]
port 28 nsew
flabel metal3 s -24 2276 -16 2284 7 FreeSans 16 0 0 0 DO[6]
port 29 nsew
flabel metal3 s -24 4196 -16 4204 7 FreeSans 16 0 0 0 DO[5]
port 30 nsew
flabel metal2 s 4437 -23 4443 -17 7 FreeSans 16 270 0 0 DO[4]
port 31 nsew
flabel metal2 s 4537 -23 4543 -17 7 FreeSans 16 270 0 0 DO[3]
port 32 nsew
flabel metal2 s 3337 -23 3343 -17 7 FreeSans 16 270 0 0 DO[2]
port 33 nsew
flabel metal3 s -24 2996 -16 3004 7 FreeSans 16 0 0 0 DO[1]
port 34 nsew
flabel metal2 s 3717 -23 3723 -17 7 FreeSans 16 270 0 0 DO[0]
port 35 nsew
flabel metal3 s -24 6356 -16 6364 7 FreeSans 16 0 0 0 WE
port 36 nsew
flabel metal2 s 1257 12057 1263 12063 3 FreeSans 16 90 0 0 IRQ
port 37 nsew
flabel metal3 s -24 10456 -16 10464 7 FreeSans 16 0 0 0 NMI
port 38 nsew
flabel metal3 s -24 9456 -16 9464 7 FreeSans 16 0 0 0 RDY
port 39 nsew
flabel metal3 s -24 356 -16 364 7 FreeSans 16 0 0 0 kbd_rdy
port 40 nsew
flabel metal3 s -24 116 -16 124 7 FreeSans 16 0 0 0 kbd_ack
port 41 nsew
flabel metal2 s 1817 -23 1823 -17 7 FreeSans 16 270 0 0 kbd_data[6]
port 42 nsew
flabel metal2 s 2117 -23 2123 -17 7 FreeSans 16 270 0 0 kbd_data[5]
port 43 nsew
flabel metal2 s 997 -23 1003 -17 7 FreeSans 16 270 0 0 kbd_data[4]
port 44 nsew
flabel metal2 s 1917 -23 1923 -17 7 FreeSans 16 270 0 0 kbd_data[3]
port 45 nsew
flabel metal2 s 297 -23 303 -17 7 FreeSans 16 270 0 0 kbd_data[2]
port 46 nsew
flabel metal2 s 1757 -23 1763 -17 7 FreeSans 16 270 0 0 kbd_data[1]
port 47 nsew
flabel metal2 s 2317 -23 2323 -17 7 FreeSans 16 270 0 0 kbd_data[0]
port 48 nsew
flabel metal2 s 4637 -23 4643 -17 7 FreeSans 16 270 0 0 dsp_rdy
port 49 nsew
flabel metal2 s 4677 -23 4683 -17 7 FreeSans 16 270 0 0 dsp_ack
port 50 nsew
flabel metal2 s 5197 -23 5203 -17 7 FreeSans 16 270 0 0 dsp_data[6]
port 51 nsew
flabel metal2 s 2597 -23 2603 -17 7 FreeSans 16 270 0 0 dsp_data[5]
port 52 nsew
flabel metal2 s 3897 -23 3903 -17 7 FreeSans 16 270 0 0 dsp_data[4]
port 53 nsew
flabel metal2 s 3497 -23 3503 -17 7 FreeSans 16 270 0 0 dsp_data[3]
port 54 nsew
flabel metal2 s 4297 -23 4303 -17 7 FreeSans 16 270 0 0 dsp_data[2]
port 55 nsew
flabel metal2 s 3157 -23 3163 -17 7 FreeSans 16 270 0 0 dsp_data[1]
port 56 nsew
flabel metal2 s 4997 -23 5003 -17 7 FreeSans 16 270 0 0 dsp_data[0]
port 57 nsew
<< properties >>
string FIXED_BBOX -40 -40 12260 12060
<< end >>
