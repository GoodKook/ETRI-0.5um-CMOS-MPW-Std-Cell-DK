magic
tech scmos
magscale 1 2
timestamp 1727572430
<< nwell >>
rect -12 154 112 272
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
rect 60 14 64 54
<< ptransistor >>
rect 22 166 26 246
rect 36 166 40 246
rect 56 206 60 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 42 40 54
rect 24 14 26 42
rect 38 14 40 42
rect 44 14 46 54
rect 58 14 60 54
rect 64 14 66 54
<< pdiffusion >>
rect 20 166 22 246
rect 26 166 36 246
rect 40 206 42 246
rect 54 206 56 246
rect 60 206 62 246
rect 40 166 51 206
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 42
rect 46 14 58 54
rect 66 14 78 54
<< pdcontact >>
rect 8 166 20 246
rect 42 206 54 246
rect 62 206 74 246
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 254 106 266
<< polysilicon >>
rect 22 246 26 250
rect 36 246 40 250
rect 56 246 60 250
rect 22 162 26 166
rect 12 157 26 162
rect 36 162 40 166
rect 56 162 60 206
rect 36 157 44 162
rect 56 157 66 162
rect 12 129 16 157
rect 40 123 44 157
rect 12 66 16 117
rect 36 111 44 123
rect 12 59 24 66
rect 20 54 24 59
rect 40 54 44 111
rect 60 123 66 157
rect 60 54 64 123
rect 20 10 24 14
rect 40 10 44 14
rect 60 10 64 14
<< polycontact >>
rect 4 117 16 129
rect 24 111 36 123
rect 64 111 76 123
<< metal1 >>
rect -6 266 106 268
rect -6 252 106 254
rect 8 246 20 252
rect 62 246 74 252
rect 43 117 51 206
rect 49 75 57 103
rect 49 68 74 75
rect 6 54 58 57
rect 18 48 46 54
rect 66 54 74 68
rect 26 8 38 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m2contact >>
rect 23 123 37 137
rect 3 103 17 117
rect 63 123 77 137
rect 43 103 57 117
<< metal2 >>
rect 23 137 37 157
rect 63 137 77 157
rect 3 83 17 103
rect 43 83 57 103
<< m2p >>
rect 23 143 37 157
rect 63 143 77 157
rect 3 83 17 97
rect 43 83 57 97
<< labels >>
rlabel metal2 3 83 17 97 0 A
port 0 nsew signal input
rlabel metal2 23 143 37 157 0 B
port 1 nsew signal input
rlabel metal2 63 143 77 157 0 C
port 2 nsew signal input
rlabel metal2 43 83 57 97 0 Y
port 3 nsew signal output
rlabel metal1 -6 252 106 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -6 -8 106 8 0 gnd
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
