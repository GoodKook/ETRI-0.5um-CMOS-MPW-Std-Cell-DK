magic
tech scmos
magscale 1 2
timestamp 1728304996
<< nwell >>
rect -12 134 92 252
<< ntransistor >>
rect 23 14 27 54
rect 33 14 37 54
<< ptransistor >>
rect 21 186 25 226
rect 41 186 45 226
<< ndiffusion >>
rect 21 14 23 54
rect 27 14 33 54
rect 37 14 39 54
<< pdiffusion >>
rect 19 186 21 226
rect 25 186 27 226
rect 39 186 41 226
rect 45 186 47 226
<< ndcontact >>
rect 9 14 21 54
rect 39 14 51 54
<< pdcontact >>
rect 7 186 19 226
rect 27 186 39 226
rect 47 186 59 226
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 234 86 246
<< polysilicon >>
rect 21 226 25 230
rect 41 226 45 230
rect 21 109 25 186
rect 16 97 25 109
rect 19 81 25 97
rect 41 109 45 186
rect 41 97 44 109
rect 41 81 47 97
rect 19 74 27 81
rect 23 54 27 74
rect 33 74 47 81
rect 33 54 37 74
rect 23 10 27 14
rect 33 10 37 14
<< polycontact >>
rect 4 97 16 109
rect 44 97 56 109
<< metal1 >>
rect -6 246 86 248
rect -6 232 86 234
rect 7 226 19 232
rect 47 226 59 232
rect 27 131 35 186
rect 27 68 35 117
rect 27 62 51 68
rect 39 54 51 62
rect 9 8 21 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m2contact >>
rect 3 109 17 123
rect 23 117 37 131
rect 43 109 57 123
<< metal2 >>
rect 3 123 17 137
rect 23 103 37 117
rect 43 123 57 137
<< m1p >>
rect -6 232 86 248
rect -6 -8 86 8
<< m2p >>
rect 3 123 17 137
rect 43 123 57 137
rect 23 103 37 117
<< labels >>
rlabel metal1 -6 -8 86 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 -6 232 86 248 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal2 3 123 17 137 0 A
port 0 nsew signal input
rlabel metal2 43 123 57 137 0 B
port 1 nsew signal input
rlabel metal2 23 103 37 117 0 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 80 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
