magic
tech scmos
magscale 1 6
timestamp 1537935238
<< checkpaint >>
rect -110 -155 374 298
<< metal1 >>
rect 10 132 254 178
rect 10 116 46 132
rect 114 116 150 132
rect 218 116 254 132
rect 62 -7 98 12
rect 166 -7 202 12
rect 62 -35 202 -7
use nmos4_CDNS_704676826055  nmos4_CDNS_704676826055_0
timestamp 1537935238
transform 1 0 0 0 1 0
box 10 4 254 168
<< end >>
