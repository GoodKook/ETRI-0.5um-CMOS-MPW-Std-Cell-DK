magic
tech scmos
magscale 1 2
timestamp 1718295485
<< error_s >>
rect 4 6244 6436 6256
rect 4 5984 6436 5996
rect 4 5724 6436 5736
rect 4 5464 6436 5476
rect 4 5204 6436 5216
rect 4 4944 6436 4956
rect 4 4684 6436 4696
rect 4 4424 6436 4436
rect 4 4164 6436 4176
rect 4 3904 6436 3916
rect 4 3644 6436 3656
rect 4 3384 6436 3396
rect 4 3124 6436 3136
rect 4 2864 6436 2876
rect 4 2604 6436 2616
rect 4 2344 6436 2356
rect 4 2084 6436 2096
rect 4 1824 6436 1836
rect 4 1564 6436 1576
rect 4 1304 6436 1316
rect 4 1044 6436 1056
rect 4 784 6436 796
rect 4 524 6436 536
rect 4 264 6436 276
rect 4 4 6436 16
<< nwell >>
rect 1556 4069 1563 4081
<< metal1 >>
rect -63 6242 30 6258
rect -63 5738 -3 6242
rect 3247 6173 3253 6187
rect 2367 6157 2433 6163
rect 3347 6157 3373 6163
rect 1987 6137 2013 6143
rect 2807 6137 2873 6143
rect 3187 6137 3293 6143
rect 4567 6137 4633 6143
rect 4947 6137 4973 6143
rect 6347 6137 6373 6143
rect 507 6123 520 6127
rect 3400 6123 3413 6127
rect 507 6113 523 6123
rect 517 6066 523 6113
rect 3397 6113 3413 6123
rect 3800 6123 3813 6127
rect 3797 6113 3813 6123
rect 6107 6123 6120 6127
rect 6107 6113 6123 6123
rect 3397 6087 3403 6113
rect 3797 6087 3803 6113
rect 3397 6077 3413 6087
rect 3400 6073 3413 6077
rect 3797 6077 3813 6087
rect 3800 6073 3813 6077
rect 6117 6083 6123 6113
rect 6117 6077 6153 6083
rect 1607 6057 1643 6063
rect 1637 6043 1643 6057
rect 1767 6057 1813 6063
rect 2527 6057 2613 6063
rect 3187 6057 3293 6063
rect 4187 6057 4253 6063
rect 1637 6037 1713 6043
rect 2607 6037 2673 6043
rect 2407 6017 2433 6023
rect 6443 5998 6503 6258
rect 6410 5982 6503 5998
rect 627 5957 673 5963
rect 4337 5937 4373 5943
rect 581 5917 593 5923
rect 2247 5917 2313 5923
rect 3707 5917 3753 5923
rect 337 5867 343 5913
rect 500 5903 513 5907
rect 497 5893 513 5903
rect 3867 5903 3880 5907
rect 4060 5903 4073 5907
rect 3867 5893 3883 5903
rect 497 5867 503 5893
rect 3877 5867 3883 5893
rect 4057 5893 4073 5903
rect 4337 5903 4343 5937
rect 4367 5917 4413 5923
rect 5187 5917 5333 5923
rect 4660 5903 4673 5907
rect 4337 5897 4363 5903
rect 4057 5867 4063 5893
rect 4357 5867 4363 5897
rect 4657 5893 4673 5903
rect 4657 5867 4663 5893
rect 327 5857 343 5867
rect 327 5853 340 5857
rect 487 5857 503 5867
rect 487 5853 500 5857
rect 3567 5857 3593 5863
rect 3867 5857 3883 5867
rect 3867 5853 3880 5857
rect 4047 5857 4063 5867
rect 4047 5853 4060 5857
rect 4347 5857 4363 5867
rect 4347 5853 4360 5857
rect 4647 5857 4663 5867
rect 4647 5853 4660 5857
rect 947 5837 999 5843
rect 1067 5837 1113 5843
rect 2227 5837 2293 5843
rect 2507 5837 2553 5843
rect 2647 5837 2753 5843
rect 3427 5837 3453 5843
rect 3847 5837 3953 5843
rect 847 5817 873 5823
rect 2173 5823 2187 5831
rect 2173 5820 2213 5823
rect 2177 5817 2213 5820
rect 3367 5817 3473 5823
rect -63 5722 30 5738
rect -63 5218 -3 5722
rect 1727 5657 1773 5663
rect 967 5637 1053 5643
rect 1747 5637 1773 5643
rect 3227 5637 3253 5643
rect 4647 5637 4693 5643
rect 527 5617 553 5623
rect 567 5617 593 5623
rect 1187 5617 1233 5623
rect 1427 5617 1493 5623
rect 3187 5617 3253 5623
rect 3517 5617 3573 5623
rect 160 5603 173 5607
rect 157 5593 173 5603
rect 3517 5603 3523 5617
rect 4127 5617 4173 5623
rect 6047 5617 6173 5623
rect 6280 5603 6293 5607
rect 3497 5597 3523 5603
rect 157 5563 163 5593
rect 3497 5567 3503 5597
rect 6277 5593 6293 5603
rect 6387 5603 6400 5607
rect 6387 5593 6403 5603
rect 6277 5567 6283 5593
rect 157 5560 183 5563
rect 157 5557 187 5560
rect 173 5547 187 5557
rect 3487 5557 3503 5567
rect 3487 5553 3500 5557
rect 6267 5557 6283 5567
rect 6267 5553 6280 5557
rect 1727 5537 1773 5543
rect 5687 5537 5753 5543
rect 6047 5537 6133 5543
rect 6397 5543 6403 5593
rect 6367 5537 6403 5543
rect 6443 5478 6503 5982
rect 6410 5462 6503 5478
rect 1947 5437 1973 5443
rect 940 5383 953 5387
rect 937 5373 953 5383
rect 1240 5383 1253 5387
rect 1237 5373 1253 5383
rect 1647 5383 1660 5387
rect 1647 5373 1663 5383
rect 1947 5377 1973 5383
rect 2913 5383 2927 5393
rect 2913 5380 2973 5383
rect 2917 5377 2973 5380
rect 5320 5383 5333 5387
rect 5317 5373 5333 5383
rect 6200 5383 6213 5387
rect 6197 5373 6213 5383
rect 937 5367 943 5373
rect 920 5366 943 5367
rect 927 5357 943 5366
rect 927 5353 940 5357
rect 1237 5343 1243 5373
rect 1207 5337 1243 5343
rect 1657 5347 1663 5373
rect 5317 5347 5323 5373
rect 1657 5337 1673 5347
rect 1660 5333 1673 5337
rect 3987 5337 4013 5343
rect 5307 5337 5323 5347
rect 6197 5347 6203 5373
rect 6197 5337 6213 5347
rect 5307 5333 5320 5337
rect 6200 5333 6213 5337
rect 1047 5317 1093 5323
rect 1447 5317 1553 5323
rect 1907 5317 1979 5323
rect 3427 5317 3453 5323
rect 3627 5317 3753 5323
rect 3927 5317 4013 5323
rect 4107 5317 4133 5323
rect 5547 5317 5613 5323
rect 5867 5317 5919 5323
rect 6027 5317 6073 5323
rect 2187 5297 2273 5303
rect 3273 5243 3287 5253
rect 3247 5240 3287 5243
rect 3247 5237 3283 5240
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 627 5117 663 5123
rect 167 5097 273 5103
rect 567 5097 633 5103
rect 487 5083 500 5087
rect 657 5083 663 5117
rect 2297 5117 2333 5123
rect 867 5097 953 5103
rect 1007 5097 1113 5103
rect 1307 5097 1333 5103
rect 487 5073 503 5083
rect 497 5047 503 5073
rect 637 5077 663 5083
rect 497 5037 513 5047
rect 500 5033 513 5037
rect 637 5026 643 5077
rect 1447 5083 1460 5087
rect 1720 5083 1733 5087
rect 1447 5073 1463 5083
rect 1457 5047 1463 5073
rect 1717 5073 1733 5083
rect 2140 5083 2153 5087
rect 2137 5073 2153 5083
rect 2253 5083 2267 5093
rect 2253 5080 2283 5083
rect 2257 5077 2283 5080
rect 1457 5037 1473 5047
rect 1460 5033 1473 5037
rect 1717 5043 1723 5073
rect 1687 5037 1723 5043
rect 2137 5047 2143 5073
rect 2277 5047 2283 5077
rect 2137 5037 2153 5047
rect 2140 5033 2153 5037
rect 2267 5037 2283 5047
rect 2267 5033 2280 5037
rect 2297 5027 2303 5117
rect 3007 5117 3053 5123
rect 2387 5093 2393 5107
rect 2987 5097 3073 5103
rect 3287 5097 3353 5103
rect 3447 5097 3493 5103
rect 4447 5097 4493 5103
rect 5521 5097 5633 5103
rect 6207 5103 6220 5107
rect 6207 5093 6223 5103
rect 2727 5077 2773 5083
rect 3340 5086 3360 5087
rect 3340 5083 3353 5086
rect 3337 5073 3353 5083
rect 3337 5047 3343 5073
rect 4147 5083 4160 5087
rect 4147 5073 4163 5083
rect 4157 5047 4163 5073
rect 3337 5037 3353 5047
rect 3340 5033 3353 5037
rect 4147 5037 4163 5047
rect 4717 5047 4723 5093
rect 4827 5083 4840 5087
rect 5940 5083 5953 5087
rect 4827 5073 4843 5083
rect 4837 5047 4843 5073
rect 5937 5073 5953 5083
rect 6077 5077 6113 5083
rect 5937 5047 5943 5073
rect 6077 5047 6083 5077
rect 6217 5083 6223 5093
rect 6217 5077 6243 5083
rect 6237 5047 6243 5077
rect 4717 5037 4733 5047
rect 4147 5033 4160 5037
rect 4720 5033 4733 5037
rect 4827 5037 4843 5047
rect 4827 5033 4840 5037
rect 5927 5037 5943 5047
rect 5927 5033 5940 5037
rect 6067 5037 6083 5047
rect 6067 5033 6080 5037
rect 6227 5037 6243 5047
rect 6227 5033 6240 5037
rect 1587 5017 1633 5023
rect 2280 5026 2303 5027
rect 2287 5017 2303 5026
rect 2287 5013 2300 5017
rect 5947 5017 6013 5023
rect 6443 4958 6503 5462
rect 6410 4942 6503 4958
rect 1647 4897 1673 4903
rect 4207 4897 4253 4903
rect 47 4877 93 4883
rect 4987 4877 5093 4883
rect 167 4863 180 4867
rect 167 4853 183 4863
rect 177 4827 183 4853
rect 337 4827 343 4873
rect 360 4863 373 4867
rect 167 4817 183 4827
rect 167 4813 180 4817
rect 327 4817 343 4827
rect 357 4853 373 4863
rect 1167 4857 1193 4863
rect 2020 4863 2033 4867
rect 2017 4853 2033 4863
rect 2580 4863 2593 4867
rect 2577 4853 2593 4863
rect 3920 4863 3933 4867
rect 3917 4853 3933 4863
rect 4047 4863 4060 4867
rect 4047 4853 4063 4863
rect 5847 4863 5860 4867
rect 5847 4853 5863 4863
rect 5987 4863 6000 4867
rect 5987 4853 6003 4863
rect 6127 4863 6140 4867
rect 6160 4863 6173 4867
rect 6127 4853 6143 4863
rect 357 4827 363 4853
rect 357 4817 373 4827
rect 327 4813 340 4817
rect 360 4813 373 4817
rect 2017 4823 2023 4853
rect 1987 4817 2023 4823
rect 2577 4827 2583 4853
rect 3917 4827 3923 4853
rect 4057 4827 4063 4853
rect 5857 4827 5863 4853
rect 2577 4817 2593 4827
rect 2580 4813 2593 4817
rect 3917 4817 3933 4827
rect 3920 4813 3933 4817
rect 4047 4817 4063 4827
rect 4047 4813 4060 4817
rect 4367 4817 4393 4823
rect 5857 4817 5873 4827
rect 5860 4813 5873 4817
rect 5997 4823 6003 4853
rect 5997 4817 6023 4823
rect 6017 4807 6023 4817
rect 6137 4807 6143 4853
rect 6157 4853 6173 4863
rect 6247 4863 6260 4867
rect 6247 4853 6263 4863
rect 6157 4827 6163 4853
rect 6257 4827 6263 4853
rect 6157 4817 6173 4827
rect 6160 4813 6173 4817
rect 6247 4817 6263 4827
rect 6247 4813 6260 4817
rect 1747 4797 1793 4803
rect 1847 4797 1913 4803
rect 2547 4797 2653 4803
rect 3867 4797 3973 4803
rect 4927 4797 4953 4803
rect 4967 4797 5073 4803
rect 5567 4797 5613 4803
rect 5867 4797 5933 4803
rect 6017 4797 6033 4807
rect 6020 4793 6033 4797
rect 2727 4777 2753 4783
rect 4047 4757 4093 4763
rect 5987 4737 6013 4743
rect 1167 4717 1213 4723
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 5827 4657 5853 4663
rect 2047 4617 2113 4623
rect 2667 4617 2713 4623
rect 1607 4597 1653 4603
rect 207 4577 293 4583
rect 537 4577 593 4583
rect 377 4527 383 4573
rect 537 4563 543 4577
rect 1287 4577 1413 4583
rect 1467 4577 1493 4583
rect 1607 4577 1653 4583
rect 2120 4583 2133 4587
rect 517 4557 543 4563
rect 377 4517 393 4527
rect 380 4513 393 4517
rect 517 4507 523 4557
rect 1487 4563 1500 4567
rect 1487 4553 1503 4563
rect 1627 4563 1640 4567
rect 1753 4563 1767 4573
rect 2117 4573 2133 4583
rect 2307 4577 2453 4583
rect 3437 4577 3493 4583
rect 2117 4563 2123 4573
rect 1627 4553 1643 4563
rect 1753 4560 1783 4563
rect 1757 4557 1783 4560
rect 1497 4523 1503 4553
rect 1637 4527 1643 4553
rect 1777 4527 1783 4557
rect 1497 4517 1533 4523
rect 1627 4517 1643 4527
rect 1627 4513 1640 4517
rect 1767 4517 1783 4527
rect 2097 4557 2123 4563
rect 2097 4527 2103 4557
rect 2367 4563 2380 4567
rect 2367 4553 2383 4563
rect 2907 4563 2920 4567
rect 3080 4563 3093 4567
rect 2907 4553 2923 4563
rect 2377 4527 2383 4553
rect 2097 4517 2113 4527
rect 1767 4513 1780 4517
rect 2100 4513 2113 4517
rect 2367 4517 2383 4527
rect 2917 4527 2923 4553
rect 3077 4553 3093 4563
rect 3077 4527 3083 4553
rect 3437 4527 3443 4577
rect 4127 4577 4193 4583
rect 4420 4583 4433 4587
rect 4417 4573 4433 4583
rect 5087 4577 5113 4583
rect 5287 4577 5333 4583
rect 5447 4577 5473 4583
rect 3460 4563 3473 4567
rect 2917 4517 2933 4527
rect 2367 4513 2380 4517
rect 2920 4513 2933 4517
rect 3077 4517 3093 4527
rect 3080 4513 3093 4517
rect 3427 4517 3443 4527
rect 3457 4553 3473 4563
rect 3457 4527 3463 4553
rect 3977 4527 3983 4573
rect 3457 4517 3473 4527
rect 3427 4513 3440 4517
rect 3460 4513 3473 4517
rect 3977 4517 3993 4527
rect 3980 4513 3993 4517
rect 4417 4523 4423 4573
rect 5000 4563 5013 4567
rect 4997 4553 5013 4563
rect 5407 4557 5443 4563
rect 4997 4527 5003 4553
rect 4387 4517 4423 4523
rect 4987 4517 5003 4527
rect 5437 4527 5443 4557
rect 5687 4563 5700 4567
rect 5860 4563 5873 4567
rect 5687 4553 5703 4563
rect 5697 4527 5703 4553
rect 5437 4517 5453 4527
rect 4987 4513 5000 4517
rect 5440 4513 5453 4517
rect 5687 4517 5703 4527
rect 5857 4553 5873 4563
rect 5947 4563 5960 4567
rect 5947 4553 5963 4563
rect 6267 4563 6280 4567
rect 6267 4553 6283 4563
rect 5687 4513 5700 4517
rect 5857 4507 5863 4553
rect 1467 4497 1493 4503
rect 2307 4497 2393 4503
rect 3687 4497 3733 4503
rect 3787 4497 3853 4503
rect 3927 4497 4033 4503
rect 5547 4497 5613 4503
rect 5847 4497 5863 4507
rect 5957 4507 5963 4553
rect 6277 4527 6283 4553
rect 6267 4517 6283 4527
rect 6267 4513 6280 4517
rect 5957 4506 5980 4507
rect 5957 4497 5973 4506
rect 5847 4493 5860 4497
rect 5960 4493 5973 4497
rect 2517 4480 2573 4483
rect 2513 4477 2573 4480
rect 2513 4467 2527 4477
rect 6443 4438 6503 4942
rect 6410 4422 6503 4438
rect 2587 4397 2633 4403
rect 3907 4357 3953 4363
rect 4667 4357 4713 4363
rect 4727 4357 4773 4363
rect 4847 4357 4893 4363
rect 5687 4357 5773 4363
rect 6367 4357 6413 4363
rect 1767 4343 1780 4347
rect 1767 4333 1783 4343
rect 1907 4343 1920 4347
rect 1907 4333 1923 4343
rect 2207 4343 2220 4347
rect 2240 4343 2253 4347
rect 2207 4333 2223 4343
rect 1777 4307 1783 4333
rect 1467 4297 1493 4303
rect 1767 4297 1783 4307
rect 1767 4293 1780 4297
rect 1087 4277 1173 4283
rect 1227 4277 1353 4283
rect 1407 4277 1513 4283
rect 1707 4277 1793 4283
rect 1917 4283 1923 4333
rect 2217 4307 2223 4333
rect 2207 4297 2223 4307
rect 2237 4333 2253 4343
rect 2237 4307 2243 4333
rect 2377 4307 2383 4353
rect 2780 4343 2793 4347
rect 2777 4333 2793 4343
rect 4527 4337 4563 4343
rect 2777 4307 2783 4333
rect 4557 4307 4563 4337
rect 5167 4343 5180 4347
rect 5167 4333 5183 4343
rect 5177 4307 5183 4333
rect 2237 4297 2253 4307
rect 2207 4293 2220 4297
rect 2240 4293 2253 4297
rect 2377 4297 2393 4307
rect 2380 4293 2393 4297
rect 2777 4297 2793 4307
rect 2780 4293 2793 4297
rect 4557 4297 4573 4307
rect 4560 4293 4573 4297
rect 5167 4297 5183 4307
rect 5167 4293 5180 4297
rect 5547 4297 5573 4303
rect 1867 4277 1923 4283
rect 3767 4277 3813 4283
rect 4827 4277 4853 4283
rect 5147 4277 5233 4283
rect 2607 4257 2633 4263
rect 3027 4257 3113 4263
rect 5187 4257 5233 4263
rect 2747 4217 2793 4223
rect 3907 4197 3933 4203
rect -63 4162 30 4178
rect -63 3658 -3 4162
rect 3247 4117 3273 4123
rect 1547 4097 1633 4103
rect 1581 4077 1613 4083
rect 187 4057 253 4063
rect 467 4057 593 4063
rect 1077 4057 1113 4063
rect 927 4043 940 4047
rect 1077 4043 1083 4057
rect 1547 4057 1573 4063
rect 3147 4057 3193 4063
rect 3627 4063 3640 4067
rect 3627 4054 3643 4063
rect 3620 4053 3643 4054
rect 4767 4057 4793 4063
rect 5007 4057 5053 4063
rect 5207 4057 5233 4063
rect 1200 4043 1213 4047
rect 927 4033 943 4043
rect 937 4007 943 4033
rect 1057 4037 1083 4043
rect 937 3997 953 4007
rect 940 3993 953 3997
rect 1057 4003 1063 4037
rect 1197 4033 1213 4043
rect 1340 4043 1353 4047
rect 1337 4033 1353 4043
rect 1447 4043 1460 4047
rect 2600 4043 2613 4047
rect 1447 4033 1463 4043
rect 1197 4007 1203 4033
rect 1027 3997 1063 4003
rect 1187 3997 1203 4007
rect 1337 4007 1343 4033
rect 1337 3997 1353 4007
rect 1187 3993 1200 3997
rect 1340 3993 1353 3997
rect 1457 4006 1463 4033
rect 2597 4033 2613 4043
rect 2727 4043 2740 4047
rect 2727 4033 2743 4043
rect 2887 4043 2900 4047
rect 2887 4033 2903 4043
rect 2987 4043 3000 4047
rect 2987 4033 3003 4043
rect 3527 4043 3540 4047
rect 3637 4043 3643 4053
rect 4060 4043 4073 4047
rect 3527 4033 3543 4043
rect 3637 4037 3663 4043
rect 2597 4007 2603 4033
rect 2737 4007 2743 4033
rect 2597 3997 2613 4007
rect 2600 3993 2613 3997
rect 2727 3997 2743 4007
rect 2897 4007 2903 4033
rect 2997 4027 3003 4033
rect 2997 4026 3020 4027
rect 2997 4017 3013 4026
rect 3000 4013 3013 4017
rect 3537 4007 3543 4033
rect 3657 4007 3663 4037
rect 2897 3997 2913 4007
rect 2727 3993 2740 3997
rect 2900 3993 2913 3997
rect 3537 3997 3553 4007
rect 3540 3993 3553 3997
rect 3647 3997 3663 4007
rect 4057 4033 4073 4043
rect 4220 4043 4233 4047
rect 4217 4033 4233 4043
rect 6040 4043 6053 4047
rect 6037 4033 6053 4043
rect 4057 4007 4063 4033
rect 4217 4007 4223 4033
rect 6037 4007 6043 4033
rect 4057 3997 4073 4007
rect 3647 3993 3660 3997
rect 4060 3993 4073 3997
rect 4217 3997 4233 4007
rect 4220 3993 4233 3997
rect 6037 3997 6053 4007
rect 6040 3993 6053 3997
rect 2327 3977 2353 3983
rect 2907 3977 2933 3983
rect 5907 3977 5959 3983
rect 6443 3918 6503 4422
rect 6410 3902 6503 3918
rect 27 3877 73 3883
rect 4947 3857 4973 3863
rect 5267 3857 5313 3863
rect 407 3837 453 3843
rect 5687 3837 5733 3843
rect 167 3823 180 3827
rect 167 3813 183 3823
rect 177 3787 183 3813
rect 1040 3823 1053 3827
rect 733 3803 747 3813
rect 1037 3813 1053 3823
rect 1740 3823 1753 3827
rect 1737 3813 1753 3823
rect 733 3800 763 3803
rect 737 3797 763 3800
rect 167 3777 183 3787
rect 167 3773 180 3777
rect 757 3766 763 3797
rect 1037 3787 1043 3813
rect 1737 3787 1743 3813
rect 1037 3777 1053 3787
rect 1040 3773 1053 3777
rect 1737 3777 1767 3787
rect 1740 3773 1767 3777
rect 2017 3766 2023 3833
rect 2267 3823 2280 3827
rect 2300 3823 2313 3827
rect 2267 3820 2283 3823
rect 2267 3813 2287 3820
rect 2273 3806 2287 3813
rect 2297 3813 2313 3823
rect 2797 3817 2833 3823
rect 2297 3783 2303 3813
rect 2797 3787 2803 3817
rect 4040 3826 4060 3827
rect 4047 3823 4060 3826
rect 4047 3813 4063 3823
rect 4627 3823 4640 3827
rect 4627 3813 4643 3823
rect 5847 3823 5860 3827
rect 5847 3813 5863 3823
rect 6127 3817 6163 3823
rect 2267 3777 2303 3783
rect 2647 3777 2673 3783
rect 2787 3777 2803 3787
rect 4057 3787 4063 3813
rect 4637 3787 4643 3813
rect 4057 3777 4073 3787
rect 2787 3773 2800 3777
rect 4060 3773 4073 3777
rect 4627 3777 4643 3787
rect 4627 3773 4640 3777
rect 5857 3767 5863 3813
rect 6157 3787 6163 3817
rect 6287 3823 6300 3827
rect 6287 3813 6303 3823
rect 6157 3777 6173 3787
rect 6160 3773 6173 3777
rect 6297 3783 6303 3813
rect 6277 3777 6303 3783
rect 2107 3757 2173 3763
rect 3087 3757 3133 3763
rect 3867 3757 3913 3763
rect 3927 3757 3973 3763
rect 4347 3757 4413 3763
rect 5547 3757 5633 3763
rect 5857 3757 5873 3767
rect 5860 3753 5873 3757
rect 5967 3757 6073 3763
rect 6277 3763 6283 3777
rect 6227 3757 6283 3763
rect 3747 3720 3803 3723
rect 3747 3717 3807 3720
rect 3793 3707 3807 3717
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 1607 3597 1633 3603
rect 547 3577 573 3583
rect 1707 3577 1773 3583
rect 1267 3557 1333 3563
rect 5447 3557 5473 3563
rect 5487 3557 5513 3563
rect 687 3537 813 3543
rect 1427 3537 1493 3543
rect 1847 3543 1860 3547
rect 1847 3534 1863 3543
rect 1840 3533 1863 3534
rect 1887 3537 1913 3543
rect 1967 3537 2003 3543
rect 717 3517 753 3523
rect 257 3487 263 3513
rect 717 3487 723 3517
rect 1037 3517 1073 3523
rect 1037 3487 1043 3517
rect 1160 3523 1173 3527
rect 1157 3513 1173 3523
rect 1760 3523 1773 3527
rect 1757 3513 1773 3523
rect 1857 3523 1863 3533
rect 1997 3523 2003 3537
rect 2987 3537 3013 3543
rect 1857 3517 1883 3523
rect 1997 3517 2023 3523
rect 707 3477 723 3487
rect 707 3473 720 3477
rect 1027 3477 1043 3487
rect 1157 3487 1163 3513
rect 1157 3477 1173 3487
rect 1027 3473 1040 3477
rect 1160 3473 1173 3477
rect 1607 3477 1633 3483
rect 1757 3483 1763 3513
rect 1877 3483 1883 3517
rect 2017 3483 2023 3517
rect 2147 3523 2160 3527
rect 2460 3523 2473 3527
rect 2147 3513 2163 3523
rect 1757 3477 1783 3483
rect 1877 3480 1903 3483
rect 1877 3477 1907 3480
rect 2017 3477 2053 3483
rect 1777 3467 1783 3477
rect 1893 3467 1907 3477
rect 727 3457 753 3463
rect 1707 3457 1733 3463
rect 1777 3457 1793 3467
rect 1780 3453 1793 3457
rect 2157 3463 2163 3513
rect 2457 3513 2473 3523
rect 6007 3523 6020 3527
rect 6007 3513 6023 3523
rect 2457 3483 2463 3513
rect 2427 3477 2463 3483
rect 6017 3483 6023 3513
rect 6017 3477 6053 3483
rect 2127 3457 2163 3463
rect 1047 3437 1073 3443
rect 6443 3398 6503 3902
rect 6410 3382 6503 3398
rect 2037 3337 2073 3343
rect 467 3317 533 3323
rect 1227 3317 1313 3323
rect 1407 3317 1433 3323
rect 300 3303 313 3307
rect 297 3293 313 3303
rect 427 3297 463 3303
rect 297 3267 303 3293
rect 297 3257 313 3267
rect 300 3253 313 3257
rect 457 3263 463 3297
rect 897 3267 903 3313
rect 997 3267 1003 3313
rect 1020 3303 1033 3307
rect 457 3257 483 3263
rect 897 3257 913 3267
rect 367 3237 433 3243
rect 477 3243 483 3257
rect 900 3253 913 3257
rect 987 3257 1003 3267
rect 1017 3293 1033 3303
rect 1160 3303 1173 3307
rect 1157 3293 1173 3303
rect 1647 3303 1660 3307
rect 2037 3303 2043 3337
rect 5167 3337 5213 3343
rect 2167 3317 2233 3323
rect 1647 3293 1663 3303
rect 2037 3297 2073 3303
rect 2207 3303 2220 3307
rect 2207 3293 2223 3303
rect 4007 3293 4013 3307
rect 4860 3303 4873 3307
rect 4857 3293 4873 3303
rect 4987 3303 5000 3307
rect 4987 3293 5003 3303
rect 1017 3267 1023 3293
rect 1157 3267 1163 3293
rect 1017 3257 1033 3267
rect 987 3253 1000 3257
rect 1020 3253 1033 3257
rect 1157 3257 1173 3267
rect 1160 3253 1173 3257
rect 1657 3263 1663 3293
rect 2217 3267 2223 3293
rect 4857 3267 4863 3293
rect 1657 3257 1693 3263
rect 2217 3257 2233 3267
rect 2220 3253 2233 3257
rect 4857 3257 4873 3267
rect 4860 3253 4873 3257
rect 4997 3263 5003 3293
rect 5867 3297 5913 3303
rect 4997 3257 5033 3263
rect 477 3237 533 3243
rect 687 3237 813 3243
rect 2287 3237 2393 3243
rect 3867 3237 3953 3243
rect 4027 3237 4073 3243
rect -63 3122 30 3138
rect -63 2618 -3 3122
rect 1720 3066 1733 3067
rect 1727 3053 1733 3066
rect 2327 3037 2413 3043
rect 287 3017 313 3023
rect 427 3017 473 3023
rect 917 3017 973 3023
rect 37 2994 67 3008
rect 37 2946 43 2994
rect 917 2967 923 3017
rect 5827 3017 5933 3023
rect 1047 3003 1060 3007
rect 1047 2993 1063 3003
rect 1667 3003 1680 3007
rect 1960 3003 1973 3007
rect 1667 2993 1683 3003
rect 917 2957 933 2967
rect 920 2953 933 2957
rect 1057 2963 1063 2993
rect 1057 2957 1093 2963
rect 1677 2963 1683 2993
rect 1957 2993 1973 3003
rect 2347 3003 2360 3007
rect 2640 3003 2653 3007
rect 2347 2993 2363 3003
rect 1957 2967 1963 2993
rect 1677 2957 1713 2963
rect 1957 2957 1973 2967
rect 1960 2953 1973 2957
rect 2357 2963 2363 2993
rect 2637 2993 2653 3003
rect 4060 3003 4073 3007
rect 4057 2993 4073 3003
rect 5140 3003 5153 3007
rect 5137 2993 5153 3003
rect 2637 2983 2643 2993
rect 2617 2977 2643 2983
rect 2617 2967 2623 2977
rect 2357 2957 2393 2963
rect 2607 2957 2623 2967
rect 4057 2967 4063 2993
rect 4057 2957 4073 2967
rect 2607 2953 2620 2957
rect 4060 2953 4073 2957
rect 287 2937 373 2943
rect 1787 2937 1813 2943
rect 2113 2943 2127 2953
rect 2047 2940 2127 2943
rect 2047 2937 2123 2940
rect 2387 2937 2413 2943
rect 5137 2943 5143 2993
rect 5107 2937 5143 2943
rect 6443 2878 6503 3382
rect 6410 2862 6503 2878
rect 1247 2797 1273 2803
rect 1107 2783 1120 2787
rect 1107 2773 1123 2783
rect 1117 2743 1123 2773
rect 1397 2777 1433 2783
rect 1397 2747 1403 2777
rect 1557 2777 1593 2783
rect 1557 2747 1563 2777
rect 3407 2777 3453 2783
rect 5227 2777 5273 2783
rect 1097 2737 1123 2743
rect 207 2717 273 2723
rect 447 2717 513 2723
rect 527 2717 573 2723
rect 1097 2723 1103 2737
rect 1387 2737 1403 2747
rect 1387 2733 1400 2737
rect 1547 2737 1563 2747
rect 1547 2733 1560 2737
rect 1067 2717 1103 2723
rect 1367 2717 1393 2723
rect 1487 2717 1513 2723
rect 2727 2717 2753 2723
rect 2807 2717 2913 2723
rect 3153 2723 3167 2733
rect 3107 2720 3167 2723
rect 3107 2717 3163 2720
rect 4047 2717 4073 2723
rect 1487 2697 1553 2703
rect -63 2602 30 2618
rect -63 2098 -3 2602
rect 507 2517 593 2523
rect 1227 2517 1253 2523
rect 427 2497 553 2503
rect 1187 2497 1253 2503
rect 2527 2497 2593 2503
rect 937 2477 973 2483
rect 937 2426 943 2477
rect 1220 2483 1233 2487
rect 1217 2473 1233 2483
rect 1217 2447 1223 2473
rect 1207 2437 1223 2447
rect 1207 2433 1220 2437
rect 1357 2407 1363 2493
rect 1740 2483 1753 2487
rect 1737 2473 1753 2483
rect 2267 2483 2280 2487
rect 2267 2473 2283 2483
rect 2647 2483 2660 2487
rect 2647 2473 2663 2483
rect 3527 2477 3553 2483
rect 1737 2447 1743 2473
rect 2277 2447 2283 2473
rect 2657 2447 2663 2473
rect 1727 2437 1743 2447
rect 1727 2433 1740 2437
rect 2107 2437 2153 2443
rect 2267 2437 2283 2447
rect 2267 2433 2280 2437
rect 2647 2437 2663 2447
rect 2647 2433 2660 2437
rect 6287 2417 6333 2423
rect 1347 2397 1363 2407
rect 1347 2393 1360 2397
rect 6443 2358 6503 2862
rect 6410 2342 6503 2358
rect 2047 2323 2060 2327
rect 2047 2313 2063 2323
rect 847 2297 873 2303
rect 2021 2297 2033 2303
rect 1167 2277 1253 2283
rect 197 2227 203 2273
rect 2057 2283 2063 2313
rect 2007 2277 2063 2283
rect 2527 2277 2573 2283
rect 767 2263 780 2267
rect 767 2253 783 2263
rect 1307 2257 1343 2263
rect 777 2227 783 2253
rect 197 2217 213 2227
rect 200 2213 213 2217
rect 767 2217 783 2227
rect 1337 2227 1343 2257
rect 1467 2263 1480 2267
rect 1500 2263 1513 2267
rect 1467 2253 1483 2263
rect 1477 2227 1483 2253
rect 1337 2217 1353 2227
rect 767 2213 780 2217
rect 1340 2213 1353 2217
rect 1467 2217 1483 2227
rect 1497 2253 1513 2263
rect 1727 2263 1740 2267
rect 1727 2253 1743 2263
rect 2287 2263 2300 2267
rect 2580 2263 2593 2267
rect 2287 2253 2303 2263
rect 1467 2213 1480 2217
rect 1497 2207 1503 2253
rect 1737 2227 1743 2253
rect 2297 2227 2303 2253
rect 2577 2253 2593 2263
rect 2667 2263 2680 2267
rect 2667 2253 2683 2263
rect 2807 2263 2820 2267
rect 2807 2253 2823 2263
rect 3447 2263 3460 2267
rect 3447 2253 3463 2263
rect 4187 2257 4223 2263
rect 2577 2227 2583 2253
rect 2677 2227 2683 2253
rect 2817 2227 2823 2253
rect 3457 2227 3463 2253
rect 1737 2217 1753 2227
rect 1740 2213 1753 2217
rect 2297 2217 2313 2227
rect 2300 2213 2313 2217
rect 2577 2217 2593 2227
rect 2580 2213 2593 2217
rect 2677 2217 2693 2227
rect 2680 2213 2693 2217
rect 2807 2217 2823 2227
rect 2807 2213 2820 2217
rect 3447 2217 3463 2227
rect 4217 2227 4223 2257
rect 4217 2217 4233 2227
rect 3447 2213 3460 2217
rect 4220 2213 4233 2217
rect 307 2197 433 2203
rect 1347 2197 1393 2203
rect 1480 2206 1503 2207
rect 1487 2197 1503 2206
rect 1487 2193 1500 2197
rect 1567 2197 1653 2203
rect 1827 2197 1893 2203
rect 1653 2143 1667 2153
rect 1627 2140 1667 2143
rect 1627 2137 1663 2140
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 507 2017 533 2023
rect 1447 2017 1513 2023
rect 2067 2017 2093 2023
rect 327 1977 393 1983
rect 507 1977 573 1983
rect 787 1977 853 1983
rect 1380 1983 1393 1987
rect 1287 1977 1393 1983
rect 1377 1973 1393 1977
rect 3087 1977 3253 1983
rect 3587 1977 3673 1983
rect 5247 1977 5273 1983
rect 1377 1963 1383 1973
rect 1357 1957 1383 1963
rect 1357 1927 1363 1957
rect 1587 1963 1600 1967
rect 2360 1963 2373 1967
rect 1587 1953 1603 1963
rect 1597 1927 1603 1953
rect 2357 1953 2373 1963
rect 2720 1963 2733 1967
rect 2717 1953 2733 1963
rect 2357 1927 2363 1953
rect 2717 1927 2723 1953
rect 3613 1927 3627 1933
rect 167 1917 193 1923
rect 1347 1917 1363 1927
rect 1347 1913 1360 1917
rect 1587 1917 1603 1927
rect 1587 1913 1600 1917
rect 2207 1917 2233 1923
rect 2357 1917 2373 1927
rect 2360 1913 2373 1917
rect 2717 1917 2733 1927
rect 2720 1913 2733 1917
rect 3613 1920 3633 1927
rect 3617 1917 3633 1920
rect 3620 1913 3633 1917
rect 367 1897 393 1903
rect 907 1897 933 1903
rect 1747 1897 1773 1903
rect 6443 1838 6503 2342
rect 6410 1822 6503 1838
rect 6127 1797 6153 1803
rect 787 1757 853 1763
rect 1007 1757 1053 1763
rect 1687 1757 1733 1763
rect 2667 1757 2713 1763
rect 2357 1707 2363 1753
rect 2817 1707 2823 1733
rect 2357 1697 2373 1707
rect 2360 1693 2373 1697
rect 2817 1697 2833 1707
rect 2820 1693 2833 1697
rect 687 1677 813 1683
rect 1847 1677 1953 1683
rect 3627 1677 3653 1683
rect 5167 1677 5233 1683
rect 3533 1663 3547 1671
rect 3507 1660 3547 1663
rect 3507 1657 3543 1660
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 127 1457 273 1463
rect 567 1457 693 1463
rect 747 1457 873 1463
rect 927 1457 953 1463
rect 1827 1457 1913 1463
rect 1927 1457 1993 1463
rect 2427 1457 2493 1463
rect 5287 1457 5333 1463
rect 340 1443 353 1447
rect 337 1433 353 1443
rect 1467 1443 1480 1447
rect 1467 1433 1483 1443
rect 337 1407 343 1433
rect 327 1397 343 1407
rect 1477 1407 1483 1433
rect 2057 1437 2093 1443
rect 2057 1407 2063 1437
rect 1477 1397 1493 1407
rect 327 1393 340 1397
rect 1480 1393 1493 1397
rect 2047 1397 2063 1407
rect 2047 1393 2060 1397
rect 2867 1400 2923 1403
rect 2867 1397 2927 1400
rect 2913 1387 2927 1397
rect 6443 1318 6503 1822
rect 6410 1302 6503 1318
rect 1987 1257 2033 1263
rect 3447 1237 3533 1243
rect 1297 1217 1333 1223
rect 1297 1187 1303 1217
rect 1987 1223 2000 1227
rect 2020 1223 2033 1227
rect 1987 1213 2003 1223
rect 1287 1177 1303 1187
rect 1997 1183 2003 1213
rect 1977 1177 2003 1183
rect 2017 1213 2033 1223
rect 2160 1223 2173 1227
rect 2157 1213 2173 1223
rect 2260 1223 2273 1227
rect 2257 1213 2273 1223
rect 2017 1187 2023 1213
rect 2017 1177 2033 1187
rect 1287 1173 1300 1177
rect 407 1157 473 1163
rect 497 1147 503 1173
rect 1227 1157 1313 1163
rect 1977 1163 1983 1177
rect 2020 1173 2033 1177
rect 2157 1183 2163 1213
rect 2137 1177 2163 1183
rect 2257 1183 2263 1213
rect 2557 1183 2563 1233
rect 2940 1223 2953 1227
rect 2937 1213 2953 1223
rect 2937 1187 2943 1213
rect 2257 1177 2283 1183
rect 1947 1157 1983 1163
rect 2137 1163 2143 1177
rect 2107 1157 2143 1163
rect 2277 1167 2283 1177
rect 2537 1177 2563 1183
rect 2277 1157 2293 1167
rect 2280 1153 2293 1157
rect 2537 1163 2543 1177
rect 2927 1177 2943 1187
rect 3637 1183 3643 1233
rect 6240 1223 6253 1227
rect 6237 1213 6253 1223
rect 6237 1187 6243 1213
rect 3617 1177 3643 1183
rect 2927 1173 2940 1177
rect 2487 1157 2573 1163
rect 3617 1163 3623 1177
rect 6227 1177 6243 1187
rect 6227 1173 6240 1177
rect 3587 1157 3623 1163
rect 6067 1157 6153 1163
rect 6247 1157 6293 1163
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 567 937 713 943
rect 987 937 1113 943
rect 3007 937 3033 943
rect 3187 937 3233 943
rect 167 923 180 927
rect 167 913 183 923
rect 2907 923 2920 927
rect 2907 913 2923 923
rect 4667 917 4693 923
rect 177 887 183 913
rect 2917 887 2923 913
rect 167 877 183 887
rect 167 873 180 877
rect 2907 877 2923 887
rect 2907 873 2920 877
rect 2647 857 2733 863
rect 5927 857 5973 863
rect 1067 817 1093 823
rect 6443 798 6503 1302
rect 6410 782 6503 798
rect 287 717 313 723
rect 2227 717 2293 723
rect 3247 717 3273 723
rect 1373 703 1387 713
rect 1373 700 1433 703
rect 1377 697 1433 700
rect 1397 667 1403 697
rect 1667 697 1693 703
rect 3400 703 3413 707
rect 3397 693 3413 703
rect 1387 657 1403 667
rect 3397 667 3403 693
rect 3397 657 3413 667
rect 1387 653 1400 657
rect 3400 653 3413 657
rect 1427 637 1473 643
rect 1907 637 1973 643
rect -63 522 30 538
rect -63 18 -3 522
rect 627 417 653 423
rect 1047 417 1113 423
rect 1527 417 1613 423
rect 5107 417 5193 423
rect 6107 417 6133 423
rect 6187 417 6233 423
rect 667 357 693 363
rect 827 357 853 363
rect 1227 337 1313 343
rect 2247 337 2273 343
rect 6443 278 6503 782
rect 6410 262 6503 278
rect 2847 197 2873 203
rect 287 183 300 187
rect 287 173 303 183
rect 1313 183 1327 193
rect 1980 183 1993 187
rect 1287 180 1327 183
rect 1287 177 1323 180
rect 1977 173 1993 183
rect 297 147 303 173
rect 1977 147 1983 173
rect 297 137 313 147
rect 300 133 313 137
rect 1967 137 1983 147
rect 1967 133 1980 137
rect 887 117 953 123
rect 2327 117 2393 123
rect 6327 117 6393 123
rect -63 2 30 18
rect 6443 2 6503 262
<< m2contact >>
rect 3233 6173 3247 6187
rect 3253 6173 3267 6187
rect 2353 6153 2367 6167
rect 2433 6153 2447 6167
rect 3333 6153 3347 6167
rect 3373 6153 3387 6167
rect 1973 6133 1987 6147
rect 2013 6133 2027 6147
rect 2793 6133 2807 6147
rect 2873 6133 2887 6147
rect 3173 6133 3187 6147
rect 3293 6134 3307 6148
rect 4553 6134 4567 6148
rect 4633 6133 4647 6147
rect 4933 6133 4947 6147
rect 4973 6133 4987 6147
rect 6333 6133 6347 6147
rect 6373 6133 6387 6147
rect 493 6113 507 6127
rect 3413 6113 3427 6127
rect 3813 6113 3827 6127
rect 6093 6113 6107 6127
rect 3413 6073 3427 6087
rect 3813 6073 3827 6087
rect 6153 6073 6167 6087
rect 513 6052 527 6066
rect 1593 6053 1607 6067
rect 1753 6053 1767 6067
rect 1813 6053 1827 6067
rect 2513 6053 2527 6067
rect 2613 6053 2627 6067
rect 3173 6053 3187 6067
rect 3293 6053 3307 6067
rect 4173 6053 4187 6067
rect 4253 6053 4267 6067
rect 1713 6033 1727 6047
rect 2593 6033 2607 6047
rect 2673 6033 2687 6047
rect 2393 6012 2407 6026
rect 2433 6013 2447 6027
rect 613 5953 627 5967
rect 673 5952 687 5966
rect 333 5913 347 5927
rect 567 5914 581 5928
rect 593 5913 607 5927
rect 2233 5913 2247 5927
rect 2313 5914 2327 5928
rect 3693 5913 3707 5927
rect 3753 5913 3767 5927
rect 513 5893 527 5907
rect 3853 5893 3867 5907
rect 4073 5893 4087 5907
rect 4373 5933 4387 5947
rect 4353 5913 4367 5927
rect 4413 5913 4427 5927
rect 5173 5913 5187 5927
rect 5333 5912 5347 5926
rect 4673 5893 4687 5907
rect 313 5853 327 5867
rect 473 5853 487 5867
rect 3553 5853 3567 5867
rect 3593 5853 3607 5867
rect 3853 5853 3867 5867
rect 4033 5853 4047 5867
rect 4333 5853 4347 5867
rect 4633 5853 4647 5867
rect 933 5833 947 5847
rect 999 5833 1013 5847
rect 1053 5833 1067 5847
rect 1113 5833 1127 5847
rect 2173 5831 2187 5845
rect 2213 5833 2227 5847
rect 2293 5831 2307 5845
rect 2493 5833 2507 5847
rect 2553 5833 2567 5847
rect 2633 5833 2647 5847
rect 2753 5833 2767 5847
rect 3413 5833 3427 5847
rect 3453 5833 3467 5847
rect 3833 5833 3847 5847
rect 3953 5833 3967 5847
rect 833 5813 847 5827
rect 873 5812 887 5826
rect 2213 5812 2227 5826
rect 3353 5813 3367 5827
rect 3473 5813 3487 5827
rect 1713 5653 1727 5667
rect 1773 5653 1787 5667
rect 953 5633 967 5647
rect 1053 5633 1067 5647
rect 1733 5633 1747 5647
rect 1773 5632 1787 5646
rect 3213 5633 3227 5647
rect 3253 5633 3267 5647
rect 4633 5633 4647 5647
rect 4693 5633 4707 5647
rect 513 5614 527 5628
rect 553 5613 567 5627
rect 593 5613 607 5627
rect 1173 5613 1187 5627
rect 1233 5613 1247 5627
rect 1413 5613 1427 5627
rect 1493 5613 1507 5627
rect 3173 5613 3187 5627
rect 3253 5612 3267 5626
rect 173 5593 187 5607
rect 3573 5613 3587 5627
rect 4113 5613 4127 5627
rect 4173 5613 4187 5627
rect 6033 5613 6047 5627
rect 6173 5613 6187 5627
rect 6293 5593 6307 5607
rect 6373 5593 6387 5607
rect 3473 5553 3487 5567
rect 6253 5553 6267 5567
rect 173 5533 187 5547
rect 1713 5533 1727 5547
rect 1773 5533 1787 5547
rect 5673 5533 5687 5547
rect 5753 5533 5767 5547
rect 6033 5533 6047 5547
rect 6133 5533 6147 5547
rect 6353 5533 6367 5547
rect 1933 5433 1947 5447
rect 1973 5432 1987 5446
rect 2913 5393 2927 5407
rect 953 5373 967 5387
rect 1253 5373 1267 5387
rect 1633 5373 1647 5387
rect 1933 5373 1947 5387
rect 1973 5373 1987 5387
rect 2973 5373 2987 5387
rect 5333 5373 5347 5387
rect 6213 5373 6227 5387
rect 913 5352 927 5366
rect 1193 5333 1207 5347
rect 1673 5333 1687 5347
rect 3973 5333 3987 5347
rect 4013 5333 4027 5347
rect 5293 5333 5307 5347
rect 6213 5333 6227 5347
rect 1033 5313 1047 5327
rect 1093 5313 1107 5327
rect 1433 5313 1447 5327
rect 1553 5313 1567 5327
rect 1893 5313 1907 5327
rect 1979 5313 1993 5327
rect 3413 5313 3427 5327
rect 3453 5313 3467 5327
rect 3613 5313 3627 5327
rect 3753 5313 3767 5327
rect 3913 5313 3927 5327
rect 4013 5312 4027 5326
rect 4093 5313 4107 5327
rect 4133 5313 4147 5327
rect 5533 5313 5547 5327
rect 5613 5313 5627 5327
rect 5853 5313 5867 5327
rect 5919 5313 5933 5327
rect 6013 5313 6027 5327
rect 6073 5311 6087 5325
rect 2173 5293 2187 5307
rect 2273 5293 2287 5307
rect 3273 5253 3287 5267
rect 3233 5233 3247 5247
rect 613 5113 627 5127
rect 153 5093 167 5107
rect 273 5093 287 5107
rect 553 5094 567 5108
rect 633 5093 647 5107
rect 473 5073 487 5087
rect 853 5093 867 5107
rect 953 5093 967 5107
rect 993 5093 1007 5107
rect 1113 5093 1127 5107
rect 1293 5093 1307 5107
rect 1333 5093 1347 5107
rect 2253 5093 2267 5107
rect 513 5033 527 5047
rect 1433 5073 1447 5087
rect 1733 5073 1747 5087
rect 2153 5073 2167 5087
rect 1473 5033 1487 5047
rect 1673 5033 1687 5047
rect 2153 5033 2167 5047
rect 2253 5033 2267 5047
rect 2333 5113 2347 5127
rect 2993 5113 3007 5127
rect 3053 5113 3067 5127
rect 2373 5093 2387 5107
rect 2393 5093 2407 5107
rect 2973 5093 2987 5107
rect 3073 5093 3087 5107
rect 3273 5093 3287 5107
rect 3353 5093 3367 5107
rect 3433 5093 3447 5107
rect 3493 5093 3507 5107
rect 4433 5093 4447 5107
rect 4493 5093 4507 5107
rect 4713 5093 4727 5107
rect 5507 5093 5521 5107
rect 5633 5093 5647 5107
rect 6193 5093 6207 5107
rect 2713 5073 2727 5087
rect 2773 5073 2787 5087
rect 3353 5072 3367 5086
rect 4133 5073 4147 5087
rect 3353 5033 3367 5047
rect 4133 5033 4147 5047
rect 4813 5073 4827 5087
rect 5953 5073 5967 5087
rect 6113 5073 6127 5087
rect 4733 5033 4747 5047
rect 4813 5033 4827 5047
rect 5913 5033 5927 5047
rect 6053 5033 6067 5047
rect 6213 5033 6227 5047
rect 633 5012 647 5026
rect 1573 5013 1587 5027
rect 1633 5013 1647 5027
rect 2273 5012 2287 5026
rect 5933 5013 5947 5027
rect 6013 5013 6027 5027
rect 1633 4893 1647 4907
rect 1673 4893 1687 4907
rect 4193 4893 4207 4907
rect 4253 4893 4267 4907
rect 33 4873 47 4887
rect 93 4874 107 4888
rect 333 4873 347 4887
rect 4973 4873 4987 4887
rect 5093 4873 5107 4887
rect 153 4853 167 4867
rect 153 4813 167 4827
rect 313 4813 327 4827
rect 373 4853 387 4867
rect 1153 4853 1167 4867
rect 1193 4853 1207 4867
rect 2033 4853 2047 4867
rect 2593 4853 2607 4867
rect 3933 4853 3947 4867
rect 4033 4853 4047 4867
rect 5833 4853 5847 4867
rect 5973 4853 5987 4867
rect 6113 4853 6127 4867
rect 373 4813 387 4827
rect 1973 4813 1987 4827
rect 2593 4813 2607 4827
rect 3933 4813 3947 4827
rect 4033 4813 4047 4827
rect 4353 4813 4367 4827
rect 4393 4813 4407 4827
rect 5873 4813 5887 4827
rect 6173 4853 6187 4867
rect 6233 4853 6247 4867
rect 6173 4813 6187 4827
rect 6233 4813 6247 4827
rect 1733 4793 1747 4807
rect 1793 4793 1807 4807
rect 1833 4793 1847 4807
rect 1913 4793 1927 4807
rect 2533 4793 2547 4807
rect 2653 4793 2667 4807
rect 3853 4793 3867 4807
rect 3973 4793 3987 4807
rect 4913 4793 4927 4807
rect 4953 4793 4967 4807
rect 5073 4793 5087 4807
rect 5553 4791 5567 4805
rect 5613 4793 5627 4807
rect 5853 4793 5867 4807
rect 5933 4793 5947 4807
rect 6033 4793 6047 4807
rect 6133 4793 6147 4807
rect 2713 4772 2727 4786
rect 2753 4773 2767 4787
rect 4033 4753 4047 4767
rect 4093 4753 4107 4767
rect 5973 4732 5987 4746
rect 6013 4733 6027 4747
rect 1153 4713 1167 4727
rect 1213 4712 1227 4726
rect 5813 4653 5827 4667
rect 5853 4653 5867 4667
rect 2033 4613 2047 4627
rect 2113 4613 2127 4627
rect 2653 4613 2667 4627
rect 2713 4613 2727 4627
rect 1593 4593 1607 4607
rect 1653 4593 1667 4607
rect 193 4573 207 4587
rect 293 4573 307 4587
rect 373 4573 387 4587
rect 593 4573 607 4587
rect 1273 4573 1287 4587
rect 1413 4574 1427 4588
rect 1453 4574 1467 4588
rect 1493 4573 1507 4587
rect 1593 4573 1607 4587
rect 1653 4572 1667 4586
rect 1753 4573 1767 4587
rect 393 4513 407 4527
rect 1473 4553 1487 4567
rect 1613 4553 1627 4567
rect 2133 4573 2147 4587
rect 2293 4574 2307 4588
rect 2453 4573 2467 4587
rect 1533 4513 1547 4527
rect 1613 4513 1627 4527
rect 1753 4513 1767 4527
rect 2353 4553 2367 4567
rect 2893 4553 2907 4567
rect 2113 4513 2127 4527
rect 2353 4513 2367 4527
rect 3093 4553 3107 4567
rect 3493 4573 3507 4587
rect 3973 4573 3987 4587
rect 4113 4573 4127 4587
rect 4193 4573 4207 4587
rect 4433 4573 4447 4587
rect 5073 4573 5087 4587
rect 5113 4573 5127 4587
rect 5273 4573 5287 4587
rect 5333 4573 5347 4587
rect 5433 4573 5447 4587
rect 5473 4573 5487 4587
rect 2933 4513 2947 4527
rect 3093 4513 3107 4527
rect 3413 4513 3427 4527
rect 3473 4553 3487 4567
rect 3473 4513 3487 4527
rect 3993 4513 4007 4527
rect 4373 4513 4387 4527
rect 5013 4553 5027 4567
rect 5393 4553 5407 4567
rect 4973 4513 4987 4527
rect 5673 4553 5687 4567
rect 5453 4513 5467 4527
rect 5673 4513 5687 4527
rect 5873 4553 5887 4567
rect 5933 4553 5947 4567
rect 6253 4553 6267 4567
rect 513 4493 527 4507
rect 1453 4493 1467 4507
rect 1493 4493 1507 4507
rect 2293 4493 2307 4507
rect 2393 4492 2407 4506
rect 3673 4493 3687 4507
rect 3733 4493 3747 4507
rect 3773 4493 3787 4507
rect 3853 4493 3867 4507
rect 3913 4493 3927 4507
rect 4033 4491 4047 4505
rect 5533 4493 5547 4507
rect 5613 4493 5627 4507
rect 5833 4493 5847 4507
rect 6253 4513 6267 4527
rect 5973 4492 5987 4506
rect 2573 4473 2587 4487
rect 2513 4453 2527 4467
rect 2573 4393 2587 4407
rect 2633 4393 2647 4407
rect 2373 4353 2387 4367
rect 3893 4353 3907 4367
rect 3953 4353 3967 4367
rect 4653 4353 4667 4367
rect 4713 4353 4727 4367
rect 4773 4353 4787 4367
rect 4833 4353 4847 4367
rect 4893 4353 4907 4367
rect 5673 4353 5687 4367
rect 5773 4353 5787 4367
rect 6353 4353 6367 4367
rect 6413 4353 6427 4367
rect 1753 4333 1767 4347
rect 1893 4333 1907 4347
rect 2193 4333 2207 4347
rect 1453 4293 1467 4307
rect 1493 4293 1507 4307
rect 1753 4293 1767 4307
rect 1073 4273 1087 4287
rect 1173 4273 1187 4287
rect 1213 4273 1227 4287
rect 1353 4273 1367 4287
rect 1393 4273 1407 4287
rect 1513 4273 1527 4287
rect 1693 4273 1707 4287
rect 1793 4273 1807 4287
rect 1853 4273 1867 4287
rect 2193 4293 2207 4307
rect 2253 4333 2267 4347
rect 2793 4333 2807 4347
rect 4513 4333 4527 4347
rect 5153 4333 5167 4347
rect 2253 4293 2267 4307
rect 2393 4293 2407 4307
rect 2793 4293 2807 4307
rect 4573 4293 4587 4307
rect 5153 4293 5167 4307
rect 5533 4293 5547 4307
rect 5573 4293 5587 4307
rect 3753 4273 3767 4287
rect 3813 4273 3827 4287
rect 4813 4273 4827 4287
rect 4853 4273 4867 4287
rect 5133 4271 5147 4285
rect 5233 4273 5247 4287
rect 2593 4252 2607 4266
rect 2633 4253 2647 4267
rect 3013 4253 3027 4267
rect 3113 4253 3127 4267
rect 5173 4253 5187 4267
rect 5233 4252 5247 4266
rect 2733 4212 2747 4226
rect 2793 4213 2807 4227
rect 3893 4193 3907 4207
rect 3933 4193 3947 4207
rect 3233 4113 3247 4127
rect 3273 4113 3287 4127
rect 1533 4093 1547 4107
rect 1633 4093 1647 4107
rect 1567 4076 1581 4090
rect 1613 4072 1627 4086
rect 173 4053 187 4067
rect 253 4053 267 4067
rect 453 4053 467 4067
rect 593 4053 607 4067
rect 913 4033 927 4047
rect 1113 4053 1127 4067
rect 1533 4053 1547 4067
rect 1573 4053 1587 4067
rect 3133 4053 3147 4067
rect 3193 4053 3207 4067
rect 3613 4054 3627 4068
rect 4753 4053 4767 4067
rect 4793 4053 4807 4067
rect 4993 4053 5007 4067
rect 5053 4053 5067 4067
rect 5193 4053 5207 4067
rect 5233 4053 5247 4067
rect 953 3993 967 4007
rect 1013 3993 1027 4007
rect 1213 4033 1227 4047
rect 1353 4033 1367 4047
rect 1433 4033 1447 4047
rect 1173 3993 1187 4007
rect 1353 3993 1367 4007
rect 2613 4033 2627 4047
rect 2713 4033 2727 4047
rect 2873 4033 2887 4047
rect 2973 4033 2987 4047
rect 3513 4033 3527 4047
rect 1453 3992 1467 4006
rect 2613 3993 2627 4007
rect 2713 3993 2727 4007
rect 3013 4012 3027 4026
rect 2913 3993 2927 4007
rect 3553 3993 3567 4007
rect 3633 3993 3647 4007
rect 4073 4033 4087 4047
rect 4233 4033 4247 4047
rect 6053 4033 6067 4047
rect 4073 3993 4087 4007
rect 4233 3993 4247 4007
rect 6053 3993 6067 4007
rect 2313 3973 2327 3987
rect 2353 3973 2367 3987
rect 2893 3973 2907 3987
rect 2933 3973 2947 3987
rect 5893 3973 5907 3987
rect 5959 3973 5973 3987
rect 13 3873 27 3887
rect 73 3873 87 3887
rect 4933 3853 4947 3867
rect 4973 3853 4987 3867
rect 5253 3853 5267 3867
rect 5313 3853 5327 3867
rect 393 3833 407 3847
rect 453 3833 467 3847
rect 2013 3833 2027 3847
rect 5673 3833 5687 3847
rect 5733 3833 5747 3847
rect 153 3813 167 3827
rect 733 3813 747 3827
rect 1053 3813 1067 3827
rect 1753 3813 1767 3827
rect 153 3773 167 3787
rect 1053 3773 1067 3787
rect 753 3752 767 3766
rect 1753 3759 1767 3773
rect 2253 3813 2267 3827
rect 2273 3792 2287 3806
rect 2313 3813 2327 3827
rect 2253 3773 2267 3787
rect 2833 3813 2847 3827
rect 4033 3812 4047 3826
rect 4613 3813 4627 3827
rect 5833 3813 5847 3827
rect 6113 3813 6127 3827
rect 2633 3773 2647 3787
rect 2673 3773 2687 3787
rect 2773 3773 2787 3787
rect 4073 3773 4087 3787
rect 4613 3773 4627 3787
rect 6273 3813 6287 3827
rect 6173 3773 6187 3787
rect 2013 3752 2027 3766
rect 2093 3753 2107 3767
rect 2173 3753 2187 3767
rect 3073 3753 3087 3767
rect 3133 3753 3147 3767
rect 3853 3753 3867 3767
rect 3913 3753 3927 3767
rect 3973 3753 3987 3767
rect 4333 3753 4347 3767
rect 4413 3753 4427 3767
rect 5533 3752 5547 3766
rect 5633 3753 5647 3767
rect 5873 3753 5887 3767
rect 5953 3753 5967 3767
rect 6073 3753 6087 3767
rect 6213 3753 6227 3767
rect 3733 3713 3747 3727
rect 3793 3693 3807 3707
rect 1593 3593 1607 3607
rect 1633 3593 1647 3607
rect 533 3573 547 3587
rect 573 3573 587 3587
rect 1693 3573 1707 3587
rect 1773 3573 1787 3587
rect 1253 3553 1267 3567
rect 1333 3553 1347 3567
rect 5433 3553 5447 3567
rect 5473 3553 5487 3567
rect 5513 3553 5527 3567
rect 673 3533 687 3547
rect 813 3533 827 3547
rect 1413 3534 1427 3548
rect 1493 3533 1507 3547
rect 1833 3534 1847 3548
rect 1873 3533 1887 3547
rect 1913 3533 1927 3547
rect 1953 3534 1967 3548
rect 253 3513 267 3527
rect 753 3513 767 3527
rect 1073 3513 1087 3527
rect 1173 3513 1187 3527
rect 1773 3513 1787 3527
rect 2973 3533 2987 3547
rect 3013 3533 3027 3547
rect 253 3473 267 3487
rect 693 3473 707 3487
rect 1013 3473 1027 3487
rect 1173 3473 1187 3487
rect 1593 3473 1607 3487
rect 1633 3473 1647 3487
rect 2133 3513 2147 3527
rect 2053 3473 2067 3487
rect 713 3453 727 3467
rect 753 3453 767 3467
rect 1693 3453 1707 3467
rect 1733 3453 1747 3467
rect 1793 3453 1807 3467
rect 1893 3453 1907 3467
rect 2113 3453 2127 3467
rect 2473 3513 2487 3527
rect 5993 3513 6007 3527
rect 2413 3473 2427 3487
rect 6053 3473 6067 3487
rect 1033 3433 1047 3447
rect 1073 3433 1087 3447
rect 453 3313 467 3327
rect 533 3313 547 3327
rect 893 3313 907 3327
rect 993 3313 1007 3327
rect 1213 3313 1227 3327
rect 1313 3313 1327 3327
rect 1393 3313 1407 3327
rect 313 3293 327 3307
rect 413 3294 427 3308
rect 313 3253 327 3267
rect 1433 3312 1447 3326
rect 353 3231 367 3245
rect 433 3233 447 3247
rect 913 3253 927 3267
rect 973 3253 987 3267
rect 1033 3293 1047 3307
rect 1173 3293 1187 3307
rect 1633 3293 1647 3307
rect 2073 3333 2087 3347
rect 5153 3333 5167 3347
rect 5213 3333 5227 3347
rect 2153 3313 2167 3327
rect 2233 3313 2247 3327
rect 2073 3293 2087 3307
rect 2193 3293 2207 3307
rect 3993 3293 4007 3307
rect 4013 3293 4027 3307
rect 4873 3293 4887 3307
rect 4973 3293 4987 3307
rect 1033 3253 1047 3267
rect 1173 3253 1187 3267
rect 1693 3253 1707 3267
rect 2233 3253 2247 3267
rect 4873 3253 4887 3267
rect 5853 3292 5867 3306
rect 5913 3292 5927 3306
rect 5033 3253 5047 3267
rect 533 3233 547 3247
rect 673 3233 687 3247
rect 813 3233 827 3247
rect 2273 3233 2287 3247
rect 2393 3233 2407 3247
rect 3853 3233 3867 3247
rect 3953 3233 3967 3247
rect 4013 3233 4027 3247
rect 4073 3233 4087 3247
rect 1713 3052 1727 3066
rect 1733 3053 1747 3067
rect 2313 3033 2327 3047
rect 2413 3033 2427 3047
rect 53 3008 67 3022
rect 273 3013 287 3027
rect 313 3013 327 3027
rect 413 3013 427 3027
rect 473 3013 487 3027
rect 973 3013 987 3027
rect 5813 3013 5827 3027
rect 5933 3013 5947 3027
rect 1033 2993 1047 3007
rect 1653 2993 1667 3007
rect 933 2953 947 2967
rect 1093 2953 1107 2967
rect 1973 2993 1987 3007
rect 2333 2993 2347 3007
rect 1713 2953 1727 2967
rect 1973 2953 1987 2967
rect 2113 2953 2127 2967
rect 2653 2993 2667 3007
rect 4073 2993 4087 3007
rect 5153 2993 5167 3007
rect 2393 2953 2407 2967
rect 2593 2953 2607 2967
rect 4073 2953 4087 2967
rect 33 2932 47 2946
rect 273 2933 287 2947
rect 373 2933 387 2947
rect 1773 2933 1787 2947
rect 1813 2933 1827 2947
rect 2033 2933 2047 2947
rect 2373 2933 2387 2947
rect 2413 2933 2427 2947
rect 5093 2933 5107 2947
rect 1233 2794 1247 2808
rect 1273 2793 1287 2807
rect 1093 2773 1107 2787
rect 1433 2773 1447 2787
rect 1593 2773 1607 2787
rect 3393 2773 3407 2787
rect 3453 2773 3467 2787
rect 5213 2773 5227 2787
rect 5273 2773 5287 2787
rect 193 2713 207 2727
rect 273 2713 287 2727
rect 433 2713 447 2727
rect 513 2713 527 2727
rect 573 2713 587 2727
rect 1053 2713 1067 2727
rect 1373 2733 1387 2747
rect 1533 2733 1547 2747
rect 3153 2733 3167 2747
rect 1353 2713 1367 2727
rect 1393 2713 1407 2727
rect 1473 2713 1487 2727
rect 1513 2713 1527 2727
rect 2713 2713 2727 2727
rect 2753 2711 2767 2725
rect 2793 2713 2807 2727
rect 2913 2713 2927 2727
rect 3093 2713 3107 2727
rect 4033 2711 4047 2725
rect 4073 2713 4087 2727
rect 1473 2692 1487 2706
rect 1553 2693 1567 2707
rect 493 2513 507 2527
rect 593 2513 607 2527
rect 1213 2513 1227 2527
rect 1253 2513 1267 2527
rect 413 2493 427 2507
rect 553 2493 567 2507
rect 1173 2493 1187 2507
rect 1253 2492 1267 2506
rect 1353 2493 1367 2507
rect 2513 2493 2527 2507
rect 2593 2493 2607 2507
rect 973 2473 987 2487
rect 1233 2473 1247 2487
rect 1193 2433 1207 2447
rect 933 2412 947 2426
rect 1753 2473 1767 2487
rect 2253 2473 2267 2487
rect 2633 2473 2647 2487
rect 3513 2473 3527 2487
rect 3553 2473 3567 2487
rect 1713 2433 1727 2447
rect 2093 2433 2107 2447
rect 2153 2433 2167 2447
rect 2253 2433 2267 2447
rect 2633 2433 2647 2447
rect 6273 2413 6287 2427
rect 6333 2413 6347 2427
rect 1333 2393 1347 2407
rect 2033 2313 2047 2327
rect 833 2293 847 2307
rect 873 2293 887 2307
rect 2007 2293 2021 2307
rect 2033 2292 2047 2306
rect 193 2273 207 2287
rect 1153 2273 1167 2287
rect 1253 2273 1267 2287
rect 1993 2272 2007 2286
rect 2513 2273 2527 2287
rect 2573 2273 2587 2287
rect 753 2253 767 2267
rect 1293 2253 1307 2267
rect 213 2213 227 2227
rect 753 2213 767 2227
rect 1453 2253 1467 2267
rect 1353 2213 1367 2227
rect 1453 2213 1467 2227
rect 1513 2253 1527 2267
rect 1713 2253 1727 2267
rect 2273 2253 2287 2267
rect 2593 2253 2607 2267
rect 2653 2253 2667 2267
rect 2793 2253 2807 2267
rect 3433 2253 3447 2267
rect 4173 2253 4187 2267
rect 1753 2213 1767 2227
rect 2313 2213 2327 2227
rect 2593 2213 2607 2227
rect 2693 2213 2707 2227
rect 2793 2213 2807 2227
rect 3433 2213 3447 2227
rect 4233 2213 4247 2227
rect 293 2193 307 2207
rect 433 2193 447 2207
rect 1333 2193 1347 2207
rect 1393 2193 1407 2207
rect 1473 2192 1487 2206
rect 1553 2193 1567 2207
rect 1653 2193 1667 2207
rect 1813 2193 1827 2207
rect 1893 2193 1907 2207
rect 1653 2153 1667 2167
rect 1613 2133 1627 2147
rect 493 2013 507 2027
rect 533 2013 547 2027
rect 1433 2013 1447 2027
rect 1513 2013 1527 2027
rect 2053 2012 2067 2026
rect 2093 2013 2107 2027
rect 313 1973 327 1987
rect 393 1972 407 1986
rect 493 1973 507 1987
rect 573 1973 587 1987
rect 773 1973 787 1987
rect 853 1973 867 1987
rect 1273 1974 1287 1988
rect 1393 1973 1407 1987
rect 3073 1973 3087 1987
rect 3253 1973 3267 1987
rect 3573 1973 3587 1987
rect 3673 1973 3687 1987
rect 5233 1973 5247 1987
rect 5273 1973 5287 1987
rect 1573 1953 1587 1967
rect 2373 1953 2387 1967
rect 2733 1953 2747 1967
rect 3613 1933 3627 1947
rect 153 1913 167 1927
rect 193 1913 207 1927
rect 1333 1913 1347 1927
rect 1573 1913 1587 1927
rect 2193 1913 2207 1927
rect 2233 1913 2247 1927
rect 2373 1913 2387 1927
rect 2733 1913 2747 1927
rect 3633 1913 3647 1927
rect 353 1893 367 1907
rect 393 1893 407 1907
rect 893 1893 907 1907
rect 933 1893 947 1907
rect 1733 1893 1747 1907
rect 1773 1893 1787 1907
rect 6113 1793 6127 1807
rect 6153 1793 6167 1807
rect 773 1753 787 1767
rect 853 1753 867 1767
rect 993 1753 1007 1767
rect 1053 1753 1067 1767
rect 1673 1754 1687 1768
rect 1733 1753 1747 1767
rect 2353 1753 2367 1767
rect 2653 1753 2667 1767
rect 2713 1753 2727 1767
rect 2813 1733 2827 1747
rect 2373 1693 2387 1707
rect 2833 1693 2847 1707
rect 673 1673 687 1687
rect 813 1673 827 1687
rect 1833 1673 1847 1687
rect 1953 1673 1967 1687
rect 3533 1671 3547 1685
rect 3613 1673 3627 1687
rect 3653 1673 3667 1687
rect 5153 1673 5167 1687
rect 5233 1671 5247 1685
rect 3493 1653 3507 1667
rect 113 1453 127 1467
rect 273 1453 287 1467
rect 553 1453 567 1467
rect 693 1453 707 1467
rect 733 1453 747 1467
rect 873 1453 887 1467
rect 913 1453 927 1467
rect 953 1453 967 1467
rect 1813 1453 1827 1467
rect 1913 1453 1927 1467
rect 1993 1453 2007 1467
rect 2413 1453 2427 1467
rect 2493 1454 2507 1468
rect 5273 1453 5287 1467
rect 5333 1453 5347 1467
rect 353 1433 367 1447
rect 1453 1433 1467 1447
rect 313 1393 327 1407
rect 2093 1433 2107 1447
rect 1493 1393 1507 1407
rect 2033 1393 2047 1407
rect 2853 1393 2867 1407
rect 2913 1373 2927 1387
rect 1973 1253 1987 1267
rect 2033 1253 2047 1267
rect 2553 1233 2567 1247
rect 3433 1233 3447 1247
rect 3533 1233 3547 1247
rect 3633 1233 3647 1247
rect 1333 1212 1347 1226
rect 1973 1213 1987 1227
rect 493 1173 507 1187
rect 1273 1173 1287 1187
rect 2033 1213 2047 1227
rect 2173 1213 2187 1227
rect 2273 1213 2287 1227
rect 393 1153 407 1167
rect 473 1153 487 1167
rect 1213 1153 1227 1167
rect 1313 1153 1327 1167
rect 1933 1153 1947 1167
rect 2033 1173 2047 1187
rect 2953 1213 2967 1227
rect 2093 1153 2107 1167
rect 2293 1153 2307 1167
rect 2473 1153 2487 1167
rect 2913 1173 2927 1187
rect 6253 1213 6267 1227
rect 2573 1153 2587 1167
rect 3573 1153 3587 1167
rect 6213 1173 6227 1187
rect 6053 1153 6067 1167
rect 6153 1153 6167 1167
rect 6233 1153 6247 1167
rect 6293 1153 6307 1167
rect 493 1133 507 1147
rect 553 933 567 947
rect 713 933 727 947
rect 973 933 987 947
rect 1113 933 1127 947
rect 2993 933 3007 947
rect 3033 933 3047 947
rect 3173 933 3187 947
rect 3233 933 3247 947
rect 153 913 167 927
rect 2893 913 2907 927
rect 4653 913 4667 927
rect 4693 913 4707 927
rect 153 873 167 887
rect 2893 873 2907 887
rect 2633 853 2647 867
rect 2733 853 2747 867
rect 5913 853 5927 867
rect 5973 853 5987 867
rect 1053 813 1067 827
rect 1093 813 1107 827
rect 273 713 287 727
rect 313 712 327 726
rect 1373 713 1387 727
rect 2213 713 2227 727
rect 2293 713 2307 727
rect 3233 713 3247 727
rect 3273 713 3287 727
rect 1433 693 1447 707
rect 1653 693 1667 707
rect 1693 693 1707 707
rect 3413 693 3427 707
rect 1373 653 1387 667
rect 3413 653 3427 667
rect 1413 633 1427 647
rect 1473 633 1487 647
rect 1893 633 1907 647
rect 1973 633 1987 647
rect 613 413 627 427
rect 653 413 667 427
rect 1033 413 1047 427
rect 1113 413 1127 427
rect 1513 413 1527 427
rect 1613 413 1627 427
rect 5093 413 5107 427
rect 5193 413 5207 427
rect 6093 413 6107 427
rect 6133 413 6147 427
rect 6173 413 6187 427
rect 6233 413 6247 427
rect 653 353 667 367
rect 693 353 707 367
rect 813 353 827 367
rect 853 353 867 367
rect 1213 333 1227 347
rect 1313 333 1327 347
rect 2233 333 2247 347
rect 2273 333 2287 347
rect 1313 193 1327 207
rect 2833 193 2847 207
rect 2873 193 2887 207
rect 273 173 287 187
rect 1273 173 1287 187
rect 1993 173 2007 187
rect 313 133 327 147
rect 1953 133 1967 147
rect 873 113 887 127
rect 953 113 967 127
rect 2313 113 2327 127
rect 2393 113 2407 127
rect 6313 113 6327 127
rect 6393 113 6407 127
<< metal2 >>
rect 2136 6267 2143 6303
rect 2176 6296 2203 6303
rect 416 6176 453 6183
rect 156 6116 163 6153
rect 256 6116 263 6153
rect 96 6080 103 6083
rect 93 6067 107 6080
rect 136 6007 143 6083
rect 56 5807 63 5933
rect 96 5860 103 5863
rect 93 5847 107 5860
rect 136 5807 143 5863
rect 156 5427 163 5833
rect 176 5607 183 5853
rect 196 5847 203 6114
rect 236 6047 243 6073
rect 276 6007 283 6083
rect 316 6063 323 6083
rect 316 6056 343 6063
rect 236 5896 243 5933
rect 276 5896 283 5933
rect 316 5903 323 6033
rect 336 5927 343 6056
rect 356 6007 363 6133
rect 376 6087 383 6153
rect 416 6147 423 6176
rect 436 6116 443 6153
rect 496 6127 503 6153
rect 516 6087 523 6173
rect 596 6116 603 6193
rect 456 5987 463 6083
rect 536 6083 543 6114
rect 536 6076 563 6083
rect 496 6007 503 6053
rect 436 5976 453 5983
rect 316 5896 343 5903
rect 336 5867 343 5896
rect 193 5608 207 5614
rect 256 5556 283 5563
rect 173 5547 187 5552
rect 216 5507 223 5552
rect 256 5376 263 5533
rect 276 5387 283 5556
rect 296 5547 303 5852
rect 316 5608 323 5853
rect 356 5807 363 5953
rect 436 5896 443 5976
rect 476 5907 483 5933
rect 460 5863 473 5867
rect 456 5856 473 5863
rect 460 5853 473 5856
rect 496 5627 503 5993
rect 516 5907 523 6052
rect 536 5896 543 5953
rect 556 5928 563 6076
rect 616 6067 623 6083
rect 616 6056 633 6067
rect 620 6053 633 6056
rect 613 5967 627 5973
rect 656 5967 663 6073
rect 676 5987 683 6193
rect 1036 6167 1043 6193
rect 696 6087 703 6153
rect 776 6116 783 6153
rect 916 6128 923 6153
rect 1036 6116 1043 6153
rect 1276 6116 1283 6213
rect 1416 6187 1423 6213
rect 653 5943 667 5953
rect 636 5940 667 5943
rect 673 5947 687 5952
rect 636 5936 663 5940
rect 607 5913 613 5927
rect 516 5628 523 5853
rect 636 5863 643 5936
rect 716 5896 723 5993
rect 736 5907 743 6053
rect 796 6027 803 6083
rect 836 5987 843 6114
rect 936 6027 943 6083
rect 596 5856 643 5863
rect 696 5707 703 5863
rect 756 5847 763 5973
rect 796 5907 803 5973
rect 816 5896 823 5933
rect 856 5896 863 5993
rect 876 5860 883 5863
rect 836 5827 843 5852
rect 873 5847 887 5860
rect 393 5600 407 5613
rect 396 5596 403 5600
rect 456 5566 463 5613
rect 553 5600 567 5613
rect 556 5596 563 5600
rect 596 5566 603 5613
rect 696 5596 703 5693
rect 336 5507 343 5552
rect 16 4747 23 5133
rect 56 5107 63 5333
rect 156 5107 163 5374
rect 56 5046 63 5093
rect 153 5080 167 5093
rect 196 5088 203 5343
rect 296 5167 303 5473
rect 416 5427 423 5563
rect 496 5507 503 5563
rect 536 5487 543 5552
rect 616 5447 623 5594
rect 776 5567 783 5633
rect 376 5376 383 5413
rect 156 5076 163 5080
rect 233 5080 247 5093
rect 273 5088 287 5093
rect 236 5076 243 5080
rect 316 5083 323 5373
rect 356 5107 363 5343
rect 456 5343 463 5374
rect 456 5336 483 5343
rect 376 5083 383 5153
rect 316 5076 343 5083
rect 196 5047 203 5074
rect 16 3967 23 4733
rect 36 4526 43 4873
rect 56 4867 63 4993
rect 96 4888 103 5043
rect 140 4863 153 4867
rect 136 4856 153 4863
rect 140 4854 153 4856
rect 156 4607 163 4813
rect 176 4787 183 4854
rect 196 4826 203 4953
rect 256 4927 263 5032
rect 296 4907 303 5043
rect 316 4947 323 5033
rect 336 4887 343 5076
rect 356 5076 383 5083
rect 416 5076 423 5133
rect 456 5076 463 5213
rect 476 5087 483 5336
rect 516 5087 523 5343
rect 556 5108 563 5343
rect 576 5223 583 5333
rect 596 5267 603 5413
rect 676 5407 683 5552
rect 876 5527 883 5812
rect 916 5807 923 5894
rect 936 5847 943 5992
rect 996 5908 1003 6093
rect 1056 6080 1063 6083
rect 1053 6067 1067 6080
rect 1096 6047 1103 6083
rect 1196 5967 1203 6083
rect 1296 6007 1303 6083
rect 1316 5983 1323 6053
rect 1296 5976 1323 5983
rect 1036 5896 1043 5953
rect 976 5827 983 5863
rect 1016 5860 1023 5863
rect 1013 5847 1027 5860
rect 1047 5833 1053 5847
rect 1076 5827 1083 5894
rect 1236 5866 1243 5953
rect 1296 5896 1303 5976
rect 1336 5927 1343 5993
rect 1336 5896 1343 5913
rect 1116 5860 1123 5863
rect 1113 5847 1127 5860
rect 1156 5807 1163 5863
rect 1396 5863 1403 6153
rect 1496 6086 1503 6153
rect 1436 5947 1443 5993
rect 1456 5987 1463 6083
rect 1516 6067 1523 6233
rect 1576 6116 1583 6173
rect 1596 6080 1603 6083
rect 1593 6067 1607 6080
rect 1656 6067 1663 6114
rect 1676 6086 1683 6193
rect 1736 6116 1743 6153
rect 1976 6147 1983 6193
rect 1996 6187 2003 6213
rect 1796 6087 1803 6114
rect 1996 6116 2003 6173
rect 2013 6147 2027 6153
rect 2036 6128 2043 6193
rect 1936 6083 1943 6113
rect 1753 6067 1767 6072
rect 1856 6063 1863 6083
rect 1856 6056 1883 6063
rect 1727 6033 1733 6047
rect 1696 6007 1703 6033
rect 1396 5856 1423 5863
rect 1476 5860 1483 5863
rect 1473 5847 1487 5860
rect 1496 5807 1503 5894
rect 947 5633 953 5647
rect 976 5596 983 5653
rect 1007 5603 1020 5607
rect 1007 5593 1023 5603
rect 696 5376 703 5473
rect 576 5216 593 5223
rect 316 4607 323 4813
rect 116 4568 123 4593
rect 336 4587 343 4852
rect 193 4568 207 4573
rect 253 4560 267 4573
rect 293 4560 307 4573
rect 256 4556 263 4560
rect 296 4556 303 4560
rect 56 4347 63 4393
rect 76 4336 83 4513
rect 136 4407 143 4523
rect 176 4387 183 4513
rect 13 3887 27 3893
rect 16 3627 23 3852
rect 16 2707 23 3133
rect 36 2967 43 4073
rect 56 4006 63 4293
rect 136 4267 143 4303
rect 176 4067 183 4333
rect 196 4087 203 4554
rect 276 4520 283 4523
rect 273 4507 287 4520
rect 276 4348 283 4493
rect 316 4487 323 4523
rect 336 4407 343 4513
rect 356 4447 363 5076
rect 596 5076 603 5213
rect 616 5127 623 5373
rect 656 5187 663 5253
rect 716 5207 723 5343
rect 396 5007 403 5043
rect 376 4867 383 4893
rect 396 4887 403 4993
rect 436 4987 443 5043
rect 416 4856 423 4933
rect 456 4856 463 4893
rect 376 4587 383 4813
rect 396 4747 403 4823
rect 496 4823 503 5073
rect 636 5047 643 5093
rect 516 4967 523 5033
rect 576 5007 583 5043
rect 596 4907 603 5013
rect 596 4856 603 4893
rect 496 4816 543 4823
rect 376 4487 383 4552
rect 516 4523 523 4816
rect 593 4560 607 4573
rect 636 4568 643 5012
rect 656 4887 663 5173
rect 756 5147 763 5373
rect 776 5207 783 5433
rect 916 5387 923 5563
rect 956 5560 963 5563
rect 953 5547 967 5560
rect 676 5087 683 5133
rect 753 5080 767 5093
rect 756 5076 763 5080
rect 736 5040 743 5043
rect 696 5007 703 5032
rect 733 5027 747 5040
rect 796 5007 803 5313
rect 836 5267 843 5343
rect 876 5307 883 5343
rect 916 5227 923 5352
rect 936 5327 943 5513
rect 1016 5447 1023 5593
rect 1036 5563 1043 5793
rect 1516 5727 1523 5913
rect 1596 5896 1603 5933
rect 1576 5807 1583 5863
rect 1616 5860 1643 5863
rect 1613 5856 1643 5860
rect 1613 5847 1627 5856
rect 1056 5647 1063 5673
rect 1096 5596 1103 5653
rect 1036 5556 1063 5563
rect 1056 5487 1063 5556
rect 1076 5527 1083 5563
rect 1116 5553 1124 5563
rect 1113 5547 1127 5553
rect 1176 5527 1183 5613
rect 1196 5608 1203 5633
rect 1233 5600 1247 5613
rect 1236 5596 1243 5600
rect 1356 5607 1363 5713
rect 1196 5563 1203 5594
rect 1336 5567 1343 5594
rect 1396 5596 1403 5633
rect 1416 5627 1423 5673
rect 1436 5608 1443 5653
rect 1496 5627 1503 5653
rect 1576 5596 1623 5603
rect 1196 5556 1223 5563
rect 1076 5456 1123 5463
rect 967 5383 980 5387
rect 967 5376 983 5383
rect 967 5374 980 5376
rect 996 5340 1003 5343
rect 1036 5340 1043 5343
rect 993 5327 1007 5340
rect 1033 5327 1047 5340
rect 1076 5327 1083 5456
rect 1096 5387 1103 5433
rect 1116 5427 1123 5456
rect 1216 5347 1223 5556
rect 1036 5267 1043 5313
rect 1093 5307 1107 5313
rect 853 5088 867 5093
rect 893 5088 907 5094
rect 696 4856 703 4953
rect 676 4787 683 4823
rect 596 4556 603 4560
rect 393 4507 407 4513
rect 416 4503 423 4523
rect 456 4520 463 4523
rect 453 4507 467 4520
rect 416 4496 443 4503
rect 336 4303 343 4393
rect 416 4336 423 4393
rect 436 4367 443 4496
rect 496 4516 523 4523
rect 456 4336 463 4373
rect 256 4267 263 4303
rect 296 4296 343 4303
rect 133 4040 147 4053
rect 136 4036 143 4040
rect 196 4003 203 4034
rect 56 3827 63 3893
rect 76 3887 83 3913
rect 113 3820 127 3833
rect 156 3827 163 4003
rect 176 3996 203 4003
rect 176 3847 183 3996
rect 216 3983 223 4253
rect 253 4040 267 4053
rect 296 4048 303 4213
rect 256 4036 263 4040
rect 196 3976 223 3983
rect 116 3816 123 3820
rect 196 3823 203 3976
rect 176 3816 203 3823
rect 216 3816 223 3953
rect 96 3780 103 3783
rect 76 3667 83 3773
rect 93 3767 107 3780
rect 136 3727 143 3783
rect 156 3607 163 3773
rect 176 3747 183 3816
rect 276 3747 283 3783
rect 196 3528 203 3713
rect 176 3516 193 3523
rect 216 3503 223 3733
rect 196 3496 223 3503
rect 116 3367 123 3443
rect 56 3022 63 3353
rect 93 3300 107 3313
rect 136 3307 143 3353
rect 96 3296 103 3300
rect 116 3227 123 3263
rect 136 3087 143 3253
rect 156 3147 163 3333
rect 196 3296 203 3496
rect 236 3367 243 3553
rect 256 3527 263 3633
rect 316 3567 323 4003
rect 356 3907 363 4133
rect 416 4048 423 4273
rect 436 4087 443 4303
rect 496 4303 503 4516
rect 576 4520 583 4523
rect 513 4487 527 4493
rect 536 4387 543 4513
rect 573 4507 587 4520
rect 616 4467 623 4523
rect 656 4507 663 4593
rect 756 4587 763 4873
rect 816 4856 823 4973
rect 836 4887 843 5043
rect 876 5040 883 5043
rect 873 5027 887 5040
rect 936 4987 943 5193
rect 967 5093 973 5107
rect 993 5080 1007 5093
rect 1033 5080 1047 5093
rect 996 5076 1003 5080
rect 1036 5076 1043 5080
rect 1076 5046 1083 5113
rect 976 5007 983 5043
rect 1013 5026 1027 5032
rect 896 4827 903 4854
rect 713 4560 727 4573
rect 760 4563 773 4567
rect 716 4556 723 4560
rect 756 4556 773 4563
rect 760 4553 773 4556
rect 696 4447 703 4523
rect 496 4296 523 4303
rect 476 4227 483 4293
rect 453 4040 467 4053
rect 456 4036 463 4040
rect 396 3847 403 4003
rect 496 3947 503 4153
rect 416 3827 423 3873
rect 396 3816 413 3823
rect 336 3783 343 3814
rect 336 3776 363 3783
rect 356 3707 363 3776
rect 356 3647 363 3693
rect 256 3427 263 3473
rect 396 3483 403 3753
rect 387 3476 403 3483
rect 176 3167 183 3253
rect 216 3227 223 3263
rect 256 3147 263 3263
rect 276 3047 283 3253
rect 133 3008 147 3014
rect 16 1706 23 2513
rect 36 2488 43 2932
rect 76 2927 83 2963
rect 176 2827 183 3033
rect 273 3027 287 3033
rect 296 3027 303 3313
rect 316 3307 323 3373
rect 336 3347 343 3443
rect 376 3327 383 3413
rect 376 3296 383 3313
rect 416 3308 423 3733
rect 456 3527 463 3833
rect 516 3816 523 4296
rect 596 4067 603 4293
rect 616 4067 623 4373
rect 716 4336 723 4493
rect 736 4427 743 4523
rect 796 4507 803 4812
rect 836 4667 843 4823
rect 916 4823 923 4913
rect 916 4816 943 4823
rect 996 4820 1003 4823
rect 993 4807 1007 4820
rect 876 4587 883 4653
rect 896 4556 903 4693
rect 936 4567 943 4793
rect 1016 4747 1023 4973
rect 1096 4967 1103 5293
rect 1136 5127 1143 5313
rect 1156 5287 1163 5343
rect 1196 5307 1203 5333
rect 1236 5303 1243 5513
rect 1256 5487 1263 5563
rect 1296 5543 1303 5563
rect 1276 5536 1303 5543
rect 1276 5423 1283 5536
rect 1476 5427 1483 5594
rect 1256 5416 1283 5423
rect 1256 5387 1263 5416
rect 1293 5380 1307 5393
rect 1296 5376 1303 5380
rect 1216 5296 1243 5303
rect 1127 5103 1140 5107
rect 1127 5093 1143 5103
rect 1136 5076 1143 5093
rect 1196 4987 1203 5113
rect 1216 5088 1223 5296
rect 1276 5227 1283 5332
rect 1316 5287 1323 5332
rect 1376 5287 1383 5374
rect 1516 5346 1523 5413
rect 1436 5340 1443 5343
rect 1433 5327 1447 5340
rect 1536 5323 1543 5453
rect 1556 5387 1563 5563
rect 1616 5467 1623 5596
rect 1636 5387 1643 5856
rect 1656 5827 1663 5933
rect 1676 5707 1683 5953
rect 1756 5896 1763 5953
rect 1667 5656 1713 5663
rect 1736 5647 1743 5863
rect 1776 5827 1783 5863
rect 1816 5767 1823 6053
rect 1876 5908 1883 6056
rect 1896 6047 1903 6083
rect 1916 6076 1943 6083
rect 1916 5896 1923 6076
rect 1976 6023 1983 6073
rect 2016 6047 2023 6083
rect 2056 6047 2063 6083
rect 1956 6016 1983 6023
rect 1856 5827 1863 5863
rect 1896 5767 1903 5863
rect 1956 5827 1963 6016
rect 1996 5827 2003 5863
rect 2036 5827 2043 5863
rect 1787 5653 1793 5667
rect 1676 5596 1683 5633
rect 1696 5547 1703 5563
rect 1696 5536 1713 5547
rect 1700 5533 1713 5536
rect 1656 5343 1663 5493
rect 1676 5387 1683 5533
rect 1756 5507 1763 5633
rect 1776 5608 1783 5632
rect 1856 5596 1863 5693
rect 1916 5627 1923 5813
rect 1776 5547 1783 5594
rect 1696 5376 1703 5413
rect 1536 5316 1553 5323
rect 1233 5080 1247 5093
rect 1293 5080 1307 5093
rect 1236 5076 1243 5080
rect 1296 5076 1303 5080
rect 1216 5046 1223 5074
rect 1256 4927 1263 5043
rect 1316 4923 1323 5074
rect 1336 4987 1343 5093
rect 1436 5087 1443 5213
rect 1500 5103 1513 5107
rect 1496 5093 1513 5103
rect 1496 5076 1503 5093
rect 1536 5076 1543 5113
rect 1556 5087 1563 5313
rect 1576 5207 1583 5343
rect 1616 5336 1663 5343
rect 1673 5323 1687 5333
rect 1673 5320 1703 5323
rect 1676 5316 1703 5320
rect 1396 4967 1403 5043
rect 1456 4987 1463 5074
rect 1307 4916 1323 4923
rect 816 4487 823 4554
rect 916 4520 923 4523
rect 913 4507 927 4520
rect 836 4336 843 4373
rect 876 4307 883 4473
rect 787 4296 823 4303
rect 596 4036 603 4053
rect 676 4006 683 4053
rect 776 4047 783 4193
rect 876 4087 883 4293
rect 896 4187 903 4433
rect 936 4407 943 4513
rect 956 4467 963 4633
rect 976 4447 983 4733
rect 996 4556 1003 4673
rect 1036 4647 1043 4893
rect 1140 4863 1153 4867
rect 1136 4856 1153 4863
rect 1140 4854 1153 4856
rect 1076 4787 1083 4823
rect 1056 4523 1063 4733
rect 1116 4727 1123 4823
rect 1156 4727 1163 4773
rect 1176 4767 1183 4854
rect 1207 4854 1213 4867
rect 1296 4856 1303 4913
rect 1207 4853 1220 4854
rect 1336 4826 1343 4853
rect 1456 4827 1463 4854
rect 1036 4516 1063 4523
rect 953 4340 967 4353
rect 956 4336 963 4340
rect 996 4287 1003 4353
rect 1036 4343 1043 4516
rect 1076 4447 1083 4673
rect 1096 4527 1103 4613
rect 1156 4583 1163 4713
rect 1176 4687 1183 4753
rect 1216 4747 1223 4793
rect 1236 4787 1243 4823
rect 1136 4576 1163 4583
rect 1136 4556 1143 4576
rect 1176 4556 1183 4673
rect 1196 4563 1203 4653
rect 1216 4587 1223 4712
rect 1196 4556 1223 4563
rect 1273 4560 1287 4573
rect 1276 4556 1283 4560
rect 1216 4523 1223 4556
rect 1216 4516 1263 4523
rect 1296 4503 1303 4523
rect 1276 4496 1303 4503
rect 1016 4336 1043 4343
rect 1056 4336 1063 4393
rect 496 3516 503 3593
rect 516 3587 523 3653
rect 536 3587 543 3783
rect 316 3043 323 3253
rect 436 3247 443 3472
rect 476 3347 483 3483
rect 536 3327 543 3453
rect 556 3427 563 3473
rect 576 3447 583 3573
rect 596 3527 603 3873
rect 616 3787 623 4003
rect 696 3996 723 4003
rect 696 3967 703 3996
rect 636 3887 643 3913
rect 656 3816 663 3893
rect 636 3747 643 3783
rect 696 3780 703 3783
rect 693 3767 707 3780
rect 716 3727 723 3973
rect 796 3967 803 4073
rect 853 4040 867 4053
rect 900 4043 913 4047
rect 856 4036 863 4040
rect 896 4036 913 4043
rect 900 4033 913 4036
rect 836 3907 843 4003
rect 733 3827 747 3833
rect 756 3787 763 3893
rect 616 3667 623 3693
rect 673 3520 687 3533
rect 676 3516 683 3520
rect 616 3447 623 3483
rect 656 3447 663 3483
rect 696 3383 703 3473
rect 716 3467 723 3514
rect 676 3376 703 3383
rect 456 3266 463 3313
rect 513 3300 527 3313
rect 516 3296 523 3300
rect 556 3296 563 3373
rect 576 3307 583 3333
rect 676 3327 683 3376
rect 600 3303 613 3307
rect 596 3293 613 3303
rect 696 3296 703 3353
rect 716 3307 723 3413
rect 736 3407 743 3773
rect 833 3766 847 3772
rect 756 3527 763 3752
rect 876 3707 883 3873
rect 896 3786 903 3853
rect 916 3827 923 3992
rect 936 3947 943 4053
rect 1016 4043 1023 4336
rect 1076 4300 1083 4303
rect 1073 4287 1087 4300
rect 1116 4287 1123 4303
rect 1016 4036 1043 4043
rect 956 3927 963 3993
rect 956 3816 963 3853
rect 976 3847 983 3873
rect 996 3828 1003 3973
rect 1016 3907 1023 3993
rect 813 3528 827 3533
rect 467 3256 503 3263
rect 536 3260 543 3263
rect 533 3247 547 3260
rect 316 3036 343 3043
rect 313 3003 327 3013
rect 296 3000 327 3003
rect 296 2996 323 3000
rect 196 2887 203 2994
rect 236 2927 243 2963
rect 276 2960 283 2963
rect 273 2947 287 2960
rect 187 2816 203 2823
rect 136 2776 143 2813
rect 56 2446 63 2773
rect 116 2627 123 2743
rect 196 2727 203 2816
rect 216 2787 223 2833
rect 256 2827 263 2873
rect 276 2847 283 2933
rect 256 2776 263 2813
rect 296 2788 303 2933
rect 336 2867 343 3036
rect 356 2847 363 3231
rect 473 3027 487 3033
rect 413 3000 427 3013
rect 453 3000 467 3013
rect 416 2996 423 3000
rect 456 2996 463 3000
rect 396 2947 403 2963
rect 436 2960 443 2963
rect 387 2936 403 2947
rect 433 2947 447 2960
rect 387 2933 400 2936
rect 347 2823 360 2827
rect 347 2813 363 2823
rect 276 2740 283 2743
rect 273 2727 287 2740
rect 196 2627 203 2653
rect 156 2476 163 2553
rect 36 1926 43 2353
rect 56 1968 63 2293
rect 76 2263 83 2353
rect 96 2287 103 2443
rect 196 2287 203 2613
rect 216 2527 223 2573
rect 276 2476 283 2553
rect 296 2387 303 2443
rect 336 2427 343 2773
rect 356 2746 363 2813
rect 456 2776 463 2893
rect 496 2807 503 3153
rect 596 3047 603 3293
rect 553 3000 567 3013
rect 556 2996 563 3000
rect 596 2996 603 3033
rect 616 3003 623 3253
rect 636 3207 643 3263
rect 676 3260 683 3263
rect 673 3247 687 3260
rect 616 2996 643 3003
rect 536 2907 543 2963
rect 576 2947 583 2963
rect 436 2740 443 2743
rect 76 2256 103 2263
rect 236 2256 243 2293
rect 276 2256 283 2293
rect 296 2287 303 2373
rect 156 2216 173 2223
rect 76 1987 83 2033
rect 116 1983 123 2212
rect 96 1976 123 1983
rect 96 1956 103 1976
rect 136 1956 143 1993
rect 56 1406 63 1773
rect 116 1736 123 1773
rect 156 1736 163 1913
rect 176 1903 183 2212
rect 196 2127 203 2252
rect 216 2103 223 2213
rect 293 2207 307 2212
rect 196 2096 223 2103
rect 196 1927 203 2096
rect 236 1956 243 2013
rect 336 2007 343 2392
rect 313 1967 327 1973
rect 176 1896 203 1903
rect 96 1683 103 1692
rect 96 1676 123 1683
rect 116 1467 123 1676
rect 136 1647 143 1703
rect 116 1436 123 1453
rect 16 467 23 1313
rect 96 1247 103 1403
rect 136 1367 143 1392
rect 196 1343 203 1896
rect 216 1847 223 1913
rect 296 1920 303 1923
rect 293 1907 307 1920
rect 216 1667 223 1773
rect 276 1736 323 1743
rect 256 1647 263 1703
rect 316 1683 323 1736
rect 336 1703 343 1993
rect 356 1907 363 2732
rect 433 2727 447 2740
rect 416 2507 423 2693
rect 476 2567 483 2733
rect 496 2547 503 2793
rect 516 2727 523 2853
rect 536 2783 543 2893
rect 576 2867 583 2933
rect 636 2887 643 2996
rect 536 2776 563 2783
rect 593 2780 607 2793
rect 596 2776 603 2780
rect 576 2740 583 2743
rect 416 2476 423 2493
rect 456 2476 463 2533
rect 493 2527 507 2533
rect 396 2367 403 2443
rect 436 2440 443 2443
rect 433 2427 447 2440
rect 416 2307 423 2353
rect 416 2256 423 2293
rect 456 2256 463 2313
rect 396 2007 403 2223
rect 436 2220 443 2223
rect 433 2207 447 2220
rect 436 2027 443 2153
rect 496 2027 503 2473
rect 516 2407 523 2513
rect 536 2487 543 2733
rect 573 2727 587 2740
rect 616 2667 623 2743
rect 656 2647 663 3233
rect 716 2996 723 3073
rect 736 3027 743 3313
rect 756 3308 763 3453
rect 796 3447 803 3483
rect 876 3427 883 3653
rect 936 3647 943 3772
rect 1036 3747 1043 4036
rect 1056 3987 1063 4173
rect 1116 4067 1123 4273
rect 1156 4067 1163 4433
rect 1276 4367 1283 4496
rect 1296 4303 1303 4393
rect 1216 4287 1223 4303
rect 1256 4296 1303 4303
rect 1187 4273 1193 4287
rect 1176 4047 1183 4213
rect 1160 4003 1173 4006
rect 1116 3927 1123 4003
rect 1156 3996 1173 4003
rect 1160 3993 1173 3996
rect 1067 3823 1080 3827
rect 1067 3816 1083 3823
rect 1067 3813 1080 3816
rect 1056 3607 1063 3773
rect 1156 3667 1163 3973
rect 1176 3787 1183 3873
rect 1196 3807 1203 4053
rect 1216 4047 1223 4273
rect 1316 4167 1323 4473
rect 1336 4407 1343 4513
rect 1356 4463 1363 4693
rect 1376 4627 1383 4812
rect 1396 4563 1403 4673
rect 1416 4667 1423 4823
rect 1427 4578 1453 4585
rect 1476 4567 1483 5033
rect 1576 5027 1583 5193
rect 1496 4823 1503 4893
rect 1496 4816 1523 4823
rect 1516 4747 1523 4816
rect 1516 4627 1523 4733
rect 1556 4727 1563 4793
rect 1576 4667 1583 4791
rect 1596 4727 1603 5133
rect 1656 5076 1663 5293
rect 1636 5040 1643 5043
rect 1633 5027 1647 5040
rect 1616 4707 1623 4913
rect 1676 4907 1683 5033
rect 1696 4967 1703 5316
rect 1716 5307 1723 5332
rect 1756 5247 1763 5343
rect 1796 5287 1803 5513
rect 1836 5427 1843 5563
rect 1876 5527 1883 5563
rect 1876 5376 1883 5492
rect 1916 5427 1923 5613
rect 1936 5447 1943 5793
rect 1996 5596 2003 5693
rect 1976 5467 1983 5563
rect 2036 5527 2043 5753
rect 2096 5707 2103 6253
rect 2136 6023 2143 6153
rect 2196 6116 2203 6296
rect 2767 6236 2803 6243
rect 2356 6167 2363 6213
rect 2116 6016 2143 6023
rect 2116 5727 2123 6016
rect 2216 6007 2223 6153
rect 2353 6120 2367 6132
rect 2356 6116 2363 6120
rect 2256 6083 2263 6114
rect 2256 6076 2283 6083
rect 2156 5896 2163 5933
rect 2236 5927 2243 6073
rect 2256 5987 2263 6033
rect 2276 6027 2283 6076
rect 2296 6047 2303 6083
rect 2396 6047 2403 6193
rect 2416 6047 2423 6233
rect 2436 6027 2443 6153
rect 2456 6087 2463 6193
rect 2476 6116 2483 6233
rect 2760 6223 2773 6227
rect 2756 6220 2773 6223
rect 2753 6213 2773 6220
rect 2753 6207 2767 6213
rect 2736 6176 2773 6183
rect 2516 6080 2523 6083
rect 2576 6080 2583 6083
rect 2513 6067 2527 6080
rect 2573 6067 2587 6080
rect 2616 6067 2623 6153
rect 2736 6147 2743 6176
rect 2756 6116 2763 6153
rect 2796 6147 2803 6236
rect 2873 6120 2887 6133
rect 2876 6116 2883 6120
rect 2276 5907 2283 5953
rect 2327 5914 2333 5927
rect 2356 5896 2363 6013
rect 2316 5891 2324 5894
rect 2136 5747 2143 5853
rect 2213 5847 2227 5852
rect 2173 5827 2187 5831
rect 2196 5767 2203 5833
rect 2220 5826 2240 5827
rect 2227 5813 2233 5826
rect 2256 5747 2263 5852
rect 2133 5600 2147 5613
rect 2136 5596 2143 5600
rect 1976 5387 1983 5432
rect 1896 5327 1903 5343
rect 1896 5247 1903 5313
rect 1936 5287 1943 5373
rect 1956 5267 1963 5374
rect 2056 5376 2063 5553
rect 2076 5467 2083 5563
rect 2116 5507 2123 5563
rect 2176 5487 2183 5693
rect 2296 5567 2303 5831
rect 2336 5767 2343 5863
rect 2396 5787 2403 6012
rect 2476 5967 2483 6053
rect 2580 6046 2593 6047
rect 2587 6033 2593 6046
rect 2616 6027 2623 6053
rect 2696 6047 2703 6083
rect 2736 6080 2743 6083
rect 2733 6067 2747 6080
rect 2676 6007 2683 6033
rect 2316 5587 2323 5713
rect 2196 5467 2203 5553
rect 2236 5527 2243 5563
rect 2316 5507 2323 5573
rect 2136 5376 2143 5413
rect 1996 5340 2003 5343
rect 1993 5327 2007 5340
rect 1716 5127 1723 5173
rect 1736 5087 1743 5113
rect 1716 4907 1723 5074
rect 1936 5076 1943 5113
rect 1976 5087 1983 5233
rect 1736 5036 1763 5043
rect 1796 5040 1803 5043
rect 1736 4987 1743 5036
rect 1793 5027 1807 5040
rect 1636 4827 1643 4893
rect 1713 4860 1727 4872
rect 1716 4856 1723 4860
rect 1733 4807 1747 4813
rect 1376 4556 1403 4563
rect 1376 4487 1383 4556
rect 1396 4487 1403 4513
rect 1496 4507 1503 4573
rect 1516 4527 1523 4613
rect 1556 4596 1593 4603
rect 1556 4556 1563 4596
rect 1587 4573 1593 4587
rect 1616 4567 1623 4653
rect 1636 4527 1643 4773
rect 1756 4723 1763 5013
rect 1856 4827 1863 5074
rect 1916 5040 1923 5043
rect 1913 5027 1927 5040
rect 1776 4787 1783 4813
rect 1916 4820 1923 4823
rect 1913 4807 1927 4820
rect 1807 4796 1833 4803
rect 1756 4716 1783 4723
rect 1656 4607 1663 4653
rect 1653 4567 1667 4572
rect 1676 4556 1683 4613
rect 1696 4583 1703 4713
rect 1716 4627 1723 4673
rect 1753 4587 1767 4593
rect 1696 4576 1723 4583
rect 1716 4556 1723 4576
rect 1753 4567 1767 4573
rect 1776 4527 1783 4716
rect 1356 4456 1383 4463
rect 1376 4336 1383 4456
rect 1416 4336 1423 4453
rect 1436 4347 1443 4490
rect 1456 4307 1463 4493
rect 1356 4300 1363 4303
rect 1396 4300 1403 4303
rect 1336 4187 1343 4293
rect 1353 4287 1367 4300
rect 1393 4287 1407 4300
rect 1353 4047 1367 4053
rect 1216 3887 1223 3993
rect 1236 3983 1243 4003
rect 1336 3987 1343 4034
rect 1376 4036 1383 4113
rect 1413 4040 1427 4053
rect 1436 4047 1443 4173
rect 1416 4036 1423 4040
rect 1456 4027 1463 4293
rect 1476 4203 1483 4473
rect 1516 4367 1523 4473
rect 1536 4427 1543 4513
rect 1576 4336 1583 4453
rect 1507 4303 1520 4307
rect 1507 4296 1523 4303
rect 1507 4293 1520 4296
rect 1553 4287 1567 4293
rect 1527 4273 1533 4287
rect 1476 4196 1503 4203
rect 1476 4047 1483 4133
rect 1496 4087 1503 4196
rect 1516 4107 1523 4213
rect 1596 4207 1603 4253
rect 1616 4163 1623 4513
rect 1636 4303 1643 4413
rect 1736 4367 1743 4523
rect 1756 4347 1763 4513
rect 1796 4507 1803 4772
rect 1976 4767 1983 4813
rect 1996 4787 2003 5253
rect 2036 5207 2043 5343
rect 2136 5047 2143 5253
rect 2156 5207 2163 5343
rect 2193 5327 2207 5333
rect 2236 5327 2243 5473
rect 2296 5376 2303 5433
rect 2276 5307 2283 5343
rect 2173 5287 2187 5293
rect 2186 5280 2187 5287
rect 2196 5167 2203 5273
rect 2233 5123 2247 5133
rect 2196 5120 2247 5123
rect 2193 5116 2243 5120
rect 2193 5107 2207 5116
rect 2253 5088 2267 5093
rect 2167 5083 2180 5087
rect 2167 5076 2183 5083
rect 2167 5073 2180 5076
rect 2276 5047 2283 5293
rect 2036 4867 2043 5013
rect 2056 4927 2063 5043
rect 2096 4967 2103 5043
rect 2116 5007 2123 5033
rect 2076 4868 2083 4893
rect 2096 4887 2103 4913
rect 2116 4867 2123 4913
rect 2016 4787 2023 4853
rect 2056 4820 2063 4823
rect 2053 4807 2067 4820
rect 2136 4807 2143 4933
rect 1876 4687 1883 4753
rect 1816 4556 1843 4563
rect 1896 4556 1903 4753
rect 1636 4296 1663 4303
rect 1696 4300 1703 4303
rect 1656 4227 1663 4296
rect 1693 4287 1707 4300
rect 1733 4286 1747 4292
rect 1676 4247 1683 4273
rect 1607 4156 1623 4163
rect 1596 4127 1603 4153
rect 1633 4107 1647 4113
rect 1516 4093 1533 4107
rect 1516 4063 1523 4093
rect 1620 4086 1640 4087
rect 1496 4056 1523 4063
rect 1496 4036 1503 4056
rect 1533 4040 1547 4053
rect 1556 4047 1563 4076
rect 1627 4073 1633 4086
rect 1587 4053 1593 4067
rect 1536 4036 1543 4040
rect 1696 4036 1703 4153
rect 1396 4000 1403 4003
rect 1236 3976 1263 3983
rect 1236 3867 1243 3913
rect 1256 3887 1263 3976
rect 796 3296 803 3353
rect 836 3296 843 3413
rect 896 3327 903 3514
rect 936 3323 943 3483
rect 1013 3463 1027 3473
rect 996 3460 1027 3463
rect 1036 3463 1043 3514
rect 1056 3483 1063 3593
rect 1076 3527 1083 3653
rect 1156 3483 1163 3573
rect 1176 3527 1183 3733
rect 1216 3707 1223 3733
rect 1276 3707 1283 3783
rect 1256 3567 1263 3613
rect 1276 3607 1283 3693
rect 1296 3647 1303 3873
rect 1316 3687 1323 3953
rect 1336 3947 1343 3973
rect 1356 3923 1363 3993
rect 1393 3987 1407 4000
rect 1456 3967 1463 3992
rect 1336 3916 1363 3923
rect 1336 3727 1343 3916
rect 1516 3907 1523 4003
rect 1576 3987 1583 4013
rect 1587 3883 1600 3887
rect 1587 3880 1603 3883
rect 1587 3873 1607 3880
rect 1593 3867 1607 3873
rect 1536 3816 1543 3853
rect 1316 3623 1323 3673
rect 1296 3616 1323 3623
rect 1253 3520 1267 3532
rect 1256 3516 1263 3520
rect 1056 3476 1083 3483
rect 996 3456 1023 3460
rect 1036 3456 1063 3463
rect 956 3327 963 3353
rect 996 3327 1003 3456
rect 1056 3447 1063 3456
rect 1076 3447 1083 3476
rect 916 3316 943 3323
rect 916 3303 923 3316
rect 896 3296 923 3303
rect 756 3207 763 3294
rect 816 3247 823 3263
rect 676 2956 703 2963
rect 676 2927 683 2956
rect 676 2627 683 2813
rect 696 2707 703 2933
rect 736 2827 743 2963
rect 733 2780 747 2792
rect 736 2776 743 2780
rect 716 2587 723 2743
rect 553 2480 567 2493
rect 556 2476 563 2480
rect 596 2476 603 2513
rect 736 2476 743 2513
rect 576 2440 583 2443
rect 573 2427 587 2440
rect 616 2367 623 2432
rect 656 2387 663 2474
rect 796 2443 803 3193
rect 816 3107 823 3233
rect 896 3063 903 3296
rect 913 3247 927 3253
rect 896 3056 923 3063
rect 896 2927 903 3033
rect 816 2746 823 2813
rect 836 2567 843 2873
rect 916 2867 923 3056
rect 976 3027 983 3253
rect 1016 3047 1023 3393
rect 1036 3307 1043 3433
rect 1056 3296 1063 3433
rect 1096 3367 1103 3483
rect 1136 3476 1163 3483
rect 1096 3296 1103 3353
rect 1136 3347 1143 3476
rect 1036 3007 1043 3253
rect 1116 3207 1123 3263
rect 936 2787 943 2953
rect 956 2827 963 2873
rect 956 2746 963 2813
rect 1016 2807 1023 2963
rect 1056 2927 1063 2994
rect 1036 2776 1043 2833
rect 1076 2827 1083 3013
rect 1136 2996 1143 3173
rect 1156 3107 1163 3393
rect 1176 3307 1183 3473
rect 1196 3447 1203 3483
rect 1256 3387 1263 3433
rect 1226 3333 1227 3340
rect 1213 3327 1227 3333
rect 1236 3296 1243 3333
rect 1276 3307 1283 3473
rect 1176 3167 1183 3253
rect 1216 3207 1223 3263
rect 1296 3263 1303 3616
rect 1336 3567 1343 3613
rect 1376 3587 1383 3772
rect 1407 3756 1433 3763
rect 1516 3707 1523 3783
rect 1556 3780 1563 3783
rect 1553 3767 1567 3780
rect 1407 3534 1413 3547
rect 1400 3533 1420 3534
rect 1316 3427 1323 3533
rect 1336 3383 1343 3473
rect 1356 3427 1363 3483
rect 1396 3447 1403 3483
rect 1336 3376 1353 3383
rect 1327 3313 1333 3327
rect 1356 3296 1363 3373
rect 1436 3347 1443 3473
rect 1456 3447 1463 3653
rect 1476 3327 1483 3593
rect 1496 3547 1503 3573
rect 1516 3547 1523 3672
rect 1493 3520 1507 3533
rect 1556 3523 1563 3713
rect 1576 3607 1583 3693
rect 1596 3667 1603 3733
rect 1496 3516 1503 3520
rect 1556 3516 1583 3523
rect 1576 3487 1583 3516
rect 1596 3487 1603 3593
rect 1616 3567 1623 4013
rect 1676 3947 1683 4003
rect 1716 3983 1723 4213
rect 1736 4007 1743 4233
rect 1756 4048 1763 4293
rect 1776 4187 1783 4413
rect 1796 4383 1803 4472
rect 1816 4407 1823 4556
rect 1796 4376 1823 4383
rect 1816 4336 1823 4376
rect 1836 4367 1843 4493
rect 1876 4427 1883 4523
rect 1896 4347 1903 4493
rect 1916 4427 1923 4713
rect 1936 4547 1943 4633
rect 1796 4227 1803 4273
rect 1816 4207 1823 4273
rect 1836 4247 1843 4303
rect 1776 4127 1783 4152
rect 1796 4067 1803 4113
rect 1796 4036 1803 4053
rect 1836 4036 1843 4093
rect 1856 4087 1863 4273
rect 1876 4227 1883 4303
rect 1916 4303 1923 4353
rect 1936 4347 1943 4533
rect 1956 4507 1963 4693
rect 1996 4556 2003 4733
rect 2036 4627 2043 4653
rect 1956 4336 1963 4453
rect 1996 4336 2003 4453
rect 2016 4387 2023 4473
rect 2056 4343 2063 4413
rect 2076 4367 2083 4613
rect 2096 4607 2103 4653
rect 2127 4613 2133 4627
rect 2116 4563 2123 4592
rect 2156 4587 2163 5033
rect 2196 4907 2203 5032
rect 2253 5027 2267 5033
rect 2216 4856 2223 4993
rect 2276 4983 2283 5012
rect 2236 4976 2283 4983
rect 2236 4947 2243 4976
rect 2256 4856 2263 4933
rect 2196 4787 2203 4823
rect 2236 4807 2243 4823
rect 2247 4796 2263 4803
rect 2107 4556 2123 4563
rect 2133 4560 2147 4573
rect 2136 4556 2143 4560
rect 2096 4427 2103 4554
rect 2116 4407 2123 4513
rect 2196 4520 2203 4523
rect 2193 4507 2207 4520
rect 2176 4496 2193 4503
rect 2136 4407 2143 4473
rect 2056 4336 2083 4343
rect 2116 4336 2123 4393
rect 2176 4367 2183 4496
rect 2216 4487 2223 4513
rect 2236 4483 2243 4573
rect 2256 4567 2263 4796
rect 2296 4727 2303 5313
rect 2316 5267 2323 5343
rect 2356 5287 2363 5533
rect 2376 5527 2383 5563
rect 2416 5487 2423 5913
rect 2476 5896 2483 5953
rect 2456 5827 2463 5863
rect 2496 5847 2503 5863
rect 2476 5836 2493 5843
rect 2436 5687 2443 5713
rect 2456 5707 2463 5813
rect 2436 5447 2443 5652
rect 2476 5608 2483 5836
rect 2536 5707 2543 5993
rect 2636 5896 2643 5993
rect 2556 5847 2563 5894
rect 2616 5847 2623 5863
rect 2616 5836 2633 5847
rect 2620 5833 2633 5836
rect 2676 5827 2683 5953
rect 2776 5896 2783 5953
rect 2796 5947 2803 6112
rect 2856 6080 2863 6083
rect 2896 6080 2903 6083
rect 2853 6067 2867 6080
rect 2893 6067 2907 6080
rect 2696 5847 2703 5894
rect 2756 5860 2763 5863
rect 2753 5847 2767 5860
rect 2736 5767 2743 5833
rect 2796 5827 2803 5863
rect 2656 5596 2663 5693
rect 2536 5560 2543 5563
rect 2533 5547 2547 5560
rect 2456 5427 2463 5533
rect 2476 5376 2483 5453
rect 2316 5107 2323 5213
rect 2336 5127 2343 5193
rect 2356 5103 2363 5233
rect 2376 5187 2383 5374
rect 2456 5340 2463 5343
rect 2453 5327 2467 5340
rect 2516 5267 2523 5473
rect 2576 5427 2583 5594
rect 2716 5566 2723 5713
rect 2636 5547 2643 5563
rect 2636 5376 2643 5533
rect 2676 5527 2683 5552
rect 2616 5340 2623 5343
rect 2396 5107 2403 5193
rect 2416 5167 2423 5213
rect 2336 5096 2363 5103
rect 2336 5076 2343 5096
rect 2373 5080 2387 5093
rect 2376 5076 2383 5080
rect 2356 5040 2363 5043
rect 2316 4887 2323 5033
rect 2353 5027 2367 5040
rect 2366 5020 2367 5027
rect 2336 4856 2343 4893
rect 2376 4868 2383 5013
rect 2396 4987 2403 5043
rect 2396 4947 2403 4973
rect 2416 4867 2423 4993
rect 2316 4767 2323 4813
rect 2356 4787 2363 4823
rect 2316 4707 2323 4732
rect 2296 4588 2303 4692
rect 2340 4563 2353 4567
rect 2336 4556 2353 4563
rect 2340 4553 2353 4556
rect 2293 4487 2307 4493
rect 2236 4476 2263 4483
rect 1916 4296 1943 4303
rect 1876 4047 1883 4153
rect 1716 3976 1743 3983
rect 1667 3933 1683 3947
rect 1676 3927 1683 3933
rect 1676 3816 1683 3853
rect 1656 3763 1663 3783
rect 1656 3756 1683 3763
rect 1636 3607 1643 3653
rect 1676 3643 1683 3756
rect 1696 3667 1703 3783
rect 1736 3747 1743 3976
rect 1756 3827 1763 4034
rect 1767 3823 1780 3827
rect 1767 3816 1783 3823
rect 1767 3813 1780 3816
rect 1793 3766 1807 3772
rect 1736 3643 1743 3673
rect 1676 3636 1743 3643
rect 1673 3587 1687 3593
rect 1673 3580 1693 3587
rect 1676 3576 1693 3580
rect 1680 3573 1693 3576
rect 1387 3313 1393 3327
rect 1440 3326 1460 3327
rect 1447 3313 1453 3326
rect 1496 3303 1503 3413
rect 1516 3387 1523 3433
rect 1536 3303 1543 3472
rect 1616 3467 1623 3553
rect 1653 3520 1667 3533
rect 1693 3520 1707 3533
rect 1656 3516 1663 3520
rect 1696 3516 1703 3520
rect 1476 3296 1503 3303
rect 1516 3296 1543 3303
rect 1556 3296 1563 3333
rect 1276 3256 1303 3263
rect 1176 3008 1183 3113
rect 1096 2907 1103 2953
rect 1096 2787 1103 2893
rect 1116 2887 1123 2963
rect 856 2507 863 2693
rect 976 2647 983 2773
rect 1056 2740 1063 2743
rect 1053 2727 1067 2740
rect 876 2476 883 2513
rect 936 2447 943 2633
rect 976 2487 983 2633
rect 1096 2587 1103 2733
rect 1116 2563 1123 2813
rect 1136 2783 1143 2933
rect 1156 2867 1163 2963
rect 1136 2776 1153 2783
rect 1196 2776 1203 2952
rect 1236 2808 1243 3153
rect 1276 3027 1283 3256
rect 1296 2996 1303 3153
rect 1356 3147 1363 3173
rect 1347 3123 1360 3127
rect 1347 3120 1363 3123
rect 1347 3113 1367 3120
rect 1353 3107 1367 3113
rect 1276 2960 1283 2963
rect 1273 2947 1287 2960
rect 1316 2867 1323 2963
rect 1376 2947 1383 3253
rect 1456 3207 1463 3263
rect 1516 3167 1523 3296
rect 1636 3307 1643 3473
rect 1396 2927 1403 3153
rect 1436 2996 1443 3033
rect 1516 2967 1523 3132
rect 1536 3067 1543 3253
rect 1656 3263 1663 3453
rect 1676 3427 1683 3483
rect 1736 3467 1743 3636
rect 1696 3307 1703 3453
rect 1756 3443 1763 3759
rect 1776 3587 1783 3613
rect 1836 3548 1843 3973
rect 1896 3967 1903 4293
rect 1856 3687 1863 3953
rect 1916 3867 1923 4193
rect 1936 3987 1943 4296
rect 1976 4267 1983 4292
rect 2016 4283 2023 4303
rect 2016 4276 2043 4283
rect 2036 4247 2043 4276
rect 2036 4187 2043 4233
rect 2056 4207 2063 4313
rect 1956 4036 1963 4073
rect 2016 4048 2023 4113
rect 1913 3820 1927 3832
rect 1916 3816 1923 3820
rect 1976 3823 1983 3913
rect 1996 3887 2003 4003
rect 2016 3847 2023 3973
rect 2036 3967 2043 4173
rect 2076 4167 2083 4336
rect 2196 4347 2203 4393
rect 2136 4247 2143 4303
rect 2096 4147 2103 4213
rect 2056 3927 2063 4073
rect 2136 4036 2143 4212
rect 2116 3967 2123 4003
rect 2176 3887 2183 4113
rect 2196 3947 2203 4293
rect 2216 4127 2223 4413
rect 2236 4347 2243 4453
rect 2256 4347 2263 4476
rect 2356 4467 2363 4513
rect 2376 4503 2383 4793
rect 2396 4527 2403 4753
rect 2436 4588 2443 5253
rect 2576 5247 2583 5332
rect 2613 5327 2627 5340
rect 2496 5107 2503 5133
rect 2516 5076 2523 5232
rect 2656 5076 2663 5113
rect 2676 5107 2683 5433
rect 2736 5376 2743 5753
rect 2756 5596 2763 5793
rect 2856 5727 2863 6053
rect 2936 5967 2943 6233
rect 3716 6227 3723 6303
rect 3816 6296 3843 6303
rect 2956 6007 2963 6193
rect 3056 6116 3063 6193
rect 2996 6047 3003 6083
rect 2956 5947 2963 5993
rect 2896 5908 2903 5933
rect 3036 5908 3043 6083
rect 3096 6067 3103 6153
rect 3173 6147 3187 6153
rect 3196 6116 3203 6213
rect 3227 6173 3233 6187
rect 3267 6173 3273 6187
rect 3296 6160 3333 6163
rect 3293 6156 3333 6160
rect 3176 6080 3183 6083
rect 3173 6067 3187 6080
rect 2916 5807 2923 5863
rect 2956 5623 2963 5893
rect 3016 5667 3023 5852
rect 3096 5827 3103 6032
rect 3236 5987 3243 6152
rect 3293 6148 3307 6156
rect 3256 5967 3263 6113
rect 3316 6080 3323 6083
rect 3116 5863 3123 5933
rect 3216 5896 3263 5903
rect 3116 5856 3143 5863
rect 2956 5616 2983 5623
rect 2816 5596 2843 5603
rect 2776 5387 2783 5563
rect 2836 5543 2843 5596
rect 2976 5596 2983 5616
rect 3116 5596 3123 5793
rect 3136 5687 3143 5856
rect 3196 5807 3203 5863
rect 3156 5596 3163 5713
rect 3173 5627 3187 5633
rect 3196 5607 3203 5693
rect 3256 5647 3263 5896
rect 3276 5767 3283 6073
rect 3313 6067 3327 6080
rect 3293 6043 3307 6053
rect 3293 6040 3343 6043
rect 3296 6036 3343 6040
rect 3316 5928 3323 6013
rect 3336 6007 3343 6036
rect 3376 6027 3383 6153
rect 3396 6128 3403 6173
rect 3416 6127 3423 6213
rect 3476 6128 3483 6153
rect 3396 6087 3403 6114
rect 3306 5896 3324 5904
rect 3356 5896 3363 5973
rect 3416 5863 3423 6073
rect 3456 5947 3463 6083
rect 3516 6027 3523 6173
rect 3613 6120 3627 6133
rect 3616 6116 3623 6120
rect 3716 6116 3723 6153
rect 3816 6127 3823 6296
rect 5756 6247 5763 6303
rect 5916 6296 5943 6303
rect 3556 6007 3563 6083
rect 3596 6080 3603 6083
rect 3593 6067 3607 6080
rect 3636 6047 3643 6073
rect 3736 6047 3743 6072
rect 3796 6047 3803 6114
rect 3876 6116 3923 6123
rect 3816 5987 3823 6073
rect 3916 6083 3923 6116
rect 3896 6076 3923 6083
rect 3936 6116 3963 6123
rect 3896 6067 3903 6076
rect 3556 5867 3563 5972
rect 3540 5866 3553 5867
rect 3416 5856 3443 5863
rect 3456 5860 3463 5863
rect 3347 5813 3353 5827
rect 3216 5566 3223 5633
rect 3253 5600 3267 5612
rect 3336 5608 3343 5653
rect 3256 5596 3263 5600
rect 3356 5587 3363 5693
rect 3376 5647 3383 5852
rect 3416 5687 3423 5833
rect 3436 5807 3443 5856
rect 3453 5847 3467 5860
rect 3547 5853 3553 5866
rect 3453 5827 3467 5833
rect 3476 5767 3483 5813
rect 3436 5687 3443 5753
rect 3456 5596 3463 5713
rect 3576 5687 3583 5973
rect 3636 5896 3643 5973
rect 3667 5916 3693 5923
rect 3596 5727 3603 5853
rect 3613 5846 3627 5852
rect 3547 5683 3560 5687
rect 3547 5680 3563 5683
rect 3547 5673 3567 5680
rect 3553 5667 3567 5673
rect 3636 5627 3643 5653
rect 3573 5600 3587 5613
rect 3576 5596 3583 5600
rect 2816 5536 2843 5543
rect 2816 5387 2823 5536
rect 2896 5376 2903 5473
rect 2956 5423 2963 5563
rect 2936 5416 2963 5423
rect 2913 5388 2927 5393
rect 2716 5123 2723 5332
rect 2716 5116 2743 5123
rect 2700 5083 2713 5087
rect 2696 5076 2713 5083
rect 2536 5040 2543 5043
rect 2533 5027 2547 5040
rect 2596 5007 2603 5074
rect 2700 5073 2713 5076
rect 2476 4856 2483 4973
rect 2636 4967 2643 5043
rect 2596 4867 2603 4893
rect 2456 4587 2463 4773
rect 2496 4747 2503 4823
rect 2536 4820 2543 4823
rect 2533 4807 2547 4820
rect 2576 4747 2583 4854
rect 2676 4856 2683 4993
rect 2473 4560 2487 4573
rect 2516 4567 2523 4613
rect 2476 4556 2483 4560
rect 2376 4496 2393 4503
rect 2347 4436 2383 4443
rect 2356 4343 2363 4413
rect 2376 4367 2383 4436
rect 2396 4427 2403 4492
rect 2456 4487 2463 4523
rect 2513 4467 2527 4473
rect 2536 4467 2543 4713
rect 2596 4587 2603 4813
rect 2616 4767 2623 4812
rect 2656 4807 2663 4823
rect 2716 4807 2723 4953
rect 2736 4867 2743 5116
rect 2756 4907 2763 5113
rect 2816 5107 2823 5332
rect 2836 5323 2843 5343
rect 2836 5316 2863 5323
rect 2787 5076 2803 5083
rect 2856 5076 2863 5316
rect 2776 5007 2783 5073
rect 2836 4987 2843 5043
rect 2876 5007 2883 5153
rect 2816 4887 2823 4953
rect 2756 4843 2763 4872
rect 2813 4860 2827 4873
rect 2816 4856 2823 4860
rect 2736 4836 2763 4843
rect 2653 4787 2667 4793
rect 2646 4773 2647 4780
rect 2633 4763 2647 4773
rect 2633 4760 2663 4763
rect 2636 4756 2663 4760
rect 2556 4507 2563 4573
rect 2616 4556 2623 4732
rect 2636 4667 2643 4733
rect 2656 4627 2663 4756
rect 2696 4647 2703 4693
rect 2716 4627 2723 4772
rect 2736 4687 2743 4836
rect 2756 4816 2773 4823
rect 2756 4787 2763 4816
rect 2856 4823 2863 4933
rect 2836 4816 2863 4823
rect 2876 4787 2883 4972
rect 2896 4747 2903 5193
rect 2916 4887 2923 5332
rect 2936 5087 2943 5416
rect 2956 5367 2963 5393
rect 2987 5383 3000 5387
rect 2987 5376 3003 5383
rect 2987 5374 3000 5376
rect 3096 5347 3103 5413
rect 3176 5376 3183 5413
rect 3216 5376 3223 5493
rect 3276 5383 3283 5563
rect 3256 5376 3283 5383
rect 3313 5380 3327 5393
rect 3316 5376 3323 5380
rect 3056 5287 3063 5343
rect 3116 5167 3123 5374
rect 3156 5287 3163 5343
rect 3196 5267 3203 5332
rect 2993 5127 3007 5133
rect 3076 5120 3113 5123
rect 3073 5116 3113 5120
rect 2973 5080 2987 5093
rect 2976 5076 2983 5080
rect 2996 4927 3003 5043
rect 2656 4527 2663 4573
rect 2716 4556 2723 4592
rect 2796 4568 2803 4713
rect 2856 4607 2863 4733
rect 2896 4627 2903 4693
rect 2880 4563 2893 4567
rect 2876 4556 2893 4563
rect 2593 4507 2607 4513
rect 2336 4336 2363 4343
rect 2236 4306 2243 4333
rect 2256 4063 2263 4293
rect 2316 4187 2323 4303
rect 2316 4107 2323 4173
rect 2376 4147 2383 4332
rect 2476 4303 2483 4453
rect 2496 4307 2503 4413
rect 2516 4348 2523 4413
rect 2556 4387 2563 4493
rect 2576 4407 2583 4473
rect 2696 4447 2703 4473
rect 2596 4363 2603 4413
rect 2616 4407 2623 4433
rect 2647 4404 2660 4407
rect 2647 4400 2663 4404
rect 2647 4393 2667 4400
rect 2653 4387 2667 4393
rect 2716 4387 2723 4453
rect 2776 4427 2783 4513
rect 2596 4356 2623 4363
rect 2396 4147 2403 4293
rect 2416 4267 2423 4303
rect 2456 4296 2483 4303
rect 2256 4056 2283 4063
rect 1976 3816 2003 3823
rect 1936 3780 1943 3783
rect 1933 3767 1947 3780
rect 1876 3687 1883 3713
rect 1936 3567 1943 3753
rect 1956 3548 1963 3633
rect 1996 3567 2003 3816
rect 2016 3787 2023 3812
rect 2096 3780 2103 3783
rect 2093 3767 2107 3780
rect 1773 3527 1787 3533
rect 1796 3536 1833 3543
rect 1796 3516 1803 3536
rect 1876 3487 1883 3533
rect 1913 3520 1927 3533
rect 1916 3516 1923 3520
rect 1776 3447 1783 3473
rect 1893 3467 1907 3473
rect 1736 3436 1763 3443
rect 1616 3227 1623 3263
rect 1636 3256 1663 3263
rect 1576 3047 1583 3173
rect 1456 2907 1463 2963
rect 1536 2927 1543 3013
rect 1576 2996 1583 3033
rect 1636 3027 1643 3256
rect 1626 3013 1627 3020
rect 1613 3000 1627 3013
rect 1656 3007 1663 3093
rect 1616 2996 1623 3000
rect 1136 2567 1143 2733
rect 1176 2687 1183 2743
rect 1216 2707 1223 2743
rect 1096 2556 1123 2563
rect 556 2256 563 2313
rect 696 2256 703 2313
rect 736 2287 743 2413
rect 756 2407 763 2443
rect 776 2436 803 2443
rect 740 2263 753 2267
rect 736 2256 753 2263
rect 740 2254 753 2256
rect 740 2253 744 2254
rect 536 2127 543 2223
rect 576 2220 583 2223
rect 573 2207 587 2220
rect 393 1960 407 1972
rect 396 1956 403 1960
rect 436 1956 443 2013
rect 496 1927 503 1973
rect 396 1736 403 1893
rect 416 1847 423 1923
rect 516 1907 523 1993
rect 536 1967 543 2013
rect 573 1960 587 1973
rect 576 1956 583 1960
rect 636 1963 643 2253
rect 673 2206 687 2212
rect 716 2127 723 2212
rect 756 2067 763 2213
rect 776 2087 783 2436
rect 836 2256 843 2293
rect 856 2287 863 2443
rect 816 2220 823 2223
rect 813 2207 827 2220
rect 876 2167 883 2293
rect 636 1956 663 1963
rect 556 1920 563 1923
rect 436 1736 443 1773
rect 336 1696 363 1703
rect 376 1700 383 1703
rect 316 1676 333 1683
rect 273 1440 287 1453
rect 336 1448 343 1673
rect 276 1436 283 1440
rect 356 1447 363 1696
rect 373 1687 387 1700
rect 476 1627 483 1813
rect 536 1787 543 1913
rect 553 1907 567 1920
rect 596 1827 603 1923
rect 656 1907 663 1956
rect 676 1926 683 2053
rect 856 2047 863 2113
rect 736 1956 743 1993
rect 896 1987 903 2293
rect 936 2256 943 2412
rect 956 2407 963 2474
rect 996 2167 1003 2443
rect 867 1983 880 1987
rect 867 1973 883 1983
rect 773 1960 787 1973
rect 776 1956 783 1960
rect 336 1407 343 1434
rect 396 1436 403 1513
rect 436 1436 443 1473
rect 256 1367 263 1403
rect 276 1343 283 1373
rect 176 1336 203 1343
rect 256 1336 283 1343
rect 56 1186 63 1233
rect 116 1216 123 1253
rect 156 1216 163 1273
rect 176 1227 183 1336
rect 96 928 103 1172
rect 136 1147 143 1183
rect 147 1136 163 1143
rect 133 920 147 933
rect 156 927 163 1136
rect 136 916 143 920
rect 36 827 43 913
rect 116 880 123 883
rect 76 703 83 872
rect 113 867 127 880
rect 153 867 167 873
rect 176 867 183 1173
rect 196 947 203 1253
rect 216 1227 223 1273
rect 236 1247 243 1313
rect 256 1216 263 1336
rect 296 1307 303 1403
rect 313 1387 327 1393
rect 476 1347 483 1533
rect 496 1406 503 1553
rect 536 1467 543 1703
rect 576 1527 583 1703
rect 596 1567 603 1693
rect 553 1440 567 1453
rect 556 1436 563 1440
rect 596 1436 603 1553
rect 616 1447 623 1773
rect 696 1736 703 1813
rect 716 1807 723 1923
rect 676 1700 683 1703
rect 716 1700 723 1703
rect 673 1687 687 1700
rect 713 1687 727 1700
rect 536 1383 543 1403
rect 536 1376 563 1383
rect 287 1256 323 1263
rect 293 1220 307 1233
rect 316 1227 323 1256
rect 356 1247 363 1333
rect 296 1216 303 1220
rect 416 1216 423 1253
rect 236 947 243 1183
rect 396 1180 403 1183
rect 196 923 203 933
rect 196 916 223 923
rect 166 860 167 867
rect 156 787 163 853
rect 56 696 103 703
rect 16 188 23 453
rect 56 408 63 696
rect 216 696 223 853
rect 236 827 243 883
rect 276 727 283 883
rect 316 747 323 1173
rect 393 1167 407 1180
rect 476 1167 483 1273
rect 496 1187 503 1293
rect 556 1267 563 1376
rect 576 1367 583 1403
rect 556 1243 563 1253
rect 556 1236 583 1243
rect 576 1216 583 1236
rect 616 1227 623 1393
rect 636 1367 643 1513
rect 656 1407 663 1653
rect 676 1487 683 1613
rect 756 1547 763 1873
rect 816 1767 823 1953
rect 836 1887 843 1973
rect 876 1956 883 1973
rect 936 1947 943 2073
rect 1016 1987 1023 2373
rect 1076 2347 1083 2433
rect 1096 2387 1103 2556
rect 1116 2407 1123 2533
rect 1156 2476 1163 2513
rect 1176 2507 1183 2633
rect 1136 2287 1143 2373
rect 1176 2347 1183 2443
rect 1196 2323 1203 2433
rect 1176 2316 1203 2323
rect 1176 2287 1183 2316
rect 1216 2283 1223 2513
rect 1236 2487 1243 2533
rect 1256 2527 1263 2733
rect 1276 2687 1283 2793
rect 1336 2776 1343 2873
rect 1376 2787 1383 2853
rect 1316 2723 1323 2743
rect 1356 2727 1363 2743
rect 1316 2716 1343 2723
rect 1336 2687 1343 2716
rect 1276 2647 1283 2673
rect 1253 2480 1267 2492
rect 1256 2476 1263 2480
rect 1276 2307 1283 2443
rect 1196 2276 1223 2283
rect 996 1920 1003 1923
rect 893 1907 907 1912
rect 993 1907 1007 1920
rect 693 1448 707 1453
rect 733 1440 747 1453
rect 776 1443 783 1753
rect 836 1736 843 1813
rect 867 1763 880 1767
rect 867 1753 883 1763
rect 876 1736 883 1753
rect 816 1687 823 1703
rect 853 1687 867 1693
rect 827 1676 843 1683
rect 836 1663 843 1676
rect 836 1656 873 1663
rect 736 1436 743 1440
rect 776 1436 803 1443
rect 796 1406 803 1436
rect 396 916 403 953
rect 336 887 343 914
rect 156 427 163 693
rect 136 416 153 423
rect 136 396 143 416
rect 233 400 247 413
rect 276 408 283 663
rect 236 396 243 400
rect 316 403 323 712
rect 336 666 343 873
rect 476 847 483 914
rect 436 696 443 733
rect 316 396 343 403
rect 56 366 63 394
rect 116 360 123 363
rect 113 347 127 360
rect 156 356 183 363
rect 16 107 23 174
rect 156 147 163 333
rect 176 247 183 356
rect 196 347 203 394
rect 336 366 343 396
rect 436 396 443 453
rect 476 408 483 693
rect 496 666 503 1133
rect 553 920 567 933
rect 556 916 563 920
rect 596 916 603 1013
rect 576 880 583 883
rect 516 723 523 753
rect 536 747 543 872
rect 573 867 587 880
rect 636 867 643 1233
rect 656 1227 663 1273
rect 693 1220 707 1233
rect 696 1216 703 1220
rect 736 1216 743 1353
rect 816 1267 823 1473
rect 876 1467 883 1553
rect 916 1527 923 1733
rect 936 1627 943 1893
rect 996 1767 1003 1893
rect 1036 1823 1043 1953
rect 1056 1827 1063 1993
rect 1096 1956 1103 1993
rect 1156 1983 1163 2273
rect 1196 2263 1203 2276
rect 1267 2283 1280 2287
rect 1267 2273 1283 2283
rect 1136 1976 1163 1983
rect 1176 2256 1203 2263
rect 1136 1968 1143 1976
rect 1176 1963 1183 2256
rect 1276 2256 1283 2273
rect 1296 2267 1303 2393
rect 1316 2387 1323 2433
rect 1336 2423 1343 2673
rect 1356 2507 1363 2713
rect 1376 2547 1383 2733
rect 1396 2727 1403 2813
rect 1436 2787 1443 2833
rect 1516 2803 1523 2913
rect 1516 2800 1543 2803
rect 1516 2796 1547 2800
rect 1493 2780 1507 2793
rect 1533 2787 1547 2796
rect 1496 2776 1503 2780
rect 1520 2743 1533 2747
rect 1476 2740 1483 2743
rect 1473 2727 1487 2740
rect 1516 2736 1533 2743
rect 1520 2733 1533 2736
rect 1473 2687 1487 2692
rect 1516 2687 1523 2713
rect 1556 2707 1563 2933
rect 1576 2727 1583 2913
rect 1616 2787 1623 2933
rect 1636 2867 1643 2963
rect 1607 2776 1623 2787
rect 1607 2773 1620 2776
rect 1416 2507 1423 2553
rect 1436 2488 1443 2573
rect 1356 2447 1363 2472
rect 1336 2416 1363 2423
rect 1196 2147 1203 2193
rect 1176 1956 1203 1963
rect 1156 1920 1163 1923
rect 1153 1907 1167 1920
rect 1016 1816 1043 1823
rect 1016 1787 1023 1816
rect 1016 1743 1023 1773
rect 996 1736 1023 1743
rect 976 1667 983 1703
rect 1036 1627 1043 1793
rect 1056 1706 1063 1753
rect 1156 1736 1163 1773
rect 1136 1700 1143 1703
rect 1133 1687 1147 1700
rect 876 1436 883 1453
rect 913 1440 927 1453
rect 916 1436 923 1440
rect 956 1407 963 1453
rect 896 1287 903 1403
rect 676 1147 683 1183
rect 776 1067 783 1253
rect 836 1216 843 1253
rect 916 1216 923 1353
rect 976 1347 983 1613
rect 1196 1443 1203 1956
rect 1216 1887 1223 2173
rect 1316 2167 1323 2293
rect 1336 2207 1343 2393
rect 1356 2347 1363 2416
rect 1416 2387 1423 2443
rect 1456 2436 1473 2443
rect 1396 2268 1403 2293
rect 1440 2263 1453 2267
rect 1436 2256 1453 2263
rect 1440 2254 1453 2256
rect 1476 2227 1483 2433
rect 1496 2407 1503 2573
rect 1596 2443 1603 2513
rect 1616 2487 1623 2613
rect 1636 2587 1643 2743
rect 1676 2587 1683 3294
rect 1716 3296 1723 3433
rect 1736 3327 1743 3436
rect 1756 3347 1763 3413
rect 1796 3387 1803 3453
rect 1936 3463 1943 3483
rect 1916 3456 1943 3463
rect 1776 3323 1783 3353
rect 1756 3316 1783 3323
rect 1756 3296 1763 3316
rect 1693 3243 1707 3253
rect 1693 3240 1723 3243
rect 1696 3236 1723 3240
rect 1716 3087 1723 3236
rect 1736 3127 1743 3252
rect 1776 3227 1783 3263
rect 1707 3066 1720 3067
rect 1707 3053 1713 3066
rect 1696 2927 1703 3013
rect 1716 3008 1723 3032
rect 1736 3023 1743 3053
rect 1756 3023 1763 3153
rect 1796 3043 1803 3253
rect 1876 3147 1883 3452
rect 1896 3187 1903 3432
rect 1916 3307 1923 3456
rect 1976 3447 1983 3483
rect 1936 3387 1943 3433
rect 2016 3367 2023 3752
rect 2036 3607 2043 3693
rect 2056 3587 2063 3613
rect 2116 3547 2123 3772
rect 2136 3707 2143 3853
rect 2216 3848 2223 4003
rect 2236 3847 2243 3913
rect 2256 3827 2263 3973
rect 2276 3827 2283 4056
rect 2316 3987 2323 4093
rect 2456 4087 2463 4296
rect 2596 4287 2603 4334
rect 2616 4327 2623 4356
rect 2476 4036 2483 4093
rect 2496 4067 2503 4233
rect 2516 4036 2523 4273
rect 2636 4267 2643 4372
rect 2656 4287 2663 4303
rect 2536 4087 2543 4173
rect 2596 4007 2603 4252
rect 2656 4227 2663 4273
rect 2716 4227 2723 4303
rect 2736 4247 2743 4334
rect 2616 4047 2623 4173
rect 2656 4063 2663 4213
rect 2636 4056 2663 4063
rect 2636 4036 2643 4056
rect 2676 4036 2683 4113
rect 2716 4047 2723 4133
rect 2356 4000 2363 4003
rect 2353 3987 2367 4000
rect 2156 3747 2163 3772
rect 2156 3703 2163 3733
rect 2176 3727 2183 3753
rect 2156 3696 2183 3703
rect 2113 3520 2127 3533
rect 2136 3527 2143 3553
rect 2116 3516 2123 3520
rect 2016 3307 2023 3332
rect 1996 3227 2003 3263
rect 2036 3187 2043 3513
rect 2096 3476 2135 3484
rect 2056 3447 2063 3473
rect 2107 3453 2113 3467
rect 2076 3347 2083 3393
rect 2096 3307 2103 3432
rect 2156 3407 2163 3553
rect 2176 3447 2183 3696
rect 2256 3528 2263 3773
rect 2276 3563 2283 3792
rect 2296 3747 2303 3933
rect 2316 3827 2323 3952
rect 2336 3927 2343 3973
rect 2396 3967 2403 4003
rect 2496 3987 2503 4003
rect 2496 3973 2513 3987
rect 2400 3943 2413 3947
rect 2396 3933 2413 3943
rect 2396 3847 2403 3933
rect 2496 3907 2503 3973
rect 2576 3947 2583 3993
rect 2413 3820 2427 3833
rect 2416 3816 2423 3820
rect 2336 3647 2343 3783
rect 2276 3556 2303 3563
rect 2296 3527 2303 3556
rect 2356 3547 2363 3653
rect 2376 3567 2383 3772
rect 2416 3667 2423 3753
rect 2476 3687 2483 3813
rect 2116 3296 2123 3373
rect 2153 3300 2167 3313
rect 2196 3307 2203 3473
rect 2236 3367 2243 3483
rect 2276 3427 2283 3483
rect 2296 3363 2303 3473
rect 2316 3427 2323 3533
rect 2353 3520 2367 3533
rect 2356 3516 2363 3520
rect 2413 3467 2427 3473
rect 2436 3427 2443 3514
rect 2276 3356 2303 3363
rect 2156 3296 2163 3300
rect 1796 3036 1823 3043
rect 1736 3016 1763 3023
rect 1736 2996 1743 3016
rect 1756 2960 1763 2963
rect 1713 2947 1727 2953
rect 1753 2947 1767 2960
rect 1816 2947 1823 3036
rect 1776 2847 1783 2933
rect 1796 2827 1803 2913
rect 1836 2887 1843 3113
rect 1856 3008 1863 3073
rect 1916 2996 1923 3033
rect 1896 2927 1903 2963
rect 1753 2807 1767 2813
rect 1753 2800 1773 2807
rect 1756 2796 1773 2800
rect 1760 2794 1773 2796
rect 1816 2783 1823 2853
rect 1896 2808 1903 2913
rect 1796 2776 1823 2783
rect 1936 2776 1943 3053
rect 1956 2867 1963 3073
rect 1976 3007 1983 3133
rect 1996 2996 2003 3153
rect 2056 3087 2063 3293
rect 2036 2996 2043 3033
rect 2076 2987 2083 3293
rect 2116 3008 2123 3133
rect 2176 3107 2183 3263
rect 2176 2996 2183 3072
rect 1976 2927 1983 2953
rect 1956 2787 1963 2853
rect 1976 2788 1983 2813
rect 1696 2583 1703 2753
rect 1716 2707 1723 2732
rect 1716 2647 1723 2693
rect 1736 2627 1743 2743
rect 1756 2647 1763 2713
rect 1836 2687 1843 2753
rect 1876 2723 1883 2743
rect 1876 2716 1903 2723
rect 1696 2576 1723 2583
rect 1653 2480 1667 2493
rect 1656 2476 1663 2480
rect 1696 2476 1703 2553
rect 1716 2527 1723 2576
rect 1756 2487 1763 2593
rect 1556 2436 1603 2443
rect 1636 2440 1643 2443
rect 1633 2427 1647 2440
rect 1516 2267 1523 2413
rect 1676 2407 1683 2443
rect 1713 2427 1727 2433
rect 1736 2367 1743 2473
rect 1576 2256 1583 2293
rect 1716 2267 1723 2333
rect 1756 2327 1763 2433
rect 1776 2387 1783 2443
rect 1836 2387 1843 2573
rect 1896 2547 1903 2716
rect 1916 2687 1923 2743
rect 1953 2723 1967 2733
rect 1953 2720 1983 2723
rect 1956 2716 1987 2720
rect 1973 2707 1987 2716
rect 1916 2647 1923 2673
rect 1936 2627 1943 2653
rect 1776 2307 1783 2373
rect 1856 2347 1863 2513
rect 1896 2488 1903 2533
rect 1936 2476 1943 2613
rect 1956 2527 1963 2693
rect 1916 2440 1923 2443
rect 1876 2403 1883 2433
rect 1913 2427 1927 2440
rect 1876 2396 1903 2403
rect 1276 1988 1283 2133
rect 1336 1963 1343 2153
rect 1356 2087 1363 2213
rect 1376 2103 1383 2212
rect 1396 2123 1403 2193
rect 1416 2147 1423 2212
rect 1396 2116 1443 2123
rect 1376 2096 1413 2103
rect 1316 1956 1343 1963
rect 1256 1767 1263 1923
rect 1296 1887 1303 1923
rect 1336 1847 1343 1913
rect 1216 1567 1223 1753
rect 1276 1736 1283 1813
rect 1256 1700 1263 1703
rect 1253 1687 1267 1700
rect 1196 1436 1223 1443
rect 876 1167 883 1213
rect 1016 1183 1023 1213
rect 976 1176 1023 1183
rect 1036 1183 1043 1333
rect 1076 1267 1083 1434
rect 1176 1327 1183 1403
rect 1096 1243 1103 1313
rect 1216 1287 1223 1436
rect 1236 1367 1243 1413
rect 1276 1367 1283 1403
rect 1076 1236 1103 1243
rect 1076 1228 1083 1236
rect 1036 1176 1063 1183
rect 676 916 683 1013
rect 713 928 727 933
rect 776 887 783 953
rect 696 880 703 883
rect 693 867 707 880
rect 916 886 923 973
rect 976 947 983 1153
rect 976 916 983 933
rect 1016 916 1023 973
rect 736 787 743 872
rect 516 716 543 723
rect 536 696 543 716
rect 636 663 643 773
rect 596 656 643 663
rect 656 663 663 733
rect 713 700 727 713
rect 716 696 723 700
rect 756 696 763 733
rect 776 707 783 833
rect 956 827 963 883
rect 996 880 1003 883
rect 993 867 1007 880
rect 1056 827 1063 1176
rect 1096 1147 1103 1172
rect 1136 947 1143 1213
rect 1156 1047 1163 1273
rect 1276 1227 1283 1253
rect 1216 1180 1223 1183
rect 1213 1167 1227 1180
rect 1276 1027 1283 1173
rect 1296 1087 1303 1233
rect 1316 1186 1323 1393
rect 1336 1247 1343 1733
rect 1356 1247 1363 2033
rect 1376 1967 1383 2053
rect 1436 2027 1443 2116
rect 1456 2003 1463 2213
rect 1476 2047 1483 2192
rect 1496 2187 1503 2253
rect 1556 2220 1563 2223
rect 1553 2207 1567 2220
rect 1596 2216 1623 2223
rect 1496 2027 1503 2113
rect 1513 2027 1527 2033
rect 1427 1996 1463 2003
rect 1393 1960 1407 1973
rect 1433 1960 1447 1973
rect 1396 1956 1403 1960
rect 1436 1956 1443 1960
rect 1416 1920 1423 1923
rect 1376 1748 1383 1913
rect 1413 1907 1427 1920
rect 1396 1436 1403 1593
rect 1416 1567 1423 1703
rect 1436 1507 1443 1813
rect 1436 1436 1443 1493
rect 1456 1447 1463 1893
rect 1476 1827 1483 1973
rect 1516 1956 1523 2013
rect 1536 2007 1543 2073
rect 1576 1967 1583 2193
rect 1536 1920 1543 1923
rect 1533 1907 1547 1920
rect 1596 1926 1603 2173
rect 1616 2147 1623 2216
rect 1616 2107 1623 2133
rect 1636 2127 1643 2254
rect 1836 2256 1843 2293
rect 1676 2207 1683 2223
rect 1667 2196 1683 2207
rect 1667 2193 1680 2196
rect 1653 2147 1667 2153
rect 1716 2147 1723 2213
rect 1736 2167 1743 2253
rect 1656 1956 1663 2093
rect 1756 2067 1763 2213
rect 1776 2127 1783 2223
rect 1816 2220 1823 2223
rect 1813 2207 1827 2220
rect 1876 2207 1883 2373
rect 1896 2247 1903 2396
rect 1896 2207 1903 2233
rect 1827 2196 1843 2203
rect 1796 2147 1803 2173
rect 1816 2067 1823 2153
rect 1836 2107 1843 2196
rect 1716 1987 1723 2033
rect 1756 1968 1763 2032
rect 1836 2027 1843 2053
rect 1896 2047 1903 2172
rect 1916 2127 1923 2373
rect 1936 2287 1943 2393
rect 1976 2307 1983 2633
rect 2036 2627 2043 2933
rect 2056 2847 2063 2873
rect 2076 2827 2083 2973
rect 2116 2967 2123 2994
rect 2136 2943 2143 2963
rect 2136 2936 2163 2943
rect 2156 2807 2163 2936
rect 2056 2587 2063 2793
rect 2176 2787 2183 2933
rect 2196 2927 2203 3213
rect 2216 3087 2223 3333
rect 2276 3327 2283 3356
rect 2456 3347 2463 3653
rect 2496 3647 2503 3872
rect 2616 3843 2623 3993
rect 2616 3836 2633 3843
rect 2636 3787 2643 3833
rect 2656 3827 2663 4003
rect 2696 3983 2703 4003
rect 2676 3976 2703 3983
rect 2676 3827 2683 3976
rect 2716 3967 2723 3993
rect 2736 3947 2743 4212
rect 2756 4003 2763 4373
rect 2776 4187 2783 4413
rect 2796 4347 2803 4554
rect 2880 4553 2893 4556
rect 2916 4527 2923 4693
rect 2936 4567 2943 4753
rect 2956 4707 2963 4823
rect 2976 4556 2983 4693
rect 2996 4687 3003 4823
rect 3016 4767 3023 4813
rect 3016 4556 3023 4753
rect 3036 4647 3043 5033
rect 3036 4568 3043 4593
rect 2836 4423 2843 4453
rect 2856 4447 2863 4523
rect 2836 4416 2863 4423
rect 2816 4336 2823 4373
rect 2856 4336 2863 4416
rect 2896 4407 2903 4513
rect 2936 4307 2943 4513
rect 2996 4447 3003 4523
rect 3036 4427 3043 4473
rect 3056 4467 3063 5113
rect 3073 5107 3087 5116
rect 3093 5088 3107 5094
rect 3156 4987 3163 5252
rect 3233 5227 3247 5233
rect 3256 5207 3263 5376
rect 3316 5263 3323 5313
rect 3396 5287 3403 5413
rect 3476 5376 3483 5553
rect 3496 5447 3503 5594
rect 3636 5567 3643 5613
rect 3656 5587 3663 5831
rect 3696 5787 3703 5853
rect 3716 5747 3723 5933
rect 3767 5923 3780 5927
rect 3767 5913 3783 5923
rect 3776 5896 3783 5913
rect 3856 5907 3863 5973
rect 3796 5827 3803 5863
rect 3836 5860 3843 5863
rect 3833 5847 3847 5860
rect 3736 5596 3743 5793
rect 3836 5727 3843 5833
rect 3556 5507 3563 5563
rect 3456 5340 3463 5343
rect 3453 5327 3467 5340
rect 3316 5256 3343 5263
rect 3273 5247 3287 5253
rect 3273 5107 3287 5113
rect 3273 5080 3287 5093
rect 3276 5076 3283 5080
rect 3176 5043 3183 5074
rect 3316 5046 3323 5093
rect 3176 5036 3203 5043
rect 3136 4856 3143 4953
rect 3176 4867 3183 4993
rect 3076 4527 3083 4673
rect 3096 4567 3103 4773
rect 3116 4607 3123 4823
rect 3196 4823 3203 5036
rect 3153 4806 3167 4812
rect 3176 4816 3203 4823
rect 3176 4727 3183 4816
rect 3196 4647 3203 4753
rect 3216 4687 3223 5032
rect 3256 4987 3263 5043
rect 3236 4707 3243 4854
rect 3256 4727 3263 4823
rect 3287 4803 3300 4807
rect 3287 4793 3303 4803
rect 3136 4587 3143 4633
rect 3156 4556 3163 4613
rect 3056 4347 3063 4432
rect 2836 4300 2843 4303
rect 2796 4227 2803 4293
rect 2833 4287 2847 4300
rect 2836 4127 2843 4273
rect 2876 4263 2883 4303
rect 2976 4283 2983 4303
rect 3016 4283 3023 4292
rect 2976 4276 3003 4283
rect 3016 4280 3043 4283
rect 3016 4276 3047 4280
rect 2876 4260 2903 4263
rect 2876 4256 2907 4260
rect 2893 4247 2907 4256
rect 2876 4147 2883 4233
rect 2816 4036 2823 4073
rect 2876 4047 2883 4133
rect 2756 3996 2783 4003
rect 2776 3927 2783 3996
rect 2696 3816 2703 3873
rect 2516 3776 2543 3783
rect 2516 3707 2523 3776
rect 2596 3627 2603 3783
rect 2656 3767 2663 3792
rect 2796 3787 2803 4003
rect 2896 3987 2903 4193
rect 2956 4036 2963 4073
rect 2976 4067 2983 4213
rect 2996 4107 3003 4276
rect 3033 4267 3047 4276
rect 2973 4047 2987 4053
rect 2927 4003 2940 4007
rect 2927 3996 2943 4003
rect 2927 3993 2940 3996
rect 2833 3827 2847 3833
rect 2616 3667 2623 3713
rect 2487 3523 2500 3527
rect 2487 3516 2503 3523
rect 2487 3513 2500 3516
rect 2596 3516 2603 3613
rect 2676 3587 2683 3773
rect 2760 3783 2773 3787
rect 2756 3776 2773 3783
rect 2760 3773 2773 3776
rect 2653 3520 2667 3533
rect 2656 3516 2663 3520
rect 2516 3407 2523 3483
rect 2556 3427 2563 3483
rect 2596 3387 2603 3453
rect 2676 3367 2683 3473
rect 2696 3407 2703 3533
rect 2716 3487 2723 3772
rect 2816 3707 2823 3813
rect 2836 3667 2843 3773
rect 2856 3707 2863 3783
rect 2896 3780 2903 3783
rect 2893 3767 2907 3780
rect 2936 3767 2943 3973
rect 2816 3528 2823 3553
rect 2247 3323 2260 3327
rect 2247 3313 2263 3323
rect 2256 3296 2263 3313
rect 2296 3296 2303 3333
rect 2276 3260 2283 3263
rect 2316 3260 2323 3263
rect 2236 3063 2243 3253
rect 2273 3247 2287 3260
rect 2313 3247 2327 3260
rect 2216 3056 2243 3063
rect 2216 2903 2223 3056
rect 2276 3008 2283 3173
rect 2316 3047 2323 3233
rect 2356 3227 2363 3273
rect 2336 3147 2343 3173
rect 2320 3003 2333 3007
rect 2316 2996 2333 3003
rect 2320 2993 2333 2996
rect 2256 2907 2263 2963
rect 2356 2963 2363 3213
rect 2376 3127 2383 3313
rect 2416 3247 2423 3263
rect 2407 3236 2423 3247
rect 2407 3233 2420 3236
rect 2476 3207 2483 3263
rect 2536 3260 2543 3263
rect 2533 3247 2547 3260
rect 2416 3143 2423 3173
rect 2416 3140 2463 3143
rect 2416 3136 2467 3140
rect 2453 3127 2467 3136
rect 2336 2956 2363 2963
rect 2196 2896 2223 2903
rect 2196 2787 2203 2896
rect 2216 2776 2223 2813
rect 2156 2736 2183 2743
rect 1996 2307 2003 2573
rect 2076 2567 2083 2693
rect 2036 2507 2043 2553
rect 2096 2507 2103 2593
rect 2076 2476 2103 2483
rect 2096 2447 2103 2476
rect 2036 2347 2043 2443
rect 2116 2443 2123 2613
rect 2107 2436 2123 2443
rect 2033 2327 2047 2333
rect 2136 2307 2143 2593
rect 2156 2487 2163 2713
rect 2176 2607 2183 2736
rect 2196 2587 2203 2733
rect 2173 2480 2187 2493
rect 2216 2488 2223 2513
rect 2176 2476 2183 2480
rect 2256 2487 2263 2553
rect 2276 2527 2283 2853
rect 2296 2607 2303 2913
rect 2316 2787 2323 2893
rect 2336 2847 2343 2956
rect 2376 2947 2383 3053
rect 2416 3047 2423 3073
rect 2436 3067 2443 3113
rect 2436 3023 2443 3053
rect 2416 3016 2443 3023
rect 2416 2996 2423 3016
rect 2536 2996 2543 3053
rect 2556 3047 2563 3253
rect 2576 3247 2583 3353
rect 2576 3087 2583 3173
rect 2573 3000 2587 3013
rect 2596 3007 2603 3352
rect 2576 2996 2583 3000
rect 2393 2947 2407 2953
rect 2416 2787 2423 2933
rect 2496 2887 2503 2994
rect 2436 2783 2443 2833
rect 2436 2776 2463 2783
rect 2336 2740 2343 2743
rect 2316 2647 2323 2733
rect 2333 2727 2347 2740
rect 2296 2487 2303 2572
rect 2316 2476 2323 2633
rect 2396 2607 2403 2743
rect 2416 2627 2423 2733
rect 2516 2727 2523 2753
rect 2536 2743 2543 2933
rect 2596 2907 2603 2953
rect 2616 2927 2623 3013
rect 2636 2867 2643 3153
rect 2656 3007 2663 3233
rect 2696 3223 2703 3333
rect 2716 3247 2723 3433
rect 2836 3347 2843 3653
rect 2856 3647 2863 3693
rect 2896 3607 2903 3633
rect 2956 3567 2963 3933
rect 2996 3923 3003 4093
rect 3016 4043 3023 4253
rect 3036 4147 3043 4213
rect 3076 4087 3083 4433
rect 3096 4427 3103 4513
rect 3136 4336 3143 4413
rect 3176 4343 3183 4453
rect 3196 4447 3203 4573
rect 3233 4560 3247 4573
rect 3236 4556 3243 4560
rect 3276 4556 3283 4733
rect 3296 4727 3303 4793
rect 3316 4607 3323 4812
rect 3336 4787 3343 5256
rect 3396 5207 3403 5252
rect 3416 5167 3423 5313
rect 3496 5167 3503 5332
rect 3616 5327 3623 5343
rect 3616 5203 3623 5313
rect 3616 5196 3643 5203
rect 3367 5093 3373 5107
rect 3360 5086 3380 5087
rect 3367 5083 3380 5086
rect 3367 5076 3383 5083
rect 3416 5076 3423 5153
rect 3433 5107 3447 5113
rect 3453 5088 3467 5094
rect 3367 5073 3380 5076
rect 3496 5067 3503 5093
rect 3356 4927 3363 5033
rect 3436 5040 3443 5043
rect 3433 5027 3447 5040
rect 3476 4947 3483 5033
rect 3516 5027 3523 5193
rect 3553 5080 3567 5093
rect 3556 5076 3563 5080
rect 3596 5076 3603 5193
rect 3416 4856 3423 4913
rect 3456 4868 3463 4913
rect 3496 4827 3503 4973
rect 3436 4820 3443 4823
rect 3433 4807 3447 4820
rect 3486 4813 3487 4820
rect 3473 4803 3487 4813
rect 3473 4800 3503 4803
rect 3476 4796 3503 4800
rect 3316 4527 3323 4593
rect 3356 4556 3363 4633
rect 3396 4556 3443 4563
rect 3256 4387 3263 4523
rect 3416 4487 3423 4513
rect 3276 4407 3283 4473
rect 3176 4336 3203 4343
rect 3116 4267 3123 4303
rect 3156 4247 3163 4303
rect 3016 4036 3033 4043
rect 3016 3947 3023 4012
rect 2976 3916 3003 3923
rect 2976 3827 2983 3916
rect 3116 3823 3123 4053
rect 3136 3847 3143 4053
rect 3156 4007 3163 4113
rect 3176 4047 3183 4093
rect 3196 4067 3203 4336
rect 3216 4067 3223 4373
rect 3233 4343 3247 4353
rect 3233 4340 3263 4343
rect 3236 4336 3263 4340
rect 3296 4336 3303 4433
rect 3236 4127 3243 4273
rect 3276 4127 3283 4303
rect 3356 4167 3363 4473
rect 3436 4467 3443 4556
rect 3456 4527 3463 4693
rect 3476 4567 3483 4733
rect 3496 4587 3503 4796
rect 3516 4707 3523 4793
rect 3487 4563 3500 4567
rect 3487 4556 3503 4563
rect 3536 4556 3543 4653
rect 3556 4567 3563 4673
rect 3487 4553 3500 4556
rect 3416 4348 3423 4433
rect 3436 4367 3443 4453
rect 3456 4347 3463 4393
rect 3476 4367 3483 4513
rect 3496 4343 3503 4473
rect 3476 4336 3503 4343
rect 3536 4336 3543 4493
rect 3576 4347 3583 4773
rect 3396 4227 3403 4303
rect 3236 4043 3243 4113
rect 3216 4036 3263 4043
rect 3156 3867 3163 3953
rect 3176 3843 3183 3913
rect 3156 3836 3183 3843
rect 3096 3816 3123 3823
rect 3156 3816 3163 3836
rect 3196 3816 3203 3953
rect 3256 3887 3263 4036
rect 2996 3780 3003 3783
rect 2993 3767 3007 3780
rect 3036 3776 3053 3783
rect 2856 3483 2863 3553
rect 2976 3487 2983 3533
rect 3013 3520 3027 3533
rect 3056 3528 3063 3772
rect 3076 3767 3083 3813
rect 3096 3747 3103 3816
rect 3136 3780 3143 3783
rect 3133 3767 3147 3780
rect 3116 3567 3123 3613
rect 3016 3516 3023 3520
rect 3116 3516 3123 3553
rect 3216 3547 3223 3773
rect 2856 3476 2873 3483
rect 3036 3480 3043 3483
rect 2696 3216 2723 3223
rect 2716 3008 2723 3216
rect 2736 3107 2743 3313
rect 2756 3308 2763 3333
rect 2856 3323 2863 3413
rect 2793 3300 2807 3313
rect 2836 3316 2863 3323
rect 2796 3296 2803 3300
rect 2836 3296 2843 3316
rect 2776 3207 2783 3263
rect 2536 2736 2563 2743
rect 2576 2740 2583 2743
rect 2396 2567 2403 2593
rect 1973 2260 1987 2272
rect 1976 2256 1983 2260
rect 1936 2220 1943 2223
rect 1933 2207 1947 2220
rect 1916 1985 1923 2092
rect 1936 2067 1943 2113
rect 1976 2067 1983 2153
rect 1996 2107 2003 2272
rect 2016 2187 2023 2254
rect 2036 2087 2043 2292
rect 2056 2147 2063 2293
rect 2076 2123 2083 2212
rect 2056 2116 2083 2123
rect 1936 2007 1943 2032
rect 1916 1978 1953 1985
rect 1696 1956 1743 1963
rect 1573 1907 1587 1913
rect 1416 1327 1423 1403
rect 1416 1243 1423 1313
rect 1396 1236 1423 1243
rect 1340 1226 1360 1227
rect 1347 1223 1360 1226
rect 1347 1216 1363 1223
rect 1396 1216 1403 1236
rect 1347 1214 1360 1216
rect 1313 1167 1327 1172
rect 1076 886 1083 933
rect 1113 920 1127 933
rect 1116 916 1123 920
rect 1156 916 1163 973
rect 1316 928 1323 1033
rect 1456 1007 1463 1233
rect 1476 1027 1483 1533
rect 1496 1507 1503 1703
rect 1536 1487 1543 1703
rect 1576 1547 1583 1753
rect 1596 1523 1603 1833
rect 1676 1768 1683 1923
rect 1736 1907 1743 1956
rect 1896 1927 1903 1973
rect 2016 1956 2023 2013
rect 2036 1987 2043 2073
rect 2056 2047 2063 2116
rect 2096 2027 2103 2113
rect 2116 2067 2123 2193
rect 1633 1740 1647 1753
rect 1636 1736 1643 1740
rect 1736 1706 1743 1753
rect 1587 1516 1603 1523
rect 1576 1436 1583 1512
rect 1656 1467 1663 1692
rect 1496 1307 1503 1393
rect 1516 1263 1523 1403
rect 1616 1267 1623 1453
rect 1676 1448 1683 1633
rect 1716 1436 1723 1513
rect 1736 1447 1743 1593
rect 1756 1587 1763 1913
rect 1776 1907 1783 1923
rect 1776 1787 1783 1893
rect 1816 1807 1823 1913
rect 1836 1787 1843 1923
rect 1896 1807 1903 1833
rect 1916 1827 1923 1953
rect 1816 1700 1823 1703
rect 1776 1563 1783 1693
rect 1813 1687 1827 1700
rect 1836 1587 1843 1673
rect 1767 1556 1783 1563
rect 1756 1406 1763 1552
rect 1813 1440 1827 1453
rect 1856 1448 1863 1703
rect 1816 1436 1823 1440
rect 1876 1443 1883 1693
rect 1896 1687 1903 1793
rect 1936 1787 1943 1913
rect 1896 1567 1903 1613
rect 1916 1467 1923 1773
rect 1956 1763 1963 1893
rect 2056 1787 2063 2012
rect 2136 1988 2143 2223
rect 2156 2167 2163 2433
rect 2240 2443 2253 2447
rect 2236 2436 2253 2443
rect 2240 2433 2253 2436
rect 2156 2047 2163 2073
rect 2176 2027 2183 2293
rect 2196 2287 2203 2333
rect 2236 2256 2243 2293
rect 2276 2267 2283 2473
rect 2376 2367 2383 2513
rect 2296 2227 2303 2353
rect 2356 2256 2363 2353
rect 2076 1867 2083 1973
rect 2096 1847 2103 1913
rect 2116 1807 2123 1923
rect 2136 1787 2143 1853
rect 2156 1827 2163 1923
rect 1956 1756 1983 1763
rect 1976 1748 1983 1756
rect 2016 1736 2023 1773
rect 2076 1703 2083 1733
rect 1956 1700 1963 1703
rect 1953 1687 1967 1700
rect 1956 1627 1963 1673
rect 1936 1507 1943 1593
rect 1956 1448 1963 1573
rect 1996 1507 2003 1703
rect 2036 1667 2043 1703
rect 2076 1696 2103 1703
rect 2076 1627 2083 1673
rect 2016 1487 2023 1533
rect 2096 1523 2103 1696
rect 2116 1627 2123 1703
rect 2156 1687 2163 1703
rect 2147 1676 2163 1687
rect 2147 1673 2160 1676
rect 2196 1667 2203 1913
rect 2136 1607 2143 1652
rect 2216 1567 2223 2173
rect 2296 2167 2303 2192
rect 2236 1927 2243 2153
rect 2316 2007 2323 2213
rect 2356 2087 2363 2173
rect 2296 1956 2323 1963
rect 2256 1787 2263 1923
rect 2316 1867 2323 1956
rect 2316 1767 2323 1853
rect 2336 1807 2343 1933
rect 2356 1767 2363 2073
rect 2396 1983 2403 2493
rect 2436 2476 2443 2653
rect 2456 2547 2463 2673
rect 2496 2476 2503 2593
rect 2516 2447 2523 2493
rect 2456 2287 2463 2432
rect 2476 2256 2483 2353
rect 2513 2287 2527 2293
rect 2516 2256 2523 2273
rect 2536 2267 2543 2473
rect 2556 2347 2563 2736
rect 2573 2727 2587 2740
rect 2636 2667 2643 2743
rect 2676 2727 2683 2813
rect 2696 2767 2703 2963
rect 2716 2727 2723 2933
rect 2736 2927 2743 2963
rect 2756 2807 2763 2933
rect 2776 2887 2783 3013
rect 2816 3007 2823 3263
rect 2776 2776 2783 2813
rect 2796 2807 2803 2994
rect 2836 2996 2843 3193
rect 2876 3127 2883 3472
rect 3033 3467 3047 3480
rect 2916 3296 2923 3373
rect 2976 3267 2983 3393
rect 2936 3127 2943 3263
rect 2996 3187 3003 3433
rect 3076 3427 3083 3483
rect 3016 3227 3023 3333
rect 2936 3008 2943 3073
rect 3016 3027 3023 3093
rect 3016 2996 3023 3013
rect 2936 2967 2943 2994
rect 2856 2960 2863 2963
rect 2896 2960 2903 2963
rect 2853 2947 2867 2960
rect 2893 2947 2907 2960
rect 3036 2960 3043 2963
rect 2996 2943 3003 2952
rect 3033 2947 3047 2960
rect 2996 2936 3023 2943
rect 2816 2776 2823 2873
rect 2716 2647 2723 2673
rect 2596 2507 2603 2633
rect 2736 2627 2743 2733
rect 2796 2740 2803 2743
rect 2793 2727 2807 2740
rect 2616 2476 2623 2613
rect 2636 2487 2643 2593
rect 2416 2127 2423 2213
rect 2436 2047 2443 2093
rect 2376 1980 2403 1983
rect 2373 1976 2403 1980
rect 2373 1967 2387 1976
rect 2436 1956 2443 2033
rect 2456 1987 2463 2223
rect 2273 1740 2287 1753
rect 2376 1747 2383 1913
rect 2476 1907 2483 1923
rect 2276 1736 2283 1740
rect 2316 1736 2363 1743
rect 2256 1667 2263 1703
rect 2296 1700 2303 1703
rect 2293 1687 2307 1700
rect 2256 1547 2263 1653
rect 2076 1516 2103 1523
rect 1876 1436 1903 1443
rect 1656 1367 1663 1403
rect 1496 1256 1523 1263
rect 1496 1227 1503 1256
rect 1533 1243 1547 1253
rect 1516 1240 1547 1243
rect 1516 1236 1543 1240
rect 1516 1216 1523 1236
rect 1693 1220 1707 1233
rect 1696 1216 1703 1220
rect 1576 1180 1583 1183
rect 1573 1167 1587 1180
rect 1236 916 1263 923
rect 656 656 703 663
rect 613 400 627 413
rect 616 396 623 400
rect 296 307 303 363
rect 316 356 333 363
rect 260 183 273 187
rect 256 176 273 183
rect 260 174 273 176
rect 296 146 303 213
rect 316 188 323 356
rect 336 203 343 233
rect 356 227 363 393
rect 516 367 523 394
rect 656 367 663 413
rect 556 307 563 363
rect 596 267 603 363
rect 676 327 683 453
rect 696 407 703 433
rect 736 408 743 573
rect 796 447 803 693
rect 816 423 823 733
rect 896 696 903 733
rect 936 703 943 773
rect 956 727 963 813
rect 936 696 963 703
rect 956 666 963 696
rect 1056 696 1063 733
rect 876 547 883 663
rect 916 423 923 652
rect 996 627 1003 663
rect 816 416 843 423
rect 776 396 823 403
rect 716 366 722 369
rect 816 367 823 396
rect 707 365 722 366
rect 707 363 720 365
rect 707 356 723 363
rect 707 353 720 356
rect 336 196 363 203
rect 356 176 363 196
rect 393 180 407 193
rect 396 176 403 180
rect 196 107 203 143
rect 327 143 340 147
rect 327 136 343 143
rect 376 140 383 143
rect 327 133 340 136
rect 373 127 387 140
rect 436 127 443 173
rect 496 87 503 143
rect 536 107 543 143
rect 596 87 603 232
rect 676 188 683 313
rect 736 107 743 333
rect 756 327 763 363
rect 796 287 803 353
rect 836 347 843 416
rect 896 416 923 423
rect 896 396 903 416
rect 936 396 943 533
rect 1096 527 1103 813
rect 1176 807 1183 883
rect 1236 847 1243 916
rect 1336 886 1343 993
rect 1456 916 1463 993
rect 1153 723 1167 733
rect 1176 723 1183 793
rect 1153 720 1183 723
rect 1156 716 1183 720
rect 1156 696 1163 716
rect 1236 707 1243 833
rect 1316 727 1323 753
rect 1396 727 1403 813
rect 1373 708 1387 713
rect 1256 696 1303 703
rect 1116 487 1123 693
rect 856 303 863 353
rect 876 323 883 363
rect 916 360 923 363
rect 913 347 927 360
rect 876 316 903 323
rect 856 296 873 303
rect 836 176 843 273
rect 856 207 863 253
rect 816 107 823 143
rect 876 127 883 293
rect 896 247 903 316
rect 976 307 983 473
rect 1033 400 1047 413
rect 1076 408 1083 433
rect 1036 396 1043 400
rect 1016 327 1023 363
rect 1056 307 1063 363
rect 1116 307 1123 413
rect 1156 396 1163 473
rect 1196 396 1203 573
rect 1256 447 1263 696
rect 1396 666 1403 713
rect 1376 627 1383 653
rect 1416 647 1423 793
rect 1436 707 1443 883
rect 1447 696 1463 703
rect 1496 696 1503 1113
rect 1516 747 1523 1073
rect 1556 916 1563 1073
rect 1596 987 1603 1173
rect 1656 886 1663 1153
rect 1676 928 1683 1183
rect 1736 1047 1743 1293
rect 1796 1247 1803 1403
rect 1816 1223 1823 1273
rect 1896 1247 1903 1436
rect 1993 1440 2007 1453
rect 1996 1436 2003 1440
rect 1796 1216 1843 1223
rect 1836 1186 1843 1216
rect 1776 1087 1783 1183
rect 1856 1087 1863 1233
rect 1956 1216 1963 1253
rect 1976 1227 1983 1253
rect 1936 1180 1943 1183
rect 1933 1167 1947 1180
rect 1776 943 1783 1073
rect 1756 936 1783 943
rect 1756 916 1763 936
rect 1876 916 1883 1013
rect 1976 923 1983 1173
rect 1996 1027 2003 1213
rect 2016 1167 2023 1392
rect 2036 1267 2043 1393
rect 2056 1243 2063 1493
rect 2076 1347 2083 1516
rect 2093 1447 2107 1453
rect 2076 1267 2083 1333
rect 2036 1240 2063 1243
rect 2033 1236 2063 1240
rect 2033 1227 2047 1236
rect 2116 1216 2123 1253
rect 2176 1227 2183 1373
rect 2196 1228 2203 1453
rect 2236 1347 2243 1403
rect 2236 1227 2243 1293
rect 2056 1180 2063 1183
rect 2096 1180 2103 1183
rect 1956 916 1983 923
rect 1476 660 1483 663
rect 1473 647 1487 660
rect 1556 567 1563 733
rect 1233 400 1247 413
rect 1236 396 1243 400
rect 1216 360 1223 363
rect 1213 347 1227 360
rect 936 176 943 233
rect 956 207 963 233
rect 1016 147 1023 174
rect 956 140 963 143
rect 953 127 967 140
rect 1033 143 1047 153
rect 1033 140 1063 143
rect 1036 136 1063 140
rect 1056 87 1063 136
rect 1116 67 1123 143
rect 1136 107 1143 213
rect 1216 176 1223 253
rect 1276 227 1283 513
rect 1296 366 1303 413
rect 1396 396 1403 493
rect 1336 347 1343 363
rect 1327 336 1343 347
rect 1327 333 1340 336
rect 1267 173 1273 187
rect 1156 146 1163 173
rect 1296 146 1303 313
rect 1313 188 1327 193
rect 1393 180 1407 193
rect 1396 176 1403 180
rect 1196 87 1203 143
rect 1356 67 1363 113
rect 1376 87 1383 143
rect 1436 27 1443 553
rect 1513 400 1527 413
rect 1516 396 1523 400
rect 1556 396 1563 493
rect 1576 487 1583 793
rect 1616 747 1623 883
rect 1736 880 1743 883
rect 1733 867 1747 880
rect 1896 807 1903 883
rect 1640 703 1653 707
rect 1636 696 1653 703
rect 1640 693 1653 696
rect 1773 700 1787 713
rect 1776 696 1783 700
rect 1616 660 1623 663
rect 1613 647 1627 660
rect 1576 408 1583 473
rect 1616 427 1623 633
rect 1633 400 1647 413
rect 1636 396 1643 400
rect 1676 396 1683 673
rect 1696 427 1703 693
rect 1756 660 1763 663
rect 1753 647 1767 660
rect 1456 366 1463 393
rect 1496 307 1503 363
rect 1516 176 1523 313
rect 1656 307 1663 363
rect 1736 307 1743 533
rect 1796 507 1803 663
rect 1836 527 1843 713
rect 1916 696 1923 733
rect 1956 707 1963 916
rect 2036 923 2043 1173
rect 2053 1167 2067 1180
rect 2093 1167 2107 1180
rect 2156 1167 2163 1213
rect 2036 916 2063 923
rect 1976 876 1993 883
rect 1896 660 1903 663
rect 1893 647 1907 660
rect 1936 587 1943 652
rect 1976 647 1983 876
rect 2056 787 2063 916
rect 2076 886 2083 1013
rect 2116 916 2123 953
rect 2156 928 2163 1073
rect 2136 747 2143 883
rect 2056 696 2063 733
rect 2156 696 2163 773
rect 2196 767 2203 913
rect 2216 727 2223 1033
rect 2256 967 2263 1233
rect 2276 1227 2283 1333
rect 2296 1247 2303 1593
rect 2316 1406 2323 1493
rect 2356 1467 2363 1736
rect 2416 1736 2423 1853
rect 2476 1823 2483 1893
rect 2536 1847 2543 2212
rect 2556 1987 2563 2293
rect 2576 1963 2583 2273
rect 2596 2267 2603 2432
rect 2616 2256 2623 2333
rect 2636 2327 2643 2419
rect 2656 2267 2663 2613
rect 2596 2067 2603 2213
rect 2636 2187 2643 2223
rect 2656 2127 2663 2213
rect 2676 2207 2683 2573
rect 2756 2507 2763 2711
rect 2796 2587 2803 2713
rect 2836 2627 2843 2733
rect 2856 2527 2863 2793
rect 2916 2776 2923 2873
rect 2896 2740 2903 2743
rect 2893 2727 2907 2740
rect 2913 2707 2927 2713
rect 2896 2647 2903 2673
rect 2736 2407 2743 2443
rect 2696 2267 2703 2373
rect 2836 2363 2843 2493
rect 2856 2446 2863 2513
rect 2956 2476 2963 2553
rect 2996 2488 3003 2773
rect 3016 2607 3023 2936
rect 3076 2927 3083 3213
rect 3096 3107 3103 3473
rect 3196 3427 3203 3472
rect 3216 3467 3223 3512
rect 3116 3308 3123 3373
rect 3236 3347 3243 3853
rect 3276 3847 3283 4073
rect 3296 4047 3303 4153
rect 3316 4036 3323 4133
rect 3356 4036 3363 4093
rect 3396 4067 3403 4153
rect 3436 4087 3443 4292
rect 3456 4107 3463 4292
rect 3476 4187 3483 4336
rect 3516 4267 3523 4303
rect 3476 4127 3483 4173
rect 3396 3987 3403 4053
rect 3453 4040 3467 4053
rect 3456 4036 3463 4040
rect 3516 4047 3523 4253
rect 3416 3996 3443 4003
rect 3336 3828 3343 3971
rect 3356 3847 3363 3913
rect 3416 3907 3423 3996
rect 3436 3847 3443 3973
rect 3496 3907 3503 3973
rect 3536 3967 3543 4113
rect 3556 4047 3563 4133
rect 3596 4067 3603 4893
rect 3616 4867 3623 5033
rect 3636 4987 3643 5196
rect 3656 4967 3663 5173
rect 3676 4927 3683 5253
rect 3656 4888 3663 4913
rect 3696 4907 3703 5563
rect 3776 5487 3783 5653
rect 3856 5596 3863 5853
rect 3876 5807 3883 6033
rect 3896 5707 3903 6053
rect 3936 6023 3943 6116
rect 3996 6063 4003 6083
rect 3916 6016 3943 6023
rect 3976 6056 4003 6063
rect 3916 5967 3923 6016
rect 3916 5907 3923 5953
rect 3976 5927 3983 6056
rect 4036 6047 4043 6173
rect 4136 6116 4143 6153
rect 3960 5923 3973 5927
rect 3956 5913 3973 5923
rect 3956 5896 3963 5913
rect 3996 5896 4003 5953
rect 3816 5447 3823 5563
rect 3876 5507 3883 5594
rect 3816 5376 3823 5412
rect 3896 5376 3903 5693
rect 3916 5647 3923 5833
rect 3936 5667 3943 5852
rect 3953 5827 3967 5833
rect 3976 5767 3983 5863
rect 4056 5866 4063 6113
rect 4196 6107 4203 6153
rect 4276 6116 4283 6153
rect 4116 6063 4123 6083
rect 4116 6056 4143 6063
rect 4136 5908 4143 6056
rect 4087 5903 4100 5907
rect 4087 5896 4103 5903
rect 4087 5894 4100 5896
rect 4176 5907 4183 6053
rect 4216 6047 4223 6114
rect 4316 6087 4323 6173
rect 4413 6120 4427 6133
rect 4416 6116 4423 6120
rect 4256 6080 4263 6083
rect 4253 6067 4267 6080
rect 4236 6007 4243 6033
rect 3996 5767 4003 5813
rect 4016 5747 4023 5852
rect 4033 5847 4047 5853
rect 4156 5727 4163 5863
rect 4176 5667 4183 5853
rect 4196 5727 4203 5953
rect 3973 5600 3987 5613
rect 3976 5596 3983 5600
rect 4016 5567 4023 5653
rect 4216 5627 4223 5913
rect 4236 5907 4243 5993
rect 4256 5967 4263 6053
rect 4276 5896 4283 5973
rect 4316 5896 4323 5933
rect 4336 5907 4343 6093
rect 4376 5947 4383 5973
rect 4396 5927 4403 6083
rect 4187 5623 4200 5627
rect 4187 5613 4203 5623
rect 4113 5600 4127 5613
rect 4116 5596 4123 5600
rect 4196 5596 4203 5613
rect 3756 5340 3763 5343
rect 3753 5327 3767 5340
rect 3716 5076 3723 5153
rect 3796 5127 3803 5332
rect 3856 5167 3863 5374
rect 3960 5343 3973 5347
rect 3916 5340 3923 5343
rect 3913 5327 3927 5340
rect 3956 5336 3973 5343
rect 3960 5333 3973 5336
rect 3876 5047 3883 5074
rect 3756 5023 3763 5043
rect 3807 5043 3820 5046
rect 3807 5040 3823 5043
rect 3807 5033 3827 5040
rect 3813 5027 3827 5033
rect 3756 5016 3783 5023
rect 3716 4863 3723 4993
rect 3696 4856 3723 4863
rect 3736 4826 3743 4913
rect 3636 4687 3643 4812
rect 3656 4647 3663 4733
rect 3636 4556 3643 4593
rect 3676 4567 3683 4812
rect 3736 4707 3743 4812
rect 3756 4683 3763 4953
rect 3776 4867 3783 5016
rect 3876 5007 3883 5033
rect 3896 4967 3903 5113
rect 3936 5076 3943 5153
rect 3956 5023 3963 5032
rect 3936 5016 3963 5023
rect 3793 4860 3807 4873
rect 3796 4856 3803 4860
rect 3836 4856 3843 4933
rect 3936 4867 3943 5016
rect 3996 4907 4003 5433
rect 4016 5347 4023 5413
rect 4076 5376 4083 5533
rect 4096 5507 4103 5563
rect 4156 5527 4163 5573
rect 4216 5556 4243 5563
rect 4176 5383 4183 5533
rect 4236 5427 4243 5556
rect 4256 5507 4263 5793
rect 4336 5767 4343 5853
rect 4356 5707 4363 5913
rect 4413 5900 4427 5913
rect 4456 5908 4463 5933
rect 4416 5896 4423 5900
rect 4356 5627 4363 5693
rect 4376 5647 4383 5853
rect 4396 5807 4403 5863
rect 4396 5747 4403 5793
rect 4436 5787 4443 5863
rect 4476 5827 4483 5853
rect 4496 5847 4503 6213
rect 4687 6176 4713 6183
rect 4547 6134 4553 6147
rect 4547 6133 4560 6134
rect 4536 5947 4543 6033
rect 4556 5967 4563 6053
rect 4576 6007 4583 6083
rect 4616 6027 4623 6073
rect 4636 6067 4643 6133
rect 4696 6128 4703 6153
rect 4736 6116 4743 6153
rect 4876 6116 4883 6153
rect 4976 6147 4983 6213
rect 5616 6187 5623 6213
rect 4676 6080 4683 6083
rect 4673 6067 4687 6080
rect 4573 5900 4587 5913
rect 4616 5908 4623 5973
rect 4576 5896 4583 5900
rect 4496 5787 4503 5833
rect 4516 5727 4523 5893
rect 4556 5747 4563 5863
rect 4596 5860 4603 5863
rect 4593 5847 4607 5860
rect 4656 5866 4663 5933
rect 4687 5903 4700 5907
rect 4687 5896 4703 5903
rect 4736 5896 4743 6033
rect 4687 5893 4700 5896
rect 4636 5827 4643 5853
rect 4316 5467 4323 5563
rect 4356 5547 4363 5592
rect 4416 5527 4423 5563
rect 4176 5376 4203 5383
rect 4056 5340 4063 5343
rect 4053 5327 4067 5340
rect 4096 5327 4103 5343
rect 4136 5327 4143 5374
rect 4016 4987 4023 5312
rect 4096 5107 4103 5313
rect 4116 5076 4123 5113
rect 4136 5087 4143 5292
rect 4176 5083 4183 5376
rect 4316 5346 4323 5453
rect 4476 5443 4483 5633
rect 4536 5608 4543 5633
rect 4496 5527 4503 5594
rect 4476 5436 4503 5443
rect 4416 5376 4423 5413
rect 4296 5336 4313 5343
rect 4336 5287 4343 5374
rect 4476 5346 4483 5413
rect 4156 5076 4183 5083
rect 4056 5040 4063 5043
rect 4096 5040 4103 5043
rect 4053 5027 4067 5040
rect 4093 5027 4107 5040
rect 4133 5027 4147 5033
rect 4036 4867 4043 4953
rect 3816 4803 3823 4823
rect 3853 4807 3867 4812
rect 3816 4796 3843 4803
rect 3736 4676 3763 4683
rect 3616 4068 3623 4493
rect 3656 4383 3663 4453
rect 3676 4447 3683 4493
rect 3696 4467 3703 4613
rect 3736 4607 3743 4676
rect 3756 4627 3763 4653
rect 3776 4587 3783 4673
rect 3816 4526 3823 4753
rect 3836 4707 3843 4796
rect 3916 4767 3923 4853
rect 3976 4820 3983 4823
rect 3736 4520 3743 4523
rect 3733 4507 3747 4520
rect 3776 4516 3803 4523
rect 3773 4487 3787 4493
rect 3656 4376 3683 4383
rect 3676 4363 3683 4376
rect 3716 4363 3723 4393
rect 3676 4356 3723 4363
rect 3567 4043 3580 4047
rect 3567 4036 3583 4043
rect 3567 4033 3580 4036
rect 3636 4043 3643 4333
rect 3656 4267 3663 4303
rect 3696 4187 3703 4213
rect 3636 4036 3663 4043
rect 3556 3907 3563 3993
rect 3316 3747 3323 3783
rect 3316 3627 3323 3733
rect 3336 3587 3343 3753
rect 3296 3447 3303 3483
rect 3096 2947 3103 2993
rect 3116 2963 3123 3294
rect 3136 3266 3143 3333
rect 3296 3303 3303 3433
rect 3356 3308 3363 3773
rect 3376 3567 3383 3783
rect 3276 3296 3303 3303
rect 3256 3263 3263 3293
rect 3216 3256 3263 3263
rect 3276 3227 3283 3296
rect 3336 3260 3343 3263
rect 3216 3167 3223 3193
rect 3296 3167 3303 3253
rect 3333 3247 3347 3260
rect 3376 3187 3383 3532
rect 3396 3516 3403 3693
rect 3436 3387 3443 3483
rect 3456 3367 3463 3753
rect 3476 3727 3483 3873
rect 3496 3707 3503 3893
rect 3556 3816 3563 3853
rect 3476 3447 3483 3613
rect 3496 3483 3503 3633
rect 3516 3527 3523 3673
rect 3556 3516 3563 3713
rect 3596 3687 3603 3833
rect 3616 3767 3623 3893
rect 3636 3847 3643 3993
rect 3656 3823 3663 4036
rect 3676 4007 3683 4093
rect 3716 4067 3723 4292
rect 3736 4207 3743 4334
rect 3756 4287 3763 4353
rect 3776 4307 3783 4433
rect 3796 4427 3803 4516
rect 3816 4363 3823 4512
rect 3836 4507 3843 4693
rect 3856 4607 3863 4733
rect 3916 4556 3923 4673
rect 3936 4647 3943 4813
rect 3973 4807 3987 4820
rect 4016 4807 4023 4823
rect 3996 4796 4013 4803
rect 3996 4783 4003 4796
rect 4036 4783 4043 4813
rect 3956 4776 4003 4783
rect 4016 4776 4043 4783
rect 3853 4507 3867 4512
rect 3896 4427 3903 4523
rect 3847 4403 3860 4407
rect 3847 4393 3863 4403
rect 3796 4356 3823 4363
rect 3736 4087 3743 4113
rect 3736 4036 3743 4073
rect 3776 4036 3783 4093
rect 3796 4087 3803 4356
rect 3856 4348 3863 4393
rect 3896 4303 3903 4353
rect 3816 4287 3823 4303
rect 3876 4296 3903 4303
rect 3827 4276 3843 4283
rect 3816 4047 3823 4173
rect 3836 4147 3843 4276
rect 3893 4207 3907 4213
rect 3916 4207 3923 4493
rect 3956 4367 3963 4776
rect 4016 4763 4023 4776
rect 3976 4756 4023 4763
rect 3976 4587 3983 4756
rect 4033 4743 4047 4753
rect 4016 4740 4047 4743
rect 4016 4736 4043 4740
rect 3996 4563 4003 4733
rect 4016 4607 4023 4736
rect 4056 4667 4063 4893
rect 4116 4856 4123 4973
rect 4156 4907 4163 5076
rect 4236 5023 4243 5032
rect 4216 5016 4243 5023
rect 4216 4947 4223 5016
rect 4196 4868 4203 4893
rect 4076 4826 4083 4853
rect 4107 4763 4120 4767
rect 4107 4753 4123 4763
rect 4076 4687 4083 4713
rect 3987 4556 4003 4563
rect 4056 4556 4063 4632
rect 4076 4583 4083 4673
rect 4096 4627 4103 4732
rect 4116 4587 4123 4753
rect 4076 4576 4103 4583
rect 4096 4556 4103 4576
rect 3976 4447 3983 4552
rect 3996 4423 4003 4513
rect 4036 4467 4043 4491
rect 4076 4467 4083 4523
rect 4136 4487 4143 4613
rect 3976 4416 4003 4423
rect 3976 4336 3983 4416
rect 4016 4347 4023 4433
rect 3956 4267 3963 4303
rect 3893 4167 3907 4172
rect 3893 4160 3913 4167
rect 3896 4156 3913 4160
rect 3900 4153 3913 4156
rect 3896 4087 3903 4133
rect 3807 4036 3823 4047
rect 3807 4033 3820 4036
rect 3716 4000 3723 4003
rect 3713 3987 3727 4000
rect 3756 3983 3763 4003
rect 3756 3976 3783 3983
rect 3636 3816 3663 3823
rect 3693 3820 3707 3833
rect 3696 3816 3703 3820
rect 3596 3516 3603 3652
rect 3636 3607 3643 3816
rect 3676 3647 3683 3783
rect 3716 3747 3723 3783
rect 3736 3687 3743 3713
rect 3636 3528 3643 3553
rect 3693 3520 3707 3533
rect 3716 3527 3723 3633
rect 3696 3516 3703 3520
rect 3736 3507 3743 3553
rect 3496 3476 3523 3483
rect 3436 3296 3443 3333
rect 3416 3207 3423 3263
rect 3456 3260 3463 3263
rect 3453 3247 3467 3260
rect 3116 2956 3133 2963
rect 3053 2780 3067 2793
rect 3056 2776 3063 2780
rect 3096 2776 3103 2933
rect 3156 2747 3163 2913
rect 3196 2907 3203 3093
rect 3196 2776 3203 2893
rect 3216 2827 3223 3113
rect 3276 2996 3283 3073
rect 3316 3008 3323 3173
rect 3360 3143 3373 3147
rect 3356 3140 3373 3143
rect 3353 3133 3373 3140
rect 3353 3127 3367 3133
rect 3256 2960 3263 2963
rect 3236 2867 3243 2952
rect 3253 2947 3267 2960
rect 2816 2356 2843 2363
rect 3016 2363 3023 2432
rect 3076 2363 3083 2593
rect 3096 2407 3103 2713
rect 3216 2707 3223 2743
rect 3256 2727 3263 2933
rect 3276 2743 3283 2813
rect 3296 2787 3303 2963
rect 3347 2963 3360 2967
rect 3347 2956 3363 2963
rect 3347 2953 3360 2956
rect 3336 2776 3343 2913
rect 3416 2827 3423 3172
rect 3476 3127 3483 3193
rect 3496 3087 3503 3213
rect 3516 3187 3523 3476
rect 3576 3427 3583 3483
rect 3756 3483 3763 3933
rect 3776 3923 3783 3976
rect 3796 3947 3803 3993
rect 3816 3923 3823 3953
rect 3776 3916 3823 3923
rect 3776 3707 3783 3853
rect 3836 3816 3843 3913
rect 3896 3903 3903 3973
rect 3916 3927 3923 4034
rect 3936 3927 3943 4193
rect 3976 4147 3983 4273
rect 3996 4227 4003 4303
rect 4016 4207 4023 4253
rect 3996 4087 4003 4173
rect 4036 4167 4043 4303
rect 4096 4296 4123 4303
rect 4116 4167 4123 4296
rect 4136 4207 4143 4473
rect 4016 4067 4023 4133
rect 3996 3996 4023 4003
rect 3973 3983 3987 3993
rect 3973 3980 4003 3983
rect 3976 3976 4003 3980
rect 3896 3896 3923 3903
rect 3876 3847 3883 3893
rect 3896 3823 3903 3853
rect 3876 3816 3903 3823
rect 3816 3780 3823 3783
rect 3856 3780 3863 3783
rect 3813 3767 3827 3780
rect 3806 3753 3807 3760
rect 3853 3767 3867 3780
rect 3916 3767 3923 3896
rect 3996 3843 4003 3976
rect 4016 3947 4023 3996
rect 4036 3907 4043 4034
rect 4056 3883 4063 4053
rect 4076 4047 4083 4153
rect 4156 4067 4163 4653
rect 4176 4567 4183 4812
rect 4193 4587 4207 4593
rect 4216 4587 4223 4893
rect 4236 4827 4243 4993
rect 4267 4893 4273 4907
rect 4296 4887 4303 5273
rect 4356 5007 4363 5043
rect 4416 5007 4423 5173
rect 4496 5107 4503 5436
rect 4516 5387 4523 5553
rect 4556 5376 4563 5493
rect 4596 5387 4603 5531
rect 4636 5507 4643 5633
rect 4656 5607 4663 5653
rect 4707 5633 4713 5647
rect 4676 5596 4683 5633
rect 4776 5563 4783 5594
rect 4756 5556 4783 5563
rect 4696 5376 4703 5473
rect 4756 5347 4763 5556
rect 4796 5383 4803 5893
rect 4816 5866 4823 5973
rect 4896 5947 4903 6083
rect 4936 6047 4943 6133
rect 4973 6120 4987 6133
rect 4976 6116 4983 6120
rect 5196 6116 5203 6173
rect 5356 6116 5403 6123
rect 5096 6047 5103 6114
rect 4956 5866 4963 5933
rect 5036 5896 5043 5953
rect 5076 5907 5083 6013
rect 4876 5707 4883 5863
rect 5096 5863 5103 5993
rect 5136 5987 5143 6072
rect 5056 5856 5103 5863
rect 5116 5827 5123 5953
rect 5156 5896 5163 6033
rect 5176 6027 5183 6083
rect 5176 5927 5183 6013
rect 5336 5947 5343 6083
rect 5376 6047 5383 6073
rect 5396 6027 5403 6116
rect 5416 6087 5423 6153
rect 5476 6116 5483 6173
rect 5513 6120 5527 6133
rect 5516 6116 5523 6120
rect 5616 6116 5623 6173
rect 5653 6120 5667 6133
rect 5656 6116 5663 6120
rect 5333 5900 5347 5912
rect 5336 5896 5343 5900
rect 4876 5596 4883 5633
rect 4916 5587 4923 5613
rect 4776 5376 4803 5383
rect 4576 5336 4593 5343
rect 4676 5340 4683 5343
rect 4533 5326 4547 5332
rect 4356 4927 4363 4993
rect 4316 4856 4323 4893
rect 4340 4823 4353 4827
rect 4296 4707 4303 4823
rect 4336 4816 4353 4823
rect 4340 4813 4353 4816
rect 4376 4807 4383 4893
rect 4396 4827 4403 4973
rect 4436 4947 4443 5093
rect 4576 5047 4583 5153
rect 4407 4823 4420 4827
rect 4496 4823 4503 4993
rect 4407 4816 4423 4823
rect 4476 4816 4503 4823
rect 4407 4813 4420 4816
rect 4347 4763 4360 4767
rect 4347 4753 4363 4763
rect 4336 4707 4343 4732
rect 4193 4560 4207 4573
rect 4196 4556 4203 4560
rect 4236 4556 4243 4613
rect 4256 4307 4263 4413
rect 4073 3987 4087 3993
rect 4156 4000 4163 4003
rect 4153 3987 4167 4000
rect 4036 3876 4063 3883
rect 4036 3847 4043 3876
rect 3976 3836 4003 3843
rect 3793 3743 3807 3753
rect 3853 3747 3867 3753
rect 3793 3740 3823 3743
rect 3796 3736 3823 3740
rect 3793 3707 3807 3713
rect 3816 3687 3823 3736
rect 3936 3647 3943 3833
rect 3976 3816 3983 3836
rect 4020 3826 4040 3827
rect 4020 3823 4033 3826
rect 4016 3816 4033 3823
rect 4020 3813 4033 3816
rect 3736 3476 3763 3483
rect 3616 3387 3623 3473
rect 3536 3107 3543 3353
rect 3556 3003 3563 3333
rect 3696 3308 3703 3433
rect 3676 3296 3693 3303
rect 3556 2996 3583 3003
rect 3436 2927 3443 2994
rect 3380 2783 3393 2787
rect 3376 2776 3393 2783
rect 3380 2773 3393 2776
rect 3276 2736 3303 2743
rect 3196 2476 3203 2553
rect 3256 2407 3263 2474
rect 3016 2356 3043 2363
rect 2716 2287 2723 2313
rect 2736 2256 2743 2293
rect 2776 2256 2783 2333
rect 2793 2267 2807 2273
rect 2696 2147 2703 2213
rect 2716 2107 2723 2223
rect 2756 2220 2763 2223
rect 2753 2207 2767 2220
rect 2556 1956 2583 1963
rect 2593 1960 2607 1973
rect 2596 1956 2603 1960
rect 2656 1956 2663 2013
rect 2556 1827 2563 1956
rect 2696 1907 2703 1954
rect 2476 1816 2503 1823
rect 2376 1587 2383 1693
rect 2396 1667 2403 1703
rect 2436 1700 2443 1703
rect 2433 1687 2447 1700
rect 2496 1647 2503 1816
rect 2576 1763 2583 1793
rect 2716 1767 2723 1993
rect 2736 1967 2743 2113
rect 2776 1956 2783 2153
rect 2796 2047 2803 2213
rect 2816 2167 2823 2356
rect 2836 2187 2843 2313
rect 2856 2267 2863 2293
rect 2916 2256 2923 2313
rect 2976 2268 2983 2293
rect 2856 2143 2863 2213
rect 2896 2187 2903 2223
rect 2856 2136 2883 2143
rect 2816 1956 2823 1993
rect 2747 1923 2760 1927
rect 2747 1916 2763 1923
rect 2747 1913 2760 1916
rect 2736 1807 2743 1913
rect 2796 1863 2803 1923
rect 2856 1867 2863 2093
rect 2876 1927 2883 2136
rect 2936 1956 2943 2173
rect 2996 1967 3003 1993
rect 2956 1867 2963 1923
rect 2796 1856 2823 1863
rect 2556 1756 2583 1763
rect 2556 1736 2563 1756
rect 2516 1507 2523 1733
rect 2656 1706 2663 1753
rect 2536 1607 2543 1633
rect 2376 1436 2383 1473
rect 2507 1456 2543 1463
rect 2413 1447 2427 1453
rect 2536 1448 2543 1456
rect 2356 1307 2363 1403
rect 2393 1386 2407 1392
rect 2376 1376 2393 1383
rect 2356 1247 2363 1293
rect 2376 1223 2383 1376
rect 2436 1307 2443 1413
rect 2476 1400 2483 1403
rect 2473 1387 2487 1400
rect 2356 1216 2383 1223
rect 2296 1180 2303 1183
rect 2276 1147 2283 1173
rect 2293 1167 2307 1180
rect 2396 1107 2403 1233
rect 2453 1220 2467 1233
rect 2496 1228 2503 1293
rect 2556 1247 2563 1353
rect 2576 1267 2583 1513
rect 2596 1287 2603 1593
rect 2616 1507 2623 1703
rect 2676 1527 2683 1733
rect 2716 1647 2723 1692
rect 2756 1627 2763 1703
rect 2736 1616 2753 1623
rect 2636 1436 2643 1473
rect 2656 1367 2663 1403
rect 2696 1367 2703 1393
rect 2456 1216 2463 1220
rect 2416 1147 2423 1214
rect 2636 1216 2643 1293
rect 2676 1227 2683 1313
rect 2476 1180 2483 1183
rect 2473 1167 2487 1180
rect 2396 1096 2413 1107
rect 2400 1093 2413 1096
rect 2276 943 2283 1013
rect 2256 936 2283 943
rect 2256 916 2263 936
rect 2296 916 2303 1053
rect 2356 887 2363 933
rect 2376 927 2383 1013
rect 2396 916 2403 1053
rect 2433 920 2447 933
rect 2436 916 2443 920
rect 2276 863 2283 872
rect 2256 856 2283 863
rect 2236 667 2243 694
rect 1973 627 1987 633
rect 1756 366 1763 493
rect 1876 366 1883 413
rect 1956 396 1963 473
rect 1996 427 2003 653
rect 2036 587 2043 663
rect 2076 627 2083 663
rect 2176 507 2183 663
rect 2196 483 2203 533
rect 2176 476 2203 483
rect 2016 367 2023 473
rect 2036 307 2043 394
rect 1536 227 1543 253
rect 1556 176 1563 233
rect 1676 176 1683 233
rect 1796 227 1803 293
rect 2096 287 2103 363
rect 1816 207 1823 233
rect 1813 180 1827 193
rect 1816 176 1823 180
rect 1496 140 1503 143
rect 1493 127 1507 140
rect 1576 107 1583 132
rect 1616 107 1623 153
rect 1876 47 1883 173
rect 1940 143 1953 147
rect 1936 136 1953 143
rect 1940 133 1953 136
rect 1976 107 1983 174
rect 2007 183 2020 187
rect 2007 176 2023 183
rect 2007 173 2020 176
rect 2176 176 2183 476
rect 2236 467 2243 653
rect 2256 547 2263 856
rect 2316 827 2323 883
rect 2293 700 2307 713
rect 2296 696 2303 700
rect 2336 696 2343 733
rect 2496 696 2503 1093
rect 2556 987 2563 1212
rect 2573 1147 2587 1153
rect 2656 1147 2663 1183
rect 2696 1007 2703 1253
rect 2716 1228 2723 1553
rect 2736 1387 2743 1616
rect 2776 1587 2783 1692
rect 2796 1607 2803 1833
rect 2816 1747 2823 1856
rect 3016 1847 3023 2113
rect 3036 2007 3043 2356
rect 3056 2356 3083 2363
rect 3056 2187 3063 2356
rect 3096 2220 3103 2223
rect 3056 2087 3063 2173
rect 3076 2167 3083 2212
rect 3093 2207 3107 2220
rect 3156 2127 3163 2223
rect 3196 2207 3203 2293
rect 3216 2187 3223 2393
rect 3276 2367 3283 2693
rect 3296 2647 3303 2736
rect 3356 2707 3363 2743
rect 3416 2547 3423 2773
rect 3436 2727 3443 2853
rect 3456 2527 3463 2773
rect 3476 2607 3483 2893
rect 3496 2667 3503 2743
rect 3516 2487 3523 2713
rect 3536 2567 3543 2933
rect 3556 2747 3563 2953
rect 3576 2547 3583 2996
rect 3596 2667 3603 3033
rect 3616 2967 3623 3233
rect 3716 3147 3723 3473
rect 3736 3387 3743 3476
rect 3816 3407 3823 3483
rect 3836 3427 3843 3473
rect 3676 2827 3683 2963
rect 3716 2907 3723 3093
rect 3736 3047 3743 3373
rect 3796 3207 3803 3263
rect 3836 3167 3843 3253
rect 3856 3247 3863 3533
rect 3876 3486 3883 3593
rect 3976 3527 3983 3753
rect 3876 3247 3883 3433
rect 3916 3347 3923 3472
rect 3956 3463 3963 3472
rect 3936 3456 3963 3463
rect 3936 3308 3943 3456
rect 3996 3447 4003 3751
rect 4036 3647 4043 3773
rect 4056 3687 4063 3814
rect 4073 3767 4087 3773
rect 4156 3767 4163 3814
rect 4016 3407 4023 3533
rect 4116 3527 4123 3753
rect 4176 3727 4183 3893
rect 4196 3887 4203 4033
rect 4216 3967 4223 4053
rect 4236 4047 4243 4133
rect 4276 4087 4283 4573
rect 4356 4556 4363 4753
rect 4376 4567 4383 4733
rect 4296 4043 4303 4453
rect 4376 4427 4383 4513
rect 4396 4487 4403 4773
rect 4416 4563 4423 4793
rect 4436 4707 4443 4793
rect 4496 4767 4503 4816
rect 4433 4587 4447 4593
rect 4416 4556 4443 4563
rect 4496 4556 4503 4633
rect 4416 4367 4423 4512
rect 4493 4483 4507 4493
rect 4476 4480 4507 4483
rect 4476 4476 4503 4480
rect 4396 4306 4403 4333
rect 4416 4303 4423 4353
rect 4476 4336 4483 4476
rect 4516 4347 4523 4933
rect 4536 4467 4543 4873
rect 4596 4856 4603 5333
rect 4673 5327 4687 5340
rect 4676 5083 4683 5193
rect 4716 5107 4723 5332
rect 4776 5147 4783 5376
rect 4876 5376 4883 5513
rect 4816 5307 4823 5343
rect 4856 5323 4863 5343
rect 4836 5316 4863 5323
rect 4693 5083 4707 5093
rect 4676 5080 4707 5083
rect 4676 5076 4703 5080
rect 4696 5046 4703 5076
rect 4793 5080 4807 5093
rect 4816 5087 4823 5133
rect 4796 5076 4803 5080
rect 4636 4987 4643 5043
rect 4696 4907 4703 5032
rect 4716 4987 4723 5072
rect 4736 4967 4743 5033
rect 4776 5007 4783 5043
rect 4676 4896 4693 4903
rect 4656 4827 4663 4854
rect 4576 4783 4583 4812
rect 4616 4787 4623 4823
rect 4556 4776 4583 4783
rect 4556 4567 4563 4776
rect 4576 4556 4583 4593
rect 4616 4556 4623 4633
rect 4636 4587 4643 4633
rect 4536 4306 4543 4333
rect 4416 4296 4443 4303
rect 4287 4036 4303 4043
rect 4316 4006 4323 4073
rect 4356 4063 4363 4292
rect 4376 4127 4383 4173
rect 4396 4063 4403 4173
rect 4336 4056 4363 4063
rect 4376 4056 4403 4063
rect 4236 3856 4243 3993
rect 4256 3947 4263 3992
rect 4336 3967 4343 4056
rect 4376 4036 4383 4056
rect 4436 4048 4443 4296
rect 4556 4267 4563 4512
rect 4596 4487 4603 4523
rect 4656 4367 4663 4433
rect 4633 4340 4647 4353
rect 4676 4347 4683 4896
rect 4776 4823 4783 4953
rect 4696 4787 4703 4823
rect 4756 4816 4783 4823
rect 4696 4527 4703 4752
rect 4756 4556 4763 4793
rect 4716 4516 4743 4523
rect 4636 4336 4643 4340
rect 4336 3767 4343 3793
rect 4356 3786 4363 4033
rect 4416 3967 4423 4003
rect 4456 3967 4463 4193
rect 4376 3887 4383 3913
rect 4376 3827 4383 3873
rect 4396 3816 4403 3893
rect 4436 3816 4443 3893
rect 4476 3827 4483 4173
rect 4516 4167 4523 4253
rect 4576 4127 4583 4293
rect 4616 4267 4623 4303
rect 4660 4283 4673 4286
rect 4656 4273 4673 4283
rect 4516 4048 4523 4113
rect 4656 4048 4663 4273
rect 4696 4167 4703 4473
rect 4716 4407 4723 4516
rect 4756 4367 4763 4493
rect 4776 4427 4783 4523
rect 4816 4387 4823 5033
rect 4836 4967 4843 5316
rect 4916 5307 4923 5552
rect 4936 5487 4943 5733
rect 5116 5667 5123 5753
rect 5176 5727 5183 5863
rect 5216 5787 5223 5863
rect 5256 5807 5263 5873
rect 5316 5827 5323 5863
rect 5356 5860 5363 5863
rect 5353 5847 5367 5860
rect 5136 5596 5143 5633
rect 5176 5627 5183 5713
rect 5116 5543 5123 5563
rect 5096 5536 5123 5543
rect 5096 5376 5103 5536
rect 4976 5340 4983 5343
rect 4973 5327 4987 5340
rect 5016 5267 5023 5343
rect 5056 5227 5063 5374
rect 4893 5080 4907 5093
rect 4896 5076 4903 5080
rect 4876 4987 4883 5043
rect 4956 4927 4963 5213
rect 5116 5167 5123 5343
rect 5033 5080 5047 5093
rect 5036 5076 5043 5080
rect 5136 5083 5143 5313
rect 5156 5267 5163 5343
rect 5196 5307 5203 5633
rect 5216 5567 5223 5773
rect 5236 5596 5263 5603
rect 5316 5596 5323 5633
rect 5236 5567 5243 5596
rect 5296 5527 5303 5563
rect 5256 5376 5263 5413
rect 5296 5387 5303 5513
rect 5127 5076 5143 5083
rect 4976 5007 4983 5053
rect 5116 5047 5123 5074
rect 5256 5047 5263 5293
rect 5296 5083 5303 5333
rect 5316 5227 5323 5393
rect 5336 5387 5343 5653
rect 5356 5447 5363 5613
rect 5396 5596 5403 5853
rect 5416 5627 5423 5933
rect 5436 5667 5443 5993
rect 5496 5947 5503 6013
rect 5496 5896 5503 5933
rect 5576 5896 5583 6072
rect 5596 5947 5603 6083
rect 5696 6083 5703 6233
rect 5756 6116 5763 6173
rect 5793 6120 5807 6133
rect 5796 6116 5803 6120
rect 5936 6116 5943 6296
rect 6093 6127 6107 6133
rect 5676 6076 5703 6083
rect 5736 6080 5743 6083
rect 5476 5860 5483 5863
rect 5473 5847 5487 5860
rect 5536 5807 5543 5894
rect 5536 5703 5543 5793
rect 5596 5727 5603 5863
rect 5636 5787 5643 5863
rect 5527 5696 5543 5703
rect 5496 5567 5503 5594
rect 5353 5380 5367 5393
rect 5356 5376 5363 5380
rect 5396 5376 5403 5433
rect 5416 5407 5423 5563
rect 5456 5507 5463 5563
rect 5516 5527 5523 5693
rect 5596 5527 5603 5563
rect 5416 5307 5423 5343
rect 5276 5076 5303 5083
rect 5316 5076 5323 5153
rect 5356 5088 5363 5113
rect 5016 4947 5023 5043
rect 5216 5023 5223 5043
rect 5276 5027 5283 5076
rect 5396 5087 5403 5253
rect 5196 5020 5223 5023
rect 5196 5016 5227 5020
rect 4876 4856 4883 4913
rect 4916 4856 4963 4863
rect 4856 4807 4863 4823
rect 4956 4807 4963 4856
rect 4976 4847 4983 4873
rect 5036 4868 5043 4893
rect 5093 4860 5107 4873
rect 5096 4856 5103 4860
rect 4996 4807 5003 4854
rect 5196 4827 5203 5016
rect 5213 5007 5227 5016
rect 5236 4856 5243 4893
rect 5276 4856 5283 4933
rect 5316 4863 5323 5013
rect 5336 4987 5343 5043
rect 5376 5007 5383 5043
rect 5416 4907 5423 5213
rect 5476 5147 5483 5393
rect 5556 5376 5563 5513
rect 5536 5340 5543 5343
rect 5533 5327 5547 5340
rect 5616 5327 5623 5373
rect 5636 5347 5643 5553
rect 5656 5387 5663 5594
rect 5676 5547 5683 6076
rect 5733 6067 5747 6080
rect 5736 5896 5743 6032
rect 5876 5967 5883 6113
rect 6116 6087 6123 6153
rect 6216 6116 6223 6153
rect 6333 6120 6347 6133
rect 6336 6116 6343 6120
rect 5896 6007 5903 6083
rect 6036 6047 6043 6083
rect 6076 6027 6083 6072
rect 6136 6043 6143 6114
rect 6153 6067 6167 6073
rect 6256 6083 6263 6114
rect 6256 6076 6283 6083
rect 6127 6036 6143 6043
rect 5876 5903 5883 5953
rect 5876 5896 5903 5903
rect 5956 5896 5963 6013
rect 5696 5607 5703 5753
rect 5716 5707 5723 5863
rect 5756 5787 5763 5863
rect 5796 5747 5803 5894
rect 5716 5596 5723 5633
rect 5676 5427 5683 5453
rect 5676 5376 5683 5413
rect 5756 5307 5763 5533
rect 5776 5447 5783 5563
rect 5816 5507 5823 5633
rect 5856 5608 5863 5863
rect 5836 5596 5853 5603
rect 5836 5566 5843 5596
rect 5896 5596 5903 5896
rect 5936 5767 5943 5863
rect 5976 5747 5983 5852
rect 6016 5827 6023 6013
rect 6073 5900 6087 5913
rect 6076 5896 6083 5900
rect 6116 5896 6123 6033
rect 6216 5896 6223 5973
rect 6096 5827 6103 5863
rect 5916 5527 5923 5563
rect 5956 5507 5963 5553
rect 5976 5547 5983 5633
rect 6033 5608 6047 5613
rect 6076 5596 6083 5633
rect 6016 5560 6023 5563
rect 5896 5367 5903 5433
rect 5956 5376 5963 5493
rect 5996 5467 6003 5553
rect 6013 5547 6027 5560
rect 6033 5523 6047 5533
rect 6056 5527 6063 5563
rect 6016 5520 6047 5523
rect 6016 5516 6043 5520
rect 5856 5340 5863 5343
rect 5853 5327 5867 5340
rect 5936 5327 5943 5343
rect 5976 5323 5983 5332
rect 6016 5327 6023 5516
rect 6116 5487 6123 5833
rect 6136 5547 6143 5793
rect 6156 5607 6163 5893
rect 6196 5860 6203 5863
rect 6193 5847 6207 5860
rect 6236 5807 6243 5863
rect 6173 5600 6187 5613
rect 6176 5596 6183 5600
rect 6216 5596 6223 5633
rect 6256 5607 6263 5653
rect 6156 5523 6163 5553
rect 6156 5516 6183 5523
rect 6136 5487 6143 5512
rect 6036 5327 6043 5473
rect 6136 5376 6143 5473
rect 6156 5387 6163 5493
rect 5956 5316 5983 5323
rect 5696 5187 5703 5293
rect 5436 5043 5443 5093
rect 5493 5080 5507 5093
rect 5496 5076 5503 5080
rect 5436 5036 5463 5043
rect 5316 4856 5343 4863
rect 5076 4820 5083 4823
rect 5073 4807 5087 4820
rect 4856 4747 4863 4793
rect 4876 4556 4883 4613
rect 4916 4556 4923 4793
rect 5073 4787 5087 4793
rect 5256 4787 5263 4812
rect 5296 4787 5303 4823
rect 4956 4568 4963 4713
rect 5036 4627 5043 4673
rect 5016 4616 5033 4623
rect 4836 4367 4843 4533
rect 4896 4487 4903 4523
rect 4936 4503 4943 4523
rect 4936 4496 4963 4503
rect 4716 4247 4723 4353
rect 4773 4340 4787 4353
rect 4876 4348 4883 4433
rect 4776 4336 4783 4340
rect 4756 4187 4763 4292
rect 4796 4267 4803 4303
rect 4836 4300 4843 4303
rect 4833 4287 4847 4300
rect 4816 4247 4823 4273
rect 4696 4048 4703 4153
rect 4756 4067 4763 4173
rect 4836 4087 4843 4273
rect 4856 4247 4863 4273
rect 4876 4207 4883 4334
rect 4896 4187 4903 4353
rect 4576 4036 4603 4043
rect 4496 3786 4503 3853
rect 4416 3780 4423 3783
rect 4153 3520 4167 3533
rect 4156 3516 4163 3520
rect 4196 3516 4203 3613
rect 4276 3516 4283 3553
rect 4316 3516 4323 3633
rect 4356 3627 4363 3772
rect 4413 3767 4427 3780
rect 4056 3407 4063 3483
rect 3980 3303 3993 3307
rect 3976 3296 3993 3303
rect 3980 3294 3993 3296
rect 4027 3293 4033 3307
rect 4053 3300 4067 3313
rect 4056 3296 4063 3300
rect 4096 3296 4103 3413
rect 4116 3327 4123 3513
rect 4356 3487 4363 3514
rect 4176 3427 4183 3483
rect 4333 3300 4347 3313
rect 4336 3296 4343 3300
rect 3956 3260 3963 3263
rect 3953 3247 3967 3260
rect 4016 3247 4023 3272
rect 3796 2996 3803 3133
rect 3836 3008 3843 3113
rect 3736 2867 3743 2973
rect 3776 2907 3783 2963
rect 3776 2787 3783 2893
rect 3856 2847 3863 3093
rect 3876 2963 3883 3153
rect 3936 3047 3943 3213
rect 4016 3003 4023 3033
rect 4007 2996 4023 3003
rect 3876 2956 3903 2963
rect 3616 2647 3623 2743
rect 3356 2440 3363 2443
rect 3353 2427 3367 2440
rect 3236 2287 3243 2333
rect 3276 2256 3283 2293
rect 3316 2256 3323 2313
rect 3336 2267 3343 2353
rect 3116 2007 3123 2033
rect 3073 1987 3087 1993
rect 3073 1960 3087 1973
rect 3076 1956 3083 1960
rect 3116 1956 3123 1993
rect 3156 1967 3163 2013
rect 3176 1926 3183 2033
rect 3216 1956 3223 1993
rect 3253 1960 3267 1973
rect 3256 1956 3263 1960
rect 2896 1736 2903 1773
rect 2816 1667 2823 1712
rect 2836 1627 2843 1693
rect 2776 1436 2783 1473
rect 2816 1436 2823 1533
rect 2876 1406 2883 1593
rect 2956 1487 2963 1773
rect 2856 1367 2863 1393
rect 2896 1367 2903 1473
rect 2976 1467 2983 1813
rect 3056 1807 3063 1923
rect 3096 1887 3103 1923
rect 3236 1887 3243 1923
rect 3056 1743 3063 1793
rect 3047 1736 3063 1743
rect 3076 1607 3083 1833
rect 3113 1740 3127 1753
rect 3116 1736 3123 1740
rect 3176 1667 3183 1692
rect 3216 1607 3223 1773
rect 3276 1767 3283 1923
rect 3316 1787 3323 1953
rect 3336 1883 3343 2073
rect 3356 2047 3363 2413
rect 3436 2407 3443 2443
rect 3456 2287 3463 2353
rect 3476 2347 3483 2443
rect 3536 2427 3543 2473
rect 3556 2407 3563 2473
rect 3616 2407 3623 2443
rect 3420 2263 3433 2267
rect 3416 2256 3433 2263
rect 3420 2253 3433 2256
rect 3456 2223 3463 2273
rect 3476 2267 3483 2333
rect 3513 2260 3527 2273
rect 3516 2256 3523 2260
rect 3456 2216 3503 2223
rect 3436 2187 3443 2213
rect 3556 2207 3563 2393
rect 3636 2383 3643 2733
rect 3676 2587 3683 2743
rect 3616 2376 3643 2383
rect 3616 2256 3623 2376
rect 3656 2267 3663 2533
rect 3676 2307 3683 2573
rect 3716 2476 3723 2553
rect 3756 2267 3763 2713
rect 3796 2367 3803 2793
rect 3856 2776 3863 2833
rect 3916 2727 3923 2893
rect 3836 2547 3843 2633
rect 3836 2476 3843 2533
rect 3936 2487 3943 2923
rect 4016 2907 4023 2953
rect 4036 2807 4043 3252
rect 4073 3247 4087 3252
rect 4116 3127 4123 3263
rect 4076 3007 4083 3113
rect 4136 3008 4143 3252
rect 4156 3227 4163 3263
rect 4376 3227 4383 3573
rect 4396 3267 4403 3733
rect 4496 3303 4503 3713
rect 4516 3486 4523 3893
rect 4556 3887 4563 3992
rect 4596 3987 4603 4036
rect 4576 3816 4583 3853
rect 4616 3827 4623 4034
rect 4793 4040 4807 4053
rect 4833 4056 4875 4064
rect 4833 4048 4847 4056
rect 4916 4048 4923 4373
rect 4956 4348 4963 4496
rect 4976 4387 4983 4513
rect 4996 4423 5003 4593
rect 5016 4567 5023 4616
rect 5036 4556 5043 4613
rect 5116 4587 5123 4613
rect 5073 4560 5087 4573
rect 5076 4556 5083 4560
rect 5016 4483 5023 4513
rect 5016 4476 5043 4483
rect 4996 4416 5023 4423
rect 4996 4300 5003 4303
rect 4936 4227 4943 4292
rect 4993 4287 5007 4300
rect 4796 4036 4803 4040
rect 4956 4036 4963 4113
rect 5016 4087 5023 4416
rect 5036 4287 5043 4476
rect 5056 4427 5063 4523
rect 5116 4487 5123 4573
rect 5156 4556 5163 4673
rect 5196 4556 5203 4673
rect 5236 4556 5243 4593
rect 5056 4107 5063 4373
rect 5116 4336 5123 4452
rect 5156 4347 5163 4493
rect 5176 4348 5183 4523
rect 5216 4487 5223 4523
rect 5120 4285 5140 4287
rect 5120 4282 5133 4285
rect 5116 4273 5133 4282
rect 5116 4067 5123 4273
rect 5136 4207 5143 4233
rect 4993 4048 5007 4053
rect 4596 3707 4603 3772
rect 4616 3747 4623 3773
rect 4556 3627 4563 3673
rect 4576 3516 4583 3653
rect 4616 3627 4623 3653
rect 4613 3543 4627 3553
rect 4636 3543 4643 3973
rect 4676 3847 4683 4003
rect 4756 3987 4763 4032
rect 4776 3907 4783 3993
rect 4856 3883 4863 4003
rect 4976 3927 4983 4003
rect 4856 3876 4883 3883
rect 4676 3816 4683 3833
rect 4716 3828 4723 3853
rect 4696 3780 4703 3783
rect 4693 3767 4707 3780
rect 4756 3567 4763 3853
rect 4813 3820 4827 3833
rect 4816 3816 4823 3820
rect 4856 3816 4863 3853
rect 4876 3847 4883 3876
rect 4896 3816 4903 3873
rect 4987 3853 4993 3867
rect 4776 3786 4783 3813
rect 4936 3767 4943 3853
rect 4956 3786 4963 3833
rect 4993 3820 5007 3832
rect 4996 3816 5003 3820
rect 5036 3816 5043 3853
rect 5056 3827 5063 4053
rect 5136 4036 5143 4093
rect 5156 4047 5163 4293
rect 5176 4267 5183 4334
rect 5196 4083 5203 4413
rect 5256 4336 5263 4493
rect 5276 4367 5283 4573
rect 5296 4467 5303 4773
rect 5316 4563 5323 4713
rect 5336 4587 5343 4856
rect 5356 4587 5363 4893
rect 5456 4787 5463 5036
rect 5576 5007 5583 5074
rect 5376 4568 5383 4633
rect 5316 4556 5343 4563
rect 5396 4567 5403 4673
rect 5476 4587 5483 4953
rect 5496 4867 5503 4993
rect 5596 4967 5603 5133
rect 5633 5080 5647 5093
rect 5636 5076 5643 5080
rect 5736 5047 5743 5113
rect 5656 5007 5663 5043
rect 5756 5036 5783 5043
rect 5536 4856 5543 4913
rect 5696 4856 5703 4973
rect 5516 4667 5523 4823
rect 5616 4807 5623 4854
rect 5356 4367 5363 4523
rect 5236 4300 5243 4303
rect 5233 4287 5247 4300
rect 5233 4247 5247 4252
rect 5176 4076 5203 4083
rect 5176 4027 5183 4076
rect 5236 4067 5243 4233
rect 5076 3667 5083 3993
rect 4613 3540 4643 3543
rect 4616 3536 4643 3540
rect 4616 3516 4623 3536
rect 4476 3296 4503 3303
rect 4233 3008 4247 3014
rect 4056 2923 4063 2994
rect 4073 2947 4087 2953
rect 4056 2916 4083 2923
rect 3973 2780 3987 2793
rect 3976 2776 3983 2780
rect 3996 2740 4003 2743
rect 3993 2727 4007 2740
rect 4076 2727 4083 2916
rect 4176 2883 4183 2994
rect 4316 2963 4323 3153
rect 4176 2876 4203 2883
rect 4096 2787 4103 2833
rect 4133 2780 4147 2793
rect 4136 2776 4143 2780
rect 4116 2727 4123 2743
rect 4196 2727 4203 2876
rect 4216 2867 4223 2963
rect 4256 2927 4263 2963
rect 4296 2956 4323 2963
rect 3976 2488 3983 2513
rect 3776 2226 3783 2313
rect 3376 1968 3383 2173
rect 3396 1887 3403 1923
rect 3336 1876 3363 1883
rect 3276 1736 3283 1753
rect 3236 1667 3243 1733
rect 3336 1707 3343 1833
rect 3356 1807 3363 1876
rect 3436 1787 3443 1923
rect 3296 1647 3303 1703
rect 2913 1387 2927 1392
rect 2896 1327 2903 1353
rect 2936 1303 2943 1403
rect 2936 1296 2963 1303
rect 2816 1228 2823 1273
rect 2876 1216 2883 1253
rect 2716 1027 2723 1214
rect 2776 1147 2783 1183
rect 2553 920 2567 933
rect 2556 916 2563 920
rect 2596 916 2603 993
rect 2516 827 2523 913
rect 2533 863 2547 873
rect 2533 860 2563 863
rect 2536 856 2563 860
rect 2536 707 2543 833
rect 2556 823 2563 856
rect 2576 847 2583 883
rect 2616 880 2623 883
rect 2613 867 2627 880
rect 2636 827 2643 853
rect 2556 816 2593 823
rect 2656 767 2663 973
rect 2696 916 2703 993
rect 2736 928 2743 953
rect 2716 847 2723 883
rect 2736 827 2743 853
rect 2756 807 2763 883
rect 2236 360 2243 363
rect 2233 347 2247 360
rect 2276 347 2283 433
rect 2336 396 2343 513
rect 2376 487 2383 694
rect 2436 527 2443 663
rect 2376 396 2383 473
rect 2476 447 2483 663
rect 2556 543 2563 753
rect 2616 696 2623 733
rect 2536 536 2563 543
rect 2233 327 2247 333
rect 2236 167 2243 233
rect 2336 176 2343 213
rect 2156 87 2163 143
rect 2196 47 2203 143
rect 2216 27 2223 133
rect 2236 127 2243 153
rect 2256 87 2263 173
rect 2396 146 2403 273
rect 2316 140 2323 143
rect 2356 140 2363 143
rect 2313 127 2327 140
rect 2353 127 2367 140
rect 2393 127 2407 132
rect 2536 47 2543 536
rect 2556 407 2563 473
rect 2556 327 2563 393
rect 2576 366 2583 693
rect 2636 627 2643 663
rect 2716 627 2723 753
rect 2756 696 2763 733
rect 2796 708 2803 1093
rect 2816 947 2823 1214
rect 2900 1183 2913 1187
rect 2856 1107 2863 1183
rect 2896 1173 2913 1183
rect 2896 927 2903 1173
rect 2936 923 2943 1273
rect 2956 1227 2963 1296
rect 3036 1267 3043 1493
rect 3216 1436 3223 1533
rect 3276 1406 3283 1453
rect 3416 1443 3423 1593
rect 3436 1527 3443 1733
rect 3456 1706 3463 1813
rect 3476 1747 3483 2173
rect 3496 1767 3503 2193
rect 3596 2187 3603 2223
rect 3616 2167 3623 2193
rect 3636 2087 3643 2212
rect 3676 2127 3683 2223
rect 3796 2127 3803 2293
rect 3876 2127 3883 2213
rect 3556 1987 3563 2013
rect 3556 1973 3573 1987
rect 3556 1956 3563 1973
rect 3616 1947 3623 2033
rect 3676 2027 3683 2113
rect 3673 1960 3687 1973
rect 3676 1956 3683 1960
rect 3816 1927 3823 1954
rect 3647 1923 3660 1927
rect 3647 1916 3663 1923
rect 3647 1913 3660 1916
rect 3536 1887 3543 1912
rect 3756 1887 3763 1923
rect 3836 1907 3843 2113
rect 3896 2107 3903 2473
rect 4036 2447 4043 2711
rect 4116 2507 4123 2713
rect 4236 2587 4243 2873
rect 4296 2816 4303 2956
rect 4336 2887 4343 3113
rect 4356 3047 4363 3173
rect 4373 3000 4387 3013
rect 4376 2996 4383 3000
rect 4416 2996 4423 3293
rect 4447 3256 4463 3263
rect 4436 3087 4443 3253
rect 4456 2996 4463 3113
rect 4516 3087 4523 3333
rect 4536 3266 4543 3373
rect 4556 3307 4563 3453
rect 4596 3347 4603 3483
rect 4636 3480 4643 3483
rect 4633 3467 4647 3480
rect 4636 3336 4643 3373
rect 4556 2966 4563 3293
rect 4436 2927 4443 2953
rect 4576 2847 4583 3073
rect 4696 3008 4703 3513
rect 4736 3303 4743 3483
rect 4716 3296 4743 3303
rect 4776 3296 4783 3333
rect 4796 3327 4803 3553
rect 4956 3487 4963 3553
rect 4987 3516 5003 3523
rect 4816 3296 4823 3433
rect 4976 3427 4983 3514
rect 4836 3307 4843 3373
rect 4716 3107 4723 3296
rect 4756 3187 4763 3263
rect 4796 3227 4803 3263
rect 4856 3207 4863 3333
rect 4876 3307 4883 3353
rect 4913 3300 4927 3313
rect 4916 3296 4923 3300
rect 4956 3296 4963 3353
rect 5096 3328 5103 3913
rect 5116 3887 5123 4003
rect 5196 3907 5203 4053
rect 5233 4040 5247 4053
rect 5236 4036 5243 4040
rect 5276 4036 5283 4073
rect 5156 3847 5163 3873
rect 5136 3516 5143 3553
rect 5236 3543 5243 3793
rect 5216 3536 5243 3543
rect 4986 3313 4987 3320
rect 4973 3307 4987 3313
rect 4856 2963 4863 3073
rect 4876 3067 4883 3253
rect 4896 3207 4903 3263
rect 4936 3187 4943 3263
rect 4956 3087 4963 3233
rect 4836 2956 4863 2963
rect 4376 2727 4383 2773
rect 4093 2480 4107 2493
rect 4096 2476 4103 2480
rect 4296 2476 4303 2573
rect 4353 2480 4367 2493
rect 4376 2487 4383 2713
rect 4396 2707 4403 2813
rect 4436 2740 4443 2743
rect 4433 2727 4447 2740
rect 4476 2707 4483 2743
rect 4356 2476 4363 2480
rect 3916 2187 3923 2273
rect 3976 2256 3983 2313
rect 4013 2260 4027 2273
rect 4036 2267 4043 2433
rect 4176 2443 4183 2474
rect 4116 2387 4123 2443
rect 4176 2436 4203 2443
rect 4016 2256 4023 2260
rect 3916 2087 3923 2113
rect 3936 2067 3943 2213
rect 3956 2203 3963 2223
rect 3956 2196 3983 2203
rect 3976 2127 3983 2196
rect 3996 2167 4003 2223
rect 3956 2047 3963 2113
rect 3873 1960 3887 1973
rect 3876 1956 3883 1960
rect 3936 1956 3943 1993
rect 3516 1736 3523 1833
rect 3976 1827 3983 1953
rect 3996 1847 4003 1993
rect 4036 1968 4043 2173
rect 4056 2167 4063 2273
rect 4096 2256 4103 2333
rect 4173 2267 4187 2273
rect 4116 2220 4123 2223
rect 4113 2207 4127 2220
rect 4196 2207 4203 2436
rect 4376 2347 4383 2433
rect 4216 2226 4223 2333
rect 4336 2256 4343 2333
rect 4236 2187 4243 2213
rect 4296 2207 4303 2223
rect 4116 1947 4123 2113
rect 4216 1968 4223 2153
rect 4296 2003 4303 2193
rect 4396 2167 4403 2533
rect 4416 2387 4423 2493
rect 4516 2488 4523 2833
rect 4596 2740 4603 2743
rect 4593 2727 4607 2740
rect 4636 2727 4643 2853
rect 4716 2776 4723 2853
rect 4796 2827 4803 2923
rect 4876 2867 4883 3032
rect 4956 2996 4963 3073
rect 4853 2780 4867 2793
rect 4856 2776 4863 2780
rect 4656 2707 4663 2773
rect 4673 2743 4687 2753
rect 4916 2743 4923 2833
rect 4996 2807 5003 3313
rect 5053 3300 5067 3313
rect 5136 3307 5143 3433
rect 5216 3347 5223 3536
rect 5256 3523 5263 3853
rect 5276 3783 5283 3933
rect 5316 3867 5323 4353
rect 5376 4336 5383 4413
rect 5336 3887 5343 4053
rect 5396 4036 5403 4153
rect 5416 4067 5423 4573
rect 5436 4347 5443 4573
rect 5467 4523 5480 4527
rect 5467 4513 5483 4523
rect 5476 4427 5483 4513
rect 5536 4507 5543 4553
rect 5453 4340 5467 4353
rect 5456 4336 5463 4340
rect 5536 4347 5543 4472
rect 5436 4043 5443 4293
rect 5476 4227 5483 4303
rect 5496 4043 5503 4273
rect 5536 4227 5543 4293
rect 5556 4283 5563 4791
rect 5676 4567 5683 4812
rect 5716 4747 5723 4823
rect 5756 4807 5763 5036
rect 5776 4867 5783 5013
rect 5836 4867 5843 5293
rect 5856 5087 5863 5233
rect 5893 5088 5907 5094
rect 5876 4947 5883 5043
rect 5776 4707 5783 4813
rect 5796 4747 5803 4823
rect 5716 4647 5723 4673
rect 5813 4667 5827 4673
rect 5836 4667 5843 4813
rect 5856 4807 5863 4913
rect 5896 4887 5903 5013
rect 5916 4967 5923 5033
rect 5936 5027 5943 5313
rect 5956 5087 5963 5316
rect 6013 5080 6027 5093
rect 6016 5076 6023 5080
rect 5976 4963 5983 5013
rect 5996 4983 6003 5043
rect 6013 5007 6027 5013
rect 5996 4976 6023 4983
rect 5976 4956 6003 4963
rect 5916 4856 5923 4893
rect 5960 4863 5973 4867
rect 5956 4856 5973 4863
rect 5960 4854 5973 4856
rect 5960 4853 5964 4854
rect 5853 4647 5867 4653
rect 5660 4523 5673 4526
rect 5616 4520 5623 4523
rect 5613 4507 5627 4520
rect 5656 4516 5673 4523
rect 5660 4513 5673 4516
rect 5696 4507 5703 4554
rect 5836 4523 5843 4593
rect 5876 4567 5883 4813
rect 5996 4823 6003 4956
rect 6016 4907 6023 4976
rect 6016 4867 6023 4893
rect 6056 4887 6063 5033
rect 6076 5023 6083 5311
rect 6096 5043 6103 5313
rect 6116 5247 6123 5343
rect 6176 5147 6183 5516
rect 6196 5487 6203 5563
rect 6196 5267 6203 5393
rect 6216 5387 6223 5533
rect 6236 5487 6243 5563
rect 6236 5376 6243 5433
rect 6256 5407 6263 5553
rect 6276 5527 6283 6076
rect 6296 5607 6303 6053
rect 6316 5907 6323 6083
rect 6376 6067 6383 6133
rect 6336 5667 6343 5863
rect 6376 5607 6383 5633
rect 6296 5447 6303 5553
rect 6336 5547 6343 5563
rect 6336 5536 6353 5547
rect 6340 5533 6353 5536
rect 6116 5087 6123 5133
rect 6193 5107 6207 5113
rect 6133 5080 6147 5093
rect 6136 5076 6143 5080
rect 6216 5083 6223 5333
rect 6216 5076 6243 5083
rect 6096 5036 6123 5043
rect 6076 5016 6103 5023
rect 6096 4963 6103 5016
rect 6116 4983 6123 5036
rect 6156 5023 6163 5043
rect 6136 5020 6163 5023
rect 6133 5016 6163 5020
rect 6133 5007 6147 5016
rect 6213 5023 6227 5033
rect 6173 5003 6187 5013
rect 6156 5000 6187 5003
rect 6196 5020 6227 5023
rect 6196 5016 6223 5020
rect 6156 4996 6183 5000
rect 6116 4976 6143 4983
rect 6096 4956 6123 4963
rect 6073 4943 6087 4953
rect 6073 4940 6103 4943
rect 6076 4936 6103 4940
rect 6047 4876 6063 4887
rect 6047 4874 6060 4876
rect 6096 4856 6103 4936
rect 6116 4867 6123 4956
rect 5936 4820 5943 4823
rect 5933 4807 5947 4820
rect 5976 4816 6003 4823
rect 5936 4767 5943 4793
rect 5916 4587 5923 4673
rect 5936 4567 5943 4693
rect 5796 4516 5843 4523
rect 5756 4503 5763 4512
rect 5856 4507 5863 4553
rect 5756 4496 5793 4503
rect 5836 4467 5843 4493
rect 5576 4307 5583 4413
rect 5556 4276 5573 4283
rect 5576 4063 5583 4272
rect 5596 4247 5603 4453
rect 5616 4267 5623 4373
rect 5673 4340 5687 4353
rect 5733 4340 5747 4353
rect 5676 4336 5683 4340
rect 5736 4336 5743 4340
rect 5636 4300 5643 4303
rect 5633 4287 5647 4300
rect 5616 4187 5623 4213
rect 5556 4056 5583 4063
rect 5436 4036 5463 4043
rect 5456 3887 5463 4036
rect 5476 4036 5503 4043
rect 5356 3816 5363 3853
rect 5276 3776 5303 3783
rect 5236 3516 5263 3523
rect 5296 3516 5303 3776
rect 5236 3367 5243 3516
rect 5336 3487 5343 3693
rect 5396 3528 5403 3873
rect 5416 3783 5423 3853
rect 5476 3843 5483 4036
rect 5556 4036 5563 4056
rect 5596 4047 5603 4153
rect 5496 3867 5503 3993
rect 5456 3836 5483 3843
rect 5456 3828 5463 3836
rect 5416 3776 5443 3783
rect 5496 3780 5503 3783
rect 5493 3767 5507 3780
rect 5436 3516 5443 3553
rect 5356 3367 5363 3513
rect 5056 3296 5063 3300
rect 5016 3027 5023 3293
rect 5036 3207 5043 3253
rect 5076 3187 5083 3263
rect 5116 3260 5123 3263
rect 5113 3247 5127 3260
rect 5156 3247 5163 3333
rect 5213 3300 5227 3312
rect 5253 3300 5267 3313
rect 5216 3296 5223 3300
rect 5256 3296 5263 3300
rect 5176 3187 5183 3293
rect 5236 3207 5243 3263
rect 4673 2740 4703 2743
rect 4676 2736 4703 2740
rect 4756 2687 4763 2743
rect 4436 2216 4463 2223
rect 4436 2187 4443 2216
rect 4276 1996 4303 2003
rect 3487 1653 3493 1667
rect 3416 1436 3443 1443
rect 3473 1440 3487 1453
rect 3476 1436 3483 1440
rect 3096 1367 3103 1403
rect 3196 1400 3203 1403
rect 3193 1387 3207 1400
rect 3176 1376 3193 1383
rect 3036 1187 3043 1214
rect 3096 1107 3103 1183
rect 3156 1147 3163 1214
rect 3176 947 3183 1376
rect 3256 1216 3263 1253
rect 3316 1183 3323 1392
rect 3376 1216 3383 1433
rect 3433 1247 3447 1253
rect 3456 1247 3463 1403
rect 3516 1387 3523 1673
rect 3533 1667 3547 1671
rect 3576 1647 3583 1692
rect 3616 1687 3623 1733
rect 3656 1700 3663 1703
rect 3653 1687 3667 1700
rect 3696 1667 3703 1703
rect 3536 1406 3543 1453
rect 3556 1436 3563 1473
rect 3416 1216 3463 1223
rect 3276 1176 3323 1183
rect 3356 1107 3363 1183
rect 3396 1087 3403 1183
rect 2916 916 2943 923
rect 2953 920 2967 933
rect 2993 920 3007 933
rect 2956 916 2963 920
rect 2996 916 3003 920
rect 2916 886 2923 916
rect 2776 660 2783 663
rect 2773 647 2787 660
rect 2836 627 2843 853
rect 2876 723 2883 793
rect 2896 767 2903 873
rect 2916 856 2963 863
rect 2916 827 2923 856
rect 2876 716 2913 723
rect 2936 696 2943 833
rect 2956 827 2963 856
rect 2976 847 2983 883
rect 3036 867 3043 933
rect 3056 847 3063 914
rect 3096 827 3103 883
rect 2976 666 2983 753
rect 2876 660 2883 663
rect 2873 647 2887 660
rect 3116 663 3123 853
rect 3136 827 3143 883
rect 3176 880 3183 883
rect 3173 867 3187 880
rect 3216 827 3223 953
rect 3236 727 3243 933
rect 3153 700 3167 713
rect 3156 696 3163 700
rect 3036 627 3043 663
rect 3076 656 3123 663
rect 2596 396 2623 403
rect 2596 267 2603 396
rect 2776 366 2783 433
rect 2836 396 2843 473
rect 2876 408 2883 612
rect 2656 327 2663 363
rect 2716 360 2723 363
rect 2713 347 2727 360
rect 2596 227 2603 253
rect 2916 247 2923 453
rect 2956 267 2963 363
rect 2556 147 2563 173
rect 2576 136 2603 143
rect 2576 27 2583 136
rect 2716 87 2723 213
rect 2820 203 2833 207
rect 2816 193 2833 203
rect 2736 107 2743 174
rect 2756 147 2763 193
rect 2816 176 2823 193
rect 2856 187 2863 233
rect 2876 146 2883 193
rect 2913 180 2927 193
rect 2916 176 2923 180
rect 2956 176 2963 232
rect 2996 187 3003 213
rect 3016 207 3023 533
rect 3096 507 3103 656
rect 3216 660 3223 663
rect 3213 647 3227 660
rect 3156 547 3163 593
rect 3096 467 3103 493
rect 3036 367 3043 413
rect 3113 400 3127 413
rect 3116 396 3123 400
rect 3156 396 3163 533
rect 3236 403 3243 653
rect 3216 396 3243 403
rect 3076 207 3083 233
rect 3096 183 3103 363
rect 3256 327 3263 633
rect 3096 176 3123 183
rect 2796 107 2803 143
rect 3116 107 3123 176
rect 3136 147 3143 213
rect 3193 188 3207 194
rect 3276 183 3283 713
rect 3316 567 3323 663
rect 3356 660 3363 663
rect 3353 647 3367 660
rect 3256 176 3283 183
rect 3236 147 3243 173
rect 3107 76 3133 83
rect 3256 63 3263 176
rect 3376 146 3383 433
rect 3396 287 3403 993
rect 3436 983 3443 1173
rect 3456 1167 3463 1216
rect 3476 1007 3483 1373
rect 3636 1247 3643 1513
rect 3676 1367 3683 1473
rect 3716 1448 3723 1693
rect 3736 1467 3743 1773
rect 3776 1736 3783 1793
rect 3796 1507 3803 1692
rect 3747 1456 3763 1463
rect 3756 1436 3763 1456
rect 3796 1367 3803 1434
rect 3676 1287 3683 1353
rect 3856 1287 3863 1403
rect 3916 1247 3923 1813
rect 3956 1700 3963 1703
rect 3953 1687 3967 1700
rect 4056 1667 4063 1734
rect 4076 1706 4083 1833
rect 4096 1743 4103 1913
rect 4136 1907 4143 1953
rect 4256 1907 4263 1954
rect 4136 1827 4143 1893
rect 4276 1807 4283 1996
rect 4336 1956 4343 2033
rect 4436 1983 4443 2093
rect 4516 2067 4523 2223
rect 4516 2007 4523 2053
rect 4436 1976 4463 1983
rect 4456 1956 4463 1976
rect 4536 1927 4543 1954
rect 4296 1916 4323 1923
rect 4296 1847 4303 1916
rect 4096 1736 4113 1743
rect 4296 1743 4303 1833
rect 4156 1736 4203 1743
rect 4276 1736 4303 1743
rect 4016 1448 4023 1653
rect 4096 1448 4103 1653
rect 4196 1647 4203 1736
rect 4316 1667 4323 1893
rect 4356 1747 4363 1923
rect 4436 1920 4443 1923
rect 4433 1907 4447 1920
rect 4476 1867 4483 1923
rect 4376 1736 4383 1793
rect 4556 1787 4563 2593
rect 4836 2488 4843 2743
rect 4896 2736 4923 2743
rect 4916 2547 4923 2736
rect 4956 2587 4963 2793
rect 5016 2776 5023 2992
rect 5076 2947 5083 2963
rect 5076 2936 5093 2947
rect 5080 2933 5093 2936
rect 5136 2847 5143 3173
rect 5156 3036 5223 3043
rect 5156 3007 5163 3036
rect 5216 3023 5223 3036
rect 5216 3016 5243 3023
rect 5193 3000 5207 3013
rect 5196 2996 5203 3000
rect 5236 2996 5243 3016
rect 5276 2963 5283 2994
rect 5176 2803 5183 2952
rect 5176 2796 5203 2803
rect 5196 2776 5203 2796
rect 5216 2787 5223 2963
rect 5256 2956 5283 2963
rect 4996 2707 5003 2743
rect 5036 2687 5043 2743
rect 4956 2476 4963 2533
rect 4716 2387 4723 2474
rect 5016 2446 5023 2573
rect 5096 2547 5103 2773
rect 5136 2687 5143 2743
rect 5196 2483 5203 2533
rect 5176 2476 5203 2483
rect 4656 2256 4663 2373
rect 4776 2226 4783 2443
rect 5036 2436 5083 2443
rect 5036 2407 5043 2436
rect 4636 2127 4643 2223
rect 4596 1987 4603 2113
rect 4676 2007 4683 2212
rect 4896 2127 4903 2223
rect 4593 1960 4607 1973
rect 4596 1956 4603 1960
rect 4736 1956 4743 2053
rect 4936 1967 4943 2153
rect 4956 2127 4963 2223
rect 5016 2216 5043 2223
rect 5036 2167 5043 2216
rect 4256 1507 4263 1633
rect 4436 1547 4443 1703
rect 4256 1443 4263 1493
rect 4236 1436 4263 1443
rect 3533 1220 3547 1233
rect 3536 1216 3543 1220
rect 3636 1186 3643 1212
rect 3516 1180 3523 1183
rect 3513 1167 3527 1180
rect 3556 1147 3563 1183
rect 3596 1176 3623 1183
rect 3416 976 3443 983
rect 3416 707 3423 976
rect 3436 923 3443 953
rect 3436 916 3463 923
rect 3516 916 3523 1013
rect 3576 827 3583 1153
rect 3616 1087 3623 1176
rect 3836 1176 3863 1183
rect 3616 923 3623 1073
rect 3676 1047 3683 1172
rect 3836 1147 3843 1176
rect 3916 1067 3923 1183
rect 3956 1127 3963 1433
rect 3976 1400 3983 1403
rect 3973 1387 3987 1400
rect 3596 916 3623 923
rect 3596 867 3603 916
rect 3676 883 3683 993
rect 3756 916 3763 1033
rect 3836 1027 3843 1053
rect 3976 1027 3983 1233
rect 3996 1186 4003 1273
rect 4036 1247 4043 1433
rect 4136 1367 4143 1403
rect 4036 1216 4043 1233
rect 4096 1147 4103 1183
rect 4136 1107 4143 1183
rect 4216 1107 4223 1153
rect 4136 1067 4143 1093
rect 3836 916 3843 1013
rect 3656 876 3683 883
rect 3596 727 3603 853
rect 3493 700 3507 713
rect 3496 696 3503 700
rect 3416 627 3423 653
rect 3476 627 3483 663
rect 3536 607 3543 663
rect 3516 596 3533 603
rect 3436 408 3443 473
rect 3476 396 3483 433
rect 3516 396 3523 596
rect 3636 523 3643 813
rect 3696 807 3703 914
rect 3736 880 3743 883
rect 3733 867 3747 880
rect 3747 856 3763 863
rect 3656 647 3663 694
rect 3756 666 3763 856
rect 3856 696 3863 793
rect 3916 663 3923 713
rect 3876 656 3923 663
rect 3756 567 3763 652
rect 3616 516 3643 523
rect 3456 327 3463 363
rect 3396 143 3403 193
rect 3516 146 3523 173
rect 3396 136 3443 143
rect 3196 56 3263 63
rect 1396 -24 1403 13
rect 3196 -17 3203 56
rect 3476 47 3483 143
rect 3176 -24 3203 -17
rect 3216 -24 3223 33
rect 3536 -17 3543 193
rect 3596 176 3603 353
rect 3616 207 3623 516
rect 3636 188 3643 493
rect 3676 47 3683 173
rect 3696 146 3703 193
rect 3736 176 3743 433
rect 3756 207 3763 393
rect 3776 176 3783 233
rect 3816 187 3823 293
rect 3856 287 3863 363
rect 3916 267 3923 393
rect 3756 87 3763 143
rect 3936 27 3943 1013
rect 4236 1007 4243 1353
rect 4356 1347 4363 1403
rect 4416 1400 4423 1403
rect 4413 1387 4427 1400
rect 4476 1387 4483 1533
rect 4496 1327 4503 1773
rect 4656 1706 4663 1853
rect 4676 1748 4683 1953
rect 4576 1627 4583 1693
rect 4576 1527 4583 1613
rect 4516 1487 4523 1513
rect 4516 1443 4523 1473
rect 4596 1448 4603 1533
rect 4516 1436 4543 1443
rect 4496 1287 4503 1313
rect 3956 886 3963 913
rect 4096 887 4103 933
rect 4116 883 4123 993
rect 4176 916 4203 923
rect 4116 876 4143 883
rect 4016 727 4023 872
rect 4196 867 4203 916
rect 4216 907 4223 953
rect 4256 916 4263 1273
rect 4356 1207 4363 1233
rect 4376 1187 4383 1214
rect 4396 1147 4403 1213
rect 4616 1186 4623 1373
rect 4636 1347 4643 1473
rect 4676 1307 4683 1734
rect 4776 1667 4783 1703
rect 4836 1667 4843 1703
rect 4747 1436 4763 1443
rect 4516 1180 4523 1183
rect 4327 1136 4353 1143
rect 4296 916 4303 1033
rect 4336 916 4343 1113
rect 4436 916 4443 1172
rect 4513 1167 4527 1180
rect 3976 627 3983 663
rect 4016 587 4023 663
rect 4056 627 4063 663
rect 4016 507 4023 573
rect 4056 407 4063 613
rect 4156 447 4163 853
rect 4236 696 4243 753
rect 4176 666 4183 693
rect 4067 396 4083 403
rect 4076 307 4083 396
rect 4156 267 4163 433
rect 3956 146 3963 233
rect 3536 -24 3563 -17
rect 4016 -24 4023 13
rect 4056 -24 4063 253
rect 4096 107 4103 213
rect 4153 180 4167 193
rect 4156 176 4163 180
rect 4176 140 4183 143
rect 4136 107 4143 132
rect 4173 127 4187 140
rect 4216 127 4223 253
rect 4256 143 4263 573
rect 4276 367 4283 883
rect 4296 408 4303 793
rect 4316 767 4323 883
rect 4396 696 4403 913
rect 4456 707 4463 883
rect 4516 807 4523 1013
rect 4596 916 4603 953
rect 4640 923 4653 927
rect 4636 916 4653 923
rect 4496 696 4503 753
rect 4536 727 4543 914
rect 4640 913 4653 916
rect 4676 886 4683 953
rect 4736 916 4743 1293
rect 4756 1027 4763 1436
rect 4796 1167 4803 1533
rect 4856 1436 4863 1533
rect 4936 1448 4943 1953
rect 4876 1183 4883 1373
rect 4956 1223 4963 1533
rect 4936 1216 4963 1223
rect 4856 1176 4883 1183
rect 4796 923 4803 1153
rect 4896 1107 4903 1214
rect 4893 943 4907 953
rect 4876 940 4907 943
rect 4876 936 4903 940
rect 4796 916 4823 923
rect 4876 916 4883 936
rect 4576 880 4583 883
rect 4573 867 4587 880
rect 4696 823 4703 913
rect 4916 887 4923 1073
rect 4936 1007 4943 1216
rect 4996 1147 5003 1183
rect 4676 816 4703 823
rect 4676 747 4683 816
rect 4936 807 4943 953
rect 5016 928 5023 1313
rect 5036 967 5043 1433
rect 5056 1228 5063 2293
rect 5216 2268 5223 2474
rect 5236 2307 5243 2793
rect 5256 2487 5263 2956
rect 5296 2807 5303 3353
rect 5416 3327 5423 3483
rect 5436 3266 5443 3353
rect 5476 3347 5483 3553
rect 5496 3296 5503 3573
rect 5516 3567 5523 3873
rect 5536 3787 5543 4003
rect 5616 3967 5623 4173
rect 5556 3807 5563 3853
rect 5616 3816 5623 3932
rect 5636 3927 5643 4233
rect 5776 4167 5783 4353
rect 5796 4306 5803 4413
rect 5836 4336 5843 4413
rect 5876 4336 5883 4453
rect 5896 4387 5903 4493
rect 5916 4367 5923 4523
rect 5956 4403 5963 4793
rect 5976 4767 5983 4816
rect 6036 4820 6043 4823
rect 6016 4747 6023 4813
rect 6033 4807 6047 4820
rect 6136 4823 6143 4976
rect 6116 4816 6143 4823
rect 6056 4767 6063 4793
rect 5976 4527 5983 4732
rect 5996 4567 6003 4733
rect 6036 4556 6043 4593
rect 5936 4396 5963 4403
rect 5796 4207 5803 4233
rect 5696 4036 5703 4133
rect 5733 4040 5747 4053
rect 5736 4036 5743 4040
rect 5676 3967 5683 4003
rect 5716 3867 5723 4003
rect 5776 3947 5783 4132
rect 5816 4036 5823 4193
rect 5856 4167 5863 4303
rect 5916 4006 5923 4053
rect 5796 3907 5803 3993
rect 5876 3987 5883 4003
rect 5876 3976 5893 3987
rect 5880 3973 5893 3976
rect 5936 3947 5943 4396
rect 5956 4067 5963 4373
rect 5976 4147 5983 4492
rect 6056 4407 6063 4473
rect 6096 4467 6103 4513
rect 6116 4443 6123 4816
rect 6096 4436 6123 4443
rect 5996 4227 6003 4303
rect 6056 4207 6063 4292
rect 6076 4183 6083 4413
rect 6056 4176 6083 4183
rect 5996 4036 6003 4073
rect 6056 4047 6063 4176
rect 6096 4067 6103 4436
rect 6136 4427 6143 4793
rect 6156 4727 6163 4996
rect 6176 4867 6183 4953
rect 6196 4868 6203 5016
rect 6236 4867 6243 5076
rect 6176 4687 6183 4813
rect 6167 4676 6183 4687
rect 6167 4673 6180 4676
rect 6176 4556 6183 4653
rect 6196 4587 6203 4793
rect 6216 4556 6223 4593
rect 6236 4587 6243 4813
rect 6256 4567 6263 5293
rect 6276 5087 6283 5253
rect 6296 5187 6303 5332
rect 6336 5307 6343 5513
rect 6376 5507 6383 5553
rect 6356 5346 6363 5473
rect 6376 5127 6383 5373
rect 6396 5247 6403 5933
rect 6416 5103 6423 5973
rect 6436 5267 6443 5894
rect 6396 5096 6423 5103
rect 6287 5043 6300 5046
rect 6287 5036 6303 5043
rect 6287 5033 6300 5036
rect 6296 4947 6303 5013
rect 6276 4568 6283 4873
rect 6296 4867 6303 4933
rect 6336 4887 6343 5043
rect 6333 4860 6347 4873
rect 6373 4860 6387 4873
rect 6396 4867 6403 5096
rect 6416 4987 6423 5074
rect 6336 4856 6343 4860
rect 6376 4856 6383 4860
rect 6356 4787 6363 4823
rect 6336 4587 6343 4713
rect 6356 4667 6363 4752
rect 6356 4556 6363 4653
rect 6276 4527 6283 4554
rect 6156 4336 6163 4513
rect 6196 4467 6203 4523
rect 6253 4503 6267 4513
rect 6236 4500 6267 4503
rect 6236 4496 6263 4500
rect 6216 4387 6223 4493
rect 6216 4306 6223 4333
rect 6236 4303 6243 4496
rect 6336 4347 6343 4512
rect 6236 4296 6263 4303
rect 5976 4000 5983 4003
rect 5973 3987 5987 4000
rect 5673 3847 5687 3853
rect 5747 3836 5823 3843
rect 5816 3816 5823 3836
rect 5836 3827 5843 3933
rect 5636 3780 5643 3783
rect 5540 3766 5560 3767
rect 5547 3753 5553 3766
rect 5596 3607 5603 3772
rect 5633 3767 5647 3780
rect 5716 3747 5723 3813
rect 5716 3567 5723 3733
rect 5756 3707 5763 3783
rect 5536 3516 5543 3553
rect 5716 3543 5723 3553
rect 5716 3536 5743 3543
rect 5736 3516 5743 3536
rect 5636 3487 5643 3514
rect 5596 3407 5603 3483
rect 5576 3303 5583 3333
rect 5576 3296 5603 3303
rect 5633 3300 5647 3313
rect 5636 3296 5643 3300
rect 5596 3266 5603 3296
rect 5356 3260 5363 3263
rect 5353 3247 5367 3260
rect 5476 3207 5483 3263
rect 5516 3243 5523 3263
rect 5516 3236 5543 3243
rect 5376 2996 5383 3173
rect 5356 2803 5363 2963
rect 5436 2827 5443 3093
rect 5456 2966 5463 3133
rect 5496 2996 5503 3053
rect 5536 3008 5543 3236
rect 5656 3147 5663 3263
rect 5716 3167 5723 3472
rect 5756 3447 5763 3483
rect 5796 3347 5803 3553
rect 5816 3527 5823 3593
rect 5836 3543 5843 3772
rect 5856 3567 5863 3933
rect 5876 3783 5883 3913
rect 5936 3816 5943 3893
rect 5876 3776 5903 3783
rect 5836 3536 5853 3543
rect 5856 3516 5863 3532
rect 5876 3527 5883 3753
rect 5856 3347 5863 3393
rect 5736 3127 5743 3333
rect 5813 3300 5827 3313
rect 5816 3296 5823 3300
rect 5753 3263 5767 3273
rect 5753 3260 5783 3263
rect 5756 3256 5783 3260
rect 5836 3207 5843 3263
rect 5856 3107 5863 3292
rect 5847 3096 5863 3107
rect 5847 3093 5860 3096
rect 5596 2966 5603 3053
rect 5813 3000 5827 3013
rect 5853 3000 5867 3013
rect 5876 3007 5883 3473
rect 5816 2996 5823 3000
rect 5856 2996 5863 3000
rect 5736 2967 5743 2994
rect 5356 2796 5383 2803
rect 5276 2743 5283 2773
rect 5276 2736 5293 2743
rect 5356 2667 5363 2743
rect 5296 2476 5303 2613
rect 5356 2483 5363 2653
rect 5336 2476 5363 2483
rect 5276 2307 5283 2443
rect 5316 2407 5323 2443
rect 5176 2187 5183 2254
rect 5216 2203 5223 2254
rect 5316 2226 5323 2293
rect 5376 2287 5383 2796
rect 5436 2788 5443 2813
rect 5516 2783 5523 2963
rect 5696 2847 5703 2963
rect 5836 2927 5843 2963
rect 5896 2907 5903 3776
rect 5916 3747 5923 3783
rect 5953 3767 5967 3772
rect 5916 3327 5923 3533
rect 5996 3527 6003 3913
rect 6016 3827 6023 3993
rect 6036 3947 6043 4033
rect 6056 3927 6063 3993
rect 6056 3816 6063 3853
rect 6096 3827 6103 4003
rect 6136 3987 6143 4053
rect 6196 4036 6203 4073
rect 6236 4036 6243 4153
rect 6256 4103 6263 4296
rect 6276 4287 6283 4303
rect 6276 4127 6283 4273
rect 6316 4227 6323 4303
rect 6256 4096 6283 4103
rect 6096 3816 6113 3827
rect 6100 3814 6113 3816
rect 5956 3447 5963 3483
rect 6016 3447 6023 3773
rect 6036 3747 6043 3783
rect 6076 3780 6083 3783
rect 6073 3767 6087 3780
rect 6116 3567 6123 3773
rect 6136 3687 6143 3973
rect 6176 3947 6183 4003
rect 5967 3436 5983 3443
rect 5976 3387 5983 3436
rect 5920 3306 5940 3307
rect 5927 3303 5940 3306
rect 5927 3296 5943 3303
rect 5976 3296 5983 3373
rect 5927 3294 5940 3296
rect 5936 3293 5940 3294
rect 5936 3027 5943 3073
rect 6036 3027 6043 3553
rect 6136 3516 6143 3593
rect 6156 3587 6163 3873
rect 6216 3867 6223 4003
rect 6276 4003 6283 4096
rect 6316 4067 6323 4093
rect 6356 4067 6363 4353
rect 6376 4167 6383 4373
rect 6376 4036 6383 4093
rect 6396 4043 6403 4813
rect 6416 4787 6423 4973
rect 6436 4907 6443 5113
rect 6416 4367 6423 4752
rect 6436 4667 6443 4872
rect 6436 4527 6443 4613
rect 6436 4387 6443 4433
rect 6416 4063 6423 4332
rect 6436 4247 6443 4333
rect 6416 4056 6443 4063
rect 6396 4036 6423 4043
rect 6276 3996 6303 4003
rect 6256 3947 6263 3993
rect 6276 3827 6283 3853
rect 6216 3780 6223 3783
rect 6256 3780 6263 3783
rect 6176 3663 6183 3773
rect 6213 3767 6227 3780
rect 6253 3767 6267 3780
rect 6216 3727 6223 3753
rect 6176 3656 6203 3663
rect 6053 3467 6067 3473
rect 6076 3347 6083 3483
rect 6076 3296 6083 3333
rect 6176 3327 6183 3613
rect 6196 3403 6203 3656
rect 6256 3607 6263 3753
rect 6216 3527 6223 3593
rect 6256 3516 6263 3553
rect 6196 3396 6223 3403
rect 6096 3207 6103 3263
rect 5936 2996 5943 3013
rect 5996 2996 6023 3003
rect 5916 2927 5923 2993
rect 5516 2776 5543 2783
rect 5456 2707 5463 2732
rect 5496 2627 5503 2743
rect 5516 2483 5523 2733
rect 5536 2527 5543 2776
rect 5656 2746 5663 2813
rect 5576 2707 5583 2743
rect 5656 2527 5663 2693
rect 5716 2667 5723 2743
rect 5796 2627 5803 2773
rect 5816 2767 5823 2833
rect 5516 2476 5543 2483
rect 5656 2483 5663 2513
rect 5656 2476 5683 2483
rect 5796 2443 5803 2533
rect 5416 2407 5423 2443
rect 5556 2327 5563 2443
rect 5776 2436 5803 2443
rect 5216 2196 5243 2203
rect 5096 1963 5103 2113
rect 5096 1956 5123 1963
rect 5196 1956 5203 1993
rect 5236 1987 5243 2196
rect 5296 2027 5303 2223
rect 5356 2216 5383 2223
rect 5356 2187 5363 2216
rect 5356 2047 5363 2173
rect 5233 1960 5247 1973
rect 5236 1956 5243 1960
rect 5076 1287 5083 1833
rect 5116 1768 5123 1956
rect 5136 1687 5143 1703
rect 5136 1676 5153 1687
rect 5140 1673 5153 1676
rect 5116 1587 5123 1653
rect 5116 1448 5123 1573
rect 5076 1223 5083 1273
rect 5156 1247 5163 1613
rect 5176 1387 5183 1773
rect 5216 1743 5223 1923
rect 5276 1783 5283 1973
rect 5376 1956 5383 2193
rect 5416 2087 5423 2223
rect 5456 2167 5463 2253
rect 5536 2147 5543 2223
rect 5576 2087 5583 2213
rect 5276 1776 5293 1783
rect 5316 1783 5323 1923
rect 5307 1776 5323 1783
rect 5196 1736 5223 1743
rect 5196 1706 5203 1736
rect 5296 1736 5303 1773
rect 5276 1687 5283 1703
rect 5247 1676 5273 1683
rect 5336 1467 5343 1733
rect 5356 1667 5363 1923
rect 5416 1887 5423 2073
rect 5436 1787 5443 2033
rect 5556 1926 5563 1973
rect 5576 1963 5583 2013
rect 5596 1987 5603 2313
rect 5616 2187 5623 2293
rect 5696 2256 5703 2293
rect 5736 2267 5743 2403
rect 5836 2387 5843 2892
rect 6016 2887 6023 2996
rect 6036 2966 6043 3013
rect 6096 2996 6103 3113
rect 6136 3107 6143 3313
rect 6196 3296 6203 3373
rect 6216 3347 6223 3396
rect 6236 3296 6243 3433
rect 6216 3207 6223 3263
rect 6136 2996 6143 3093
rect 6276 3067 6283 3473
rect 6236 2966 6243 3053
rect 6296 3047 6303 3996
rect 6316 3907 6323 4003
rect 6336 3847 6343 3973
rect 6356 3967 6363 4003
rect 6356 3887 6363 3953
rect 6356 3816 6363 3852
rect 6396 3827 6403 3893
rect 6327 3776 6343 3783
rect 6316 3303 6323 3773
rect 6376 3727 6383 3783
rect 6336 3527 6343 3673
rect 6356 3516 6363 3553
rect 6396 3547 6403 3773
rect 6416 3627 6423 4036
rect 6436 3967 6443 4056
rect 6436 3603 6443 3853
rect 6416 3596 6443 3603
rect 6416 3523 6423 3596
rect 6396 3516 6423 3523
rect 6336 3327 6343 3473
rect 6376 3407 6383 3483
rect 6436 3423 6443 3573
rect 6416 3416 6443 3423
rect 6316 3296 6343 3303
rect 6376 3296 6383 3333
rect 6416 3307 6423 3416
rect 6376 3003 6383 3093
rect 6436 3087 6443 3393
rect 6356 2996 6383 3003
rect 5856 2736 5873 2743
rect 5856 2443 5863 2736
rect 5976 2547 5983 2873
rect 6016 2776 6023 2833
rect 6036 2827 6043 2952
rect 6056 2788 6063 2953
rect 6247 2956 6263 2963
rect 6036 2488 6043 2743
rect 6116 2446 6123 2913
rect 6196 2776 6203 2873
rect 6296 2776 6303 2813
rect 6376 2747 6383 2973
rect 6156 2707 6163 2743
rect 6216 2488 6223 2743
rect 6316 2483 6323 2732
rect 6296 2476 6323 2483
rect 5856 2436 5883 2443
rect 5856 2226 5863 2293
rect 5756 2167 5763 2223
rect 5816 2220 5823 2223
rect 5813 2207 5827 2220
rect 5876 2207 5883 2373
rect 5916 2347 5923 2403
rect 5576 1956 5603 1963
rect 5636 1956 5643 1993
rect 5676 1956 5683 2073
rect 5716 1968 5723 2153
rect 5773 1960 5787 1973
rect 5836 1968 5843 2013
rect 5776 1956 5783 1960
rect 5476 1807 5483 1923
rect 5656 1887 5663 1923
rect 5396 1627 5403 1703
rect 5436 1700 5443 1703
rect 5433 1687 5447 1700
rect 5476 1547 5483 1733
rect 5496 1707 5503 1773
rect 5596 1747 5603 1873
rect 5233 1440 5247 1453
rect 5236 1436 5243 1440
rect 5216 1347 5223 1403
rect 5076 1216 5103 1223
rect 5156 1143 5163 1183
rect 5136 1136 5163 1143
rect 5116 1047 5123 1093
rect 5027 916 5043 923
rect 4996 880 5003 883
rect 4993 867 5007 880
rect 4536 663 4543 713
rect 4633 700 4647 713
rect 4636 696 4643 700
rect 4536 656 4563 663
rect 4316 176 4323 273
rect 4256 136 4283 143
rect 4336 27 4343 393
rect 4436 287 4443 363
rect 4456 207 4463 613
rect 4516 396 4523 473
rect 4556 408 4563 656
rect 4616 587 4623 663
rect 4676 627 4683 663
rect 4696 396 4703 493
rect 4776 483 4783 793
rect 4856 696 4863 753
rect 4976 708 4983 793
rect 4756 476 4783 483
rect 4756 427 4763 476
rect 4936 447 4943 694
rect 5036 687 5043 916
rect 5056 867 5063 953
rect 5136 916 5143 1136
rect 5176 928 5183 1113
rect 5196 1067 5203 1273
rect 5216 1186 5223 1293
rect 5276 1267 5283 1453
rect 5353 1440 5367 1453
rect 5356 1436 5363 1440
rect 5396 1436 5403 1533
rect 5536 1487 5543 1613
rect 5576 1607 5583 1703
rect 5616 1527 5623 1753
rect 5616 1436 5623 1513
rect 5516 1407 5523 1434
rect 5336 1400 5343 1403
rect 5333 1387 5347 1400
rect 5436 1347 5443 1403
rect 5233 1223 5247 1233
rect 5233 1220 5263 1223
rect 5236 1216 5263 1220
rect 5296 1216 5303 1293
rect 5336 1227 5343 1333
rect 5356 1186 5363 1253
rect 5376 1216 5403 1223
rect 5296 987 5303 1133
rect 5376 1047 5383 1216
rect 5576 1187 5583 1313
rect 5656 1307 5663 1793
rect 5716 1736 5743 1743
rect 5736 1567 5743 1736
rect 5756 1706 5763 1813
rect 5836 1767 5843 1954
rect 5876 1736 5883 1793
rect 5836 1696 5863 1703
rect 5436 1127 5443 1183
rect 5116 880 5123 883
rect 5113 867 5127 880
rect 5116 696 5123 753
rect 5136 747 5143 833
rect 5156 807 5163 883
rect 5216 696 5223 933
rect 5256 916 5263 953
rect 5296 916 5303 973
rect 5276 847 5283 883
rect 5253 700 5267 713
rect 5256 696 5263 700
rect 4996 507 5003 663
rect 5096 587 5103 663
rect 5193 647 5207 653
rect 4756 396 4763 413
rect 4476 327 4483 393
rect 4616 367 4623 394
rect 4976 367 4983 433
rect 5093 400 5107 413
rect 5096 396 5103 400
rect 5176 367 5183 593
rect 5236 587 5243 663
rect 5316 607 5323 713
rect 5336 707 5343 913
rect 5376 867 5383 1033
rect 5416 916 5423 993
rect 5436 927 5443 1113
rect 5576 916 5583 1073
rect 5596 947 5603 1293
rect 5656 1216 5663 1272
rect 5676 1227 5683 1513
rect 5836 1436 5843 1673
rect 5856 1667 5863 1696
rect 5856 1607 5863 1653
rect 5716 1287 5723 1403
rect 5816 1186 5823 1273
rect 5836 1127 5843 1373
rect 5856 1347 5863 1403
rect 5896 1400 5903 1403
rect 5893 1387 5907 1400
rect 5476 883 5483 913
rect 5456 876 5483 883
rect 5376 696 5383 753
rect 5396 607 5403 663
rect 5436 660 5443 663
rect 5433 647 5447 660
rect 5456 527 5463 653
rect 5207 423 5220 427
rect 5207 413 5223 423
rect 5216 396 5223 413
rect 4716 327 4723 363
rect 5036 327 5043 353
rect 5116 360 5123 363
rect 5113 347 5127 360
rect 5247 356 5283 363
rect 4487 316 4503 323
rect 4496 146 4503 316
rect 4416 107 4423 143
rect 4516 127 4523 213
rect 4556 176 4563 253
rect 4756 146 4763 173
rect 4576 140 4583 143
rect 4536 87 4543 133
rect 4573 127 4587 140
rect 4616 107 4623 143
rect 4876 107 4883 173
rect 4996 140 5003 143
rect 4956 107 4963 132
rect 4993 127 5007 140
rect 5036 127 5043 233
rect 5096 176 5103 313
rect 5256 188 5263 333
rect 5356 188 5363 513
rect 5476 423 5483 663
rect 5576 663 5583 853
rect 5596 667 5603 883
rect 5653 700 5667 713
rect 5656 696 5663 700
rect 5556 656 5583 663
rect 5467 416 5483 423
rect 5453 400 5467 413
rect 5456 396 5463 400
rect 5496 203 5503 413
rect 5556 363 5563 656
rect 5696 403 5703 872
rect 5716 447 5723 933
rect 5736 916 5743 1093
rect 5776 787 5783 883
rect 5773 700 5787 713
rect 5776 696 5783 700
rect 5816 667 5823 914
rect 5836 727 5843 1113
rect 5916 928 5923 1153
rect 5936 1107 5943 2193
rect 5976 2147 5983 2333
rect 6116 2327 6123 2432
rect 6076 2256 6083 2293
rect 6196 2283 6203 2443
rect 6276 2427 6283 2473
rect 6296 2446 6303 2476
rect 6336 2440 6343 2443
rect 6376 2440 6383 2443
rect 6333 2427 6347 2440
rect 6373 2427 6387 2440
rect 6196 2276 6223 2283
rect 6216 2256 6223 2276
rect 6396 2256 6403 2313
rect 6416 2287 6423 2473
rect 6016 2227 6023 2254
rect 6036 1983 6043 2013
rect 6056 2007 6063 2212
rect 6096 2087 6103 2223
rect 6236 2047 6243 2223
rect 6276 2207 6283 2223
rect 6276 2087 6283 2193
rect 6316 2147 6323 2254
rect 6376 2220 6383 2223
rect 6373 2207 6387 2220
rect 6036 1976 6063 1983
rect 6056 1956 6063 1976
rect 6136 1963 6143 2033
rect 6376 2027 6383 2133
rect 6116 1956 6143 1963
rect 5956 1887 5963 1953
rect 5956 1127 5963 1873
rect 6156 1807 6163 1993
rect 6376 1956 6383 2013
rect 6116 1707 6123 1793
rect 5976 1696 6003 1703
rect 5976 1647 5983 1696
rect 6056 1587 6063 1703
rect 6136 1523 6143 1773
rect 6316 1736 6323 1773
rect 6256 1706 6263 1733
rect 6216 1683 6223 1692
rect 6196 1676 6223 1683
rect 6196 1667 6203 1676
rect 6136 1516 6163 1523
rect 6036 1436 6043 1473
rect 6076 1436 6083 1513
rect 6156 1443 6163 1516
rect 6136 1436 6163 1443
rect 6016 1247 6023 1403
rect 6176 1307 6183 1473
rect 6196 1387 6203 1653
rect 6336 1448 6343 1703
rect 5976 1186 5983 1233
rect 6036 1216 6043 1253
rect 6076 1228 6083 1293
rect 6053 1167 6067 1172
rect 5956 886 5963 1053
rect 5896 867 5903 883
rect 5896 856 5913 867
rect 5900 853 5913 856
rect 5896 696 5903 773
rect 5956 703 5963 872
rect 5976 867 5983 933
rect 6016 916 6023 1013
rect 6116 943 6123 1253
rect 6256 1227 6263 1392
rect 6316 1216 6323 1273
rect 6156 1180 6163 1183
rect 6153 1167 6167 1180
rect 6196 1167 6203 1183
rect 6176 1156 6193 1163
rect 6176 987 6183 1156
rect 6116 936 6143 943
rect 6116 887 6123 914
rect 6036 847 6043 883
rect 6087 876 6103 883
rect 5936 696 5963 703
rect 6096 696 6103 876
rect 6136 666 6143 936
rect 6173 920 6187 933
rect 6176 916 6183 920
rect 6216 916 6223 1173
rect 6236 1167 6243 1213
rect 6256 1167 6263 1192
rect 6296 1180 6303 1183
rect 6293 1167 6307 1180
rect 5876 587 5883 663
rect 5916 567 5923 663
rect 6036 607 6043 663
rect 5696 396 5713 403
rect 5756 396 5763 433
rect 6036 408 6043 473
rect 5556 356 5583 363
rect 5576 287 5583 356
rect 5796 347 5803 393
rect 5476 196 5503 203
rect 5076 107 5083 143
rect 5156 127 5163 174
rect 5476 146 5483 196
rect 5856 147 5863 363
rect 5896 360 5903 363
rect 5893 347 5907 360
rect 5956 287 5963 394
rect 6076 343 6083 553
rect 6236 487 6243 872
rect 6276 667 6283 693
rect 6096 367 6103 413
rect 6133 400 6147 413
rect 6296 423 6303 1113
rect 6336 847 6343 883
rect 6313 700 6327 713
rect 6316 696 6323 700
rect 6296 416 6323 423
rect 6173 400 6187 413
rect 6136 396 6143 400
rect 6176 396 6183 400
rect 6076 340 6103 343
rect 6076 336 6107 340
rect 6093 327 6107 336
rect 6156 327 6163 363
rect 5876 147 5883 273
rect 5196 87 5203 143
rect 5516 140 5523 143
rect 5513 127 5527 140
rect 5633 127 5647 133
rect 6076 146 6083 293
rect 6236 187 6243 413
rect 6273 400 6287 413
rect 6276 396 6283 400
rect 6316 396 6323 416
rect 6296 307 6303 363
rect 6336 327 6343 363
rect 6376 267 6383 413
rect 6396 327 6403 1193
rect 6436 1186 6443 2013
rect 6196 147 6203 174
rect 6296 176 6303 253
rect 6396 227 6403 313
rect 5976 140 5983 143
rect 5973 127 5987 140
rect 6316 140 6323 143
rect 6313 127 6327 140
rect 6396 127 6403 213
rect 4607 76 4633 83
rect 4947 76 4973 83
rect 5067 76 5093 83
rect 4136 -24 4143 13
<< m3contact >>
rect 2093 6253 2107 6267
rect 2133 6253 2147 6267
rect 1513 6233 1527 6247
rect 1273 6213 1287 6227
rect 1413 6213 1427 6227
rect 593 6193 607 6207
rect 673 6193 687 6207
rect 1033 6193 1047 6207
rect 153 6153 167 6167
rect 253 6153 267 6167
rect 373 6153 387 6167
rect 113 6114 127 6128
rect 193 6114 207 6128
rect 353 6133 367 6147
rect 293 6114 307 6128
rect 93 6053 107 6067
rect 133 5993 147 6007
rect 53 5933 67 5947
rect 113 5894 127 5908
rect 153 5894 167 5908
rect 93 5833 107 5847
rect 173 5853 187 5867
rect 153 5833 167 5847
rect 53 5793 67 5807
rect 133 5793 147 5807
rect 113 5594 127 5608
rect 93 5552 107 5566
rect 233 6073 247 6087
rect 233 6033 247 6047
rect 313 6033 327 6047
rect 273 5993 287 6007
rect 233 5933 247 5947
rect 273 5933 287 5947
rect 453 6173 467 6187
rect 513 6173 527 6187
rect 433 6153 447 6167
rect 493 6153 507 6167
rect 413 6133 427 6147
rect 473 6114 487 6128
rect 533 6114 547 6128
rect 633 6114 647 6128
rect 373 6073 387 6087
rect 413 6072 427 6086
rect 353 5993 367 6007
rect 513 6073 527 6087
rect 493 6053 507 6067
rect 493 5993 507 6007
rect 353 5953 367 5967
rect 253 5852 267 5866
rect 293 5852 307 5866
rect 333 5853 347 5867
rect 193 5833 207 5847
rect 193 5614 207 5628
rect 193 5594 207 5608
rect 233 5594 247 5608
rect 173 5552 187 5566
rect 213 5552 227 5566
rect 253 5533 267 5547
rect 213 5493 227 5507
rect 153 5413 167 5427
rect 73 5374 87 5388
rect 153 5374 167 5388
rect 213 5374 227 5388
rect 393 5894 407 5908
rect 453 5973 467 5987
rect 473 5933 487 5947
rect 473 5893 487 5907
rect 413 5852 427 5866
rect 353 5793 367 5807
rect 533 5953 547 5967
rect 573 6072 587 6086
rect 653 6073 667 6087
rect 633 6053 647 6067
rect 613 5973 627 5987
rect 693 6153 707 6167
rect 773 6153 787 6167
rect 913 6153 927 6167
rect 1033 6153 1047 6167
rect 733 6114 747 6128
rect 833 6114 847 6128
rect 873 6114 887 6128
rect 913 6114 927 6128
rect 1073 6114 1087 6128
rect 1173 6114 1187 6128
rect 1413 6173 1427 6187
rect 1393 6153 1407 6167
rect 1493 6153 1507 6167
rect 1313 6114 1327 6128
rect 693 6073 707 6087
rect 753 6072 767 6086
rect 733 6053 747 6067
rect 713 5993 727 6007
rect 673 5973 687 5987
rect 653 5953 667 5967
rect 553 5914 567 5928
rect 613 5913 627 5927
rect 573 5894 587 5908
rect 513 5853 527 5867
rect 553 5852 567 5866
rect 673 5933 687 5947
rect 793 6013 807 6027
rect 993 6093 1007 6107
rect 893 6072 907 6086
rect 933 6013 947 6027
rect 853 5993 867 6007
rect 753 5973 767 5987
rect 793 5973 807 5987
rect 833 5973 847 5987
rect 733 5893 747 5907
rect 813 5933 827 5947
rect 793 5893 807 5907
rect 933 5992 947 6006
rect 913 5894 927 5908
rect 833 5852 847 5866
rect 753 5833 767 5847
rect 873 5833 887 5847
rect 693 5693 707 5707
rect 393 5613 407 5627
rect 453 5613 467 5627
rect 493 5613 507 5627
rect 313 5594 327 5608
rect 353 5594 367 5608
rect 513 5593 527 5607
rect 613 5594 627 5608
rect 653 5594 667 5608
rect 773 5633 787 5647
rect 333 5552 347 5566
rect 373 5552 387 5566
rect 293 5533 307 5547
rect 333 5493 347 5507
rect 293 5473 307 5487
rect 53 5333 67 5347
rect 13 5133 27 5147
rect 93 5332 107 5346
rect 273 5373 287 5387
rect 53 5093 67 5107
rect 113 5074 127 5088
rect 233 5332 247 5346
rect 453 5552 467 5566
rect 533 5552 547 5566
rect 593 5552 607 5566
rect 493 5493 507 5507
rect 533 5473 547 5487
rect 813 5594 827 5608
rect 673 5552 687 5566
rect 713 5552 727 5566
rect 773 5553 787 5567
rect 833 5552 847 5566
rect 613 5433 627 5447
rect 373 5413 387 5427
rect 413 5413 427 5427
rect 593 5413 607 5427
rect 313 5373 327 5387
rect 413 5374 427 5388
rect 453 5374 467 5388
rect 493 5374 507 5388
rect 533 5374 547 5388
rect 293 5153 307 5167
rect 233 5093 247 5107
rect 193 5074 207 5088
rect 273 5074 287 5088
rect 393 5332 407 5346
rect 453 5213 467 5227
rect 373 5153 387 5167
rect 353 5093 367 5107
rect 413 5133 427 5147
rect 53 5032 67 5046
rect 53 4993 67 5007
rect 13 4733 27 4747
rect 133 5032 147 5046
rect 193 5033 207 5047
rect 253 5032 267 5046
rect 193 4953 207 4967
rect 53 4853 67 4867
rect 93 4854 107 4868
rect 173 4854 187 4868
rect 73 4812 87 4826
rect 113 4812 127 4826
rect 253 4913 267 4927
rect 313 5033 327 5047
rect 313 4933 327 4947
rect 293 4893 307 4907
rect 573 5333 587 5347
rect 1053 6053 1067 6067
rect 1093 6033 1107 6047
rect 1333 6072 1347 6086
rect 1313 6053 1327 6067
rect 1293 5993 1307 6007
rect 1333 5993 1347 6007
rect 1033 5953 1047 5967
rect 1193 5953 1207 5967
rect 1233 5953 1247 5967
rect 993 5894 1007 5908
rect 1073 5894 1087 5908
rect 1133 5894 1147 5908
rect 1173 5894 1187 5908
rect 1013 5833 1027 5847
rect 1033 5833 1047 5847
rect 1333 5913 1347 5927
rect 973 5813 987 5827
rect 1073 5813 1087 5827
rect 1233 5852 1247 5866
rect 1273 5852 1287 5866
rect 1313 5852 1327 5866
rect 1433 6114 1447 6128
rect 1433 5993 1447 6007
rect 1493 6072 1507 6086
rect 1993 6213 2007 6227
rect 1673 6193 1687 6207
rect 1973 6193 1987 6207
rect 1573 6173 1587 6187
rect 1613 6114 1627 6128
rect 1653 6114 1667 6128
rect 1553 6072 1567 6086
rect 1733 6153 1747 6167
rect 2033 6193 2047 6207
rect 1993 6173 2007 6187
rect 1793 6114 1807 6128
rect 1833 6114 1847 6128
rect 1873 6114 1887 6128
rect 1933 6113 1947 6127
rect 2013 6153 2027 6167
rect 2033 6114 2047 6128
rect 1673 6072 1687 6086
rect 1713 6072 1727 6086
rect 1753 6072 1767 6086
rect 1793 6073 1807 6087
rect 1513 6053 1527 6067
rect 1653 6053 1667 6067
rect 1693 6033 1707 6047
rect 1733 6033 1747 6047
rect 1693 5993 1707 6007
rect 1453 5973 1467 5987
rect 1673 5953 1687 5967
rect 1753 5953 1767 5967
rect 1433 5933 1447 5947
rect 1593 5933 1607 5947
rect 1653 5933 1667 5947
rect 1513 5913 1527 5927
rect 1433 5894 1447 5908
rect 1493 5894 1507 5908
rect 1473 5833 1487 5847
rect 913 5793 927 5807
rect 1033 5793 1047 5807
rect 1153 5793 1167 5807
rect 1493 5793 1507 5807
rect 973 5653 987 5667
rect 933 5633 947 5647
rect 933 5594 947 5608
rect 993 5593 1007 5607
rect 873 5513 887 5527
rect 693 5473 707 5487
rect 673 5393 687 5407
rect 613 5373 627 5387
rect 653 5374 667 5388
rect 773 5433 787 5447
rect 753 5373 767 5387
rect 593 5253 607 5267
rect 593 5213 607 5227
rect 253 4854 267 4868
rect 293 4854 307 4868
rect 333 4852 347 4866
rect 193 4812 207 4826
rect 233 4812 247 4826
rect 273 4812 287 4826
rect 173 4773 187 4787
rect 113 4593 127 4607
rect 153 4593 167 4607
rect 313 4593 327 4607
rect 113 4554 127 4568
rect 153 4554 167 4568
rect 193 4554 207 4568
rect 253 4573 267 4587
rect 333 4573 347 4587
rect 33 4512 47 4526
rect 73 4513 87 4527
rect 53 4393 67 4407
rect 53 4333 67 4347
rect 93 4512 107 4526
rect 173 4513 187 4527
rect 133 4393 147 4407
rect 173 4373 187 4387
rect 113 4334 127 4348
rect 173 4333 187 4347
rect 53 4293 67 4307
rect 33 4073 47 4087
rect 13 3953 27 3967
rect 13 3893 27 3907
rect 13 3852 27 3866
rect 13 3613 27 3627
rect 13 3133 27 3147
rect 93 4292 107 4306
rect 133 4253 147 4267
rect 273 4493 287 4507
rect 333 4513 347 4527
rect 313 4473 327 4487
rect 493 5073 507 5087
rect 513 5073 527 5087
rect 553 5073 567 5087
rect 673 5332 687 5346
rect 653 5253 667 5267
rect 713 5193 727 5207
rect 653 5173 667 5187
rect 393 4993 407 5007
rect 373 4893 387 4907
rect 433 4973 447 4987
rect 413 4933 427 4947
rect 393 4873 407 4887
rect 453 4893 467 4907
rect 433 4812 447 4826
rect 533 5032 547 5046
rect 633 5033 647 5047
rect 593 5013 607 5027
rect 573 4993 587 5007
rect 513 4953 527 4967
rect 593 4893 607 4907
rect 553 4854 567 4868
rect 393 4733 407 4747
rect 373 4552 387 4566
rect 433 4554 447 4568
rect 473 4554 487 4568
rect 573 4812 587 4826
rect 553 4554 567 4568
rect 813 5374 827 5388
rect 853 5374 867 5388
rect 953 5533 967 5547
rect 933 5513 947 5527
rect 913 5373 927 5387
rect 793 5313 807 5327
rect 773 5193 787 5207
rect 673 5133 687 5147
rect 753 5133 767 5147
rect 753 5093 767 5107
rect 673 5073 687 5087
rect 713 5074 727 5088
rect 693 5032 707 5046
rect 733 5013 747 5027
rect 873 5293 887 5307
rect 833 5253 847 5267
rect 1613 5833 1627 5847
rect 1573 5793 1587 5807
rect 1353 5713 1367 5727
rect 1513 5713 1527 5727
rect 1053 5673 1067 5687
rect 1093 5653 1107 5667
rect 1193 5633 1207 5647
rect 1133 5594 1147 5608
rect 1113 5533 1127 5547
rect 1193 5594 1207 5608
rect 1273 5594 1287 5608
rect 1332 5594 1346 5608
rect 1413 5673 1427 5687
rect 1393 5633 1407 5647
rect 1353 5593 1367 5607
rect 1433 5653 1447 5667
rect 1493 5653 1507 5667
rect 1433 5594 1447 5608
rect 1473 5594 1487 5608
rect 1533 5594 1547 5608
rect 1073 5513 1087 5527
rect 1173 5513 1187 5527
rect 1053 5473 1067 5487
rect 1013 5433 1027 5447
rect 1013 5374 1027 5388
rect 933 5313 947 5327
rect 993 5313 1007 5327
rect 1093 5433 1107 5447
rect 1113 5413 1127 5427
rect 1093 5373 1107 5387
rect 1133 5374 1147 5388
rect 1173 5374 1187 5388
rect 1233 5513 1247 5527
rect 1113 5332 1127 5346
rect 1073 5313 1087 5327
rect 1133 5313 1147 5327
rect 1093 5293 1107 5307
rect 1033 5253 1047 5267
rect 913 5213 927 5227
rect 933 5193 947 5207
rect 853 5074 867 5088
rect 893 5094 907 5108
rect 893 5074 907 5088
rect 693 4993 707 5007
rect 793 4993 807 5007
rect 813 4973 827 4987
rect 693 4953 707 4967
rect 653 4873 667 4887
rect 753 4873 767 4887
rect 713 4812 727 4826
rect 673 4773 687 4787
rect 653 4593 667 4607
rect 633 4554 647 4568
rect 393 4493 407 4507
rect 373 4473 387 4487
rect 353 4433 367 4447
rect 333 4393 347 4407
rect 413 4393 427 4407
rect 233 4334 247 4348
rect 273 4334 287 4348
rect 453 4493 467 4507
rect 453 4373 467 4387
rect 433 4353 447 4367
rect 393 4292 407 4306
rect 413 4273 427 4287
rect 213 4253 227 4267
rect 253 4253 267 4267
rect 193 4073 207 4087
rect 133 4053 147 4067
rect 159 4053 173 4067
rect 93 4034 107 4048
rect 193 4034 207 4048
rect 53 3992 67 4006
rect 113 3992 127 4006
rect 73 3913 87 3927
rect 53 3893 67 3907
rect 113 3833 127 3847
rect 53 3813 67 3827
rect 293 4213 307 4227
rect 353 4133 367 4147
rect 293 4034 307 4048
rect 273 3992 287 4006
rect 173 3833 187 3847
rect 213 3953 227 3967
rect 73 3773 87 3787
rect 93 3753 107 3767
rect 133 3713 147 3727
rect 73 3653 87 3667
rect 253 3814 267 3828
rect 233 3772 247 3786
rect 173 3733 187 3747
rect 213 3733 227 3747
rect 273 3733 287 3747
rect 193 3713 207 3727
rect 153 3593 167 3607
rect 193 3514 207 3528
rect 253 3633 267 3647
rect 233 3553 247 3567
rect 73 3472 87 3486
rect 53 3353 67 3367
rect 112 3353 126 3367
rect 133 3353 147 3367
rect 93 3313 107 3327
rect 153 3333 167 3347
rect 133 3293 147 3307
rect 133 3253 147 3267
rect 113 3213 127 3227
rect 473 4293 487 4307
rect 533 4513 547 4527
rect 513 4473 527 4487
rect 573 4493 587 4507
rect 873 5013 887 5027
rect 1073 5113 1087 5127
rect 973 5093 987 5107
rect 1033 5093 1047 5107
rect 1013 5032 1027 5046
rect 1073 5032 1087 5046
rect 1013 5012 1027 5026
rect 973 4993 987 5007
rect 933 4973 947 4987
rect 1013 4973 1027 4987
rect 913 4913 927 4927
rect 833 4873 847 4887
rect 893 4854 907 4868
rect 793 4812 807 4826
rect 713 4573 727 4587
rect 753 4573 767 4587
rect 773 4553 787 4567
rect 653 4493 667 4507
rect 613 4453 627 4467
rect 713 4493 727 4507
rect 693 4433 707 4447
rect 533 4373 547 4387
rect 613 4373 627 4387
rect 533 4334 547 4348
rect 473 4213 487 4227
rect 493 4153 507 4167
rect 433 4073 447 4087
rect 413 4034 427 4048
rect 353 3893 367 3907
rect 433 3992 447 4006
rect 493 3933 507 3947
rect 413 3873 427 3887
rect 333 3814 347 3828
rect 413 3813 427 3827
rect 373 3772 387 3786
rect 393 3753 407 3767
rect 353 3693 367 3707
rect 353 3633 367 3647
rect 313 3553 327 3567
rect 273 3514 287 3528
rect 373 3472 387 3486
rect 413 3733 427 3747
rect 253 3413 267 3427
rect 313 3373 327 3387
rect 233 3353 247 3367
rect 293 3313 307 3327
rect 233 3294 247 3308
rect 173 3253 187 3267
rect 213 3213 227 3227
rect 173 3153 187 3167
rect 273 3253 287 3267
rect 153 3133 167 3147
rect 253 3133 267 3147
rect 133 3073 147 3087
rect 173 3033 187 3047
rect 273 3033 287 3047
rect 133 3014 147 3028
rect 53 2994 67 3008
rect 93 2994 107 3008
rect 133 2994 147 3008
rect 33 2953 47 2967
rect 13 2693 27 2707
rect 13 2513 27 2527
rect 113 2952 127 2966
rect 73 2913 87 2927
rect 373 3413 387 3427
rect 333 3333 347 3347
rect 373 3313 387 3327
rect 333 3294 347 3308
rect 553 4292 567 4306
rect 593 4293 607 4307
rect 673 4334 687 4348
rect 893 4813 907 4827
rect 953 4854 967 4868
rect 933 4793 947 4807
rect 993 4793 1007 4807
rect 893 4693 907 4707
rect 833 4653 847 4667
rect 873 4653 887 4667
rect 873 4573 887 4587
rect 813 4554 827 4568
rect 853 4554 867 4568
rect 1213 5333 1227 5347
rect 1193 5293 1207 5307
rect 1333 5553 1347 5567
rect 1373 5552 1387 5566
rect 1413 5552 1427 5566
rect 1253 5473 1267 5487
rect 1513 5552 1527 5566
rect 1533 5453 1547 5467
rect 1473 5413 1487 5427
rect 1513 5413 1527 5427
rect 1293 5393 1307 5407
rect 1333 5374 1347 5388
rect 1373 5374 1387 5388
rect 1413 5374 1427 5388
rect 1453 5374 1467 5388
rect 1273 5332 1287 5346
rect 1313 5332 1327 5346
rect 1153 5273 1167 5287
rect 1133 5113 1147 5127
rect 1193 5113 1207 5127
rect 1153 5032 1167 5046
rect 1473 5332 1487 5346
rect 1513 5332 1527 5346
rect 1613 5453 1627 5467
rect 1553 5373 1567 5387
rect 1593 5374 1607 5388
rect 1653 5813 1667 5827
rect 1713 5894 1727 5908
rect 1673 5693 1687 5707
rect 1653 5653 1667 5667
rect 1773 5813 1787 5827
rect 1893 6033 1907 6047
rect 1873 5894 1887 5908
rect 1973 6073 1987 6087
rect 2013 6033 2027 6047
rect 2053 6033 2067 6047
rect 1853 5813 1867 5827
rect 2013 5894 2027 5908
rect 2053 5894 2067 5908
rect 1913 5813 1927 5827
rect 1953 5813 1967 5827
rect 1993 5813 2007 5827
rect 2033 5813 2047 5827
rect 1813 5753 1827 5767
rect 1893 5753 1907 5767
rect 1853 5693 1867 5707
rect 1793 5653 1807 5667
rect 1673 5633 1687 5647
rect 1753 5633 1767 5647
rect 1713 5594 1727 5608
rect 1673 5533 1687 5547
rect 1653 5493 1667 5507
rect 1773 5594 1787 5608
rect 1813 5594 1827 5608
rect 1933 5793 1947 5807
rect 1913 5613 1927 5627
rect 1793 5513 1807 5527
rect 1753 5493 1767 5507
rect 1693 5413 1707 5427
rect 1673 5373 1687 5387
rect 1733 5374 1747 5388
rect 1313 5273 1327 5287
rect 1373 5273 1387 5287
rect 1273 5213 1287 5227
rect 1433 5213 1447 5227
rect 1233 5093 1247 5107
rect 1213 5074 1227 5088
rect 1313 5074 1327 5088
rect 1213 5032 1227 5046
rect 1193 4973 1207 4987
rect 1093 4953 1107 4967
rect 1253 4913 1267 4927
rect 1293 4913 1307 4927
rect 1373 5074 1387 5088
rect 1413 5074 1427 5088
rect 1533 5113 1547 5127
rect 1513 5093 1527 5107
rect 1453 5074 1467 5088
rect 1713 5332 1727 5346
rect 1653 5293 1667 5307
rect 1573 5193 1587 5207
rect 1333 4973 1347 4987
rect 1553 5073 1567 5087
rect 1453 4973 1467 4987
rect 1393 4953 1407 4967
rect 1033 4893 1047 4907
rect 973 4733 987 4747
rect 1013 4733 1027 4747
rect 953 4633 967 4647
rect 793 4493 807 4507
rect 933 4553 947 4567
rect 873 4512 887 4526
rect 933 4513 947 4527
rect 913 4493 927 4507
rect 813 4473 827 4487
rect 873 4473 887 4487
rect 733 4413 747 4427
rect 833 4373 847 4387
rect 893 4433 907 4447
rect 653 4292 667 4306
rect 693 4292 707 4306
rect 773 4292 787 4306
rect 873 4293 887 4307
rect 773 4193 787 4207
rect 613 4053 627 4067
rect 673 4053 687 4067
rect 553 4034 567 4048
rect 733 4034 747 4048
rect 953 4453 967 4467
rect 993 4673 1007 4687
rect 1093 4854 1107 4868
rect 1173 4854 1187 4868
rect 1073 4773 1087 4787
rect 1053 4733 1067 4747
rect 1033 4633 1047 4647
rect 1153 4773 1167 4787
rect 1213 4854 1227 4868
rect 1253 4854 1267 4868
rect 1333 4853 1347 4867
rect 1393 4854 1407 4868
rect 1453 4854 1467 4868
rect 1213 4793 1227 4807
rect 1173 4753 1187 4767
rect 1113 4713 1127 4727
rect 1073 4673 1087 4687
rect 973 4433 987 4447
rect 933 4393 947 4407
rect 953 4353 967 4367
rect 993 4353 1007 4367
rect 933 4292 947 4306
rect 1093 4613 1107 4627
rect 1273 4812 1287 4826
rect 1333 4812 1347 4826
rect 1373 4812 1387 4826
rect 1233 4773 1247 4787
rect 1213 4733 1227 4747
rect 1173 4673 1187 4687
rect 1193 4653 1207 4667
rect 1353 4693 1367 4707
rect 1213 4573 1227 4587
rect 1093 4513 1107 4527
rect 1153 4512 1167 4526
rect 1313 4554 1327 4568
rect 1333 4513 1347 4527
rect 1073 4433 1087 4447
rect 1153 4433 1167 4447
rect 1053 4393 1067 4407
rect 993 4273 1007 4287
rect 893 4173 907 4187
rect 793 4073 807 4087
rect 873 4073 887 4087
rect 773 4033 787 4047
rect 573 3992 587 4006
rect 593 3873 607 3887
rect 553 3814 567 3828
rect 493 3772 507 3786
rect 513 3653 527 3667
rect 493 3593 507 3607
rect 453 3513 467 3527
rect 513 3573 527 3587
rect 533 3514 547 3528
rect 433 3472 447 3486
rect 399 3294 413 3308
rect 353 3252 367 3266
rect 393 3252 407 3266
rect 513 3472 527 3486
rect 553 3473 567 3487
rect 533 3453 547 3467
rect 473 3333 487 3347
rect 673 3992 687 4006
rect 753 3992 767 4006
rect 713 3973 727 3987
rect 693 3953 707 3967
rect 633 3913 647 3927
rect 653 3893 667 3907
rect 633 3873 647 3887
rect 613 3773 627 3787
rect 693 3753 707 3767
rect 633 3733 647 3747
rect 853 4053 867 4067
rect 933 4053 947 4067
rect 793 3953 807 3967
rect 873 3992 887 4006
rect 913 3992 927 4006
rect 753 3893 767 3907
rect 833 3893 847 3907
rect 733 3833 747 3847
rect 873 3873 887 3887
rect 813 3814 827 3828
rect 732 3773 746 3787
rect 753 3773 767 3787
rect 713 3713 727 3727
rect 613 3693 627 3707
rect 613 3653 627 3667
rect 593 3513 607 3527
rect 633 3514 647 3528
rect 713 3514 727 3528
rect 573 3433 587 3447
rect 613 3433 627 3447
rect 653 3433 667 3447
rect 553 3413 567 3427
rect 553 3373 567 3387
rect 713 3413 727 3427
rect 513 3313 527 3327
rect 573 3333 587 3347
rect 693 3353 707 3367
rect 673 3313 687 3327
rect 573 3293 587 3307
rect 613 3293 627 3307
rect 653 3294 667 3308
rect 793 3772 807 3786
rect 833 3772 847 3786
rect 833 3752 847 3766
rect 893 3853 907 3867
rect 993 4034 1007 4048
rect 1093 4334 1107 4348
rect 1113 4273 1127 4287
rect 1053 4173 1067 4187
rect 933 3933 947 3947
rect 973 3992 987 4006
rect 993 3973 1007 3987
rect 953 3913 967 3927
rect 973 3873 987 3887
rect 953 3853 967 3867
rect 913 3813 927 3827
rect 973 3833 987 3847
rect 1013 3893 1027 3907
rect 993 3814 1007 3828
rect 893 3772 907 3786
rect 933 3772 947 3786
rect 973 3772 987 3786
rect 873 3693 887 3707
rect 873 3653 887 3667
rect 773 3514 787 3528
rect 813 3514 827 3528
rect 733 3393 747 3407
rect 733 3313 747 3327
rect 713 3293 727 3307
rect 453 3252 467 3266
rect 293 3013 307 3027
rect 193 2994 207 3008
rect 253 2994 267 3008
rect 293 2933 307 2947
rect 233 2913 247 2927
rect 193 2873 207 2887
rect 253 2873 267 2887
rect 213 2833 227 2847
rect 133 2813 147 2827
rect 173 2813 187 2827
rect 53 2773 67 2787
rect 93 2774 107 2788
rect 33 2474 47 2488
rect 153 2732 167 2746
rect 273 2833 287 2847
rect 253 2813 267 2827
rect 213 2773 227 2787
rect 333 2853 347 2867
rect 493 3153 507 3167
rect 473 3033 487 3047
rect 453 3013 467 3027
rect 433 2933 447 2947
rect 453 2893 467 2907
rect 353 2833 367 2847
rect 333 2813 347 2827
rect 293 2774 307 2788
rect 333 2773 347 2787
rect 233 2732 247 2746
rect 193 2653 207 2667
rect 113 2613 127 2627
rect 193 2613 207 2627
rect 153 2553 167 2567
rect 113 2474 127 2488
rect 53 2432 67 2446
rect 33 2353 47 2367
rect 73 2353 87 2367
rect 53 2293 67 2307
rect 133 2432 147 2446
rect 213 2573 227 2587
rect 273 2553 287 2567
rect 213 2513 227 2527
rect 233 2474 247 2488
rect 253 2432 267 2446
rect 413 2774 427 2788
rect 613 3253 627 3267
rect 593 3033 607 3047
rect 553 3013 567 3027
rect 653 3233 667 3247
rect 633 3193 647 3207
rect 573 2933 587 2947
rect 533 2893 547 2907
rect 513 2853 527 2867
rect 493 2793 507 2807
rect 353 2732 367 2746
rect 393 2732 407 2746
rect 333 2413 347 2427
rect 333 2392 347 2406
rect 293 2373 307 2387
rect 233 2293 247 2307
rect 273 2293 287 2307
rect 93 2273 107 2287
rect 133 2254 147 2268
rect 193 2252 207 2266
rect 293 2273 307 2287
rect 113 2212 127 2226
rect 173 2212 187 2226
rect 73 2033 87 2047
rect 73 1973 87 1987
rect 133 1993 147 2007
rect 53 1954 67 1968
rect 33 1912 47 1926
rect 73 1912 87 1926
rect 113 1912 127 1926
rect 53 1773 67 1787
rect 113 1773 127 1787
rect 13 1692 27 1706
rect 193 2113 207 2127
rect 253 2212 267 2226
rect 293 2212 307 2226
rect 233 2013 247 2027
rect 333 1993 347 2007
rect 273 1954 287 1968
rect 313 1953 327 1967
rect 213 1913 227 1927
rect 93 1692 107 1706
rect 133 1633 147 1647
rect 153 1434 167 1448
rect 53 1392 67 1406
rect 13 1313 27 1327
rect 133 1392 147 1406
rect 133 1353 147 1367
rect 253 1912 267 1926
rect 293 1893 307 1907
rect 213 1833 227 1847
rect 213 1773 227 1787
rect 213 1653 227 1667
rect 473 2733 487 2747
rect 413 2693 427 2707
rect 473 2553 487 2567
rect 633 2873 647 2887
rect 573 2853 587 2867
rect 593 2793 607 2807
rect 533 2733 547 2747
rect 453 2533 467 2547
rect 493 2533 507 2547
rect 513 2513 527 2527
rect 493 2473 507 2487
rect 433 2413 447 2427
rect 392 2353 406 2367
rect 413 2353 427 2367
rect 453 2313 467 2327
rect 413 2293 427 2307
rect 433 2153 447 2167
rect 613 2653 627 2667
rect 713 3073 727 3087
rect 833 3472 847 3486
rect 793 3433 807 3447
rect 1313 4473 1327 4487
rect 1293 4393 1307 4407
rect 1273 4353 1287 4367
rect 1193 4334 1207 4348
rect 1233 4334 1247 4348
rect 1193 4273 1207 4287
rect 1173 4213 1187 4227
rect 1153 4053 1167 4067
rect 1093 4034 1107 4048
rect 1133 4034 1147 4048
rect 1193 4053 1207 4067
rect 1173 4033 1187 4047
rect 1053 3973 1067 3987
rect 1153 3973 1167 3987
rect 1113 3913 1127 3927
rect 1113 3814 1127 3828
rect 1033 3733 1047 3747
rect 933 3633 947 3647
rect 1093 3772 1107 3786
rect 1173 3873 1187 3887
rect 1393 4673 1407 4687
rect 1373 4613 1387 4627
rect 1453 4813 1467 4827
rect 1413 4653 1427 4667
rect 1513 5032 1527 5046
rect 1593 5133 1607 5147
rect 1493 4893 1507 4907
rect 1553 4854 1567 4868
rect 1573 4812 1587 4826
rect 1552 4793 1566 4807
rect 1513 4733 1527 4747
rect 1573 4791 1587 4805
rect 1553 4713 1567 4727
rect 1613 4913 1627 4927
rect 1593 4713 1607 4727
rect 1713 5293 1727 5307
rect 1873 5513 1887 5527
rect 1873 5492 1887 5506
rect 1833 5413 1847 5427
rect 2033 5753 2047 5767
rect 1993 5693 2007 5707
rect 2133 6153 2147 6167
rect 2413 6233 2427 6247
rect 2473 6233 2487 6247
rect 2753 6233 2767 6247
rect 2353 6213 2367 6227
rect 2393 6193 2407 6207
rect 2213 6153 2227 6167
rect 2153 6072 2167 6086
rect 2353 6132 2367 6146
rect 2253 6114 2267 6128
rect 2313 6114 2327 6128
rect 2233 6073 2247 6087
rect 2213 5993 2227 6007
rect 2153 5933 2167 5947
rect 2253 6033 2267 6047
rect 2333 6072 2347 6086
rect 2453 6193 2467 6207
rect 2293 6033 2307 6047
rect 2392 6033 2406 6047
rect 2413 6033 2427 6047
rect 2773 6213 2787 6227
rect 2753 6193 2767 6207
rect 2613 6153 2627 6167
rect 2533 6114 2547 6128
rect 2453 6073 2467 6087
rect 2473 6053 2487 6067
rect 2773 6173 2787 6187
rect 2753 6153 2767 6167
rect 2733 6133 2747 6147
rect 2713 6114 2727 6128
rect 2933 6233 2947 6247
rect 2793 6112 2807 6126
rect 2833 6114 2847 6128
rect 2573 6053 2587 6067
rect 2273 6013 2287 6027
rect 2353 6013 2367 6027
rect 2253 5973 2267 5987
rect 2273 5953 2287 5967
rect 2193 5894 2207 5908
rect 2333 5913 2347 5927
rect 2273 5893 2287 5907
rect 2313 5894 2327 5908
rect 2133 5853 2147 5867
rect 2173 5852 2187 5866
rect 2213 5852 2227 5866
rect 2253 5852 2267 5866
rect 2293 5852 2307 5866
rect 2193 5833 2207 5847
rect 2173 5813 2187 5827
rect 2233 5812 2247 5826
rect 2193 5753 2207 5767
rect 2133 5733 2147 5747
rect 2253 5733 2267 5747
rect 2113 5713 2127 5727
rect 2093 5693 2107 5707
rect 2173 5693 2187 5707
rect 2133 5613 2147 5627
rect 2093 5594 2107 5608
rect 2053 5553 2067 5567
rect 2033 5513 2047 5527
rect 1973 5453 1987 5467
rect 1913 5413 1927 5427
rect 1953 5374 1967 5388
rect 1853 5332 1867 5346
rect 1793 5273 1807 5287
rect 1933 5273 1947 5287
rect 2013 5374 2027 5388
rect 2113 5493 2127 5507
rect 2213 5594 2227 5608
rect 2253 5594 2267 5608
rect 2573 6032 2587 6046
rect 2733 6053 2747 6067
rect 2693 6033 2707 6047
rect 2613 6013 2627 6027
rect 2533 5993 2547 6007
rect 2633 5993 2647 6007
rect 2673 5993 2687 6007
rect 2473 5953 2487 5967
rect 2413 5913 2427 5927
rect 2393 5773 2407 5787
rect 2333 5753 2347 5767
rect 2313 5713 2327 5727
rect 2353 5594 2367 5608
rect 2313 5573 2327 5587
rect 2193 5553 2207 5567
rect 2173 5473 2187 5487
rect 2293 5553 2307 5567
rect 2233 5513 2247 5527
rect 2353 5533 2367 5547
rect 2313 5493 2327 5507
rect 2233 5473 2247 5487
rect 2073 5453 2087 5467
rect 2193 5453 2207 5467
rect 2133 5413 2147 5427
rect 2173 5374 2187 5388
rect 1993 5313 2007 5327
rect 1953 5253 1967 5267
rect 1993 5253 2007 5267
rect 1753 5233 1767 5247
rect 1893 5233 1907 5247
rect 1973 5233 1987 5247
rect 1713 5173 1727 5187
rect 1712 5113 1726 5127
rect 1733 5113 1747 5127
rect 1933 5113 1947 5127
rect 1713 5074 1727 5088
rect 1693 4953 1707 4967
rect 1773 5074 1787 5088
rect 1813 5074 1827 5088
rect 1853 5074 1867 5088
rect 1893 5074 1907 5088
rect 1753 5013 1767 5027
rect 1793 5013 1807 5027
rect 1733 4973 1747 4987
rect 1713 4893 1727 4907
rect 1713 4872 1727 4886
rect 1673 4854 1687 4868
rect 1633 4813 1647 4827
rect 1693 4812 1707 4826
rect 1733 4813 1747 4827
rect 1633 4773 1647 4787
rect 1613 4693 1627 4707
rect 1573 4653 1587 4667
rect 1613 4653 1627 4667
rect 1513 4613 1527 4627
rect 1413 4553 1427 4567
rect 1453 4553 1467 4567
rect 1393 4513 1407 4527
rect 1433 4512 1447 4526
rect 1573 4573 1587 4587
rect 1593 4553 1607 4567
rect 1693 4713 1707 4727
rect 1793 4854 1807 4868
rect 1973 5073 1987 5087
rect 1953 5032 1967 5046
rect 1913 5013 1927 5027
rect 1893 4854 1907 4868
rect 1933 4854 1947 4868
rect 1773 4813 1787 4827
rect 1813 4812 1827 4826
rect 1853 4813 1867 4827
rect 1953 4812 1967 4826
rect 1772 4773 1786 4787
rect 1793 4772 1807 4786
rect 1653 4653 1667 4667
rect 1673 4613 1687 4627
rect 1653 4553 1667 4567
rect 1713 4673 1727 4687
rect 1713 4613 1727 4627
rect 1753 4593 1767 4607
rect 1753 4553 1767 4567
rect 1513 4513 1527 4527
rect 1433 4490 1447 4504
rect 1372 4473 1386 4487
rect 1393 4473 1407 4487
rect 1333 4393 1347 4407
rect 1413 4453 1427 4467
rect 1433 4333 1447 4347
rect 1473 4473 1487 4487
rect 1513 4473 1527 4487
rect 1333 4293 1347 4307
rect 1333 4173 1347 4187
rect 1433 4173 1447 4187
rect 1313 4153 1327 4167
rect 1373 4113 1387 4127
rect 1353 4053 1367 4067
rect 1253 4034 1267 4048
rect 1293 4034 1307 4048
rect 1333 4034 1347 4048
rect 1213 3993 1227 4007
rect 1273 3992 1287 4006
rect 1413 4053 1427 4067
rect 1573 4512 1587 4526
rect 1633 4513 1647 4527
rect 1573 4453 1587 4467
rect 1533 4413 1547 4427
rect 1513 4353 1527 4367
rect 1533 4334 1547 4348
rect 1553 4293 1567 4307
rect 1533 4273 1547 4287
rect 1553 4273 1567 4287
rect 1593 4253 1607 4267
rect 1513 4213 1527 4227
rect 1473 4133 1487 4147
rect 1593 4193 1607 4207
rect 1593 4153 1607 4167
rect 1693 4512 1707 4526
rect 1633 4413 1647 4427
rect 1773 4513 1787 4527
rect 1733 4353 1747 4367
rect 1673 4334 1687 4348
rect 1713 4334 1727 4348
rect 2133 5253 2147 5267
rect 2033 5193 2047 5207
rect 2033 5074 2047 5088
rect 2073 5074 2087 5088
rect 2193 5333 2207 5347
rect 2293 5433 2307 5447
rect 2193 5313 2207 5327
rect 2233 5313 2247 5327
rect 2293 5313 2307 5327
rect 2172 5273 2186 5287
rect 2193 5273 2207 5287
rect 2153 5193 2167 5207
rect 2193 5153 2207 5167
rect 2233 5133 2247 5147
rect 2193 5093 2207 5107
rect 2213 5074 2227 5088
rect 2253 5074 2267 5088
rect 2033 5013 2047 5027
rect 2112 5033 2126 5047
rect 2133 5033 2147 5047
rect 2113 4993 2127 5007
rect 2093 4953 2107 4967
rect 2133 4933 2147 4947
rect 2053 4913 2067 4927
rect 2092 4913 2106 4927
rect 2113 4913 2127 4927
rect 2073 4893 2087 4907
rect 2093 4873 2107 4887
rect 2013 4853 2027 4867
rect 2073 4854 2087 4868
rect 2113 4853 2127 4867
rect 2093 4812 2107 4826
rect 2053 4793 2067 4807
rect 2133 4793 2147 4807
rect 1992 4773 2006 4787
rect 2013 4773 2027 4787
rect 1872 4753 1886 4767
rect 1893 4753 1907 4767
rect 1973 4753 1987 4767
rect 1873 4673 1887 4687
rect 1993 4733 2007 4747
rect 1913 4713 1927 4727
rect 1793 4493 1807 4507
rect 1793 4472 1807 4486
rect 1773 4413 1787 4427
rect 1673 4273 1687 4287
rect 1733 4292 1747 4306
rect 1733 4272 1747 4286
rect 1673 4233 1687 4247
rect 1733 4233 1747 4247
rect 1653 4213 1667 4227
rect 1713 4213 1727 4227
rect 1693 4153 1707 4167
rect 1593 4113 1607 4127
rect 1633 4113 1647 4127
rect 1493 4073 1507 4087
rect 1553 4076 1567 4090
rect 1473 4033 1487 4047
rect 1633 4072 1647 4086
rect 1593 4053 1607 4067
rect 1553 4033 1567 4047
rect 1633 4034 1647 4048
rect 1453 4013 1467 4027
rect 1573 4013 1587 4027
rect 1613 4013 1627 4027
rect 1233 3913 1247 3927
rect 1213 3873 1227 3887
rect 1333 3973 1347 3987
rect 1313 3953 1327 3967
rect 1253 3873 1267 3887
rect 1293 3873 1307 3887
rect 1233 3853 1247 3867
rect 1233 3814 1247 3828
rect 1193 3793 1207 3807
rect 1173 3773 1187 3787
rect 1213 3772 1227 3786
rect 1173 3733 1187 3747
rect 1213 3733 1227 3747
rect 1073 3653 1087 3667
rect 1153 3653 1167 3667
rect 1053 3593 1067 3607
rect 893 3514 907 3528
rect 953 3514 967 3528
rect 993 3514 1007 3528
rect 1033 3514 1047 3528
rect 833 3413 847 3427
rect 873 3413 887 3427
rect 793 3353 807 3367
rect 753 3294 767 3308
rect 973 3472 987 3486
rect 1153 3573 1167 3587
rect 1113 3514 1127 3528
rect 1213 3693 1227 3707
rect 1273 3693 1287 3707
rect 1253 3613 1267 3627
rect 1333 3933 1347 3947
rect 1393 3973 1407 3987
rect 1453 3953 1467 3967
rect 1573 3973 1587 3987
rect 1513 3893 1527 3907
rect 1573 3873 1587 3887
rect 1533 3853 1547 3867
rect 1593 3853 1607 3867
rect 1393 3814 1407 3828
rect 1573 3814 1587 3828
rect 1373 3772 1387 3786
rect 1413 3772 1427 3786
rect 1333 3713 1347 3727
rect 1313 3673 1327 3687
rect 1293 3633 1307 3647
rect 1273 3593 1287 3607
rect 1253 3532 1267 3546
rect 1213 3514 1227 3528
rect 953 3353 967 3367
rect 1053 3433 1067 3447
rect 1013 3393 1027 3407
rect 953 3313 967 3327
rect 853 3252 867 3266
rect 753 3193 767 3207
rect 793 3193 807 3207
rect 733 3013 747 3027
rect 753 2994 767 3008
rect 693 2933 707 2947
rect 673 2913 687 2927
rect 673 2813 687 2827
rect 653 2633 667 2647
rect 733 2813 747 2827
rect 733 2792 747 2806
rect 693 2693 707 2707
rect 673 2613 687 2627
rect 773 2732 787 2746
rect 713 2573 727 2587
rect 733 2513 747 2527
rect 533 2473 547 2487
rect 653 2474 667 2488
rect 693 2474 707 2488
rect 613 2432 627 2446
rect 573 2413 587 2427
rect 513 2393 527 2407
rect 713 2432 727 2446
rect 813 3093 827 3107
rect 933 3294 947 3308
rect 953 3252 967 3266
rect 913 3233 927 3247
rect 893 3033 907 3047
rect 833 2994 847 3008
rect 853 2952 867 2966
rect 893 2913 907 2927
rect 833 2873 847 2887
rect 813 2813 827 2827
rect 813 2732 827 2746
rect 1093 3353 1107 3367
rect 1153 3393 1167 3407
rect 1133 3333 1147 3347
rect 1013 3033 1027 3047
rect 953 2994 967 3008
rect 993 2994 1007 3008
rect 1073 3252 1087 3266
rect 1113 3193 1127 3207
rect 1133 3173 1147 3187
rect 1073 3013 1087 3027
rect 1053 2994 1067 3008
rect 913 2853 927 2867
rect 893 2774 907 2788
rect 973 2952 987 2966
rect 953 2873 967 2887
rect 953 2813 967 2827
rect 933 2773 947 2787
rect 1053 2913 1067 2927
rect 1033 2833 1047 2847
rect 1013 2793 1027 2807
rect 973 2773 987 2787
rect 1233 3472 1247 3486
rect 1273 3473 1287 3487
rect 1193 3433 1207 3447
rect 1253 3433 1267 3447
rect 1253 3373 1267 3387
rect 1212 3333 1226 3347
rect 1233 3333 1247 3347
rect 1193 3294 1207 3308
rect 1273 3293 1287 3307
rect 1253 3252 1267 3266
rect 1333 3613 1347 3627
rect 1393 3753 1407 3767
rect 1433 3753 1447 3767
rect 1553 3753 1567 3767
rect 1593 3733 1607 3747
rect 1553 3713 1567 3727
rect 1513 3693 1527 3707
rect 1513 3672 1527 3686
rect 1453 3653 1467 3667
rect 1373 3573 1387 3587
rect 1313 3533 1327 3547
rect 1393 3534 1407 3548
rect 1373 3514 1387 3528
rect 1413 3513 1427 3527
rect 1333 3473 1347 3487
rect 1313 3413 1327 3427
rect 1433 3473 1447 3487
rect 1393 3433 1407 3447
rect 1353 3413 1367 3427
rect 1353 3373 1367 3387
rect 1333 3313 1347 3327
rect 1473 3593 1487 3607
rect 1453 3433 1467 3447
rect 1433 3333 1447 3347
rect 1493 3573 1507 3587
rect 1513 3533 1527 3547
rect 1573 3693 1587 3707
rect 1593 3653 1607 3667
rect 1573 3593 1587 3607
rect 1833 4493 1847 4507
rect 1813 4393 1827 4407
rect 1893 4493 1907 4507
rect 1873 4413 1887 4427
rect 1833 4353 1847 4367
rect 1853 4334 1867 4348
rect 1953 4693 1967 4707
rect 1933 4633 1947 4647
rect 1933 4533 1947 4547
rect 1913 4413 1927 4427
rect 1913 4353 1927 4367
rect 1813 4273 1827 4287
rect 1793 4213 1807 4227
rect 1833 4233 1847 4247
rect 1813 4193 1827 4207
rect 1773 4173 1787 4187
rect 1773 4152 1787 4166
rect 1772 4113 1786 4127
rect 1793 4113 1807 4127
rect 1833 4093 1847 4107
rect 1793 4053 1807 4067
rect 1753 4034 1767 4048
rect 1893 4293 1907 4307
rect 2033 4653 2047 4667
rect 2093 4653 2107 4667
rect 2073 4613 2087 4627
rect 2033 4554 2047 4568
rect 2013 4512 2027 4526
rect 1953 4493 1967 4507
rect 2013 4473 2027 4487
rect 1953 4453 1967 4467
rect 1993 4453 2007 4467
rect 1933 4333 1947 4347
rect 2053 4413 2067 4427
rect 2013 4373 2027 4387
rect 2133 4613 2147 4627
rect 2092 4593 2106 4607
rect 2113 4592 2127 4606
rect 2093 4554 2107 4568
rect 2193 5032 2207 5046
rect 2233 5032 2247 5046
rect 2273 5033 2287 5047
rect 2253 5013 2267 5027
rect 2213 4993 2227 5007
rect 2193 4893 2207 4907
rect 2232 4933 2246 4947
rect 2253 4933 2267 4947
rect 2233 4793 2247 4807
rect 2193 4773 2207 4787
rect 2153 4573 2167 4587
rect 2233 4573 2247 4587
rect 2173 4554 2187 4568
rect 2093 4413 2107 4427
rect 2153 4512 2167 4526
rect 2213 4513 2227 4527
rect 2133 4473 2147 4487
rect 2112 4393 2126 4407
rect 2133 4393 2147 4407
rect 2073 4353 2087 4367
rect 2193 4493 2207 4507
rect 2213 4473 2227 4487
rect 2373 5513 2387 5527
rect 2453 5813 2467 5827
rect 2433 5713 2447 5727
rect 2453 5693 2467 5707
rect 2433 5673 2447 5687
rect 2433 5652 2447 5666
rect 2413 5473 2427 5487
rect 2553 5894 2567 5908
rect 2593 5894 2607 5908
rect 2673 5953 2687 5967
rect 2773 5953 2787 5967
rect 2693 5894 2707 5908
rect 2733 5894 2747 5908
rect 2853 6053 2867 6067
rect 2893 6053 2907 6067
rect 2793 5933 2807 5947
rect 2693 5833 2707 5847
rect 2733 5833 2747 5847
rect 2673 5813 2687 5827
rect 2793 5813 2807 5827
rect 2753 5793 2767 5807
rect 2733 5753 2747 5767
rect 2713 5713 2727 5727
rect 2533 5693 2547 5707
rect 2653 5693 2667 5707
rect 2473 5594 2487 5608
rect 2513 5594 2527 5608
rect 2573 5594 2587 5608
rect 2493 5552 2507 5566
rect 2453 5533 2467 5547
rect 2533 5533 2547 5547
rect 2433 5433 2447 5447
rect 2513 5473 2527 5487
rect 2473 5453 2487 5467
rect 2453 5413 2467 5427
rect 2373 5374 2387 5388
rect 2433 5374 2447 5388
rect 2353 5273 2367 5287
rect 2313 5253 2327 5267
rect 2353 5233 2367 5247
rect 2313 5213 2327 5227
rect 2333 5193 2347 5207
rect 2313 5093 2327 5107
rect 2413 5332 2427 5346
rect 2453 5313 2467 5327
rect 2673 5552 2687 5566
rect 2713 5552 2727 5566
rect 2633 5533 2647 5547
rect 2573 5413 2587 5427
rect 2593 5374 2607 5388
rect 2673 5513 2687 5527
rect 2673 5433 2687 5447
rect 2573 5332 2587 5346
rect 2433 5253 2447 5267
rect 2513 5253 2527 5267
rect 2413 5213 2427 5227
rect 2393 5193 2407 5207
rect 2373 5173 2387 5187
rect 2413 5153 2427 5167
rect 2313 5033 2327 5047
rect 2352 5013 2366 5027
rect 2373 5013 2387 5027
rect 2333 4893 2347 4907
rect 2313 4873 2327 4887
rect 2413 4993 2427 5007
rect 2393 4973 2407 4987
rect 2393 4933 2407 4947
rect 2373 4854 2387 4868
rect 2413 4853 2427 4867
rect 2313 4813 2327 4827
rect 2393 4812 2407 4826
rect 2373 4793 2387 4807
rect 2353 4773 2367 4787
rect 2313 4753 2327 4767
rect 2313 4732 2327 4746
rect 2293 4713 2307 4727
rect 2292 4692 2306 4706
rect 2313 4693 2327 4707
rect 2253 4553 2267 4567
rect 2293 4553 2307 4567
rect 2273 4512 2287 4526
rect 2313 4512 2327 4526
rect 2233 4453 2247 4467
rect 2213 4413 2227 4427
rect 2193 4393 2207 4407
rect 2173 4353 2187 4367
rect 2053 4313 2067 4327
rect 1873 4213 1887 4227
rect 1873 4153 1887 4167
rect 1853 4073 1867 4087
rect 1733 3993 1747 4007
rect 1653 3933 1667 3947
rect 1673 3913 1687 3927
rect 1673 3853 1687 3867
rect 1633 3653 1647 3667
rect 1873 4033 1887 4047
rect 1813 3992 1827 4006
rect 1853 3992 1867 4006
rect 1833 3973 1847 3987
rect 1753 3773 1767 3787
rect 1793 3772 1807 3786
rect 1733 3733 1747 3747
rect 1733 3673 1747 3687
rect 1693 3653 1707 3667
rect 1673 3593 1687 3607
rect 1613 3553 1627 3567
rect 1533 3472 1547 3486
rect 1573 3473 1587 3487
rect 1513 3433 1527 3447
rect 1493 3413 1507 3427
rect 1373 3313 1387 3327
rect 1453 3312 1467 3326
rect 1473 3313 1487 3327
rect 1513 3373 1527 3387
rect 1653 3533 1667 3547
rect 1693 3533 1707 3547
rect 1613 3453 1627 3467
rect 1553 3333 1567 3347
rect 1213 3193 1227 3207
rect 1173 3153 1187 3167
rect 1233 3153 1247 3167
rect 1173 3113 1187 3127
rect 1153 3093 1167 3107
rect 1173 2994 1187 3008
rect 1093 2893 1107 2907
rect 1073 2813 1087 2827
rect 1073 2774 1087 2788
rect 1133 2933 1147 2947
rect 1113 2873 1127 2887
rect 1113 2813 1127 2827
rect 873 2732 887 2746
rect 913 2732 927 2746
rect 953 2732 967 2746
rect 853 2693 867 2707
rect 833 2553 847 2567
rect 1013 2732 1027 2746
rect 1093 2733 1107 2747
rect 933 2633 947 2647
rect 973 2633 987 2647
rect 873 2513 887 2527
rect 853 2493 867 2507
rect 833 2474 847 2488
rect 953 2474 967 2488
rect 1093 2573 1107 2587
rect 1193 2952 1207 2966
rect 1153 2853 1167 2867
rect 1153 2774 1167 2788
rect 1333 3252 1347 3266
rect 1373 3253 1387 3267
rect 1353 3173 1367 3187
rect 1293 3153 1307 3167
rect 1273 3013 1287 3027
rect 1353 3133 1367 3147
rect 1333 3113 1347 3127
rect 1353 3093 1367 3107
rect 1333 2994 1347 3008
rect 1273 2933 1287 2947
rect 1453 3193 1467 3207
rect 1593 3294 1607 3308
rect 1653 3453 1667 3467
rect 1533 3253 1547 3267
rect 1393 3153 1407 3167
rect 1513 3153 1527 3167
rect 1373 2933 1387 2947
rect 1513 3132 1527 3146
rect 1433 3033 1447 3047
rect 1473 2994 1487 3008
rect 1573 3252 1587 3266
rect 1673 3413 1687 3427
rect 1672 3294 1686 3308
rect 1713 3433 1727 3447
rect 1793 3752 1807 3766
rect 1773 3613 1787 3627
rect 1913 4193 1927 4207
rect 1853 3953 1867 3967
rect 1893 3953 1907 3967
rect 1973 4292 1987 4306
rect 1973 4253 1987 4267
rect 2033 4233 2047 4247
rect 2053 4193 2067 4207
rect 2033 4173 2047 4187
rect 2013 4113 2027 4127
rect 1953 4073 1967 4087
rect 2013 4034 2027 4048
rect 1933 3973 1947 3987
rect 1973 3913 1987 3927
rect 1913 3853 1927 3867
rect 1913 3832 1927 3846
rect 1953 3814 1967 3828
rect 2013 3973 2027 3987
rect 1993 3873 2007 3887
rect 2153 4334 2167 4348
rect 2173 4292 2187 4306
rect 2133 4233 2147 4247
rect 2093 4213 2107 4227
rect 2073 4153 2087 4167
rect 2133 4212 2147 4226
rect 2093 4133 2107 4147
rect 2053 4073 2067 4087
rect 2033 3953 2047 3967
rect 2093 4034 2107 4048
rect 2173 4113 2187 4127
rect 2113 3953 2127 3967
rect 2053 3913 2067 3927
rect 2293 4473 2307 4487
rect 2393 4753 2407 4767
rect 2613 5313 2627 5327
rect 2513 5232 2527 5246
rect 2573 5233 2587 5247
rect 2493 5133 2507 5147
rect 2493 5093 2507 5107
rect 2653 5113 2667 5127
rect 2553 5074 2567 5088
rect 2593 5074 2607 5088
rect 3193 6213 3207 6227
rect 3413 6213 3427 6227
rect 3713 6213 3727 6227
rect 2953 6193 2967 6207
rect 3053 6193 3067 6207
rect 3013 6114 3027 6128
rect 3093 6153 3107 6167
rect 3173 6153 3187 6167
rect 2993 6033 3007 6047
rect 2953 5993 2967 6007
rect 2933 5953 2947 5967
rect 2893 5933 2907 5947
rect 2953 5933 2967 5947
rect 3153 6114 3167 6128
rect 3213 6173 3227 6187
rect 3273 6173 3287 6187
rect 3393 6173 3407 6187
rect 3233 6152 3247 6166
rect 3133 6072 3147 6086
rect 3093 6053 3107 6067
rect 3093 6032 3107 6046
rect 2893 5894 2907 5908
rect 2953 5893 2967 5907
rect 2993 5894 3007 5908
rect 3033 5894 3047 5908
rect 2913 5793 2927 5807
rect 2853 5713 2867 5727
rect 3013 5852 3027 5866
rect 3053 5852 3067 5866
rect 3253 6113 3267 6127
rect 3293 6113 3307 6127
rect 3333 6114 3347 6128
rect 3233 5973 3247 5987
rect 3273 6073 3287 6087
rect 3253 5953 3267 5967
rect 3113 5933 3127 5947
rect 3173 5894 3187 5908
rect 3093 5813 3107 5827
rect 3113 5793 3127 5807
rect 3013 5653 3027 5667
rect 2933 5594 2947 5608
rect 3153 5852 3167 5866
rect 3193 5793 3207 5807
rect 3153 5713 3167 5727
rect 3133 5673 3147 5687
rect 3193 5693 3207 5707
rect 3173 5633 3187 5647
rect 3313 6053 3327 6067
rect 3313 6013 3327 6027
rect 3393 6114 3407 6128
rect 3513 6173 3527 6187
rect 3473 6153 3487 6167
rect 3433 6114 3447 6128
rect 3473 6114 3487 6128
rect 3393 6073 3407 6087
rect 3373 6013 3387 6027
rect 3333 5993 3347 6007
rect 3353 5973 3367 5987
rect 3313 5914 3327 5928
rect 3292 5893 3306 5907
rect 3333 5852 3347 5866
rect 3373 5852 3387 5866
rect 3713 6153 3727 6167
rect 3613 6133 3627 6147
rect 3573 6114 3587 6128
rect 3793 6114 3807 6128
rect 5693 6233 5707 6247
rect 5753 6233 5767 6247
rect 4493 6213 4507 6227
rect 4973 6213 4987 6227
rect 5613 6213 5627 6227
rect 4033 6173 4047 6187
rect 4313 6173 4327 6187
rect 3513 6013 3527 6027
rect 3633 6073 3647 6087
rect 3593 6053 3607 6067
rect 3693 6072 3707 6086
rect 3733 6072 3747 6086
rect 3833 6114 3847 6128
rect 3633 6033 3647 6047
rect 3733 6033 3747 6047
rect 3793 6033 3807 6047
rect 3553 5993 3567 6007
rect 3853 6072 3867 6086
rect 3893 6053 3907 6067
rect 3873 6033 3887 6047
rect 3552 5972 3566 5986
rect 3573 5973 3587 5987
rect 3633 5973 3647 5987
rect 3813 5973 3827 5987
rect 3853 5973 3867 5987
rect 3453 5933 3467 5947
rect 3473 5894 3487 5908
rect 3513 5894 3527 5908
rect 3333 5813 3347 5827
rect 3273 5753 3287 5767
rect 3353 5693 3367 5707
rect 3333 5653 3347 5667
rect 3193 5593 3207 5607
rect 3293 5594 3307 5608
rect 3333 5594 3347 5608
rect 3493 5852 3507 5866
rect 3533 5852 3547 5866
rect 3453 5813 3467 5827
rect 3433 5793 3447 5807
rect 3433 5753 3447 5767
rect 3473 5753 3487 5767
rect 3453 5713 3467 5727
rect 3412 5673 3426 5687
rect 3433 5673 3447 5687
rect 3373 5633 3387 5647
rect 3413 5594 3427 5608
rect 3713 5933 3727 5947
rect 3653 5913 3667 5927
rect 3673 5894 3687 5908
rect 3613 5852 3627 5866
rect 3653 5852 3667 5866
rect 3693 5853 3707 5867
rect 3613 5832 3627 5846
rect 3653 5831 3667 5845
rect 3593 5713 3607 5727
rect 3533 5673 3547 5687
rect 3573 5673 3587 5687
rect 3553 5653 3567 5667
rect 3633 5653 3647 5667
rect 3633 5613 3647 5627
rect 3493 5594 3507 5608
rect 3533 5594 3547 5608
rect 3353 5573 3367 5587
rect 2913 5552 2927 5566
rect 2893 5473 2907 5487
rect 2773 5373 2787 5387
rect 2813 5373 2827 5387
rect 2853 5374 2867 5388
rect 2993 5552 3007 5566
rect 3093 5552 3107 5566
rect 3133 5552 3147 5566
rect 3213 5552 3227 5566
rect 3213 5493 3227 5507
rect 2913 5374 2927 5388
rect 2713 5332 2727 5346
rect 2753 5332 2767 5346
rect 2813 5332 2827 5346
rect 2673 5093 2687 5107
rect 2493 5032 2507 5046
rect 2533 5013 2547 5027
rect 2593 4993 2607 5007
rect 2473 4973 2487 4987
rect 2673 5032 2687 5046
rect 2673 4993 2687 5007
rect 2633 4953 2647 4967
rect 2593 4893 2607 4907
rect 2513 4854 2527 4868
rect 2573 4854 2587 4868
rect 2453 4773 2467 4787
rect 2433 4574 2447 4588
rect 2633 4854 2647 4868
rect 2713 4953 2727 4967
rect 2493 4733 2507 4747
rect 2573 4733 2587 4747
rect 2533 4713 2547 4727
rect 2513 4613 2527 4627
rect 2473 4573 2487 4587
rect 2433 4553 2447 4567
rect 2513 4553 2527 4567
rect 2393 4513 2407 4527
rect 2353 4453 2367 4467
rect 2333 4433 2347 4447
rect 2353 4413 2367 4427
rect 2233 4333 2247 4347
rect 2293 4334 2307 4348
rect 2493 4512 2507 4526
rect 2453 4473 2467 4487
rect 2513 4473 2527 4487
rect 2613 4812 2627 4826
rect 2753 5113 2767 5127
rect 2873 5332 2887 5346
rect 2913 5332 2927 5346
rect 2813 5093 2827 5107
rect 2893 5193 2907 5207
rect 2873 5153 2887 5167
rect 2773 4993 2787 5007
rect 2873 4993 2887 5007
rect 2833 4973 2847 4987
rect 2873 4972 2887 4986
rect 2813 4953 2827 4967
rect 2753 4893 2767 4907
rect 2853 4933 2867 4947
rect 2753 4872 2767 4886
rect 2813 4873 2827 4887
rect 2733 4853 2747 4867
rect 2713 4793 2727 4807
rect 2632 4773 2646 4787
rect 2653 4773 2667 4787
rect 2613 4753 2627 4767
rect 2612 4732 2626 4746
rect 2633 4733 2647 4747
rect 2553 4573 2567 4587
rect 2593 4573 2607 4587
rect 2633 4653 2647 4667
rect 2693 4693 2707 4707
rect 2693 4633 2707 4647
rect 2773 4812 2787 4826
rect 2873 4773 2887 4787
rect 3093 5413 3107 5427
rect 3173 5413 3187 5427
rect 2953 5393 2967 5407
rect 3033 5374 3047 5388
rect 2953 5353 2967 5367
rect 3113 5374 3127 5388
rect 3313 5552 3327 5566
rect 3393 5552 3407 5566
rect 3433 5552 3447 5566
rect 3393 5413 3407 5427
rect 3313 5393 3327 5407
rect 3013 5332 3027 5346
rect 3093 5333 3107 5347
rect 3053 5273 3067 5287
rect 3193 5332 3207 5346
rect 3153 5273 3167 5287
rect 3153 5252 3167 5266
rect 3193 5253 3207 5267
rect 3113 5153 3127 5167
rect 2993 5133 3007 5147
rect 2933 5073 2947 5087
rect 3013 5074 3027 5088
rect 2953 5032 2967 5046
rect 3033 5033 3047 5047
rect 2993 4913 3007 4927
rect 2913 4873 2927 4887
rect 2933 4854 2947 4868
rect 2973 4854 2987 4868
rect 2933 4753 2947 4767
rect 2853 4733 2867 4747
rect 2893 4733 2907 4747
rect 2793 4713 2807 4727
rect 2733 4673 2747 4687
rect 2713 4592 2727 4606
rect 2653 4573 2667 4587
rect 2892 4693 2906 4707
rect 2913 4693 2927 4707
rect 2893 4613 2907 4627
rect 2853 4593 2867 4607
rect 2753 4554 2767 4568
rect 2793 4554 2807 4568
rect 2833 4554 2847 4568
rect 2593 4513 2607 4527
rect 2653 4513 2667 4527
rect 2733 4512 2747 4526
rect 2773 4513 2787 4527
rect 2553 4493 2567 4507
rect 2593 4493 2607 4507
rect 2473 4453 2487 4467
rect 2533 4453 2547 4467
rect 2393 4413 2407 4427
rect 2373 4332 2387 4346
rect 2433 4334 2447 4348
rect 2233 4292 2247 4306
rect 2213 4113 2227 4127
rect 2273 4292 2287 4306
rect 2313 4173 2327 4187
rect 2492 4413 2506 4427
rect 2513 4413 2527 4427
rect 2693 4473 2707 4487
rect 2713 4453 2727 4467
rect 2613 4433 2627 4447
rect 2693 4433 2707 4447
rect 2593 4413 2607 4427
rect 2553 4373 2567 4387
rect 2613 4393 2627 4407
rect 2773 4413 2787 4427
rect 2632 4372 2646 4386
rect 2653 4373 2667 4387
rect 2713 4373 2727 4387
rect 2753 4373 2767 4387
rect 2513 4334 2527 4348
rect 2553 4334 2567 4348
rect 2593 4334 2607 4348
rect 2413 4253 2427 4267
rect 2372 4133 2386 4147
rect 2393 4133 2407 4147
rect 2313 4093 2327 4107
rect 2253 4034 2267 4048
rect 2193 3933 2207 3947
rect 2173 3873 2187 3887
rect 2133 3853 2147 3867
rect 1893 3772 1907 3786
rect 1933 3753 1947 3767
rect 1873 3713 1887 3727
rect 1852 3673 1866 3687
rect 1873 3673 1887 3687
rect 1953 3633 1967 3647
rect 1933 3553 1947 3567
rect 2013 3812 2027 3826
rect 2073 3814 2087 3828
rect 2013 3773 2027 3787
rect 2053 3772 2067 3786
rect 2113 3772 2127 3786
rect 1993 3553 2007 3567
rect 1773 3533 1787 3547
rect 1833 3513 1847 3527
rect 1953 3513 1967 3527
rect 1773 3473 1787 3487
rect 1813 3472 1827 3486
rect 1872 3473 1886 3487
rect 1893 3473 1907 3487
rect 1613 3213 1627 3227
rect 1573 3173 1587 3187
rect 1533 3053 1547 3067
rect 1573 3033 1587 3047
rect 1533 3013 1547 3027
rect 1393 2913 1407 2927
rect 1513 2953 1527 2967
rect 1653 3093 1667 3107
rect 1612 3013 1626 3027
rect 1633 3013 1647 3027
rect 1593 2952 1607 2966
rect 1553 2933 1567 2947
rect 1613 2933 1627 2947
rect 1512 2913 1526 2927
rect 1533 2913 1547 2927
rect 1453 2893 1467 2907
rect 1333 2873 1347 2887
rect 1313 2853 1327 2867
rect 1233 2774 1247 2788
rect 1133 2733 1147 2747
rect 1253 2733 1267 2747
rect 1213 2693 1227 2707
rect 1173 2673 1187 2687
rect 1173 2633 1187 2647
rect 733 2413 747 2427
rect 653 2373 667 2387
rect 613 2353 627 2367
rect 553 2313 567 2327
rect 693 2313 707 2327
rect 593 2254 607 2268
rect 633 2253 647 2267
rect 753 2393 767 2407
rect 733 2273 747 2287
rect 573 2193 587 2207
rect 533 2113 547 2127
rect 433 2013 447 2027
rect 393 1993 407 2007
rect 513 1993 527 2007
rect 453 1912 467 1926
rect 493 1913 507 1927
rect 533 1953 547 1967
rect 613 1954 627 1968
rect 673 2212 687 2226
rect 713 2212 727 2226
rect 673 2192 687 2206
rect 713 2113 727 2127
rect 893 2432 907 2446
rect 933 2433 947 2447
rect 893 2293 907 2307
rect 853 2273 867 2287
rect 813 2193 827 2207
rect 873 2153 887 2167
rect 853 2113 867 2127
rect 773 2073 787 2087
rect 673 2053 687 2067
rect 753 2053 767 2067
rect 533 1913 547 1927
rect 513 1893 527 1907
rect 413 1833 427 1847
rect 473 1813 487 1827
rect 433 1773 447 1787
rect 333 1673 347 1687
rect 253 1633 267 1647
rect 233 1434 247 1448
rect 333 1434 347 1448
rect 413 1692 427 1706
rect 373 1673 387 1687
rect 553 1893 567 1907
rect 853 2033 867 2047
rect 733 1993 747 2007
rect 1013 2474 1027 2488
rect 1053 2474 1067 2488
rect 953 2393 967 2407
rect 953 2212 967 2226
rect 1033 2432 1047 2446
rect 1073 2433 1087 2447
rect 1013 2373 1027 2387
rect 993 2153 1007 2167
rect 933 2073 947 2087
rect 833 1973 847 1987
rect 893 1973 907 1987
rect 813 1953 827 1967
rect 673 1912 687 1926
rect 653 1893 667 1907
rect 593 1813 607 1827
rect 693 1813 707 1827
rect 533 1773 547 1787
rect 613 1773 627 1787
rect 513 1734 527 1748
rect 553 1734 567 1748
rect 473 1613 487 1627
rect 493 1553 507 1567
rect 473 1533 487 1547
rect 393 1513 407 1527
rect 433 1473 447 1487
rect 273 1373 287 1387
rect 253 1353 267 1367
rect 153 1273 167 1287
rect 113 1253 127 1267
rect 53 1233 67 1247
rect 93 1233 107 1247
rect 233 1313 247 1327
rect 213 1273 227 1287
rect 193 1253 207 1267
rect 173 1213 187 1227
rect 53 1172 67 1186
rect 93 1172 107 1186
rect 173 1173 187 1187
rect 133 1133 147 1147
rect 133 933 147 947
rect 33 913 47 927
rect 93 914 107 928
rect 73 872 87 886
rect 33 813 47 827
rect 233 1233 247 1247
rect 213 1213 227 1227
rect 333 1393 347 1407
rect 373 1392 387 1406
rect 413 1392 427 1406
rect 313 1373 327 1387
rect 593 1693 607 1707
rect 593 1553 607 1567
rect 573 1513 587 1527
rect 533 1453 547 1467
rect 653 1734 667 1748
rect 753 1912 767 1926
rect 753 1873 767 1887
rect 713 1793 727 1807
rect 713 1673 727 1687
rect 653 1653 667 1667
rect 633 1513 647 1527
rect 613 1433 627 1447
rect 493 1392 507 1406
rect 353 1333 367 1347
rect 473 1333 487 1347
rect 293 1293 307 1307
rect 273 1253 287 1267
rect 293 1233 307 1247
rect 493 1293 507 1307
rect 473 1273 487 1287
rect 413 1253 427 1267
rect 353 1233 367 1247
rect 313 1213 327 1227
rect 373 1214 387 1228
rect 273 1172 287 1186
rect 313 1173 327 1187
rect 193 933 207 947
rect 233 933 247 947
rect 253 914 267 928
rect 113 853 127 867
rect 152 853 166 867
rect 173 853 187 867
rect 213 853 227 867
rect 153 773 167 787
rect 13 453 27 467
rect 153 693 167 707
rect 233 813 247 827
rect 433 1172 447 1186
rect 613 1393 627 1407
rect 573 1353 587 1367
rect 553 1253 567 1267
rect 533 1214 547 1228
rect 673 1613 687 1627
rect 1133 2553 1147 2567
rect 1113 2533 1127 2547
rect 1153 2513 1167 2527
rect 1233 2533 1247 2547
rect 1113 2393 1127 2407
rect 1093 2373 1107 2387
rect 1133 2373 1147 2387
rect 1073 2333 1087 2347
rect 1073 2293 1087 2307
rect 1173 2333 1187 2347
rect 1133 2273 1147 2287
rect 1173 2273 1187 2287
rect 1373 2853 1387 2867
rect 1433 2833 1447 2847
rect 1393 2813 1407 2827
rect 1373 2773 1387 2787
rect 1273 2673 1287 2687
rect 1333 2673 1347 2687
rect 1273 2633 1287 2647
rect 1293 2474 1307 2488
rect 1313 2433 1327 2447
rect 1293 2393 1307 2407
rect 1273 2293 1287 2307
rect 1033 2254 1047 2268
rect 1133 2212 1147 2226
rect 1053 1993 1067 2007
rect 1093 1993 1107 2007
rect 1013 1973 1027 1987
rect 973 1954 987 1968
rect 1033 1953 1047 1967
rect 933 1933 947 1947
rect 893 1912 907 1926
rect 993 1893 1007 1907
rect 833 1873 847 1887
rect 833 1813 847 1827
rect 813 1753 827 1767
rect 753 1533 767 1547
rect 673 1473 687 1487
rect 693 1434 707 1448
rect 913 1733 927 1747
rect 853 1693 867 1707
rect 853 1673 867 1687
rect 873 1653 887 1667
rect 873 1553 887 1567
rect 813 1473 827 1487
rect 653 1393 667 1407
rect 713 1392 727 1406
rect 753 1392 767 1406
rect 793 1392 807 1406
rect 633 1353 647 1367
rect 733 1353 747 1367
rect 653 1273 667 1287
rect 633 1233 647 1247
rect 613 1213 627 1227
rect 553 1172 567 1186
rect 593 1172 607 1186
rect 393 953 407 967
rect 333 914 347 928
rect 433 914 447 928
rect 473 914 487 928
rect 333 873 347 887
rect 313 733 327 747
rect 253 694 267 708
rect 113 652 127 666
rect 233 652 247 666
rect 53 394 67 408
rect 93 394 107 408
rect 153 413 167 427
rect 233 413 247 427
rect 193 394 207 408
rect 273 394 287 408
rect 373 872 387 886
rect 413 872 427 886
rect 473 833 487 847
rect 433 733 447 747
rect 393 694 407 708
rect 473 693 487 707
rect 333 652 347 666
rect 373 652 387 666
rect 413 652 427 666
rect 433 453 447 467
rect 53 352 67 366
rect 113 333 127 347
rect 153 333 167 347
rect 13 174 27 188
rect 113 174 127 188
rect 353 393 367 407
rect 393 394 407 408
rect 593 1013 607 1027
rect 533 872 547 886
rect 513 753 527 767
rect 693 1233 707 1247
rect 653 1213 667 1227
rect 1133 1954 1147 1968
rect 1233 2254 1247 2268
rect 1493 2793 1507 2807
rect 1453 2774 1467 2788
rect 1533 2773 1547 2787
rect 1573 2913 1587 2927
rect 1633 2853 1647 2867
rect 1573 2713 1587 2727
rect 1473 2673 1487 2687
rect 1513 2673 1527 2687
rect 1613 2613 1627 2627
rect 1433 2573 1447 2587
rect 1493 2573 1507 2587
rect 1413 2553 1427 2567
rect 1373 2533 1387 2547
rect 1413 2493 1427 2507
rect 1353 2472 1367 2486
rect 1393 2474 1407 2488
rect 1433 2474 1447 2488
rect 1353 2433 1367 2447
rect 1313 2373 1327 2387
rect 1313 2293 1327 2307
rect 1213 2212 1227 2226
rect 1253 2212 1267 2226
rect 1193 2193 1207 2207
rect 1213 2173 1227 2187
rect 1193 2133 1207 2147
rect 1113 1912 1127 1926
rect 1153 1893 1167 1907
rect 1053 1813 1067 1827
rect 1033 1793 1047 1807
rect 1013 1773 1027 1787
rect 973 1653 987 1667
rect 1153 1773 1167 1787
rect 1113 1734 1127 1748
rect 1053 1692 1067 1706
rect 1093 1692 1107 1706
rect 1133 1673 1147 1687
rect 933 1613 947 1627
rect 973 1613 987 1627
rect 1033 1613 1047 1627
rect 913 1513 927 1527
rect 899 1453 913 1467
rect 853 1392 867 1406
rect 953 1393 967 1407
rect 913 1353 927 1367
rect 893 1273 907 1287
rect 773 1253 787 1267
rect 812 1253 826 1267
rect 833 1253 847 1267
rect 713 1172 727 1186
rect 673 1133 687 1147
rect 873 1213 887 1227
rect 1013 1434 1027 1448
rect 1073 1434 1087 1448
rect 1113 1434 1127 1448
rect 1153 1434 1167 1448
rect 1473 2433 1487 2447
rect 1413 2373 1427 2387
rect 1353 2333 1367 2347
rect 1393 2293 1407 2307
rect 1393 2254 1407 2268
rect 1593 2513 1607 2527
rect 1533 2474 1547 2488
rect 1693 3293 1707 3307
rect 1773 3433 1787 3447
rect 1753 3413 1767 3427
rect 1873 3452 1887 3466
rect 1793 3373 1807 3387
rect 1773 3353 1787 3367
rect 1753 3333 1767 3347
rect 1733 3313 1747 3327
rect 1813 3294 1827 3308
rect 1733 3252 1747 3266
rect 1793 3253 1807 3267
rect 1773 3213 1787 3227
rect 1753 3153 1767 3167
rect 1733 3113 1747 3127
rect 1713 3073 1727 3087
rect 1693 3053 1707 3067
rect 1713 3032 1727 3046
rect 1693 3013 1707 3027
rect 1893 3432 1907 3446
rect 1933 3433 1947 3447
rect 1973 3433 1987 3447
rect 1933 3373 1947 3387
rect 2033 3693 2047 3707
rect 2053 3613 2067 3627
rect 2033 3593 2047 3607
rect 2053 3573 2067 3587
rect 2253 3973 2267 3987
rect 2233 3913 2247 3927
rect 2212 3834 2226 3848
rect 2233 3833 2247 3847
rect 2173 3814 2187 3828
rect 2493 4293 2507 4307
rect 2533 4292 2547 4306
rect 2613 4313 2627 4327
rect 2513 4273 2527 4287
rect 2593 4273 2607 4287
rect 2493 4233 2507 4247
rect 2473 4093 2487 4107
rect 2453 4073 2467 4087
rect 2373 4034 2387 4048
rect 2493 4053 2507 4067
rect 2673 4334 2687 4348
rect 2733 4334 2747 4348
rect 2653 4273 2667 4287
rect 2533 4173 2547 4187
rect 2533 4073 2547 4087
rect 2553 4034 2567 4048
rect 2733 4233 2747 4247
rect 2653 4213 2667 4227
rect 2713 4213 2727 4227
rect 2613 4173 2627 4187
rect 2713 4133 2727 4147
rect 2673 4113 2687 4127
rect 2333 3973 2347 3987
rect 2313 3952 2327 3966
rect 2293 3933 2307 3947
rect 2213 3813 2227 3827
rect 2273 3813 2287 3827
rect 2153 3772 2167 3786
rect 2193 3772 2207 3786
rect 2233 3772 2247 3786
rect 2153 3733 2167 3747
rect 2133 3693 2147 3707
rect 2173 3713 2187 3727
rect 2132 3553 2146 3567
rect 2153 3553 2167 3567
rect 2113 3533 2127 3547
rect 2033 3513 2047 3527
rect 2073 3514 2087 3528
rect 2013 3353 2027 3367
rect 2013 3332 2027 3346
rect 1913 3293 1927 3307
rect 2013 3293 2027 3307
rect 1933 3252 1947 3266
rect 1993 3213 2007 3227
rect 2135 3473 2149 3487
rect 2093 3453 2107 3467
rect 2053 3433 2067 3447
rect 2093 3432 2107 3446
rect 2073 3393 2087 3407
rect 2533 3992 2547 4006
rect 2572 3993 2586 4007
rect 2593 3993 2607 4007
rect 2513 3973 2527 3987
rect 2393 3953 2407 3967
rect 2413 3933 2427 3947
rect 2333 3913 2347 3927
rect 2573 3933 2587 3947
rect 2493 3893 2507 3907
rect 2493 3872 2507 3886
rect 2392 3833 2406 3847
rect 2413 3833 2427 3847
rect 2353 3814 2367 3828
rect 2473 3813 2487 3827
rect 2293 3733 2307 3747
rect 2373 3772 2387 3786
rect 2353 3653 2367 3667
rect 2333 3633 2347 3647
rect 2213 3514 2227 3528
rect 2253 3514 2267 3528
rect 2413 3753 2427 3767
rect 2473 3673 2487 3687
rect 2413 3653 2427 3667
rect 2453 3653 2467 3667
rect 2373 3553 2387 3567
rect 2313 3533 2327 3547
rect 2353 3533 2367 3547
rect 2293 3513 2307 3527
rect 2193 3473 2207 3487
rect 2173 3433 2187 3447
rect 2153 3393 2167 3407
rect 2113 3373 2127 3387
rect 2053 3293 2067 3307
rect 2093 3293 2107 3307
rect 2293 3473 2307 3487
rect 2273 3413 2287 3427
rect 2233 3353 2247 3367
rect 2393 3514 2407 3528
rect 2433 3514 2447 3528
rect 2373 3472 2387 3486
rect 2413 3453 2427 3467
rect 2313 3413 2327 3427
rect 2433 3413 2447 3427
rect 2213 3333 2227 3347
rect 1893 3173 1907 3187
rect 2033 3173 2047 3187
rect 1993 3153 2007 3167
rect 1873 3133 1887 3147
rect 1973 3133 1987 3147
rect 1833 3113 1847 3127
rect 1713 2994 1727 3008
rect 1773 2994 1787 3008
rect 1713 2933 1727 2947
rect 1753 2933 1767 2947
rect 1693 2913 1707 2927
rect 1793 2913 1807 2927
rect 1773 2833 1787 2847
rect 1853 3073 1867 3087
rect 1953 3073 1967 3087
rect 1933 3053 1947 3067
rect 1913 3033 1927 3047
rect 1853 2994 1867 3008
rect 1893 2913 1907 2927
rect 1833 2873 1847 2887
rect 1813 2853 1827 2867
rect 1753 2813 1767 2827
rect 1793 2813 1807 2827
rect 1773 2793 1787 2807
rect 1753 2774 1767 2788
rect 1893 2794 1907 2808
rect 1893 2773 1907 2787
rect 2053 3073 2067 3087
rect 2033 3033 2047 3047
rect 2133 3252 2147 3266
rect 2113 3133 2127 3147
rect 2193 3213 2207 3227
rect 2173 3093 2187 3107
rect 2173 3072 2187 3086
rect 2113 2994 2127 3008
rect 2073 2973 2087 2987
rect 2013 2952 2027 2966
rect 1973 2913 1987 2927
rect 1953 2853 1967 2867
rect 1973 2813 1987 2827
rect 1952 2773 1966 2787
rect 1973 2774 1987 2788
rect 1693 2753 1707 2767
rect 1833 2753 1847 2767
rect 1633 2573 1647 2587
rect 1673 2573 1687 2587
rect 1713 2732 1727 2746
rect 1713 2693 1727 2707
rect 1713 2633 1727 2647
rect 1773 2732 1787 2746
rect 1753 2713 1767 2727
rect 1833 2673 1847 2687
rect 1753 2633 1767 2647
rect 1733 2613 1747 2627
rect 1753 2593 1767 2607
rect 1693 2553 1707 2567
rect 1653 2493 1667 2507
rect 1613 2473 1627 2487
rect 1713 2513 1727 2527
rect 1833 2573 1847 2587
rect 1733 2473 1747 2487
rect 1793 2474 1807 2488
rect 1513 2413 1527 2427
rect 1633 2413 1647 2427
rect 1493 2393 1507 2407
rect 1713 2413 1727 2427
rect 1673 2393 1687 2407
rect 1753 2433 1767 2447
rect 1733 2353 1747 2367
rect 1713 2333 1727 2347
rect 1573 2293 1587 2307
rect 1493 2253 1507 2267
rect 1533 2254 1547 2268
rect 1633 2254 1647 2268
rect 1693 2254 1707 2268
rect 1953 2733 1967 2747
rect 1952 2693 1966 2707
rect 1973 2693 1987 2707
rect 1913 2673 1927 2687
rect 1933 2653 1947 2667
rect 1913 2633 1927 2647
rect 1933 2613 1947 2627
rect 1893 2533 1907 2547
rect 1853 2513 1867 2527
rect 1773 2373 1787 2387
rect 1833 2373 1847 2387
rect 1753 2313 1767 2327
rect 1893 2474 1907 2488
rect 1973 2633 1987 2647
rect 1953 2513 1967 2527
rect 1873 2433 1887 2447
rect 1913 2413 1927 2427
rect 1873 2373 1887 2387
rect 1853 2333 1867 2347
rect 1773 2293 1787 2307
rect 1833 2293 1847 2307
rect 1312 2153 1326 2167
rect 1333 2153 1347 2167
rect 1273 2133 1287 2147
rect 1273 1953 1287 1967
rect 1373 2212 1387 2226
rect 1413 2212 1427 2226
rect 1473 2213 1487 2227
rect 1413 2133 1427 2147
rect 1413 2093 1427 2107
rect 1353 2073 1367 2087
rect 1373 2053 1387 2067
rect 1353 2033 1367 2047
rect 1213 1873 1227 1887
rect 1293 1873 1307 1887
rect 1333 1833 1347 1847
rect 1273 1813 1287 1827
rect 1213 1753 1227 1767
rect 1253 1753 1267 1767
rect 1333 1733 1347 1747
rect 1253 1673 1267 1687
rect 1213 1553 1227 1567
rect 1033 1392 1047 1406
rect 973 1333 987 1347
rect 1033 1333 1047 1347
rect 953 1214 967 1228
rect 1013 1213 1027 1227
rect 813 1172 827 1186
rect 933 1172 947 1186
rect 1133 1392 1147 1406
rect 1093 1313 1107 1327
rect 1173 1313 1187 1327
rect 1073 1253 1087 1267
rect 1293 1434 1307 1448
rect 1233 1413 1247 1427
rect 1313 1393 1327 1407
rect 1233 1353 1247 1367
rect 1273 1353 1287 1367
rect 1153 1273 1167 1287
rect 1213 1273 1227 1287
rect 1073 1214 1087 1228
rect 1133 1213 1147 1227
rect 873 1153 887 1167
rect 973 1153 987 1167
rect 773 1053 787 1067
rect 673 1013 687 1027
rect 913 973 927 987
rect 773 953 787 967
rect 713 914 727 928
rect 833 914 847 928
rect 733 872 747 886
rect 773 873 787 887
rect 1013 973 1027 987
rect 853 872 867 886
rect 913 872 927 886
rect 573 853 587 867
rect 633 853 647 867
rect 693 853 707 867
rect 773 833 787 847
rect 633 773 647 787
rect 733 773 747 787
rect 533 733 547 747
rect 573 694 587 708
rect 493 652 507 666
rect 553 652 567 666
rect 653 733 667 747
rect 753 733 767 747
rect 713 713 727 727
rect 993 853 1007 867
rect 1093 1172 1107 1186
rect 1093 1133 1107 1147
rect 1273 1253 1287 1267
rect 1193 1214 1207 1228
rect 1233 1214 1247 1228
rect 1293 1233 1307 1247
rect 1273 1213 1287 1227
rect 1253 1172 1267 1186
rect 1153 1033 1167 1047
rect 1413 1993 1427 2007
rect 1573 2193 1587 2207
rect 1493 2173 1507 2187
rect 1493 2113 1507 2127
rect 1473 2033 1487 2047
rect 1533 2073 1547 2087
rect 1513 2033 1527 2047
rect 1493 2013 1507 2027
rect 1373 1953 1387 1967
rect 1433 1973 1447 1987
rect 1473 1973 1487 1987
rect 1373 1913 1387 1927
rect 1413 1893 1427 1907
rect 1453 1893 1467 1907
rect 1433 1813 1447 1827
rect 1373 1734 1387 1748
rect 1393 1593 1407 1607
rect 1413 1553 1427 1567
rect 1433 1493 1447 1507
rect 1533 1993 1547 2007
rect 1553 1954 1567 1968
rect 1593 2173 1607 2187
rect 1533 1893 1547 1907
rect 1733 2253 1747 2267
rect 1793 2254 1807 2268
rect 1713 2213 1727 2227
rect 1733 2153 1747 2167
rect 1653 2133 1667 2147
rect 1713 2133 1727 2147
rect 1633 2113 1647 2127
rect 1613 2093 1627 2107
rect 1653 2093 1667 2107
rect 1933 2393 1947 2407
rect 1913 2373 1927 2387
rect 1893 2233 1907 2247
rect 1793 2173 1807 2187
rect 1813 2153 1827 2167
rect 1793 2133 1807 2147
rect 1773 2113 1787 2127
rect 1873 2193 1887 2207
rect 1893 2172 1907 2186
rect 1833 2093 1847 2107
rect 1753 2053 1767 2067
rect 1812 2053 1826 2067
rect 1833 2053 1847 2067
rect 1713 2033 1727 2047
rect 1753 2032 1767 2046
rect 1713 1973 1727 1987
rect 2053 2873 2067 2887
rect 2053 2833 2067 2847
rect 2073 2813 2087 2827
rect 2173 2933 2187 2947
rect 2053 2793 2067 2807
rect 2153 2793 2167 2807
rect 2033 2613 2047 2627
rect 2633 3833 2647 3847
rect 2713 3953 2727 3967
rect 2952 4693 2966 4707
rect 2973 4693 2987 4707
rect 2933 4553 2947 4567
rect 3013 4813 3027 4827
rect 3013 4753 3027 4767
rect 2993 4673 3007 4687
rect 3033 4633 3047 4647
rect 3033 4593 3047 4607
rect 3033 4554 3047 4568
rect 2833 4453 2847 4467
rect 2892 4513 2906 4527
rect 2913 4513 2927 4527
rect 2853 4433 2867 4447
rect 2813 4373 2827 4387
rect 2893 4393 2907 4407
rect 2953 4512 2967 4526
rect 3033 4473 3047 4487
rect 2993 4433 3007 4447
rect 3113 5113 3127 5127
rect 3093 5094 3107 5108
rect 3093 5074 3107 5088
rect 3113 5032 3127 5046
rect 3233 5213 3247 5227
rect 3353 5374 3367 5388
rect 3293 5332 3307 5346
rect 3333 5332 3347 5346
rect 3313 5313 3327 5327
rect 3693 5773 3707 5787
rect 3813 5894 3827 5908
rect 3793 5813 3807 5827
rect 3733 5793 3747 5807
rect 3713 5733 3727 5747
rect 3833 5713 3847 5727
rect 3773 5653 3787 5667
rect 3653 5573 3667 5587
rect 3593 5552 3607 5566
rect 3633 5553 3647 5567
rect 3553 5493 3567 5507
rect 3493 5433 3507 5447
rect 3513 5374 3527 5388
rect 3593 5374 3607 5388
rect 3633 5374 3647 5388
rect 3493 5332 3507 5346
rect 3393 5273 3407 5287
rect 3273 5233 3287 5247
rect 3253 5193 3267 5207
rect 3273 5113 3287 5127
rect 3313 5093 3327 5107
rect 3173 5074 3187 5088
rect 3233 5074 3247 5088
rect 3173 4993 3187 5007
rect 3153 4973 3167 4987
rect 3133 4953 3147 4967
rect 3093 4854 3107 4868
rect 3173 4853 3187 4867
rect 3093 4773 3107 4787
rect 3073 4673 3087 4687
rect 3153 4812 3167 4826
rect 3213 5032 3227 5046
rect 3153 4792 3167 4806
rect 3193 4753 3207 4767
rect 3173 4713 3187 4727
rect 3313 5032 3327 5046
rect 3253 4973 3267 4987
rect 3233 4854 3247 4868
rect 3273 4854 3287 4868
rect 3313 4812 3327 4826
rect 3273 4793 3287 4807
rect 3273 4733 3287 4747
rect 3253 4713 3267 4727
rect 3233 4693 3247 4707
rect 3213 4673 3227 4687
rect 3133 4633 3147 4647
rect 3193 4633 3207 4647
rect 3113 4593 3127 4607
rect 3153 4613 3167 4627
rect 3133 4573 3147 4587
rect 3113 4554 3127 4568
rect 3193 4573 3207 4587
rect 3233 4573 3247 4587
rect 3073 4513 3087 4527
rect 3053 4453 3067 4467
rect 3052 4432 3066 4446
rect 3073 4433 3087 4447
rect 3033 4413 3047 4427
rect 2993 4334 3007 4348
rect 3053 4333 3067 4347
rect 2833 4273 2847 4287
rect 2773 4173 2787 4187
rect 2933 4293 2947 4307
rect 3013 4292 3027 4306
rect 2872 4233 2886 4247
rect 2893 4233 2907 4247
rect 2973 4213 2987 4227
rect 2893 4193 2907 4207
rect 2873 4133 2887 4147
rect 2833 4113 2847 4127
rect 2813 4073 2827 4087
rect 2853 4034 2867 4048
rect 2733 3933 2747 3947
rect 2773 3913 2787 3927
rect 2693 3873 2707 3887
rect 2652 3813 2666 3827
rect 2673 3813 2687 3827
rect 2733 3814 2747 3828
rect 2653 3792 2667 3806
rect 2513 3693 2527 3707
rect 2493 3633 2507 3647
rect 2833 3992 2847 4006
rect 2953 4073 2967 4087
rect 3033 4253 3047 4267
rect 2993 4093 3007 4107
rect 2973 4053 2987 4067
rect 2833 3833 2847 3847
rect 2812 3813 2826 3827
rect 2873 3814 2887 3828
rect 2653 3753 2667 3767
rect 2613 3713 2627 3727
rect 2613 3653 2627 3667
rect 2593 3613 2607 3627
rect 2533 3514 2547 3528
rect 2713 3772 2727 3786
rect 2793 3773 2807 3787
rect 2673 3573 2687 3587
rect 2653 3533 2667 3547
rect 2693 3533 2707 3547
rect 2673 3473 2687 3487
rect 2593 3453 2607 3467
rect 2553 3413 2567 3427
rect 2513 3393 2527 3407
rect 2593 3373 2607 3387
rect 2833 3773 2847 3787
rect 2813 3693 2827 3707
rect 2953 3933 2967 3947
rect 2893 3753 2907 3767
rect 2933 3753 2947 3767
rect 2853 3693 2867 3707
rect 2833 3653 2847 3667
rect 2813 3553 2827 3567
rect 2813 3514 2827 3528
rect 2713 3473 2727 3487
rect 2773 3472 2787 3486
rect 2713 3433 2727 3447
rect 2693 3393 2707 3407
rect 2572 3353 2586 3367
rect 2293 3333 2307 3347
rect 2453 3333 2467 3347
rect 2273 3313 2287 3327
rect 2373 3313 2387 3327
rect 2353 3273 2367 3287
rect 2213 3073 2227 3087
rect 2313 3233 2327 3247
rect 2273 3173 2287 3187
rect 2193 2913 2207 2927
rect 2353 3213 2367 3227
rect 2333 3173 2347 3187
rect 2333 3133 2347 3147
rect 2273 2994 2287 3008
rect 2293 2952 2307 2966
rect 2433 3294 2447 3308
rect 2553 3253 2567 3267
rect 2533 3233 2547 3247
rect 2473 3193 2487 3207
rect 2413 3173 2427 3187
rect 2373 3113 2387 3127
rect 2432 3113 2446 3127
rect 2453 3113 2467 3127
rect 2413 3073 2427 3087
rect 2373 3053 2387 3067
rect 2293 2913 2307 2927
rect 2253 2893 2267 2907
rect 2273 2853 2287 2867
rect 2213 2813 2227 2827
rect 2172 2773 2186 2787
rect 2193 2773 2207 2787
rect 2093 2732 2107 2746
rect 2153 2713 2167 2727
rect 2073 2693 2087 2707
rect 1993 2573 2007 2587
rect 2053 2573 2067 2587
rect 2113 2613 2127 2627
rect 2093 2593 2107 2607
rect 2033 2553 2047 2567
rect 2073 2553 2087 2567
rect 2033 2493 2047 2507
rect 2093 2493 2107 2507
rect 2013 2474 2027 2488
rect 2133 2593 2147 2607
rect 2033 2333 2047 2347
rect 2193 2733 2207 2747
rect 2173 2593 2187 2607
rect 2193 2573 2207 2587
rect 2253 2553 2267 2567
rect 2213 2513 2227 2527
rect 2173 2493 2187 2507
rect 2153 2473 2167 2487
rect 2213 2474 2227 2488
rect 2313 2893 2327 2907
rect 2433 3053 2447 3067
rect 2533 3053 2547 3067
rect 2453 2994 2467 3008
rect 2493 2994 2507 3008
rect 2593 3352 2607 3366
rect 2673 3353 2687 3367
rect 2573 3233 2587 3247
rect 2573 3173 2587 3187
rect 2573 3073 2587 3087
rect 2553 3033 2567 3047
rect 2573 3013 2587 3027
rect 2693 3333 2707 3347
rect 2653 3294 2667 3308
rect 2653 3233 2667 3247
rect 2633 3153 2647 3167
rect 2613 3013 2627 3027
rect 2433 2952 2447 2966
rect 2393 2933 2407 2947
rect 2333 2833 2347 2847
rect 2593 2993 2607 3007
rect 2553 2952 2567 2966
rect 2533 2933 2547 2947
rect 2493 2873 2507 2887
rect 2433 2833 2447 2847
rect 2313 2773 2327 2787
rect 2413 2773 2427 2787
rect 2513 2753 2527 2767
rect 2313 2733 2327 2747
rect 2333 2713 2347 2727
rect 2313 2633 2327 2647
rect 2293 2593 2307 2607
rect 2293 2572 2307 2586
rect 2273 2513 2287 2527
rect 2273 2473 2287 2487
rect 2293 2473 2307 2487
rect 2413 2733 2427 2747
rect 2613 2913 2627 2927
rect 2593 2893 2607 2907
rect 2853 3633 2867 3647
rect 2893 3633 2907 3647
rect 2893 3593 2907 3607
rect 3033 4213 3047 4227
rect 3033 4133 3047 4147
rect 3133 4512 3147 4526
rect 3173 4453 3187 4467
rect 3093 4413 3107 4427
rect 3133 4413 3147 4427
rect 3293 4713 3307 4727
rect 3393 5252 3407 5266
rect 3393 5193 3407 5207
rect 3653 5332 3667 5346
rect 3513 5193 3527 5207
rect 3593 5193 3607 5207
rect 3673 5253 3687 5267
rect 3413 5153 3427 5167
rect 3493 5153 3507 5167
rect 3373 5093 3387 5107
rect 3433 5113 3447 5127
rect 3453 5094 3467 5108
rect 3453 5074 3467 5088
rect 3493 5053 3507 5067
rect 3393 5032 3407 5046
rect 3473 5033 3487 5047
rect 3433 5013 3447 5027
rect 3553 5093 3567 5107
rect 3573 5032 3587 5046
rect 3613 5033 3627 5047
rect 3513 5013 3527 5027
rect 3493 4973 3507 4987
rect 3473 4933 3487 4947
rect 3353 4913 3367 4927
rect 3413 4913 3427 4927
rect 3453 4913 3467 4927
rect 3453 4854 3467 4868
rect 3593 4893 3607 4907
rect 3553 4854 3567 4868
rect 3393 4812 3407 4826
rect 3472 4813 3486 4827
rect 3493 4813 3507 4827
rect 3433 4793 3447 4807
rect 3533 4812 3547 4826
rect 3333 4773 3347 4787
rect 3473 4733 3487 4747
rect 3453 4693 3467 4707
rect 3353 4633 3367 4647
rect 3313 4593 3327 4607
rect 3193 4433 3207 4447
rect 3313 4513 3327 4527
rect 3373 4512 3387 4526
rect 3273 4473 3287 4487
rect 3353 4473 3367 4487
rect 3413 4473 3427 4487
rect 3293 4433 3307 4447
rect 3273 4393 3287 4407
rect 3213 4373 3227 4387
rect 3253 4373 3267 4387
rect 3153 4233 3167 4247
rect 3153 4113 3167 4127
rect 3073 4073 3087 4087
rect 3113 4053 3127 4067
rect 3033 4034 3047 4048
rect 3093 4034 3107 4048
rect 3053 3992 3067 4006
rect 3013 3933 3027 3947
rect 2973 3813 2987 3827
rect 3013 3814 3027 3828
rect 3073 3813 3087 3827
rect 3173 4093 3187 4107
rect 3233 4353 3247 4367
rect 3233 4273 3247 4287
rect 3313 4292 3327 4306
rect 3513 4793 3527 4807
rect 3573 4773 3587 4787
rect 3513 4693 3527 4707
rect 3553 4673 3567 4687
rect 3533 4653 3547 4667
rect 3553 4553 3567 4567
rect 3453 4513 3467 4527
rect 3433 4453 3447 4467
rect 3413 4433 3427 4447
rect 3453 4393 3467 4407
rect 3433 4353 3447 4367
rect 3413 4334 3427 4348
rect 3513 4512 3527 4526
rect 3533 4493 3547 4507
rect 3493 4473 3507 4487
rect 3473 4353 3487 4367
rect 3453 4333 3467 4347
rect 3432 4292 3446 4306
rect 3453 4292 3467 4306
rect 3393 4213 3407 4227
rect 3293 4153 3307 4167
rect 3353 4153 3367 4167
rect 3393 4153 3407 4167
rect 3213 4053 3227 4067
rect 3173 4033 3187 4047
rect 3273 4073 3287 4087
rect 3153 3993 3167 4007
rect 3193 3992 3207 4006
rect 3153 3953 3167 3967
rect 3193 3953 3207 3967
rect 3173 3913 3187 3927
rect 3153 3853 3167 3867
rect 3133 3833 3147 3847
rect 3253 3873 3267 3887
rect 3233 3853 3247 3867
rect 3053 3772 3067 3786
rect 2993 3753 3007 3767
rect 2853 3553 2867 3567
rect 2953 3553 2967 3567
rect 2893 3514 2907 3528
rect 2933 3514 2947 3528
rect 3173 3772 3187 3786
rect 3213 3773 3227 3787
rect 3093 3733 3107 3747
rect 3113 3613 3127 3627
rect 3113 3553 3127 3567
rect 3053 3514 3067 3528
rect 3213 3533 3227 3547
rect 3173 3514 3187 3528
rect 3213 3512 3227 3526
rect 2873 3472 2887 3486
rect 2913 3472 2927 3486
rect 2973 3473 2987 3487
rect 2853 3413 2867 3427
rect 2753 3333 2767 3347
rect 2833 3333 2847 3347
rect 2733 3313 2747 3327
rect 2713 3233 2727 3247
rect 2793 3313 2807 3327
rect 2753 3294 2767 3308
rect 2773 3193 2787 3207
rect 2733 3093 2747 3107
rect 2773 3013 2787 3027
rect 2673 2994 2687 3008
rect 2713 2994 2727 3008
rect 2633 2853 2647 2867
rect 2673 2813 2687 2827
rect 2513 2713 2527 2727
rect 2453 2673 2467 2687
rect 2433 2653 2447 2667
rect 2413 2613 2427 2627
rect 2393 2593 2407 2607
rect 2393 2553 2407 2567
rect 2373 2513 2387 2527
rect 1972 2293 1986 2307
rect 1993 2293 2007 2307
rect 2053 2293 2067 2307
rect 2133 2293 2147 2307
rect 1933 2273 1947 2287
rect 1973 2272 1987 2286
rect 1933 2193 1947 2207
rect 1973 2153 1987 2167
rect 1912 2113 1926 2127
rect 1933 2113 1947 2127
rect 1913 2092 1927 2106
rect 1893 2033 1907 2047
rect 1833 2013 1847 2027
rect 1893 1973 1907 1987
rect 2013 2254 2027 2268
rect 2013 2173 2027 2187
rect 1993 2093 2007 2107
rect 2113 2254 2127 2268
rect 2073 2212 2087 2226
rect 2053 2133 2067 2147
rect 2113 2193 2127 2207
rect 2033 2073 2047 2087
rect 1933 2053 1947 2067
rect 1973 2053 1987 2067
rect 1933 2032 1947 2046
rect 2013 2013 2027 2027
rect 1933 1993 1947 2007
rect 1953 1974 1967 1988
rect 1593 1912 1607 1926
rect 1633 1912 1647 1926
rect 1573 1893 1587 1907
rect 1593 1833 1607 1847
rect 1473 1813 1487 1827
rect 1573 1753 1587 1767
rect 1513 1734 1527 1748
rect 1473 1533 1487 1547
rect 1413 1313 1427 1327
rect 1332 1233 1346 1247
rect 1353 1233 1367 1247
rect 1453 1233 1467 1247
rect 1313 1172 1327 1186
rect 1373 1172 1387 1186
rect 1413 1172 1427 1186
rect 1293 1073 1307 1087
rect 1313 1033 1327 1047
rect 1273 1013 1287 1027
rect 1153 973 1167 987
rect 1073 933 1087 947
rect 1133 933 1147 947
rect 1493 1493 1507 1507
rect 1573 1533 1587 1547
rect 1573 1512 1587 1526
rect 1753 1954 1767 1968
rect 1793 1954 1807 1968
rect 1913 1953 1927 1967
rect 1953 1953 1967 1967
rect 2093 2113 2107 2127
rect 2053 2033 2067 2047
rect 2113 2053 2127 2067
rect 2033 1973 2047 1987
rect 1753 1913 1767 1927
rect 1633 1753 1647 1767
rect 1673 1734 1687 1748
rect 1653 1692 1667 1706
rect 1693 1692 1707 1706
rect 1733 1692 1747 1706
rect 1533 1473 1547 1487
rect 1533 1434 1547 1448
rect 1673 1633 1687 1647
rect 1613 1453 1627 1467
rect 1653 1453 1667 1467
rect 1493 1293 1507 1307
rect 1553 1392 1567 1406
rect 1733 1593 1747 1607
rect 1713 1513 1727 1527
rect 1673 1434 1687 1448
rect 1813 1913 1827 1927
rect 1813 1793 1827 1807
rect 1893 1913 1907 1927
rect 1893 1833 1907 1847
rect 1933 1913 1947 1927
rect 1913 1813 1927 1827
rect 1893 1793 1907 1807
rect 1773 1773 1787 1787
rect 1833 1773 1847 1787
rect 1793 1734 1807 1748
rect 1833 1734 1847 1748
rect 1773 1693 1787 1707
rect 1753 1573 1767 1587
rect 1753 1552 1767 1566
rect 1813 1673 1827 1687
rect 1833 1573 1847 1587
rect 1733 1433 1747 1447
rect 1873 1693 1887 1707
rect 1853 1434 1867 1448
rect 1953 1893 1967 1907
rect 1912 1773 1926 1787
rect 1933 1773 1947 1787
rect 1893 1673 1907 1687
rect 1893 1613 1907 1627
rect 1893 1553 1907 1567
rect 2193 2432 2207 2446
rect 2193 2333 2207 2347
rect 2173 2293 2187 2307
rect 2153 2153 2167 2167
rect 2153 2073 2167 2087
rect 2153 2033 2167 2047
rect 2233 2293 2247 2307
rect 2193 2273 2207 2287
rect 2333 2432 2347 2446
rect 2393 2493 2407 2507
rect 2293 2353 2307 2367
rect 2352 2353 2366 2367
rect 2373 2353 2387 2367
rect 2213 2212 2227 2226
rect 2253 2212 2267 2226
rect 2293 2213 2307 2227
rect 2293 2192 2307 2206
rect 2213 2173 2227 2187
rect 2173 2013 2187 2027
rect 2073 1973 2087 1987
rect 2133 1974 2147 1988
rect 2133 1953 2147 1967
rect 2173 1954 2187 1968
rect 2093 1913 2107 1927
rect 2073 1853 2087 1867
rect 2093 1833 2107 1847
rect 2133 1853 2147 1867
rect 2113 1793 2127 1807
rect 2153 1813 2167 1827
rect 2013 1773 2027 1787
rect 2053 1773 2067 1787
rect 2133 1773 2147 1787
rect 1973 1734 1987 1748
rect 2073 1733 2087 1747
rect 2133 1734 2147 1748
rect 1953 1613 1967 1627
rect 1933 1593 1947 1607
rect 1953 1573 1967 1587
rect 1933 1493 1947 1507
rect 2073 1673 2087 1687
rect 2033 1653 2047 1667
rect 2073 1613 2087 1627
rect 2013 1533 2027 1547
rect 1993 1493 2007 1507
rect 2133 1673 2147 1687
rect 2133 1652 2147 1666
rect 2193 1653 2207 1667
rect 2113 1613 2127 1627
rect 2133 1593 2147 1607
rect 2233 2153 2247 2167
rect 2293 2153 2307 2167
rect 2333 2212 2347 2226
rect 2353 2173 2367 2187
rect 2353 2073 2367 2087
rect 2313 1993 2327 2007
rect 2333 1933 2347 1947
rect 2313 1853 2327 1867
rect 2253 1773 2267 1787
rect 2333 1793 2347 1807
rect 2493 2593 2507 2607
rect 2453 2533 2467 2547
rect 2533 2473 2547 2487
rect 2453 2432 2467 2446
rect 2513 2433 2527 2447
rect 2473 2353 2487 2367
rect 2453 2273 2467 2287
rect 2433 2254 2447 2268
rect 2513 2293 2527 2307
rect 2573 2713 2587 2727
rect 2713 2933 2727 2947
rect 2693 2753 2707 2767
rect 2753 2933 2767 2947
rect 2733 2913 2747 2927
rect 2792 2994 2806 3008
rect 2833 3193 2847 3207
rect 2773 2873 2787 2887
rect 2773 2813 2787 2827
rect 2753 2793 2767 2807
rect 2813 2993 2827 3007
rect 3033 3453 3047 3467
rect 2993 3433 3007 3447
rect 2973 3393 2987 3407
rect 2913 3373 2927 3387
rect 2973 3253 2987 3267
rect 3093 3473 3107 3487
rect 3073 3413 3087 3427
rect 3013 3333 3027 3347
rect 3073 3294 3087 3308
rect 3033 3252 3047 3266
rect 3013 3213 3027 3227
rect 3073 3213 3087 3227
rect 2993 3173 3007 3187
rect 2873 3113 2887 3127
rect 2933 3113 2947 3127
rect 3013 3093 3027 3107
rect 2933 3073 2947 3087
rect 3013 3013 3027 3027
rect 2873 2994 2887 3008
rect 2933 2994 2947 3008
rect 2853 2933 2867 2947
rect 2933 2953 2947 2967
rect 2993 2952 3007 2966
rect 2893 2933 2907 2947
rect 2813 2873 2827 2887
rect 2913 2873 2927 2887
rect 2793 2793 2807 2807
rect 2853 2793 2867 2807
rect 2732 2733 2746 2747
rect 2673 2713 2687 2727
rect 2713 2673 2727 2687
rect 2633 2653 2647 2667
rect 2593 2633 2607 2647
rect 2713 2633 2727 2647
rect 2753 2732 2767 2746
rect 2833 2733 2847 2747
rect 2613 2613 2627 2627
rect 2653 2613 2667 2627
rect 2733 2613 2747 2627
rect 2633 2593 2647 2607
rect 2593 2432 2607 2446
rect 2553 2333 2567 2347
rect 2553 2293 2567 2307
rect 2533 2253 2547 2267
rect 2413 2213 2427 2227
rect 2413 2113 2427 2127
rect 2433 2093 2447 2107
rect 2433 2033 2447 2047
rect 2393 1954 2407 1968
rect 2493 2212 2507 2226
rect 2533 2212 2547 2226
rect 2453 1973 2467 1987
rect 2273 1753 2287 1767
rect 2313 1753 2327 1767
rect 2413 1912 2427 1926
rect 2473 1893 2487 1907
rect 2413 1853 2427 1867
rect 2293 1673 2307 1687
rect 2253 1653 2267 1667
rect 2213 1553 2227 1567
rect 2293 1593 2307 1607
rect 2253 1533 2267 1547
rect 2053 1493 2067 1507
rect 2013 1473 2027 1487
rect 1693 1392 1707 1406
rect 1753 1392 1767 1406
rect 1653 1353 1667 1367
rect 1733 1293 1747 1307
rect 1533 1253 1547 1267
rect 1613 1253 1627 1267
rect 1493 1213 1507 1227
rect 1693 1233 1707 1247
rect 1553 1214 1567 1228
rect 1533 1172 1547 1186
rect 1593 1173 1607 1187
rect 1573 1153 1587 1167
rect 1493 1113 1507 1127
rect 1473 1013 1487 1027
rect 1333 993 1347 1007
rect 1453 993 1467 1007
rect 1073 872 1087 886
rect 1133 872 1147 886
rect 953 813 967 827
rect 933 773 947 787
rect 813 733 827 747
rect 893 733 907 747
rect 772 693 786 707
rect 793 693 807 707
rect 733 652 747 666
rect 733 573 747 587
rect 673 453 687 467
rect 473 394 487 408
rect 513 394 527 408
rect 573 394 587 408
rect 253 352 267 366
rect 193 333 207 347
rect 293 293 307 307
rect 173 233 187 247
rect 293 213 307 227
rect 213 174 227 188
rect 93 132 107 146
rect 153 133 167 147
rect 333 352 347 366
rect 333 233 347 247
rect 413 352 427 366
rect 453 352 467 366
rect 513 353 527 367
rect 553 293 567 307
rect 693 433 707 447
rect 793 433 807 447
rect 853 694 867 708
rect 1053 733 1067 747
rect 953 713 967 727
rect 1013 694 1027 708
rect 913 652 927 666
rect 953 652 967 666
rect 873 533 887 547
rect 1033 652 1047 666
rect 993 613 1007 627
rect 933 533 947 547
rect 693 393 707 407
rect 733 394 747 408
rect 733 333 747 347
rect 673 313 687 327
rect 593 253 607 267
rect 593 232 607 246
rect 353 213 367 227
rect 313 174 327 188
rect 393 193 407 207
rect 433 173 447 187
rect 513 174 527 188
rect 553 174 567 188
rect 233 132 247 146
rect 293 132 307 146
rect 373 113 387 127
rect 433 113 447 127
rect 13 93 27 107
rect 193 93 207 107
rect 533 93 547 107
rect 673 174 687 188
rect 653 132 667 146
rect 793 353 807 367
rect 753 313 767 327
rect 1313 914 1327 928
rect 1413 914 1427 928
rect 1273 872 1287 886
rect 1333 872 1347 886
rect 1233 833 1247 847
rect 1173 793 1187 807
rect 1153 733 1167 747
rect 1113 693 1127 707
rect 1193 694 1207 708
rect 1393 813 1407 827
rect 1313 753 1327 767
rect 1413 793 1427 807
rect 1313 713 1327 727
rect 1393 713 1407 727
rect 1233 693 1247 707
rect 1093 513 1107 527
rect 1173 652 1187 666
rect 1213 652 1227 666
rect 1193 573 1207 587
rect 973 473 987 487
rect 1113 473 1127 487
rect 1153 473 1167 487
rect 833 333 847 347
rect 913 333 927 347
rect 873 293 887 307
rect 793 273 807 287
rect 833 273 847 287
rect 793 174 807 188
rect 853 253 867 267
rect 853 193 867 207
rect 773 132 787 146
rect 1073 433 1087 447
rect 1073 394 1087 408
rect 1013 313 1027 327
rect 1333 694 1347 708
rect 1373 694 1387 708
rect 1313 652 1327 666
rect 1353 652 1367 666
rect 1393 652 1407 666
rect 1513 1073 1527 1087
rect 1553 1073 1567 1087
rect 1653 1153 1667 1167
rect 1593 973 1607 987
rect 1593 914 1607 928
rect 1833 1392 1847 1406
rect 1813 1273 1827 1287
rect 1793 1233 1807 1247
rect 1953 1434 1967 1448
rect 1973 1392 1987 1406
rect 2013 1392 2027 1406
rect 1953 1253 1967 1267
rect 1853 1233 1867 1247
rect 1893 1233 1907 1247
rect 1833 1172 1847 1186
rect 1913 1214 1927 1228
rect 1993 1213 2007 1227
rect 1893 1172 1907 1186
rect 1973 1173 1987 1187
rect 1773 1073 1787 1087
rect 1853 1073 1867 1087
rect 1733 1033 1747 1047
rect 1873 1013 1887 1027
rect 1673 914 1687 928
rect 1713 914 1727 928
rect 1913 914 1927 928
rect 2093 1453 2107 1467
rect 2193 1453 2207 1467
rect 2133 1434 2147 1448
rect 2113 1392 2127 1406
rect 2173 1373 2187 1387
rect 2073 1333 2087 1347
rect 2073 1253 2087 1267
rect 2113 1253 2127 1267
rect 2073 1214 2087 1228
rect 2253 1434 2267 1448
rect 2233 1333 2247 1347
rect 2273 1333 2287 1347
rect 2233 1293 2247 1307
rect 2153 1213 2167 1227
rect 2193 1214 2207 1228
rect 2253 1233 2267 1247
rect 2233 1213 2247 1227
rect 2013 1153 2027 1167
rect 1993 1013 2007 1027
rect 1573 872 1587 886
rect 1573 793 1587 807
rect 1513 733 1527 747
rect 1553 733 1567 747
rect 1513 652 1527 666
rect 1373 613 1387 627
rect 1433 553 1447 567
rect 1553 553 1567 567
rect 1273 513 1287 527
rect 1253 433 1267 447
rect 1233 413 1247 427
rect 1173 352 1187 366
rect 973 293 987 307
rect 1053 293 1067 307
rect 1113 293 1127 307
rect 1213 253 1227 267
rect 893 233 907 247
rect 932 233 946 247
rect 953 233 967 247
rect 1133 213 1147 227
rect 953 193 967 207
rect 973 174 987 188
rect 1013 174 1027 188
rect 1093 174 1107 188
rect 1033 153 1047 167
rect 913 132 927 146
rect 1013 133 1027 147
rect 733 93 747 107
rect 813 93 827 107
rect 493 73 507 87
rect 593 73 607 87
rect 1053 73 1067 87
rect 1153 173 1167 187
rect 1393 493 1407 507
rect 1293 413 1307 427
rect 1353 394 1367 408
rect 1293 352 1307 366
rect 1373 352 1387 366
rect 1293 313 1307 327
rect 1273 213 1287 227
rect 1253 173 1267 187
rect 1393 193 1407 207
rect 1313 174 1327 188
rect 1353 174 1367 188
rect 1153 132 1167 146
rect 1133 93 1147 107
rect 1233 132 1247 146
rect 1293 132 1307 146
rect 1333 132 1347 146
rect 1353 113 1367 127
rect 1193 73 1207 87
rect 1373 73 1387 87
rect 1113 53 1127 67
rect 1353 53 1367 67
rect 1553 493 1567 507
rect 1453 393 1467 407
rect 1653 872 1667 886
rect 1773 872 1787 886
rect 1853 872 1867 886
rect 1733 853 1747 867
rect 1893 793 1907 807
rect 1613 733 1627 747
rect 1913 733 1927 747
rect 1773 713 1787 727
rect 1833 713 1847 727
rect 1733 694 1747 708
rect 1673 673 1687 687
rect 1613 633 1627 647
rect 1573 473 1587 487
rect 1633 413 1647 427
rect 1573 394 1587 408
rect 1753 633 1767 647
rect 1733 533 1747 547
rect 1693 413 1707 427
rect 1453 352 1467 366
rect 1533 352 1547 366
rect 1513 313 1527 327
rect 1493 293 1507 307
rect 1693 352 1707 366
rect 1873 694 1887 708
rect 2013 914 2027 928
rect 2053 1153 2067 1167
rect 2213 1172 2227 1186
rect 2153 1153 2167 1167
rect 2153 1073 2167 1087
rect 2073 1013 2087 1027
rect 1953 693 1967 707
rect 1933 652 1947 666
rect 1993 872 2007 886
rect 2113 953 2127 967
rect 2213 1033 2227 1047
rect 2153 914 2167 928
rect 2193 913 2207 927
rect 2073 872 2087 886
rect 2053 773 2067 787
rect 2153 773 2167 787
rect 2053 733 2067 747
rect 2133 733 2147 747
rect 2013 694 2027 708
rect 2193 753 2207 767
rect 2313 1493 2327 1507
rect 2373 1733 2387 1747
rect 2553 1973 2567 1987
rect 2633 2419 2647 2433
rect 2613 2333 2627 2347
rect 2633 2313 2647 2327
rect 2673 2573 2687 2587
rect 2653 2213 2667 2227
rect 2633 2173 2647 2187
rect 2833 2613 2847 2627
rect 2793 2573 2807 2587
rect 2953 2774 2967 2788
rect 2993 2773 3007 2787
rect 2933 2732 2947 2746
rect 2893 2713 2907 2727
rect 2913 2693 2927 2707
rect 2893 2673 2907 2687
rect 2893 2633 2907 2647
rect 2953 2553 2967 2567
rect 2853 2513 2867 2527
rect 2753 2493 2767 2507
rect 2833 2493 2847 2507
rect 2713 2474 2727 2488
rect 2773 2432 2787 2446
rect 2733 2393 2747 2407
rect 2693 2373 2707 2387
rect 2893 2474 2907 2488
rect 3033 2933 3047 2947
rect 3193 3472 3207 3486
rect 3213 3453 3227 3467
rect 3193 3413 3207 3427
rect 3113 3373 3127 3387
rect 3313 4133 3327 4147
rect 3293 4033 3307 4047
rect 3353 4093 3367 4107
rect 3573 4333 3587 4347
rect 3553 4292 3567 4306
rect 3513 4253 3527 4267
rect 3473 4173 3487 4187
rect 3473 4113 3487 4127
rect 3453 4093 3467 4107
rect 3433 4073 3447 4087
rect 3393 4053 3407 4067
rect 3453 4053 3467 4067
rect 3333 3992 3347 4006
rect 3493 4034 3507 4048
rect 3553 4133 3567 4147
rect 3533 4113 3547 4127
rect 3333 3971 3347 3985
rect 3393 3973 3407 3987
rect 3273 3833 3287 3847
rect 3353 3913 3367 3927
rect 3473 3992 3487 4006
rect 3433 3973 3447 3987
rect 3493 3973 3507 3987
rect 3413 3893 3427 3907
rect 3653 5173 3667 5187
rect 3633 4973 3647 4987
rect 3653 4953 3667 4967
rect 3652 4913 3666 4927
rect 3673 4913 3687 4927
rect 3873 5793 3887 5807
rect 4013 6114 4027 6128
rect 3913 5953 3927 5967
rect 4133 6153 4147 6167
rect 4193 6153 4207 6167
rect 4273 6153 4287 6167
rect 4053 6113 4067 6127
rect 4093 6114 4107 6128
rect 4033 6033 4047 6047
rect 3993 5953 4007 5967
rect 3973 5913 3987 5927
rect 3913 5893 3927 5907
rect 3933 5852 3947 5866
rect 3913 5833 3927 5847
rect 3893 5693 3907 5707
rect 3873 5594 3887 5608
rect 3773 5473 3787 5487
rect 3873 5493 3887 5507
rect 3813 5433 3827 5447
rect 3813 5412 3827 5426
rect 3773 5374 3787 5388
rect 3853 5374 3867 5388
rect 3953 5813 3967 5827
rect 4013 5852 4027 5866
rect 4213 6114 4227 6128
rect 4193 6093 4207 6107
rect 4153 6072 4167 6086
rect 4133 5894 4147 5908
rect 4413 6133 4427 6147
rect 4373 6114 4387 6128
rect 4333 6093 4347 6107
rect 4313 6073 4327 6087
rect 4212 6033 4226 6047
rect 4233 6033 4247 6047
rect 4233 5993 4247 6007
rect 4193 5953 4207 5967
rect 4173 5893 4187 5907
rect 3993 5813 4007 5827
rect 3972 5753 3986 5767
rect 3993 5753 4007 5767
rect 4053 5852 4067 5866
rect 4113 5852 4127 5866
rect 4033 5833 4047 5847
rect 4013 5733 4027 5747
rect 4173 5853 4187 5867
rect 4153 5713 4167 5727
rect 4213 5913 4227 5927
rect 4193 5713 4207 5727
rect 3933 5653 3947 5667
rect 4013 5653 4027 5667
rect 4173 5653 4187 5667
rect 3913 5633 3927 5647
rect 3973 5613 3987 5627
rect 3933 5594 3947 5608
rect 4273 5973 4287 5987
rect 4253 5953 4267 5967
rect 4233 5893 4247 5907
rect 4313 5933 4327 5947
rect 4373 5973 4387 5987
rect 4433 6072 4447 6086
rect 4453 5933 4467 5947
rect 4392 5913 4406 5927
rect 4427 5913 4441 5927
rect 4333 5893 4347 5907
rect 4253 5852 4267 5866
rect 4293 5852 4307 5866
rect 4253 5793 4267 5807
rect 4213 5613 4227 5627
rect 4073 5594 4087 5608
rect 4153 5573 4167 5587
rect 3953 5552 3967 5566
rect 4013 5553 4027 5567
rect 4073 5533 4087 5547
rect 3993 5433 4007 5447
rect 3933 5374 3947 5388
rect 3793 5332 3807 5346
rect 3713 5153 3727 5167
rect 3853 5153 3867 5167
rect 3933 5153 3947 5167
rect 3793 5113 3807 5127
rect 3893 5113 3907 5127
rect 3773 5074 3787 5088
rect 3873 5074 3887 5088
rect 3793 5033 3807 5047
rect 3873 5033 3887 5047
rect 3713 4993 3727 5007
rect 3693 4893 3707 4907
rect 3653 4874 3667 4888
rect 3613 4853 3627 4867
rect 3653 4853 3667 4867
rect 3753 4953 3767 4967
rect 3733 4913 3747 4927
rect 3633 4812 3647 4826
rect 3673 4812 3687 4826
rect 3733 4812 3747 4826
rect 3653 4733 3667 4747
rect 3633 4673 3647 4687
rect 3653 4633 3667 4647
rect 3633 4593 3647 4607
rect 3733 4693 3747 4707
rect 3813 5013 3827 5027
rect 3873 4993 3887 5007
rect 3953 5032 3967 5046
rect 3893 4953 3907 4967
rect 3833 4933 3847 4947
rect 3793 4873 3807 4887
rect 3773 4853 3787 4867
rect 3873 4854 3887 4868
rect 4013 5413 4027 5427
rect 4173 5533 4187 5547
rect 4153 5513 4167 5527
rect 4093 5493 4107 5507
rect 4133 5374 4147 5388
rect 4333 5753 4347 5767
rect 4453 5894 4467 5908
rect 4373 5853 4387 5867
rect 4353 5693 4367 5707
rect 4393 5793 4407 5807
rect 4473 5853 4487 5867
rect 4673 6173 4687 6187
rect 4713 6173 4727 6187
rect 4693 6153 4707 6167
rect 4733 6153 4747 6167
rect 4873 6153 4887 6167
rect 4533 6133 4547 6147
rect 4553 6113 4567 6127
rect 4593 6114 4607 6128
rect 4533 6072 4547 6086
rect 4553 6053 4567 6067
rect 4533 6033 4547 6047
rect 4613 6073 4627 6087
rect 4693 6114 4707 6128
rect 4833 6114 4847 6128
rect 5193 6173 5207 6187
rect 5473 6173 5487 6187
rect 5613 6173 5627 6187
rect 4713 6072 4727 6086
rect 4853 6072 4867 6086
rect 4633 6053 4647 6067
rect 4673 6053 4687 6067
rect 4733 6033 4747 6047
rect 4613 6013 4627 6027
rect 4573 5993 4587 6007
rect 4613 5973 4627 5987
rect 4553 5953 4567 5967
rect 4533 5933 4547 5947
rect 4573 5913 4587 5927
rect 4513 5893 4527 5907
rect 4653 5933 4667 5947
rect 4613 5894 4627 5908
rect 4493 5833 4507 5847
rect 4473 5813 4487 5827
rect 4433 5773 4447 5787
rect 4493 5773 4507 5787
rect 4393 5733 4407 5747
rect 4813 5973 4827 5987
rect 4793 5893 4807 5907
rect 4593 5833 4607 5847
rect 4653 5852 4667 5866
rect 4713 5852 4727 5866
rect 4753 5852 4767 5866
rect 4633 5813 4647 5827
rect 4553 5733 4567 5747
rect 4513 5713 4527 5727
rect 4653 5653 4667 5667
rect 4373 5633 4387 5647
rect 4473 5633 4487 5647
rect 4533 5633 4547 5647
rect 4353 5613 4367 5627
rect 4293 5594 4307 5608
rect 4353 5592 4367 5606
rect 4393 5594 4407 5608
rect 4433 5594 4447 5608
rect 4253 5493 4267 5507
rect 4353 5533 4367 5547
rect 4413 5513 4427 5527
rect 4313 5453 4327 5467
rect 4233 5413 4247 5427
rect 4027 5312 4041 5326
rect 4053 5313 4067 5327
rect 4133 5292 4147 5306
rect 4113 5113 4127 5127
rect 4093 5093 4107 5107
rect 4073 5074 4087 5088
rect 4493 5594 4507 5608
rect 4533 5594 4547 5608
rect 4573 5594 4587 5608
rect 4513 5553 4527 5567
rect 4493 5513 4507 5527
rect 4413 5413 4427 5427
rect 4473 5413 4487 5427
rect 4333 5374 4347 5388
rect 4373 5374 4387 5388
rect 4313 5332 4327 5346
rect 4393 5332 4407 5346
rect 4433 5332 4447 5346
rect 4473 5332 4487 5346
rect 4293 5273 4307 5287
rect 4333 5273 4347 5287
rect 4053 5013 4067 5027
rect 4093 5013 4107 5027
rect 4133 5013 4147 5027
rect 4013 4973 4027 4987
rect 4113 4973 4127 4987
rect 4033 4953 4047 4967
rect 3993 4893 4007 4907
rect 3913 4853 3927 4867
rect 3953 4854 3967 4868
rect 3993 4854 4007 4868
rect 4053 4893 4067 4907
rect 3853 4812 3867 4826
rect 3813 4753 3827 4767
rect 3693 4613 3707 4627
rect 3673 4553 3687 4567
rect 3653 4512 3667 4526
rect 3613 4493 3627 4507
rect 3653 4453 3667 4467
rect 3773 4673 3787 4687
rect 3753 4653 3767 4667
rect 3753 4613 3767 4627
rect 3733 4593 3747 4607
rect 3773 4573 3787 4587
rect 3753 4554 3767 4568
rect 3913 4753 3927 4767
rect 3853 4733 3867 4747
rect 3833 4693 3847 4707
rect 3773 4473 3787 4487
rect 3693 4453 3707 4467
rect 3673 4433 3687 4447
rect 3773 4433 3787 4447
rect 3713 4393 3727 4407
rect 3753 4353 3767 4367
rect 3633 4333 3647 4347
rect 3673 4334 3687 4348
rect 3733 4334 3747 4348
rect 3593 4053 3607 4067
rect 3553 4033 3567 4047
rect 3613 4033 3627 4047
rect 3713 4292 3727 4306
rect 3653 4253 3667 4267
rect 3693 4213 3707 4227
rect 3693 4173 3707 4187
rect 3673 4093 3687 4107
rect 3533 3953 3547 3967
rect 3593 3992 3607 4006
rect 3493 3893 3507 3907
rect 3553 3893 3567 3907
rect 3613 3893 3627 3907
rect 3473 3873 3487 3887
rect 3353 3833 3367 3847
rect 3433 3833 3447 3847
rect 3293 3814 3307 3828
rect 3333 3814 3347 3828
rect 3273 3772 3287 3786
rect 3353 3773 3367 3787
rect 3333 3753 3347 3767
rect 3313 3733 3327 3747
rect 3313 3613 3327 3627
rect 3333 3573 3347 3587
rect 3293 3433 3307 3447
rect 3133 3333 3147 3347
rect 3233 3333 3247 3347
rect 3113 3294 3127 3308
rect 3093 3093 3107 3107
rect 3093 2993 3107 3007
rect 3193 3294 3207 3308
rect 3253 3293 3267 3307
rect 3433 3772 3447 3786
rect 3453 3753 3467 3767
rect 3393 3693 3407 3707
rect 3373 3553 3387 3567
rect 3373 3532 3387 3546
rect 3133 3252 3147 3266
rect 3173 3252 3187 3266
rect 3313 3294 3327 3308
rect 3353 3294 3367 3308
rect 3293 3253 3307 3267
rect 3273 3213 3287 3227
rect 3213 3193 3227 3207
rect 3333 3233 3347 3247
rect 3433 3373 3447 3387
rect 3473 3713 3487 3727
rect 3553 3853 3567 3867
rect 3593 3833 3607 3847
rect 3553 3713 3567 3727
rect 3493 3693 3507 3707
rect 3513 3673 3527 3687
rect 3493 3633 3507 3647
rect 3473 3613 3487 3627
rect 3513 3513 3527 3527
rect 3633 3833 3647 3847
rect 3813 4512 3827 4526
rect 3793 4413 3807 4427
rect 3913 4673 3927 4687
rect 3853 4593 3867 4607
rect 3873 4554 3887 4568
rect 4013 4793 4027 4807
rect 3933 4633 3947 4647
rect 3853 4512 3867 4526
rect 3833 4493 3847 4507
rect 3893 4413 3907 4427
rect 3833 4393 3847 4407
rect 3773 4293 3787 4307
rect 3733 4193 3747 4207
rect 3733 4113 3747 4127
rect 3773 4093 3787 4107
rect 3733 4073 3747 4087
rect 3713 4053 3727 4067
rect 3853 4334 3867 4348
rect 3813 4173 3827 4187
rect 3793 4073 3807 4087
rect 3893 4213 3907 4227
rect 3993 4733 4007 4747
rect 3973 4552 3987 4566
rect 4073 4853 4087 4867
rect 4213 5074 4227 5088
rect 4253 5074 4267 5088
rect 4193 5032 4207 5046
rect 4233 5032 4247 5046
rect 4233 4993 4247 5007
rect 4213 4933 4227 4947
rect 4153 4893 4167 4907
rect 4213 4893 4227 4907
rect 4153 4854 4167 4868
rect 4193 4854 4207 4868
rect 4073 4812 4087 4826
rect 4133 4812 4147 4826
rect 4173 4812 4187 4826
rect 4093 4732 4107 4746
rect 4073 4713 4087 4727
rect 4073 4673 4087 4687
rect 4053 4653 4067 4667
rect 4053 4632 4067 4646
rect 4013 4593 4027 4607
rect 4013 4554 4027 4568
rect 4093 4613 4107 4627
rect 4153 4653 4167 4667
rect 4133 4613 4147 4627
rect 3973 4433 3987 4447
rect 4033 4512 4047 4526
rect 4133 4473 4147 4487
rect 4033 4453 4047 4467
rect 4073 4453 4087 4467
rect 4013 4433 4027 4447
rect 4013 4333 4027 4347
rect 3973 4273 3987 4287
rect 3953 4253 3967 4267
rect 3913 4193 3927 4207
rect 3893 4172 3907 4186
rect 3913 4153 3927 4167
rect 3833 4133 3847 4147
rect 3893 4133 3907 4147
rect 3893 4073 3907 4087
rect 3793 4033 3807 4047
rect 3873 4034 3887 4048
rect 3913 4034 3927 4048
rect 3673 3993 3687 4007
rect 3713 3973 3727 3987
rect 3793 3993 3807 4007
rect 3753 3933 3767 3947
rect 3693 3833 3707 3847
rect 3613 3753 3627 3767
rect 3593 3673 3607 3687
rect 3593 3652 3607 3666
rect 3713 3733 3727 3747
rect 3733 3673 3747 3687
rect 3673 3633 3687 3647
rect 3713 3633 3727 3647
rect 3633 3593 3647 3607
rect 3633 3553 3647 3567
rect 3693 3533 3707 3547
rect 3633 3514 3647 3528
rect 3733 3553 3747 3567
rect 3713 3513 3727 3527
rect 3733 3493 3747 3507
rect 3473 3433 3487 3447
rect 3453 3353 3467 3367
rect 3433 3333 3447 3347
rect 3473 3294 3487 3308
rect 3453 3233 3467 3247
rect 3493 3213 3507 3227
rect 3413 3193 3427 3207
rect 3473 3193 3487 3207
rect 3313 3173 3327 3187
rect 3373 3173 3387 3187
rect 3213 3153 3227 3167
rect 3293 3153 3307 3167
rect 3213 3113 3227 3127
rect 3193 3093 3207 3107
rect 3173 2994 3187 3008
rect 3133 2952 3147 2966
rect 3093 2933 3107 2947
rect 3073 2913 3087 2927
rect 3053 2793 3067 2807
rect 3153 2913 3167 2927
rect 3193 2893 3207 2907
rect 3273 3073 3287 3087
rect 3413 3172 3427 3186
rect 3373 3133 3387 3147
rect 3353 3113 3367 3127
rect 3313 2994 3327 3008
rect 3233 2952 3247 2966
rect 3253 2933 3267 2947
rect 3233 2853 3247 2867
rect 3213 2813 3227 2827
rect 3073 2732 3087 2746
rect 3013 2593 3027 2607
rect 3073 2593 3087 2607
rect 2993 2474 3007 2488
rect 2853 2432 2867 2446
rect 3013 2432 3027 2446
rect 3273 2813 3287 2827
rect 3333 2953 3347 2967
rect 3333 2913 3347 2927
rect 3293 2773 3307 2787
rect 3473 3113 3487 3127
rect 3533 3472 3547 3486
rect 3613 3473 3627 3487
rect 3713 3473 3727 3487
rect 3893 3973 3907 3987
rect 3813 3953 3827 3967
rect 3793 3933 3807 3947
rect 3833 3913 3847 3927
rect 3773 3853 3787 3867
rect 3873 3893 3887 3907
rect 4013 4253 4027 4267
rect 3993 4213 4007 4227
rect 4013 4193 4027 4207
rect 3993 4173 4007 4187
rect 3973 4133 3987 4147
rect 4133 4193 4147 4207
rect 4033 4153 4047 4167
rect 4073 4153 4087 4167
rect 4113 4153 4127 4167
rect 4013 4133 4027 4147
rect 3993 4073 4007 4087
rect 4013 4053 4027 4067
rect 4053 4053 4067 4067
rect 4033 4034 4047 4048
rect 3973 3993 3987 4007
rect 3912 3913 3926 3927
rect 3933 3913 3947 3927
rect 3893 3853 3907 3867
rect 3873 3833 3887 3847
rect 3792 3753 3806 3767
rect 3813 3753 3827 3767
rect 3933 3833 3947 3847
rect 4013 3933 4027 3947
rect 4033 3893 4047 3907
rect 4193 4593 4207 4607
rect 4273 4893 4287 4907
rect 4413 5173 4427 5187
rect 4373 5074 4387 5088
rect 4553 5552 4567 5566
rect 4593 5552 4607 5566
rect 4593 5531 4607 5545
rect 4553 5493 4567 5507
rect 4513 5373 4527 5387
rect 4673 5633 4687 5647
rect 4713 5633 4727 5647
rect 4653 5593 4667 5607
rect 4713 5594 4727 5608
rect 4773 5594 4787 5608
rect 4693 5552 4707 5566
rect 4733 5552 4747 5566
rect 4633 5493 4647 5507
rect 4693 5473 4707 5487
rect 4593 5373 4607 5387
rect 5013 6114 5027 6128
rect 5093 6114 5107 6128
rect 5153 6114 5167 6128
rect 5413 6153 5427 6167
rect 5313 6114 5327 6128
rect 4993 6072 5007 6086
rect 5033 6072 5047 6086
rect 5133 6072 5147 6086
rect 4933 6033 4947 6047
rect 5093 6033 5107 6047
rect 5073 6013 5087 6027
rect 5033 5953 5047 5967
rect 4893 5933 4907 5947
rect 4953 5933 4967 5947
rect 4853 5894 4867 5908
rect 4893 5894 4907 5908
rect 4993 5894 5007 5908
rect 5093 5993 5107 6007
rect 5073 5893 5087 5907
rect 4813 5852 4827 5866
rect 4913 5852 4927 5866
rect 4953 5852 4967 5866
rect 5013 5852 5027 5866
rect 5153 6033 5167 6047
rect 5133 5973 5147 5987
rect 5113 5953 5127 5967
rect 5293 6072 5307 6086
rect 5173 6013 5187 6027
rect 5373 6073 5387 6087
rect 5373 6033 5387 6047
rect 5513 6133 5527 6147
rect 5653 6133 5667 6147
rect 5413 6073 5427 6087
rect 5453 6072 5467 6086
rect 5493 6072 5507 6086
rect 5573 6072 5587 6086
rect 5393 6013 5407 6027
rect 5493 6013 5507 6027
rect 5433 5993 5447 6007
rect 5333 5933 5347 5947
rect 5413 5933 5427 5947
rect 5193 5894 5207 5908
rect 5373 5894 5387 5908
rect 5253 5873 5267 5887
rect 5113 5813 5127 5827
rect 5113 5753 5127 5767
rect 4933 5733 4947 5747
rect 4873 5693 4887 5707
rect 4873 5633 4887 5647
rect 4833 5594 4847 5608
rect 4913 5613 4927 5627
rect 4913 5573 4927 5587
rect 4853 5552 4867 5566
rect 4913 5552 4927 5566
rect 4873 5513 4887 5527
rect 4533 5332 4547 5346
rect 4593 5333 4607 5347
rect 4533 5312 4547 5326
rect 4573 5153 4587 5167
rect 4353 4993 4367 5007
rect 4413 4993 4427 5007
rect 4393 4973 4407 4987
rect 4353 4913 4367 4927
rect 4313 4893 4327 4907
rect 4373 4893 4387 4907
rect 4293 4873 4307 4887
rect 4273 4854 4287 4868
rect 4233 4813 4247 4827
rect 4473 5074 4487 5088
rect 4513 5074 4527 5088
rect 4493 5032 4507 5046
rect 4533 5032 4547 5046
rect 4573 5033 4587 5047
rect 4493 4993 4507 5007
rect 4433 4933 4447 4947
rect 4433 4854 4447 4868
rect 4513 4933 4527 4947
rect 4373 4793 4387 4807
rect 4412 4793 4426 4807
rect 4433 4793 4447 4807
rect 4393 4773 4407 4787
rect 4333 4753 4347 4767
rect 4333 4732 4347 4746
rect 4293 4693 4307 4707
rect 4333 4693 4347 4707
rect 4233 4613 4247 4627
rect 4213 4573 4227 4587
rect 4173 4553 4187 4567
rect 4273 4573 4287 4587
rect 4213 4512 4227 4526
rect 4253 4413 4267 4427
rect 4213 4334 4227 4348
rect 4253 4293 4267 4307
rect 4233 4133 4247 4147
rect 4153 4053 4167 4067
rect 4213 4053 4227 4067
rect 4093 4034 4107 4048
rect 4133 4034 4147 4048
rect 4193 4033 4207 4047
rect 4113 3992 4127 4006
rect 4073 3973 4087 3987
rect 4153 3973 4167 3987
rect 4173 3893 4187 3907
rect 3793 3713 3807 3727
rect 3773 3693 3787 3707
rect 3853 3733 3867 3747
rect 3813 3673 3827 3687
rect 4033 3833 4047 3847
rect 4053 3814 4067 3828
rect 4113 3814 4127 3828
rect 4153 3814 4167 3828
rect 3993 3772 4007 3786
rect 4033 3773 4047 3787
rect 3933 3633 3947 3647
rect 3873 3593 3887 3607
rect 3853 3533 3867 3547
rect 3573 3413 3587 3427
rect 3693 3433 3707 3447
rect 3613 3373 3627 3387
rect 3533 3353 3547 3367
rect 3513 3173 3527 3187
rect 3553 3333 3567 3347
rect 3633 3333 3647 3347
rect 3533 3093 3547 3107
rect 3493 3073 3507 3087
rect 3433 2994 3447 3008
rect 3473 2994 3487 3008
rect 3533 2994 3547 3008
rect 3693 3294 3707 3308
rect 3573 3252 3587 3266
rect 3613 3233 3627 3247
rect 3593 3033 3607 3047
rect 3553 2953 3567 2967
rect 3533 2933 3547 2947
rect 3433 2913 3447 2927
rect 3473 2893 3487 2907
rect 3433 2853 3447 2867
rect 3413 2813 3427 2827
rect 3413 2773 3427 2787
rect 3253 2713 3267 2727
rect 3213 2693 3227 2707
rect 3273 2693 3287 2707
rect 3193 2553 3207 2567
rect 3133 2474 3147 2488
rect 3253 2474 3267 2488
rect 3093 2393 3107 2407
rect 3213 2393 3227 2407
rect 3253 2393 3267 2407
rect 2773 2333 2787 2347
rect 2713 2313 2727 2327
rect 2733 2293 2747 2307
rect 2713 2273 2727 2287
rect 2693 2253 2707 2267
rect 2793 2273 2807 2287
rect 2673 2193 2687 2207
rect 2693 2133 2707 2147
rect 2653 2113 2667 2127
rect 2753 2193 2767 2207
rect 2773 2153 2787 2167
rect 2733 2113 2747 2127
rect 2713 2093 2727 2107
rect 2593 2053 2607 2067
rect 2653 2013 2667 2027
rect 2593 1973 2607 1987
rect 2713 1993 2727 2007
rect 2533 1833 2547 1847
rect 2693 1954 2707 1968
rect 2693 1893 2707 1907
rect 2453 1734 2467 1748
rect 2433 1673 2447 1687
rect 2393 1653 2407 1667
rect 2553 1813 2567 1827
rect 2573 1793 2587 1807
rect 2833 2313 2847 2327
rect 2913 2313 2927 2327
rect 2853 2293 2867 2307
rect 2852 2253 2866 2267
rect 2873 2254 2887 2268
rect 2973 2293 2987 2307
rect 2973 2254 2987 2268
rect 2853 2213 2867 2227
rect 2833 2173 2847 2187
rect 2813 2153 2827 2167
rect 2933 2212 2947 2226
rect 2893 2173 2907 2187
rect 2933 2173 2947 2187
rect 2853 2093 2867 2107
rect 2793 2033 2807 2047
rect 2813 1993 2827 2007
rect 3013 2113 3027 2127
rect 2993 1993 3007 2007
rect 2972 1954 2986 1968
rect 2993 1953 3007 1967
rect 2873 1913 2887 1927
rect 2913 1912 2927 1926
rect 2793 1833 2807 1847
rect 2733 1793 2747 1807
rect 2513 1733 2527 1747
rect 2593 1734 2607 1748
rect 2493 1633 2507 1647
rect 2373 1573 2387 1587
rect 2673 1733 2687 1747
rect 2733 1734 2747 1748
rect 2573 1692 2587 1706
rect 2533 1633 2547 1647
rect 2533 1593 2547 1607
rect 2593 1593 2607 1607
rect 2573 1513 2587 1527
rect 2513 1493 2527 1507
rect 2373 1473 2387 1487
rect 2353 1453 2367 1467
rect 2413 1433 2427 1447
rect 2493 1433 2507 1447
rect 2533 1434 2547 1448
rect 2433 1413 2447 1427
rect 2313 1392 2327 1406
rect 2393 1392 2407 1406
rect 2353 1293 2367 1307
rect 2293 1233 2307 1247
rect 2353 1233 2367 1247
rect 2313 1214 2327 1228
rect 2393 1372 2407 1386
rect 2513 1392 2527 1406
rect 2473 1373 2487 1387
rect 2553 1353 2567 1367
rect 2433 1293 2447 1307
rect 2493 1293 2507 1307
rect 2393 1233 2407 1247
rect 2453 1233 2467 1247
rect 2273 1173 2287 1187
rect 2333 1172 2347 1186
rect 2273 1133 2287 1147
rect 2413 1214 2427 1228
rect 2653 1692 2667 1706
rect 2713 1692 2727 1706
rect 2713 1633 2727 1647
rect 2773 1692 2787 1706
rect 2713 1553 2727 1567
rect 2673 1513 2687 1527
rect 2613 1493 2627 1507
rect 2633 1473 2647 1487
rect 2673 1434 2687 1448
rect 2693 1393 2707 1407
rect 2653 1353 2667 1367
rect 2693 1353 2707 1367
rect 2673 1313 2687 1327
rect 2633 1293 2647 1307
rect 2593 1273 2607 1287
rect 2573 1253 2587 1267
rect 2493 1214 2507 1228
rect 2553 1212 2567 1226
rect 2593 1214 2607 1228
rect 2693 1253 2707 1267
rect 2673 1213 2687 1227
rect 2513 1172 2527 1186
rect 2413 1133 2427 1147
rect 2413 1093 2427 1107
rect 2493 1093 2507 1107
rect 2293 1053 2307 1067
rect 2393 1053 2407 1067
rect 2273 1013 2287 1027
rect 2253 953 2267 967
rect 2373 1013 2387 1027
rect 2353 933 2367 947
rect 2373 913 2387 927
rect 2433 933 2447 947
rect 2273 872 2287 886
rect 2193 694 2207 708
rect 2233 694 2247 708
rect 1993 653 2007 667
rect 1973 613 1987 627
rect 1933 573 1947 587
rect 1833 513 1847 527
rect 1753 493 1767 507
rect 1793 493 1807 507
rect 1953 473 1967 487
rect 1873 413 1887 427
rect 1793 394 1807 408
rect 1913 394 1927 408
rect 2073 613 2087 627
rect 2033 573 2047 587
rect 2233 653 2247 667
rect 2193 533 2207 547
rect 2173 493 2187 507
rect 2013 473 2027 487
rect 1993 413 2007 427
rect 2033 394 2047 408
rect 2073 394 2087 408
rect 2113 394 2127 408
rect 1753 352 1767 366
rect 1813 352 1827 366
rect 1873 352 1887 366
rect 1933 352 1947 366
rect 1973 352 1987 366
rect 2013 353 2027 367
rect 1653 293 1667 307
rect 1733 293 1747 307
rect 1793 293 1807 307
rect 2033 293 2047 307
rect 1533 253 1547 267
rect 1553 233 1567 247
rect 1673 233 1687 247
rect 1533 213 1547 227
rect 2093 273 2107 287
rect 1813 233 1827 247
rect 1793 213 1807 227
rect 1813 193 1827 207
rect 1713 174 1727 188
rect 1873 173 1887 187
rect 1913 174 1927 188
rect 1973 174 1987 188
rect 1613 153 1627 167
rect 1533 132 1547 146
rect 1573 132 1587 146
rect 1493 113 1507 127
rect 1653 132 1667 146
rect 1693 132 1707 146
rect 1793 132 1807 146
rect 1573 93 1587 107
rect 1613 93 1627 107
rect 2053 174 2067 188
rect 2133 174 2147 188
rect 2353 873 2367 887
rect 2413 872 2427 886
rect 2453 872 2467 886
rect 2313 813 2327 827
rect 2333 733 2347 747
rect 2373 694 2387 708
rect 2453 694 2467 708
rect 2613 1172 2627 1186
rect 2573 1133 2587 1147
rect 2653 1133 2667 1147
rect 2753 1613 2767 1627
rect 2853 1853 2867 1867
rect 2953 1853 2967 1867
rect 3193 2293 3207 2307
rect 3073 2212 3087 2226
rect 3053 2173 3067 2187
rect 3093 2193 3107 2207
rect 3073 2153 3087 2167
rect 3193 2193 3207 2207
rect 3313 2732 3327 2746
rect 3353 2693 3367 2707
rect 3293 2633 3307 2647
rect 3433 2713 3447 2727
rect 3413 2533 3427 2547
rect 3513 2713 3527 2727
rect 3493 2653 3507 2667
rect 3473 2593 3487 2607
rect 3453 2513 3467 2527
rect 3333 2474 3347 2488
rect 3453 2474 3467 2488
rect 3493 2474 3507 2488
rect 3553 2733 3567 2747
rect 3533 2553 3547 2567
rect 3833 3473 3847 3487
rect 3833 3413 3847 3427
rect 3813 3393 3827 3407
rect 3733 3373 3747 3387
rect 3713 3133 3727 3147
rect 3713 3093 3727 3107
rect 3653 2994 3667 3008
rect 3613 2953 3627 2967
rect 3773 3294 3787 3308
rect 3813 3294 3827 3308
rect 3833 3253 3847 3267
rect 3793 3193 3807 3207
rect 3933 3514 3947 3528
rect 3993 3751 4007 3765
rect 3973 3513 3987 3527
rect 3873 3472 3887 3486
rect 3913 3472 3927 3486
rect 3953 3472 3967 3486
rect 3873 3433 3887 3447
rect 3913 3333 3927 3347
rect 4093 3772 4107 3786
rect 4073 3753 4087 3767
rect 4113 3753 4127 3767
rect 4153 3753 4167 3767
rect 4053 3673 4067 3687
rect 4033 3633 4047 3647
rect 4013 3533 4027 3547
rect 3993 3433 4007 3447
rect 4073 3514 4087 3528
rect 4313 4554 4327 4568
rect 4373 4733 4387 4747
rect 4373 4553 4387 4567
rect 4333 4512 4347 4526
rect 4293 4453 4307 4467
rect 4273 4073 4287 4087
rect 4273 4034 4287 4048
rect 4493 4753 4507 4767
rect 4433 4693 4447 4707
rect 4493 4633 4507 4647
rect 4433 4593 4447 4607
rect 4413 4512 4427 4526
rect 4473 4512 4487 4526
rect 4393 4473 4407 4487
rect 4373 4413 4387 4427
rect 4493 4493 4507 4507
rect 4413 4353 4427 4367
rect 4333 4334 4347 4348
rect 4393 4333 4407 4347
rect 4353 4292 4367 4306
rect 4393 4292 4407 4306
rect 4533 4873 4547 4887
rect 4713 5332 4727 5346
rect 4753 5333 4767 5347
rect 4673 5313 4687 5327
rect 4673 5193 4687 5207
rect 4613 5074 4627 5088
rect 4833 5374 4847 5388
rect 4813 5293 4827 5307
rect 4773 5133 4787 5147
rect 4813 5133 4827 5147
rect 4693 5093 4707 5107
rect 4793 5093 4807 5107
rect 4713 5072 4727 5086
rect 4753 5074 4767 5088
rect 4693 5032 4707 5046
rect 4633 4973 4647 4987
rect 4713 4973 4727 4987
rect 4773 4993 4787 5007
rect 4733 4953 4747 4967
rect 4773 4953 4787 4967
rect 4653 4854 4667 4868
rect 4573 4812 4587 4826
rect 4653 4813 4667 4827
rect 4613 4773 4627 4787
rect 4612 4633 4626 4647
rect 4633 4633 4647 4647
rect 4573 4593 4587 4607
rect 4553 4553 4567 4567
rect 4633 4573 4647 4587
rect 4553 4512 4567 4526
rect 4533 4453 4547 4467
rect 4533 4333 4547 4347
rect 4313 4073 4327 4087
rect 4372 4173 4386 4187
rect 4393 4173 4407 4187
rect 4373 4113 4387 4127
rect 4213 3953 4227 3967
rect 4193 3873 4207 3887
rect 4253 3992 4267 4006
rect 4313 3992 4327 4006
rect 4353 4033 4367 4047
rect 4453 4292 4467 4306
rect 4493 4292 4507 4306
rect 4533 4292 4547 4306
rect 4633 4512 4647 4526
rect 4593 4473 4607 4487
rect 4653 4433 4667 4447
rect 4633 4353 4647 4367
rect 4593 4334 4607 4348
rect 4693 4893 4707 4907
rect 4733 4854 4747 4868
rect 4753 4793 4767 4807
rect 4693 4773 4707 4787
rect 4693 4752 4707 4766
rect 4693 4513 4707 4527
rect 4693 4473 4707 4487
rect 4673 4333 4687 4347
rect 4513 4253 4527 4267
rect 4553 4253 4567 4267
rect 4453 4193 4467 4207
rect 4433 4034 4447 4048
rect 4333 3953 4347 3967
rect 4253 3933 4267 3947
rect 4193 3814 4207 3828
rect 4333 3793 4347 3807
rect 4293 3772 4307 3786
rect 4473 4173 4487 4187
rect 4413 3953 4427 3967
rect 4453 3953 4467 3967
rect 4373 3913 4387 3927
rect 4393 3893 4407 3907
rect 4433 3893 4447 3907
rect 4373 3873 4387 3887
rect 4373 3813 4387 3827
rect 4513 4153 4527 4167
rect 4653 4292 4667 4306
rect 4673 4273 4687 4287
rect 4613 4253 4627 4267
rect 4513 4113 4527 4127
rect 4573 4113 4587 4127
rect 4753 4493 4767 4507
rect 4713 4393 4727 4407
rect 4773 4413 4787 4427
rect 5393 5853 5407 5867
rect 5353 5833 5367 5847
rect 5313 5813 5327 5827
rect 5253 5793 5267 5807
rect 5213 5773 5227 5787
rect 5173 5713 5187 5727
rect 5113 5653 5127 5667
rect 5133 5633 5147 5647
rect 4993 5594 5007 5608
rect 5093 5594 5107 5608
rect 5193 5633 5207 5647
rect 5173 5613 5187 5627
rect 4973 5552 4987 5566
rect 5153 5552 5167 5566
rect 4933 5473 4947 5487
rect 4953 5374 4967 5388
rect 4993 5374 5007 5388
rect 5053 5374 5067 5388
rect 5133 5374 5147 5388
rect 4973 5313 4987 5327
rect 4913 5293 4927 5307
rect 5013 5253 5027 5267
rect 4953 5213 4967 5227
rect 5053 5213 5067 5227
rect 4893 5093 4907 5107
rect 4913 5032 4927 5046
rect 4873 4973 4887 4987
rect 4833 4953 4847 4967
rect 5133 5313 5147 5327
rect 5113 5153 5127 5167
rect 5033 5093 5047 5107
rect 5073 5074 5087 5088
rect 5113 5074 5127 5088
rect 5333 5653 5347 5667
rect 5313 5633 5327 5647
rect 5213 5553 5227 5567
rect 5233 5553 5247 5567
rect 5293 5513 5307 5527
rect 5253 5413 5267 5427
rect 5313 5393 5327 5407
rect 5293 5373 5307 5387
rect 5233 5332 5247 5346
rect 5273 5332 5287 5346
rect 5193 5293 5207 5307
rect 5253 5293 5267 5307
rect 5153 5253 5167 5267
rect 5153 5074 5167 5088
rect 5193 5074 5207 5088
rect 4973 5053 4987 5067
rect 5353 5613 5367 5627
rect 5493 5933 5507 5947
rect 5533 5894 5547 5908
rect 5633 6072 5647 6086
rect 5753 6173 5767 6187
rect 5793 6133 5807 6147
rect 5873 6113 5887 6127
rect 6113 6153 6127 6167
rect 6213 6153 6227 6167
rect 6093 6133 6107 6147
rect 6053 6114 6067 6128
rect 5593 5933 5607 5947
rect 5613 5894 5627 5908
rect 5473 5833 5487 5847
rect 5533 5793 5547 5807
rect 5513 5693 5527 5707
rect 5633 5773 5647 5787
rect 5593 5713 5607 5727
rect 5433 5653 5447 5667
rect 5413 5613 5427 5627
rect 5433 5594 5447 5608
rect 5493 5594 5507 5608
rect 5353 5433 5367 5447
rect 5393 5433 5407 5447
rect 5353 5393 5367 5407
rect 5493 5553 5507 5567
rect 5573 5594 5587 5608
rect 5613 5594 5627 5608
rect 5653 5594 5667 5608
rect 5553 5552 5567 5566
rect 5633 5553 5647 5567
rect 5513 5513 5527 5527
rect 5553 5513 5567 5527
rect 5593 5513 5607 5527
rect 5453 5493 5467 5507
rect 5413 5393 5427 5407
rect 5473 5393 5487 5407
rect 5373 5332 5387 5346
rect 5413 5293 5427 5307
rect 5393 5253 5407 5267
rect 5313 5213 5327 5227
rect 5313 5153 5327 5167
rect 5353 5113 5367 5127
rect 4973 4993 4987 5007
rect 5053 5032 5067 5046
rect 5113 5033 5127 5047
rect 5173 5032 5187 5046
rect 5253 5033 5267 5047
rect 5353 5074 5367 5088
rect 5413 5213 5427 5227
rect 5393 5073 5407 5087
rect 5013 4933 5027 4947
rect 4873 4913 4887 4927
rect 4953 4913 4967 4927
rect 5033 4893 5047 4907
rect 4893 4812 4907 4826
rect 4993 4854 5007 4868
rect 5033 4854 5047 4868
rect 4973 4833 4987 4847
rect 5273 5013 5287 5027
rect 5313 5013 5327 5027
rect 5213 4993 5227 5007
rect 5273 4933 5287 4947
rect 5233 4893 5247 4907
rect 5373 4993 5387 5007
rect 5333 4973 5347 4987
rect 5513 5374 5527 5388
rect 5613 5373 5627 5387
rect 5573 5332 5587 5346
rect 5773 6072 5787 6086
rect 5733 6053 5747 6067
rect 5733 6032 5747 6046
rect 6133 6114 6147 6128
rect 6173 6114 6187 6128
rect 6253 6114 6267 6128
rect 6293 6114 6307 6128
rect 6073 6072 6087 6086
rect 6113 6073 6127 6087
rect 6033 6033 6047 6047
rect 6113 6033 6127 6047
rect 6193 6072 6207 6086
rect 6153 6053 6167 6067
rect 5953 6013 5967 6027
rect 6013 6013 6027 6027
rect 6073 6013 6087 6027
rect 5893 5993 5907 6007
rect 5873 5953 5887 5967
rect 5793 5894 5807 5908
rect 5833 5894 5847 5908
rect 5693 5753 5707 5767
rect 5753 5773 5767 5787
rect 5793 5733 5807 5747
rect 5713 5693 5727 5707
rect 5713 5633 5727 5647
rect 5813 5633 5827 5647
rect 5693 5593 5707 5607
rect 5753 5594 5767 5608
rect 5733 5552 5747 5566
rect 5673 5453 5687 5467
rect 5673 5413 5687 5427
rect 5653 5373 5667 5387
rect 5633 5333 5647 5347
rect 5693 5332 5707 5346
rect 5853 5594 5867 5608
rect 5973 5852 5987 5866
rect 5933 5753 5947 5767
rect 6073 5913 6087 5927
rect 6213 5973 6227 5987
rect 6153 5893 6167 5907
rect 6053 5852 6067 5866
rect 6113 5833 6127 5847
rect 6013 5813 6027 5827
rect 6093 5813 6107 5827
rect 5973 5733 5987 5747
rect 5973 5633 5987 5647
rect 6073 5633 6087 5647
rect 5933 5594 5947 5608
rect 5833 5552 5847 5566
rect 5873 5552 5887 5566
rect 5953 5553 5967 5567
rect 5913 5513 5927 5527
rect 6033 5594 6047 5608
rect 5993 5553 6007 5567
rect 5973 5533 5987 5547
rect 5813 5493 5827 5507
rect 5953 5493 5967 5507
rect 5773 5433 5787 5447
rect 5893 5433 5907 5447
rect 5793 5374 5807 5388
rect 5833 5374 5847 5388
rect 6013 5533 6027 5547
rect 5993 5453 6007 5467
rect 5893 5353 5907 5367
rect 5813 5332 5827 5346
rect 5973 5332 5987 5346
rect 5933 5313 5947 5327
rect 6053 5513 6067 5527
rect 6133 5793 6147 5807
rect 6193 5833 6207 5847
rect 6233 5793 6247 5807
rect 6253 5653 6267 5667
rect 6213 5633 6227 5647
rect 6153 5593 6167 5607
rect 6253 5593 6267 5607
rect 6153 5553 6167 5567
rect 6133 5512 6147 5526
rect 6153 5493 6167 5507
rect 6033 5473 6047 5487
rect 6112 5473 6126 5487
rect 6133 5473 6147 5487
rect 6093 5374 6107 5388
rect 6153 5373 6167 5387
rect 6073 5332 6087 5346
rect 5693 5293 5707 5307
rect 5753 5293 5767 5307
rect 5833 5293 5847 5307
rect 5693 5173 5707 5187
rect 5473 5133 5487 5147
rect 5593 5133 5607 5147
rect 5433 5093 5447 5107
rect 5493 5093 5507 5107
rect 5533 5074 5547 5088
rect 5573 5074 5587 5088
rect 5353 4893 5367 4907
rect 5413 4893 5427 4907
rect 5133 4812 5147 4826
rect 5193 4813 5207 4827
rect 5253 4812 5267 4826
rect 4853 4793 4867 4807
rect 4993 4793 5007 4807
rect 4853 4733 4867 4747
rect 4873 4613 4887 4627
rect 5073 4773 5087 4787
rect 5253 4773 5267 4787
rect 5293 4773 5307 4787
rect 4953 4713 4967 4727
rect 5033 4673 5047 4687
rect 5153 4673 5167 4687
rect 5193 4673 5207 4687
rect 4993 4593 5007 4607
rect 4953 4554 4967 4568
rect 4833 4533 4847 4547
rect 4813 4373 4827 4387
rect 4893 4473 4907 4487
rect 4873 4433 4887 4447
rect 4753 4353 4767 4367
rect 4913 4373 4927 4387
rect 4813 4334 4827 4348
rect 4873 4334 4887 4348
rect 4753 4292 4767 4306
rect 4713 4233 4727 4247
rect 4833 4273 4847 4287
rect 4793 4253 4807 4267
rect 4813 4233 4827 4247
rect 4753 4173 4767 4187
rect 4693 4153 4707 4167
rect 4853 4233 4867 4247
rect 4873 4193 4887 4207
rect 4893 4173 4907 4187
rect 4833 4073 4847 4087
rect 4513 4034 4527 4048
rect 4553 3992 4567 4006
rect 4513 3893 4527 3907
rect 4493 3853 4507 3867
rect 4473 3813 4487 3827
rect 4353 3772 4367 3786
rect 4173 3713 4187 3727
rect 4313 3633 4327 3647
rect 4193 3613 4207 3627
rect 4153 3533 4167 3547
rect 4113 3513 4127 3527
rect 4273 3553 4287 3567
rect 4453 3772 4467 3786
rect 4493 3772 4507 3786
rect 4393 3733 4407 3747
rect 4353 3613 4367 3627
rect 4373 3573 4387 3587
rect 4353 3514 4367 3528
rect 4093 3413 4107 3427
rect 4013 3393 4027 3407
rect 4053 3393 4067 3407
rect 4053 3313 4067 3327
rect 3933 3294 3947 3308
rect 4033 3293 4047 3307
rect 4293 3472 4307 3486
rect 4353 3473 4367 3487
rect 4173 3413 4187 3427
rect 4113 3313 4127 3327
rect 4333 3313 4347 3327
rect 4013 3272 4027 3286
rect 3913 3252 3927 3266
rect 4033 3252 4047 3266
rect 4073 3252 4087 3266
rect 3873 3233 3887 3247
rect 3933 3213 3947 3227
rect 3833 3153 3847 3167
rect 3873 3153 3887 3167
rect 3793 3133 3807 3147
rect 3733 3033 3747 3047
rect 3833 3113 3847 3127
rect 3853 3093 3867 3107
rect 3833 2994 3847 3008
rect 3733 2973 3747 2987
rect 3713 2893 3727 2907
rect 3773 2893 3787 2907
rect 3733 2853 3747 2867
rect 3673 2813 3687 2827
rect 3933 3033 3947 3047
rect 4013 3033 4027 3047
rect 3993 2994 4007 3008
rect 4013 2953 4027 2967
rect 3913 2893 3927 2907
rect 3853 2833 3867 2847
rect 3793 2793 3807 2807
rect 3773 2773 3787 2787
rect 3593 2653 3607 2667
rect 3633 2733 3647 2747
rect 3613 2633 3627 2647
rect 3573 2533 3587 2547
rect 3533 2473 3547 2487
rect 3573 2474 3587 2488
rect 3313 2432 3327 2446
rect 3353 2413 3367 2427
rect 3273 2353 3287 2367
rect 3333 2353 3347 2367
rect 3233 2333 3247 2347
rect 3313 2313 3327 2327
rect 3273 2293 3287 2307
rect 3233 2273 3247 2287
rect 3333 2253 3347 2267
rect 3253 2212 3267 2226
rect 3293 2212 3307 2226
rect 3213 2173 3227 2187
rect 3153 2113 3167 2127
rect 3053 2073 3067 2087
rect 3333 2073 3347 2087
rect 3113 2033 3127 2047
rect 3173 2033 3187 2047
rect 3153 2013 3167 2027
rect 3033 1993 3047 2007
rect 3073 1993 3087 2007
rect 3113 1993 3127 2007
rect 3153 1953 3167 1967
rect 3213 1993 3227 2007
rect 3313 1953 3327 1967
rect 3013 1833 3027 1847
rect 2973 1813 2987 1827
rect 2893 1773 2907 1787
rect 2953 1773 2967 1787
rect 2853 1734 2867 1748
rect 2813 1712 2827 1726
rect 2813 1653 2827 1667
rect 2873 1692 2887 1706
rect 2913 1692 2927 1706
rect 2833 1613 2847 1627
rect 2793 1593 2807 1607
rect 2873 1593 2887 1607
rect 2773 1573 2787 1587
rect 2813 1533 2827 1547
rect 2773 1473 2787 1487
rect 2793 1392 2807 1406
rect 2833 1392 2847 1406
rect 2893 1473 2907 1487
rect 2953 1473 2967 1487
rect 2733 1373 2747 1387
rect 2873 1392 2887 1406
rect 3173 1912 3187 1926
rect 3093 1873 3107 1887
rect 3233 1873 3247 1887
rect 3073 1833 3087 1847
rect 3053 1793 3067 1807
rect 3033 1734 3047 1748
rect 3013 1692 3027 1706
rect 3213 1773 3227 1787
rect 3113 1753 3127 1767
rect 3153 1734 3167 1748
rect 3133 1692 3147 1706
rect 3173 1692 3187 1706
rect 3173 1653 3187 1667
rect 3433 2393 3447 2407
rect 3453 2353 3467 2367
rect 3533 2413 3547 2427
rect 3553 2393 3567 2407
rect 3613 2393 3627 2407
rect 3473 2333 3487 2347
rect 3453 2273 3467 2287
rect 3393 2212 3407 2226
rect 3513 2273 3527 2287
rect 3473 2253 3487 2267
rect 3733 2732 3747 2746
rect 3753 2713 3767 2727
rect 3673 2573 3687 2587
rect 3653 2533 3667 2547
rect 3713 2553 3727 2567
rect 3673 2293 3687 2307
rect 3913 2713 3927 2727
rect 3833 2633 3847 2647
rect 3833 2533 3847 2547
rect 4013 2893 4027 2907
rect 4133 3252 4147 3266
rect 4073 3113 4087 3127
rect 4113 3113 4127 3127
rect 4053 2994 4067 3008
rect 4213 3252 4227 3266
rect 4493 3713 4507 3727
rect 4413 3514 4427 3528
rect 4473 3514 4487 3528
rect 4453 3472 4467 3486
rect 4413 3293 4427 3307
rect 4613 4034 4627 4048
rect 4653 4034 4667 4048
rect 4693 4034 4707 4048
rect 4593 3973 4607 3987
rect 4553 3873 4567 3887
rect 4573 3853 4587 3867
rect 4753 4032 4767 4046
rect 4875 4053 4889 4067
rect 5033 4613 5047 4627
rect 5113 4613 5127 4627
rect 5013 4513 5027 4527
rect 4973 4373 4987 4387
rect 4953 4334 4967 4348
rect 4933 4292 4947 4306
rect 4993 4273 5007 4287
rect 4933 4213 4947 4227
rect 4953 4113 4967 4127
rect 4833 4034 4847 4048
rect 4913 4034 4927 4048
rect 5233 4593 5247 4607
rect 5153 4493 5167 4507
rect 5113 4473 5127 4487
rect 5113 4452 5127 4466
rect 5053 4413 5067 4427
rect 5053 4373 5067 4387
rect 5033 4273 5047 4287
rect 5253 4493 5267 4507
rect 5213 4473 5227 4487
rect 5193 4413 5207 4427
rect 5173 4334 5187 4348
rect 5093 4292 5107 4306
rect 5133 4293 5147 4307
rect 5053 4093 5067 4107
rect 5013 4073 5027 4087
rect 5133 4233 5147 4247
rect 5133 4193 5147 4207
rect 5133 4093 5147 4107
rect 5113 4053 5127 4067
rect 4993 4034 5007 4048
rect 4633 3973 4647 3987
rect 4553 3772 4567 3786
rect 4593 3772 4607 3786
rect 4613 3733 4627 3747
rect 4593 3693 4607 3707
rect 4553 3673 4567 3687
rect 4573 3653 4587 3667
rect 4613 3653 4627 3667
rect 4553 3613 4567 3627
rect 4613 3613 4627 3627
rect 4613 3553 4627 3567
rect 4773 3993 4787 4007
rect 4753 3973 4767 3987
rect 4813 3992 4827 4006
rect 4773 3893 4787 3907
rect 4973 3913 4987 3927
rect 4713 3853 4727 3867
rect 4753 3853 4767 3867
rect 4853 3853 4867 3867
rect 4673 3833 4687 3847
rect 4713 3814 4727 3828
rect 4693 3753 4707 3767
rect 4813 3833 4827 3847
rect 4773 3813 4787 3827
rect 4893 3873 4907 3887
rect 4873 3833 4887 3847
rect 4993 3853 5007 3867
rect 5033 3853 5047 3867
rect 4773 3772 4787 3786
rect 4833 3772 4847 3786
rect 4873 3772 4887 3786
rect 4953 3833 4967 3847
rect 4993 3832 5007 3846
rect 5093 4034 5107 4048
rect 5313 4713 5327 4727
rect 5393 4854 5407 4868
rect 5413 4812 5427 4826
rect 5473 5032 5487 5046
rect 5513 5032 5527 5046
rect 5493 4993 5507 5007
rect 5573 4993 5587 5007
rect 5473 4953 5487 4967
rect 5453 4773 5467 4787
rect 5393 4673 5407 4687
rect 5373 4633 5387 4647
rect 5353 4573 5367 4587
rect 5373 4554 5387 4568
rect 5733 5113 5747 5127
rect 5673 5074 5687 5088
rect 5793 5074 5807 5088
rect 5693 5032 5707 5046
rect 5733 5033 5747 5047
rect 5653 4993 5667 5007
rect 5693 4973 5707 4987
rect 5593 4953 5607 4967
rect 5533 4913 5547 4927
rect 5493 4853 5507 4867
rect 5573 4854 5587 4868
rect 5613 4854 5627 4868
rect 5653 4854 5667 4868
rect 5553 4812 5567 4826
rect 5673 4812 5687 4826
rect 5513 4653 5527 4667
rect 5413 4573 5427 4587
rect 5293 4453 5307 4467
rect 5373 4413 5387 4427
rect 5273 4353 5287 4367
rect 5313 4353 5327 4367
rect 5353 4353 5367 4367
rect 5273 4292 5287 4306
rect 5233 4233 5247 4247
rect 5153 4033 5167 4047
rect 5273 4073 5287 4087
rect 5173 4013 5187 4027
rect 5073 3993 5087 4007
rect 5053 3813 5067 3827
rect 4953 3772 4967 3786
rect 5013 3772 5027 3786
rect 4933 3753 4947 3767
rect 5093 3913 5107 3927
rect 5073 3653 5087 3667
rect 4753 3553 4767 3567
rect 4793 3553 4807 3567
rect 4953 3553 4967 3567
rect 4693 3513 4707 3527
rect 4753 3514 4767 3528
rect 4513 3472 4527 3486
rect 4553 3453 4567 3467
rect 4533 3373 4547 3387
rect 4513 3333 4527 3347
rect 4393 3253 4407 3267
rect 4153 3213 4167 3227
rect 4373 3213 4387 3227
rect 4353 3173 4367 3187
rect 4313 3153 4327 3167
rect 4233 3014 4247 3028
rect 4093 2994 4107 3008
rect 4133 2994 4147 3008
rect 4173 2994 4187 3008
rect 4233 2994 4247 3008
rect 4273 2994 4287 3008
rect 4113 2952 4127 2966
rect 4073 2933 4087 2947
rect 3973 2793 3987 2807
rect 4033 2793 4047 2807
rect 4013 2774 4027 2788
rect 4033 2732 4047 2746
rect 4333 3113 4347 3127
rect 4093 2833 4107 2847
rect 4133 2793 4147 2807
rect 4093 2773 4107 2787
rect 4153 2732 4167 2746
rect 4253 2913 4267 2927
rect 4233 2873 4247 2887
rect 4213 2853 4227 2867
rect 3993 2713 4007 2727
rect 4113 2713 4127 2727
rect 4193 2713 4207 2727
rect 3973 2513 3987 2527
rect 3893 2473 3907 2487
rect 3933 2473 3947 2487
rect 3973 2474 3987 2488
rect 3793 2353 3807 2367
rect 3773 2313 3787 2327
rect 3653 2253 3667 2267
rect 3753 2253 3767 2267
rect 3793 2293 3807 2307
rect 3493 2193 3507 2207
rect 3553 2193 3567 2207
rect 3373 2173 3387 2187
rect 3433 2173 3447 2187
rect 3473 2173 3487 2187
rect 3353 2033 3367 2047
rect 3373 1954 3387 1968
rect 3413 1954 3427 1968
rect 3333 1833 3347 1847
rect 3313 1773 3327 1787
rect 3273 1753 3287 1767
rect 3233 1733 3247 1747
rect 3393 1873 3407 1887
rect 3353 1793 3367 1807
rect 3453 1813 3467 1827
rect 3433 1773 3447 1787
rect 3373 1734 3387 1748
rect 3433 1733 3447 1747
rect 3233 1653 3247 1667
rect 3333 1693 3347 1707
rect 3393 1692 3407 1706
rect 3293 1633 3307 1647
rect 3073 1593 3087 1607
rect 3213 1593 3227 1607
rect 3413 1593 3427 1607
rect 3213 1533 3227 1547
rect 3033 1493 3047 1507
rect 2973 1453 2987 1467
rect 2953 1434 2967 1448
rect 2993 1434 3007 1448
rect 2913 1392 2927 1406
rect 2853 1353 2867 1367
rect 2893 1353 2907 1367
rect 2893 1313 2907 1327
rect 2973 1392 2987 1406
rect 2813 1273 2827 1287
rect 2933 1273 2947 1287
rect 2873 1253 2887 1267
rect 2713 1214 2727 1228
rect 2753 1214 2767 1228
rect 2813 1214 2827 1228
rect 2773 1133 2787 1147
rect 2793 1093 2807 1107
rect 2713 1013 2727 1027
rect 2593 993 2607 1007
rect 2693 993 2707 1007
rect 2553 973 2567 987
rect 2553 933 2567 947
rect 2513 913 2527 927
rect 2653 973 2667 987
rect 2533 873 2547 887
rect 2533 833 2547 847
rect 2513 813 2527 827
rect 2613 853 2627 867
rect 2573 833 2587 847
rect 2593 813 2607 827
rect 2633 813 2647 827
rect 2733 953 2747 967
rect 2733 914 2747 928
rect 2713 833 2727 847
rect 2733 813 2747 827
rect 2753 793 2767 807
rect 2553 753 2567 767
rect 2653 753 2667 767
rect 2713 753 2727 767
rect 2313 652 2327 666
rect 2253 533 2267 547
rect 2333 513 2347 527
rect 2233 453 2247 467
rect 2273 433 2287 447
rect 2213 394 2227 408
rect 2533 693 2547 707
rect 2433 513 2447 527
rect 2373 473 2387 487
rect 2513 652 2527 666
rect 2613 733 2627 747
rect 2573 693 2587 707
rect 2653 694 2667 708
rect 2473 433 2487 447
rect 2473 394 2487 408
rect 2353 352 2367 366
rect 2453 352 2467 366
rect 2493 352 2507 366
rect 2233 313 2247 327
rect 2393 273 2407 287
rect 2233 233 2247 247
rect 2333 213 2347 227
rect 2253 173 2267 187
rect 2293 174 2307 188
rect 2233 153 2247 167
rect 2033 132 2047 146
rect 1973 93 1987 107
rect 2153 73 2167 87
rect 2213 133 2227 147
rect 1873 33 1887 47
rect 2193 33 2207 47
rect 2233 113 2247 127
rect 2453 174 2467 188
rect 2493 174 2507 188
rect 2353 113 2367 127
rect 2393 132 2407 146
rect 2433 132 2447 146
rect 2473 132 2487 146
rect 2253 73 2267 87
rect 2553 473 2567 487
rect 2553 393 2567 407
rect 2673 652 2687 666
rect 2753 733 2767 747
rect 2853 1093 2867 1107
rect 2813 933 2827 947
rect 2853 914 2867 928
rect 3073 1434 3087 1448
rect 3273 1453 3287 1467
rect 3333 1434 3347 1448
rect 3373 1433 3387 1447
rect 3633 2212 3647 2226
rect 3613 2193 3627 2207
rect 3593 2173 3607 2187
rect 3613 2153 3627 2167
rect 3733 2212 3747 2226
rect 3773 2212 3787 2226
rect 3853 2254 3867 2268
rect 3873 2213 3887 2227
rect 3673 2113 3687 2127
rect 3793 2113 3807 2127
rect 3833 2113 3847 2127
rect 3873 2113 3887 2127
rect 3633 2073 3647 2087
rect 3613 2033 3627 2047
rect 3553 2013 3567 2027
rect 3673 2013 3687 2027
rect 3713 1954 3727 1968
rect 3813 1954 3827 1968
rect 3533 1912 3547 1926
rect 3693 1912 3707 1926
rect 3813 1913 3827 1927
rect 4353 3033 4367 3047
rect 4373 3013 4387 3027
rect 4433 3253 4447 3267
rect 4453 3113 4467 3127
rect 4433 3073 4447 3087
rect 4633 3453 4647 3467
rect 4633 3373 4647 3387
rect 4593 3333 4607 3347
rect 4553 3293 4567 3307
rect 4673 3294 4687 3308
rect 4533 3252 4547 3266
rect 4513 3073 4527 3087
rect 4513 2994 4527 3008
rect 4393 2952 4407 2966
rect 4433 2953 4447 2967
rect 4573 3252 4587 3266
rect 4573 3073 4587 3087
rect 4553 2952 4567 2966
rect 4433 2913 4447 2927
rect 4333 2873 4347 2887
rect 4773 3333 4787 3347
rect 4853 3514 4867 3528
rect 4893 3514 4907 3528
rect 4973 3514 4987 3528
rect 5053 3514 5067 3528
rect 4873 3472 4887 3486
rect 4953 3473 4967 3487
rect 4813 3433 4827 3447
rect 4793 3313 4807 3327
rect 5013 3472 5027 3486
rect 4973 3413 4987 3427
rect 4833 3373 4847 3387
rect 4873 3353 4887 3367
rect 4953 3353 4967 3367
rect 4853 3333 4867 3347
rect 4833 3293 4847 3307
rect 4793 3213 4807 3227
rect 4913 3313 4927 3327
rect 5253 3992 5267 4006
rect 5273 3933 5287 3947
rect 5193 3893 5207 3907
rect 5113 3873 5127 3887
rect 5153 3873 5167 3887
rect 5173 3853 5187 3867
rect 5153 3833 5167 3847
rect 5213 3814 5227 3828
rect 5233 3793 5247 3807
rect 5113 3772 5127 3786
rect 5133 3553 5147 3567
rect 5173 3514 5187 3528
rect 5153 3472 5167 3486
rect 5133 3433 5147 3447
rect 4972 3313 4986 3327
rect 4993 3313 5007 3327
rect 5053 3313 5067 3327
rect 5093 3314 5107 3328
rect 4853 3193 4867 3207
rect 4753 3173 4767 3187
rect 4713 3093 4727 3107
rect 4853 3073 4867 3087
rect 4693 2994 4707 3008
rect 4733 2994 4747 3008
rect 4633 2952 4647 2966
rect 4893 3193 4907 3207
rect 4953 3233 4967 3247
rect 4933 3173 4947 3187
rect 4953 3073 4967 3087
rect 4873 3053 4887 3067
rect 4873 3032 4887 3046
rect 4633 2853 4647 2867
rect 4713 2853 4727 2867
rect 4513 2833 4527 2847
rect 4573 2833 4587 2847
rect 4393 2813 4407 2827
rect 4253 2774 4267 2788
rect 4373 2773 4387 2787
rect 4353 2732 4367 2746
rect 4373 2713 4387 2727
rect 4233 2573 4247 2587
rect 4293 2573 4307 2587
rect 4093 2493 4107 2507
rect 4113 2493 4127 2507
rect 4133 2474 4147 2488
rect 4173 2474 4187 2488
rect 4213 2474 4227 2488
rect 4253 2474 4267 2488
rect 4353 2493 4367 2507
rect 4453 2774 4467 2788
rect 4433 2713 4447 2727
rect 4393 2693 4407 2707
rect 4473 2693 4487 2707
rect 4393 2533 4407 2547
rect 3953 2432 3967 2446
rect 4033 2433 4047 2447
rect 3973 2313 3987 2327
rect 3913 2273 3927 2287
rect 4013 2273 4027 2287
rect 4073 2432 4087 2446
rect 4373 2473 4387 2487
rect 4113 2373 4127 2387
rect 4093 2333 4107 2347
rect 4053 2273 4067 2287
rect 4033 2253 4047 2267
rect 3933 2213 3947 2227
rect 3913 2173 3927 2187
rect 3913 2113 3927 2127
rect 3893 2093 3907 2107
rect 3913 2073 3927 2087
rect 4033 2173 4047 2187
rect 3993 2153 4007 2167
rect 3952 2113 3966 2127
rect 3973 2113 3987 2127
rect 3933 2053 3947 2067
rect 3953 2033 3967 2047
rect 3933 1993 3947 2007
rect 3993 1993 4007 2007
rect 3873 1973 3887 1987
rect 3973 1953 3987 1967
rect 3833 1893 3847 1907
rect 3533 1873 3547 1887
rect 3753 1873 3767 1887
rect 3513 1833 3527 1847
rect 3493 1753 3507 1767
rect 3473 1733 3487 1747
rect 4173 2273 4187 2287
rect 4133 2254 4147 2268
rect 4153 2212 4167 2226
rect 4233 2432 4247 2446
rect 4373 2433 4387 2447
rect 4213 2333 4227 2347
rect 4333 2333 4347 2347
rect 4373 2333 4387 2347
rect 4273 2254 4287 2268
rect 4213 2212 4227 2226
rect 4113 2193 4127 2207
rect 4193 2193 4207 2207
rect 4253 2212 4267 2226
rect 4293 2193 4307 2207
rect 4233 2173 4247 2187
rect 4053 2153 4067 2167
rect 4213 2153 4227 2167
rect 4113 2113 4127 2127
rect 4033 1954 4047 1968
rect 4073 1954 4087 1968
rect 4413 2493 4427 2507
rect 4573 2774 4587 2788
rect 4553 2732 4567 2746
rect 4653 2773 4667 2787
rect 4913 2994 4927 3008
rect 4933 2952 4947 2966
rect 4873 2853 4887 2867
rect 4913 2833 4927 2847
rect 4793 2813 4807 2827
rect 4853 2793 4867 2807
rect 4593 2713 4607 2727
rect 4633 2713 4647 2727
rect 4673 2753 4687 2767
rect 5013 3293 5027 3307
rect 5353 4292 5367 4306
rect 5393 4153 5407 4167
rect 5333 4053 5347 4067
rect 5493 4554 5507 4568
rect 5533 4553 5547 4567
rect 5533 4472 5547 4486
rect 5473 4413 5487 4427
rect 5453 4353 5467 4367
rect 5433 4333 5447 4347
rect 5493 4334 5507 4348
rect 5533 4333 5547 4347
rect 5433 4293 5447 4307
rect 5413 4053 5427 4067
rect 5513 4292 5527 4306
rect 5493 4273 5507 4287
rect 5473 4213 5487 4227
rect 5593 4554 5607 4568
rect 5633 4554 5647 4568
rect 5773 5013 5787 5027
rect 5773 4853 5787 4867
rect 5813 4854 5827 4868
rect 5853 5233 5867 5247
rect 5893 5094 5907 5108
rect 5853 5073 5867 5087
rect 5893 5074 5907 5088
rect 5893 5013 5907 5027
rect 5873 4933 5887 4947
rect 5853 4913 5867 4927
rect 5773 4813 5787 4827
rect 5753 4793 5767 4807
rect 5713 4733 5727 4747
rect 5833 4813 5847 4827
rect 5793 4733 5807 4747
rect 5773 4693 5787 4707
rect 5713 4673 5727 4687
rect 5813 4673 5827 4687
rect 6033 5313 6047 5327
rect 6093 5313 6107 5327
rect 6013 5093 6027 5107
rect 5973 5074 5987 5088
rect 5973 5013 5987 5027
rect 5913 4953 5927 4967
rect 6033 5032 6047 5046
rect 6013 4993 6027 5007
rect 5913 4893 5927 4907
rect 5893 4873 5907 4887
rect 5833 4653 5847 4667
rect 5713 4633 5727 4647
rect 5853 4633 5867 4647
rect 5833 4593 5847 4607
rect 5693 4554 5707 4568
rect 5733 4554 5747 4568
rect 5773 4554 5787 4568
rect 5753 4512 5767 4526
rect 5893 4812 5907 4826
rect 6013 4893 6027 4907
rect 6113 5233 6127 5247
rect 6213 5533 6227 5547
rect 6193 5473 6207 5487
rect 6193 5393 6207 5407
rect 6233 5473 6247 5487
rect 6233 5433 6247 5447
rect 6293 6053 6307 6067
rect 6373 6053 6387 6067
rect 6413 5973 6427 5987
rect 6393 5933 6407 5947
rect 6313 5893 6327 5907
rect 6353 5894 6367 5908
rect 6333 5653 6347 5667
rect 6373 5633 6387 5647
rect 6313 5594 6327 5608
rect 6353 5594 6367 5608
rect 6293 5553 6307 5567
rect 6273 5513 6287 5527
rect 6373 5553 6387 5567
rect 6333 5513 6347 5527
rect 6293 5433 6307 5447
rect 6253 5393 6267 5407
rect 6273 5374 6287 5388
rect 6193 5253 6207 5267
rect 6113 5133 6127 5147
rect 6173 5133 6187 5147
rect 6193 5113 6207 5127
rect 6133 5093 6147 5107
rect 6173 5074 6187 5088
rect 6253 5332 6267 5346
rect 6293 5332 6307 5346
rect 6253 5293 6267 5307
rect 6073 4953 6087 4967
rect 6193 5032 6207 5046
rect 6133 4993 6147 5007
rect 6173 5013 6187 5027
rect 6033 4873 6047 4887
rect 6013 4853 6027 4867
rect 6053 4854 6067 4868
rect 5953 4793 5967 4807
rect 5933 4753 5947 4767
rect 5933 4693 5947 4707
rect 5913 4673 5927 4687
rect 5913 4573 5927 4587
rect 5853 4553 5867 4567
rect 5893 4554 5907 4568
rect 5627 4493 5641 4507
rect 5693 4493 5707 4507
rect 5793 4493 5807 4507
rect 5853 4493 5867 4507
rect 5893 4493 5907 4507
rect 5593 4453 5607 4467
rect 5833 4453 5847 4467
rect 5873 4453 5887 4467
rect 5573 4413 5587 4427
rect 5573 4272 5587 4286
rect 5533 4213 5547 4227
rect 5793 4413 5807 4427
rect 5833 4413 5847 4427
rect 5613 4373 5627 4387
rect 5733 4353 5747 4367
rect 5693 4292 5707 4306
rect 5633 4273 5647 4287
rect 5613 4253 5627 4267
rect 5593 4233 5607 4247
rect 5633 4233 5647 4247
rect 5613 4213 5627 4227
rect 5613 4173 5627 4187
rect 5593 4153 5607 4167
rect 5373 3992 5387 4006
rect 5413 3992 5427 4006
rect 5333 3873 5347 3887
rect 5393 3873 5407 3887
rect 5453 3873 5467 3887
rect 5353 3853 5367 3867
rect 5313 3814 5327 3828
rect 5333 3772 5347 3786
rect 5333 3693 5347 3707
rect 5413 3853 5427 3867
rect 5513 4034 5527 4048
rect 5593 4033 5607 4047
rect 5493 3993 5507 4007
rect 5513 3873 5527 3887
rect 5493 3853 5507 3867
rect 5453 3814 5467 3828
rect 5493 3753 5507 3767
rect 5493 3573 5507 3587
rect 5353 3513 5367 3527
rect 5393 3514 5407 3528
rect 5273 3472 5287 3486
rect 5333 3473 5347 3487
rect 5233 3353 5247 3367
rect 5293 3353 5307 3367
rect 5353 3353 5367 3367
rect 5093 3293 5107 3307
rect 5133 3293 5147 3307
rect 5033 3193 5047 3207
rect 5213 3312 5227 3326
rect 5173 3293 5187 3307
rect 5253 3313 5267 3327
rect 5113 3233 5127 3247
rect 5153 3233 5167 3247
rect 5233 3193 5247 3207
rect 5073 3173 5087 3187
rect 5133 3173 5147 3187
rect 5173 3173 5187 3187
rect 5013 3013 5027 3027
rect 5013 2992 5027 3006
rect 5053 2994 5067 3008
rect 5093 2994 5107 3008
rect 4953 2793 4967 2807
rect 4993 2793 5007 2807
rect 4653 2693 4667 2707
rect 4753 2673 4767 2687
rect 4553 2593 4567 2607
rect 4513 2474 4527 2488
rect 4473 2432 4487 2446
rect 4413 2373 4427 2387
rect 4433 2173 4447 2187
rect 4393 2153 4407 2167
rect 4433 2093 4447 2107
rect 4333 2033 4347 2047
rect 4133 1953 4147 1967
rect 4173 1954 4187 1968
rect 4213 1954 4227 1968
rect 4253 1954 4267 1968
rect 4113 1933 4127 1947
rect 4053 1912 4067 1926
rect 4093 1913 4107 1927
rect 3993 1833 4007 1847
rect 4073 1833 4087 1847
rect 3913 1813 3927 1827
rect 3973 1813 3987 1827
rect 3773 1793 3787 1807
rect 3733 1773 3747 1787
rect 3553 1734 3567 1748
rect 3613 1733 3627 1747
rect 3673 1734 3687 1748
rect 3453 1692 3467 1706
rect 3493 1692 3507 1706
rect 3533 1692 3547 1706
rect 3573 1692 3587 1706
rect 3513 1673 3527 1687
rect 3473 1653 3487 1667
rect 3433 1513 3447 1527
rect 3473 1453 3487 1467
rect 3273 1392 3287 1406
rect 3313 1392 3327 1406
rect 3093 1353 3107 1367
rect 3033 1253 3047 1267
rect 2993 1214 3007 1228
rect 3033 1214 3047 1228
rect 3073 1214 3087 1228
rect 3113 1214 3127 1228
rect 3153 1214 3167 1228
rect 2973 1172 2987 1186
rect 3033 1173 3047 1187
rect 3153 1133 3167 1147
rect 3093 1093 3107 1107
rect 3193 1373 3207 1387
rect 3253 1253 3267 1267
rect 3213 1214 3227 1228
rect 3233 1172 3247 1186
rect 3433 1253 3447 1267
rect 3533 1653 3547 1667
rect 3713 1693 3727 1707
rect 3693 1653 3707 1667
rect 3573 1633 3587 1647
rect 3633 1513 3647 1527
rect 3553 1473 3567 1487
rect 3533 1453 3547 1467
rect 3613 1434 3627 1448
rect 3533 1392 3547 1406
rect 3593 1392 3607 1406
rect 3473 1373 3487 1387
rect 3513 1373 3527 1387
rect 3453 1233 3467 1247
rect 3353 1093 3367 1107
rect 3433 1173 3447 1187
rect 3393 1073 3407 1087
rect 3393 993 3407 1007
rect 3213 953 3227 967
rect 2953 933 2967 947
rect 2873 872 2887 886
rect 2833 853 2847 867
rect 2793 694 2807 708
rect 2773 633 2787 647
rect 2873 793 2887 807
rect 2913 872 2927 886
rect 2933 833 2947 847
rect 2913 813 2927 827
rect 2893 753 2907 767
rect 2913 713 2927 727
rect 2893 694 2907 708
rect 3053 914 3067 928
rect 3113 914 3127 928
rect 3153 914 3167 928
rect 3033 853 3047 867
rect 2973 833 2987 847
rect 3053 833 3067 847
rect 3113 853 3127 867
rect 2953 813 2967 827
rect 3093 813 3107 827
rect 2973 753 2987 767
rect 3053 694 3067 708
rect 2913 652 2927 666
rect 2973 652 2987 666
rect 3173 853 3187 867
rect 3133 813 3147 827
rect 3213 813 3227 827
rect 3273 914 3287 928
rect 3293 872 3307 886
rect 3333 872 3347 886
rect 3153 713 3167 727
rect 3193 694 3207 708
rect 2873 633 2887 647
rect 2633 613 2647 627
rect 2713 613 2727 627
rect 2833 613 2847 627
rect 2873 612 2887 626
rect 3033 613 3047 627
rect 2833 473 2847 487
rect 2773 433 2787 447
rect 2573 352 2587 366
rect 2553 313 2567 327
rect 2673 394 2687 408
rect 3013 533 3027 547
rect 2913 453 2927 467
rect 2873 394 2887 408
rect 2773 352 2787 366
rect 2813 352 2827 366
rect 2853 352 2867 366
rect 2713 333 2727 347
rect 2653 313 2667 327
rect 2593 253 2607 267
rect 2973 394 2987 408
rect 2953 253 2967 267
rect 2853 233 2867 247
rect 2913 233 2927 247
rect 2593 213 2607 227
rect 2653 213 2667 227
rect 2713 213 2727 227
rect 2553 173 2567 187
rect 2693 174 2707 188
rect 2553 133 2567 147
rect 2533 33 2547 47
rect 2753 193 2767 207
rect 2733 174 2747 188
rect 2953 232 2967 246
rect 2913 193 2927 207
rect 2853 173 2867 187
rect 2753 133 2767 147
rect 2993 213 3007 227
rect 3173 652 3187 666
rect 3233 653 3247 667
rect 3213 633 3227 647
rect 3153 593 3167 607
rect 3153 533 3167 547
rect 3093 493 3107 507
rect 3093 453 3107 467
rect 3033 413 3047 427
rect 3113 413 3127 427
rect 3073 394 3087 408
rect 3253 633 3267 647
rect 3033 353 3047 367
rect 3073 233 3087 247
rect 3013 193 3027 207
rect 3073 193 3087 207
rect 2993 173 3007 187
rect 3253 313 3267 327
rect 3133 213 3147 227
rect 2833 132 2847 146
rect 2873 132 2887 146
rect 2933 132 2947 146
rect 2973 132 2987 146
rect 3013 132 3027 146
rect 3073 132 3087 146
rect 3193 194 3207 208
rect 3193 174 3207 188
rect 3233 173 3247 187
rect 3333 694 3347 708
rect 3353 633 3367 647
rect 3313 553 3327 567
rect 3373 433 3387 447
rect 3333 352 3347 366
rect 3133 133 3147 147
rect 3233 133 3247 147
rect 2733 93 2747 107
rect 2793 93 2807 107
rect 3113 93 3127 107
rect 2713 73 2727 87
rect 3093 73 3107 87
rect 3133 73 3147 87
rect 3313 174 3327 188
rect 3453 1153 3467 1167
rect 3673 1473 3687 1487
rect 3833 1734 3847 1748
rect 3793 1692 3807 1706
rect 3793 1493 3807 1507
rect 3733 1453 3747 1467
rect 3713 1434 3727 1448
rect 3793 1434 3807 1448
rect 3833 1434 3847 1448
rect 3873 1434 3887 1448
rect 3733 1392 3747 1406
rect 3673 1353 3687 1367
rect 3793 1353 3807 1367
rect 3673 1273 3687 1287
rect 3853 1273 3867 1287
rect 4053 1734 4067 1748
rect 4013 1692 4027 1706
rect 3953 1673 3967 1687
rect 4193 1912 4207 1926
rect 4133 1893 4147 1907
rect 4253 1893 4267 1907
rect 4133 1813 4147 1827
rect 4513 2053 4527 2067
rect 4513 1993 4527 2007
rect 4493 1954 4507 1968
rect 4533 1954 4547 1968
rect 4313 1893 4327 1907
rect 4293 1833 4307 1847
rect 4273 1793 4287 1807
rect 4113 1734 4127 1748
rect 4073 1692 4087 1706
rect 4133 1692 4147 1706
rect 4013 1653 4027 1667
rect 4053 1653 4067 1667
rect 4093 1653 4107 1667
rect 4253 1692 4267 1706
rect 4433 1893 4447 1907
rect 4533 1913 4547 1927
rect 4473 1853 4487 1867
rect 4373 1793 4387 1807
rect 4353 1733 4367 1747
rect 5193 3013 5207 3027
rect 5273 2994 5287 3008
rect 5173 2952 5187 2966
rect 5133 2833 5147 2847
rect 5093 2773 5107 2787
rect 5153 2774 5167 2788
rect 5233 2793 5247 2807
rect 4993 2693 5007 2707
rect 5033 2673 5047 2687
rect 4953 2573 4967 2587
rect 5013 2573 5027 2587
rect 4913 2533 4927 2547
rect 4953 2533 4967 2547
rect 4673 2474 4687 2488
rect 4713 2474 4727 2488
rect 4753 2474 4767 2488
rect 4793 2474 4807 2488
rect 4833 2474 4847 2488
rect 4913 2474 4927 2488
rect 4573 2432 4587 2446
rect 4613 2393 4627 2407
rect 5173 2732 5187 2746
rect 5133 2673 5147 2687
rect 5093 2533 5107 2547
rect 5193 2533 5207 2547
rect 5213 2474 5227 2488
rect 4653 2373 4667 2387
rect 4713 2373 4727 2387
rect 4713 2254 4727 2268
rect 4813 2432 4827 2446
rect 4933 2432 4947 2446
rect 4973 2432 4987 2446
rect 5013 2432 5027 2446
rect 5033 2393 5047 2407
rect 5113 2393 5127 2407
rect 5053 2293 5067 2307
rect 4673 2212 4687 2226
rect 4773 2212 4787 2226
rect 4833 2212 4847 2226
rect 4593 2113 4607 2127
rect 4633 2113 4647 2127
rect 4933 2153 4947 2167
rect 4893 2113 4907 2127
rect 4733 2053 4747 2067
rect 4673 1993 4687 2007
rect 4593 1973 4607 1987
rect 4633 1954 4647 1968
rect 4673 1953 4687 1967
rect 4853 1954 4867 1968
rect 5033 2153 5047 2167
rect 4953 2113 4967 2127
rect 4933 1953 4947 1967
rect 4973 1954 4987 1968
rect 4613 1912 4627 1926
rect 4653 1853 4667 1867
rect 4493 1773 4507 1787
rect 4553 1773 4567 1787
rect 4413 1734 4427 1748
rect 4393 1692 4407 1706
rect 4313 1653 4327 1667
rect 4193 1633 4207 1647
rect 4253 1633 4267 1647
rect 4433 1533 4447 1547
rect 4473 1533 4487 1547
rect 4253 1493 4267 1507
rect 3953 1433 3967 1447
rect 4012 1434 4026 1448
rect 4033 1433 4047 1447
rect 4093 1434 4107 1448
rect 4173 1434 4187 1448
rect 3913 1233 3927 1247
rect 3573 1214 3587 1228
rect 3633 1212 3647 1226
rect 3693 1214 3707 1228
rect 3733 1214 3747 1228
rect 3513 1153 3527 1167
rect 3553 1133 3567 1147
rect 3513 1013 3527 1027
rect 3473 993 3487 1007
rect 3433 953 3447 967
rect 3633 1172 3647 1186
rect 3673 1172 3687 1186
rect 3613 1073 3627 1087
rect 3833 1133 3847 1147
rect 3973 1373 3987 1387
rect 3993 1273 4007 1287
rect 3973 1233 3987 1247
rect 3953 1113 3967 1127
rect 3833 1053 3847 1067
rect 3913 1053 3927 1067
rect 3673 1033 3687 1047
rect 3753 1033 3767 1047
rect 3673 993 3687 1007
rect 3693 914 3707 928
rect 4133 1353 4147 1367
rect 4233 1353 4247 1367
rect 4033 1233 4047 1247
rect 4073 1214 4087 1228
rect 3993 1172 4007 1186
rect 4053 1172 4067 1186
rect 4093 1133 4107 1147
rect 4193 1172 4207 1186
rect 4213 1153 4227 1167
rect 4133 1093 4147 1107
rect 4213 1093 4227 1107
rect 4133 1053 4147 1067
rect 3833 1013 3847 1027
rect 3933 1013 3947 1027
rect 3973 1013 3987 1027
rect 3793 914 3807 928
rect 3893 914 3907 928
rect 3593 853 3607 867
rect 3573 813 3587 827
rect 3633 813 3647 827
rect 3493 713 3507 727
rect 3593 713 3607 727
rect 3453 694 3467 708
rect 3433 652 3447 666
rect 3413 613 3427 627
rect 3473 613 3487 627
rect 3593 652 3607 666
rect 3433 473 3447 487
rect 3473 433 3487 447
rect 3433 394 3447 408
rect 3533 593 3547 607
rect 3773 872 3787 886
rect 3733 853 3747 867
rect 3693 793 3707 807
rect 3653 694 3667 708
rect 3713 694 3727 708
rect 3853 793 3867 807
rect 3913 713 3927 727
rect 3753 652 3767 666
rect 3833 652 3847 666
rect 3653 633 3667 647
rect 3753 553 3767 567
rect 3573 394 3587 408
rect 3593 353 3607 367
rect 3453 313 3467 327
rect 3393 273 3407 287
rect 3393 193 3407 207
rect 3533 193 3547 207
rect 3293 132 3307 146
rect 3333 132 3347 146
rect 3373 132 3387 146
rect 3453 174 3467 188
rect 3513 173 3527 187
rect 1393 13 1407 27
rect 1433 13 1447 27
rect 2213 13 2227 27
rect 2573 13 2587 27
rect 3513 132 3527 146
rect 3213 33 3227 47
rect 3473 33 3487 47
rect 3633 493 3647 507
rect 3613 193 3627 207
rect 3733 433 3747 447
rect 3693 352 3707 366
rect 3693 193 3707 207
rect 3633 174 3647 188
rect 3673 173 3687 187
rect 3573 132 3587 146
rect 3613 132 3627 146
rect 3753 393 3767 407
rect 3813 394 3827 408
rect 3913 393 3927 407
rect 3793 352 3807 366
rect 3813 293 3827 307
rect 3773 233 3787 247
rect 3753 193 3767 207
rect 3853 273 3867 287
rect 3913 253 3927 267
rect 3813 173 3827 187
rect 3693 132 3707 146
rect 3793 132 3807 146
rect 3833 132 3847 146
rect 3893 132 3907 146
rect 3753 73 3767 87
rect 3673 33 3687 47
rect 4413 1373 4427 1387
rect 4473 1373 4487 1387
rect 4353 1333 4367 1347
rect 4553 1734 4567 1748
rect 4593 1734 4607 1748
rect 4533 1692 4547 1706
rect 4573 1693 4587 1707
rect 4673 1734 4687 1748
rect 4653 1692 4667 1706
rect 4573 1613 4587 1627
rect 4593 1533 4607 1547
rect 4513 1513 4527 1527
rect 4573 1513 4587 1527
rect 4513 1473 4527 1487
rect 4633 1473 4647 1487
rect 4593 1434 4607 1448
rect 4613 1373 4627 1387
rect 4493 1313 4507 1327
rect 4253 1273 4267 1287
rect 4493 1273 4507 1287
rect 4113 993 4127 1007
rect 4233 993 4247 1007
rect 4093 933 4107 947
rect 3953 913 3967 927
rect 3953 872 3967 886
rect 4013 872 4027 886
rect 4093 873 4107 887
rect 4213 953 4227 967
rect 4353 1233 4367 1247
rect 4313 1214 4327 1228
rect 4372 1214 4386 1228
rect 4353 1193 4367 1207
rect 4393 1213 4407 1227
rect 4453 1214 4467 1228
rect 4373 1173 4387 1187
rect 4633 1333 4647 1347
rect 4713 1692 4727 1706
rect 4893 1692 4907 1706
rect 4773 1653 4787 1667
rect 4833 1653 4847 1667
rect 4793 1533 4807 1547
rect 4853 1533 4867 1547
rect 4733 1434 4747 1448
rect 4673 1293 4687 1307
rect 4733 1293 4747 1307
rect 4693 1214 4707 1228
rect 4433 1172 4447 1186
rect 4473 1172 4487 1186
rect 4313 1133 4327 1147
rect 4353 1133 4367 1147
rect 4393 1133 4407 1147
rect 4333 1113 4347 1127
rect 4293 1033 4307 1047
rect 4393 913 4407 927
rect 4573 1172 4587 1186
rect 4613 1172 4627 1186
rect 4513 1153 4527 1167
rect 4513 1013 4527 1027
rect 4473 914 4487 928
rect 4213 893 4227 907
rect 4153 853 4167 867
rect 4193 853 4207 867
rect 4013 713 4027 727
rect 3993 694 4007 708
rect 3973 613 3987 627
rect 4113 652 4127 666
rect 4053 613 4067 627
rect 4013 573 4027 587
rect 4013 493 4027 507
rect 3973 394 3987 408
rect 4033 394 4047 408
rect 4233 753 4247 767
rect 4173 693 4187 707
rect 4173 652 4187 666
rect 4253 573 4267 587
rect 4153 433 4167 447
rect 4053 393 4067 407
rect 4073 293 4087 307
rect 4173 394 4187 408
rect 4053 253 4067 267
rect 4153 253 4167 267
rect 4213 253 4227 267
rect 3953 233 3967 247
rect 4013 174 4027 188
rect 3953 132 3967 146
rect 3933 13 3947 27
rect 4013 13 4027 27
rect 4093 213 4107 227
rect 4153 193 4167 207
rect 4133 132 4147 146
rect 4293 793 4307 807
rect 4313 753 4327 767
rect 4353 694 4367 708
rect 4593 953 4607 967
rect 4673 953 4687 967
rect 4533 914 4547 928
rect 4513 793 4527 807
rect 4493 753 4507 767
rect 4453 693 4467 707
rect 5013 1734 5027 1748
rect 4953 1533 4967 1547
rect 4933 1434 4947 1448
rect 4873 1373 4887 1387
rect 4813 1214 4827 1228
rect 4893 1214 4907 1228
rect 4993 1434 5007 1448
rect 5033 1433 5047 1447
rect 5013 1313 5027 1327
rect 4793 1153 4807 1167
rect 4753 1013 4767 1027
rect 4773 914 4787 928
rect 4893 1093 4907 1107
rect 4913 1073 4927 1087
rect 4893 953 4907 967
rect 4613 872 4627 886
rect 4673 872 4687 886
rect 4573 853 4587 867
rect 4993 1133 5007 1147
rect 4933 993 4947 1007
rect 4933 953 4947 967
rect 4753 872 4767 886
rect 4913 873 4927 887
rect 5433 3353 5447 3367
rect 5413 3313 5427 3327
rect 5373 3294 5387 3308
rect 5473 3333 5487 3347
rect 5573 3992 5587 4006
rect 5613 3953 5627 3967
rect 5613 3932 5627 3946
rect 5553 3853 5567 3867
rect 5893 4373 5907 4387
rect 6013 4813 6027 4827
rect 5973 4753 5987 4767
rect 6073 4812 6087 4826
rect 6053 4793 6067 4807
rect 6053 4753 6067 4767
rect 5993 4733 6007 4747
rect 6033 4593 6047 4607
rect 5993 4553 6007 4567
rect 6073 4554 6087 4568
rect 5973 4513 5987 4527
rect 6013 4512 6027 4526
rect 6053 4512 6067 4526
rect 6093 4513 6107 4527
rect 5913 4353 5927 4367
rect 5793 4292 5807 4306
rect 5793 4233 5807 4247
rect 5792 4193 5806 4207
rect 5813 4193 5827 4207
rect 5773 4153 5787 4167
rect 5693 4133 5707 4147
rect 5773 4132 5787 4146
rect 5733 4053 5747 4067
rect 5673 3953 5687 3967
rect 5633 3913 5647 3927
rect 5893 4292 5907 4306
rect 5853 4153 5867 4167
rect 5913 4053 5927 4067
rect 5853 4034 5867 4048
rect 5793 3993 5807 4007
rect 5773 3933 5787 3947
rect 5833 3992 5847 4006
rect 5913 3992 5927 4006
rect 5953 4373 5967 4387
rect 6053 4473 6067 4487
rect 6093 4453 6107 4467
rect 6073 4413 6087 4427
rect 6053 4393 6067 4407
rect 6013 4334 6027 4348
rect 6053 4292 6067 4306
rect 5993 4213 6007 4227
rect 6053 4193 6067 4207
rect 5973 4133 5987 4147
rect 5993 4073 6007 4087
rect 5953 4053 5967 4067
rect 6173 4953 6187 4967
rect 6193 4854 6207 4868
rect 6153 4713 6167 4727
rect 6213 4812 6227 4826
rect 6193 4793 6207 4807
rect 6153 4673 6167 4687
rect 6173 4653 6187 4667
rect 6213 4593 6227 4607
rect 6193 4573 6207 4587
rect 6233 4573 6247 4587
rect 6273 5253 6287 5267
rect 6373 5493 6387 5507
rect 6353 5473 6367 5487
rect 6373 5373 6387 5387
rect 6353 5332 6367 5346
rect 6333 5293 6347 5307
rect 6293 5173 6307 5187
rect 6393 5233 6407 5247
rect 6373 5113 6387 5127
rect 6433 5894 6447 5908
rect 6433 5253 6447 5267
rect 6433 5113 6447 5127
rect 6273 5073 6287 5087
rect 6313 5074 6327 5088
rect 6353 5074 6367 5088
rect 6273 5032 6287 5046
rect 6293 5013 6307 5027
rect 6293 4933 6307 4947
rect 6273 4873 6287 4887
rect 6333 4873 6347 4887
rect 6293 4853 6307 4867
rect 6373 4873 6387 4887
rect 6413 5074 6427 5088
rect 6413 4973 6427 4987
rect 6393 4853 6407 4867
rect 6313 4812 6327 4826
rect 6393 4813 6407 4827
rect 6353 4773 6367 4787
rect 6353 4752 6367 4766
rect 6333 4713 6347 4727
rect 6353 4653 6367 4667
rect 6333 4573 6347 4587
rect 6273 4554 6287 4568
rect 6313 4554 6327 4568
rect 6153 4513 6167 4527
rect 6133 4413 6147 4427
rect 6233 4512 6247 4526
rect 6273 4513 6287 4527
rect 6213 4493 6227 4507
rect 6333 4512 6347 4526
rect 6193 4453 6207 4467
rect 6213 4373 6227 4387
rect 6213 4333 6227 4347
rect 6133 4292 6147 4306
rect 6173 4292 6187 4306
rect 6213 4292 6227 4306
rect 6293 4334 6307 4348
rect 6373 4373 6387 4387
rect 6333 4333 6347 4347
rect 6233 4153 6247 4167
rect 6193 4073 6207 4087
rect 6093 4053 6107 4067
rect 6133 4053 6147 4067
rect 6033 4033 6047 4047
rect 6073 4034 6087 4048
rect 6013 3993 6027 4007
rect 5973 3973 5987 3987
rect 5832 3933 5846 3947
rect 5853 3933 5867 3947
rect 5933 3933 5947 3947
rect 5793 3893 5807 3907
rect 5673 3853 5687 3867
rect 5713 3853 5727 3867
rect 5653 3814 5667 3828
rect 5713 3813 5727 3827
rect 5773 3814 5787 3828
rect 5553 3793 5567 3807
rect 5533 3773 5547 3787
rect 5593 3772 5607 3786
rect 5553 3752 5567 3766
rect 5713 3733 5727 3747
rect 5593 3593 5607 3607
rect 5793 3772 5807 3786
rect 5833 3772 5847 3786
rect 5753 3693 5767 3707
rect 5813 3593 5827 3607
rect 5533 3553 5547 3567
rect 5713 3553 5727 3567
rect 5793 3553 5807 3567
rect 5573 3514 5587 3528
rect 5633 3514 5647 3528
rect 5693 3514 5707 3528
rect 5553 3472 5567 3486
rect 5633 3473 5647 3487
rect 5713 3472 5727 3486
rect 5593 3393 5607 3407
rect 5573 3333 5587 3347
rect 5533 3294 5547 3308
rect 5633 3313 5647 3327
rect 5673 3294 5687 3308
rect 5393 3252 5407 3266
rect 5433 3252 5447 3266
rect 5353 3233 5367 3247
rect 5553 3252 5567 3266
rect 5593 3252 5607 3266
rect 5473 3193 5487 3207
rect 5373 3173 5387 3187
rect 5333 2994 5347 3008
rect 5453 3133 5467 3147
rect 5433 3093 5447 3107
rect 5293 2793 5307 2807
rect 5393 2952 5407 2966
rect 5493 3053 5507 3067
rect 5753 3433 5767 3447
rect 5873 3913 5887 3927
rect 5993 3913 6007 3927
rect 5933 3893 5947 3907
rect 5853 3553 5867 3567
rect 5853 3532 5867 3546
rect 5813 3513 5827 3527
rect 5873 3513 5887 3527
rect 5833 3472 5847 3486
rect 5873 3473 5887 3487
rect 5853 3393 5867 3407
rect 5733 3333 5747 3347
rect 5793 3333 5807 3347
rect 5853 3333 5867 3347
rect 5713 3153 5727 3167
rect 5653 3133 5667 3147
rect 5813 3313 5827 3327
rect 5753 3273 5767 3287
rect 5833 3193 5847 3207
rect 5733 3113 5747 3127
rect 5833 3093 5847 3107
rect 5593 3053 5607 3067
rect 5533 2994 5547 3008
rect 5633 2994 5647 3008
rect 5673 2994 5687 3008
rect 5733 2994 5747 3008
rect 5853 3013 5867 3027
rect 5873 2993 5887 3007
rect 5453 2952 5467 2966
rect 5433 2813 5447 2827
rect 5313 2774 5327 2788
rect 5293 2732 5307 2746
rect 5353 2653 5367 2667
rect 5293 2613 5307 2627
rect 5253 2473 5267 2487
rect 5313 2393 5327 2407
rect 5233 2293 5247 2307
rect 5273 2293 5287 2307
rect 5313 2293 5327 2307
rect 5133 2254 5147 2268
rect 5173 2254 5187 2268
rect 5213 2254 5227 2268
rect 5273 2254 5287 2268
rect 5433 2774 5447 2788
rect 5473 2774 5487 2788
rect 5593 2952 5607 2966
rect 5653 2952 5667 2966
rect 5733 2953 5747 2967
rect 5793 2952 5807 2966
rect 5833 2913 5847 2927
rect 5953 3772 5967 3786
rect 5913 3733 5927 3747
rect 5913 3533 5927 3547
rect 5973 3514 5987 3528
rect 6033 3933 6047 3947
rect 6053 3913 6067 3927
rect 6053 3853 6067 3867
rect 6013 3813 6027 3827
rect 6273 4273 6287 4287
rect 6313 4213 6327 4227
rect 6273 4113 6287 4127
rect 6133 3973 6147 3987
rect 6013 3773 6027 3787
rect 6113 3773 6127 3787
rect 6033 3733 6047 3747
rect 6173 3933 6187 3947
rect 6153 3873 6167 3887
rect 6133 3673 6147 3687
rect 6133 3593 6147 3607
rect 6033 3553 6047 3567
rect 6113 3553 6127 3567
rect 5953 3433 5967 3447
rect 6013 3433 6027 3447
rect 5973 3373 5987 3387
rect 5913 3313 5927 3327
rect 5953 3252 5967 3266
rect 5993 3252 6007 3266
rect 5933 3073 5947 3087
rect 6093 3514 6107 3528
rect 6253 3993 6267 4007
rect 6313 4093 6327 4107
rect 6373 4153 6387 4167
rect 6373 4093 6387 4107
rect 6313 4053 6327 4067
rect 6353 4053 6367 4067
rect 6333 4034 6347 4048
rect 6433 4893 6447 4907
rect 6433 4872 6447 4886
rect 6413 4773 6427 4787
rect 6413 4752 6427 4766
rect 6433 4653 6447 4667
rect 6433 4613 6447 4627
rect 6433 4513 6447 4527
rect 6433 4433 6447 4447
rect 6433 4373 6447 4387
rect 6412 4332 6426 4346
rect 6433 4333 6447 4347
rect 6433 4233 6447 4247
rect 6253 3933 6267 3947
rect 6213 3853 6227 3867
rect 6273 3853 6287 3867
rect 6193 3814 6207 3828
rect 6233 3814 6247 3828
rect 6253 3753 6267 3767
rect 6213 3713 6227 3727
rect 6173 3613 6187 3627
rect 6153 3573 6167 3587
rect 6053 3453 6067 3467
rect 6113 3472 6127 3486
rect 6073 3333 6087 3347
rect 6213 3593 6227 3607
rect 6253 3593 6267 3607
rect 6253 3553 6267 3567
rect 6213 3513 6227 3527
rect 6233 3472 6247 3486
rect 6273 3473 6287 3487
rect 6233 3433 6247 3447
rect 6193 3373 6207 3387
rect 6133 3313 6147 3327
rect 6173 3313 6187 3327
rect 6093 3193 6107 3207
rect 6093 3113 6107 3127
rect 6033 3013 6047 3027
rect 5913 2993 5927 3007
rect 5973 2952 5987 2966
rect 5913 2913 5927 2927
rect 5833 2892 5847 2906
rect 5893 2893 5907 2907
rect 5693 2833 5707 2847
rect 5813 2833 5827 2847
rect 5653 2813 5667 2827
rect 5453 2732 5467 2746
rect 5453 2693 5467 2707
rect 5513 2733 5527 2747
rect 5493 2613 5507 2627
rect 5433 2474 5447 2488
rect 5593 2774 5607 2788
rect 5753 2774 5767 2788
rect 5793 2773 5807 2787
rect 5613 2732 5627 2746
rect 5653 2732 5667 2746
rect 5573 2693 5587 2707
rect 5653 2693 5667 2707
rect 5773 2732 5787 2746
rect 5713 2653 5727 2667
rect 5813 2753 5827 2767
rect 5793 2613 5807 2627
rect 5793 2533 5807 2547
rect 5533 2513 5547 2527
rect 5653 2513 5667 2527
rect 5573 2474 5587 2488
rect 5413 2393 5427 2407
rect 5553 2313 5567 2327
rect 5593 2313 5607 2327
rect 5373 2273 5387 2287
rect 5393 2254 5407 2268
rect 5453 2253 5467 2267
rect 5513 2254 5527 2268
rect 5553 2254 5567 2268
rect 5233 2212 5247 2226
rect 5173 2173 5187 2187
rect 5093 2113 5107 2127
rect 5193 1993 5207 2007
rect 5313 2212 5327 2226
rect 5373 2193 5387 2207
rect 5353 2173 5367 2187
rect 5353 2033 5367 2047
rect 5293 2013 5307 2027
rect 5073 1833 5087 1847
rect 5173 1773 5187 1787
rect 5113 1754 5127 1768
rect 5113 1733 5127 1747
rect 5113 1653 5127 1667
rect 5153 1613 5167 1627
rect 5113 1573 5127 1587
rect 5113 1434 5127 1448
rect 5073 1273 5087 1287
rect 5053 1214 5067 1228
rect 5333 1954 5347 1968
rect 5493 2212 5507 2226
rect 5453 2153 5467 2167
rect 5573 2213 5587 2227
rect 5533 2133 5547 2147
rect 5413 2073 5427 2087
rect 5573 2073 5587 2087
rect 5293 1773 5307 1787
rect 5253 1734 5267 1748
rect 5333 1733 5347 1747
rect 5193 1692 5207 1706
rect 5233 1692 5247 1706
rect 5273 1673 5287 1687
rect 5433 2033 5447 2047
rect 5413 1873 5427 1887
rect 5573 2013 5587 2027
rect 5553 1973 5567 1987
rect 5493 1954 5507 1968
rect 5613 2293 5627 2307
rect 5693 2293 5707 2307
rect 5653 2254 5667 2268
rect 6213 3333 6227 3347
rect 6173 3252 6187 3266
rect 6213 3193 6227 3207
rect 6133 3093 6147 3107
rect 6233 3053 6247 3067
rect 6273 3053 6287 3067
rect 6032 2952 6046 2966
rect 6053 2953 6067 2967
rect 6333 3973 6347 3987
rect 6313 3893 6327 3907
rect 6353 3953 6367 3967
rect 6393 3893 6407 3907
rect 6353 3873 6367 3887
rect 6353 3852 6367 3866
rect 6333 3833 6347 3847
rect 6393 3813 6407 3827
rect 6313 3773 6327 3787
rect 6393 3773 6407 3787
rect 6373 3713 6387 3727
rect 6333 3673 6347 3687
rect 6353 3553 6367 3567
rect 6333 3513 6347 3527
rect 6433 3953 6447 3967
rect 6433 3853 6447 3867
rect 6413 3613 6427 3627
rect 6393 3533 6407 3547
rect 6433 3573 6447 3587
rect 6333 3473 6347 3487
rect 6373 3393 6387 3407
rect 6373 3333 6387 3347
rect 6333 3313 6347 3327
rect 6433 3393 6447 3407
rect 6413 3293 6427 3307
rect 6353 3252 6367 3266
rect 6393 3252 6407 3266
rect 6373 3093 6387 3107
rect 6293 3033 6307 3047
rect 6433 3073 6447 3087
rect 6373 2973 6387 2987
rect 5973 2873 5987 2887
rect 6013 2873 6027 2887
rect 5893 2774 5907 2788
rect 5933 2774 5947 2788
rect 5873 2732 5887 2746
rect 5913 2732 5927 2746
rect 6013 2833 6027 2847
rect 6033 2813 6047 2827
rect 6113 2952 6127 2966
rect 6153 2952 6167 2966
rect 6233 2952 6247 2966
rect 6113 2913 6127 2927
rect 6293 2913 6307 2927
rect 6053 2774 6067 2788
rect 5973 2533 5987 2547
rect 5973 2474 5987 2488
rect 6033 2474 6047 2488
rect 6073 2474 6087 2488
rect 6193 2873 6207 2887
rect 6293 2813 6307 2827
rect 6153 2693 6167 2707
rect 6313 2732 6327 2746
rect 6373 2733 6387 2747
rect 6173 2474 6187 2488
rect 6213 2474 6227 2488
rect 6273 2473 6287 2487
rect 6053 2432 6067 2446
rect 6113 2432 6127 2446
rect 5833 2373 5847 2387
rect 5873 2373 5887 2387
rect 5853 2293 5867 2307
rect 5733 2253 5747 2267
rect 5673 2212 5687 2226
rect 5713 2212 5727 2226
rect 5613 2173 5627 2187
rect 5853 2212 5867 2226
rect 5913 2333 5927 2347
rect 5973 2333 5987 2347
rect 5933 2254 5947 2268
rect 5813 2193 5827 2207
rect 5873 2193 5887 2207
rect 5933 2193 5947 2207
rect 5713 2153 5727 2167
rect 5753 2153 5767 2167
rect 5673 2073 5687 2087
rect 5633 1993 5647 2007
rect 5593 1973 5607 1987
rect 5833 2013 5847 2027
rect 5773 1973 5787 1987
rect 5713 1954 5727 1968
rect 5833 1954 5847 1968
rect 5553 1912 5567 1926
rect 5613 1912 5627 1926
rect 5593 1873 5607 1887
rect 5653 1873 5667 1887
rect 5473 1793 5487 1807
rect 5433 1773 5447 1787
rect 5493 1773 5507 1787
rect 5413 1734 5427 1748
rect 5473 1733 5487 1747
rect 5353 1653 5367 1667
rect 5433 1673 5447 1687
rect 5393 1613 5407 1627
rect 5553 1734 5567 1748
rect 5753 1813 5767 1827
rect 5653 1793 5667 1807
rect 5613 1753 5627 1767
rect 5593 1733 5607 1747
rect 5493 1693 5507 1707
rect 5533 1692 5547 1706
rect 5533 1613 5547 1627
rect 5393 1533 5407 1547
rect 5473 1533 5487 1547
rect 5233 1453 5247 1467
rect 5353 1453 5367 1467
rect 5173 1373 5187 1387
rect 5213 1333 5227 1347
rect 5213 1293 5227 1307
rect 5193 1273 5207 1287
rect 5153 1233 5167 1247
rect 5133 1214 5147 1228
rect 5113 1172 5127 1186
rect 5113 1093 5127 1107
rect 5113 1033 5127 1047
rect 5032 953 5046 967
rect 5053 953 5067 967
rect 5013 914 5027 928
rect 4993 853 5007 867
rect 4773 793 4787 807
rect 4933 793 4947 807
rect 4973 793 4987 807
rect 4673 733 4687 747
rect 4533 713 4547 727
rect 4633 713 4647 727
rect 4333 652 4347 666
rect 4373 652 4387 666
rect 4473 652 4487 666
rect 4593 694 4607 708
rect 4453 613 4467 627
rect 4293 394 4307 408
rect 4333 393 4347 407
rect 4393 394 4407 408
rect 4273 353 4287 367
rect 4313 273 4327 287
rect 4173 113 4187 127
rect 4213 113 4227 127
rect 4093 93 4107 107
rect 4133 93 4147 107
rect 4433 273 4447 287
rect 4513 473 4527 487
rect 4473 393 4487 407
rect 4573 652 4587 666
rect 4733 652 4747 666
rect 4673 613 4687 627
rect 4613 573 4627 587
rect 4693 493 4707 507
rect 4553 394 4567 408
rect 4613 394 4627 408
rect 4653 394 4667 408
rect 4853 753 4867 767
rect 4933 694 4947 708
rect 4973 694 4987 708
rect 5093 914 5107 928
rect 5173 1113 5187 1127
rect 5573 1593 5587 1607
rect 5613 1513 5627 1527
rect 5533 1473 5547 1487
rect 5513 1434 5527 1448
rect 5553 1434 5567 1448
rect 5373 1392 5387 1406
rect 5333 1373 5347 1387
rect 5513 1393 5527 1407
rect 5333 1333 5347 1347
rect 5433 1333 5447 1347
rect 5293 1293 5307 1307
rect 5273 1253 5287 1267
rect 5233 1233 5247 1247
rect 5573 1313 5587 1327
rect 5353 1253 5367 1267
rect 5333 1213 5347 1227
rect 5213 1172 5227 1186
rect 5273 1172 5287 1186
rect 5313 1172 5327 1186
rect 5353 1172 5367 1186
rect 5293 1133 5307 1147
rect 5193 1053 5207 1067
rect 5673 1692 5687 1706
rect 5893 1912 5907 1926
rect 5873 1793 5887 1807
rect 5833 1753 5847 1767
rect 5813 1734 5827 1748
rect 5753 1692 5767 1706
rect 5793 1692 5807 1706
rect 5833 1673 5847 1687
rect 5733 1553 5747 1567
rect 5673 1513 5687 1527
rect 5593 1293 5607 1307
rect 5653 1293 5667 1307
rect 5473 1172 5487 1186
rect 5533 1172 5547 1186
rect 5573 1173 5587 1187
rect 5433 1113 5447 1127
rect 5373 1033 5387 1047
rect 5293 973 5307 987
rect 5253 953 5267 967
rect 5213 933 5227 947
rect 5173 914 5187 928
rect 5053 853 5067 867
rect 5113 853 5127 867
rect 5133 833 5147 847
rect 5113 753 5127 767
rect 5153 793 5167 807
rect 5133 733 5147 747
rect 5333 913 5347 927
rect 5273 833 5287 847
rect 5253 713 5267 727
rect 5313 713 5327 727
rect 5033 673 5047 687
rect 5193 653 5207 667
rect 5193 633 5207 647
rect 5173 593 5187 607
rect 5093 573 5107 587
rect 4993 493 5007 507
rect 4933 433 4947 447
rect 4973 433 4987 447
rect 4753 413 4767 427
rect 4813 394 4827 408
rect 5053 394 5067 408
rect 5273 652 5287 666
rect 5413 993 5427 1007
rect 5573 1073 5587 1087
rect 5433 913 5447 927
rect 5473 913 5487 927
rect 5653 1272 5667 1286
rect 5733 1434 5747 1448
rect 5853 1653 5867 1667
rect 5853 1593 5867 1607
rect 5873 1434 5887 1448
rect 5833 1373 5847 1387
rect 5713 1273 5727 1287
rect 5813 1273 5827 1287
rect 5673 1213 5687 1227
rect 5713 1172 5727 1186
rect 5773 1172 5787 1186
rect 5813 1172 5827 1186
rect 5893 1373 5907 1387
rect 5853 1333 5867 1347
rect 5893 1214 5907 1228
rect 5913 1153 5927 1167
rect 5833 1113 5847 1127
rect 5733 1093 5747 1107
rect 5593 933 5607 947
rect 5713 933 5727 947
rect 5613 914 5627 928
rect 5373 853 5387 867
rect 5573 853 5587 867
rect 5373 753 5387 767
rect 5333 693 5347 707
rect 5413 694 5427 708
rect 5353 652 5367 666
rect 5453 653 5467 667
rect 5433 633 5447 647
rect 5313 593 5327 607
rect 5393 593 5407 607
rect 5233 573 5247 587
rect 5353 513 5367 527
rect 5453 513 5467 527
rect 4533 352 4547 366
rect 4613 353 4627 367
rect 4673 352 4687 366
rect 4933 352 4947 366
rect 4973 353 4987 367
rect 5033 353 5047 367
rect 5073 352 5087 366
rect 5173 353 5187 367
rect 5233 352 5247 366
rect 5113 333 5127 347
rect 5253 333 5267 347
rect 4473 313 4487 327
rect 4453 193 4467 207
rect 4433 174 4447 188
rect 4713 313 4727 327
rect 5033 313 5047 327
rect 5093 313 5107 327
rect 4553 253 4567 267
rect 4513 213 4527 227
rect 4453 132 4467 146
rect 4493 132 4507 146
rect 5033 233 5047 247
rect 4593 174 4607 188
rect 4753 173 4767 187
rect 4833 174 4847 188
rect 4873 173 4887 187
rect 4973 174 4987 188
rect 4533 133 4547 147
rect 4513 113 4527 127
rect 4413 93 4427 107
rect 4573 113 4587 127
rect 4653 132 4667 146
rect 4713 132 4727 146
rect 4753 132 4767 146
rect 4953 132 4967 146
rect 5453 413 5467 427
rect 5533 652 5547 666
rect 5633 872 5647 886
rect 5693 872 5707 886
rect 5653 713 5667 727
rect 5493 413 5507 427
rect 5393 394 5407 408
rect 5593 653 5607 667
rect 5613 394 5627 408
rect 5813 914 5827 928
rect 5773 773 5787 787
rect 5773 713 5787 727
rect 6113 2313 6127 2327
rect 6073 2293 6087 2307
rect 6013 2254 6027 2268
rect 6233 2432 6247 2446
rect 6353 2474 6367 2488
rect 6413 2473 6427 2487
rect 6293 2432 6307 2446
rect 6373 2413 6387 2427
rect 6393 2313 6407 2327
rect 6253 2254 6267 2268
rect 6313 2254 6327 2268
rect 6353 2254 6367 2268
rect 6413 2273 6427 2287
rect 6013 2213 6027 2227
rect 6053 2212 6067 2226
rect 5973 2133 5987 2147
rect 6033 2013 6047 2027
rect 6193 2212 6207 2226
rect 6093 2073 6107 2087
rect 6273 2193 6287 2207
rect 6413 2212 6427 2226
rect 6373 2193 6387 2207
rect 6313 2133 6327 2147
rect 6373 2133 6387 2147
rect 6273 2073 6287 2087
rect 6133 2033 6147 2047
rect 6233 2033 6247 2047
rect 6053 1993 6067 2007
rect 5953 1953 5967 1967
rect 6013 1954 6027 1968
rect 6373 2013 6387 2027
rect 6433 2013 6447 2027
rect 6153 1993 6167 2007
rect 5993 1912 6007 1926
rect 5953 1873 5967 1887
rect 6233 1912 6247 1926
rect 6353 1912 6367 1926
rect 6133 1773 6147 1787
rect 6313 1773 6327 1787
rect 5973 1633 5987 1647
rect 6113 1693 6127 1707
rect 6053 1573 6067 1587
rect 6073 1513 6087 1527
rect 6193 1734 6207 1748
rect 6253 1733 6267 1747
rect 6353 1734 6367 1748
rect 6173 1692 6187 1706
rect 6213 1692 6227 1706
rect 6253 1692 6267 1706
rect 6293 1692 6307 1706
rect 6193 1653 6207 1667
rect 6033 1473 6047 1487
rect 5993 1434 6007 1448
rect 6173 1473 6187 1487
rect 6333 1434 6347 1448
rect 6393 1434 6407 1448
rect 6253 1392 6267 1406
rect 6373 1392 6387 1406
rect 6193 1373 6207 1387
rect 6073 1293 6087 1307
rect 6173 1293 6187 1307
rect 6033 1253 6047 1267
rect 5973 1233 5987 1247
rect 6013 1233 6027 1247
rect 6113 1253 6127 1267
rect 6073 1214 6087 1228
rect 5973 1172 5987 1186
rect 6013 1172 6027 1186
rect 6053 1172 6067 1186
rect 5953 1113 5967 1127
rect 5933 1093 5947 1107
rect 5953 1053 5967 1067
rect 5873 914 5887 928
rect 5913 914 5927 928
rect 6013 1013 6027 1027
rect 5973 933 5987 947
rect 5953 872 5967 886
rect 5893 773 5907 787
rect 5833 713 5847 727
rect 6173 1214 6187 1228
rect 6313 1273 6327 1287
rect 6233 1213 6247 1227
rect 6353 1214 6367 1228
rect 6193 1153 6207 1167
rect 6173 973 6187 987
rect 6053 914 6067 928
rect 6113 914 6127 928
rect 6073 872 6087 886
rect 6033 833 6047 847
rect 6053 694 6067 708
rect 6113 873 6127 887
rect 5753 652 5767 666
rect 5813 653 5827 667
rect 6173 933 6187 947
rect 6253 1192 6267 1206
rect 6393 1193 6407 1207
rect 6333 1172 6347 1186
rect 6253 1153 6267 1167
rect 6293 1113 6307 1127
rect 6193 872 6207 886
rect 6233 872 6247 886
rect 6173 694 6187 708
rect 5873 573 5887 587
rect 6073 652 6087 666
rect 6133 652 6147 666
rect 6213 652 6227 666
rect 6033 593 6047 607
rect 5913 553 5927 567
rect 6073 553 6087 567
rect 6033 473 6047 487
rect 5713 433 5727 447
rect 5753 433 5767 447
rect 5713 394 5727 408
rect 5793 393 5807 407
rect 5833 394 5847 408
rect 5873 394 5887 408
rect 5953 394 5967 408
rect 5993 394 6007 408
rect 6033 394 6047 408
rect 5733 352 5747 366
rect 5793 333 5807 347
rect 5573 273 5587 287
rect 5153 174 5167 188
rect 5213 174 5227 188
rect 5253 174 5267 188
rect 5353 174 5367 188
rect 5393 174 5407 188
rect 4993 113 5007 127
rect 5033 113 5047 127
rect 5113 132 5127 146
rect 5813 174 5827 188
rect 5893 333 5907 347
rect 6013 352 6027 366
rect 6273 693 6287 707
rect 6273 653 6287 667
rect 6233 473 6247 487
rect 6273 413 6287 427
rect 6373 914 6387 928
rect 6333 833 6347 847
rect 6313 713 6327 727
rect 6353 652 6367 666
rect 6093 353 6107 367
rect 6193 352 6207 366
rect 6093 313 6107 327
rect 6153 313 6167 327
rect 6073 293 6087 307
rect 5873 273 5887 287
rect 5953 273 5967 287
rect 5913 174 5927 188
rect 5153 113 5167 127
rect 4613 93 4627 107
rect 4873 93 4887 107
rect 4953 93 4967 107
rect 5073 93 5087 107
rect 5233 132 5247 146
rect 5333 132 5347 146
rect 5473 132 5487 146
rect 5573 132 5587 146
rect 5633 133 5647 147
rect 5513 113 5527 127
rect 5693 132 5707 146
rect 5852 133 5866 147
rect 5873 133 5887 147
rect 6153 174 6167 188
rect 6193 174 6207 188
rect 6373 413 6387 427
rect 6333 313 6347 327
rect 6293 293 6307 307
rect 6433 1172 6447 1186
rect 6393 313 6407 327
rect 6293 253 6307 267
rect 6373 253 6387 267
rect 6233 173 6247 187
rect 6393 213 6407 227
rect 5933 132 5947 146
rect 5633 113 5647 127
rect 6033 132 6047 146
rect 6073 132 6087 146
rect 6193 133 6207 147
rect 6273 132 6287 146
rect 5973 113 5987 127
rect 4533 73 4547 87
rect 4593 73 4607 87
rect 4633 73 4647 87
rect 4933 73 4947 87
rect 4973 73 4987 87
rect 5053 73 5067 87
rect 5093 73 5107 87
rect 5193 73 5207 87
rect 4133 13 4147 27
rect 4333 13 4347 27
<< metal3 >>
rect 2107 6256 2133 6264
rect 1527 6236 2413 6244
rect 2487 6236 2753 6244
rect 2947 6236 3904 6244
rect 1287 6216 1413 6224
rect 2007 6216 2353 6224
rect 2787 6216 3193 6224
rect 3427 6216 3713 6224
rect 3896 6224 3904 6236
rect 5707 6236 5753 6244
rect 3896 6216 4493 6224
rect 4987 6216 5613 6224
rect 607 6196 673 6204
rect 687 6196 1033 6204
rect 1687 6196 1973 6204
rect 2047 6196 2393 6204
rect 2467 6196 2753 6204
rect 2967 6196 3053 6204
rect 467 6176 513 6184
rect 1427 6176 1573 6184
rect 1587 6176 1993 6184
rect 2787 6176 3213 6184
rect 3287 6176 3393 6184
rect 3527 6176 4033 6184
rect 4327 6176 4673 6184
rect 4727 6176 5193 6184
rect 5207 6176 5473 6184
rect 5627 6176 5753 6184
rect 167 6156 253 6164
rect 267 6156 373 6164
rect 447 6156 493 6164
rect 507 6156 693 6164
rect 787 6156 913 6164
rect 1047 6156 1393 6164
rect 1507 6156 1733 6164
rect 2027 6156 2133 6164
rect 2227 6156 2613 6164
rect 2627 6156 2753 6164
rect 3107 6156 3173 6164
rect 3247 6156 3473 6164
rect 3727 6156 4133 6164
rect 4147 6156 4193 6164
rect 4287 6156 4693 6164
rect 4747 6156 4873 6164
rect 4887 6156 5413 6164
rect 6127 6156 6213 6164
rect 367 6136 413 6144
rect 2367 6136 2733 6144
rect 3627 6136 3804 6144
rect 3796 6128 3804 6136
rect 4427 6136 4533 6144
rect 5527 6136 5653 6144
rect 5667 6136 5793 6144
rect 5807 6136 6093 6144
rect 127 6117 193 6125
rect 487 6117 533 6125
rect 847 6117 873 6125
rect 927 6116 1024 6124
rect 296 6084 304 6114
rect 636 6087 644 6114
rect 736 6104 744 6114
rect 736 6096 993 6104
rect 1016 6104 1024 6116
rect 1087 6116 1173 6124
rect 1327 6116 1433 6124
rect 1627 6117 1653 6125
rect 1807 6117 1833 6125
rect 1876 6104 1884 6114
rect 1947 6116 2004 6124
rect 1016 6096 1524 6104
rect 247 6076 304 6084
rect 387 6076 413 6084
rect 527 6076 573 6084
rect 636 6076 653 6087
rect 640 6073 653 6076
rect 707 6076 753 6084
rect 776 6076 893 6084
rect 107 6056 493 6064
rect 647 6056 733 6064
rect 776 6064 784 6076
rect 907 6076 1024 6084
rect 747 6056 784 6064
rect 1016 6064 1024 6076
rect 1347 6075 1493 6083
rect 1516 6084 1524 6096
rect 1776 6096 1884 6104
rect 1996 6104 2004 6116
rect 2267 6117 2313 6125
rect 2547 6116 2713 6124
rect 2036 6104 2044 6114
rect 1996 6096 2044 6104
rect 2716 6104 2724 6114
rect 2807 6117 2833 6125
rect 3016 6104 3024 6114
rect 2716 6096 2784 6104
rect 1516 6076 1553 6084
rect 1687 6075 1713 6083
rect 1776 6084 1784 6096
rect 1767 6076 1784 6084
rect 1807 6076 1973 6084
rect 2167 6076 2233 6084
rect 2347 6076 2453 6084
rect 2776 6084 2784 6096
rect 2856 6096 3024 6104
rect 2856 6084 2864 6096
rect 2776 6076 2864 6084
rect 3016 6084 3024 6096
rect 3016 6076 3133 6084
rect 1016 6056 1053 6064
rect 1327 6056 1513 6064
rect 1667 6056 2473 6064
rect 2587 6056 2704 6064
rect 2696 6047 2704 6056
rect 2747 6056 2853 6064
rect 2907 6056 3093 6064
rect 3156 6064 3164 6114
rect 3267 6116 3293 6124
rect 3407 6117 3433 6125
rect 3487 6116 3573 6124
rect 3807 6117 3833 6125
rect 4027 6116 4053 6124
rect 3336 6084 3344 6114
rect 3576 6104 3584 6114
rect 4067 6116 4093 6124
rect 4227 6117 4373 6125
rect 4707 6116 4833 6124
rect 4847 6116 5004 6124
rect 3576 6096 3704 6104
rect 3287 6076 3344 6084
rect 3407 6076 3633 6084
rect 3696 6086 3704 6096
rect 4207 6096 4333 6104
rect 3747 6076 3853 6084
rect 4167 6076 4313 6084
rect 4447 6076 4533 6084
rect 4556 6067 4564 6113
rect 4596 6087 4604 6114
rect 4996 6104 5004 6116
rect 5027 6116 5093 6124
rect 5107 6117 5153 6125
rect 5316 6104 5324 6114
rect 5887 6116 6053 6124
rect 6147 6117 6173 6125
rect 6267 6117 6293 6125
rect 4996 6096 5304 6104
rect 5316 6096 5344 6104
rect 4596 6076 4613 6087
rect 4600 6073 4613 6076
rect 5296 6086 5304 6096
rect 4727 6076 4853 6084
rect 4867 6076 4993 6084
rect 5047 6076 5133 6084
rect 5336 6084 5344 6096
rect 5336 6076 5373 6084
rect 5427 6076 5453 6084
rect 5507 6076 5573 6084
rect 5587 6075 5633 6083
rect 5647 6076 5773 6084
rect 6087 6076 6113 6084
rect 6156 6080 6193 6084
rect 6153 6076 6193 6080
rect 6153 6067 6167 6076
rect 3156 6056 3313 6064
rect 3327 6056 3384 6064
rect 247 6036 313 6044
rect 1107 6036 1693 6044
rect 1747 6036 1893 6044
rect 1907 6036 2013 6044
rect 2067 6036 2253 6044
rect 2307 6036 2392 6044
rect 2427 6036 2573 6044
rect 2707 6036 2993 6044
rect 3007 6036 3093 6044
rect 3376 6044 3384 6056
rect 3607 6056 3893 6064
rect 4647 6056 4673 6064
rect 5656 6056 5733 6064
rect 3376 6036 3604 6044
rect 807 6016 933 6024
rect 947 6016 2273 6024
rect 2287 6016 2353 6024
rect 2627 6016 3313 6024
rect 3387 6016 3513 6024
rect 3596 6024 3604 6036
rect 3647 6036 3733 6044
rect 3807 6036 3873 6044
rect 4047 6036 4212 6044
rect 4247 6036 4533 6044
rect 4747 6036 4933 6044
rect 5107 6036 5153 6044
rect 5656 6044 5664 6056
rect 6307 6056 6373 6064
rect 5387 6036 5664 6044
rect 5747 6036 6033 6044
rect 6047 6036 6113 6044
rect 3596 6016 3864 6024
rect 147 5996 273 6004
rect 287 5996 353 6004
rect 507 5996 713 6004
rect 867 5996 933 6004
rect 947 5996 1293 6004
rect 1347 5996 1433 6004
rect 1707 5996 2213 6004
rect 2547 5996 2633 6004
rect 2687 5996 2953 6004
rect 3347 5996 3553 6004
rect 3856 6004 3864 6016
rect 4627 6016 5073 6024
rect 5087 6016 5173 6024
rect 5407 6016 5493 6024
rect 5967 6016 6013 6024
rect 6027 6016 6073 6024
rect 3856 5996 4233 6004
rect 4587 5996 5093 6004
rect 5396 6004 5404 6013
rect 5107 5996 5404 6004
rect 5447 5996 5893 6004
rect 467 5976 613 5984
rect 687 5976 753 5984
rect 807 5976 833 5984
rect 1467 5976 2104 5984
rect 367 5956 533 5964
rect 667 5956 1033 5964
rect 1047 5956 1193 5964
rect 1207 5956 1233 5964
rect 1687 5956 1753 5964
rect 2096 5964 2104 5976
rect 2267 5976 3233 5984
rect 3367 5976 3552 5984
rect 3587 5976 3633 5984
rect 3827 5976 3853 5984
rect 4287 5976 4373 5984
rect 4627 5976 4813 5984
rect 5147 5984 5160 5987
rect 5147 5973 5164 5984
rect 6227 5976 6413 5984
rect 2096 5956 2273 5964
rect 2487 5956 2673 5964
rect 2787 5956 2933 5964
rect 3267 5956 3913 5964
rect 4007 5956 4193 5964
rect 4267 5956 4553 5964
rect 4567 5956 5033 5964
rect 5047 5956 5113 5964
rect 5156 5964 5164 5973
rect 5156 5956 5873 5964
rect 67 5936 233 5944
rect 287 5936 473 5944
rect 687 5936 813 5944
rect 1447 5936 1593 5944
rect 1667 5936 2153 5944
rect 2807 5936 2893 5944
rect 2967 5936 3113 5944
rect 3467 5936 3713 5944
rect 4327 5936 4453 5944
rect 4547 5936 4653 5944
rect 4907 5936 4953 5944
rect 5347 5936 5413 5944
rect 5507 5936 5593 5944
rect 6336 5936 6393 5944
rect 416 5916 553 5924
rect 127 5896 144 5904
rect 136 5864 144 5896
rect 167 5896 393 5904
rect 136 5856 173 5864
rect 256 5866 264 5896
rect 307 5856 333 5864
rect 416 5866 424 5916
rect 627 5916 1333 5924
rect 1527 5916 1564 5924
rect 487 5896 524 5904
rect 516 5867 524 5896
rect 576 5884 584 5894
rect 927 5897 993 5905
rect 1087 5897 1133 5905
rect 1187 5896 1324 5904
rect 733 5884 747 5893
rect 576 5880 747 5884
rect 576 5876 744 5880
rect 796 5864 804 5893
rect 1316 5866 1324 5896
rect 1447 5897 1493 5905
rect 1556 5904 1564 5916
rect 2347 5916 2413 5924
rect 3327 5924 3340 5927
rect 3327 5914 3344 5924
rect 3320 5913 3344 5914
rect 3987 5916 4213 5924
rect 4380 5924 4392 5927
rect 4376 5913 4392 5924
rect 4441 5916 4573 5924
rect 6336 5924 6344 5936
rect 6087 5916 6344 5924
rect 1556 5896 1713 5904
rect 1727 5896 1873 5904
rect 2067 5896 2184 5904
rect 1876 5884 1884 5894
rect 2016 5884 2024 5894
rect 1876 5876 2024 5884
rect 567 5856 584 5864
rect 796 5856 833 5864
rect 107 5836 153 5844
rect 167 5836 193 5844
rect 576 5844 584 5856
rect 1247 5855 1273 5863
rect 2176 5866 2184 5896
rect 2147 5856 2173 5864
rect 2196 5847 2204 5894
rect 2287 5896 2313 5904
rect 2567 5897 2593 5905
rect 2707 5897 2733 5905
rect 2316 5884 2324 5894
rect 2236 5876 2324 5884
rect 2896 5884 2904 5894
rect 2967 5896 2993 5904
rect 3047 5896 3173 5904
rect 3196 5896 3292 5904
rect 3196 5884 3204 5896
rect 2896 5876 2944 5884
rect 2236 5864 2244 5876
rect 2227 5856 2244 5864
rect 2267 5855 2293 5863
rect 2936 5864 2944 5876
rect 3156 5876 3204 5884
rect 3156 5866 3164 5876
rect 3336 5866 3344 5913
rect 3527 5896 3624 5904
rect 2936 5856 3013 5864
rect 3067 5856 3153 5864
rect 3476 5864 3484 5894
rect 3616 5866 3624 5896
rect 3656 5866 3664 5913
rect 3676 5867 3684 5894
rect 3387 5856 3484 5864
rect 3507 5855 3533 5863
rect 3676 5856 3693 5867
rect 3680 5853 3693 5856
rect 3816 5864 3824 5894
rect 4036 5896 4133 5904
rect 3916 5864 3924 5893
rect 3816 5856 3864 5864
rect 3916 5856 3933 5864
rect 576 5836 753 5844
rect 887 5836 984 5844
rect 976 5827 984 5836
rect 1027 5833 1033 5847
rect 1487 5836 1613 5844
rect 2707 5836 2733 5844
rect 3627 5836 3653 5844
rect 3856 5844 3864 5856
rect 4036 5864 4044 5896
rect 4247 5904 4260 5907
rect 4247 5893 4264 5904
rect 4176 5867 4184 5893
rect 4027 5856 4044 5864
rect 4067 5855 4113 5863
rect 4256 5866 4264 5893
rect 4296 5896 4333 5904
rect 4296 5866 4304 5896
rect 4376 5867 4384 5913
rect 4456 5867 4464 5894
rect 4527 5896 4613 5904
rect 4807 5896 4853 5904
rect 4907 5896 4993 5904
rect 5016 5896 5073 5904
rect 4456 5856 4473 5867
rect 4460 5853 4473 5856
rect 5016 5866 5024 5896
rect 5387 5896 5404 5904
rect 5196 5884 5204 5894
rect 5196 5876 5253 5884
rect 5396 5867 5404 5896
rect 5547 5897 5613 5905
rect 5807 5897 5833 5905
rect 6167 5896 6313 5904
rect 6367 5897 6433 5905
rect 4667 5855 4713 5863
rect 4767 5855 4813 5863
rect 4927 5855 4953 5863
rect 5987 5856 6053 5864
rect 3856 5836 3913 5844
rect 3927 5836 4033 5844
rect 4507 5836 4593 5844
rect 5367 5836 5473 5844
rect 6127 5836 6193 5844
rect 987 5816 1073 5824
rect 1087 5816 1653 5824
rect 1787 5816 1853 5824
rect 1867 5816 1913 5824
rect 1927 5816 1953 5824
rect 1967 5816 1993 5824
rect 2047 5816 2173 5824
rect 2247 5816 2453 5824
rect 2687 5816 2793 5824
rect 3107 5816 3333 5824
rect 3467 5816 3793 5824
rect 3967 5816 3993 5824
rect 4487 5816 4633 5824
rect 5127 5816 5313 5824
rect 6027 5816 6093 5824
rect 67 5796 133 5804
rect 147 5796 353 5804
rect 927 5796 1033 5804
rect 1047 5796 1153 5804
rect 1507 5796 1573 5804
rect 1587 5796 1933 5804
rect 2476 5796 2753 5804
rect 2476 5784 2484 5796
rect 2927 5796 3113 5804
rect 3127 5796 3193 5804
rect 3447 5796 3733 5804
rect 3887 5796 4253 5804
rect 4267 5796 4393 5804
rect 5267 5796 5533 5804
rect 6147 5796 6233 5804
rect 2407 5776 2484 5784
rect 3196 5784 3204 5793
rect 3196 5776 3693 5784
rect 4447 5776 4493 5784
rect 5227 5776 5633 5784
rect 5647 5776 5753 5784
rect 1827 5756 1893 5764
rect 1907 5756 2033 5764
rect 2207 5756 2333 5764
rect 2347 5756 2733 5764
rect 3287 5756 3433 5764
rect 3487 5756 3972 5764
rect 4007 5756 4333 5764
rect 5127 5756 5693 5764
rect 5707 5756 5933 5764
rect 2147 5736 2253 5744
rect 3727 5736 4013 5744
rect 4407 5736 4553 5744
rect 4947 5736 5793 5744
rect 5807 5736 5973 5744
rect 1367 5716 1513 5724
rect 2127 5716 2313 5724
rect 2447 5716 2713 5724
rect 2867 5716 3153 5724
rect 3167 5716 3453 5724
rect 3607 5716 3833 5724
rect 4167 5716 4193 5724
rect 4207 5716 4513 5724
rect 5187 5716 5593 5724
rect 707 5696 1544 5704
rect 1067 5676 1413 5684
rect 1536 5684 1544 5696
rect 1687 5696 1853 5704
rect 1867 5696 1993 5704
rect 2107 5696 2173 5704
rect 2467 5696 2533 5704
rect 2547 5696 2653 5704
rect 3207 5696 3353 5704
rect 3907 5696 4353 5704
rect 4636 5696 4873 5704
rect 1536 5676 2433 5684
rect 3147 5676 3412 5684
rect 3447 5676 3533 5684
rect 4636 5684 4644 5696
rect 5527 5696 5713 5704
rect 3587 5676 4644 5684
rect 987 5656 1093 5664
rect 1107 5656 1433 5664
rect 1507 5656 1653 5664
rect 1807 5656 2424 5664
rect 787 5636 933 5644
rect 1207 5636 1393 5644
rect 1687 5636 1753 5644
rect 2416 5644 2424 5656
rect 2447 5656 3013 5664
rect 3027 5656 3333 5664
rect 3567 5656 3633 5664
rect 3787 5656 3933 5664
rect 4027 5656 4173 5664
rect 4667 5656 5113 5664
rect 5347 5656 5433 5664
rect 6267 5656 6333 5664
rect 2416 5636 3173 5644
rect 3387 5636 3913 5644
rect 4387 5636 4473 5644
rect 4547 5636 4673 5644
rect 4727 5636 4873 5644
rect 5147 5636 5193 5644
rect 5327 5636 5713 5644
rect 5827 5636 5973 5644
rect 6087 5636 6213 5644
rect 6227 5636 6373 5644
rect 207 5616 393 5624
rect 467 5616 493 5624
rect 1927 5616 2133 5624
rect 3647 5616 3973 5624
rect 3987 5616 4213 5624
rect 4367 5616 4704 5624
rect 127 5596 193 5604
rect 247 5596 313 5604
rect 327 5597 353 5605
rect 376 5596 513 5604
rect 376 5584 384 5596
rect 527 5596 613 5604
rect 627 5597 653 5605
rect 827 5596 933 5604
rect 947 5596 993 5604
rect 1036 5596 1133 5604
rect 1036 5584 1044 5596
rect 1147 5597 1193 5605
rect 1287 5597 1332 5605
rect 1367 5596 1424 5604
rect 1416 5584 1424 5596
rect 1487 5597 1533 5605
rect 1787 5597 1813 5605
rect 2267 5596 2353 5604
rect 2587 5597 2933 5605
rect 3136 5596 3193 5604
rect 96 5576 384 5584
rect 1016 5576 1044 5584
rect 1116 5576 1424 5584
rect 96 5566 104 5576
rect 187 5555 213 5563
rect 347 5555 373 5563
rect 467 5555 533 5563
rect 607 5555 673 5563
rect 727 5556 773 5564
rect 1016 5564 1024 5576
rect 847 5556 1024 5564
rect 1116 5547 1124 5576
rect 1416 5566 1424 5576
rect 1347 5556 1373 5564
rect 1436 5564 1444 5594
rect 1436 5556 1513 5564
rect 267 5536 293 5544
rect 967 5536 1113 5544
rect 1716 5544 1724 5594
rect 2096 5564 2104 5594
rect 2216 5567 2224 5594
rect 2476 5584 2484 5594
rect 2327 5576 2484 5584
rect 2067 5556 2104 5564
rect 2207 5556 2224 5567
rect 2207 5553 2220 5556
rect 2307 5556 2493 5564
rect 2516 5564 2524 5594
rect 3136 5566 3144 5596
rect 3347 5597 3413 5605
rect 3507 5597 3533 5605
rect 3887 5597 3933 5605
rect 4307 5596 4344 5604
rect 3296 5584 3304 5594
rect 3296 5576 3344 5584
rect 2516 5556 2673 5564
rect 2727 5555 2913 5563
rect 3007 5556 3093 5564
rect 3227 5555 3313 5563
rect 3336 5564 3344 5576
rect 3367 5576 3653 5584
rect 3436 5566 3444 5576
rect 3336 5556 3393 5564
rect 3607 5556 3633 5564
rect 3967 5556 4013 5564
rect 4076 5547 4084 5594
rect 4336 5584 4344 5596
rect 4367 5597 4393 5605
rect 4507 5597 4533 5605
rect 4436 5584 4444 5594
rect 4167 5576 4444 5584
rect 4556 5566 4564 5616
rect 4527 5556 4553 5564
rect 1687 5536 1724 5544
rect 2367 5536 2453 5544
rect 2547 5536 2633 5544
rect 4187 5536 4353 5544
rect 4576 5546 4584 5594
rect 4656 5564 4664 5593
rect 4696 5566 4704 5616
rect 4927 5616 5173 5624
rect 5367 5616 5413 5624
rect 4727 5597 4773 5605
rect 5007 5596 5093 5604
rect 5447 5597 5493 5605
rect 5627 5597 5653 5605
rect 4607 5556 4664 5564
rect 4836 5564 4844 5594
rect 4900 5584 4913 5587
rect 4896 5573 4913 5584
rect 4747 5556 4844 5564
rect 4896 5564 4904 5573
rect 4867 5556 4904 5564
rect 4927 5555 4973 5563
rect 5167 5556 5213 5564
rect 5227 5556 5233 5564
rect 5507 5556 5553 5564
rect 5576 5564 5584 5594
rect 5707 5596 5744 5604
rect 5576 5556 5633 5564
rect 5736 5566 5744 5596
rect 5767 5597 5853 5605
rect 5936 5567 5944 5594
rect 5847 5555 5873 5563
rect 5936 5556 5953 5567
rect 5940 5553 5953 5556
rect 6036 5564 6044 5594
rect 6216 5596 6253 5604
rect 6156 5567 6164 5593
rect 6007 5556 6044 5564
rect 6216 5547 6224 5596
rect 6316 5567 6324 5594
rect 6307 5556 6324 5567
rect 6356 5567 6364 5594
rect 6356 5556 6373 5567
rect 6307 5553 6320 5556
rect 6360 5553 6373 5556
rect 4576 5545 4600 5546
rect 4576 5536 4593 5545
rect 4580 5533 4593 5536
rect 887 5516 933 5524
rect 1087 5516 1173 5524
rect 1187 5516 1233 5524
rect 1807 5516 1873 5524
rect 2047 5516 2233 5524
rect 2536 5524 2544 5533
rect 5987 5536 6013 5544
rect 2387 5516 2544 5524
rect 2687 5516 4153 5524
rect 4427 5516 4493 5524
rect 4887 5516 5293 5524
rect 5307 5516 5513 5524
rect 5567 5516 5593 5524
rect 5607 5516 5913 5524
rect 6067 5516 6133 5524
rect 6287 5516 6333 5524
rect 227 5496 333 5504
rect 356 5496 493 5504
rect 356 5484 364 5496
rect 1667 5496 1753 5504
rect 1767 5496 1873 5504
rect 2127 5496 2313 5504
rect 3227 5496 3553 5504
rect 3567 5496 3873 5504
rect 4107 5496 4253 5504
rect 4567 5496 4633 5504
rect 5467 5496 5813 5504
rect 5967 5496 6153 5504
rect 6167 5496 6373 5504
rect 307 5476 364 5484
rect 547 5476 693 5484
rect 1067 5476 1253 5484
rect 2187 5476 2233 5484
rect 2427 5476 2513 5484
rect 2907 5476 3773 5484
rect 4707 5476 4933 5484
rect 6047 5476 6112 5484
rect 6147 5476 6193 5484
rect 6247 5476 6353 5484
rect 1547 5456 1613 5464
rect 1627 5456 1973 5464
rect 1987 5456 2073 5464
rect 2207 5456 2473 5464
rect 2487 5456 4313 5464
rect 5687 5456 5993 5464
rect 627 5436 773 5444
rect 1027 5436 1093 5444
rect 2307 5436 2433 5444
rect 2687 5436 3493 5444
rect 3827 5436 3993 5444
rect 5367 5436 5393 5444
rect 5787 5436 5893 5444
rect 5907 5436 6233 5444
rect 6247 5436 6293 5444
rect 167 5416 373 5424
rect 427 5416 593 5424
rect 1127 5416 1204 5424
rect 1196 5404 1204 5416
rect 1487 5416 1513 5424
rect 1527 5416 1693 5424
rect 1847 5416 1913 5424
rect 1927 5416 2133 5424
rect 2467 5416 2573 5424
rect 3107 5416 3173 5424
rect 3407 5416 3813 5424
rect 4027 5416 4233 5424
rect 4427 5416 4473 5424
rect 5267 5416 5673 5424
rect 1196 5396 1293 5404
rect 2967 5396 3313 5404
rect 5327 5396 5353 5404
rect 5427 5396 5473 5404
rect 6207 5396 6253 5404
rect 167 5377 213 5385
rect 76 5347 84 5374
rect 287 5376 313 5384
rect 427 5377 453 5385
rect 476 5376 493 5384
rect 476 5364 484 5376
rect 67 5336 84 5347
rect 396 5356 484 5364
rect 396 5346 404 5356
rect 67 5333 80 5336
rect 107 5336 233 5344
rect 536 5344 544 5374
rect 627 5376 653 5384
rect 536 5336 573 5344
rect 676 5346 684 5393
rect 767 5376 813 5384
rect 867 5377 913 5385
rect 927 5376 1013 5384
rect 1187 5376 1333 5384
rect 1347 5377 1373 5385
rect 1396 5376 1413 5384
rect 1093 5364 1107 5373
rect 1093 5360 1124 5364
rect 1096 5356 1124 5360
rect 1116 5346 1124 5356
rect 1136 5327 1144 5374
rect 1396 5364 1404 5376
rect 1467 5376 1553 5384
rect 1567 5376 1593 5384
rect 1747 5376 1953 5384
rect 1316 5356 1404 5364
rect 1316 5346 1324 5356
rect 1227 5336 1273 5344
rect 1487 5335 1513 5343
rect 1676 5344 1684 5373
rect 1856 5346 1864 5376
rect 1967 5377 2013 5385
rect 2027 5376 2173 5384
rect 2387 5377 2433 5385
rect 2447 5376 2593 5384
rect 2867 5377 2913 5385
rect 3047 5377 3113 5385
rect 3367 5376 3513 5384
rect 3527 5376 3593 5384
rect 3647 5376 3773 5384
rect 3787 5377 3853 5385
rect 3947 5377 4133 5385
rect 4347 5377 4373 5385
rect 4436 5376 4513 5384
rect 2773 5364 2787 5373
rect 2736 5360 2787 5364
rect 2736 5356 2784 5360
rect 1676 5336 1713 5344
rect 2207 5336 2413 5344
rect 2427 5336 2573 5344
rect 2736 5344 2744 5356
rect 2816 5346 2824 5373
rect 2876 5356 2953 5364
rect 2876 5346 2884 5356
rect 2727 5336 2744 5344
rect 2767 5335 2813 5343
rect 2927 5335 3013 5343
rect 3027 5336 3093 5344
rect 4436 5346 4444 5376
rect 4847 5376 4953 5384
rect 4967 5376 4984 5384
rect 4596 5347 4604 5373
rect 4976 5364 4984 5376
rect 5007 5377 5053 5385
rect 5067 5376 5133 5384
rect 5280 5384 5293 5387
rect 5276 5373 5293 5384
rect 5376 5376 5513 5384
rect 4976 5356 5124 5364
rect 3207 5336 3293 5344
rect 3347 5336 3493 5344
rect 3667 5336 3793 5344
rect 4327 5335 4393 5343
rect 4487 5335 4533 5343
rect 4727 5336 4753 5344
rect 5116 5344 5124 5356
rect 5276 5346 5284 5373
rect 5376 5346 5384 5376
rect 5627 5376 5653 5384
rect 5667 5376 5793 5384
rect 5847 5376 6093 5384
rect 5816 5356 5893 5364
rect 5116 5336 5233 5344
rect 5587 5336 5633 5344
rect 5816 5346 5824 5356
rect 6096 5364 6104 5374
rect 6167 5384 6180 5387
rect 6167 5373 6184 5384
rect 6287 5376 6373 5384
rect 5996 5356 6104 5364
rect 6176 5364 6184 5373
rect 6176 5356 6264 5364
rect 5647 5336 5693 5344
rect 5996 5344 6004 5356
rect 6256 5346 6264 5356
rect 5987 5336 6004 5344
rect 6016 5336 6073 5344
rect 807 5316 933 5324
rect 1007 5316 1073 5324
rect 2007 5316 2193 5324
rect 2247 5316 2293 5324
rect 2467 5316 2613 5324
rect 2627 5316 3313 5324
rect 996 5304 1004 5313
rect 4041 5316 4053 5324
rect 4547 5316 4673 5324
rect 4987 5316 5133 5324
rect 6016 5324 6024 5336
rect 6307 5335 6353 5343
rect 5947 5316 6024 5324
rect 6047 5316 6093 5324
rect 887 5296 1004 5304
rect 1107 5296 1193 5304
rect 1667 5296 1713 5304
rect 4147 5296 4813 5304
rect 4827 5296 4913 5304
rect 5207 5296 5253 5304
rect 5427 5296 5693 5304
rect 5767 5296 5833 5304
rect 6267 5296 6333 5304
rect 1167 5276 1313 5284
rect 1387 5276 1793 5284
rect 1947 5276 2172 5284
rect 2207 5276 2353 5284
rect 3067 5276 3153 5284
rect 3167 5276 3393 5284
rect 4307 5276 4333 5284
rect 607 5256 653 5264
rect 847 5256 1033 5264
rect 1967 5256 1993 5264
rect 2147 5256 2313 5264
rect 2447 5256 2513 5264
rect 3167 5256 3193 5264
rect 3236 5256 3393 5264
rect 1767 5236 1893 5244
rect 1987 5236 2353 5244
rect 2367 5236 2513 5244
rect 3236 5244 3244 5256
rect 3476 5256 3673 5264
rect 2587 5236 3244 5244
rect 3476 5244 3484 5256
rect 5027 5256 5153 5264
rect 5167 5256 5393 5264
rect 6096 5256 6193 5264
rect 3287 5236 3484 5244
rect 6096 5244 6104 5256
rect 6287 5256 6433 5264
rect 5867 5236 6104 5244
rect 6127 5236 6393 5244
rect 467 5216 593 5224
rect 607 5216 913 5224
rect 1287 5216 1433 5224
rect 2156 5216 2313 5224
rect 2156 5207 2164 5216
rect 2427 5216 3233 5224
rect 4967 5216 5053 5224
rect 5327 5216 5413 5224
rect 727 5196 773 5204
rect 787 5196 933 5204
rect 1587 5196 2033 5204
rect 2047 5196 2153 5204
rect 2347 5196 2393 5204
rect 2907 5196 3253 5204
rect 3407 5196 3504 5204
rect 667 5176 1704 5184
rect 307 5156 373 5164
rect 1696 5164 1704 5176
rect 1727 5176 2373 5184
rect 3496 5184 3504 5196
rect 3527 5196 3593 5204
rect 3607 5196 4673 5204
rect 3496 5176 3653 5184
rect 3667 5176 4413 5184
rect 5707 5176 6293 5184
rect 1696 5156 2193 5164
rect 2216 5156 2413 5164
rect 27 5136 413 5144
rect 687 5136 753 5144
rect 2216 5144 2224 5156
rect 2436 5156 2873 5164
rect 1607 5136 2224 5144
rect 2436 5144 2444 5156
rect 3127 5156 3413 5164
rect 3507 5156 3713 5164
rect 3867 5156 3933 5164
rect 4587 5156 5113 5164
rect 5127 5156 5313 5164
rect 2247 5136 2444 5144
rect 2507 5136 2993 5144
rect 4787 5136 4813 5144
rect 5487 5136 5593 5144
rect 6127 5136 6173 5144
rect 1087 5116 1133 5124
rect 1207 5116 1533 5124
rect 1547 5116 1712 5124
rect 1747 5116 1933 5124
rect 2667 5116 2753 5124
rect 3127 5116 3273 5124
rect 3807 5116 3893 5124
rect 3907 5116 4113 5124
rect 5367 5116 5733 5124
rect 6387 5116 6433 5124
rect 67 5096 233 5104
rect 247 5096 353 5104
rect 367 5096 404 5104
rect 127 5077 193 5085
rect 396 5084 404 5096
rect 767 5096 893 5104
rect 987 5096 1033 5104
rect 1047 5096 1233 5104
rect 1527 5096 2193 5104
rect 2327 5096 2493 5104
rect 3107 5096 3313 5104
rect 3433 5104 3447 5113
rect 3387 5100 3447 5104
rect 3387 5096 3444 5100
rect 3467 5096 3553 5104
rect 4707 5096 4793 5104
rect 4907 5096 5033 5104
rect 5447 5096 5493 5104
rect 5907 5096 6013 5104
rect 6193 5104 6207 5113
rect 6147 5100 6207 5104
rect 6147 5096 6204 5100
rect 396 5076 424 5084
rect 67 5035 133 5043
rect 207 5036 253 5044
rect 276 5044 284 5074
rect 416 5064 424 5076
rect 507 5076 513 5084
rect 527 5076 553 5084
rect 596 5076 673 5084
rect 416 5056 444 5064
rect 276 5036 313 5044
rect 436 5044 444 5056
rect 436 5036 533 5044
rect 596 5027 604 5076
rect 727 5076 853 5084
rect 907 5077 1213 5085
rect 1327 5077 1373 5085
rect 1427 5077 1453 5085
rect 1727 5077 1773 5085
rect 1827 5076 1853 5084
rect 1867 5077 1893 5085
rect 2227 5077 2253 5085
rect 2567 5077 2593 5085
rect 647 5036 693 5044
rect 1027 5035 1073 5043
rect 1167 5035 1213 5043
rect 1556 5044 1564 5073
rect 1527 5036 1564 5044
rect 1976 5044 1984 5073
rect 1967 5036 1984 5044
rect 2036 5027 2044 5074
rect 2076 5044 2084 5074
rect 2076 5036 2112 5044
rect 2147 5036 2193 5044
rect 2247 5036 2273 5044
rect 2676 5046 2684 5093
rect 2327 5036 2493 5044
rect 2816 5044 2824 5093
rect 2947 5076 3004 5084
rect 2996 5064 3004 5076
rect 3027 5076 3093 5084
rect 3187 5077 3233 5085
rect 3787 5077 3873 5085
rect 3887 5076 4073 5084
rect 2996 5060 3044 5064
rect 2996 5056 3047 5060
rect 3033 5047 3047 5056
rect 2816 5036 2953 5044
rect 3456 5047 3464 5074
rect 3507 5056 3544 5064
rect 3127 5036 3213 5044
rect 3327 5035 3393 5043
rect 3456 5036 3473 5047
rect 3460 5033 3473 5036
rect 3536 5044 3544 5056
rect 3536 5036 3573 5044
rect 3627 5036 3793 5044
rect 3887 5036 3953 5044
rect 4096 5044 4104 5093
rect 4267 5076 4373 5084
rect 4387 5076 4473 5084
rect 4527 5076 4613 5084
rect 4096 5036 4193 5044
rect 747 5016 873 5024
rect 887 5016 1013 5024
rect 1767 5016 1793 5024
rect 1807 5016 1913 5024
rect 2267 5016 2352 5024
rect 2387 5016 2533 5024
rect 3447 5016 3513 5024
rect 3827 5016 4053 5024
rect 4107 5016 4133 5024
rect 4216 5024 4224 5074
rect 4727 5077 4753 5085
rect 5127 5077 5153 5085
rect 5207 5076 5353 5084
rect 5076 5064 5084 5074
rect 5547 5077 5573 5085
rect 5596 5076 5673 5084
rect 4987 5056 5084 5064
rect 4247 5036 4493 5044
rect 4547 5036 4573 5044
rect 4707 5035 4913 5043
rect 5067 5036 5113 5044
rect 5187 5036 5253 5044
rect 5396 5044 5404 5073
rect 5396 5036 5473 5044
rect 5596 5044 5604 5076
rect 5687 5076 5793 5084
rect 6156 5076 6173 5084
rect 5527 5036 5604 5044
rect 5707 5036 5733 5044
rect 4216 5016 4784 5024
rect 4776 5007 4784 5016
rect 5287 5016 5313 5024
rect 5856 5024 5864 5073
rect 5896 5027 5904 5074
rect 5976 5027 5984 5074
rect 6156 5044 6164 5076
rect 6367 5077 6413 5085
rect 6273 5064 6287 5073
rect 6047 5036 6164 5044
rect 6176 5060 6287 5064
rect 6176 5056 6284 5060
rect 6176 5027 6184 5056
rect 6207 5035 6273 5043
rect 6316 5027 6324 5074
rect 5787 5016 5864 5024
rect 6307 5016 6324 5027
rect 6307 5013 6320 5016
rect 67 4996 393 5004
rect 587 4996 693 5004
rect 807 4996 973 5004
rect 2127 4996 2213 5004
rect 2427 4996 2593 5004
rect 2607 4996 2673 5004
rect 2687 4996 2773 5004
rect 2887 4996 3173 5004
rect 3727 4996 3873 5004
rect 4247 4996 4353 5004
rect 4427 4996 4493 5004
rect 4787 4996 4973 5004
rect 5227 4996 5373 5004
rect 5507 4996 5573 5004
rect 5587 4996 5653 5004
rect 6027 4996 6133 5004
rect 576 4984 584 4993
rect 447 4976 584 4984
rect 827 4976 933 4984
rect 1027 4976 1193 4984
rect 1347 4976 1453 4984
rect 1467 4976 1733 4984
rect 2407 4976 2473 4984
rect 2847 4976 2873 4984
rect 3167 4976 3253 4984
rect 3507 4976 3633 4984
rect 4027 4976 4113 4984
rect 4407 4976 4633 4984
rect 4647 4976 4713 4984
rect 4727 4976 4873 4984
rect 4896 4976 5333 4984
rect 207 4956 513 4964
rect 527 4956 693 4964
rect 1107 4956 1393 4964
rect 1707 4956 2093 4964
rect 2647 4956 2713 4964
rect 2827 4956 3133 4964
rect 3667 4956 3753 4964
rect 3907 4956 4033 4964
rect 4747 4956 4773 4964
rect 4896 4964 4904 4976
rect 5707 4976 6413 4984
rect 4847 4956 4904 4964
rect 5487 4956 5593 4964
rect 5927 4956 6073 4964
rect 6087 4956 6173 4964
rect 327 4936 413 4944
rect 2147 4936 2232 4944
rect 2267 4936 2393 4944
rect 2867 4936 3473 4944
rect 3847 4936 4213 4944
rect 4447 4936 4513 4944
rect 4596 4936 5013 4944
rect 267 4916 913 4924
rect 1267 4916 1293 4924
rect 1336 4916 1613 4924
rect 307 4896 373 4904
rect 467 4896 593 4904
rect 1336 4904 1344 4916
rect 2067 4916 2092 4924
rect 2856 4924 2864 4933
rect 2127 4916 2864 4924
rect 3007 4916 3353 4924
rect 3367 4916 3413 4924
rect 3467 4916 3652 4924
rect 3687 4916 3733 4924
rect 4596 4924 4604 4936
rect 5287 4936 5873 4944
rect 5887 4936 6293 4944
rect 4367 4916 4604 4924
rect 4887 4916 4953 4924
rect 5547 4916 5853 4924
rect 1047 4896 1344 4904
rect 1507 4896 1704 4904
rect 1696 4887 1704 4896
rect 1727 4896 2073 4904
rect 2207 4896 2333 4904
rect 2607 4896 2753 4904
rect 3607 4896 3693 4904
rect 4007 4896 4053 4904
rect 4167 4896 4213 4904
rect 4287 4896 4313 4904
rect 4387 4896 4693 4904
rect 5047 4896 5233 4904
rect 5367 4896 5413 4904
rect 5927 4896 6013 4904
rect 6447 4904 6460 4907
rect 6447 4893 6464 4904
rect 356 4876 393 4884
rect 67 4864 80 4867
rect 67 4853 84 4864
rect 107 4856 173 4864
rect 187 4857 253 4865
rect 307 4856 333 4864
rect 76 4826 84 4853
rect 356 4844 364 4876
rect 667 4876 753 4884
rect 796 4876 833 4884
rect 276 4836 364 4844
rect 376 4856 553 4864
rect 276 4826 284 4836
rect 127 4816 193 4824
rect 207 4815 233 4823
rect 376 4824 384 4856
rect 796 4864 804 4876
rect 1696 4886 1720 4887
rect 1696 4876 1713 4886
rect 1700 4873 1713 4876
rect 2107 4876 2313 4884
rect 2767 4876 2813 4884
rect 2927 4876 3644 4884
rect 576 4856 804 4864
rect 576 4826 584 4856
rect 907 4857 953 4865
rect 1107 4857 1173 4865
rect 1227 4857 1253 4865
rect 1347 4856 1393 4864
rect 1467 4857 1553 4865
rect 1567 4856 1673 4864
rect 1776 4856 1793 4864
rect 1616 4840 1744 4844
rect 1616 4836 1747 4840
rect 296 4816 384 4824
rect 296 4784 304 4816
rect 447 4816 573 4824
rect 727 4816 793 4824
rect 807 4816 893 4824
rect 1287 4815 1333 4823
rect 1387 4816 1453 4824
rect 1616 4824 1624 4836
rect 1733 4827 1747 4836
rect 1776 4827 1784 4856
rect 1807 4856 1893 4864
rect 1947 4856 2013 4864
rect 2036 4856 2073 4864
rect 2036 4844 2044 4856
rect 2100 4864 2113 4867
rect 1956 4836 2044 4844
rect 2096 4853 2113 4864
rect 1587 4816 1624 4824
rect 1647 4816 1693 4824
rect 1827 4816 1853 4824
rect 1956 4826 1964 4836
rect 2096 4826 2104 4853
rect 2376 4824 2384 4854
rect 2587 4857 2633 4865
rect 2327 4816 2384 4824
rect 2416 4824 2424 4853
rect 2407 4816 2424 4824
rect 2516 4824 2524 4854
rect 2747 4856 2933 4864
rect 2987 4856 3093 4864
rect 3247 4857 3273 4865
rect 3567 4856 3613 4864
rect 2516 4816 2613 4824
rect 2787 4816 3013 4824
rect 3176 4824 3184 4853
rect 3456 4827 3464 4854
rect 3167 4816 3184 4824
rect 3327 4816 3393 4824
rect 3456 4816 3472 4827
rect 3460 4813 3472 4816
rect 3507 4816 3533 4824
rect 3556 4824 3564 4854
rect 3636 4864 3644 4876
rect 3667 4876 3793 4884
rect 3807 4876 4264 4884
rect 3636 4856 3653 4864
rect 3760 4864 3773 4867
rect 3756 4853 3773 4864
rect 3887 4856 3913 4864
rect 3927 4856 3953 4864
rect 4007 4856 4073 4864
rect 4167 4857 4193 4865
rect 4256 4864 4264 4876
rect 4307 4876 4533 4884
rect 5956 4876 6033 4884
rect 4256 4856 4273 4864
rect 4667 4857 4733 4865
rect 5007 4857 5033 4865
rect 3756 4844 3764 4853
rect 3716 4836 3764 4844
rect 3556 4816 3633 4824
rect 3716 4824 3724 4836
rect 3687 4816 3724 4824
rect 3747 4815 3853 4823
rect 4087 4815 4133 4823
rect 4187 4816 4233 4824
rect 4436 4807 4444 4854
rect 4836 4836 4973 4844
rect 4587 4816 4653 4824
rect 947 4796 993 4804
rect 1227 4796 1552 4804
rect 187 4776 304 4784
rect 936 4784 944 4793
rect 1587 4796 2053 4804
rect 2147 4796 2233 4804
rect 2387 4796 2713 4804
rect 3167 4796 3273 4804
rect 3447 4796 3513 4804
rect 4027 4796 4373 4804
rect 4387 4796 4412 4804
rect 4836 4804 4844 4836
rect 4896 4826 4904 4836
rect 5396 4844 5404 4854
rect 5587 4856 5613 4864
rect 5627 4857 5653 4865
rect 5376 4836 5404 4844
rect 5147 4816 5193 4824
rect 5376 4824 5384 4836
rect 5267 4816 5384 4824
rect 5496 4824 5504 4853
rect 5776 4827 5784 4853
rect 5816 4827 5824 4854
rect 5427 4816 5504 4824
rect 5567 4816 5673 4824
rect 5816 4816 5833 4827
rect 5820 4813 5833 4816
rect 5896 4826 5904 4873
rect 5956 4807 5964 4876
rect 6287 4876 6333 4884
rect 6387 4876 6433 4884
rect 6016 4827 6024 4853
rect 6056 4807 6064 4854
rect 6196 4844 6204 4854
rect 6307 4864 6320 4867
rect 6307 4853 6324 4864
rect 6456 4864 6464 4893
rect 6436 4856 6464 4864
rect 6196 4836 6244 4844
rect 6087 4816 6213 4824
rect 4767 4796 4844 4804
rect 4867 4796 4993 4804
rect 5007 4796 5753 4804
rect 6236 4804 6244 4836
rect 6316 4826 6324 4853
rect 6396 4827 6404 4853
rect 6207 4796 6244 4804
rect 687 4776 944 4784
rect 1087 4776 1153 4784
rect 1247 4776 1633 4784
rect 1647 4776 1772 4784
rect 1807 4776 1992 4784
rect 2027 4776 2193 4784
rect 2207 4776 2353 4784
rect 2467 4776 2632 4784
rect 2667 4776 2873 4784
rect 2887 4776 3093 4784
rect 3347 4776 3573 4784
rect 4407 4776 4613 4784
rect 4627 4776 4693 4784
rect 5087 4776 5253 4784
rect 5307 4776 5453 4784
rect 6367 4776 6413 4784
rect 6436 4767 6444 4856
rect 1187 4756 1872 4764
rect 1907 4756 1973 4764
rect 2327 4756 2393 4764
rect 2627 4756 2933 4764
rect 3027 4756 3193 4764
rect 3827 4756 3913 4764
rect 4056 4756 4333 4764
rect 27 4736 393 4744
rect 987 4736 1013 4744
rect 1067 4736 1213 4744
rect 1236 4736 1513 4744
rect 1236 4724 1244 4736
rect 2007 4736 2313 4744
rect 2507 4736 2573 4744
rect 2587 4736 2612 4744
rect 2647 4736 2853 4744
rect 2907 4736 3273 4744
rect 3376 4736 3473 4744
rect 1127 4716 1244 4724
rect 1567 4716 1593 4724
rect 1607 4716 1693 4724
rect 1856 4716 1913 4724
rect 907 4696 1353 4704
rect 1856 4704 1864 4716
rect 2307 4716 2533 4724
rect 2556 4716 2793 4724
rect 1627 4696 1864 4704
rect 1967 4696 2292 4704
rect 2556 4704 2564 4716
rect 3187 4716 3253 4724
rect 3376 4724 3384 4736
rect 3667 4736 3853 4744
rect 4056 4744 4064 4756
rect 4507 4756 4693 4764
rect 5947 4756 5973 4764
rect 6420 4766 6444 4767
rect 6067 4756 6353 4764
rect 6427 4756 6444 4766
rect 6427 4753 6440 4756
rect 4007 4736 4064 4744
rect 4107 4736 4333 4744
rect 4387 4736 4853 4744
rect 5727 4736 5793 4744
rect 5807 4736 5993 4744
rect 3307 4716 3384 4724
rect 4087 4716 4953 4724
rect 4967 4716 5313 4724
rect 6167 4716 6333 4724
rect 2327 4696 2564 4704
rect 2707 4696 2892 4704
rect 2927 4696 2952 4704
rect 2987 4696 3233 4704
rect 3247 4696 3453 4704
rect 3527 4696 3733 4704
rect 3847 4696 4293 4704
rect 4347 4696 4433 4704
rect 5787 4696 5933 4704
rect 1007 4676 1073 4684
rect 1087 4676 1173 4684
rect 1407 4676 1713 4684
rect 1887 4676 2733 4684
rect 3007 4676 3073 4684
rect 3087 4676 3213 4684
rect 3567 4676 3633 4684
rect 3787 4676 3913 4684
rect 3927 4676 4073 4684
rect 5047 4676 5153 4684
rect 5207 4676 5393 4684
rect 5727 4676 5813 4684
rect 5927 4676 6153 4684
rect 847 4656 873 4664
rect 887 4656 1193 4664
rect 1427 4656 1573 4664
rect 1587 4656 1613 4664
rect 1667 4656 2033 4664
rect 2107 4656 2633 4664
rect 2736 4664 2744 4673
rect 2736 4656 3533 4664
rect 3547 4656 3753 4664
rect 4067 4656 4153 4664
rect 4616 4656 5513 4664
rect 4616 4647 4624 4656
rect 5527 4656 5833 4664
rect 5847 4656 6173 4664
rect 6367 4656 6433 4664
rect 967 4636 1033 4644
rect 1947 4636 2693 4644
rect 3047 4636 3133 4644
rect 3207 4636 3353 4644
rect 3367 4636 3653 4644
rect 3947 4636 4053 4644
rect 4507 4636 4612 4644
rect 4647 4636 5373 4644
rect 5387 4636 5713 4644
rect 5867 4636 6464 4644
rect 1107 4616 1373 4624
rect 1527 4616 1673 4624
rect 1727 4616 2073 4624
rect 2147 4616 2513 4624
rect 2907 4616 3153 4624
rect 3167 4616 3693 4624
rect 3767 4616 4093 4624
rect 4147 4616 4233 4624
rect 4396 4616 4873 4624
rect 127 4596 153 4604
rect 327 4596 653 4604
rect 1767 4596 2092 4604
rect 2127 4596 2713 4604
rect 2867 4596 3033 4604
rect 3127 4596 3313 4604
rect 3647 4596 3733 4604
rect 3867 4596 4013 4604
rect 4396 4604 4404 4616
rect 4887 4616 5033 4624
rect 5127 4616 6433 4624
rect 6456 4624 6464 4636
rect 6456 4616 6484 4624
rect 4207 4596 4404 4604
rect 4447 4596 4573 4604
rect 5007 4596 5233 4604
rect 5847 4596 6033 4604
rect 6047 4596 6213 4604
rect 6476 4596 6484 4616
rect 267 4576 333 4584
rect 727 4576 753 4584
rect 1227 4576 1344 4584
rect 167 4557 193 4565
rect 116 4544 124 4554
rect 116 4540 184 4544
rect 116 4536 187 4540
rect 173 4527 187 4536
rect 336 4527 344 4573
rect 387 4557 433 4565
rect 567 4557 633 4565
rect 476 4544 484 4554
rect 827 4557 853 4565
rect 476 4540 544 4544
rect 476 4536 547 4540
rect 533 4527 547 4536
rect 47 4515 73 4523
rect 87 4515 93 4523
rect 287 4496 393 4504
rect 467 4500 524 4504
rect 467 4496 527 4500
rect 513 4487 527 4496
rect 587 4496 653 4504
rect 776 4504 784 4553
rect 876 4526 884 4573
rect 936 4527 944 4553
rect 1316 4527 1324 4554
rect 1336 4544 1344 4576
rect 1476 4576 1573 4584
rect 1476 4564 1484 4576
rect 2247 4576 2433 4584
rect 2487 4576 2553 4584
rect 2607 4576 2653 4584
rect 3147 4576 3193 4584
rect 3207 4576 3233 4584
rect 3416 4576 3773 4584
rect 1467 4556 1484 4564
rect 1667 4556 1753 4564
rect 2047 4557 2093 4565
rect 1336 4536 1364 4544
rect 1107 4516 1153 4524
rect 1316 4516 1333 4527
rect 1320 4513 1333 4516
rect 1356 4524 1364 4536
rect 1356 4516 1393 4524
rect 727 4496 784 4504
rect 807 4496 913 4504
rect 1416 4505 1424 4553
rect 1596 4544 1604 4553
rect 1596 4536 1933 4544
rect 1447 4516 1513 4524
rect 1587 4516 1633 4524
rect 1707 4516 1773 4524
rect 2156 4526 2164 4573
rect 2176 4544 2184 4554
rect 2307 4556 2433 4564
rect 2527 4556 2753 4564
rect 2807 4557 2833 4565
rect 2176 4540 2224 4544
rect 2176 4536 2227 4540
rect 2213 4527 2227 4536
rect 2027 4516 2144 4524
rect 1416 4504 1440 4505
rect 1416 4496 1433 4504
rect 1420 4493 1433 4496
rect 1807 4496 1833 4504
rect 1907 4496 1953 4504
rect 2136 4504 2144 4516
rect 2256 4524 2264 4553
rect 2436 4544 2444 4553
rect 2436 4536 2524 4544
rect 2256 4516 2273 4524
rect 2407 4516 2493 4524
rect 2516 4524 2524 4536
rect 2756 4527 2764 4554
rect 3047 4557 3113 4565
rect 3416 4564 3424 4576
rect 4227 4576 4273 4584
rect 4336 4576 4633 4584
rect 3540 4564 3553 4567
rect 3127 4556 3424 4564
rect 2933 4544 2947 4553
rect 2896 4540 2947 4544
rect 3536 4553 3553 4564
rect 3687 4556 3753 4564
rect 2893 4536 2944 4540
rect 2893 4527 2907 4536
rect 2516 4516 2593 4524
rect 2667 4516 2733 4524
rect 2756 4516 2773 4527
rect 2760 4513 2773 4516
rect 2906 4520 2907 4527
rect 2927 4516 2953 4524
rect 3087 4516 3133 4524
rect 3327 4516 3373 4524
rect 3467 4516 3513 4524
rect 2136 4496 2193 4504
rect 2316 4504 2324 4512
rect 3536 4507 3544 4553
rect 3667 4515 3813 4523
rect 3876 4523 3884 4554
rect 3987 4557 4013 4565
rect 4336 4564 4344 4576
rect 5367 4576 5413 4584
rect 5927 4584 5940 4587
rect 6180 4584 6193 4587
rect 5927 4573 5944 4584
rect 4327 4556 4344 4564
rect 4967 4556 5024 4564
rect 3867 4515 4033 4523
rect 4176 4524 4184 4553
rect 4176 4516 4213 4524
rect 4376 4524 4384 4553
rect 4553 4544 4567 4553
rect 4536 4536 4833 4544
rect 4347 4516 4384 4524
rect 4427 4515 4473 4523
rect 2316 4496 2553 4504
rect 2607 4496 2644 4504
rect 327 4476 373 4484
rect 827 4476 873 4484
rect 1327 4476 1372 4484
rect 1407 4476 1473 4484
rect 1527 4476 1793 4484
rect 2027 4476 2133 4484
rect 2227 4476 2293 4484
rect 2467 4476 2513 4484
rect 2636 4484 2644 4496
rect 3627 4496 3833 4504
rect 4536 4504 4544 4536
rect 5016 4527 5024 4556
rect 5507 4556 5533 4564
rect 4567 4515 4633 4523
rect 4707 4524 4720 4527
rect 4707 4513 4724 4524
rect 5376 4524 5384 4554
rect 5707 4557 5733 4565
rect 5156 4520 5384 4524
rect 5153 4516 5384 4520
rect 4507 4496 4544 4504
rect 4716 4504 4724 4513
rect 5153 4507 5167 4516
rect 4716 4496 4753 4504
rect 5596 4504 5604 4554
rect 5636 4524 5644 4554
rect 5636 4516 5753 4524
rect 5267 4496 5604 4504
rect 2636 4476 2693 4484
rect 3047 4476 3273 4484
rect 3367 4476 3413 4484
rect 3507 4476 3773 4484
rect 3876 4476 4133 4484
rect 627 4456 953 4464
rect 1427 4456 1573 4464
rect 1587 4456 1953 4464
rect 2007 4456 2233 4464
rect 2456 4464 2464 4473
rect 2367 4456 2464 4464
rect 2487 4456 2533 4464
rect 2727 4456 2833 4464
rect 3067 4456 3173 4464
rect 3447 4456 3653 4464
rect 3876 4464 3884 4476
rect 4407 4476 4593 4484
rect 4707 4476 4893 4484
rect 4907 4476 5113 4484
rect 5127 4476 5213 4484
rect 5533 4486 5547 4496
rect 5641 4496 5693 4504
rect 5776 4484 5784 4554
rect 5867 4556 5893 4564
rect 5936 4544 5944 4573
rect 6176 4573 6193 4584
rect 6220 4584 6233 4587
rect 6216 4573 6233 4584
rect 6007 4556 6064 4564
rect 5916 4536 5944 4544
rect 5916 4524 5924 4536
rect 5896 4520 5924 4524
rect 5893 4516 5924 4520
rect 5893 4507 5907 4516
rect 6056 4526 6064 4556
rect 6076 4527 6084 4554
rect 6176 4544 6184 4573
rect 6216 4564 6224 4573
rect 6156 4540 6184 4544
rect 6153 4536 6184 4540
rect 6196 4556 6224 4564
rect 6153 4527 6167 4536
rect 5987 4516 6013 4524
rect 6076 4516 6093 4527
rect 6080 4513 6093 4516
rect 5807 4496 5853 4504
rect 6196 4507 6204 4556
rect 6287 4557 6313 4565
rect 6247 4516 6273 4524
rect 6336 4526 6344 4573
rect 6476 4544 6484 4564
rect 6476 4536 6504 4544
rect 6447 4516 6484 4524
rect 6196 4496 6213 4507
rect 6200 4493 6213 4496
rect 5547 4476 5784 4484
rect 6496 4484 6504 4536
rect 6067 4476 6504 4484
rect 3707 4456 3884 4464
rect 4047 4456 4073 4464
rect 4307 4456 4533 4464
rect 5127 4456 5293 4464
rect 5607 4456 5833 4464
rect 5887 4456 6093 4464
rect 6107 4456 6193 4464
rect 367 4436 693 4444
rect 907 4436 973 4444
rect 1087 4436 1153 4444
rect 1516 4436 2333 4444
rect 1516 4424 1524 4436
rect 2376 4436 2613 4444
rect 2376 4427 2384 4436
rect 2707 4436 2853 4444
rect 3007 4436 3052 4444
rect 3087 4436 3193 4444
rect 3236 4436 3293 4444
rect 747 4416 1524 4424
rect 1547 4416 1633 4424
rect 1787 4416 1873 4424
rect 1927 4416 2053 4424
rect 2107 4416 2213 4424
rect 2367 4416 2384 4427
rect 2367 4413 2380 4416
rect 2407 4416 2492 4424
rect 2527 4416 2593 4424
rect 2787 4416 3033 4424
rect 3107 4416 3133 4424
rect 3236 4424 3244 4436
rect 3427 4436 3673 4444
rect 3787 4436 3973 4444
rect 4027 4436 4653 4444
rect 4887 4436 6433 4444
rect 3156 4416 3244 4424
rect 67 4396 133 4404
rect 347 4396 413 4404
rect 947 4396 1053 4404
rect 1307 4396 1333 4404
rect 1347 4396 1813 4404
rect 1827 4396 2112 4404
rect 2147 4396 2193 4404
rect 2627 4396 2764 4404
rect 2756 4387 2764 4396
rect 3156 4404 3164 4416
rect 3807 4416 3893 4424
rect 4267 4416 4373 4424
rect 4787 4416 5053 4424
rect 5067 4416 5193 4424
rect 5207 4416 5373 4424
rect 5487 4416 5573 4424
rect 5587 4416 5793 4424
rect 5807 4416 5833 4424
rect 6087 4416 6133 4424
rect 2907 4396 3164 4404
rect 3287 4396 3453 4404
rect 3727 4396 3833 4404
rect 3896 4404 3904 4413
rect 3896 4396 4713 4404
rect 5836 4396 6053 4404
rect 96 4376 173 4384
rect 56 4307 64 4333
rect 96 4306 104 4376
rect 467 4376 533 4384
rect 547 4376 613 4384
rect 627 4376 833 4384
rect 1756 4376 2013 4384
rect 1756 4367 1764 4376
rect 2567 4376 2632 4384
rect 2667 4376 2713 4384
rect 2767 4376 2813 4384
rect 2827 4376 3204 4384
rect 967 4356 993 4364
rect 1256 4356 1273 4364
rect 127 4336 164 4344
rect 156 4324 164 4336
rect 187 4336 233 4344
rect 433 4344 447 4353
rect 433 4340 533 4344
rect 436 4336 533 4340
rect 1107 4336 1193 4344
rect 1256 4344 1264 4356
rect 1287 4356 1513 4364
rect 1747 4356 1764 4367
rect 1747 4353 1760 4356
rect 1847 4356 1913 4364
rect 3196 4364 3204 4376
rect 3227 4376 3253 4384
rect 4827 4376 4913 4384
rect 4987 4376 5053 4384
rect 5836 4384 5844 4396
rect 5627 4376 5844 4384
rect 5907 4376 5953 4384
rect 6227 4376 6373 4384
rect 6447 4376 6484 4384
rect 2187 4356 2224 4364
rect 3196 4356 3233 4364
rect 1247 4336 1264 4344
rect 156 4316 264 4324
rect 256 4284 264 4316
rect 276 4304 284 4334
rect 536 4324 544 4334
rect 476 4320 544 4324
rect 473 4316 544 4320
rect 473 4307 487 4316
rect 276 4296 393 4304
rect 567 4296 593 4304
rect 607 4296 653 4304
rect 256 4276 413 4284
rect 147 4256 213 4264
rect 227 4256 253 4264
rect 416 4264 424 4273
rect 676 4264 684 4334
rect 1476 4336 1533 4344
rect 707 4295 773 4303
rect 887 4296 933 4304
rect 1436 4304 1444 4333
rect 1476 4324 1484 4336
rect 1556 4336 1673 4344
rect 1347 4296 1444 4304
rect 1456 4316 1484 4324
rect 1007 4276 1113 4284
rect 1456 4284 1464 4316
rect 1556 4307 1564 4336
rect 1207 4276 1464 4284
rect 1547 4273 1553 4287
rect 1716 4284 1724 4334
rect 1856 4324 1864 4334
rect 1796 4316 1864 4324
rect 1796 4304 1804 4316
rect 1747 4296 1804 4304
rect 1936 4304 1944 4333
rect 2076 4327 2084 4353
rect 2067 4316 2084 4327
rect 2067 4313 2080 4316
rect 1907 4296 1944 4304
rect 2156 4304 2164 4334
rect 2216 4324 2224 4356
rect 3276 4356 3433 4364
rect 2247 4336 2293 4344
rect 2387 4336 2433 4344
rect 2447 4337 2513 4345
rect 2567 4337 2593 4345
rect 2687 4337 2733 4345
rect 2756 4336 2993 4344
rect 2216 4316 2284 4324
rect 2276 4306 2284 4316
rect 2756 4324 2764 4336
rect 3276 4344 3284 4356
rect 3487 4356 3753 4364
rect 4427 4356 4633 4364
rect 5287 4356 5313 4364
rect 5367 4356 5453 4364
rect 5467 4356 5733 4364
rect 5747 4356 5913 4364
rect 3067 4336 3284 4344
rect 3316 4336 3413 4344
rect 2627 4316 2764 4324
rect 1987 4296 2164 4304
rect 2187 4295 2233 4303
rect 2507 4296 2533 4304
rect 3316 4306 3324 4336
rect 3587 4336 3633 4344
rect 3687 4337 3733 4345
rect 3867 4336 4013 4344
rect 3453 4324 3467 4333
rect 3436 4320 3467 4324
rect 3436 4316 3464 4320
rect 3436 4306 3444 4316
rect 2947 4296 3013 4304
rect 3467 4295 3553 4303
rect 3727 4296 3773 4304
rect 1687 4276 1724 4284
rect 1747 4276 1813 4284
rect 1896 4276 2513 4284
rect 416 4256 684 4264
rect 1896 4264 1904 4276
rect 2607 4276 2653 4284
rect 2847 4276 3233 4284
rect 3856 4284 3864 4334
rect 4347 4336 4393 4344
rect 4216 4324 4224 4334
rect 4547 4336 4593 4344
rect 4660 4344 4673 4347
rect 4656 4333 4673 4344
rect 4216 4316 4404 4324
rect 4396 4306 4404 4316
rect 4656 4306 4664 4333
rect 4756 4306 4764 4353
rect 4827 4337 4873 4345
rect 4967 4337 5173 4345
rect 5476 4336 5493 4344
rect 5436 4307 5444 4333
rect 4267 4296 4353 4304
rect 4407 4295 4453 4303
rect 4507 4295 4533 4303
rect 4947 4296 5093 4304
rect 5147 4296 5273 4304
rect 5287 4296 5353 4304
rect 5476 4287 5484 4336
rect 5520 4344 5533 4347
rect 5516 4333 5533 4344
rect 5916 4344 5924 4353
rect 5896 4336 5924 4344
rect 5516 4306 5524 4333
rect 5896 4306 5904 4336
rect 5707 4295 5793 4303
rect 3856 4276 3973 4284
rect 4687 4276 4833 4284
rect 5007 4276 5033 4284
rect 5476 4276 5493 4287
rect 5480 4273 5493 4276
rect 5587 4276 5633 4284
rect 6016 4284 6024 4334
rect 6227 4336 6293 4344
rect 6347 4336 6412 4344
rect 6447 4336 6484 4344
rect 6067 4296 6133 4304
rect 6187 4295 6213 4303
rect 6016 4276 6273 4284
rect 1607 4256 1904 4264
rect 1987 4256 2413 4264
rect 3047 4256 3513 4264
rect 3667 4256 3953 4264
rect 4027 4256 4513 4264
rect 4567 4256 4613 4264
rect 4627 4256 4793 4264
rect 5496 4256 5613 4264
rect 1687 4236 1733 4244
rect 1747 4236 1833 4244
rect 2047 4236 2133 4244
rect 2507 4236 2733 4244
rect 2747 4236 2872 4244
rect 2907 4236 3153 4244
rect 3656 4244 3664 4253
rect 3167 4236 3664 4244
rect 4727 4236 4813 4244
rect 4867 4236 5133 4244
rect 5496 4244 5504 4256
rect 5247 4236 5504 4244
rect 5607 4236 5633 4244
rect 5807 4236 6433 4244
rect 307 4216 473 4224
rect 1187 4216 1513 4224
rect 1667 4216 1713 4224
rect 1807 4216 1873 4224
rect 1887 4216 2093 4224
rect 2147 4216 2653 4224
rect 2727 4216 2973 4224
rect 3047 4216 3393 4224
rect 3707 4216 3893 4224
rect 4007 4216 4933 4224
rect 5487 4216 5533 4224
rect 5627 4216 5993 4224
rect 6007 4216 6313 4224
rect 787 4196 1593 4204
rect 1827 4196 1913 4204
rect 2067 4196 2893 4204
rect 3396 4204 3404 4213
rect 3396 4196 3733 4204
rect 3747 4196 3913 4204
rect 3927 4196 4013 4204
rect 4147 4196 4453 4204
rect 4467 4196 4873 4204
rect 5147 4196 5792 4204
rect 5827 4196 6053 4204
rect 907 4176 1053 4184
rect 1347 4176 1433 4184
rect 1787 4176 2033 4184
rect 2327 4176 2533 4184
rect 2627 4176 2773 4184
rect 3487 4176 3693 4184
rect 3827 4176 3893 4184
rect 4007 4176 4372 4184
rect 4407 4176 4473 4184
rect 4487 4176 4753 4184
rect 4907 4176 5613 4184
rect 507 4156 1313 4164
rect 1607 4156 1693 4164
rect 1787 4156 1873 4164
rect 2087 4156 3293 4164
rect 3367 4156 3393 4164
rect 3927 4156 4033 4164
rect 4087 4156 4113 4164
rect 4527 4156 4693 4164
rect 5407 4156 5593 4164
rect 5607 4156 5773 4164
rect 5787 4156 5853 4164
rect 6247 4156 6373 4164
rect 367 4136 1473 4144
rect 2107 4136 2372 4144
rect 2407 4136 2713 4144
rect 2887 4136 3033 4144
rect 3327 4136 3553 4144
rect 3847 4136 3893 4144
rect 3987 4136 4013 4144
rect 4247 4136 5693 4144
rect 1387 4116 1593 4124
rect 1647 4116 1772 4124
rect 1807 4116 2013 4124
rect 2187 4116 2213 4124
rect 2687 4116 2833 4124
rect 3167 4116 3473 4124
rect 3547 4116 3733 4124
rect 4387 4116 4513 4124
rect 4587 4116 4953 4124
rect 5696 4124 5704 4133
rect 5787 4136 5973 4144
rect 5696 4116 6273 4124
rect 1847 4096 2313 4104
rect 2487 4096 2993 4104
rect 3187 4096 3353 4104
rect 3367 4096 3453 4104
rect 3687 4096 3773 4104
rect 5067 4096 5133 4104
rect 6327 4096 6373 4104
rect 47 4076 193 4084
rect 207 4076 433 4084
rect 807 4076 873 4084
rect 1507 4076 1553 4084
rect 1647 4076 1853 4084
rect 1967 4076 2053 4084
rect 2356 4076 2453 4084
rect 147 4056 159 4064
rect 627 4056 673 4064
rect 867 4056 933 4064
rect 1167 4056 1193 4064
rect 1367 4056 1413 4064
rect 1607 4056 1793 4064
rect 107 4036 193 4044
rect 207 4037 293 4045
rect 427 4036 553 4044
rect 716 4036 733 4044
rect 67 3995 113 4003
rect 127 3996 273 4004
rect 447 3996 573 4004
rect 587 3995 673 4003
rect 716 3987 724 4036
rect 760 4044 773 4047
rect 756 4033 773 4044
rect 876 4036 993 4044
rect 756 4006 764 4033
rect 876 4006 884 4036
rect 1007 4036 1093 4044
rect 1136 4024 1144 4034
rect 1236 4036 1253 4044
rect 1016 4016 1144 4024
rect 927 3995 973 4003
rect 1016 3987 1024 4016
rect 1176 3987 1184 4033
rect 1236 4007 1244 4036
rect 1307 4037 1333 4045
rect 1567 4036 1604 4044
rect 1227 3996 1244 4007
rect 1473 4024 1487 4033
rect 1596 4027 1604 4036
rect 1647 4037 1753 4045
rect 2027 4036 2093 4044
rect 2356 4044 2364 4076
rect 2547 4076 2813 4084
rect 2827 4076 2953 4084
rect 3087 4076 3273 4084
rect 3447 4076 3644 4084
rect 2987 4056 3084 4064
rect 2267 4036 2364 4044
rect 2493 4044 2507 4053
rect 2493 4040 2544 4044
rect 2496 4036 2544 4040
rect 1473 4020 1573 4024
rect 1476 4016 1573 4020
rect 1596 4016 1613 4027
rect 1600 4013 1613 4016
rect 1873 4024 1887 4033
rect 2376 4024 2384 4034
rect 1873 4020 2384 4024
rect 1876 4016 2384 4020
rect 1227 3993 1240 3996
rect 1453 4004 1467 4013
rect 1287 4000 1467 4004
rect 1287 3996 1464 4000
rect 2536 4006 2544 4036
rect 2867 4036 3033 4044
rect 3076 4044 3084 4056
rect 3127 4056 3213 4064
rect 3407 4056 3453 4064
rect 3516 4056 3593 4064
rect 3076 4036 3093 4044
rect 3107 4036 3173 4044
rect 2556 4007 2564 4034
rect 3293 4024 3307 4033
rect 3356 4036 3493 4044
rect 3293 4020 3324 4024
rect 3296 4016 3324 4020
rect 1747 3996 1813 4004
rect 1867 3996 2044 4004
rect 1007 3976 1024 3987
rect 1007 3973 1020 3976
rect 1067 3976 1144 3984
rect 27 3956 213 3964
rect 707 3956 793 3964
rect 1136 3964 1144 3976
rect 1167 3976 1184 3987
rect 1167 3973 1180 3976
rect 1347 3976 1393 3984
rect 1587 3976 1833 3984
rect 1947 3976 2013 3984
rect 2036 3984 2044 3996
rect 2556 3996 2572 4007
rect 2560 3993 2572 3996
rect 2607 3996 2833 4004
rect 3036 3996 3053 4004
rect 2036 3976 2253 3984
rect 2267 3976 2333 3984
rect 3036 3984 3044 3996
rect 3067 3996 3153 4004
rect 3167 3996 3193 4004
rect 2527 3976 3044 3984
rect 3316 3986 3324 4016
rect 3356 4004 3364 4036
rect 3516 4024 3524 4056
rect 3636 4064 3644 4076
rect 3747 4076 3793 4084
rect 3807 4076 3864 4084
rect 3636 4056 3713 4064
rect 3636 4044 3644 4056
rect 3627 4036 3644 4044
rect 3476 4016 3524 4024
rect 3476 4006 3484 4016
rect 3347 3996 3364 4004
rect 3316 3985 3340 3986
rect 3316 3976 3333 3985
rect 3320 3973 3333 3976
rect 3407 3976 3433 3984
rect 3556 3984 3564 4033
rect 3796 4007 3804 4033
rect 3856 4024 3864 4076
rect 3907 4076 3993 4084
rect 4287 4076 4313 4084
rect 4847 4076 5013 4084
rect 5027 4076 5273 4084
rect 6007 4076 6193 4084
rect 4027 4056 4053 4064
rect 4167 4056 4213 4064
rect 4889 4056 5113 4064
rect 5347 4056 5413 4064
rect 5747 4056 5913 4064
rect 5927 4056 5953 4064
rect 6147 4056 6313 4064
rect 3887 4037 3913 4045
rect 4047 4037 4093 4045
rect 4136 4024 4144 4034
rect 4207 4036 4273 4044
rect 4367 4036 4433 4044
rect 4527 4036 4613 4044
rect 4627 4037 4653 4045
rect 4707 4036 4744 4044
rect 3856 4020 3984 4024
rect 3856 4016 3987 4020
rect 3973 4007 3987 4016
rect 3607 3996 3673 4004
rect 4056 4016 4144 4024
rect 4736 4024 4744 4036
rect 4767 4037 4833 4045
rect 4927 4037 4993 4045
rect 5107 4036 5153 4044
rect 4736 4016 4824 4024
rect 3507 3976 3713 3984
rect 4056 3984 4064 4016
rect 4076 4000 4113 4004
rect 3907 3976 4064 3984
rect 4073 3996 4113 4000
rect 4073 3987 4087 3996
rect 4267 3995 4313 4003
rect 4567 3996 4773 4004
rect 4816 4006 4824 4016
rect 5096 4007 5104 4034
rect 5580 4044 5593 4047
rect 5187 4016 5424 4024
rect 5087 3996 5104 4007
rect 5416 4006 5424 4016
rect 5516 4007 5524 4034
rect 5087 3993 5100 3996
rect 5267 3996 5373 4004
rect 5507 3996 5524 4007
rect 5576 4033 5593 4044
rect 5836 4036 5853 4044
rect 5576 4006 5584 4033
rect 5836 4024 5844 4036
rect 6047 4036 6073 4044
rect 5796 4020 5844 4024
rect 5793 4016 5844 4020
rect 5793 4007 5807 4016
rect 5507 3993 5520 3996
rect 5847 3995 5913 4003
rect 6096 4004 6104 4053
rect 6336 4024 6344 4034
rect 6276 4016 6344 4024
rect 6276 4007 6284 4016
rect 6027 3996 6104 4004
rect 6267 3996 6284 4007
rect 6356 4004 6364 4053
rect 6336 4000 6364 4004
rect 6333 3996 6364 4000
rect 6267 3993 6280 3996
rect 6333 3987 6347 3996
rect 4167 3976 4244 3984
rect 1136 3956 1313 3964
rect 1467 3956 1544 3964
rect -24 3936 493 3944
rect 947 3936 1333 3944
rect 1536 3944 1544 3956
rect 1867 3956 1893 3964
rect 2047 3956 2113 3964
rect 2327 3956 2393 3964
rect 2727 3956 3153 3964
rect 3207 3956 3533 3964
rect 3827 3956 4213 3964
rect 4236 3964 4244 3976
rect 4607 3976 4633 3984
rect 4647 3976 4753 3984
rect 5987 3976 6133 3984
rect 4236 3956 4333 3964
rect 4427 3956 4453 3964
rect 5627 3956 5673 3964
rect 6367 3956 6433 3964
rect 1536 3936 1653 3944
rect 2207 3936 2293 3944
rect 2427 3936 2573 3944
rect 2587 3936 2733 3944
rect 2967 3936 3013 3944
rect 3767 3936 3793 3944
rect 4027 3936 4253 3944
rect 5287 3936 5613 3944
rect 5787 3936 5832 3944
rect 5867 3936 5933 3944
rect 6047 3936 6173 3944
rect 6187 3936 6253 3944
rect 87 3916 633 3924
rect 967 3916 1113 3924
rect 1127 3916 1233 3924
rect 1687 3916 1973 3924
rect 2067 3916 2233 3924
rect 2347 3916 2773 3924
rect 3187 3916 3353 3924
rect 3847 3916 3912 3924
rect 3947 3916 4373 3924
rect 4987 3916 5093 3924
rect 5647 3916 5873 3924
rect 6007 3916 6053 3924
rect -24 3896 13 3904
rect 67 3896 353 3904
rect 667 3896 753 3904
rect 767 3896 833 3904
rect 1027 3896 1513 3904
rect 2356 3896 2493 3904
rect 427 3876 593 3884
rect 647 3876 873 3884
rect 987 3876 1173 3884
rect 1187 3876 1213 3884
rect 1267 3876 1293 3884
rect 1307 3876 1573 3884
rect 2007 3876 2173 3884
rect 2356 3884 2364 3896
rect 3427 3896 3493 3904
rect 3567 3896 3613 3904
rect 3887 3896 4033 3904
rect 4187 3896 4393 3904
rect 4447 3896 4513 3904
rect 4787 3896 5193 3904
rect 5807 3896 5933 3904
rect 6327 3896 6393 3904
rect 2187 3876 2364 3884
rect 2507 3876 2693 3884
rect 3267 3876 3473 3884
rect 3916 3876 4193 3884
rect 3916 3867 3924 3876
rect 4387 3876 4553 3884
rect 4907 3876 5113 3884
rect 5127 3876 5153 3884
rect 5347 3876 5393 3884
rect 5467 3876 5513 3884
rect 6167 3876 6353 3884
rect -24 3856 13 3864
rect 907 3856 953 3864
rect 1247 3856 1533 3864
rect 1607 3856 1673 3864
rect 1927 3856 2133 3864
rect 3167 3856 3233 3864
rect 3567 3856 3773 3864
rect 3907 3856 3924 3867
rect 3907 3853 3920 3856
rect 4507 3856 4573 3864
rect 4587 3856 4713 3864
rect 4767 3856 4853 3864
rect 5007 3856 5033 3864
rect 5187 3856 5353 3864
rect 5367 3856 5413 3864
rect 5427 3856 5493 3864
rect 5567 3856 5673 3864
rect 5727 3856 6053 3864
rect 6227 3856 6273 3864
rect 6367 3856 6433 3864
rect 127 3836 173 3844
rect -24 3816 53 3824
rect 267 3817 333 3825
rect 427 3824 440 3827
rect 427 3813 444 3824
rect 733 3824 747 3833
rect 567 3816 813 3824
rect 436 3804 444 3813
rect 436 3796 504 3804
rect -24 3776 73 3784
rect 496 3786 504 3796
rect 247 3776 373 3784
rect 627 3776 732 3784
rect 767 3775 793 3783
rect 847 3775 893 3783
rect 916 3784 924 3813
rect 976 3786 984 3833
rect 1927 3836 2212 3844
rect 2380 3844 2392 3847
rect 2247 3836 2392 3844
rect 2376 3833 2392 3836
rect 2427 3836 2633 3844
rect 3147 3836 3224 3844
rect 1127 3816 1233 3824
rect 1247 3816 1393 3824
rect 1587 3816 1724 3824
rect 916 3776 933 3784
rect 996 3784 1004 3814
rect 1716 3804 1724 3816
rect 1956 3804 1964 3814
rect 2027 3816 2073 3824
rect 2176 3804 2184 3814
rect 2227 3816 2273 3824
rect 2296 3816 2353 3824
rect 2296 3804 2304 3816
rect 1207 3796 1364 3804
rect 996 3776 1093 3784
rect 1187 3776 1213 3784
rect 1356 3784 1364 3796
rect 1596 3796 1644 3804
rect 1716 3796 1784 3804
rect 1956 3796 2184 3804
rect 2236 3796 2304 3804
rect 1356 3776 1373 3784
rect 1596 3784 1604 3796
rect 1427 3776 1604 3784
rect 1636 3784 1644 3796
rect 1636 3776 1753 3784
rect 1776 3784 1784 3796
rect 1776 3776 1793 3784
rect 1907 3775 2013 3783
rect 2067 3775 2113 3783
rect 2136 3784 2144 3796
rect 2236 3786 2244 3796
rect 2376 3786 2384 3833
rect 2487 3816 2652 3824
rect 2747 3816 2812 3824
rect 2833 3824 2847 3833
rect 2833 3820 2873 3824
rect 2836 3816 2873 3820
rect 3027 3816 3073 3824
rect 2673 3807 2687 3813
rect 2660 3806 2687 3807
rect 2667 3800 2687 3806
rect 2667 3796 2684 3800
rect 2667 3793 2680 3796
rect 2127 3776 2144 3784
rect 2167 3775 2193 3783
rect 2727 3776 2793 3784
rect 2976 3784 2984 3813
rect 3216 3787 3224 3836
rect 3367 3844 3380 3847
rect 3367 3833 3384 3844
rect 3447 3836 3593 3844
rect 3707 3836 3873 3844
rect 3947 3836 4033 3844
rect 4687 3836 4813 3844
rect 4887 3836 4953 3844
rect 4967 3836 4993 3844
rect 2847 3776 2984 3784
rect 3067 3775 3173 3783
rect 3276 3786 3284 3833
rect 3307 3816 3324 3824
rect 3316 3767 3324 3816
rect 3347 3816 3364 3824
rect 3356 3787 3364 3816
rect 3376 3804 3384 3833
rect 3636 3804 3644 3833
rect 4067 3817 4113 3825
rect 4167 3817 4193 3825
rect 4387 3816 4464 3824
rect 3376 3796 3404 3804
rect 3396 3784 3404 3796
rect 3596 3796 3644 3804
rect 4276 3796 4333 3804
rect 3396 3776 3433 3784
rect 3596 3784 3604 3796
rect 3476 3776 3604 3784
rect 3476 3767 3484 3776
rect 4007 3776 4033 3784
rect 4076 3780 4093 3784
rect 4073 3776 4093 3780
rect 4073 3767 4087 3776
rect 4276 3784 4284 3796
rect 4456 3804 4464 3816
rect 4487 3816 4604 3824
rect 4456 3796 4564 3804
rect 4556 3786 4564 3796
rect 4596 3786 4604 3816
rect 4727 3816 4773 3824
rect 5153 3824 5167 3833
rect 5153 3820 5213 3824
rect 5156 3816 5213 3820
rect 5327 3816 5453 3824
rect 5667 3816 5713 3824
rect 5787 3816 5964 3824
rect 5053 3804 5067 3813
rect 5053 3800 5233 3804
rect 5056 3796 5233 3800
rect 5516 3796 5553 3804
rect 4107 3776 4284 3784
rect 4307 3775 4353 3783
rect 4467 3775 4493 3783
rect 4787 3775 4833 3783
rect 4887 3775 4953 3783
rect 5027 3776 5113 3784
rect 5516 3784 5524 3796
rect 5347 3776 5524 3784
rect 5956 3786 5964 3816
rect 6116 3816 6193 3824
rect 6016 3787 6024 3813
rect 6116 3787 6124 3816
rect 5547 3775 5593 3783
rect 5807 3775 5833 3783
rect 6236 3784 6244 3814
rect 6236 3776 6313 3784
rect 107 3756 393 3764
rect 707 3756 833 3764
rect 1196 3756 1393 3764
rect 187 3736 213 3744
rect 287 3736 413 3744
rect 427 3736 633 3744
rect 1047 3736 1173 3744
rect 1196 3744 1204 3756
rect 1447 3756 1553 3764
rect 1807 3756 1933 3764
rect 2427 3756 2653 3764
rect 2907 3756 2933 3764
rect 2947 3756 2993 3764
rect 3316 3756 3333 3767
rect 3320 3753 3333 3756
rect 3467 3756 3484 3767
rect 3467 3753 3480 3756
rect 3627 3756 3792 3764
rect 3827 3756 3993 3764
rect 4127 3756 4153 3764
rect 4707 3756 4933 3764
rect 5507 3756 5553 3764
rect 6336 3764 6344 3833
rect 6396 3787 6404 3813
rect 6267 3756 6344 3764
rect 1187 3736 1204 3744
rect 1227 3736 1584 3744
rect 147 3716 193 3724
rect 207 3716 713 3724
rect 1347 3716 1553 3724
rect 1576 3724 1584 3736
rect 1607 3736 1733 3744
rect 2167 3736 2293 3744
rect 3107 3736 3313 3744
rect 3727 3736 3853 3744
rect 4407 3736 4613 3744
rect 5727 3736 5913 3744
rect 5927 3736 6033 3744
rect 1576 3716 1873 3724
rect 2187 3716 2613 3724
rect 3487 3716 3553 3724
rect 3807 3716 4173 3724
rect 4187 3716 4493 3724
rect 6227 3716 6373 3724
rect 367 3696 613 3704
rect 887 3696 1213 3704
rect 1287 3696 1513 3704
rect 1587 3696 2033 3704
rect 2147 3704 2160 3707
rect 2147 3693 2164 3704
rect 2527 3696 2813 3704
rect 2867 3696 3393 3704
rect 3407 3696 3493 3704
rect 3787 3696 4593 3704
rect 5347 3696 5753 3704
rect 1327 3676 1513 3684
rect 1747 3676 1852 3684
rect 2156 3684 2164 3693
rect 1887 3676 2124 3684
rect 2156 3676 2473 3684
rect 87 3656 513 3664
rect 627 3656 873 3664
rect 1087 3656 1153 3664
rect 1467 3656 1593 3664
rect 1647 3656 1693 3664
rect 2116 3664 2124 3676
rect 3527 3676 3593 3684
rect 3607 3676 3733 3684
rect 3827 3676 4053 3684
rect 4067 3676 4553 3684
rect 6147 3676 6333 3684
rect 2116 3656 2353 3664
rect 2427 3656 2453 3664
rect 2627 3656 2833 3664
rect 3607 3656 4044 3664
rect 4036 3647 4044 3656
rect 4316 3656 4573 3664
rect 4316 3647 4324 3656
rect 4627 3656 5073 3664
rect 267 3636 353 3644
rect 947 3636 1293 3644
rect 1476 3636 1953 3644
rect 27 3616 1253 3624
rect 1476 3624 1484 3636
rect 2347 3636 2493 3644
rect 2507 3636 2853 3644
rect 2907 3636 3493 3644
rect 3507 3636 3673 3644
rect 3727 3636 3933 3644
rect 4047 3636 4313 3644
rect 1347 3616 1484 3624
rect 1787 3616 2053 3624
rect 2607 3616 3113 3624
rect 3327 3616 3473 3624
rect 4207 3616 4353 3624
rect 4567 3616 4613 3624
rect 6187 3616 6413 3624
rect 167 3596 493 3604
rect 1067 3596 1273 3604
rect 1487 3596 1573 3604
rect 1596 3596 1673 3604
rect 527 3576 1153 3584
rect 1387 3576 1484 3584
rect 247 3556 313 3564
rect 1476 3564 1484 3576
rect 1596 3584 1604 3596
rect 2047 3596 2893 3604
rect 3647 3596 3873 3604
rect 5607 3596 5813 3604
rect 5827 3596 6133 3604
rect 6227 3596 6253 3604
rect 1507 3576 1604 3584
rect 2067 3576 2673 3584
rect 3347 3576 4373 3584
rect 4387 3576 5493 3584
rect 6167 3576 6433 3584
rect 1476 3556 1504 3564
rect 1267 3536 1313 3544
rect 1356 3536 1393 3544
rect 207 3517 273 3525
rect 467 3516 504 3524
rect 496 3504 504 3516
rect 536 3504 544 3514
rect 647 3516 713 3524
rect 727 3517 773 3525
rect 907 3517 953 3525
rect 1007 3517 1033 3525
rect 1127 3516 1213 3524
rect 1356 3524 1364 3536
rect 1256 3516 1364 3524
rect 496 3496 524 3504
rect 536 3500 564 3504
rect 536 3496 567 3500
rect 516 3486 524 3496
rect 553 3487 567 3496
rect 87 3476 373 3484
rect 387 3475 433 3483
rect 596 3484 604 3513
rect 816 3504 824 3514
rect 816 3496 864 3504
rect 576 3476 833 3484
rect 576 3464 584 3476
rect 856 3484 864 3496
rect 1256 3487 1264 3516
rect 856 3476 973 3484
rect 987 3476 1233 3484
rect 1256 3476 1273 3487
rect 1260 3473 1273 3476
rect 1376 3484 1384 3514
rect 1496 3524 1504 3556
rect 1627 3560 1704 3564
rect 1627 3556 1707 3560
rect 1693 3547 1707 3556
rect 1816 3556 1933 3564
rect 1527 3536 1653 3544
rect 1816 3544 1824 3556
rect 2007 3556 2132 3564
rect 2167 3556 2373 3564
rect 2516 3556 2813 3564
rect 1787 3536 1824 3544
rect 2127 3536 2313 3544
rect 2516 3544 2524 3556
rect 2867 3556 2953 3564
rect 3127 3556 3373 3564
rect 3387 3556 3633 3564
rect 3696 3560 3733 3564
rect 3693 3556 3733 3560
rect 3693 3547 3707 3556
rect 4287 3556 4613 3564
rect 4767 3556 4793 3564
rect 4967 3556 5133 3564
rect 5547 3556 5713 3564
rect 5807 3556 5853 3564
rect 6047 3556 6113 3564
rect 6267 3556 6353 3564
rect 2367 3536 2524 3544
rect 2667 3536 2693 3544
rect 3227 3536 3373 3544
rect 3867 3544 3880 3547
rect 3867 3533 3884 3544
rect 4027 3536 4153 3544
rect 1496 3516 1524 3524
rect 1347 3476 1384 3484
rect 1416 3487 1424 3513
rect 1416 3476 1433 3487
rect 1420 3473 1433 3476
rect 1516 3484 1524 3516
rect 1847 3516 1953 3524
rect 1967 3516 2033 3524
rect 2056 3516 2073 3524
rect 2056 3504 2064 3516
rect 2216 3504 2224 3514
rect 1896 3500 2064 3504
rect 1893 3496 2064 3500
rect 2156 3496 2224 3504
rect 1893 3487 1907 3496
rect 1516 3476 1533 3484
rect 1587 3476 1773 3484
rect 1827 3476 1872 3484
rect 2156 3484 2164 3496
rect 2149 3476 2164 3484
rect 2256 3484 2264 3514
rect 2207 3476 2264 3484
rect 2407 3517 2433 3525
rect 2827 3517 2893 3525
rect 2947 3516 3053 3524
rect 3067 3516 3084 3524
rect 2293 3504 2307 3513
rect 2536 3504 2544 3514
rect 2293 3496 2544 3504
rect 2293 3487 2307 3496
rect 2536 3484 2544 3496
rect 3076 3487 3084 3516
rect 3187 3516 3213 3524
rect 2387 3480 2424 3484
rect 2387 3476 2427 3480
rect 2536 3476 2564 3484
rect 2413 3467 2427 3476
rect 547 3456 584 3464
rect 1627 3456 1653 3464
rect 1887 3456 2093 3464
rect 2556 3464 2564 3476
rect 2687 3476 2713 3484
rect 2787 3475 2873 3483
rect 2927 3476 2973 3484
rect 3076 3476 3093 3487
rect 3080 3473 3093 3476
rect 3516 3483 3524 3513
rect 3636 3487 3644 3514
rect 3876 3524 3884 3533
rect 5867 3536 5913 3544
rect 6276 3536 6393 3544
rect 3876 3516 3933 3524
rect 4087 3516 4113 3524
rect 4367 3517 4413 3525
rect 4487 3516 4693 3524
rect 4767 3516 4853 3524
rect 4867 3516 4884 3524
rect 3716 3487 3724 3513
rect 3747 3504 3760 3507
rect 3747 3493 3764 3504
rect 3207 3475 3533 3483
rect 3627 3476 3644 3487
rect 3627 3473 3640 3476
rect 3756 3484 3764 3493
rect 3756 3476 3833 3484
rect 3887 3475 3913 3483
rect 3976 3484 3984 3513
rect 4876 3504 4884 3516
rect 4907 3517 4973 3525
rect 5067 3516 5173 3524
rect 5187 3516 5344 3524
rect 5336 3504 5344 3516
rect 5367 3516 5393 3524
rect 5587 3517 5633 3525
rect 5696 3504 5704 3514
rect 5987 3516 6093 3524
rect 6227 3524 6240 3527
rect 6227 3513 6244 3524
rect 4876 3496 5024 3504
rect 5336 3496 5704 3504
rect 3967 3476 3984 3484
rect 4307 3476 4353 3484
rect 4467 3475 4513 3483
rect 4887 3476 4953 3484
rect 5016 3486 5024 3496
rect 5167 3476 5273 3484
rect 5287 3476 5333 3484
rect 5556 3486 5564 3496
rect 5647 3476 5713 3484
rect 5816 3484 5824 3513
rect 5876 3487 5884 3513
rect 5816 3476 5833 3484
rect 6236 3486 6244 3513
rect 6276 3487 6284 3536
rect 6336 3487 6344 3513
rect 6056 3480 6113 3484
rect 6053 3476 6113 3480
rect 6053 3467 6067 3476
rect 2556 3456 2593 3464
rect 3047 3456 3213 3464
rect 4567 3456 4633 3464
rect 587 3436 613 3444
rect 667 3436 793 3444
rect 807 3436 1053 3444
rect 1207 3436 1253 3444
rect 1407 3436 1453 3444
rect 1527 3436 1713 3444
rect 1787 3436 1893 3444
rect 1947 3436 1973 3444
rect 2067 3436 2093 3444
rect 2187 3436 2713 3444
rect 3007 3436 3293 3444
rect 3487 3436 3693 3444
rect 3887 3436 3993 3444
rect 4827 3436 5133 3444
rect 5767 3436 5953 3444
rect 6027 3436 6233 3444
rect 267 3416 373 3424
rect 567 3416 713 3424
rect 847 3416 873 3424
rect 1327 3416 1353 3424
rect 1367 3416 1493 3424
rect 1507 3416 1673 3424
rect 1687 3416 1753 3424
rect 2287 3416 2313 3424
rect 2327 3416 2433 3424
rect 2447 3416 2553 3424
rect 2567 3416 2724 3424
rect 747 3396 1013 3404
rect 1167 3396 1964 3404
rect 327 3376 553 3384
rect 1267 3376 1353 3384
rect 1367 3376 1513 3384
rect 1807 3376 1933 3384
rect 1956 3384 1964 3396
rect 2087 3396 2153 3404
rect 2527 3396 2693 3404
rect 2716 3404 2724 3416
rect 2867 3416 3073 3424
rect 3087 3416 3193 3424
rect 3587 3416 3804 3424
rect 2716 3396 2973 3404
rect 1956 3376 2113 3384
rect 2607 3376 2913 3384
rect 3127 3376 3433 3384
rect 3627 3376 3733 3384
rect 3796 3384 3804 3416
rect 3847 3416 4093 3424
rect 4187 3416 4973 3424
rect 3827 3396 4013 3404
rect 4027 3396 4053 3404
rect 5607 3396 5853 3404
rect 6387 3396 6433 3404
rect 3796 3376 4533 3384
rect 4647 3376 4833 3384
rect 5987 3376 6193 3384
rect 67 3356 112 3364
rect 147 3356 233 3364
rect 707 3356 793 3364
rect 807 3356 953 3364
rect 1107 3356 1244 3364
rect 1236 3347 1244 3356
rect 1787 3356 2013 3364
rect 2027 3356 2224 3364
rect 2216 3347 2224 3356
rect 2247 3356 2572 3364
rect 2607 3356 2673 3364
rect 3467 3356 3533 3364
rect 4887 3356 4953 3364
rect 5247 3356 5293 3364
rect 5367 3356 5433 3364
rect 167 3336 333 3344
rect 487 3336 573 3344
rect 1147 3336 1212 3344
rect 1247 3336 1433 3344
rect 1447 3336 1553 3344
rect 1767 3336 2013 3344
rect 2227 3336 2293 3344
rect 2467 3336 2693 3344
rect 2767 3336 2833 3344
rect 2847 3336 3013 3344
rect 3147 3336 3233 3344
rect 3247 3336 3433 3344
rect 3567 3336 3633 3344
rect 3927 3336 4324 3344
rect 4316 3327 4324 3336
rect 4527 3336 4593 3344
rect 4787 3336 4853 3344
rect 5487 3336 5573 3344
rect 5747 3336 5793 3344
rect 5867 3336 6073 3344
rect 6227 3336 6373 3344
rect 107 3316 293 3324
rect 387 3316 513 3324
rect 687 3316 733 3324
rect 967 3324 980 3327
rect 967 3313 984 3324
rect 1347 3316 1373 3324
rect 1460 3326 1473 3327
rect 276 3296 333 3304
rect 136 3267 144 3293
rect 236 3264 244 3294
rect 276 3267 284 3296
rect 356 3296 399 3304
rect 187 3256 244 3264
rect 356 3266 364 3296
rect 587 3304 600 3307
rect 587 3293 604 3304
rect 627 3296 653 3304
rect 767 3297 933 3305
rect 976 3304 984 3313
rect 1467 3313 1473 3326
rect 976 3296 1193 3304
rect 1607 3297 1672 3305
rect 596 3284 604 3293
rect 596 3280 624 3284
rect 596 3276 627 3280
rect 613 3267 627 3276
rect 407 3255 453 3263
rect 716 3244 724 3293
rect 1273 3284 1287 3293
rect 1733 3304 1747 3313
rect 2076 3316 2273 3324
rect 1733 3300 1813 3304
rect 1736 3296 1813 3300
rect 2076 3307 2084 3316
rect 2316 3316 2373 3324
rect 1693 3284 1707 3293
rect 1273 3280 1364 3284
rect 1276 3276 1364 3280
rect 1356 3267 1364 3276
rect 1556 3280 1707 3284
rect 1556 3276 1704 3280
rect 1556 3267 1564 3276
rect 1816 3267 1824 3294
rect 2027 3304 2040 3307
rect 2027 3293 2044 3304
rect 2067 3296 2084 3307
rect 2067 3293 2080 3296
rect 2316 3304 2324 3316
rect 2747 3316 2793 3324
rect 4067 3316 4113 3324
rect 4316 3316 4333 3327
rect 4320 3313 4333 3316
rect 4927 3316 4972 3324
rect 5007 3316 5053 3324
rect 5067 3316 5093 3324
rect 5107 3316 5213 3324
rect 2107 3296 2324 3304
rect 2596 3296 2653 3304
rect 867 3256 953 3264
rect 667 3236 724 3244
rect 913 3247 927 3256
rect 1087 3256 1253 3264
rect 1267 3256 1333 3264
rect 1356 3256 1373 3267
rect 1360 3253 1373 3256
rect 1547 3256 1564 3267
rect 1547 3253 1560 3256
rect 1587 3256 1733 3264
rect 1807 3256 1824 3267
rect 1916 3264 1924 3293
rect 2036 3284 2044 3293
rect 2036 3276 2144 3284
rect 2136 3266 2144 3276
rect 2436 3284 2444 3294
rect 2596 3284 2604 3296
rect 2667 3297 2753 3305
rect 3087 3297 3113 3305
rect 2367 3276 2444 3284
rect 2556 3280 2604 3284
rect 2553 3276 2604 3280
rect 3196 3284 3204 3294
rect 3267 3296 3313 3304
rect 3327 3297 3353 3305
rect 3487 3296 3584 3304
rect 3196 3280 3304 3284
rect 3196 3276 3307 3280
rect 2553 3267 2567 3276
rect 3293 3267 3307 3276
rect 1916 3256 1933 3264
rect 1807 3253 1820 3256
rect 2987 3256 3033 3264
rect 3147 3255 3173 3263
rect 3576 3266 3584 3296
rect 3707 3297 3773 3305
rect 3816 3267 3824 3294
rect 3936 3284 3944 3294
rect 4047 3296 4224 3304
rect 3936 3276 4013 3284
rect 3816 3256 3833 3267
rect 3820 3253 3833 3256
rect 4216 3266 4224 3296
rect 4427 3296 4553 3304
rect 4567 3296 4673 3304
rect 3927 3255 4033 3263
rect 4087 3255 4133 3263
rect 4407 3256 4433 3264
rect 4547 3255 4573 3263
rect 4796 3264 4804 3313
rect 5267 3316 5413 3324
rect 5427 3316 5633 3324
rect 5647 3316 5813 3324
rect 5856 3324 5864 3333
rect 5856 3316 5904 3324
rect 4847 3296 5013 3304
rect 5107 3296 5124 3304
rect 5116 3284 5124 3296
rect 5147 3296 5173 3304
rect 5387 3296 5533 3304
rect 5896 3304 5904 3316
rect 5927 3316 5964 3324
rect 5956 3304 5964 3316
rect 6147 3316 6173 3324
rect 6347 3324 6360 3327
rect 6347 3313 6364 3324
rect 5896 3296 5944 3304
rect 5956 3296 6004 3304
rect 5676 3284 5684 3294
rect 5116 3276 5753 3284
rect 5936 3284 5944 3296
rect 5936 3276 5964 3284
rect 5956 3266 5964 3276
rect 5996 3266 6004 3296
rect 6356 3266 6364 3313
rect 6400 3304 6413 3307
rect 6396 3293 6413 3304
rect 6396 3266 6404 3293
rect 4796 3260 4964 3264
rect 4796 3256 4967 3260
rect 4953 3247 4967 3256
rect 5407 3255 5433 3263
rect 5567 3255 5593 3263
rect 6007 3256 6173 3264
rect 1956 3236 2313 3244
rect 127 3216 213 3224
rect 1627 3216 1773 3224
rect 1956 3224 1964 3236
rect 2547 3236 2573 3244
rect 2667 3236 2713 3244
rect 3347 3236 3453 3244
rect 3627 3236 3873 3244
rect 5127 3236 5153 3244
rect 5167 3236 5353 3244
rect 1787 3216 1964 3224
rect 2007 3216 2193 3224
rect 2367 3216 2544 3224
rect 647 3196 753 3204
rect 767 3196 793 3204
rect 1127 3196 1213 3204
rect 1227 3196 1453 3204
rect 2196 3204 2204 3213
rect 2196 3196 2473 3204
rect 2536 3204 2544 3216
rect 3027 3216 3073 3224
rect 3287 3216 3493 3224
rect 3947 3216 4153 3224
rect 4387 3216 4793 3224
rect 2536 3196 2773 3204
rect 2787 3196 2833 3204
rect 3227 3196 3413 3204
rect 3427 3196 3473 3204
rect 3807 3196 4853 3204
rect 4867 3196 4893 3204
rect 5047 3196 5233 3204
rect 5247 3196 5473 3204
rect 5496 3196 5833 3204
rect 1147 3176 1353 3184
rect 1587 3176 1893 3184
rect 2047 3176 2273 3184
rect 2347 3176 2413 3184
rect 2587 3176 2993 3184
rect 3327 3176 3373 3184
rect 3427 3176 3513 3184
rect 4367 3176 4753 3184
rect 4767 3176 4933 3184
rect 5087 3176 5133 3184
rect 5147 3176 5173 3184
rect 5496 3184 5504 3196
rect 6107 3196 6213 3204
rect 5387 3176 5504 3184
rect 187 3156 493 3164
rect 1187 3156 1233 3164
rect 1247 3156 1293 3164
rect 1407 3156 1513 3164
rect 1767 3156 1993 3164
rect 2647 3156 3213 3164
rect 3307 3156 3833 3164
rect 3847 3156 3873 3164
rect 4327 3156 5713 3164
rect 27 3136 153 3144
rect 167 3136 253 3144
rect 1367 3136 1513 3144
rect 1887 3136 1973 3144
rect 2127 3136 2333 3144
rect 3387 3136 3713 3144
rect 3727 3136 3793 3144
rect 5467 3136 5653 3144
rect 1187 3116 1333 3124
rect 1747 3116 1833 3124
rect 2387 3116 2432 3124
rect 2467 3116 2873 3124
rect 2887 3116 2933 3124
rect 3227 3116 3353 3124
rect 3487 3116 3833 3124
rect 4087 3116 4113 3124
rect 4347 3116 4453 3124
rect 5747 3116 6093 3124
rect 827 3096 1153 3104
rect 1367 3096 1653 3104
rect 2187 3096 2733 3104
rect 3027 3096 3093 3104
rect 3107 3096 3193 3104
rect 3547 3096 3713 3104
rect 3867 3096 4713 3104
rect 5447 3096 5833 3104
rect 6147 3096 6373 3104
rect 147 3076 713 3084
rect 1727 3076 1853 3084
rect 1967 3076 2053 3084
rect 2187 3076 2213 3084
rect 2427 3076 2573 3084
rect 2947 3076 3273 3084
rect 3507 3076 4433 3084
rect 4527 3076 4573 3084
rect 4867 3076 4953 3084
rect 5947 3076 6433 3084
rect 1547 3056 1693 3064
rect 1947 3056 2373 3064
rect 2447 3056 2533 3064
rect 4887 3056 5493 3064
rect 5507 3056 5593 3064
rect 6247 3056 6273 3064
rect 187 3036 273 3044
rect 487 3036 593 3044
rect 907 3036 1013 3044
rect 1447 3036 1573 3044
rect 1727 3036 1913 3044
rect 2047 3036 2304 3044
rect 147 3016 293 3024
rect 467 3016 553 3024
rect 567 3016 733 3024
rect 1087 3016 1273 3024
rect 1547 3016 1612 3024
rect 1647 3016 1693 3024
rect 2296 3024 2304 3036
rect 2396 3036 2553 3044
rect 2396 3024 2404 3036
rect 3607 3036 3733 3044
rect 3747 3036 3933 3044
rect 4027 3036 4353 3044
rect 4887 3036 5024 3044
rect 2296 3016 2404 3024
rect 2587 3016 2613 3024
rect 2787 3016 3013 3024
rect 5016 3027 5024 3036
rect 4247 3016 4373 3024
rect 5027 3016 5193 3024
rect 5867 3016 6033 3024
rect 67 2997 93 3005
rect 207 2997 253 3005
rect 847 2996 953 3004
rect 1007 2997 1053 3005
rect 1076 2996 1173 3004
rect 47 2956 113 2964
rect 136 2964 144 2994
rect 136 2956 164 2964
rect 156 2944 164 2956
rect 156 2936 293 2944
rect 447 2936 573 2944
rect 756 2944 764 2994
rect 1076 2984 1084 2996
rect 1347 2996 1473 3004
rect 1487 2997 1713 3005
rect 1867 2997 2113 3005
rect 2287 2996 2453 3004
rect 2467 2997 2493 3005
rect 856 2976 1084 2984
rect 1776 2984 1784 2994
rect 2727 2997 2792 3005
rect 1776 2976 2073 2984
rect 856 2966 864 2976
rect 2593 2984 2607 2993
rect 2536 2980 2607 2984
rect 2536 2976 2604 2980
rect 987 2955 1193 2963
rect 1527 2956 1593 2964
rect 1636 2956 2013 2964
rect 1636 2947 1644 2956
rect 2276 2956 2293 2964
rect 707 2936 764 2944
rect 1147 2936 1273 2944
rect 1387 2936 1553 2944
rect 1627 2936 1644 2947
rect 1627 2933 1640 2936
rect 1727 2936 1753 2944
rect 2276 2944 2284 2956
rect 2396 2960 2433 2964
rect 2393 2956 2433 2960
rect 2187 2936 2284 2944
rect 2393 2947 2407 2956
rect 2536 2947 2544 2976
rect 2676 2964 2684 2994
rect 2887 2997 2933 3005
rect 3107 2996 3173 3004
rect 3327 2996 3344 3004
rect 2813 2984 2827 2993
rect 2736 2980 2827 2984
rect 2736 2976 2824 2980
rect 2736 2964 2744 2976
rect 3336 2967 3344 2996
rect 3447 2997 3473 3005
rect 3667 2996 3704 3004
rect 2567 2956 2684 2964
rect 2716 2960 2744 2964
rect 2713 2956 2744 2960
rect 2713 2947 2727 2956
rect 2947 2956 2993 2964
rect 3147 2955 3233 2963
rect 3536 2947 3544 2994
rect 3696 2984 3704 2996
rect 3847 2997 3993 3005
rect 4067 2997 4093 3005
rect 4187 2997 4233 3005
rect 4707 2997 4733 3005
rect 4747 2996 4913 3004
rect 3696 2976 3733 2984
rect 4136 2984 4144 2994
rect 4056 2976 4144 2984
rect 3567 2956 3613 2964
rect 4056 2964 4064 2976
rect 4027 2956 4064 2964
rect 4076 2960 4113 2964
rect 4073 2956 4113 2960
rect 4073 2947 4087 2956
rect 4276 2964 4284 2994
rect 4276 2956 4393 2964
rect 4516 2964 4524 2994
rect 5027 2997 5053 3005
rect 5287 2997 5333 3005
rect 5547 2996 5633 3004
rect 5687 2997 5733 3005
rect 4447 2956 4524 2964
rect 4567 2955 4633 2963
rect 5096 2964 5104 2994
rect 5887 2996 5913 3004
rect 6296 2984 6304 3033
rect 6296 2976 6373 2984
rect 4947 2956 5173 2964
rect 5407 2955 5453 2963
rect 5607 2955 5653 2963
rect 5747 2956 5793 2964
rect 5987 2955 6032 2963
rect 6067 2956 6113 2964
rect 6167 2955 6233 2963
rect 2767 2936 2853 2944
rect 2907 2936 3033 2944
rect 3047 2936 3093 2944
rect 3107 2936 3253 2944
rect 87 2916 233 2924
rect 687 2916 893 2924
rect 1067 2916 1164 2924
rect 467 2896 533 2904
rect 1156 2904 1164 2916
rect 1407 2916 1512 2924
rect 1547 2916 1573 2924
rect 1707 2916 1793 2924
rect 1907 2916 1973 2924
rect 2207 2916 2293 2924
rect 2627 2916 2733 2924
rect 2896 2924 2904 2933
rect 2747 2916 2904 2924
rect 3087 2916 3153 2924
rect 3347 2916 3433 2924
rect 4267 2916 4433 2924
rect 5847 2916 5913 2924
rect 5927 2916 6113 2924
rect 6127 2916 6293 2924
rect 1107 2896 1144 2904
rect 1156 2896 1453 2904
rect 207 2876 253 2884
rect 647 2876 833 2884
rect 967 2876 1113 2884
rect 1136 2884 1144 2896
rect 2267 2896 2313 2904
rect 2327 2896 2593 2904
rect 3207 2896 3473 2904
rect 3727 2896 3773 2904
rect 3927 2896 4013 2904
rect 5847 2896 5893 2904
rect 1136 2876 1333 2884
rect 1847 2876 2053 2884
rect 2507 2876 2773 2884
rect 2827 2876 2913 2884
rect 2927 2876 3744 2884
rect 3736 2867 3744 2876
rect 4247 2876 4333 2884
rect 5987 2876 6013 2884
rect 6027 2876 6193 2884
rect 347 2856 513 2864
rect 587 2856 913 2864
rect 1167 2856 1313 2864
rect 1387 2856 1633 2864
rect 1647 2856 1813 2864
rect 1827 2856 1953 2864
rect 2287 2856 2633 2864
rect 3247 2856 3433 2864
rect 3747 2856 4213 2864
rect 4647 2856 4713 2864
rect 4727 2856 4873 2864
rect 227 2836 273 2844
rect 367 2836 1033 2844
rect 1447 2836 1773 2844
rect 2067 2836 2333 2844
rect 2347 2836 2433 2844
rect 3867 2836 4093 2844
rect 4527 2836 4573 2844
rect 4927 2836 5133 2844
rect 5707 2836 5813 2844
rect 5827 2836 6013 2844
rect 147 2816 173 2824
rect 267 2816 333 2824
rect 687 2816 733 2824
rect 827 2816 953 2824
rect 1087 2816 1113 2824
rect 1407 2816 1753 2824
rect 1807 2816 1973 2824
rect 2087 2816 2213 2824
rect 2227 2816 2344 2824
rect 507 2796 593 2804
rect 747 2796 1013 2804
rect 1507 2796 1624 2804
rect 67 2776 93 2784
rect 227 2784 240 2787
rect 227 2773 244 2784
rect 307 2776 333 2784
rect 427 2776 484 2784
rect 236 2746 244 2773
rect 476 2747 484 2776
rect 536 2776 893 2784
rect 536 2747 544 2776
rect 947 2776 973 2784
rect 1016 2764 1024 2793
rect 1247 2776 1373 2784
rect 876 2756 1024 2764
rect 167 2736 233 2744
rect 367 2735 393 2743
rect 876 2746 884 2756
rect 1016 2746 1024 2756
rect 1076 2747 1084 2774
rect 1156 2747 1164 2774
rect 1396 2776 1453 2784
rect 1396 2764 1404 2776
rect 1616 2784 1624 2796
rect 1547 2776 1604 2784
rect 1616 2776 1753 2784
rect 1256 2760 1404 2764
rect 787 2735 813 2743
rect 927 2735 953 2743
rect 1076 2736 1093 2747
rect 1080 2733 1093 2736
rect 1147 2736 1164 2747
rect 1253 2756 1404 2760
rect 1596 2764 1604 2776
rect 1773 2784 1787 2793
rect 1856 2796 1893 2804
rect 1856 2784 1864 2796
rect 2067 2796 2153 2804
rect 1773 2780 1864 2784
rect 1776 2776 1864 2780
rect 1876 2776 1893 2784
rect 1596 2756 1693 2764
rect 1253 2747 1267 2756
rect 1876 2764 1884 2776
rect 1847 2756 1884 2764
rect 1956 2747 1964 2773
rect 1147 2733 1160 2736
rect 1727 2735 1773 2743
rect 1276 2716 1573 2724
rect 27 2696 413 2704
rect 707 2696 853 2704
rect 1276 2704 1284 2716
rect 1587 2716 1753 2724
rect 1976 2724 1984 2774
rect 2175 2744 2183 2773
rect 2196 2747 2204 2773
rect 2316 2747 2324 2773
rect 2107 2736 2183 2744
rect 2336 2744 2344 2816
rect 2687 2816 2773 2824
rect 3227 2816 3273 2824
rect 3427 2816 3673 2824
rect 4407 2816 4793 2824
rect 5447 2816 5653 2824
rect 6047 2816 6293 2824
rect 2867 2796 3053 2804
rect 3807 2796 3973 2804
rect 3987 2796 4033 2804
rect 4056 2796 4133 2804
rect 2427 2776 2724 2784
rect 2527 2756 2693 2764
rect 2716 2747 2724 2776
rect 2336 2736 2413 2744
rect 2716 2736 2732 2747
rect 2720 2733 2732 2736
rect 2756 2746 2764 2793
rect 2796 2744 2804 2793
rect 2967 2776 2993 2784
rect 3307 2784 3320 2787
rect 3307 2773 3324 2784
rect 3427 2776 3773 2784
rect 3996 2776 4013 2784
rect 2796 2736 2833 2744
rect 3316 2746 3324 2773
rect 3996 2764 4004 2776
rect 4056 2784 4064 2796
rect 4867 2796 4953 2804
rect 4967 2796 4993 2804
rect 5247 2796 5293 2804
rect 4036 2776 4064 2784
rect 3756 2756 4004 2764
rect 2947 2736 3073 2744
rect 3567 2736 3633 2744
rect 3756 2744 3764 2756
rect 4036 2746 4044 2776
rect 4107 2776 4164 2784
rect 4156 2746 4164 2776
rect 4267 2776 4373 2784
rect 4467 2776 4504 2784
rect 4496 2764 4504 2776
rect 4587 2776 4653 2784
rect 5107 2776 5153 2784
rect 5327 2776 5433 2784
rect 5607 2776 5753 2784
rect 4496 2756 4673 2764
rect 4556 2746 4564 2756
rect 5476 2764 5484 2774
rect 5807 2776 5893 2784
rect 5947 2776 6053 2784
rect 5476 2760 5524 2764
rect 5476 2756 5527 2760
rect 5513 2747 5527 2756
rect 5827 2756 5924 2764
rect 3747 2736 3764 2744
rect 4956 2736 5173 2744
rect 1976 2716 2153 2724
rect 2347 2716 2513 2724
rect 2587 2716 2673 2724
rect 2907 2716 3253 2724
rect 3447 2716 3513 2724
rect 3767 2716 3913 2724
rect 4007 2716 4113 2724
rect 4127 2716 4193 2724
rect 1227 2696 1284 2704
rect 1727 2696 1952 2704
rect 1987 2696 2073 2704
rect 2927 2696 3213 2704
rect 3227 2696 3273 2704
rect 3287 2696 3353 2704
rect 4356 2704 4364 2732
rect 4387 2716 4433 2724
rect 4607 2716 4633 2724
rect 4956 2724 4964 2736
rect 5307 2736 5453 2744
rect 5916 2746 5924 2756
rect 5627 2735 5653 2743
rect 5787 2736 5873 2744
rect 6327 2736 6373 2744
rect 4647 2716 4964 2724
rect 4356 2696 4393 2704
rect 4407 2696 4473 2704
rect 4667 2696 4993 2704
rect 5467 2696 5573 2704
rect 5667 2696 6153 2704
rect 1187 2676 1273 2684
rect 1347 2676 1473 2684
rect 1527 2676 1833 2684
rect 1927 2676 2453 2684
rect 2727 2676 2893 2684
rect 4767 2676 5033 2684
rect 5047 2676 5133 2684
rect 207 2656 613 2664
rect 1947 2656 2433 2664
rect 2647 2656 3493 2664
rect 3507 2656 3593 2664
rect 5367 2656 5713 2664
rect 667 2636 933 2644
rect 987 2636 1173 2644
rect 1287 2636 1713 2644
rect 1767 2636 1913 2644
rect 1987 2636 2313 2644
rect 2607 2636 2713 2644
rect 2907 2636 3293 2644
rect 3627 2636 3833 2644
rect 127 2616 193 2624
rect 687 2616 1613 2624
rect 1747 2616 1933 2624
rect 2047 2616 2113 2624
rect 2427 2616 2504 2624
rect 2496 2607 2504 2616
rect 2627 2616 2653 2624
rect 2667 2616 2733 2624
rect 2747 2616 2833 2624
rect 5307 2616 5493 2624
rect 5507 2616 5793 2624
rect 1767 2596 2093 2604
rect 2147 2596 2173 2604
rect 2187 2596 2293 2604
rect 2307 2596 2393 2604
rect 2507 2596 2633 2604
rect 3027 2596 3073 2604
rect 3487 2596 4553 2604
rect 227 2576 713 2584
rect 1107 2576 1433 2584
rect 1507 2576 1633 2584
rect 1687 2576 1833 2584
rect 2007 2576 2053 2584
rect 2207 2576 2293 2584
rect 2687 2576 2793 2584
rect 3687 2576 4233 2584
rect 4247 2576 4293 2584
rect 4967 2576 5013 2584
rect 167 2556 273 2564
rect 287 2556 473 2564
rect 847 2556 1084 2564
rect 467 2536 493 2544
rect 1076 2544 1084 2556
rect 1147 2556 1413 2564
rect 1707 2556 2033 2564
rect 2087 2556 2253 2564
rect 2407 2556 2953 2564
rect 2967 2556 3193 2564
rect 3207 2556 3533 2564
rect 3547 2556 3713 2564
rect 1076 2536 1113 2544
rect 1247 2536 1373 2544
rect 1616 2536 1893 2544
rect 1616 2527 1624 2536
rect 2467 2536 3413 2544
rect 3587 2536 3653 2544
rect 3847 2536 4393 2544
rect 4927 2536 4953 2544
rect 5107 2536 5193 2544
rect 5807 2536 5973 2544
rect 27 2516 213 2524
rect 527 2516 733 2524
rect 887 2516 1153 2524
rect 1607 2516 1624 2527
rect 1607 2513 1620 2516
rect 1727 2516 1853 2524
rect 1967 2516 2213 2524
rect 2287 2516 2373 2524
rect 2696 2516 2853 2524
rect 867 2504 880 2507
rect 867 2493 884 2504
rect 1667 2496 1764 2504
rect 47 2477 113 2485
rect 127 2476 233 2484
rect 507 2476 533 2484
rect 667 2477 693 2485
rect 67 2435 133 2443
rect 147 2436 253 2444
rect 627 2436 713 2444
rect 347 2416 433 2424
rect 447 2416 573 2424
rect 836 2424 844 2474
rect 876 2444 884 2493
rect 967 2477 1013 2485
rect 1056 2447 1064 2474
rect 1296 2447 1304 2474
rect 1367 2477 1393 2485
rect 1416 2464 1424 2493
rect 1447 2476 1533 2484
rect 1627 2476 1733 2484
rect 1756 2464 1764 2496
rect 2107 2496 2173 2504
rect 2696 2504 2704 2516
rect 3467 2516 3973 2524
rect 5547 2516 5653 2524
rect 2407 2496 2704 2504
rect 2767 2496 2833 2504
rect 4107 2496 4113 2504
rect 4127 2496 4184 2504
rect 1807 2476 1884 2484
rect 1416 2456 1744 2464
rect 1756 2456 1784 2464
rect 1736 2447 1744 2456
rect 876 2436 893 2444
rect 947 2436 1033 2444
rect 1056 2436 1073 2447
rect 1060 2433 1073 2436
rect 1296 2436 1313 2447
rect 1300 2433 1313 2436
rect 1487 2440 1724 2444
rect 1487 2436 1727 2440
rect 1736 2436 1753 2447
rect 747 2416 844 2424
rect 1353 2424 1367 2433
rect 1713 2427 1727 2436
rect 1740 2433 1753 2436
rect 1353 2420 1513 2424
rect 1356 2416 1513 2420
rect 1527 2416 1633 2424
rect 1776 2424 1784 2456
rect 1876 2447 1884 2476
rect 1907 2476 2013 2484
rect 2036 2444 2044 2493
rect 4176 2488 4184 2496
rect 4367 2496 4413 2504
rect 2227 2476 2273 2484
rect 2307 2476 2533 2484
rect 2547 2476 2713 2484
rect 2907 2477 2993 2485
rect 3147 2477 3253 2485
rect 3347 2476 3453 2484
rect 3507 2476 3533 2484
rect 3547 2476 3573 2484
rect 3907 2476 3933 2484
rect 3987 2476 4084 2484
rect 2153 2464 2167 2473
rect 2153 2460 2324 2464
rect 2156 2456 2324 2460
rect 2036 2436 2193 2444
rect 2316 2444 2324 2456
rect 2316 2436 2333 2444
rect 1776 2416 1913 2424
rect 2316 2424 2324 2436
rect 2467 2436 2513 2444
rect 2633 2443 2647 2447
rect 2607 2435 2647 2443
rect 2633 2433 2647 2435
rect 2216 2416 2324 2424
rect 2787 2435 2853 2443
rect 3027 2436 3313 2444
rect 3967 2436 4033 2444
rect 4076 2446 4084 2476
rect 4187 2477 4213 2485
rect 4136 2444 4144 2474
rect 4136 2436 4233 2444
rect 4256 2444 4264 2474
rect 4527 2477 4673 2485
rect 4727 2477 4753 2485
rect 4807 2477 4833 2485
rect 4927 2477 5213 2485
rect 5227 2476 5253 2484
rect 5447 2476 5573 2484
rect 5987 2477 6033 2485
rect 6087 2476 6173 2484
rect 6227 2476 6273 2484
rect 6367 2476 6413 2484
rect 4376 2447 4384 2473
rect 4256 2436 4364 2444
rect 347 2396 513 2404
rect 767 2396 953 2404
rect 1127 2396 1293 2404
rect 1507 2396 1673 2404
rect 2216 2404 2224 2416
rect 3367 2416 3533 2424
rect 4356 2424 4364 2436
rect 4416 2436 4473 2444
rect 4416 2424 4424 2436
rect 4487 2436 4573 2444
rect 4827 2436 4933 2444
rect 4987 2435 5013 2443
rect 6067 2435 6113 2443
rect 6247 2435 6293 2443
rect 4356 2416 4424 2424
rect 6296 2424 6304 2432
rect 6296 2416 6373 2424
rect 1947 2396 2224 2404
rect 2396 2396 2684 2404
rect 307 2376 653 2384
rect 1027 2376 1093 2384
rect 1147 2376 1313 2384
rect 1327 2376 1413 2384
rect 1787 2376 1833 2384
rect 1847 2376 1873 2384
rect 2396 2384 2404 2396
rect 1927 2376 2404 2384
rect 2676 2387 2684 2396
rect 2747 2396 3093 2404
rect 3107 2396 3213 2404
rect 3267 2396 3433 2404
rect 3567 2396 3613 2404
rect 4627 2396 5033 2404
rect 5127 2396 5313 2404
rect 5327 2396 5413 2404
rect 2676 2376 2693 2387
rect 2680 2373 2693 2376
rect 4127 2376 4413 2384
rect 4667 2376 4713 2384
rect 5847 2376 5873 2384
rect 47 2356 73 2364
rect 87 2356 392 2364
rect 427 2356 613 2364
rect 1747 2356 2293 2364
rect 2307 2356 2352 2364
rect 2387 2356 2473 2364
rect 3287 2356 3333 2364
rect 3467 2356 3793 2364
rect 696 2336 1073 2344
rect 696 2327 704 2336
rect 1087 2336 1173 2344
rect 1367 2336 1713 2344
rect 1867 2336 2033 2344
rect 2207 2336 2553 2344
rect 2567 2336 2613 2344
rect 2787 2336 3233 2344
rect 3487 2336 4093 2344
rect 4227 2336 4333 2344
rect 4347 2336 4373 2344
rect 5927 2336 5973 2344
rect 467 2316 553 2324
rect 567 2316 693 2324
rect 1767 2316 2064 2324
rect 2056 2307 2064 2316
rect 2647 2316 2713 2324
rect 2847 2316 2913 2324
rect 3476 2324 3484 2333
rect 3327 2316 3484 2324
rect 3787 2316 3973 2324
rect 5567 2316 5593 2324
rect 6127 2316 6393 2324
rect 67 2296 233 2304
rect 287 2296 413 2304
rect 907 2296 1073 2304
rect 1287 2296 1313 2304
rect 1407 2296 1573 2304
rect 1587 2296 1773 2304
rect 1847 2296 1972 2304
rect 2067 2296 2124 2304
rect 1993 2287 2007 2293
rect 840 2284 853 2287
rect 836 2273 853 2284
rect 1980 2286 2007 2287
rect 96 2244 104 2273
rect 147 2256 193 2264
rect 96 2236 124 2244
rect 116 2226 124 2236
rect 296 2226 304 2273
rect 607 2256 633 2264
rect 736 2244 744 2273
rect 696 2236 744 2244
rect 187 2215 253 2223
rect 696 2224 704 2236
rect 687 2216 704 2224
rect 836 2224 844 2273
rect 996 2256 1033 2264
rect 727 2216 844 2224
rect 996 2224 1004 2256
rect 1136 2226 1144 2273
rect 967 2216 1004 2224
rect 1176 2207 1184 2273
rect 1247 2256 1393 2264
rect 1507 2256 1533 2264
rect 1647 2257 1693 2265
rect 1747 2256 1793 2264
rect 1933 2264 1947 2273
rect 1987 2280 2007 2286
rect 2116 2284 2124 2296
rect 2147 2296 2173 2304
rect 2247 2296 2513 2304
rect 2567 2296 2733 2304
rect 2867 2296 2973 2304
rect 3207 2296 3273 2304
rect 3687 2296 3793 2304
rect 5067 2296 5233 2304
rect 5287 2296 5313 2304
rect 5627 2296 5693 2304
rect 5867 2296 6073 2304
rect 1987 2276 2004 2280
rect 2116 2276 2193 2284
rect 1987 2273 2000 2276
rect 2727 2276 2793 2284
rect 3247 2276 3453 2284
rect 3527 2276 3913 2284
rect 4027 2276 4053 2284
rect 6400 2284 6413 2287
rect 6396 2273 6413 2284
rect 1856 2260 1947 2264
rect 1856 2256 1944 2260
rect 1216 2236 1304 2244
rect 1216 2226 1224 2236
rect 1296 2224 1304 2236
rect 1267 2216 1284 2224
rect 1296 2216 1373 2224
rect 587 2196 673 2204
rect 687 2196 813 2204
rect 1176 2196 1193 2207
rect 1180 2193 1193 2196
rect 1276 2204 1284 2216
rect 1396 2216 1413 2224
rect 1396 2204 1404 2216
rect 1856 2224 1864 2256
rect 2027 2257 2113 2265
rect 2436 2244 2444 2254
rect 1907 2236 2244 2244
rect 1727 2216 1864 2224
rect 1276 2196 1404 2204
rect 1473 2204 1487 2213
rect 2087 2216 2213 2224
rect 1473 2200 1573 2204
rect 1476 2196 1573 2200
rect 1887 2196 1933 2204
rect 1956 2196 2113 2204
rect 1227 2176 1493 2184
rect 1607 2176 1793 2184
rect 1956 2184 1964 2196
rect 2236 2204 2244 2236
rect 2396 2236 2444 2244
rect 2267 2215 2293 2223
rect 2396 2224 2404 2236
rect 2347 2216 2404 2224
rect 2456 2224 2464 2273
rect 2547 2256 2664 2264
rect 2656 2227 2664 2256
rect 2707 2256 2852 2264
rect 2936 2256 2973 2264
rect 2876 2227 2884 2254
rect 2427 2216 2464 2224
rect 2507 2215 2533 2223
rect 2867 2216 2884 2227
rect 2936 2226 2944 2256
rect 3296 2256 3333 2264
rect 3296 2226 3304 2256
rect 3616 2256 3653 2264
rect 2867 2213 2880 2216
rect 3087 2215 3253 2223
rect 3476 2224 3484 2253
rect 3407 2216 3484 2224
rect 3616 2207 3624 2256
rect 3936 2256 4033 2264
rect 3753 2244 3767 2253
rect 3716 2240 3767 2244
rect 3716 2236 3764 2240
rect 3716 2224 3724 2236
rect 3856 2227 3864 2254
rect 3936 2227 3944 2256
rect 4173 2264 4187 2273
rect 4147 2260 4187 2264
rect 4147 2256 4184 2260
rect 4196 2256 4273 2264
rect 4196 2244 4204 2256
rect 5147 2257 5173 2265
rect 5227 2257 5273 2265
rect 4156 2236 4204 2244
rect 3647 2216 3724 2224
rect 3747 2215 3773 2223
rect 3856 2216 3873 2227
rect 3860 2213 3873 2216
rect 4156 2226 4164 2236
rect 4227 2215 4253 2223
rect 4716 2224 4724 2254
rect 4687 2216 4724 2224
rect 4787 2215 4833 2223
rect 5247 2215 5313 2223
rect 5376 2207 5384 2273
rect 5407 2256 5444 2264
rect 5436 2244 5444 2256
rect 5467 2256 5513 2264
rect 5567 2256 5653 2264
rect 5676 2256 5733 2264
rect 5556 2244 5564 2254
rect 5436 2236 5504 2244
rect 5556 2240 5584 2244
rect 5556 2236 5587 2240
rect 5496 2226 5504 2236
rect 5573 2227 5587 2236
rect 5676 2226 5684 2256
rect 5947 2257 6013 2265
rect 6267 2257 6313 2265
rect 6356 2244 6364 2254
rect 6336 2236 6364 2244
rect 5727 2215 5853 2223
rect 6027 2216 6053 2224
rect 6336 2224 6344 2236
rect 6207 2216 6344 2224
rect 6396 2224 6404 2273
rect 6396 2216 6413 2224
rect 2236 2196 2293 2204
rect 2687 2196 2753 2204
rect 3107 2196 3193 2204
rect 3507 2196 3553 2204
rect 4127 2196 4193 2204
rect 4207 2196 4293 2204
rect 5887 2196 5933 2204
rect 6287 2196 6373 2204
rect 1907 2176 1964 2184
rect 2027 2176 2213 2184
rect 2367 2176 2633 2184
rect 2847 2184 2860 2187
rect 2847 2173 2864 2184
rect 2907 2176 2933 2184
rect 2947 2176 3053 2184
rect 3227 2176 3373 2184
rect 3447 2176 3473 2184
rect 3487 2176 3593 2184
rect 3927 2176 4033 2184
rect 4247 2176 4433 2184
rect 5187 2176 5353 2184
rect 5813 2184 5827 2193
rect 5627 2180 5827 2184
rect 5627 2176 5824 2180
rect 447 2156 873 2164
rect 887 2156 993 2164
rect 1007 2156 1312 2164
rect 1347 2156 1733 2164
rect 1827 2156 1973 2164
rect 2167 2156 2233 2164
rect 2307 2156 2773 2164
rect 2787 2156 2813 2164
rect 2856 2164 2864 2173
rect 2856 2156 3073 2164
rect 3627 2156 3993 2164
rect 4067 2156 4213 2164
rect 4407 2156 4933 2164
rect 5047 2156 5453 2164
rect 5727 2156 5753 2164
rect 1207 2136 1273 2144
rect 1427 2136 1624 2144
rect 207 2116 533 2124
rect 547 2116 713 2124
rect 867 2116 1493 2124
rect 1616 2124 1624 2136
rect 1667 2136 1713 2144
rect 1807 2136 2053 2144
rect 2707 2136 2764 2144
rect 1616 2116 1633 2124
rect 1647 2116 1773 2124
rect 1787 2116 1912 2124
rect 1947 2116 2024 2124
rect 1427 2096 1613 2104
rect 1667 2096 1833 2104
rect 1927 2096 1993 2104
rect 2016 2104 2024 2116
rect 2107 2116 2413 2124
rect 2667 2116 2733 2124
rect 2756 2124 2764 2136
rect 5547 2136 5973 2144
rect 6327 2136 6373 2144
rect 2756 2116 3013 2124
rect 3167 2116 3673 2124
rect 3687 2116 3793 2124
rect 3847 2116 3873 2124
rect 3927 2116 3952 2124
rect 3987 2116 4113 2124
rect 4607 2116 4633 2124
rect 4907 2116 4953 2124
rect 4967 2116 5093 2124
rect 2016 2096 2433 2104
rect 2727 2096 2853 2104
rect 3907 2096 4433 2104
rect 787 2076 933 2084
rect 1367 2076 1533 2084
rect 1556 2076 2033 2084
rect 687 2056 753 2064
rect 1556 2064 1564 2076
rect 2167 2076 2353 2084
rect 3067 2076 3333 2084
rect 3647 2076 3913 2084
rect 5427 2076 5573 2084
rect 5587 2076 5673 2084
rect 5687 2076 6093 2084
rect 6107 2076 6273 2084
rect 1387 2056 1564 2064
rect 1767 2056 1812 2064
rect 1847 2056 1933 2064
rect 1987 2056 2084 2064
rect 87 2036 853 2044
rect 1367 2036 1473 2044
rect 1527 2036 1713 2044
rect 1767 2036 1893 2044
rect 1947 2036 2053 2044
rect 2076 2044 2084 2056
rect 2127 2056 2593 2064
rect 2616 2056 3933 2064
rect 2076 2036 2153 2044
rect 2616 2044 2624 2056
rect 4527 2056 4733 2064
rect 2447 2036 2624 2044
rect 2807 2036 3113 2044
rect 3187 2036 3353 2044
rect 3367 2036 3613 2044
rect 3967 2036 4333 2044
rect 5367 2036 5433 2044
rect 6147 2036 6233 2044
rect 247 2016 433 2024
rect 1507 2016 1833 2024
rect 2027 2016 2173 2024
rect 2187 2016 2653 2024
rect 3167 2016 3553 2024
rect 3687 2016 3944 2024
rect 3936 2007 3944 2016
rect 5307 2016 5573 2024
rect 5847 2016 6033 2024
rect 6387 2016 6433 2024
rect 147 1996 333 2004
rect 347 1996 393 2004
rect 527 1996 733 2004
rect 1067 1996 1093 2004
rect 1107 1996 1413 2004
rect 1547 1996 1933 2004
rect 2327 1996 2713 2004
rect 2827 1996 2993 2004
rect 3047 1996 3073 2004
rect 3127 1996 3213 2004
rect 3947 1996 3993 2004
rect 4007 1996 4513 2004
rect 4687 1996 5193 2004
rect 5647 2000 5784 2004
rect 5647 1996 5787 2000
rect -24 1976 73 1984
rect -24 1956 -16 1976
rect 847 1976 893 1984
rect 1027 1976 1433 1984
rect 1447 1976 1473 1984
rect 1727 1976 1893 1984
rect 1967 1984 1980 1987
rect 1967 1974 1984 1984
rect 1960 1973 1984 1974
rect 2047 1976 2073 1984
rect 5773 1987 5787 1996
rect 6067 1996 6153 2004
rect 2147 1976 2453 1984
rect 2567 1976 2593 1984
rect 3696 1976 3873 1984
rect 67 1957 273 1965
rect 287 1956 313 1964
rect 536 1927 544 1953
rect 616 1944 624 1954
rect 827 1956 973 1964
rect 1047 1956 1133 1964
rect 1567 1957 1753 1965
rect 616 1936 784 1944
rect 47 1915 73 1923
rect 127 1916 213 1924
rect 227 1916 253 1924
rect 467 1916 493 1924
rect 687 1915 753 1923
rect 776 1924 784 1936
rect 947 1936 1024 1944
rect 776 1916 893 1924
rect 1016 1924 1024 1936
rect 1016 1916 1113 1924
rect 307 1896 513 1904
rect 567 1896 653 1904
rect 1007 1896 1153 1904
rect 1276 1904 1284 1953
rect 1376 1927 1384 1953
rect 1736 1927 1744 1957
rect 1807 1956 1824 1964
rect 1816 1927 1824 1956
rect 1927 1956 1953 1964
rect 1976 1944 1984 1973
rect 2407 1956 2424 1964
rect 1956 1936 1984 1944
rect 1607 1915 1633 1923
rect 1736 1916 1753 1927
rect 1740 1913 1753 1916
rect 1907 1916 1933 1924
rect 1956 1907 1964 1936
rect 2136 1924 2144 1953
rect 2107 1916 2144 1924
rect 2176 1924 2184 1954
rect 2416 1944 2424 1956
rect 2707 1957 2972 1965
rect 3007 1956 3153 1964
rect 3327 1956 3373 1964
rect 3427 1956 3444 1964
rect 2347 1936 2504 1944
rect 2176 1916 2413 1924
rect 2496 1924 2504 1936
rect 2496 1916 2873 1924
rect 2887 1916 2913 1924
rect 2927 1915 3173 1923
rect 3436 1924 3444 1956
rect 3696 1926 3704 1976
rect 4256 1976 4593 1984
rect 4256 1968 4264 1976
rect 5567 1976 5593 1984
rect 3727 1957 3813 1965
rect 3987 1956 4033 1964
rect 4076 1927 4084 1954
rect 4147 1956 4173 1964
rect 4227 1957 4253 1965
rect 4507 1957 4533 1965
rect 4647 1956 4673 1964
rect 4867 1956 4933 1964
rect 4947 1956 4973 1964
rect 5347 1956 5493 1964
rect 5727 1957 5833 1965
rect 5967 1956 6013 1964
rect 4127 1936 4164 1944
rect 3436 1916 3533 1924
rect 3827 1916 4053 1924
rect 4076 1916 4093 1927
rect 4080 1913 4093 1916
rect 4156 1924 4164 1936
rect 4156 1916 4193 1924
rect 4547 1916 4613 1924
rect 5567 1915 5613 1923
rect 5907 1916 5993 1924
rect 6247 1916 6353 1924
rect 1167 1896 1413 1904
rect 1467 1896 1533 1904
rect 1547 1896 1573 1904
rect 2487 1896 2693 1904
rect 3847 1896 4133 1904
rect 4267 1896 4313 1904
rect 4327 1896 4433 1904
rect 767 1876 833 1884
rect 1227 1876 1293 1884
rect 2416 1876 3093 1884
rect 2416 1867 2424 1876
rect 3107 1876 3233 1884
rect 3247 1876 3393 1884
rect 3547 1876 3753 1884
rect 5427 1876 5593 1884
rect 5667 1876 5953 1884
rect 2087 1856 2133 1864
rect 2327 1856 2413 1864
rect 2867 1856 2953 1864
rect 4487 1856 4653 1864
rect 227 1836 413 1844
rect 1347 1836 1593 1844
rect 1907 1836 2093 1844
rect 2547 1836 2793 1844
rect 3027 1836 3073 1844
rect 3347 1836 3513 1844
rect 4007 1836 4073 1844
rect 4307 1836 5073 1844
rect 487 1816 593 1824
rect 707 1816 833 1824
rect 847 1816 1053 1824
rect 1067 1816 1273 1824
rect 1447 1816 1473 1824
rect 1927 1816 2153 1824
rect 2567 1816 2973 1824
rect 3296 1816 3453 1824
rect 727 1796 1033 1804
rect 1827 1796 1893 1804
rect 2127 1796 2333 1804
rect 2587 1796 2733 1804
rect 3296 1804 3304 1816
rect 3927 1816 3973 1824
rect 4147 1816 5753 1824
rect 3067 1796 3304 1804
rect 3367 1796 3773 1804
rect 4287 1796 4373 1804
rect 5487 1796 5653 1804
rect 5667 1796 5873 1804
rect 67 1776 113 1784
rect 127 1776 213 1784
rect 447 1776 533 1784
rect 547 1776 613 1784
rect 1027 1776 1153 1784
rect 1787 1776 1833 1784
rect 1847 1776 1912 1784
rect 1947 1776 2013 1784
rect 2027 1776 2053 1784
rect 2147 1776 2253 1784
rect 2907 1776 2953 1784
rect 3227 1776 3313 1784
rect 3447 1776 3733 1784
rect 4507 1776 4553 1784
rect 5187 1776 5293 1784
rect 5447 1776 5493 1784
rect 6147 1776 6313 1784
rect 827 1756 864 1764
rect 416 1736 513 1744
rect 416 1706 424 1736
rect 567 1736 653 1744
rect 596 1707 604 1736
rect 856 1707 864 1756
rect 1227 1756 1253 1764
rect 1587 1756 1633 1764
rect 2287 1756 2313 1764
rect 2876 1756 3113 1764
rect 927 1736 1113 1744
rect 1347 1736 1373 1744
rect 1527 1736 1664 1744
rect 27 1695 93 1703
rect 1656 1706 1664 1736
rect 1687 1736 1793 1744
rect 1876 1736 1973 1744
rect 1067 1695 1093 1703
rect 1707 1695 1733 1703
rect 1836 1704 1844 1734
rect 1876 1707 1884 1736
rect 2087 1736 2133 1744
rect 2467 1736 2513 1744
rect 2607 1736 2673 1744
rect 2747 1736 2853 1744
rect 1787 1696 1844 1704
rect 347 1676 373 1684
rect 727 1676 853 1684
rect 1147 1676 1253 1684
rect 1827 1676 1893 1684
rect 2087 1676 2133 1684
rect 2376 1684 2384 1733
rect 2813 1726 2827 1736
rect 2876 1706 2884 1756
rect 3127 1756 3273 1764
rect 5127 1756 5613 1764
rect 5627 1756 5833 1764
rect 2916 1736 3033 1744
rect 2916 1706 2924 1736
rect 3167 1736 3233 1744
rect 3356 1736 3373 1744
rect 3356 1724 3364 1736
rect 3447 1736 3473 1744
rect 3316 1716 3364 1724
rect 3496 1724 3504 1753
rect 3567 1736 3613 1744
rect 3687 1736 3724 1744
rect 3496 1716 3524 1724
rect 2587 1695 2653 1703
rect 2727 1695 2773 1703
rect 3027 1696 3133 1704
rect 3316 1704 3324 1716
rect 3187 1696 3324 1704
rect 3347 1696 3393 1704
rect 3467 1695 3493 1703
rect 3516 1687 3524 1716
rect 3716 1707 3724 1736
rect 3796 1736 3833 1744
rect 3547 1695 3573 1703
rect 3796 1706 3804 1736
rect 4067 1737 4113 1745
rect 4367 1736 4413 1744
rect 4567 1736 4584 1744
rect 4416 1724 4424 1734
rect 4416 1716 4444 1724
rect 4027 1695 4073 1703
rect 4147 1696 4253 1704
rect 4267 1696 4393 1704
rect 4436 1704 4444 1716
rect 4576 1707 4584 1736
rect 4607 1737 4673 1745
rect 5027 1736 5113 1744
rect 5256 1724 5264 1734
rect 5347 1736 5413 1744
rect 5487 1736 5553 1744
rect 5827 1736 5844 1744
rect 5176 1716 5264 1724
rect 4436 1696 4533 1704
rect 4667 1695 4713 1703
rect 5176 1704 5184 1716
rect 4907 1696 5184 1704
rect 5207 1695 5233 1703
rect 5507 1696 5533 1704
rect 5596 1704 5604 1733
rect 5596 1696 5673 1704
rect 5767 1695 5793 1703
rect 5836 1687 5844 1736
rect 6207 1736 6253 1744
rect 6356 1724 6364 1734
rect 6216 1716 6364 1724
rect 6216 1706 6224 1716
rect 6127 1696 6173 1704
rect 6267 1695 6293 1703
rect 2307 1676 2433 1684
rect 5287 1676 5433 1684
rect 227 1656 653 1664
rect 887 1656 973 1664
rect 2047 1656 2133 1664
rect 2207 1656 2253 1664
rect 2267 1656 2393 1664
rect 2827 1656 3173 1664
rect 3247 1656 3473 1664
rect 3547 1656 3693 1664
rect 3953 1664 3967 1673
rect 3953 1660 4013 1664
rect 3956 1656 4013 1660
rect 4027 1656 4053 1664
rect 4107 1656 4313 1664
rect 4787 1656 4833 1664
rect 4847 1656 5113 1664
rect 5367 1656 5424 1664
rect 147 1636 253 1644
rect 1687 1636 2493 1644
rect 2547 1636 2713 1644
rect 3307 1636 3573 1644
rect 4207 1636 4253 1644
rect 5416 1644 5424 1656
rect 5867 1656 6193 1664
rect 5416 1636 5973 1644
rect 487 1616 673 1624
rect 947 1616 973 1624
rect 1047 1616 1893 1624
rect 1967 1616 2073 1624
rect 2127 1616 2753 1624
rect 2847 1616 3284 1624
rect 1407 1596 1733 1604
rect 2116 1604 2124 1613
rect 1947 1596 2124 1604
rect 2147 1596 2293 1604
rect 2307 1596 2533 1604
rect 2607 1596 2793 1604
rect 2887 1596 3073 1604
rect 3096 1596 3213 1604
rect 1767 1576 1833 1584
rect 1967 1576 2373 1584
rect 3096 1584 3104 1596
rect 3276 1604 3284 1616
rect 4587 1616 5153 1624
rect 5167 1616 5393 1624
rect 5407 1616 5533 1624
rect 3276 1596 3413 1604
rect 5587 1596 5853 1604
rect 2787 1576 3104 1584
rect 5127 1576 6053 1584
rect 507 1556 593 1564
rect 887 1556 1213 1564
rect 1427 1556 1753 1564
rect 1907 1556 2213 1564
rect 2227 1556 2713 1564
rect 5336 1556 5733 1564
rect 487 1536 753 1544
rect 1487 1536 1573 1544
rect 2027 1536 2253 1544
rect 2827 1536 3213 1544
rect 4447 1536 4473 1544
rect 4607 1536 4793 1544
rect 4807 1536 4853 1544
rect 5336 1544 5344 1556
rect 4967 1536 5344 1544
rect 5407 1536 5473 1544
rect 407 1516 573 1524
rect 587 1516 633 1524
rect 647 1516 913 1524
rect 1587 1516 1713 1524
rect 2587 1516 2673 1524
rect 3447 1516 3633 1524
rect 4527 1516 4573 1524
rect 5627 1516 5673 1524
rect 5687 1516 6073 1524
rect 1447 1496 1493 1504
rect 1507 1496 1933 1504
rect 2007 1496 2053 1504
rect 2327 1496 2513 1504
rect 2627 1496 3033 1504
rect 3807 1496 4253 1504
rect 447 1476 544 1484
rect 536 1467 544 1476
rect 687 1476 813 1484
rect 1547 1476 2013 1484
rect 2387 1476 2633 1484
rect 2647 1476 2773 1484
rect 2907 1476 2953 1484
rect 3567 1476 3673 1484
rect 4527 1476 4633 1484
rect 5547 1476 6033 1484
rect 6047 1476 6173 1484
rect 547 1456 899 1464
rect 1627 1456 1653 1464
rect 2207 1456 2353 1464
rect 2987 1456 3273 1464
rect 3487 1456 3533 1464
rect 3547 1456 3733 1464
rect 5247 1456 5353 1464
rect 167 1436 233 1444
rect 247 1437 333 1445
rect 707 1436 1013 1444
rect 1087 1437 1113 1445
rect 1307 1436 1324 1444
rect 616 1407 624 1433
rect 1156 1424 1164 1434
rect 1156 1416 1233 1424
rect 1316 1407 1324 1436
rect 1547 1436 1673 1444
rect 1747 1436 1853 1444
rect 1867 1436 1953 1444
rect 2093 1444 2107 1453
rect 2093 1440 2133 1444
rect 2096 1436 2133 1440
rect 2267 1436 2413 1444
rect 2547 1436 2673 1444
rect 2816 1436 2953 1444
rect 2496 1424 2504 1433
rect 2447 1416 2504 1424
rect 67 1395 133 1403
rect 347 1396 373 1404
rect 427 1395 493 1403
rect 667 1396 713 1404
rect 767 1395 793 1403
rect 807 1396 853 1404
rect 967 1396 1033 1404
rect 1047 1396 1133 1404
rect 1567 1396 1693 1404
rect 1707 1395 1753 1403
rect 1767 1396 1833 1404
rect 1847 1396 1973 1404
rect 2027 1396 2113 1404
rect 2327 1395 2393 1403
rect 2527 1396 2693 1404
rect 2816 1404 2824 1436
rect 3007 1436 3073 1444
rect 3347 1436 3373 1444
rect 3627 1436 3713 1444
rect 3807 1437 3833 1445
rect 2807 1396 2824 1404
rect 2847 1395 2873 1403
rect 2927 1395 2973 1403
rect 3287 1395 3313 1403
rect 3547 1395 3593 1403
rect 3876 1404 3884 1434
rect 3967 1436 4012 1444
rect 4047 1436 4093 1444
rect 4187 1436 4593 1444
rect 4747 1436 4933 1444
rect 4947 1437 4993 1445
rect 5047 1436 5113 1444
rect 5527 1437 5553 1445
rect 5747 1436 5873 1444
rect 5887 1436 5993 1444
rect 6347 1437 6393 1445
rect 3747 1396 3884 1404
rect 5387 1396 5513 1404
rect 6267 1396 6373 1404
rect 287 1376 313 1384
rect 2187 1376 2393 1384
rect 2407 1376 2473 1384
rect 2747 1376 3193 1384
rect 3487 1376 3513 1384
rect 3527 1376 3973 1384
rect 4427 1376 4473 1384
rect 4487 1376 4613 1384
rect 4887 1376 5173 1384
rect 5187 1376 5333 1384
rect 5847 1376 5893 1384
rect 5907 1376 6193 1384
rect 147 1356 253 1364
rect 587 1356 633 1364
rect 747 1356 913 1364
rect 927 1356 1233 1364
rect 1247 1356 1273 1364
rect 1287 1356 1653 1364
rect 2567 1356 2653 1364
rect 2707 1356 2853 1364
rect 2907 1356 3093 1364
rect 3687 1356 3793 1364
rect 4147 1356 4233 1364
rect 367 1336 473 1344
rect 987 1336 1033 1344
rect 2087 1336 2233 1344
rect 2247 1336 2273 1344
rect 4367 1336 4633 1344
rect 5227 1336 5333 1344
rect 5347 1336 5433 1344
rect 5576 1340 5853 1344
rect 5573 1336 5853 1340
rect 5573 1327 5587 1336
rect 27 1316 233 1324
rect 1107 1316 1173 1324
rect 1187 1316 1413 1324
rect 2687 1316 2893 1324
rect 4507 1316 5013 1324
rect 307 1296 493 1304
rect 1507 1296 1733 1304
rect 2247 1296 2353 1304
rect 2367 1296 2433 1304
rect 2507 1296 2633 1304
rect 4687 1296 4733 1304
rect 5227 1296 5293 1304
rect 5607 1296 5653 1304
rect 6087 1296 6173 1304
rect 167 1276 213 1284
rect 487 1276 653 1284
rect 667 1276 893 1284
rect 1167 1276 1213 1284
rect 1616 1276 1813 1284
rect 1616 1267 1624 1276
rect 2607 1276 2813 1284
rect 2947 1276 3673 1284
rect 3867 1276 3993 1284
rect 4267 1276 4493 1284
rect 5087 1276 5193 1284
rect 5667 1276 5713 1284
rect 5827 1276 6313 1284
rect 127 1256 193 1264
rect 207 1256 273 1264
rect 427 1256 553 1264
rect 787 1256 812 1264
rect 847 1256 1073 1264
rect 1087 1256 1273 1264
rect 1547 1256 1613 1264
rect 1796 1256 1953 1264
rect 1796 1247 1804 1256
rect 2087 1256 2113 1264
rect 2587 1256 2693 1264
rect 2887 1256 3033 1264
rect 3267 1256 3433 1264
rect 5287 1256 5353 1264
rect 6047 1256 6113 1264
rect 67 1236 93 1244
rect 247 1236 293 1244
rect 307 1236 353 1244
rect 647 1236 693 1244
rect 1307 1236 1332 1244
rect 1367 1236 1453 1244
rect 1536 1236 1693 1244
rect 227 1216 284 1224
rect 176 1187 184 1213
rect 67 1175 93 1183
rect 276 1186 284 1216
rect 327 1216 373 1224
rect 396 1216 533 1224
rect 396 1184 404 1216
rect 556 1216 613 1224
rect 556 1186 564 1216
rect 887 1216 953 1224
rect 1027 1216 1073 1224
rect 1147 1216 1193 1224
rect 1256 1216 1273 1224
rect 653 1204 667 1213
rect 596 1200 667 1204
rect 596 1196 664 1200
rect 596 1186 604 1196
rect 327 1176 404 1184
rect 447 1176 553 1184
rect 727 1176 813 1184
rect 827 1176 933 1184
rect 1236 1184 1244 1214
rect 1256 1186 1264 1216
rect 1287 1216 1493 1224
rect 1416 1186 1424 1216
rect 1536 1186 1544 1236
rect 1707 1236 1793 1244
rect 1867 1236 1893 1244
rect 2267 1236 2293 1244
rect 2340 1244 2353 1247
rect 2336 1233 2353 1244
rect 2407 1236 2453 1244
rect 3440 1244 3453 1247
rect 3436 1233 3453 1244
rect 3927 1236 3973 1244
rect 4047 1236 4353 1244
rect 5167 1236 5233 1244
rect 5987 1236 6013 1244
rect 1567 1216 1604 1224
rect 1596 1187 1604 1216
rect 1927 1216 1984 1224
rect 1976 1187 1984 1216
rect 2007 1216 2073 1224
rect 2167 1216 2193 1224
rect 2276 1216 2313 1224
rect 1107 1176 1244 1184
rect 1327 1175 1373 1183
rect 1847 1175 1893 1183
rect 2236 1184 2244 1213
rect 2276 1187 2284 1216
rect 2227 1176 2244 1184
rect 2336 1186 2344 1233
rect 2427 1217 2493 1225
rect 2567 1216 2593 1224
rect 2636 1216 2673 1224
rect 2527 1176 2613 1184
rect 2636 1184 2644 1216
rect 2727 1217 2753 1225
rect 2827 1217 2993 1225
rect 3047 1217 3073 1225
rect 3127 1217 3153 1225
rect 3167 1216 3213 1224
rect 3436 1187 3444 1233
rect 3587 1216 3633 1224
rect 3707 1216 3733 1224
rect 4087 1216 4204 1224
rect 2627 1176 2644 1184
rect 2987 1176 3033 1184
rect 3047 1176 3233 1184
rect 4196 1186 4204 1216
rect 4327 1217 4372 1225
rect 4407 1216 4453 1224
rect 4707 1216 4813 1224
rect 4827 1217 4893 1225
rect 5067 1217 5133 1225
rect 5276 1216 5333 1224
rect 4367 1196 4484 1204
rect 3647 1175 3673 1183
rect 4007 1175 4053 1183
rect 4476 1186 4484 1196
rect 5276 1186 5284 1216
rect 5687 1224 5700 1227
rect 5687 1213 5704 1224
rect 6187 1216 6233 1224
rect 5696 1204 5704 1213
rect 5476 1196 5704 1204
rect 5896 1204 5904 1214
rect 5896 1196 6044 1204
rect 5476 1186 5484 1196
rect 4387 1176 4433 1184
rect 4587 1175 4613 1183
rect 5127 1175 5213 1183
rect 5327 1175 5353 1183
rect 5547 1176 5573 1184
rect 5696 1184 5704 1196
rect 5696 1176 5713 1184
rect 5787 1175 5813 1183
rect 5987 1175 6013 1183
rect 6036 1184 6044 1196
rect 6036 1176 6053 1184
rect 887 1156 973 1164
rect 1587 1156 1653 1164
rect 1667 1156 2013 1164
rect 2067 1156 2153 1164
rect 3467 1156 3513 1164
rect 4227 1156 4513 1164
rect 4527 1156 4793 1164
rect 6076 1164 6084 1214
rect 6356 1204 6364 1214
rect 6267 1196 6393 1204
rect 6347 1175 6433 1183
rect 5927 1156 6084 1164
rect 6207 1156 6253 1164
rect 147 1136 324 1144
rect 316 1124 324 1136
rect 687 1136 1093 1144
rect 2287 1136 2413 1144
rect 2587 1136 2653 1144
rect 2787 1136 3153 1144
rect 3567 1136 3833 1144
rect 4107 1136 4313 1144
rect 4367 1136 4393 1144
rect 5007 1136 5293 1144
rect 316 1116 1493 1124
rect 3967 1116 4333 1124
rect 4347 1116 5173 1124
rect 5447 1116 5833 1124
rect 5967 1116 6293 1124
rect 2427 1096 2493 1104
rect 2507 1096 2793 1104
rect 2807 1096 2853 1104
rect 3107 1096 3353 1104
rect 4147 1096 4213 1104
rect 4907 1096 5113 1104
rect 5747 1096 5933 1104
rect 1307 1076 1513 1084
rect 1567 1076 1773 1084
rect 1867 1076 2153 1084
rect 3407 1076 3613 1084
rect 4927 1076 5573 1084
rect 787 1056 2293 1064
rect 2307 1056 2393 1064
rect 3847 1056 3913 1064
rect 3927 1056 4133 1064
rect 5207 1056 5953 1064
rect 1167 1036 1313 1044
rect 1747 1036 2213 1044
rect 3687 1036 3753 1044
rect 4307 1036 5104 1044
rect 607 1016 673 1024
rect 687 1016 1273 1024
rect 1487 1016 1873 1024
rect 2007 1016 2073 1024
rect 2287 1016 2373 1024
rect 2387 1016 2713 1024
rect 3527 1016 3833 1024
rect 3947 1016 3973 1024
rect 4527 1016 4753 1024
rect 5096 1024 5104 1036
rect 5127 1036 5373 1044
rect 5096 1016 6013 1024
rect 1347 996 1453 1004
rect 2607 996 2693 1004
rect 3407 996 3473 1004
rect 3687 996 4113 1004
rect 4127 996 4233 1004
rect 4247 996 4933 1004
rect 4947 996 5413 1004
rect 927 976 1013 984
rect 1027 976 1153 984
rect 1167 976 1593 984
rect 2567 976 2653 984
rect 5307 976 6173 984
rect 407 956 773 964
rect 2127 956 2253 964
rect 2596 956 2733 964
rect 147 936 193 944
rect 220 944 233 947
rect 216 933 233 944
rect 1087 936 1133 944
rect 2367 936 2433 944
rect 2596 944 2604 956
rect 3227 956 3433 964
rect 4227 956 4593 964
rect 4687 956 4893 964
rect 4947 956 5032 964
rect 5067 956 5253 964
rect 2567 936 2604 944
rect 2696 936 2813 944
rect 47 916 93 924
rect 216 904 224 933
rect 267 917 333 925
rect 447 917 473 925
rect 727 916 833 924
rect 1327 916 1413 924
rect 1607 916 1673 924
rect 1687 917 1713 925
rect 1927 916 2013 924
rect 2167 916 2193 924
rect 2387 916 2424 924
rect 196 896 224 904
rect 196 884 204 896
rect 87 876 204 884
rect 347 876 373 884
rect 427 876 533 884
rect 747 876 773 884
rect 867 875 913 883
rect 1087 875 1133 883
rect 1287 875 1333 883
rect 1587 875 1653 883
rect 1787 876 1853 884
rect 2007 875 2073 883
rect 2287 876 2353 884
rect 2416 886 2424 916
rect 2696 924 2704 936
rect 2827 936 2953 944
rect 4107 936 5213 944
rect 5607 936 5713 944
rect 5987 936 6173 944
rect 2527 916 2704 924
rect 2747 916 2853 924
rect 3067 917 3113 925
rect 3167 916 3273 924
rect 3287 916 3644 924
rect 3636 904 3644 916
rect 3707 917 3793 925
rect 3907 916 3953 924
rect 4407 916 4473 924
rect 4487 917 4533 925
rect 4547 916 4773 924
rect 5027 917 5093 925
rect 5187 916 5333 924
rect 5447 916 5473 924
rect 5627 916 5813 924
rect 5827 917 5873 925
rect 5927 916 6044 924
rect 3636 896 4213 904
rect 6036 904 6044 916
rect 6067 917 6113 925
rect 6387 916 6484 924
rect 6036 896 6224 904
rect 2467 876 2533 884
rect 2887 875 2913 883
rect 3307 876 3333 884
rect 3787 875 3953 883
rect 4027 876 4093 884
rect 4627 875 4673 883
rect 4767 876 4913 884
rect 5647 875 5693 883
rect 5967 875 6073 883
rect 6127 876 6193 884
rect 6216 884 6224 896
rect 6216 876 6233 884
rect 127 856 152 864
rect 187 856 213 864
rect 587 856 633 864
rect 647 856 693 864
rect 1076 864 1084 872
rect 1007 856 1084 864
rect 1656 864 1664 872
rect 1656 856 1733 864
rect 2627 856 2833 864
rect 3047 856 3113 864
rect 3127 856 3173 864
rect 3607 856 3733 864
rect 4167 856 4193 864
rect 4207 856 4573 864
rect 5007 856 5053 864
rect 5067 856 5113 864
rect 5387 856 5573 864
rect 487 836 773 844
rect 787 836 1233 844
rect 2547 836 2573 844
rect 2587 836 2713 844
rect 2727 836 2933 844
rect 2987 836 3053 844
rect 5147 836 5273 844
rect 6047 836 6333 844
rect 47 816 233 824
rect 967 816 1393 824
rect 2327 816 2513 824
rect 2607 816 2633 824
rect 2747 816 2913 824
rect 2967 816 3093 824
rect 3147 816 3213 824
rect 3587 816 3633 824
rect 1187 796 1413 804
rect 1587 796 1893 804
rect 2767 796 2873 804
rect 3707 796 3853 804
rect 4307 796 4513 804
rect 4787 796 4933 804
rect 4987 796 5153 804
rect 167 776 633 784
rect 747 776 933 784
rect 2067 776 2153 784
rect 5787 776 5893 784
rect 436 756 513 764
rect 436 747 444 756
rect 656 756 1313 764
rect 656 747 664 756
rect 2207 756 2553 764
rect 2667 756 2713 764
rect 2907 756 2973 764
rect 4247 756 4313 764
rect 4327 756 4493 764
rect 4867 756 5113 764
rect 5127 756 5373 764
rect 327 736 433 744
rect 547 736 653 744
rect 767 736 813 744
rect 827 736 893 744
rect 1067 736 1153 744
rect 1527 736 1553 744
rect 1627 736 1913 744
rect 1927 736 2053 744
rect 2147 736 2333 744
rect 2347 736 2613 744
rect 2627 736 2753 744
rect 4687 736 5133 744
rect 727 716 953 724
rect 1407 716 1524 724
rect 167 696 253 704
rect 267 696 393 704
rect 487 696 573 704
rect 736 696 772 704
rect 736 666 744 696
rect 807 696 853 704
rect 916 696 1013 704
rect 916 666 924 696
rect 1127 696 1193 704
rect 127 656 233 664
rect 347 655 373 663
rect 427 656 493 664
rect 507 655 553 663
rect 967 655 1033 663
rect 1047 656 1173 664
rect 1236 664 1244 693
rect 1316 666 1324 713
rect 1347 697 1373 705
rect 1516 666 1524 716
rect 1787 716 1833 724
rect 2927 716 3153 724
rect 3507 716 3593 724
rect 3927 716 4013 724
rect 4547 716 4633 724
rect 5267 716 5313 724
rect 5667 716 5773 724
rect 5847 716 6313 724
rect 1676 700 1733 704
rect 1673 696 1733 700
rect 1673 687 1687 696
rect 1747 696 1873 704
rect 1940 704 1953 707
rect 1936 693 1953 704
rect 1996 696 2013 704
rect 1936 666 1944 693
rect 1996 667 2004 696
rect 2207 697 2233 705
rect 2387 697 2453 705
rect 2520 704 2533 707
rect 2516 693 2533 704
rect 2587 696 2653 704
rect 2676 696 2793 704
rect 1227 656 1244 664
rect 1367 655 1393 663
rect 2516 666 2524 693
rect 2676 666 2684 696
rect 2807 697 2893 705
rect 3067 696 3184 704
rect 3176 666 3184 696
rect 3207 696 3244 704
rect 3236 667 3244 696
rect 3347 696 3444 704
rect 2247 656 2313 664
rect 2927 655 2973 663
rect 3436 666 3444 696
rect 3467 696 3604 704
rect 3596 666 3604 696
rect 3667 697 3713 705
rect 4007 696 4173 704
rect 4296 696 4353 704
rect 4296 684 4304 696
rect 4467 696 4584 704
rect 4156 676 4304 684
rect 3767 655 3833 663
rect 4156 664 4164 676
rect 4576 666 4584 696
rect 4947 697 4973 705
rect 4127 656 4164 664
rect 4187 655 4333 663
rect 4387 656 4473 664
rect 4596 664 4604 694
rect 5347 704 5360 707
rect 5347 693 5364 704
rect 6067 696 6173 704
rect 5047 684 5060 687
rect 5047 673 5064 684
rect 4596 656 4733 664
rect 5056 664 5064 673
rect 5056 656 5193 664
rect 5356 666 5364 693
rect 5416 684 5424 694
rect 6287 696 6484 704
rect 5416 680 5464 684
rect 5416 676 5467 680
rect 5453 667 5467 676
rect 5287 656 5353 664
rect 5547 656 5593 664
rect 5767 656 5813 664
rect 6087 655 6133 663
rect 6227 656 6273 664
rect 6367 656 6484 664
rect 1627 636 1753 644
rect 2787 636 2873 644
rect 3227 636 3253 644
rect 3367 636 3653 644
rect 5207 636 5433 644
rect 1007 616 1373 624
rect 1987 616 2073 624
rect 2647 616 2713 624
rect 2847 616 2873 624
rect 2887 616 3033 624
rect 3427 616 3473 624
rect 3656 624 3664 633
rect 3656 616 3973 624
rect 4067 616 4453 624
rect 4467 616 4673 624
rect 3167 596 3533 604
rect 4056 604 4064 613
rect 3547 596 4064 604
rect 5187 596 5313 604
rect 5407 596 6033 604
rect 747 576 1193 584
rect 1947 576 2033 584
rect 4027 576 4253 584
rect 4627 576 5093 584
rect 5247 576 5873 584
rect 1447 556 1553 564
rect 3327 556 3753 564
rect 5927 556 6073 564
rect 887 536 933 544
rect 947 536 1733 544
rect 2207 536 2253 544
rect 3027 536 3153 544
rect 1107 516 1273 524
rect 1847 516 2333 524
rect 2347 516 2433 524
rect 5367 516 5453 524
rect 1407 496 1553 504
rect 1567 496 1753 504
rect 1767 496 1793 504
rect 1807 496 2173 504
rect 3107 496 3633 504
rect 3647 496 4013 504
rect 4707 496 4993 504
rect 987 476 1113 484
rect 1127 476 1153 484
rect 1587 476 1953 484
rect 2027 476 2373 484
rect 2567 476 2833 484
rect 3447 476 4513 484
rect 6047 476 6233 484
rect 27 456 433 464
rect 687 456 2233 464
rect 2927 456 3093 464
rect 707 436 793 444
rect 1087 436 1253 444
rect 2287 436 2473 444
rect 2487 436 2773 444
rect 3387 436 3473 444
rect 3487 436 3733 444
rect 3747 436 4153 444
rect 4947 436 4973 444
rect 5727 436 5753 444
rect 167 416 233 424
rect 1247 416 1293 424
rect 1307 416 1633 424
rect 1647 416 1693 424
rect 1707 416 1873 424
rect 1887 416 1993 424
rect 3047 416 3113 424
rect 4767 416 5453 424
rect 5480 424 5493 427
rect 5467 416 5493 424
rect 5480 413 5493 416
rect 6287 416 6373 424
rect 67 397 93 405
rect 207 397 273 405
rect 367 396 393 404
rect 407 397 473 405
rect 527 397 573 405
rect 707 404 720 407
rect 707 393 724 404
rect 747 396 804 404
rect 67 355 253 363
rect 347 355 413 363
rect 467 356 513 364
rect 716 364 724 393
rect 796 367 804 396
rect 1087 396 1184 404
rect 716 360 744 364
rect 716 356 747 360
rect 733 347 747 356
rect 1176 366 1184 396
rect 1367 397 1453 405
rect 1467 397 1573 405
rect 1696 396 1793 404
rect 1696 366 1704 396
rect 1807 396 1913 404
rect 2047 397 2073 405
rect 2127 396 2213 404
rect 2487 396 2553 404
rect 2687 396 2873 404
rect 2987 396 3073 404
rect 3336 396 3433 404
rect 1307 355 1373 363
rect 1467 355 1533 363
rect 1767 355 1813 363
rect 1887 355 1933 363
rect 1987 356 2013 364
rect 2367 356 2453 364
rect 2507 355 2573 363
rect 2787 355 2813 363
rect 2867 356 3033 364
rect 3336 366 3344 396
rect 3576 367 3584 394
rect 3767 396 3813 404
rect 3927 396 3973 404
rect 4047 396 4053 404
rect 4067 396 4173 404
rect 4307 396 4333 404
rect 4407 396 4473 404
rect 4487 396 4553 404
rect 4627 397 4653 405
rect 4676 396 4813 404
rect 3576 356 3593 367
rect 3580 353 3593 356
rect 3707 356 3793 364
rect 3807 356 4273 364
rect 4547 356 4613 364
rect 4676 366 4684 396
rect 5076 396 5393 404
rect 5056 384 5064 394
rect 5036 380 5064 384
rect 5033 376 5064 380
rect 5033 367 5047 376
rect 4947 356 4973 364
rect 5076 366 5084 396
rect 5627 396 5713 404
rect 5727 396 5793 404
rect 5887 396 5953 404
rect 5967 397 5993 405
rect 6047 396 6184 404
rect 5187 356 5233 364
rect 5836 364 5844 394
rect 5747 356 5844 364
rect 6027 356 6093 364
rect 6176 364 6184 396
rect 6176 356 6193 364
rect 127 336 153 344
rect 167 336 193 344
rect 847 336 913 344
rect 2776 344 2784 352
rect 2727 336 2784 344
rect 5127 336 5253 344
rect 5267 336 5793 344
rect 5807 336 5893 344
rect 687 316 753 324
rect 916 316 1013 324
rect 307 296 553 304
rect 916 304 924 316
rect 1307 316 1513 324
rect 1527 316 2233 324
rect 2567 316 2653 324
rect 3267 316 3453 324
rect 4487 316 4713 324
rect 5047 316 5093 324
rect 6107 316 6153 324
rect 6347 316 6393 324
rect 887 296 924 304
rect 987 296 1053 304
rect 1127 296 1493 304
rect 1667 296 1733 304
rect 1807 296 2033 304
rect 3827 296 4073 304
rect 6087 296 6293 304
rect 807 276 833 284
rect 2107 276 2393 284
rect 3407 276 3853 284
rect 4327 276 4433 284
rect 4447 276 5573 284
rect 5887 276 5953 284
rect 607 256 853 264
rect 1227 256 1533 264
rect 2607 256 2953 264
rect 3927 256 4053 264
rect 4167 256 4213 264
rect 4227 256 4553 264
rect 6307 256 6373 264
rect 187 236 333 244
rect 607 236 893 244
rect 907 236 932 244
rect 967 236 1553 244
rect 1567 236 1673 244
rect 1827 236 2233 244
rect 2867 236 2913 244
rect 2967 236 3073 244
rect 3787 236 3953 244
rect 5047 236 5364 244
rect 307 216 353 224
rect 656 216 1133 224
rect 656 204 664 216
rect 1147 216 1273 224
rect 1547 216 1793 224
rect 2347 216 2593 224
rect 407 196 664 204
rect 867 196 953 204
rect 1407 196 1813 204
rect 27 177 113 185
rect 227 177 313 185
rect 447 176 513 184
rect 687 176 784 184
rect 107 136 153 144
rect 247 135 293 143
rect 556 144 564 174
rect 776 164 784 176
rect 807 176 964 184
rect 776 156 924 164
rect 916 146 924 156
rect 556 136 653 144
rect 667 136 773 144
rect 956 144 964 176
rect 987 176 1004 184
rect 996 164 1004 176
rect 1027 177 1093 185
rect 1107 176 1153 184
rect 1167 176 1253 184
rect 1327 177 1353 185
rect 1727 176 1873 184
rect 1887 176 1913 184
rect 1987 177 2053 185
rect 2067 176 2133 184
rect 2267 176 2293 184
rect 996 156 1033 164
rect 1536 156 1613 164
rect 956 136 1013 144
rect 1536 146 1544 156
rect 2456 164 2464 174
rect 2247 156 2464 164
rect 1167 135 1233 143
rect 1307 135 1333 143
rect 1587 136 1653 144
rect 1707 136 1793 144
rect 2047 136 2213 144
rect 2476 146 2484 216
rect 2667 216 2713 224
rect 3007 216 3133 224
rect 3796 216 4044 224
rect 2767 196 2913 204
rect 3207 196 3393 204
rect 3547 196 3613 204
rect 3707 196 3753 204
rect 2507 176 2553 184
rect 2707 177 2733 185
rect 2840 184 2853 187
rect 2836 173 2853 184
rect 2980 184 2993 187
rect 2976 173 2993 184
rect 2407 135 2433 143
rect 2567 136 2753 144
rect 2836 146 2844 173
rect 2976 146 2984 173
rect 3016 146 3024 193
rect 3076 146 3084 193
rect 3196 164 3204 174
rect 3247 176 3313 184
rect 3467 176 3513 184
rect 3647 176 3673 184
rect 3196 156 3264 164
rect 2887 135 2933 143
rect 3147 136 3233 144
rect 3256 144 3264 156
rect 3796 146 3804 216
rect 4036 204 4044 216
rect 4107 216 4513 224
rect 5356 224 5364 236
rect 5356 216 6393 224
rect 4036 196 4153 204
rect 4467 196 4564 204
rect 3827 184 3840 187
rect 3827 173 3844 184
rect 4556 184 4564 196
rect 4447 176 4544 184
rect 4556 176 4584 184
rect 3836 146 3844 173
rect 3256 136 3293 144
rect 3347 135 3373 143
rect 3527 135 3573 143
rect 3627 135 3693 143
rect 3907 135 3953 143
rect 4016 144 4024 174
rect 4536 147 4544 176
rect 4576 164 4584 176
rect 4607 176 4753 184
rect 4576 156 4664 164
rect 4016 136 4133 144
rect 4467 135 4493 143
rect 4656 146 4664 156
rect 4727 135 4753 143
rect 4836 144 4844 174
rect 4887 176 4973 184
rect 5167 177 5213 185
rect 5236 176 5253 184
rect 5236 164 5244 176
rect 5367 176 5393 184
rect 5827 176 5913 184
rect 6167 177 6193 185
rect 6207 176 6233 184
rect 5116 156 5244 164
rect 5116 146 5124 156
rect 4836 136 4953 144
rect 5247 136 5333 144
rect 5487 135 5573 143
rect 5587 136 5633 144
rect 5707 136 5852 144
rect 5887 136 5933 144
rect 6047 135 6073 143
rect 6207 136 6273 144
rect 387 116 433 124
rect 1367 116 1493 124
rect 2247 116 2353 124
rect 4187 116 4213 124
rect 4527 116 4573 124
rect 5007 116 5033 124
rect 5167 116 5513 124
rect 5647 116 5973 124
rect 27 96 193 104
rect 547 96 733 104
rect 747 96 813 104
rect 1147 96 1573 104
rect 1627 96 1973 104
rect 2256 96 2733 104
rect 2256 87 2264 96
rect 2747 96 2793 104
rect 3127 96 4093 104
rect 4147 96 4413 104
rect 4627 96 4873 104
rect 4967 96 5073 104
rect 507 76 593 84
rect 1067 76 1193 84
rect 1207 76 1373 84
rect 2167 76 2253 84
rect 2727 76 3093 84
rect 3147 76 3753 84
rect 4547 76 4593 84
rect 4647 76 4933 84
rect 4987 76 5053 84
rect 5107 76 5193 84
rect 1127 56 1353 64
rect 1887 36 2193 44
rect 2547 36 3213 44
rect 3487 36 3673 44
rect 1407 16 1433 24
rect 2227 16 2573 24
rect 3947 16 4013 24
rect 4147 16 4333 24
use NOR2X1  _922_ digital_ETRI
timestamp 1701862152
transform -1 0 4170 0 -1 1830
box -12 -8 74 272
use INVX2  _923_ digital_ETRI
timestamp 1701862152
transform 1 0 4250 0 -1 1830
box -12 -8 52 272
use INVX1  _924_ digital_ETRI
timestamp 1701862152
transform -1 0 5790 0 -1 790
box -12 -8 52 272
use NAND2X1  _925_ digital_ETRI
timestamp 1702508443
transform -1 0 5930 0 1 790
box -12 -8 72 272
use OAI21X1  _926_ digital_ETRI
timestamp 1702508443
transform -1 0 6250 0 1 790
box -12 -8 92 272
use INVX2  _927_
timestamp 1701862152
transform -1 0 3810 0 -1 1830
box -12 -8 52 272
use NOR2X1  _928_
timestamp 1701862152
transform -1 0 3050 0 1 2870
box -12 -8 74 272
use AOI22X1  _929_ digital_ETRI
timestamp 1701862152
transform -1 0 4350 0 1 790
box -14 -8 114 272
use OAI21X1  _930_
timestamp 1702508443
transform -1 0 6090 0 1 790
box -12 -8 92 272
use INVX1  _931_
timestamp 1701862152
transform 1 0 5710 0 1 1310
box -12 -8 52 272
use NAND2X1  _932_
timestamp 1702508443
transform -1 0 6050 0 1 1310
box -12 -8 72 272
use OAI21X1  _933_
timestamp 1702508443
transform -1 0 6090 0 -1 1310
box -12 -8 92 272
use AOI22X1  _934_
timestamp 1701862152
transform 1 0 5350 0 -1 790
box -14 -8 114 272
use OAI21X1  _935_
timestamp 1702508443
transform -1 0 6110 0 -1 790
box -12 -8 92 272
use INVX1  _936_
timestamp 1701862152
transform 1 0 5110 0 -1 1830
box -12 -8 52 272
use NAND2X1  _937_
timestamp 1702508443
transform 1 0 5390 0 -1 1830
box -12 -8 72 272
use OAI21X1  _938_
timestamp 1702508443
transform 1 0 5250 0 -1 1310
box -12 -8 92 272
use AOI22X1  _939_
timestamp 1701862152
transform -1 0 5190 0 1 790
box -14 -8 114 272
use OAI21X1  _940_
timestamp 1702508443
transform 1 0 5090 0 -1 1310
box -12 -8 92 272
use INVX1  _941_
timestamp 1701862152
transform 1 0 5910 0 -1 270
box -12 -8 52 272
use NAND2X1  _942_
timestamp 1702508443
transform -1 0 6050 0 1 270
box -12 -8 72 272
use OAI21X1  _943_
timestamp 1702508443
transform -1 0 6210 0 1 270
box -12 -8 92 272
use AOI22X1  _944_
timestamp 1701862152
transform -1 0 5290 0 -1 790
box -14 -8 114 272
use OAI21X1  _945_
timestamp 1702508443
transform -1 0 5950 0 -1 790
box -12 -8 92 272
use INVX1  _946_
timestamp 1701862152
transform 1 0 1770 0 -1 3910
box -12 -8 52 272
use NAND2X1  _947_
timestamp 1702508443
transform 1 0 2050 0 -1 3910
box -12 -8 72 272
use OAI21X1  _948_
timestamp 1702508443
transform -1 0 1970 0 -1 3910
box -12 -8 92 272
use INVX1  _949_
timestamp 1701862152
transform -1 0 2350 0 1 2350
box -12 -8 52 272
use NAND2X1  _950_
timestamp 1702508443
transform 1 0 2330 0 -1 3910
box -12 -8 72 272
use OAI21X1  _951_
timestamp 1702508443
transform 1 0 2170 0 -1 3910
box -12 -8 92 272
use INVX2  _952_
timestamp 1701862152
transform 1 0 4450 0 -1 3390
box -12 -8 52 272
use NAND2X1  _953_
timestamp 1702508443
transform 1 0 3310 0 1 3910
box -12 -8 72 272
use OAI21X1  _954_
timestamp 1702508443
transform 1 0 3430 0 1 3910
box -12 -8 92 272
use INVX2  _955_
timestamp 1701862152
transform 1 0 3630 0 1 4430
box -12 -8 52 272
use NAND2X1  _956_
timestamp 1702508443
transform 1 0 3570 0 1 3910
box -12 -8 72 272
use OAI21X1  _957_
timestamp 1702508443
transform 1 0 3710 0 1 3910
box -12 -8 92 272
use NAND2X1  _958_
timestamp 1702508443
transform 1 0 1790 0 1 3390
box -12 -8 72 272
use OAI21X1  _959_
timestamp 1702508443
transform -1 0 1990 0 1 3390
box -12 -8 92 272
use NAND2X1  _960_
timestamp 1702508443
transform 1 0 2410 0 1 2870
box -12 -8 72 272
use OAI21X1  _961_
timestamp 1702508443
transform 1 0 2250 0 1 2870
box -12 -8 92 272
use NAND2X1  _962_
timestamp 1702508443
transform 1 0 2890 0 1 3390
box -12 -8 72 272
use OAI21X1  _963_
timestamp 1702508443
transform -1 0 3090 0 1 3390
box -12 -8 92 272
use NAND2X1  _964_
timestamp 1702508443
transform 1 0 2990 0 -1 3910
box -12 -8 72 272
use OAI21X1  _965_
timestamp 1702508443
transform -1 0 3210 0 -1 3910
box -12 -8 92 272
use INVX1  _966_
timestamp 1701862152
transform -1 0 4510 0 -1 790
box -12 -8 52 272
use NAND2X1  _967_
timestamp 1702508443
transform 1 0 3970 0 -1 790
box -12 -8 72 272
use OAI21X1  _968_
timestamp 1702508443
transform -1 0 4410 0 -1 790
box -12 -8 92 272
use INVX1  _969_
timestamp 1701862152
transform -1 0 5130 0 -1 790
box -12 -8 52 272
use NAND2X1  _970_
timestamp 1702508443
transform -1 0 4490 0 1 790
box -12 -8 72 272
use OAI21X1  _971_
timestamp 1702508443
transform -1 0 4650 0 -1 790
box -12 -8 92 272
use INVX1  _972_
timestamp 1701862152
transform 1 0 4970 0 -1 790
box -12 -8 52 272
use NAND2X1  _973_
timestamp 1702508443
transform -1 0 4570 0 1 270
box -12 -8 72 272
use OAI21X1  _974_
timestamp 1702508443
transform -1 0 4730 0 1 270
box -12 -8 92 272
use INVX1  _975_
timestamp 1701862152
transform -1 0 5250 0 1 270
box -12 -8 52 272
use NAND2X1  _976_
timestamp 1702508443
transform -1 0 5130 0 -1 270
box -12 -8 72 272
use OAI21X1  _977_
timestamp 1702508443
transform -1 0 5130 0 1 270
box -12 -8 92 272
use INVX1  _978_
timestamp 1701862152
transform 1 0 3790 0 1 270
box -12 -8 52 272
use NAND2X1  _979_
timestamp 1702508443
transform -1 0 3490 0 -1 270
box -12 -8 72 272
use OAI21X1  _980_
timestamp 1702508443
transform -1 0 3650 0 -1 270
box -12 -8 92 272
use INVX1  _981_
timestamp 1701862152
transform -1 0 5370 0 -1 270
box -12 -8 52 272
use NAND2X1  _982_
timestamp 1702508443
transform -1 0 4470 0 -1 270
box -12 -8 72 272
use OAI21X1  _983_
timestamp 1702508443
transform -1 0 5270 0 -1 270
box -12 -8 92 272
use INVX8  _984_ digital_ETRI
timestamp 1701862152
transform -1 0 5490 0 1 790
box -12 -8 114 272
use INVX1  _985_
timestamp 1701862152
transform -1 0 3310 0 1 790
box -12 -8 52 272
use NAND2X1  _986_
timestamp 1702508443
transform 1 0 5250 0 1 790
box -12 -8 72 272
use OAI21X1  _987_
timestamp 1702508443
transform 1 0 4570 0 1 790
box -12 -8 92 272
use INVX1  _988_
timestamp 1701862152
transform -1 0 3710 0 -1 1310
box -12 -8 52 272
use NAND2X1  _989_
timestamp 1702508443
transform -1 0 3890 0 -1 790
box -12 -8 72 272
use OAI21X1  _990_
timestamp 1702508443
transform 1 0 3730 0 1 790
box -12 -8 92 272
use NAND2X1  _991_
timestamp 1702508443
transform -1 0 4790 0 1 790
box -12 -8 72 272
use OAI21X1  _992_
timestamp 1702508443
transform -1 0 5650 0 1 790
box -12 -8 92 272
use NAND2X1  _993_
timestamp 1702508443
transform -1 0 5850 0 -1 1830
box -12 -8 72 272
use OAI21X1  _994_
timestamp 1702508443
transform -1 0 5910 0 1 1310
box -12 -8 92 272
use NAND2X1  _995_
timestamp 1702508443
transform -1 0 5250 0 1 1830
box -12 -8 72 272
use OAI21X1  _996_
timestamp 1702508443
transform -1 0 5310 0 -1 1830
box -12 -8 92 272
use NAND2X1  _997_
timestamp 1702508443
transform 1 0 5710 0 1 270
box -12 -8 72 272
use OAI21X1  _998_
timestamp 1702508443
transform -1 0 5910 0 1 270
box -12 -8 92 272
use INVX1  _999_
timestamp 1701862152
transform 1 0 6370 0 1 1310
box -12 -8 52 272
use NAND2X1  _1000_
timestamp 1702508443
transform -1 0 6230 0 -1 1830
box -12 -8 72 272
use OAI21X1  _1001_
timestamp 1702508443
transform -1 0 6370 0 -1 1830
box -12 -8 92 272
use INVX1  _1002_
timestamp 1701862152
transform 1 0 6350 0 1 1830
box -12 -8 52 272
use NAND2X1  _1003_
timestamp 1702508443
transform 1 0 6150 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1004_
timestamp 1702508443
transform -1 0 6370 0 -1 1310
box -12 -8 92 272
use INVX1  _1005_
timestamp 1701862152
transform 1 0 5210 0 1 1310
box -12 -8 52 272
use NAND2X1  _1006_
timestamp 1702508443
transform -1 0 5590 0 -1 1830
box -12 -8 72 272
use OAI21X1  _1007_
timestamp 1702508443
transform 1 0 5330 0 1 1310
box -12 -8 92 272
use INVX1  _1008_
timestamp 1701862152
transform 1 0 5990 0 1 1830
box -12 -8 52 272
use NAND2X1  _1009_
timestamp 1702508443
transform 1 0 6270 0 -1 270
box -12 -8 72 272
use OAI21X1  _1010_
timestamp 1702508443
transform -1 0 6350 0 1 270
box -12 -8 92 272
use NAND3X1  _1011_ digital_ETRI
timestamp 1702508443
transform 1 0 3370 0 1 1830
box -12 -8 92 272
use INVX1  _1012_
timestamp 1701862152
transform -1 0 2750 0 1 2350
box -12 -8 52 272
use INVX1  _1013_
timestamp 1701862152
transform 1 0 1770 0 1 2350
box -12 -8 52 272
use INVX1  _1014_
timestamp 1701862152
transform 1 0 3530 0 1 1830
box -12 -8 52 272
use OAI21X1  _1015_
timestamp 1702508443
transform 1 0 2750 0 1 1830
box -12 -8 92 272
use NAND2X1  _1016_
timestamp 1702508443
transform -1 0 3490 0 1 1310
box -12 -8 72 272
use NAND2X1  _1017_
timestamp 1702508443
transform -1 0 3370 0 -1 790
box -12 -8 72 272
use OAI21X1  _1018_
timestamp 1702508443
transform -1 0 3510 0 -1 790
box -12 -8 92 272
use AOI21X1  _1019_ digital_ETRI
timestamp 1702508443
transform 1 0 3210 0 1 1830
box -12 -8 92 272
use NAND3X1  _1020_
timestamp 1702508443
transform -1 0 3130 0 1 1830
box -12 -8 92 272
use INVX1  _1021_
timestamp 1701862152
transform -1 0 3050 0 -1 1830
box -12 -8 52 272
use NAND2X1  _1022_
timestamp 1702508443
transform 1 0 2710 0 -1 1830
box -12 -8 72 272
use OAI21X1  _1023_
timestamp 1702508443
transform 1 0 3110 0 -1 1830
box -12 -8 92 272
use INVX1  _1024_
timestamp 1701862152
transform 1 0 3270 0 -1 1830
box -12 -8 52 272
use INVX1  _1025_
timestamp 1701862152
transform 1 0 3370 0 -1 1830
box -12 -8 52 272
use NAND3X1  _1026_
timestamp 1702508443
transform 1 0 3490 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1027_
timestamp 1702508443
transform 1 0 3650 0 -1 1830
box -12 -8 72 272
use OR2X2  _1028_ digital_ETRI
timestamp 1702508443
transform -1 0 3630 0 1 1310
box -12 -8 92 272
use NAND2X1  _1029_
timestamp 1702508443
transform -1 0 3770 0 1 1310
box -12 -8 72 272
use NAND2X1  _1030_
timestamp 1702508443
transform -1 0 3890 0 1 1310
box -12 -8 72 272
use NAND2X1  _1031_
timestamp 1702508443
transform 1 0 4430 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1032_
timestamp 1702508443
transform 1 0 4030 0 -1 1310
box -12 -8 92 272
use NAND2X1  _1033_
timestamp 1702508443
transform 1 0 3430 0 1 270
box -12 -8 72 272
use INVX1  _1034_
timestamp 1701862152
transform -1 0 2890 0 1 790
box -12 -8 52 272
use INVX4  _1035_ digital_ETRI
timestamp 1701862152
transform 1 0 990 0 1 4430
box -12 -8 72 272
use OAI21X1  _1036_
timestamp 1702508443
transform 1 0 2850 0 -1 1830
box -12 -8 92 272
use INVX1  _1037_
timestamp 1701862152
transform -1 0 3110 0 1 1310
box -12 -8 52 272
use INVX1  _1038_
timestamp 1701862152
transform 1 0 2590 0 1 2350
box -12 -8 52 272
use INVX1  _1039_
timestamp 1701862152
transform 1 0 3190 0 1 1310
box -12 -8 52 272
use AOI21X1  _1040_
timestamp 1702508443
transform 1 0 2390 0 -1 1830
box -12 -8 92 272
use NAND3X1  _1041_
timestamp 1702508443
transform 1 0 2250 0 -1 1830
box -12 -8 92 272
use INVX1  _1042_
timestamp 1701862152
transform 1 0 2190 0 -1 1310
box -12 -8 52 272
use NOR2X1  _1043_
timestamp 1701862152
transform -1 0 2410 0 1 1310
box -12 -8 74 272
use OAI21X1  _1044_
timestamp 1702508443
transform -1 0 2850 0 1 1310
box -12 -8 92 272
use NAND2X1  _1045_
timestamp 1702508443
transform -1 0 2170 0 -1 1830
box -12 -8 72 272
use INVX1  _1046_
timestamp 1701862152
transform 1 0 2230 0 1 1310
box -12 -8 52 272
use OAI21X1  _1047_
timestamp 1702508443
transform 1 0 2470 0 1 1310
box -12 -8 92 272
use NAND3X1  _1048_
timestamp 1702508443
transform -1 0 3010 0 1 1310
box -12 -8 92 272
use NAND2X1  _1049_
timestamp 1702508443
transform -1 0 2690 0 1 1310
box -12 -8 72 272
use OAI21X1  _1050_
timestamp 1702508443
transform -1 0 2370 0 -1 1310
box -12 -8 92 272
use NAND3X1  _1051_
timestamp 1702508443
transform -1 0 2530 0 -1 1310
box -12 -8 92 272
use NAND2X1  _1052_
timestamp 1702508443
transform 1 0 2850 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1053_
timestamp 1702508443
transform 1 0 2550 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1054_
timestamp 1702508443
transform 1 0 2110 0 1 790
box -12 -8 72 272
use INVX1  _1055_
timestamp 1701862152
transform 1 0 2750 0 -1 790
box -12 -8 52 272
use NAND3X1  _1056_
timestamp 1702508443
transform 1 0 2870 0 -1 790
box -12 -8 92 272
use AOI21X1  _1057_
timestamp 1702508443
transform 1 0 2690 0 1 790
box -12 -8 92 272
use NAND3X1  _1058_
timestamp 1702508443
transform 1 0 2550 0 1 790
box -12 -8 92 272
use NAND2X1  _1059_
timestamp 1702508443
transform -1 0 3090 0 -1 790
box -12 -8 72 272
use OAI21X1  _1060_
timestamp 1702508443
transform 1 0 3150 0 -1 790
box -12 -8 92 272
use NAND2X1  _1061_
timestamp 1702508443
transform 1 0 4950 0 -1 270
box -12 -8 72 272
use AOI21X1  _1062_
timestamp 1702508443
transform -1 0 2670 0 -1 1310
box -12 -8 92 272
use OAI21X1  _1063_
timestamp 1702508443
transform 1 0 2610 0 -1 790
box -12 -8 92 272
use NAND2X1  _1064_
timestamp 1702508443
transform -1 0 1570 0 1 1830
box -12 -8 72 272
use NOR2X1  _1065_
timestamp 1701862152
transform -1 0 2350 0 -1 790
box -12 -8 74 272
use AOI22X1  _1066_
timestamp 1701862152
transform -1 0 2050 0 -1 1830
box -14 -8 114 272
use NOR2X1  _1067_
timestamp 1701862152
transform 1 0 2150 0 -1 790
box -12 -8 74 272
use OAI21X1  _1068_
timestamp 1702508443
transform -1 0 2130 0 -1 1310
box -12 -8 92 272
use NAND2X1  _1069_
timestamp 1702508443
transform -1 0 1550 0 -1 1830
box -12 -8 72 272
use NAND3X1  _1070_
timestamp 1702508443
transform 1 0 1950 0 1 1310
box -12 -8 92 272
use INVX1  _1071_
timestamp 1701862152
transform 1 0 2110 0 1 1310
box -12 -8 52 272
use AOI21X1  _1072_
timestamp 1702508443
transform -1 0 1870 0 1 1310
box -12 -8 92 272
use OAI21X1  _1073_
timestamp 1702508443
transform -1 0 1970 0 -1 1310
box -12 -8 92 272
use INVX1  _1074_
timestamp 1701862152
transform -1 0 1810 0 -1 1310
box -12 -8 52 272
use INVX1  _1075_
timestamp 1701862152
transform -1 0 1710 0 -1 1310
box -12 -8 52 272
use NAND3X1  _1076_
timestamp 1702508443
transform 1 0 1550 0 1 790
box -12 -8 92 272
use NAND3X1  _1077_
timestamp 1702508443
transform -1 0 2090 0 -1 790
box -12 -8 92 272
use INVX1  _1078_
timestamp 1701862152
transform -1 0 1650 0 -1 790
box -12 -8 52 272
use AOI21X1  _1079_
timestamp 1702508443
transform -1 0 1950 0 -1 790
box -12 -8 92 272
use OAI21X1  _1080_
timestamp 1702508443
transform 1 0 1730 0 -1 790
box -12 -8 92 272
use INVX1  _1081_
timestamp 1701862152
transform -1 0 1830 0 1 270
box -12 -8 52 272
use INVX1  _1082_
timestamp 1701862152
transform 1 0 1990 0 1 790
box -12 -8 52 272
use AOI21X1  _1083_
timestamp 1702508443
transform 1 0 1710 0 1 790
box -12 -8 92 272
use INVX1  _1084_
timestamp 1701862152
transform 1 0 1770 0 1 1830
box -12 -8 52 272
use NAND3X1  _1085_
timestamp 1702508443
transform -1 0 1870 0 -1 1830
box -12 -8 92 272
use INVX2  _1086_
timestamp 1701862152
transform -1 0 2650 0 -1 2350
box -12 -8 52 272
use OAI21X1  _1087_
timestamp 1702508443
transform 1 0 1630 0 1 1830
box -12 -8 92 272
use AOI21X1  _1088_
timestamp 1702508443
transform -1 0 1710 0 -1 1830
box -12 -8 92 272
use OAI21X1  _1089_
timestamp 1702508443
transform 1 0 1850 0 1 790
box -12 -8 92 272
use NAND3X1  _1090_
timestamp 1702508443
transform 1 0 1910 0 1 270
box -12 -8 92 272
use NAND2X1  _1091_
timestamp 1702508443
transform -1 0 2390 0 1 270
box -12 -8 72 272
use NOR2X1  _1092_
timestamp 1701862152
transform -1 0 2510 0 1 270
box -12 -8 74 272
use AOI22X1  _1093_
timestamp 1701862152
transform -1 0 2530 0 -1 790
box -14 -8 114 272
use OAI21X1  _1094_
timestamp 1702508443
transform 1 0 2810 0 1 270
box -12 -8 92 272
use NOR3X1  _1095_ digital_ETRI
timestamp 1701862152
transform -1 0 2750 0 1 270
box -12 -8 172 272
use INVX1  _1096_
timestamp 1701862152
transform 1 0 2950 0 1 270
box -12 -8 52 272
use NAND2X1  _1097_
timestamp 1702508443
transform -1 0 3130 0 1 270
box -12 -8 72 272
use OAI21X1  _1098_
timestamp 1702508443
transform 1 0 4550 0 -1 270
box -12 -8 92 272
use NAND2X1  _1099_
timestamp 1702508443
transform 1 0 3290 0 -1 270
box -12 -8 72 272
use INVX1  _1100_
timestamp 1701862152
transform -1 0 690 0 -1 270
box -12 -8 52 272
use OAI21X1  _1101_
timestamp 1702508443
transform -1 0 1710 0 1 270
box -12 -8 92 272
use OAI21X1  _1102_
timestamp 1702508443
transform 1 0 1510 0 -1 1310
box -12 -8 92 272
use INVX1  _1103_
timestamp 1701862152
transform -1 0 870 0 1 790
box -12 -8 52 272
use AOI21X1  _1104_
timestamp 1702508443
transform -1 0 1730 0 1 1310
box -12 -8 92 272
use INVX1  _1105_
timestamp 1701862152
transform 1 0 1270 0 1 1310
box -12 -8 52 272
use NAND3X1  _1106_
timestamp 1702508443
transform -1 0 1590 0 1 1310
box -12 -8 92 272
use NAND2X1  _1107_
timestamp 1702508443
transform 1 0 1390 0 1 1310
box -12 -8 72 272
use NAND3X1  _1108_
timestamp 1702508443
transform -1 0 1430 0 -1 1310
box -12 -8 92 272
use INVX1  _1109_
timestamp 1701862152
transform -1 0 850 0 -1 1310
box -12 -8 52 272
use INVX1  _1110_
timestamp 1701862152
transform 1 0 1070 0 -1 1310
box -12 -8 52 272
use OAI21X1  _1111_
timestamp 1702508443
transform -1 0 750 0 -1 1310
box -12 -8 92 272
use NAND3X1  _1112_
timestamp 1702508443
transform -1 0 610 0 1 790
box -12 -8 92 272
use NAND3X1  _1113_
timestamp 1702508443
transform -1 0 1270 0 -1 1310
box -12 -8 92 272
use OAI21X1  _1114_
timestamp 1702508443
transform 1 0 910 0 -1 1310
box -12 -8 92 272
use NAND3X1  _1115_
timestamp 1702508443
transform -1 0 1030 0 1 790
box -12 -8 92 272
use NAND2X1  _1116_
timestamp 1702508443
transform -1 0 2050 0 1 2870
box -12 -8 72 272
use INVX1  _1117_
timestamp 1701862152
transform 1 0 1610 0 -1 2870
box -12 -8 52 272
use AND2X2  _1118_ digital_ETRI
timestamp 1701862152
transform -1 0 2510 0 1 2350
box -12 -8 94 272
use AND2X2  _1119_
timestamp 1701862152
transform -1 0 2090 0 1 2350
box -12 -8 94 272
use NAND2X1  _1120_
timestamp 1702508443
transform -1 0 1950 0 1 2350
box -12 -8 72 272
use INVX2  _1121_
timestamp 1701862152
transform -1 0 2950 0 -1 3390
box -12 -8 52 272
use OAI21X1  _1122_
timestamp 1702508443
transform -1 0 2250 0 1 2350
box -12 -8 92 272
use NAND3X1  _1123_
timestamp 1702508443
transform -1 0 1710 0 1 2350
box -12 -8 92 272
use OAI21X1  _1124_
timestamp 1702508443
transform -1 0 1810 0 -1 2870
box -12 -8 92 272
use INVX2  _1125_
timestamp 1701862152
transform -1 0 3810 0 1 2870
box -12 -8 52 272
use OAI21X1  _1126_
timestamp 1702508443
transform -1 0 1950 0 -1 2870
box -12 -8 92 272
use NAND3X1  _1127_
timestamp 1702508443
transform -1 0 1530 0 -1 2870
box -12 -8 92 272
use AND2X2  _1128_
timestamp 1701862152
transform -1 0 1330 0 1 790
box -12 -8 94 272
use NAND3X1  _1129_
timestamp 1702508443
transform 1 0 690 0 -1 790
box -12 -8 92 272
use AOI21X1  _1130_
timestamp 1702508443
transform 1 0 1110 0 1 790
box -12 -8 92 272
use AOI21X1  _1131_
timestamp 1702508443
transform 1 0 670 0 1 790
box -12 -8 92 272
use NAND2X1  _1132_
timestamp 1702508443
transform -1 0 1470 0 1 790
box -12 -8 72 272
use OAI21X1  _1133_
timestamp 1702508443
transform -1 0 1070 0 -1 790
box -12 -8 92 272
use AOI21X1  _1134_
timestamp 1702508443
transform -1 0 930 0 -1 790
box -12 -8 92 272
use NAND3X1  _1135_
timestamp 1702508443
transform -1 0 1410 0 1 270
box -12 -8 92 272
use NAND3X1  _1136_
timestamp 1702508443
transform -1 0 1370 0 -1 790
box -12 -8 92 272
use OAI21X1  _1137_
timestamp 1702508443
transform 1 0 1150 0 -1 790
box -12 -8 92 272
use AOI22X1  _1138_
timestamp 1701862152
transform -1 0 1250 0 1 270
box -14 -8 114 272
use OAI21X1  _1139_
timestamp 1702508443
transform -1 0 850 0 -1 270
box -12 -8 92 272
use AOI21X1  _1140_
timestamp 1702508443
transform -1 0 1570 0 1 270
box -12 -8 92 272
use NAND3X1  _1141_
timestamp 1702508443
transform -1 0 1090 0 1 270
box -12 -8 92 272
use NAND3X1  _1142_
timestamp 1702508443
transform -1 0 950 0 1 270
box -12 -8 92 272
use NAND3X1  _1143_
timestamp 1702508443
transform 1 0 910 0 -1 270
box -12 -8 92 272
use NAND3X1  _1144_
timestamp 1702508443
transform 1 0 1330 0 -1 270
box -12 -8 92 272
use INVX1  _1145_
timestamp 1701862152
transform -1 0 2250 0 1 270
box -12 -8 52 272
use NAND2X1  _1146_
timestamp 1702508443
transform -1 0 1250 0 -1 270
box -12 -8 72 272
use NAND2X1  _1147_
timestamp 1702508443
transform -1 0 2130 0 1 270
box -12 -8 72 272
use AOI21X1  _1148_
timestamp 1702508443
transform 1 0 2430 0 -1 270
box -12 -8 92 272
use NAND3X1  _1149_
timestamp 1702508443
transform -1 0 2370 0 -1 270
box -12 -8 92 272
use NAND2X1  _1150_
timestamp 1702508443
transform -1 0 2850 0 -1 270
box -12 -8 72 272
use OAI21X1  _1151_
timestamp 1702508443
transform 1 0 2910 0 -1 270
box -12 -8 92 272
use NAND2X1  _1152_
timestamp 1702508443
transform 1 0 4130 0 -1 270
box -12 -8 72 272
use INVX1  _1153_
timestamp 1701862152
transform -1 0 1830 0 -1 270
box -12 -8 52 272
use OAI21X1  _1154_
timestamp 1702508443
transform -1 0 570 0 -1 270
box -12 -8 92 272
use INVX1  _1155_
timestamp 1701862152
transform 1 0 2930 0 1 3910
box -12 -8 52 272
use NOR2X1  _1156_
timestamp 1701862152
transform -1 0 2410 0 1 3910
box -12 -8 74 272
use INVX1  _1157_
timestamp 1701862152
transform 1 0 930 0 -1 2350
box -12 -8 52 272
use INVX1  _1158_
timestamp 1701862152
transform -1 0 1570 0 1 2350
box -12 -8 52 272
use OAI21X1  _1159_
timestamp 1702508443
transform -1 0 1470 0 1 2350
box -12 -8 92 272
use XOR2X1  _1160_ digital_ETRI
timestamp 1702508443
transform -1 0 1150 0 -1 2350
box -12 -8 132 272
use AOI21X1  _1161_
timestamp 1702508443
transform -1 0 450 0 1 790
box -12 -8 92 272
use NAND2X1  _1162_
timestamp 1702508443
transform -1 0 1790 0 1 2870
box -12 -8 72 272
use AND2X2  _1163_
timestamp 1701862152
transform 1 0 1850 0 1 2870
box -12 -8 94 272
use OAI21X1  _1164_
timestamp 1702508443
transform 1 0 1270 0 1 2870
box -12 -8 92 272
use AND2X2  _1165_
timestamp 1701862152
transform 1 0 1490 0 1 3390
box -12 -8 94 272
use OAI21X1  _1166_
timestamp 1702508443
transform -1 0 1650 0 1 2870
box -12 -8 92 272
use NAND3X1  _1167_
timestamp 1702508443
transform -1 0 1190 0 1 2870
box -12 -8 92 272
use INVX1  _1168_
timestamp 1701862152
transform -1 0 870 0 1 2870
box -12 -8 52 272
use NAND2X1  _1169_
timestamp 1702508443
transform -1 0 1490 0 1 2870
box -12 -8 72 272
use OAI22X1  _1170_ digital_ETRI
timestamp 1701862152
transform -1 0 1250 0 -1 2870
box -12 -8 112 272
use NAND3X1  _1171_
timestamp 1702508443
transform 1 0 950 0 1 2870
box -12 -8 92 272
use NAND2X1  _1172_
timestamp 1702508443
transform 1 0 870 0 -1 2870
box -12 -8 72 272
use OAI21X1  _1173_
timestamp 1702508443
transform -1 0 1190 0 1 1310
box -12 -8 92 272
use INVX1  _1174_
timestamp 1701862152
transform -1 0 1050 0 1 1310
box -12 -8 52 272
use NAND2X1  _1175_
timestamp 1702508443
transform 1 0 1390 0 1 1830
box -12 -8 72 272
use NAND3X1  _1176_
timestamp 1702508443
transform 1 0 1370 0 -1 2350
box -12 -8 92 272
use INVX1  _1177_
timestamp 1701862152
transform -1 0 1290 0 -1 1830
box -12 -8 52 272
use AOI21X1  _1178_
timestamp 1702508443
transform 1 0 1210 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1179_
timestamp 1702508443
transform -1 0 1170 0 -1 1830
box -12 -8 92 272
use INVX1  _1180_
timestamp 1701862152
transform -1 0 1010 0 1 1830
box -12 -8 52 272
use INVX1  _1181_
timestamp 1701862152
transform -1 0 1010 0 -1 1830
box -12 -8 52 272
use NAND3X1  _1182_
timestamp 1702508443
transform -1 0 730 0 -1 1830
box -12 -8 92 272
use NAND3X1  _1183_
timestamp 1702508443
transform -1 0 610 0 1 1310
box -12 -8 92 272
use AOI21X1  _1184_
timestamp 1702508443
transform 1 0 810 0 -1 1830
box -12 -8 92 272
use INVX1  _1185_
timestamp 1701862152
transform -1 0 1710 0 -1 2350
box -12 -8 52 272
use NAND3X1  _1186_
timestamp 1702508443
transform -1 0 1610 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1187_
timestamp 1702508443
transform -1 0 1850 0 -1 2350
box -12 -8 92 272
use AOI21X1  _1188_
timestamp 1702508443
transform -1 0 1330 0 1 1830
box -12 -8 92 272
use OAI21X1  _1189_
timestamp 1702508443
transform 1 0 850 0 1 1310
box -12 -8 92 272
use NAND3X1  _1190_
timestamp 1702508443
transform -1 0 450 0 -1 1310
box -12 -8 92 272
use AND2X2  _1191_
timestamp 1701862152
transform -1 0 790 0 -1 2870
box -12 -8 94 272
use NAND3X1  _1192_
timestamp 1702508443
transform -1 0 450 0 1 1310
box -12 -8 92 272
use OAI21X1  _1193_
timestamp 1702508443
transform -1 0 770 0 1 1310
box -12 -8 92 272
use NAND3X1  _1194_
timestamp 1702508443
transform -1 0 170 0 1 1310
box -12 -8 92 272
use NAND3X1  _1195_
timestamp 1702508443
transform 1 0 210 0 1 790
box -12 -8 92 272
use OAI21X1  _1196_
timestamp 1702508443
transform 1 0 1450 0 -1 790
box -12 -8 92 272
use AOI21X1  _1197_
timestamp 1702508443
transform 1 0 230 0 1 1310
box -12 -8 92 272
use AOI21X1  _1198_
timestamp 1702508443
transform -1 0 610 0 -1 1310
box -12 -8 92 272
use OAI21X1  _1199_
timestamp 1702508443
transform 1 0 530 0 -1 790
box -12 -8 92 272
use NAND3X1  _1200_
timestamp 1702508443
transform 1 0 190 0 -1 270
box -12 -8 92 272
use INVX1  _1201_
timestamp 1701862152
transform -1 0 130 0 -1 270
box -12 -8 52 272
use NAND3X1  _1202_
timestamp 1702508443
transform -1 0 150 0 1 790
box -12 -8 92 272
use OAI21X1  _1203_
timestamp 1702508443
transform -1 0 450 0 -1 790
box -12 -8 92 272
use NAND3X1  _1204_
timestamp 1702508443
transform 1 0 90 0 1 270
box -12 -8 92 272
use NAND3X1  _1205_
timestamp 1702508443
transform 1 0 330 0 -1 270
box -12 -8 92 272
use AOI21X1  _1206_
timestamp 1702508443
transform -1 0 790 0 1 270
box -12 -8 92 272
use AOI21X1  _1207_
timestamp 1702508443
transform 1 0 230 0 1 270
box -12 -8 92 272
use AOI21X1  _1208_
timestamp 1702508443
transform 1 0 390 0 1 270
box -12 -8 92 272
use OAI21X1  _1209_
timestamp 1702508443
transform 1 0 550 0 1 270
box -12 -8 92 272
use NAND3X1  _1210_
timestamp 1702508443
transform 1 0 1650 0 -1 270
box -12 -8 92 272
use INVX1  _1211_
timestamp 1701862152
transform 1 0 1910 0 -1 270
box -12 -8 52 272
use AND2X2  _1212_
timestamp 1701862152
transform 1 0 1050 0 -1 270
box -12 -8 94 272
use AOI22X1  _1213_
timestamp 1701862152
transform 1 0 1490 0 -1 270
box -14 -8 114 272
use NOR2X1  _1214_
timestamp 1701862152
transform -1 0 2070 0 -1 270
box -12 -8 74 272
use XOR2X1  _1215_
timestamp 1702508443
transform 1 0 2590 0 -1 270
box -12 -8 132 272
use OAI21X1  _1216_
timestamp 1702508443
transform 1 0 3730 0 -1 270
box -12 -8 92 272
use OAI21X1  _1217_
timestamp 1702508443
transform 1 0 2130 0 -1 270
box -12 -8 92 272
use INVX1  _1218_
timestamp 1701862152
transform -1 0 910 0 1 1830
box -12 -8 52 272
use NAND2X1  _1219_
timestamp 1702508443
transform 1 0 1250 0 1 2350
box -12 -8 72 272
use INVX1  _1220_
timestamp 1701862152
transform 1 0 90 0 -1 790
box -12 -8 52 272
use AOI21X1  _1221_
timestamp 1702508443
transform -1 0 290 0 -1 790
box -12 -8 92 272
use AOI22X1  _1222_
timestamp 1701862152
transform 1 0 2470 0 1 3910
box -14 -8 114 272
use AND2X2  _1223_
timestamp 1701862152
transform 1 0 1950 0 1 3910
box -12 -8 94 272
use NAND2X1  _1224_
timestamp 1702508443
transform -1 0 1550 0 1 3910
box -12 -8 72 272
use INVX1  _1225_
timestamp 1701862152
transform -1 0 970 0 -1 4430
box -12 -8 52 272
use NOR2X1  _1226_
timestamp 1701862152
transform -1 0 770 0 1 3910
box -12 -8 74 272
use NAND2X1  _1227_
timestamp 1702508443
transform 1 0 1310 0 -1 2870
box -12 -8 72 272
use OAI21X1  _1228_
timestamp 1702508443
transform -1 0 1090 0 -1 2870
box -12 -8 92 272
use XNOR2X1  _1229_ digital_ETRI
timestamp 1702508443
transform -1 0 190 0 1 3390
box -12 -8 132 272
use INVX1  _1230_
timestamp 1701862152
transform -1 0 290 0 -1 1830
box -12 -8 52 272
use AOI21X1  _1231_
timestamp 1702508443
transform 1 0 90 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1232_
timestamp 1702508443
transform -1 0 1710 0 -1 3910
box -12 -8 72 272
use NAND2X1  _1233_
timestamp 1702508443
transform -1 0 1430 0 -1 3910
box -12 -8 72 272
use NOR2X1  _1234_
timestamp 1701862152
transform 1 0 1070 0 -1 3910
box -12 -8 74 272
use AND2X2  _1235_
timestamp 1701862152
transform -1 0 1290 0 -1 3910
box -12 -8 94 272
use OAI21X1  _1236_
timestamp 1702508443
transform -1 0 1010 0 -1 3910
box -12 -8 92 272
use INVX1  _1237_
timestamp 1701862152
transform 1 0 970 0 1 3910
box -12 -8 52 272
use AND2X2  _1238_
timestamp 1701862152
transform 1 0 1630 0 1 3910
box -12 -8 94 272
use NAND2X1  _1239_
timestamp 1702508443
transform -1 0 1430 0 1 3910
box -12 -8 72 272
use OAI21X1  _1240_
timestamp 1702508443
transform -1 0 1590 0 -1 3910
box -12 -8 92 272
use NAND3X1  _1241_
timestamp 1702508443
transform -1 0 910 0 1 3910
box -12 -8 92 272
use NAND2X1  _1242_
timestamp 1702508443
transform 1 0 790 0 -1 3910
box -12 -8 72 272
use OAI21X1  _1243_
timestamp 1702508443
transform -1 0 1170 0 1 1830
box -12 -8 92 272
use INVX1  _1244_
timestamp 1701862152
transform 1 0 930 0 -1 3390
box -12 -8 52 272
use NAND2X1  _1245_
timestamp 1702508443
transform -1 0 1710 0 1 3390
box -12 -8 72 272
use NAND3X1  _1246_
timestamp 1702508443
transform -1 0 1630 0 -1 3390
box -12 -8 92 272
use INVX1  _1247_
timestamp 1701862152
transform 1 0 1090 0 1 3390
box -12 -8 52 272
use AOI21X1  _1248_
timestamp 1702508443
transform -1 0 1790 0 -1 3390
box -12 -8 92 272
use OAI21X1  _1249_
timestamp 1702508443
transform 1 0 1190 0 1 3390
box -12 -8 92 272
use INVX1  _1250_
timestamp 1701862152
transform -1 0 1490 0 -1 3390
box -12 -8 52 272
use INVX1  _1251_
timestamp 1701862152
transform -1 0 1370 0 -1 3390
box -12 -8 52 272
use NAND3X1  _1252_
timestamp 1702508443
transform -1 0 1130 0 -1 3390
box -12 -8 92 272
use NAND3X1  _1253_
timestamp 1702508443
transform -1 0 1010 0 1 3390
box -12 -8 92 272
use AOI21X1  _1254_
timestamp 1702508443
transform -1 0 1270 0 -1 3390
box -12 -8 92 272
use INVX1  _1255_
timestamp 1701862152
transform -1 0 2450 0 -1 3390
box -12 -8 52 272
use NAND3X1  _1256_
timestamp 1702508443
transform -1 0 2330 0 -1 3390
box -12 -8 92 272
use OAI21X1  _1257_
timestamp 1702508443
transform -1 0 2850 0 -1 3390
box -12 -8 92 272
use AOI21X1  _1258_
timestamp 1702508443
transform -1 0 2190 0 -1 3390
box -12 -8 92 272
use OAI21X1  _1259_
timestamp 1702508443
transform -1 0 710 0 -1 3390
box -12 -8 92 272
use NAND3X1  _1260_
timestamp 1702508443
transform -1 0 470 0 1 2870
box -12 -8 92 272
use AND2X2  _1261_
timestamp 1701862152
transform -1 0 710 0 -1 3910
box -12 -8 94 272
use NAND3X1  _1262_
timestamp 1702508443
transform 1 0 770 0 1 3390
box -12 -8 92 272
use OAI21X1  _1263_
timestamp 1702508443
transform 1 0 790 0 -1 3390
box -12 -8 92 272
use NAND3X1  _1264_
timestamp 1702508443
transform -1 0 410 0 -1 3390
box -12 -8 92 272
use NAND3X1  _1265_
timestamp 1702508443
transform -1 0 170 0 -1 2870
box -12 -8 92 272
use AOI21X1  _1266_
timestamp 1702508443
transform -1 0 590 0 -1 1830
box -12 -8 92 272
use OAI21X1  _1267_
timestamp 1702508443
transform -1 0 450 0 -1 1830
box -12 -8 92 272
use AOI21X1  _1268_
timestamp 1702508443
transform 1 0 490 0 -1 3390
box -12 -8 92 272
use AOI21X1  _1269_
timestamp 1702508443
transform -1 0 610 0 1 2870
box -12 -8 92 272
use OAI21X1  _1270_
timestamp 1702508443
transform -1 0 470 0 -1 2870
box -12 -8 92 272
use NAND3X1  _1271_
timestamp 1702508443
transform 1 0 230 0 1 2350
box -12 -8 92 272
use XOR2X1  _1272_
timestamp 1702508443
transform 1 0 270 0 1 3390
box -12 -8 132 272
use NAND3X1  _1273_
timestamp 1702508443
transform 1 0 230 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1274_
timestamp 1702508443
transform 1 0 550 0 -1 2870
box -12 -8 92 272
use NAND3X1  _1275_
timestamp 1702508443
transform 1 0 550 0 1 2350
box -12 -8 92 272
use NAND3X1  _1276_
timestamp 1702508443
transform -1 0 310 0 -1 2350
box -12 -8 92 272
use AOI21X1  _1277_
timestamp 1702508443
transform 1 0 90 0 -1 1310
box -12 -8 92 272
use OAI21X1  _1278_
timestamp 1702508443
transform -1 0 310 0 -1 1310
box -12 -8 92 272
use AOI21X1  _1279_
timestamp 1702508443
transform -1 0 470 0 1 2350
box -12 -8 92 272
use AOI21X1  _1280_
timestamp 1702508443
transform -1 0 170 0 1 2350
box -12 -8 92 272
use OAI21X1  _1281_
timestamp 1702508443
transform 1 0 70 0 1 1830
box -12 -8 92 272
use NAND3X1  _1282_
timestamp 1702508443
transform 1 0 230 0 1 1830
box -12 -8 92 272
use INVX1  _1283_
timestamp 1701862152
transform -1 0 850 0 -1 2350
box -12 -8 52 272
use NAND3X1  _1284_
timestamp 1702508443
transform 1 0 390 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1285_
timestamp 1702508443
transform 1 0 90 0 -1 2350
box -12 -8 92 272
use NAND3X1  _1286_
timestamp 1702508443
transform 1 0 670 0 -1 2350
box -12 -8 92 272
use NAND3X1  _1287_
timestamp 1702508443
transform -1 0 790 0 1 1830
box -12 -8 92 272
use AOI21X1  _1288_
timestamp 1702508443
transform 1 0 530 0 -1 2350
box -12 -8 92 272
use AOI21X1  _1289_
timestamp 1702508443
transform 1 0 390 0 1 1830
box -12 -8 92 272
use OAI21X1  _1290_
timestamp 1702508443
transform 1 0 550 0 1 1830
box -12 -8 92 272
use AOI21X1  _1291_
timestamp 1702508443
transform 1 0 2390 0 1 790
box -12 -8 92 272
use NAND3X1  _1292_
timestamp 1702508443
transform 1 0 2250 0 1 790
box -12 -8 92 272
use NAND2X1  _1293_
timestamp 1702508443
transform -1 0 3010 0 1 790
box -12 -8 72 272
use OAI22X1  _1294_
timestamp 1701862152
transform -1 0 3190 0 1 790
box -12 -8 112 272
use INVX1  _1295_
timestamp 1701862152
transform 1 0 2750 0 -1 1310
box -12 -8 52 272
use INVX1  _1296_
timestamp 1701862152
transform -1 0 3010 0 -1 1310
box -12 -8 52 272
use INVX1  _1297_
timestamp 1701862152
transform -1 0 1190 0 1 2350
box -12 -8 52 272
use AOI21X1  _1298_
timestamp 1702508443
transform 1 0 830 0 1 2350
box -12 -8 92 272
use NAND2X1  _1299_
timestamp 1702508443
transform 1 0 90 0 -1 3910
box -12 -8 72 272
use INVX1  _1300_
timestamp 1701862152
transform 1 0 90 0 -1 3390
box -12 -8 52 272
use AOI21X1  _1301_
timestamp 1702508443
transform -1 0 270 0 -1 3390
box -12 -8 92 272
use NAND2X1  _1302_
timestamp 1702508443
transform 1 0 2970 0 -1 4430
box -12 -8 72 272
use INVX1  _1303_
timestamp 1701862152
transform -1 0 2450 0 -1 4430
box -12 -8 52 272
use AND2X2  _1304_
timestamp 1701862152
transform -1 0 2730 0 -1 4430
box -12 -8 94 272
use NAND2X1  _1305_
timestamp 1702508443
transform 1 0 2090 0 1 3910
box -12 -8 72 272
use NAND2X1  _1306_
timestamp 1702508443
transform 1 0 1990 0 1 4430
box -12 -8 72 272
use OAI21X1  _1307_
timestamp 1702508443
transform -1 0 2350 0 -1 4430
box -12 -8 92 272
use AOI21X1  _1308_
timestamp 1702508443
transform -1 0 2030 0 -1 4430
box -12 -8 92 272
use INVX1  _1309_
timestamp 1701862152
transform 1 0 3190 0 1 3910
box -12 -8 52 272
use OAI21X1  _1310_
timestamp 1702508443
transform -1 0 2710 0 1 3910
box -12 -8 92 272
use OAI21X1  _1311_
timestamp 1702508443
transform -1 0 1870 0 1 3910
box -12 -8 92 272
use AOI21X1  _1312_
timestamp 1702508443
transform -1 0 1750 0 -1 4430
box -12 -8 92 272
use OAI21X1  _1313_
timestamp 1702508443
transform 1 0 1230 0 1 3910
box -12 -8 92 272
use OAI21X1  _1314_
timestamp 1702508443
transform -1 0 1590 0 -1 4430
box -12 -8 92 272
use NAND3X1  _1315_
timestamp 1702508443
transform -1 0 1890 0 -1 4430
box -12 -8 92 272
use NAND3X1  _1316_
timestamp 1702508443
transform -1 0 2190 0 -1 4430
box -12 -8 92 272
use AOI21X1  _1317_
timestamp 1702508443
transform 1 0 1090 0 1 3910
box -12 -8 92 272
use NAND3X1  _1318_
timestamp 1702508443
transform -1 0 1270 0 -1 4430
box -12 -8 92 272
use NAND3X1  _1319_
timestamp 1702508443
transform -1 0 1130 0 -1 4430
box -12 -8 92 272
use NAND3X1  _1320_
timestamp 1702508443
transform -1 0 1330 0 1 4430
box -12 -8 92 272
use OAI21X1  _1321_
timestamp 1702508443
transform -1 0 1430 0 -1 4430
box -12 -8 92 272
use NAND3X1  _1322_
timestamp 1702508443
transform 1 0 850 0 1 4430
box -12 -8 92 272
use NAND2X1  _1323_
timestamp 1702508443
transform 1 0 670 0 -1 4950
box -12 -8 72 272
use INVX1  _1324_
timestamp 1701862152
transform -1 0 410 0 -1 3910
box -12 -8 52 272
use AOI21X1  _1325_
timestamp 1702508443
transform -1 0 290 0 -1 3910
box -12 -8 92 272
use NAND2X1  _1326_
timestamp 1702508443
transform 1 0 1550 0 1 4430
box -12 -8 72 272
use NAND2X1  _1327_
timestamp 1702508443
transform -1 0 1470 0 1 4430
box -12 -8 72 272
use NAND3X1  _1328_
timestamp 1702508443
transform 1 0 1070 0 -1 4950
box -12 -8 92 272
use NAND2X1  _1329_
timestamp 1702508443
transform 1 0 1130 0 1 4430
box -12 -8 72 272
use NAND2X1  _1330_
timestamp 1702508443
transform 1 0 1370 0 -1 4950
box -12 -8 72 272
use NAND3X1  _1331_
timestamp 1702508443
transform 1 0 1230 0 -1 4950
box -12 -8 92 272
use INVX1  _1332_
timestamp 1701862152
transform 1 0 1790 0 -1 4950
box -12 -8 52 272
use AND2X2  _1333_
timestamp 1701862152
transform 1 0 2770 0 -1 4950
box -12 -8 94 272
use NAND2X1  _1334_
timestamp 1702508443
transform 1 0 2050 0 -1 4950
box -12 -8 72 272
use OAI21X1  _1335_
timestamp 1702508443
transform -1 0 1750 0 1 4430
box -12 -8 92 272
use NAND3X1  _1336_
timestamp 1702508443
transform -1 0 1830 0 1 4950
box -12 -8 92 272
use NAND2X1  _1337_
timestamp 1702508443
transform 1 0 1370 0 1 4950
box -12 -8 72 272
use OAI21X1  _1338_
timestamp 1702508443
transform 1 0 1350 0 1 3390
box -12 -8 92 272
use INVX1  _1339_
timestamp 1701862152
transform -1 0 850 0 1 5470
box -12 -8 52 272
use NAND2X1  _1340_
timestamp 1702508443
transform 1 0 1490 0 1 4950
box -12 -8 72 272
use INVX1  _1341_
timestamp 1701862152
transform 1 0 1630 0 1 4950
box -12 -8 52 272
use NAND3X1  _1342_
timestamp 1702508443
transform -1 0 1770 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1343_
timestamp 1702508443
transform -1 0 1910 0 -1 5470
box -12 -8 72 272
use NAND2X1  _1344_
timestamp 1702508443
transform 1 0 1570 0 -1 5470
box -12 -8 72 272
use NAND3X1  _1345_
timestamp 1702508443
transform -1 0 1590 0 1 5470
box -12 -8 92 272
use INVX1  _1346_
timestamp 1701862152
transform 1 0 1970 0 1 5470
box -12 -8 52 272
use NAND3X1  _1347_
timestamp 1702508443
transform -1 0 2210 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1348_
timestamp 1702508443
transform -1 0 1730 0 1 5470
box -12 -8 72 272
use NAND3X1  _1349_
timestamp 1702508443
transform -1 0 1790 0 -1 5990
box -12 -8 92 272
use NAND3X1  _1350_
timestamp 1702508443
transform -1 0 990 0 1 5470
box -12 -8 92 272
use AOI21X1  _1351_
timestamp 1702508443
transform 1 0 1810 0 1 5470
box -12 -8 92 272
use AOI21X1  _1352_
timestamp 1702508443
transform -1 0 1490 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1353_
timestamp 1702508443
transform -1 0 1350 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1354_
timestamp 1702508443
transform -1 0 1050 0 -1 5470
box -12 -8 92 272
use AND2X2  _1355_
timestamp 1701862152
transform -1 0 1310 0 1 4950
box -12 -8 94 272
use NAND3X1  _1356_
timestamp 1702508443
transform -1 0 1150 0 1 5470
box -12 -8 92 272
use OAI21X1  _1357_
timestamp 1702508443
transform -1 0 1190 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1358_
timestamp 1702508443
transform -1 0 770 0 1 4950
box -12 -8 92 272
use NAND3X1  _1359_
timestamp 1702508443
transform -1 0 470 0 1 4950
box -12 -8 92 272
use AOI21X1  _1360_
timestamp 1702508443
transform -1 0 690 0 1 3390
box -12 -8 92 272
use OAI21X1  _1361_
timestamp 1702508443
transform -1 0 570 0 -1 3910
box -12 -8 92 272
use AOI21X1  _1362_
timestamp 1702508443
transform -1 0 910 0 1 4950
box -12 -8 92 272
use AOI21X1  _1363_
timestamp 1702508443
transform -1 0 890 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1364_
timestamp 1702508443
transform -1 0 610 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1365_
timestamp 1702508443
transform 1 0 230 0 -1 4950
box -12 -8 92 272
use AND2X2  _1366_
timestamp 1701862152
transform -1 0 1010 0 -1 4950
box -12 -8 94 272
use NAND3X1  _1367_
timestamp 1702508443
transform -1 0 610 0 1 4950
box -12 -8 92 272
use OAI21X1  _1368_
timestamp 1702508443
transform -1 0 470 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1369_
timestamp 1702508443
transform 1 0 230 0 1 4950
box -12 -8 92 272
use NAND3X1  _1370_
timestamp 1702508443
transform -1 0 310 0 -1 4430
box -12 -8 92 272
use AOI21X1  _1371_
timestamp 1702508443
transform -1 0 310 0 1 2870
box -12 -8 92 272
use OAI21X1  _1372_
timestamp 1702508443
transform 1 0 70 0 1 2870
box -12 -8 92 272
use AOI21X1  _1373_
timestamp 1702508443
transform -1 0 170 0 1 4950
box -12 -8 92 272
use AOI21X1  _1374_
timestamp 1702508443
transform 1 0 70 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1375_
timestamp 1702508443
transform 1 0 90 0 1 4430
box -12 -8 92 272
use AOI21X1  _1376_
timestamp 1702508443
transform 1 0 250 0 1 3910
box -12 -8 92 272
use INVX1  _1377_
timestamp 1701862152
transform 1 0 530 0 -1 4430
box -12 -8 52 272
use NAND3X1  _1378_
timestamp 1702508443
transform 1 0 390 0 -1 4430
box -12 -8 92 272
use OAI21X1  _1379_
timestamp 1702508443
transform 1 0 70 0 -1 4430
box -12 -8 92 272
use AOI21X1  _1380_
timestamp 1702508443
transform 1 0 550 0 1 3910
box -12 -8 92 272
use OAI21X1  _1381_
timestamp 1702508443
transform 1 0 690 0 1 2870
box -12 -8 92 272
use AOI21X1  _1382_
timestamp 1702508443
transform 1 0 690 0 1 2350
box -12 -8 92 272
use OAI21X1  _1383_
timestamp 1702508443
transform 1 0 990 0 1 2350
box -12 -8 92 272
use NAND3X1  _1384_
timestamp 1702508443
transform -1 0 470 0 1 3910
box -12 -8 92 272
use NAND3X1  _1385_
timestamp 1702508443
transform 1 0 90 0 1 3910
box -12 -8 92 272
use NAND3X1  _1386_
timestamp 1702508443
transform -1 0 550 0 1 3390
box -12 -8 92 272
use NAND2X1  _1387_
timestamp 1702508443
transform 1 0 2210 0 -1 2350
box -12 -8 72 272
use OAI21X1  _1388_
timestamp 1702508443
transform 1 0 3210 0 -1 1310
box -12 -8 92 272
use NOR2X1  _1389_
timestamp 1701862152
transform -1 0 3130 0 -1 1310
box -12 -8 74 272
use INVX1  _1390_
timestamp 1701862152
transform 1 0 3310 0 1 1310
box -12 -8 52 272
use AOI21X1  _1391_
timestamp 1702508443
transform 1 0 3350 0 -1 1310
box -12 -8 92 272
use AOI22X1  _1392_
timestamp 1701862152
transform -1 0 3610 0 -1 1310
box -14 -8 114 272
use NAND2X1  _1393_
timestamp 1702508443
transform -1 0 4650 0 1 1830
box -12 -8 72 272
use INVX1  _1394_
timestamp 1701862152
transform -1 0 2370 0 -1 2350
box -12 -8 52 272
use AND2X2  _1395_
timestamp 1701862152
transform 1 0 2070 0 -1 2350
box -12 -8 94 272
use OAI22X1  _1396_
timestamp 1701862152
transform 1 0 2430 0 -1 2350
box -12 -8 112 272
use AOI21X1  _1397_
timestamp 1702508443
transform 1 0 250 0 1 4430
box -12 -8 92 272
use OAI21X1  _1398_
timestamp 1702508443
transform 1 0 410 0 1 4430
box -12 -8 92 272
use NAND2X1  _1399_
timestamp 1702508443
transform -1 0 850 0 -1 4950
box -12 -8 72 272
use INVX1  _1400_
timestamp 1701862152
transform 1 0 90 0 1 5470
box -12 -8 52 272
use INVX1  _1401_
timestamp 1701862152
transform 1 0 70 0 -1 5470
box -12 -8 52 272
use AOI21X1  _1402_
timestamp 1702508443
transform 1 0 190 0 -1 5470
box -12 -8 92 272
use AND2X2  _1403_
timestamp 1701862152
transform 1 0 1830 0 1 4430
box -12 -8 94 272
use NAND2X1  _1404_
timestamp 1702508443
transform 1 0 2830 0 1 4430
box -12 -8 72 272
use INVX1  _1405_
timestamp 1701862152
transform 1 0 2590 0 1 4430
box -12 -8 52 272
use AND2X2  _1406_
timestamp 1701862152
transform -1 0 3110 0 1 3910
box -12 -8 94 272
use AND2X2  _1407_
timestamp 1701862152
transform -1 0 3730 0 -1 4430
box -12 -8 94 272
use NAND2X1  _1408_
timestamp 1702508443
transform 1 0 3110 0 -1 4430
box -12 -8 72 272
use NAND2X1  _1409_
timestamp 1702508443
transform -1 0 3450 0 -1 4430
box -12 -8 72 272
use OAI21X1  _1410_
timestamp 1702508443
transform 1 0 3250 0 -1 4430
box -12 -8 92 272
use AOI21X1  _1411_
timestamp 1702508443
transform -1 0 2550 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1412_
timestamp 1702508443
transform 1 0 2810 0 -1 4430
box -12 -8 92 272
use OAI21X1  _1413_
timestamp 1702508443
transform 1 0 2790 0 1 3910
box -12 -8 92 272
use AOI21X1  _1414_
timestamp 1702508443
transform -1 0 2350 0 1 4430
box -12 -8 92 272
use AND2X2  _1415_
timestamp 1701862152
transform 1 0 1510 0 -1 4950
box -12 -8 94 272
use OAI21X1  _1416_
timestamp 1702508443
transform 1 0 1890 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1417_
timestamp 1702508443
transform -1 0 2270 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1418_
timestamp 1702508443
transform 1 0 2430 0 1 4430
box -12 -8 92 272
use NAND3X1  _1419_
timestamp 1702508443
transform 1 0 2610 0 -1 4950
box -12 -8 92 272
use NOR2X1  _1420_
timestamp 1701862152
transform -1 0 1730 0 -1 4950
box -12 -8 74 272
use AOI21X1  _1421_
timestamp 1702508443
transform 1 0 1890 0 1 4950
box -12 -8 92 272
use NAND3X1  _1422_
timestamp 1702508443
transform -1 0 2570 0 1 4950
box -12 -8 92 272
use NAND3X1  _1423_
timestamp 1702508443
transform 1 0 2030 0 1 4950
box -12 -8 92 272
use INVX1  _1424_
timestamp 1701862152
transform -1 0 2570 0 -1 4430
box -12 -8 52 272
use OAI21X1  _1425_
timestamp 1702508443
transform -1 0 2210 0 1 4430
box -12 -8 92 272
use NAND3X1  _1426_
timestamp 1702508443
transform -1 0 2410 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1427_
timestamp 1702508443
transform -1 0 2410 0 1 4950
box -12 -8 92 272
use NAND3X1  _1428_
timestamp 1702508443
transform 1 0 2170 0 1 4950
box -12 -8 92 272
use NAND2X1  _1429_
timestamp 1702508443
transform -1 0 1630 0 -1 5990
box -12 -8 72 272
use INVX1  _1430_
timestamp 1701862152
transform -1 0 1170 0 1 4950
box -12 -8 52 272
use AOI21X1  _1431_
timestamp 1702508443
transform -1 0 1050 0 1 4950
box -12 -8 92 272
use NAND2X1  _1432_
timestamp 1702508443
transform 1 0 3110 0 1 4430
box -12 -8 72 272
use NAND2X1  _1433_
timestamp 1702508443
transform 1 0 3350 0 1 4430
box -12 -8 72 272
use NAND3X1  _1434_
timestamp 1702508443
transform -1 0 3170 0 -1 4950
box -12 -8 92 272
use NAND2X1  _1435_
timestamp 1702508443
transform 1 0 3490 0 1 4430
box -12 -8 72 272
use NAND3X1  _1436_
timestamp 1702508443
transform -1 0 3030 0 1 4430
box -12 -8 92 272
use NAND3X1  _1437_
timestamp 1702508443
transform -1 0 3010 0 -1 4950
box -12 -8 92 272
use INVX1  _1438_
timestamp 1701862152
transform -1 0 3130 0 1 4950
box -12 -8 52 272
use AND2X2  _1439_
timestamp 1701862152
transform 1 0 3810 0 -1 4430
box -12 -8 94 272
use NAND2X1  _1440_
timestamp 1702508443
transform 1 0 3550 0 1 4950
box -12 -8 72 272
use OAI21X1  _1441_
timestamp 1702508443
transform -1 0 3470 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1442_
timestamp 1702508443
transform -1 0 3030 0 1 4950
box -12 -8 92 272
use NAND2X1  _1443_
timestamp 1702508443
transform 1 0 2710 0 -1 5470
box -12 -8 72 272
use AOI21X1  _1444_
timestamp 1702508443
transform 1 0 2570 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1445_
timestamp 1702508443
transform 1 0 2410 0 -1 5470
box -12 -8 92 272
use INVX1  _1446_
timestamp 1701862152
transform -1 0 4330 0 1 5470
box -12 -8 52 272
use NOR2X1  _1447_
timestamp 1701862152
transform 1 0 2630 0 1 5470
box -12 -8 74 272
use NAND3X1  _1448_
timestamp 1702508443
transform 1 0 1990 0 -1 5990
box -12 -8 92 272
use AOI21X1  _1449_
timestamp 1702508443
transform 1 0 1990 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1450_
timestamp 1702508443
transform 1 0 2070 0 1 5470
box -12 -8 92 272
use OAI21X1  _1451_
timestamp 1702508443
transform -1 0 2550 0 1 5470
box -12 -8 92 272
use NAND3X1  _1452_
timestamp 1702508443
transform -1 0 2230 0 -1 5990
box -12 -8 92 272
use AND2X2  _1453_
timestamp 1701862152
transform -1 0 2830 0 1 5470
box -12 -8 94 272
use INVX1  _1454_
timestamp 1701862152
transform -1 0 2390 0 1 5470
box -12 -8 52 272
use NAND2X1  _1455_
timestamp 1702508443
transform 1 0 2210 0 1 5470
box -12 -8 72 272
use NOR2X1  _1456_
timestamp 1701862152
transform 1 0 1710 0 1 5990
box -12 -8 74 272
use INVX1  _1457_
timestamp 1701862152
transform -1 0 1470 0 1 5990
box -12 -8 52 272
use OAI21X1  _1458_
timestamp 1702508443
transform -1 0 1350 0 1 5990
box -12 -8 92 272
use NAND3X1  _1459_
timestamp 1702508443
transform -1 0 890 0 -1 5990
box -12 -8 92 272
use AOI21X1  _1460_
timestamp 1702508443
transform -1 0 1450 0 1 5470
box -12 -8 92 272
use OAI21X1  _1461_
timestamp 1702508443
transform -1 0 1310 0 1 5470
box -12 -8 92 272
use NAND2X1  _1462_
timestamp 1702508443
transform -1 0 2510 0 -1 5990
box -12 -8 72 272
use NAND3X1  _1463_
timestamp 1702508443
transform 1 0 1830 0 1 5990
box -12 -8 92 272
use AOI21X1  _1464_
timestamp 1702508443
transform -1 0 1630 0 1 5990
box -12 -8 92 272
use AOI21X1  _1465_
timestamp 1702508443
transform 1 0 2290 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1466_
timestamp 1702508443
transform -1 0 810 0 1 5990
box -12 -8 92 272
use NAND3X1  _1467_
timestamp 1702508443
transform -1 0 490 0 1 5990
box -12 -8 92 272
use AND2X2  _1468_
timestamp 1701862152
transform -1 0 1490 0 -1 5990
box -12 -8 94 272
use NAND3X1  _1469_
timestamp 1702508443
transform 1 0 970 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1470_
timestamp 1702508443
transform -1 0 950 0 1 5990
box -12 -8 92 272
use NAND3X1  _1471_
timestamp 1702508443
transform -1 0 650 0 1 5990
box -12 -8 92 272
use NAND3X1  _1472_
timestamp 1702508443
transform 1 0 250 0 1 5990
box -12 -8 92 272
use AOI21X1  _1473_
timestamp 1702508443
transform -1 0 570 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1474_
timestamp 1702508443
transform -1 0 430 0 -1 5470
box -12 -8 92 272
use AOI21X1  _1475_
timestamp 1702508443
transform -1 0 610 0 -1 5990
box -12 -8 92 272
use AOI21X1  _1476_
timestamp 1702508443
transform -1 0 470 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1477_
timestamp 1702508443
transform -1 0 170 0 -1 5990
box -12 -8 92 272
use NAND3X1  _1478_
timestamp 1702508443
transform 1 0 190 0 1 5470
box -12 -8 92 272
use NAND3X1  _1479_
timestamp 1702508443
transform -1 0 170 0 1 5990
box -12 -8 92 272
use OAI21X1  _1480_
timestamp 1702508443
transform 1 0 230 0 -1 5990
box -12 -8 92 272
use NAND3X1  _1481_
timestamp 1702508443
transform -1 0 730 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1482_
timestamp 1702508443
transform 1 0 550 0 1 4430
box -12 -8 92 272
use INVX1  _1483_
timestamp 1701862152
transform -1 0 850 0 -1 4430
box -12 -8 52 272
use AOI21X1  _1484_
timestamp 1702508443
transform 1 0 650 0 -1 4430
box -12 -8 92 272
use AOI21X1  _1485_
timestamp 1702508443
transform -1 0 570 0 1 5470
box -12 -8 92 272
use AOI21X1  _1486_
timestamp 1702508443
transform 1 0 350 0 1 5470
box -12 -8 92 272
use OAI21X1  _1487_
timestamp 1702508443
transform 1 0 690 0 1 4430
box -12 -8 92 272
use NAND2X1  _1488_
timestamp 1702508443
transform -1 0 3230 0 -1 3390
box -12 -8 72 272
use XOR2X1  _1489_
timestamp 1702508443
transform -1 0 4010 0 1 2870
box -12 -8 132 272
use OAI21X1  _1490_
timestamp 1702508443
transform 1 0 4430 0 1 1830
box -12 -8 92 272
use INVX1  _1491_
timestamp 1701862152
transform 1 0 3310 0 -1 3390
box -12 -8 52 272
use AOI21X1  _1492_
timestamp 1702508443
transform 1 0 3410 0 -1 3390
box -12 -8 92 272
use INVX1  _1493_
timestamp 1701862152
transform -1 0 730 0 -1 5990
box -12 -8 52 272
use AOI21X1  _1494_
timestamp 1702508443
transform 1 0 650 0 1 5470
box -12 -8 92 272
use NAND2X1  _1495_
timestamp 1702508443
transform -1 0 2330 0 -1 5470
box -12 -8 72 272
use INVX1  _1496_
timestamp 1701862152
transform 1 0 2890 0 -1 5990
box -12 -8 52 272
use INVX1  _1497_
timestamp 1701862152
transform -1 0 1210 0 1 5990
box -12 -8 52 272
use AOI21X1  _1498_
timestamp 1702508443
transform 1 0 1030 0 1 5990
box -12 -8 92 272
use AND2X2  _1499_
timestamp 1701862152
transform 1 0 2790 0 1 4950
box -12 -8 94 272
use NAND2X1  _1500_
timestamp 1702508443
transform -1 0 3570 0 -1 4430
box -12 -8 72 272
use NAND2X1  _1501_
timestamp 1702508443
transform -1 0 3930 0 1 4430
box -12 -8 72 272
use NOR2X1  _1502_
timestamp 1701862152
transform 1 0 3730 0 1 4430
box -12 -8 74 272
use AOI22X1  _1503_
timestamp 1701862152
transform -1 0 4110 0 1 4430
box -14 -8 114 272
use NOR3X1  _1504_
timestamp 1701862152
transform -1 0 3850 0 1 4950
box -12 -8 172 272
use INVX1  _1505_
timestamp 1701862152
transform -1 0 3570 0 -1 4950
box -12 -8 52 272
use AND2X2  _1506_
timestamp 1701862152
transform -1 0 5010 0 -1 4430
box -12 -8 94 272
use NAND2X1  _1507_
timestamp 1702508443
transform 1 0 3950 0 -1 4430
box -12 -8 72 272
use INVX1  _1508_
timestamp 1701862152
transform -1 0 3970 0 1 4950
box -12 -8 52 272
use AOI21X1  _1509_
timestamp 1702508443
transform -1 0 3670 0 -1 5470
box -12 -8 92 272
use AND2X2  _1510_
timestamp 1701862152
transform -1 0 3330 0 -1 4950
box -12 -8 94 272
use OAI21X1  _1511_
timestamp 1702508443
transform 1 0 3210 0 1 4950
box -12 -8 92 272
use OAI21X1  _1512_
timestamp 1702508443
transform -1 0 3370 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1513_
timestamp 1702508443
transform 1 0 3750 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1514_
timestamp 1702508443
transform -1 0 3710 0 -1 4950
box -12 -8 92 272
use AOI22X1  _1515_
timestamp 1701862152
transform -1 0 3470 0 1 4950
box -14 -8 114 272
use NAND3X1  _1516_
timestamp 1702508443
transform -1 0 3070 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1517_
timestamp 1702508443
transform 1 0 2830 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1518_
timestamp 1702508443
transform -1 0 2770 0 1 4430
box -12 -8 72 272
use OAI21X1  _1519_
timestamp 1702508443
transform 1 0 2630 0 1 4950
box -12 -8 92 272
use NAND3X1  _1520_
timestamp 1702508443
transform 1 0 3150 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1521_
timestamp 1702508443
transform -1 0 3530 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1522_
timestamp 1702508443
transform 1 0 3530 0 1 5470
box -12 -8 92 272
use NAND2X1  _1523_
timestamp 1702508443
transform 1 0 3290 0 1 5990
box -12 -8 72 272
use AOI21X1  _1524_
timestamp 1702508443
transform 1 0 1850 0 -1 5990
box -12 -8 92 272
use AOI21X1  _1525_
timestamp 1702508443
transform 1 0 1990 0 1 5990
box -12 -8 92 272
use NAND2X1  _1526_
timestamp 1702508443
transform 1 0 4190 0 1 4430
box -12 -8 72 272
use AND2X2  _1527_
timestamp 1701862152
transform -1 0 4490 0 -1 4950
box -12 -8 94 272
use OAI21X1  _1528_
timestamp 1702508443
transform 1 0 4270 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1529_
timestamp 1702508443
transform 1 0 3950 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1530_
timestamp 1702508443
transform -1 0 4190 0 -1 4950
box -12 -8 92 272
use INVX1  _1531_
timestamp 1701862152
transform 1 0 4350 0 1 4950
box -12 -8 52 272
use NAND2X1  _1532_
timestamp 1702508443
transform -1 0 4810 0 1 4950
box -12 -8 72 272
use OAI22X1  _1533_
timestamp 1701862152
transform 1 0 3790 0 -1 4950
box -12 -8 112 272
use NAND3X1  _1534_
timestamp 1702508443
transform -1 0 4270 0 1 4950
box -12 -8 92 272
use NAND2X1  _1535_
timestamp 1702508443
transform -1 0 4110 0 -1 5470
box -12 -8 72 272
use XNOR2X1  _1536_
timestamp 1702508443
transform -1 0 4310 0 -1 5470
box -12 -8 132 272
use INVX1  _1537_
timestamp 1701862152
transform -1 0 4230 0 1 5470
box -12 -8 52 272
use NAND2X1  _1538_
timestamp 1702508443
transform -1 0 4130 0 1 5470
box -12 -8 72 272
use NAND3X1  _1539_
timestamp 1702508443
transform -1 0 3970 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1540_
timestamp 1702508443
transform -1 0 3890 0 1 5990
box -12 -8 72 272
use NOR2X1  _1541_
timestamp 1701862152
transform 1 0 3690 0 1 5990
box -12 -8 74 272
use NOR2X1  _1542_
timestamp 1701862152
transform 1 0 2590 0 -1 5990
box -12 -8 74 272
use OAI21X1  _1543_
timestamp 1702508443
transform 1 0 2730 0 -1 5990
box -12 -8 92 272
use AOI21X1  _1544_
timestamp 1702508443
transform 1 0 4390 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1545_
timestamp 1702508443
transform -1 0 4330 0 -1 5990
box -12 -8 92 272
use AND2X2  _1546_
timestamp 1701862152
transform 1 0 3950 0 1 5990
box -12 -8 94 272
use NAND3X1  _1547_
timestamp 1702508443
transform 1 0 4550 0 -1 5990
box -12 -8 92 272
use NAND2X1  _1548_
timestamp 1702508443
transform -1 0 3490 0 1 5990
box -12 -8 72 272
use NAND3X1  _1549_
timestamp 1702508443
transform -1 0 4170 0 -1 5990
box -12 -8 92 272
use NAND3X1  _1550_
timestamp 1702508443
transform -1 0 3390 0 -1 5990
box -12 -8 92 272
use AOI21X1  _1551_
timestamp 1702508443
transform 1 0 1110 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1552_
timestamp 1702508443
transform -1 0 1350 0 -1 5990
box -12 -8 92 272
use AOI22X1  _1553_
timestamp 1701862152
transform 1 0 3930 0 -1 5990
box -14 -8 114 272
use NAND3X1  _1554_
timestamp 1702508443
transform -1 0 3630 0 1 5990
box -12 -8 92 272
use OAI21X1  _1555_
timestamp 1702508443
transform 1 0 2290 0 1 5990
box -12 -8 92 272
use AOI21X1  _1556_
timestamp 1702508443
transform -1 0 3210 0 1 5990
box -12 -8 92 272
use OAI21X1  _1557_
timestamp 1702508443
transform 1 0 2990 0 1 5990
box -12 -8 92 272
use AOI21X1  _1558_
timestamp 1702508443
transform 1 0 3150 0 -1 5990
box -12 -8 92 272
use NAND3X1  _1559_
timestamp 1702508443
transform 1 0 3450 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1560_
timestamp 1702508443
transform 1 0 2690 0 1 5990
box -12 -8 92 272
use AOI21X1  _1561_
timestamp 1702508443
transform -1 0 3470 0 1 5470
box -12 -8 92 272
use OAI21X1  _1562_
timestamp 1702508443
transform -1 0 3330 0 1 5470
box -12 -8 92 272
use AOI21X1  _1563_
timestamp 1702508443
transform -1 0 3170 0 1 5470
box -12 -8 92 272
use AOI21X1  _1564_
timestamp 1702508443
transform -1 0 3070 0 -1 5990
box -12 -8 92 272
use OAI22X1  _1565_
timestamp 1701862152
transform -1 0 3010 0 1 5470
box -12 -8 112 272
use NAND2X1  _1566_
timestamp 1702508443
transform -1 0 3290 0 1 4430
box -12 -8 72 272
use XNOR2X1  _1567_
timestamp 1702508443
transform 1 0 3570 0 -1 3390
box -12 -8 132 272
use NAND2X1  _1568_
timestamp 1702508443
transform 1 0 4170 0 1 1830
box -12 -8 72 272
use OAI21X1  _1569_
timestamp 1702508443
transform -1 0 4030 0 -1 2350
box -12 -8 92 272
use NAND2X1  _1570_
timestamp 1702508443
transform -1 0 4690 0 -1 2350
box -12 -8 72 272
use OAI21X1  _1571_
timestamp 1702508443
transform -1 0 3350 0 -1 3910
box -12 -8 92 272
use NOR2X1  _1572_
timestamp 1701862152
transform 1 0 3770 0 -1 3390
box -12 -8 74 272
use AOI21X1  _1573_
timestamp 1702508443
transform 1 0 4750 0 -1 3390
box -12 -8 92 272
use AOI21X1  _1574_
timestamp 1702508443
transform -1 0 3850 0 -1 5990
box -12 -8 92 272
use OAI21X1  _1575_
timestamp 1702508443
transform -1 0 3690 0 -1 5990
box -12 -8 92 272
use NAND2X1  _1576_
timestamp 1702508443
transform 1 0 3930 0 1 5470
box -12 -8 72 272
use INVX1  _1577_
timestamp 1701862152
transform 1 0 4250 0 1 5990
box -12 -8 52 272
use AOI21X1  _1578_
timestamp 1702508443
transform 1 0 4090 0 1 5990
box -12 -8 92 272
use OAI21X1  _1579_
timestamp 1702508443
transform 1 0 4050 0 1 4950
box -12 -8 92 272
use INVX1  _1580_
timestamp 1701862152
transform 1 0 4970 0 1 5470
box -12 -8 52 272
use NAND2X1  _1581_
timestamp 1702508443
transform -1 0 4370 0 1 4430
box -12 -8 72 272
use AOI22X1  _1582_
timestamp 1701862152
transform -1 0 4970 0 1 4430
box -14 -8 114 272
use NAND2X1  _1583_
timestamp 1702508443
transform 1 0 5030 0 1 4430
box -12 -8 72 272
use NOR2X1  _1584_
timestamp 1701862152
transform 1 0 4730 0 1 4430
box -12 -8 74 272
use NOR3X1  _1585_
timestamp 1701862152
transform 1 0 5010 0 -1 4950
box -12 -8 172 272
use INVX1  _1586_
timestamp 1701862152
transform 1 0 5770 0 1 4950
box -12 -8 52 272
use INVX1  _1587_
timestamp 1701862152
transform 1 0 5390 0 -1 4950
box -12 -8 52 272
use INVX1  _1588_
timestamp 1701862152
transform -1 0 5390 0 -1 4430
box -12 -8 52 272
use NAND2X1  _1589_
timestamp 1702508443
transform 1 0 5090 0 -1 4430
box -12 -8 72 272
use AOI21X1  _1590_
timestamp 1702508443
transform 1 0 5630 0 1 4950
box -12 -8 92 272
use NOR2X1  _1591_
timestamp 1701862152
transform -1 0 4930 0 1 4950
box -12 -8 74 272
use OAI21X1  _1592_
timestamp 1702508443
transform 1 0 5010 0 1 4950
box -12 -8 92 272
use OAI21X1  _1593_
timestamp 1702508443
transform -1 0 5230 0 1 4950
box -12 -8 92 272
use NAND3X1  _1594_
timestamp 1702508443
transform -1 0 5550 0 1 4950
box -12 -8 92 272
use OAI21X1  _1595_
timestamp 1702508443
transform -1 0 4930 0 -1 4950
box -12 -8 92 272
use AND2X2  _1596_
timestamp 1701862152
transform -1 0 4690 0 1 4950
box -12 -8 94 272
use AOI21X1  _1597_
timestamp 1702508443
transform 1 0 4470 0 1 4950
box -12 -8 92 272
use NAND3X1  _1598_
timestamp 1702508443
transform -1 0 5170 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1599_
timestamp 1702508443
transform 1 0 5090 0 1 5470
box -12 -8 92 272
use NAND3X1  _1600_
timestamp 1702508443
transform -1 0 5030 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1601_
timestamp 1702508443
transform -1 0 5390 0 1 4950
box -12 -8 92 272
use NAND3X1  _1602_
timestamp 1702508443
transform 1 0 4810 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1603_
timestamp 1702508443
transform 1 0 5710 0 -1 5990
box -12 -8 72 272
use INVX1  _1604_
timestamp 1701862152
transform 1 0 4250 0 1 3910
box -12 -8 52 272
use OAI21X1  _1605_
timestamp 1702508443
transform 1 0 4370 0 -1 5470
box -12 -8 92 272
use INVX1  _1606_
timestamp 1701862152
transform 1 0 4330 0 -1 4430
box -12 -8 52 272
use AND2X2  _1607_
timestamp 1701862152
transform 1 0 4370 0 1 3910
box -12 -8 94 272
use AND2X2  _1608_
timestamp 1701862152
transform 1 0 4430 0 1 4430
box -12 -8 94 272
use AOI22X1  _1609_
timestamp 1701862152
transform -1 0 4850 0 -1 4430
box -14 -8 114 272
use OAI21X1  _1610_
timestamp 1702508443
transform -1 0 4650 0 1 4430
box -12 -8 92 272
use AOI21X1  _1611_
timestamp 1702508443
transform -1 0 4670 0 -1 4430
box -12 -8 92 272
use NAND2X1  _1612_
timestamp 1702508443
transform 1 0 4450 0 -1 4430
box -12 -8 72 272
use AND2X2  _1613_
timestamp 1701862152
transform 1 0 4690 0 -1 4950
box -12 -8 94 272
use NAND2X1  _1614_
timestamp 1702508443
transform -1 0 4730 0 -1 5470
box -12 -8 72 272
use NAND2X1  _1615_
timestamp 1702508443
transform 1 0 4390 0 1 5470
box -12 -8 72 272
use NAND2X1  _1616_
timestamp 1702508443
transform 1 0 4570 0 -1 4950
box -12 -8 72 272
use NAND3X1  _1617_
timestamp 1702508443
transform 1 0 4530 0 1 5470
box -12 -8 92 272
use NAND2X1  _1618_
timestamp 1702508443
transform 1 0 5930 0 -1 5990
box -12 -8 72 272
use NAND2X1  _1619_
timestamp 1702508443
transform 1 0 6170 0 1 5990
box -12 -8 72 272
use NAND3X1  _1620_
timestamp 1702508443
transform 1 0 4670 0 1 5470
box -12 -8 92 272
use NAND2X1  _1621_
timestamp 1702508443
transform -1 0 4590 0 -1 5470
box -12 -8 72 272
use NAND2X1  _1622_
timestamp 1702508443
transform 1 0 4830 0 1 5470
box -12 -8 72 272
use NAND3X1  _1623_
timestamp 1702508443
transform -1 0 5650 0 -1 5990
box -12 -8 92 272
use NAND3X1  _1624_
timestamp 1702508443
transform -1 0 5530 0 1 5990
box -12 -8 92 272
use OAI21X1  _1625_
timestamp 1702508443
transform 1 0 4690 0 -1 5990
box -12 -8 92 272
use AOI21X1  _1626_
timestamp 1702508443
transform -1 0 5230 0 -1 5990
box -12 -8 92 272
use NOR2X1  _1627_
timestamp 1701862152
transform 1 0 6030 0 1 5990
box -12 -8 74 272
use OAI21X1  _1628_
timestamp 1702508443
transform -1 0 5050 0 1 5990
box -12 -8 92 272
use NAND3X1  _1629_
timestamp 1702508443
transform 1 0 4830 0 1 5990
box -12 -8 92 272
use NAND3X1  _1630_
timestamp 1702508443
transform -1 0 5670 0 1 5990
box -12 -8 92 272
use OAI21X1  _1631_
timestamp 1702508443
transform 1 0 5130 0 1 5990
box -12 -8 92 272
use NAND3X1  _1632_
timestamp 1702508443
transform -1 0 5070 0 -1 5990
box -12 -8 92 272
use NAND3X1  _1633_
timestamp 1702508443
transform -1 0 4930 0 -1 5990
box -12 -8 92 272
use NOR3X1  _1634_
timestamp 1701862152
transform -1 0 2610 0 1 5990
box -12 -8 172 272
use AOI21X1  _1635_
timestamp 1702508443
transform 1 0 2830 0 1 5990
box -12 -8 92 272
use AOI21X1  _1636_
timestamp 1702508443
transform -1 0 4610 0 1 5990
box -12 -8 92 272
use AOI21X1  _1637_
timestamp 1702508443
transform -1 0 4750 0 1 5990
box -12 -8 92 272
use OAI21X1  _1638_
timestamp 1702508443
transform -1 0 4450 0 1 5990
box -12 -8 92 272
use NAND2X1  _1639_
timestamp 1702508443
transform -1 0 5010 0 1 3910
box -12 -8 72 272
use AND2X2  _1640_
timestamp 1701862152
transform -1 0 4910 0 -1 2870
box -12 -8 94 272
use OAI21X1  _1641_
timestamp 1702508443
transform -1 0 4990 0 1 2350
box -12 -8 92 272
use OAI21X1  _1642_
timestamp 1702508443
transform -1 0 4830 0 1 2350
box -12 -8 92 272
use INVX1  _1643_
timestamp 1701862152
transform 1 0 5470 0 1 1830
box -12 -8 52 272
use OAI21X1  _1644_
timestamp 1702508443
transform 1 0 5050 0 -1 3390
box -12 -8 92 272
use AOI21X1  _1645_
timestamp 1702508443
transform -1 0 5810 0 1 5990
box -12 -8 92 272
use OAI21X1  _1646_
timestamp 1702508443
transform 1 0 5290 0 1 5990
box -12 -8 92 272
use NAND2X1  _1647_
timestamp 1702508443
transform 1 0 5230 0 -1 5470
box -12 -8 72 272
use INVX1  _1648_
timestamp 1701862152
transform 1 0 5670 0 -1 5470
box -12 -8 52 272
use AND2X2  _1649_
timestamp 1701862152
transform 1 0 5250 0 1 5470
box -12 -8 94 272
use INVX1  _1650_
timestamp 1701862152
transform 1 0 5830 0 -1 5990
box -12 -8 52 272
use AOI21X1  _1651_
timestamp 1702508443
transform 1 0 5710 0 1 5470
box -12 -8 92 272
use OAI21X1  _1652_
timestamp 1702508443
transform 1 0 5230 0 -1 4950
box -12 -8 92 272
use NAND2X1  _1653_
timestamp 1702508443
transform 1 0 5330 0 1 4430
box -12 -8 72 272
use INVX1  _1654_
timestamp 1701862152
transform -1 0 5930 0 1 4430
box -12 -8 52 272
use AOI22X1  _1655_
timestamp 1701862152
transform 1 0 5150 0 1 4430
box -14 -8 114 272
use INVX1  _1656_
timestamp 1701862152
transform 1 0 5470 0 1 4430
box -12 -8 52 272
use AND2X2  _1657_
timestamp 1701862152
transform 1 0 4510 0 1 3910
box -12 -8 94 272
use NAND2X1  _1658_
timestamp 1702508443
transform 1 0 5230 0 -1 4430
box -12 -8 72 272
use NAND3X1  _1659_
timestamp 1702508443
transform 1 0 5730 0 1 4430
box -12 -8 92 272
use NAND2X1  _1660_
timestamp 1702508443
transform -1 0 5290 0 1 3910
box -12 -8 72 272
use NOR2X1  _1661_
timestamp 1701862152
transform -1 0 5430 0 1 3910
box -12 -8 74 272
use OAI21X1  _1662_
timestamp 1702508443
transform 1 0 5830 0 -1 4430
box -12 -8 92 272
use NAND3X1  _1663_
timestamp 1702508443
transform 1 0 6170 0 1 4430
box -12 -8 92 272
use INVX1  _1664_
timestamp 1701862152
transform -1 0 5830 0 -1 4950
box -12 -8 52 272
use NOR3X1  _1665_
timestamp 1701862152
transform -1 0 5770 0 -1 4430
box -12 -8 172 272
use AOI21X1  _1666_
timestamp 1702508443
transform 1 0 5590 0 1 4430
box -12 -8 92 272
use OAI21X1  _1667_
timestamp 1702508443
transform 1 0 5650 0 -1 4950
box -12 -8 92 272
use AOI21X1  _1668_
timestamp 1702508443
transform -1 0 6370 0 1 4950
box -12 -8 92 272
use INVX1  _1669_
timestamp 1701862152
transform 1 0 5870 0 1 4950
box -12 -8 52 272
use OAI21X1  _1670_
timestamp 1702508443
transform -1 0 5590 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1671_
timestamp 1702508443
transform -1 0 6090 0 1 4430
box -12 -8 92 272
use AOI21X1  _1672_
timestamp 1702508443
transform 1 0 5970 0 1 4950
box -12 -8 92 272
use INVX1  _1673_
timestamp 1701862152
transform 1 0 4050 0 1 3390
box -12 -8 52 272
use XOR2X1  _1674_
timestamp 1702508443
transform -1 0 4310 0 -1 3910
box -12 -8 132 272
use OR2X2  _1675_
timestamp 1702508443
transform 1 0 5990 0 -1 4430
box -12 -8 92 272
use NAND2X1  _1676_
timestamp 1702508443
transform 1 0 6270 0 -1 4430
box -12 -8 72 272
use NAND2X1  _1677_
timestamp 1702508443
transform -1 0 6190 0 -1 4430
box -12 -8 72 272
use OAI21X1  _1678_
timestamp 1702508443
transform -1 0 6210 0 1 4950
box -12 -8 92 272
use NAND3X1  _1679_
timestamp 1702508443
transform 1 0 5890 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1680_
timestamp 1702508443
transform 1 0 6310 0 -1 4950
box -12 -8 92 272
use INVX1  _1681_
timestamp 1701862152
transform 1 0 6190 0 -1 4950
box -12 -8 52 272
use NAND3X1  _1682_
timestamp 1702508443
transform 1 0 6030 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1683_
timestamp 1702508443
transform -1 0 5870 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1684_
timestamp 1702508443
transform 1 0 5930 0 -1 5470
box -12 -8 72 272
use OAI21X1  _1685_
timestamp 1702508443
transform 1 0 5870 0 1 5470
box -12 -8 92 272
use NAND3X1  _1686_
timestamp 1702508443
transform -1 0 5590 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1687_
timestamp 1702508443
transform -1 0 6130 0 -1 5990
box -12 -8 92 272
use NAND3X1  _1688_
timestamp 1702508443
transform 1 0 6070 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1689_
timestamp 1702508443
transform -1 0 6370 0 1 5470
box -12 -8 72 272
use NAND3X1  _1690_
timestamp 1702508443
transform 1 0 6170 0 1 5470
box -12 -8 92 272
use NAND3X1  _1691_
timestamp 1702508443
transform -1 0 5430 0 -1 5470
box -12 -8 92 272
use INVX1  _1692_
timestamp 1701862152
transform -1 0 5510 0 -1 5990
box -12 -8 52 272
use AOI21X1  _1693_
timestamp 1702508443
transform 1 0 5310 0 -1 5990
box -12 -8 92 272
use AOI21X1  _1694_
timestamp 1702508443
transform -1 0 6090 0 1 5470
box -12 -8 92 272
use AOI21X1  _1695_
timestamp 1702508443
transform -1 0 5630 0 1 5470
box -12 -8 92 272
use OAI21X1  _1696_
timestamp 1702508443
transform -1 0 5470 0 1 5470
box -12 -8 92 272
use NAND2X1  _1697_
timestamp 1702508443
transform 1 0 5390 0 1 3390
box -12 -8 72 272
use AND2X2  _1698_
timestamp 1701862152
transform 1 0 5770 0 -1 3390
box -12 -8 94 272
use NOR2X1  _1699_
timestamp 1701862152
transform 1 0 5630 0 -1 3390
box -12 -8 74 272
use OAI21X1  _1700_
timestamp 1702508443
transform -1 0 5410 0 1 2870
box -12 -8 92 272
use OAI21X1  _1701_
timestamp 1702508443
transform 1 0 5310 0 1 1830
box -12 -8 92 272
use NAND2X1  _1702_
timestamp 1702508443
transform 1 0 6050 0 -1 2350
box -12 -8 72 272
use NOR2X1  _1703_
timestamp 1701862152
transform -1 0 5270 0 -1 3390
box -12 -8 74 272
use NAND3X1  _1704_
timestamp 1702508443
transform 1 0 4890 0 -1 3390
box -12 -8 92 272
use NAND2X1  _1705_
timestamp 1702508443
transform -1 0 5410 0 -1 3390
box -12 -8 72 272
use AOI22X1  _1706_
timestamp 1701862152
transform -1 0 5570 0 -1 3390
box -14 -8 114 272
use NAND2X1  _1707_
timestamp 1702508443
transform 1 0 5490 0 1 2870
box -12 -8 72 272
use OAI21X1  _1708_
timestamp 1702508443
transform 1 0 6230 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1709_
timestamp 1702508443
transform 1 0 6310 0 1 4430
box -12 -8 72 272
use OAI21X1  _1710_
timestamp 1702508443
transform 1 0 5670 0 1 3910
box -12 -8 92 272
use OAI21X1  _1711_
timestamp 1702508443
transform 1 0 5450 0 -1 4430
box -12 -8 92 272
use NAND2X1  _1712_
timestamp 1702508443
transform -1 0 5150 0 1 3910
box -12 -8 72 272
use AOI21X1  _1713_
timestamp 1702508443
transform 1 0 4790 0 1 3910
box -12 -8 92 272
use NAND2X1  _1714_
timestamp 1702508443
transform 1 0 4650 0 1 3910
box -12 -8 72 272
use NAND2X1  _1715_
timestamp 1702508443
transform -1 0 4610 0 -1 3910
box -12 -8 72 272
use NOR2X1  _1716_
timestamp 1701862152
transform 1 0 4670 0 -1 3910
box -12 -8 74 272
use NOR2X1  _1717_
timestamp 1701862152
transform -1 0 5050 0 -1 3910
box -12 -8 74 272
use XNOR2X1  _1718_
timestamp 1702508443
transform 1 0 5110 0 -1 3910
box -12 -8 132 272
use NOR2X1  _1719_
timestamp 1701862152
transform 1 0 5310 0 -1 3910
box -12 -8 74 272
use OAI21X1  _1720_
timestamp 1702508443
transform -1 0 5590 0 1 3910
box -12 -8 92 272
use INVX1  _1721_
timestamp 1701862152
transform 1 0 5830 0 1 3390
box -12 -8 52 272
use INVX1  _1722_
timestamp 1701862152
transform 1 0 4730 0 1 3390
box -12 -8 52 272
use NAND2X1  _1723_
timestamp 1702508443
transform 1 0 4150 0 1 3390
box -12 -8 72 272
use NAND2X1  _1724_
timestamp 1702508443
transform 1 0 4850 0 1 3390
box -12 -8 72 272
use OR2X2  _1725_
timestamp 1702508443
transform 1 0 4990 0 1 3390
box -12 -8 92 272
use NAND2X1  _1726_
timestamp 1702508443
transform 1 0 5130 0 1 3390
box -12 -8 72 272
use OAI21X1  _1727_
timestamp 1702508443
transform -1 0 5830 0 -1 3910
box -12 -8 92 272
use OR2X2  _1728_
timestamp 1702508443
transform 1 0 5430 0 -1 3910
box -12 -8 92 272
use INVX1  _1729_
timestamp 1701862152
transform 1 0 5270 0 1 3390
box -12 -8 52 272
use NAND3X1  _1730_
timestamp 1702508443
transform 1 0 5590 0 -1 3910
box -12 -8 92 272
use NAND3X1  _1731_
timestamp 1702508443
transform 1 0 6030 0 -1 3910
box -12 -8 92 272
use NAND2X1  _1732_
timestamp 1702508443
transform 1 0 5910 0 -1 3910
box -12 -8 72 272
use NAND3X1  _1733_
timestamp 1702508443
transform 1 0 5810 0 1 3910
box -12 -8 92 272
use NAND3X1  _1734_
timestamp 1702508443
transform -1 0 6410 0 -1 3390
box -12 -8 92 272
use INVX1  _1735_
timestamp 1701862152
transform -1 0 6370 0 -1 5990
box -12 -8 52 272
use INVX1  _1736_
timestamp 1701862152
transform -1 0 6110 0 1 3910
box -12 -8 52 272
use INVX1  _1737_
timestamp 1701862152
transform 1 0 5970 0 1 3910
box -12 -8 52 272
use OAI21X1  _1738_
timestamp 1702508443
transform 1 0 6170 0 1 3910
box -12 -8 92 272
use NAND3X1  _1739_
timestamp 1702508443
transform -1 0 6270 0 -1 3910
box -12 -8 92 272
use INVX1  _1740_
timestamp 1701862152
transform 1 0 6230 0 1 3390
box -12 -8 52 272
use NAND2X1  _1741_
timestamp 1702508443
transform 1 0 6330 0 -1 3910
box -12 -8 72 272
use NAND2X1  _1742_
timestamp 1702508443
transform 1 0 6350 0 1 3390
box -12 -8 72 272
use AND2X2  _1743_
timestamp 1701862152
transform 1 0 5930 0 1 2870
box -12 -8 94 272
use XNOR2X1  _1744_
timestamp 1702508443
transform 1 0 5670 0 1 2350
box -12 -8 132 272
use OAI21X1  _1745_
timestamp 1702508443
transform 1 0 5650 0 -1 2350
box -12 -8 92 272
use INVX1  _1746_
timestamp 1701862152
transform 1 0 6290 0 -1 2870
box -12 -8 52 272
use AND2X2  _1747_
timestamp 1701862152
transform 1 0 6150 0 -1 2870
box -12 -8 94 272
use AOI21X1  _1748_
timestamp 1702508443
transform -1 0 6390 0 1 3910
box -12 -8 92 272
use OAI22X1  _1749_
timestamp 1701862152
transform 1 0 4810 0 -1 3910
box -12 -8 112 272
use INVX1  _1750_
timestamp 1701862152
transform -1 0 4130 0 -1 3910
box -12 -8 52 272
use OAI21X1  _1751_
timestamp 1702508443
transform 1 0 4390 0 -1 3910
box -12 -8 92 272
use NOR2X1  _1752_
timestamp 1701862152
transform 1 0 3970 0 -1 3910
box -12 -8 74 272
use NAND2X1  _1753_
timestamp 1702508443
transform 1 0 4270 0 1 3390
box -12 -8 72 272
use AND2X2  _1754_
timestamp 1701862152
transform 1 0 4410 0 1 3390
box -12 -8 94 272
use XOR2X1  _1755_
timestamp 1702508443
transform 1 0 4730 0 1 2870
box -12 -8 132 272
use XNOR2X1  _1756_
timestamp 1702508443
transform -1 0 4370 0 -1 2870
box -12 -8 132 272
use AOI21X1  _1757_
timestamp 1702508443
transform 1 0 5530 0 1 3390
box -12 -8 92 272
use INVX1  _1758_
timestamp 1701862152
transform 1 0 6070 0 -1 3390
box -12 -8 52 272
use NAND3X1  _1759_
timestamp 1702508443
transform 1 0 5690 0 1 3390
box -12 -8 92 272
use NAND3X1  _1760_
timestamp 1702508443
transform 1 0 6170 0 -1 3390
box -12 -8 92 272
use INVX1  _1761_
timestamp 1701862152
transform 1 0 5950 0 1 3390
box -12 -8 52 272
use OAI21X1  _1762_
timestamp 1702508443
transform 1 0 6070 0 1 3390
box -12 -8 92 272
use NAND2X1  _1763_
timestamp 1702508443
transform 1 0 6190 0 -1 5990
box -12 -8 72 272
use XOR2X1  _1764_
timestamp 1702508443
transform -1 0 6370 0 1 2870
box -12 -8 132 272
use INVX1  _1765_
timestamp 1701862152
transform 1 0 6050 0 1 2350
box -12 -8 52 272
use OAI21X1  _1766_
timestamp 1702508443
transform -1 0 6250 0 1 2350
box -12 -8 92 272
use NOR2X1  _1767_
timestamp 1701862152
transform -1 0 6390 0 1 2350
box -12 -8 74 272
use AOI21X1  _1768_
timestamp 1702508443
transform -1 0 6430 0 -1 2350
box -12 -8 92 272
use AOI22X1  _1769_
timestamp 1701862152
transform -1 0 6290 0 -1 2350
box -14 -8 114 272
use NAND2X1  _1770_
timestamp 1702508443
transform 1 0 5370 0 -1 2350
box -12 -8 72 272
use NAND3X1  _1771_
timestamp 1702508443
transform -1 0 5870 0 1 2870
box -12 -8 92 272
use AOI21X1  _1772_
timestamp 1702508443
transform 1 0 5630 0 1 2870
box -12 -8 92 272
use NAND2X1  _1773_
timestamp 1702508443
transform -1 0 6350 0 1 5990
box -12 -8 72 272
use OAI21X1  _1774_
timestamp 1702508443
transform -1 0 6170 0 1 2870
box -12 -8 92 272
use NOR2X1  _1775_
timestamp 1701862152
transform -1 0 6070 0 -1 2870
box -12 -8 74 272
use AOI21X1  _1776_
timestamp 1702508443
transform -1 0 6010 0 -1 3390
box -12 -8 92 272
use NAND2X1  _1777_
timestamp 1702508443
transform -1 0 4970 0 1 2870
box -12 -8 72 272
use OAI21X1  _1778_
timestamp 1702508443
transform 1 0 3530 0 1 3390
box -12 -8 92 272
use XOR2X1  _1779_
timestamp 1702508443
transform 1 0 4570 0 -1 3390
box -12 -8 132 272
use NAND2X1  _1780_
timestamp 1702508443
transform 1 0 4430 0 -1 2870
box -12 -8 72 272
use OR2X2  _1781_
timestamp 1702508443
transform 1 0 4690 0 -1 2870
box -12 -8 92 272
use NAND2X1  _1782_
timestamp 1702508443
transform -1 0 4610 0 -1 2870
box -12 -8 72 272
use NAND2X1  _1783_
timestamp 1702508443
transform 1 0 4990 0 -1 2870
box -12 -8 72 272
use NAND2X1  _1784_
timestamp 1702508443
transform -1 0 5110 0 1 2870
box -12 -8 72 272
use OAI21X1  _1785_
timestamp 1702508443
transform 1 0 5170 0 1 2870
box -12 -8 92 272
use OR2X2  _1786_
timestamp 1702508443
transform 1 0 5290 0 -1 2870
box -12 -8 92 272
use NAND2X1  _1787_
timestamp 1702508443
transform -1 0 5630 0 -1 2870
box -12 -8 72 272
use AND2X2  _1788_
timestamp 1701862152
transform 1 0 5710 0 -1 2870
box -12 -8 94 272
use XOR2X1  _1789_
timestamp 1702508443
transform -1 0 5990 0 1 2350
box -12 -8 132 272
use OAI21X1  _1790_
timestamp 1702508443
transform -1 0 5570 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1791_
timestamp 1702508443
transform -1 0 5950 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1792_
timestamp 1702508443
transform 1 0 5430 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1793_
timestamp 1702508443
transform -1 0 5210 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1794_
timestamp 1702508443
transform -1 0 4650 0 1 3390
box -12 -8 92 272
use XOR2X1  _1795_
timestamp 1702508443
transform -1 0 4690 0 1 2350
box -12 -8 132 272
use XNOR2X1  _1796_
timestamp 1702508443
transform -1 0 5190 0 1 2350
box -12 -8 132 272
use INVX1  _1797_
timestamp 1701862152
transform 1 0 5410 0 1 2350
box -12 -8 52 272
use NAND2X1  _1798_
timestamp 1702508443
transform -1 0 5590 0 1 2350
box -12 -8 72 272
use NAND3X1  _1799_
timestamp 1702508443
transform -1 0 5350 0 1 2350
box -12 -8 92 272
use AND2X2  _1800_
timestamp 1701862152
transform 1 0 5230 0 -1 2350
box -12 -8 94 272
use AOI22X1  _1801_
timestamp 1701862152
transform -1 0 5690 0 1 1830
box -14 -8 114 272
use INVX1  _1802_
timestamp 1701862152
transform -1 0 3530 0 -1 2350
box -12 -8 52 272
use INVX1  _1803_
timestamp 1701862152
transform -1 0 4570 0 -1 1830
box -12 -8 52 272
use NAND3X1  _1804_
timestamp 1702508443
transform -1 0 4450 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1805_
timestamp 1702508443
transform -1 0 4170 0 -1 2870
box -12 -8 72 272
use OAI21X1  _1806_
timestamp 1702508443
transform 1 0 3970 0 -1 2870
box -12 -8 92 272
use INVX1  _1807_
timestamp 1701862152
transform -1 0 3430 0 -1 2350
box -12 -8 52 272
use NAND2X1  _1808_
timestamp 1702508443
transform 1 0 4250 0 -1 2350
box -12 -8 72 272
use OAI21X1  _1809_
timestamp 1702508443
transform 1 0 4090 0 -1 2350
box -12 -8 92 272
use INVX1  _1810_
timestamp 1701862152
transform -1 0 3690 0 1 2870
box -12 -8 52 272
use NAND2X1  _1811_
timestamp 1702508443
transform -1 0 4430 0 1 2870
box -12 -8 72 272
use OAI21X1  _1812_
timestamp 1702508443
transform 1 0 4210 0 1 2870
box -12 -8 92 272
use INVX1  _1813_
timestamp 1701862152
transform 1 0 3950 0 1 2350
box -12 -8 52 272
use NAND2X1  _1814_
timestamp 1702508443
transform -1 0 4270 0 1 2350
box -12 -8 72 272
use OAI21X1  _1815_
timestamp 1702508443
transform 1 0 4070 0 1 2350
box -12 -8 92 272
use NOR2X1  _1816_
timestamp 1701862152
transform -1 0 4370 0 1 1830
box -12 -8 74 272
use NOR2X1  _1817_
timestamp 1701862152
transform 1 0 3910 0 1 3390
box -12 -8 74 272
use AOI21X1  _1818_
timestamp 1702508443
transform 1 0 3910 0 -1 3390
box -12 -8 92 272
use NAND2X1  _1819_
timestamp 1702508443
transform 1 0 3590 0 -1 2350
box -12 -8 72 272
use OAI21X1  _1820_
timestamp 1702508443
transform -1 0 3890 0 -1 3910
box -12 -8 92 272
use NAND2X1  _1821_
timestamp 1702508443
transform 1 0 3670 0 -1 3910
box -12 -8 72 272
use OAI21X1  _1822_
timestamp 1702508443
transform -1 0 4170 0 1 3910
box -12 -8 92 272
use NAND2X1  _1823_
timestamp 1702508443
transform 1 0 4090 0 1 2870
box -12 -8 72 272
use OAI21X1  _1824_
timestamp 1702508443
transform 1 0 4050 0 -1 3390
box -12 -8 92 272
use INVX1  _1825_
timestamp 1701862152
transform 1 0 3190 0 -1 2870
box -12 -8 52 272
use OAI21X1  _1826_
timestamp 1702508443
transform 1 0 2910 0 1 1830
box -12 -8 92 272
use OAI21X1  _1827_
timestamp 1702508443
transform -1 0 2790 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1828_
timestamp 1702508443
transform 1 0 2870 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1829_
timestamp 1702508443
transform -1 0 3330 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1830_
timestamp 1702508443
transform -1 0 2910 0 1 2870
box -12 -8 92 272
use OAI21X1  _1831_
timestamp 1702508443
transform -1 0 2830 0 -1 2870
box -12 -8 92 272
use OAI21X1  _1832_
timestamp 1702508443
transform 1 0 3250 0 1 2870
box -12 -8 92 272
use OAI21X1  _1833_
timestamp 1702508443
transform -1 0 3390 0 -1 2870
box -12 -8 92 272
use NAND2X1  _1834_
timestamp 1702508443
transform -1 0 4090 0 1 1830
box -12 -8 72 272
use OAI21X1  _1835_
timestamp 1702508443
transform 1 0 3650 0 1 1830
box -12 -8 92 272
use NOR2X1  _1836_
timestamp 1701862152
transform -1 0 3370 0 1 2350
box -12 -8 74 272
use AOI21X1  _1837_
timestamp 1702508443
transform -1 0 3510 0 1 2350
box -12 -8 92 272
use NOR2X1  _1838_
timestamp 1701862152
transform -1 0 3110 0 -1 2870
box -12 -8 74 272
use AOI21X1  _1839_
timestamp 1702508443
transform 1 0 2890 0 -1 2870
box -12 -8 92 272
use NAND2X1  _1840_
timestamp 1702508443
transform 1 0 2390 0 1 1830
box -12 -8 72 272
use OAI21X1  _1841_
timestamp 1702508443
transform 1 0 2110 0 1 1830
box -12 -8 92 272
use NAND2X1  _1842_
timestamp 1702508443
transform -1 0 2130 0 1 3390
box -12 -8 72 272
use OAI21X1  _1843_
timestamp 1702508443
transform -1 0 2290 0 1 3390
box -12 -8 92 272
use NAND2X1  _1844_
timestamp 1702508443
transform -1 0 2590 0 1 2870
box -12 -8 72 272
use OAI21X1  _1845_
timestamp 1702508443
transform -1 0 2750 0 1 2870
box -12 -8 92 272
use NAND2X1  _1846_
timestamp 1702508443
transform -1 0 2410 0 1 3390
box -12 -8 72 272
use OAI21X1  _1847_
timestamp 1702508443
transform -1 0 2570 0 1 3390
box -12 -8 92 272
use NAND2X1  _1848_
timestamp 1702508443
transform 1 0 2850 0 -1 3910
box -12 -8 72 272
use OAI21X1  _1849_
timestamp 1702508443
transform 1 0 2690 0 -1 3910
box -12 -8 92 272
use DFFPOSX1  _1850_ digital_ETRI
timestamp 1702508443
transform -1 0 2030 0 -1 3390
box -13 -8 253 272
use DFFPOSX1  _1851_
timestamp 1702508443
transform -1 0 2190 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1852_
timestamp 1702508443
transform 1 0 3090 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1853_
timestamp 1702508443
transform 1 0 3350 0 -1 3910
box -13 -8 253 272
use DFFPOSX1  _1854_
timestamp 1702508443
transform 1 0 4030 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1855_
timestamp 1702508443
transform 1 0 4650 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1856_
timestamp 1702508443
transform 1 0 4730 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1857_
timestamp 1702508443
transform -1 0 5490 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1858_
timestamp 1702508443
transform 1 0 3490 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1859_
timestamp 1702508443
transform -1 0 5610 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1860_
timestamp 1702508443
transform 1 0 4790 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1861_
timestamp 1702508443
transform 1 0 3810 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1862_
timestamp 1702508443
transform 1 0 5450 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1863_
timestamp 1702508443
transform 1 0 5450 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1864_
timestamp 1702508443
transform 1 0 4810 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1865_
timestamp 1702508443
transform 1 0 5610 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1866_
timestamp 1702508443
transform 1 0 6050 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1867_
timestamp 1702508443
transform 1 0 5690 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1868_
timestamp 1702508443
transform -1 0 5650 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1869_
timestamp 1702508443
transform 1 0 5950 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1870_
timestamp 1702508443
transform 1 0 3510 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1871_
timestamp 1702508443
transform 1 0 4110 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1872_
timestamp 1702508443
transform 1 0 3130 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1873_
timestamp 1702508443
transform 1 0 4630 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1874_
timestamp 1702508443
transform 1 0 2990 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1875_
timestamp 1702508443
transform 1 0 3810 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1876_
timestamp 1702508443
transform -1 0 3550 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1877_
timestamp 1702508443
transform -1 0 3950 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1878_
timestamp 1702508443
transform -1 0 4810 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1879_
timestamp 1702508443
transform 1 0 3650 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1880_
timestamp 1702508443
transform -1 0 4930 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1881_
timestamp 1702508443
transform -1 0 6090 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1882_
timestamp 1702508443
transform 1 0 5730 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1883_
timestamp 1702508443
transform 1 0 6030 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1884_
timestamp 1702508443
transform 1 0 4930 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1885_
timestamp 1702508443
transform 1 0 5690 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1886_
timestamp 1702508443
transform 1 0 3650 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1887_
timestamp 1702508443
transform -1 0 4550 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1888_
timestamp 1702508443
transform 1 0 4430 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1889_
timestamp 1702508443
transform 1 0 4270 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1890_
timestamp 1702508443
transform 1 0 4130 0 -1 3390
box -13 -8 253 272
use DFFPOSX1  _1891_
timestamp 1702508443
transform 1 0 3790 0 1 3910
box -13 -8 253 272
use DFFPOSX1  _1892_
timestamp 1702508443
transform 1 0 4010 0 -1 4430
box -13 -8 253 272
use DFFPOSX1  _1893_
timestamp 1702508443
transform 1 0 3610 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1894_
timestamp 1702508443
transform -1 0 2690 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1895_
timestamp 1702508443
transform -1 0 3190 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1896_
timestamp 1702508443
transform -1 0 2670 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1897_
timestamp 1702508443
transform -1 0 3570 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1898_
timestamp 1702508443
transform -1 0 3970 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1899_
timestamp 1702508443
transform -1 0 3230 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1900_
timestamp 1702508443
transform -1 0 2990 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1901_
timestamp 1702508443
transform -1 0 2050 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1902_
timestamp 1702508443
transform 1 0 2450 0 -1 3390
box -13 -8 253 272
use DFFPOSX1  _1903_
timestamp 1702508443
transform -1 0 2430 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1904_
timestamp 1702508443
transform 1 0 2570 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1905_
timestamp 1702508443
transform -1 0 2630 0 -1 3910
box -13 -8 253 272
use DFFPOSX1  _1906_
timestamp 1702508443
transform -1 0 4070 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1907_
timestamp 1702508443
transform -1 0 4050 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1908_
timestamp 1702508443
transform 1 0 4150 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1909_
timestamp 1702508443
transform -1 0 4630 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1910_
timestamp 1702508443
transform 1 0 4490 0 -1 1310
box -13 -8 253 272
use BUFX2  _1911_ digital_ETRI
timestamp 1702508443
transform 1 0 6310 0 -1 790
box -12 -8 72 272
use BUFX2  _1912_
timestamp 1702508443
transform 1 0 2210 0 1 3910
box -12 -8 72 272
use BUFX2  _1913_
timestamp 1702508443
transform 1 0 2150 0 1 5990
box -12 -8 72 272
use BUFX2  _1914_
timestamp 1702508443
transform 1 0 3690 0 1 5470
box -12 -8 72 272
use BUFX2  _1915_
timestamp 1702508443
transform 1 0 3810 0 1 5470
box -12 -8 72 272
use BUFX2  _1916_
timestamp 1702508443
transform 1 0 6330 0 1 790
box -12 -8 72 272
use BUFX2  _1917_
timestamp 1702508443
transform 1 0 6170 0 -1 790
box -12 -8 72 272
use BUFX2  _1918_
timestamp 1702508443
transform 1 0 5890 0 1 5990
box -12 -8 72 272
use BUFX2  _1919_
timestamp 1702508443
transform -1 0 5790 0 1 790
box -12 -8 72 272
use BUFX2  BUFX2_insert0
timestamp 1702508443
transform 1 0 4810 0 -1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert1
timestamp 1702508443
transform -1 0 4450 0 1 270
box -12 -8 72 272
use BUFX2  BUFX2_insert2
timestamp 1702508443
transform -1 0 4330 0 -1 270
box -12 -8 72 272
use BUFX2  BUFX2_insert3
timestamp 1702508443
transform 1 0 5390 0 -1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert4
timestamp 1702508443
transform 1 0 5570 0 1 270
box -12 -8 72 272
use BUFX2  BUFX2_insert12
timestamp 1702508443
transform 1 0 2130 0 1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert13
timestamp 1702508443
transform 1 0 2250 0 1 1830
box -12 -8 72 272
use BUFX2  BUFX2_insert14
timestamp 1702508443
transform 1 0 1370 0 -1 1830
box -12 -8 72 272
use BUFX2  BUFX2_insert15
timestamp 1702508443
transform -1 0 1990 0 -1 2350
box -12 -8 72 272
use BUFX2  BUFX2_insert16
timestamp 1702508443
transform -1 0 3630 0 1 2350
box -12 -8 72 272
use BUFX2  BUFX2_insert17
timestamp 1702508443
transform 1 0 3130 0 1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert18
timestamp 1702508443
transform -1 0 3450 0 1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert19
timestamp 1702508443
transform -1 0 3090 0 -1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert20
timestamp 1702508443
transform 1 0 3970 0 1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert21
timestamp 1702508443
transform -1 0 4150 0 1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert22
timestamp 1702508443
transform -1 0 5730 0 -1 1830
box -12 -8 72 272
use BUFX2  BUFX2_insert23
timestamp 1702508443
transform -1 0 3670 0 1 790
box -12 -8 72 272
use BUFX2  BUFX2_insert24
timestamp 1702508443
transform 1 0 4130 0 1 790
box -12 -8 72 272
use BUFX2  BUFX2_insert25
timestamp 1702508443
transform 1 0 4950 0 -1 1310
box -12 -8 72 272
use CLKBUF1  CLKBUF1_insert5 digital_ETRI
timestamp 1701862152
transform 1 0 4970 0 1 1310
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert6
timestamp 1701862152
transform 1 0 4950 0 1 1830
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert7
timestamp 1701862152
transform -1 0 4330 0 1 270
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert8
timestamp 1701862152
transform -1 0 3870 0 1 2350
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert9
timestamp 1701862152
transform -1 0 3650 0 -1 2870
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert10
timestamp 1701862152
transform 1 0 4710 0 1 1310
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert11
timestamp 1701862152
transform -1 0 4890 0 1 1830
box -12 -8 192 272
use FILL  FILL94650x78150 digital_ETRI
timestamp 1701859473
transform -1 0 6330 0 -1 5470
box -12 -8 32 272
use FILL  FILL94950x150
timestamp 1701859473
transform -1 0 6350 0 -1 270
box -12 -8 32 272
use FILL  FILL94950x39150
timestamp 1701859473
transform -1 0 6350 0 -1 2870
box -12 -8 32 272
use FILL  FILL94950x62550
timestamp 1701859473
transform -1 0 6350 0 -1 4430
box -12 -8 32 272
use FILL  FILL94950x78150
timestamp 1701859473
transform -1 0 6350 0 -1 5470
box -12 -8 32 272
use FILL  FILL95250x150
timestamp 1701859473
transform -1 0 6370 0 -1 270
box -12 -8 32 272
use FILL  FILL95250x4050
timestamp 1701859473
transform 1 0 6350 0 1 270
box -12 -8 32 272
use FILL  FILL95250x39150
timestamp 1701859473
transform -1 0 6370 0 -1 2870
box -12 -8 32 272
use FILL  FILL95250x62550
timestamp 1701859473
transform -1 0 6370 0 -1 4430
box -12 -8 32 272
use FILL  FILL95250x78150
timestamp 1701859473
transform -1 0 6370 0 -1 5470
box -12 -8 32 272
use FILL  FILL95250x89850
timestamp 1701859473
transform 1 0 6350 0 1 5990
box -12 -8 32 272
use FILL  FILL95550x150
timestamp 1701859473
transform -1 0 6390 0 -1 270
box -12 -8 32 272
use FILL  FILL95550x4050
timestamp 1701859473
transform 1 0 6370 0 1 270
box -12 -8 32 272
use FILL  FILL95550x7950
timestamp 1701859473
transform -1 0 6390 0 -1 790
box -12 -8 32 272
use FILL  FILL95550x15750
timestamp 1701859473
transform -1 0 6390 0 -1 1310
box -12 -8 32 272
use FILL  FILL95550x23550
timestamp 1701859473
transform -1 0 6390 0 -1 1830
box -12 -8 32 272
use FILL  FILL95550x39150
timestamp 1701859473
transform -1 0 6390 0 -1 2870
box -12 -8 32 272
use FILL  FILL95550x43050
timestamp 1701859473
transform 1 0 6370 0 1 2870
box -12 -8 32 272
use FILL  FILL95550x62550
timestamp 1701859473
transform -1 0 6390 0 -1 4430
box -12 -8 32 272
use FILL  FILL95550x66450
timestamp 1701859473
transform 1 0 6370 0 1 4430
box -12 -8 32 272
use FILL  FILL95550x74250
timestamp 1701859473
transform 1 0 6370 0 1 4950
box -12 -8 32 272
use FILL  FILL95550x78150
timestamp 1701859473
transform -1 0 6390 0 -1 5470
box -12 -8 32 272
use FILL  FILL95550x82050
timestamp 1701859473
transform 1 0 6370 0 1 5470
box -12 -8 32 272
use FILL  FILL95550x85950
timestamp 1701859473
transform -1 0 6390 0 -1 5990
box -12 -8 32 272
use FILL  FILL95550x89850
timestamp 1701859473
transform 1 0 6370 0 1 5990
box -12 -8 32 272
use FILL  FILL95850x150
timestamp 1701859473
transform -1 0 6410 0 -1 270
box -12 -8 32 272
use FILL  FILL95850x4050
timestamp 1701859473
transform 1 0 6390 0 1 270
box -12 -8 32 272
use FILL  FILL95850x7950
timestamp 1701859473
transform -1 0 6410 0 -1 790
box -12 -8 32 272
use FILL  FILL95850x11850
timestamp 1701859473
transform 1 0 6390 0 1 790
box -12 -8 32 272
use FILL  FILL95850x15750
timestamp 1701859473
transform -1 0 6410 0 -1 1310
box -12 -8 32 272
use FILL  FILL95850x23550
timestamp 1701859473
transform -1 0 6410 0 -1 1830
box -12 -8 32 272
use FILL  FILL95850x27450
timestamp 1701859473
transform 1 0 6390 0 1 1830
box -12 -8 32 272
use FILL  FILL95850x35250
timestamp 1701859473
transform 1 0 6390 0 1 2350
box -12 -8 32 272
use FILL  FILL95850x39150
timestamp 1701859473
transform -1 0 6410 0 -1 2870
box -12 -8 32 272
use FILL  FILL95850x43050
timestamp 1701859473
transform 1 0 6390 0 1 2870
box -12 -8 32 272
use FILL  FILL95850x54750
timestamp 1701859473
transform -1 0 6410 0 -1 3910
box -12 -8 32 272
use FILL  FILL95850x58650
timestamp 1701859473
transform 1 0 6390 0 1 3910
box -12 -8 32 272
use FILL  FILL95850x62550
timestamp 1701859473
transform -1 0 6410 0 -1 4430
box -12 -8 32 272
use FILL  FILL95850x66450
timestamp 1701859473
transform 1 0 6390 0 1 4430
box -12 -8 32 272
use FILL  FILL95850x70350
timestamp 1701859473
transform -1 0 6410 0 -1 4950
box -12 -8 32 272
use FILL  FILL95850x74250
timestamp 1701859473
transform 1 0 6390 0 1 4950
box -12 -8 32 272
use FILL  FILL95850x78150
timestamp 1701859473
transform -1 0 6410 0 -1 5470
box -12 -8 32 272
use FILL  FILL95850x82050
timestamp 1701859473
transform 1 0 6390 0 1 5470
box -12 -8 32 272
use FILL  FILL95850x85950
timestamp 1701859473
transform -1 0 6410 0 -1 5990
box -12 -8 32 272
use FILL  FILL95850x89850
timestamp 1701859473
transform 1 0 6390 0 1 5990
box -12 -8 32 272
use FILL  FILL96150x150
timestamp 1701859473
transform -1 0 6430 0 -1 270
box -12 -8 32 272
use FILL  FILL96150x4050
timestamp 1701859473
transform 1 0 6410 0 1 270
box -12 -8 32 272
use FILL  FILL96150x7950
timestamp 1701859473
transform -1 0 6430 0 -1 790
box -12 -8 32 272
use FILL  FILL96150x11850
timestamp 1701859473
transform 1 0 6410 0 1 790
box -12 -8 32 272
use FILL  FILL96150x15750
timestamp 1701859473
transform -1 0 6430 0 -1 1310
box -12 -8 32 272
use FILL  FILL96150x19650
timestamp 1701859473
transform 1 0 6410 0 1 1310
box -12 -8 32 272
use FILL  FILL96150x23550
timestamp 1701859473
transform -1 0 6430 0 -1 1830
box -12 -8 32 272
use FILL  FILL96150x27450
timestamp 1701859473
transform 1 0 6410 0 1 1830
box -12 -8 32 272
use FILL  FILL96150x35250
timestamp 1701859473
transform 1 0 6410 0 1 2350
box -12 -8 32 272
use FILL  FILL96150x39150
timestamp 1701859473
transform -1 0 6430 0 -1 2870
box -12 -8 32 272
use FILL  FILL96150x43050
timestamp 1701859473
transform 1 0 6410 0 1 2870
box -12 -8 32 272
use FILL  FILL96150x46950
timestamp 1701859473
transform -1 0 6430 0 -1 3390
box -12 -8 32 272
use FILL  FILL96150x50850
timestamp 1701859473
transform 1 0 6410 0 1 3390
box -12 -8 32 272
use FILL  FILL96150x54750
timestamp 1701859473
transform -1 0 6430 0 -1 3910
box -12 -8 32 272
use FILL  FILL96150x58650
timestamp 1701859473
transform 1 0 6410 0 1 3910
box -12 -8 32 272
use FILL  FILL96150x62550
timestamp 1701859473
transform -1 0 6430 0 -1 4430
box -12 -8 32 272
use FILL  FILL96150x66450
timestamp 1701859473
transform 1 0 6410 0 1 4430
box -12 -8 32 272
use FILL  FILL96150x70350
timestamp 1701859473
transform -1 0 6430 0 -1 4950
box -12 -8 32 272
use FILL  FILL96150x74250
timestamp 1701859473
transform 1 0 6410 0 1 4950
box -12 -8 32 272
use FILL  FILL96150x78150
timestamp 1701859473
transform -1 0 6430 0 -1 5470
box -12 -8 32 272
use FILL  FILL96150x82050
timestamp 1701859473
transform 1 0 6410 0 1 5470
box -12 -8 32 272
use FILL  FILL96150x85950
timestamp 1701859473
transform -1 0 6430 0 -1 5990
box -12 -8 32 272
use FILL  FILL96150x89850
timestamp 1701859473
transform 1 0 6410 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__922_
timestamp 1701859473
transform -1 0 4070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__923_
timestamp 1701859473
transform 1 0 4170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__924_
timestamp 1701859473
transform -1 0 5710 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__925_
timestamp 1701859473
transform -1 0 5810 0 1 790
box -12 -8 32 272
use FILL  FILL_0__926_
timestamp 1701859473
transform -1 0 6110 0 1 790
box -12 -8 32 272
use FILL  FILL_0__927_
timestamp 1701859473
transform -1 0 3730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__928_
timestamp 1701859473
transform -1 0 2930 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__929_
timestamp 1701859473
transform -1 0 4210 0 1 790
box -12 -8 32 272
use FILL  FILL_0__930_
timestamp 1701859473
transform -1 0 5950 0 1 790
box -12 -8 32 272
use FILL  FILL_0__931_
timestamp 1701859473
transform 1 0 5650 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__932_
timestamp 1701859473
transform -1 0 5930 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__933_
timestamp 1701859473
transform -1 0 5950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__934_
timestamp 1701859473
transform 1 0 5290 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__935_
timestamp 1701859473
transform -1 0 5970 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__936_
timestamp 1701859473
transform 1 0 5050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__937_
timestamp 1701859473
transform 1 0 5310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__938_
timestamp 1701859473
transform 1 0 5170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__939_
timestamp 1701859473
transform -1 0 5050 0 1 790
box -12 -8 32 272
use FILL  FILL_0__940_
timestamp 1701859473
transform 1 0 5010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__941_
timestamp 1701859473
transform 1 0 5850 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__942_
timestamp 1701859473
transform -1 0 5930 0 1 270
box -12 -8 32 272
use FILL  FILL_0__943_
timestamp 1701859473
transform -1 0 6070 0 1 270
box -12 -8 32 272
use FILL  FILL_0__944_
timestamp 1701859473
transform -1 0 5150 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__945_
timestamp 1701859473
transform -1 0 5810 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__946_
timestamp 1701859473
transform 1 0 1710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__947_
timestamp 1701859473
transform 1 0 1970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__948_
timestamp 1701859473
transform -1 0 1830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__949_
timestamp 1701859473
transform -1 0 2270 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__950_
timestamp 1701859473
transform 1 0 2250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__951_
timestamp 1701859473
transform 1 0 2110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__952_
timestamp 1701859473
transform 1 0 4370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__953_
timestamp 1701859473
transform 1 0 3230 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__954_
timestamp 1701859473
transform 1 0 3370 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__955_
timestamp 1701859473
transform 1 0 3550 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__956_
timestamp 1701859473
transform 1 0 3510 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__957_
timestamp 1701859473
transform 1 0 3630 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__958_
timestamp 1701859473
transform 1 0 1710 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__959_
timestamp 1701859473
transform -1 0 1870 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__960_
timestamp 1701859473
transform 1 0 2330 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__961_
timestamp 1701859473
transform 1 0 2190 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__962_
timestamp 1701859473
transform 1 0 2810 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__963_
timestamp 1701859473
transform -1 0 2970 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__964_
timestamp 1701859473
transform 1 0 2910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__965_
timestamp 1701859473
transform -1 0 3070 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__966_
timestamp 1701859473
transform -1 0 4430 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__967_
timestamp 1701859473
transform 1 0 3890 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__968_
timestamp 1701859473
transform -1 0 4290 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__969_
timestamp 1701859473
transform -1 0 5030 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__970_
timestamp 1701859473
transform -1 0 4370 0 1 790
box -12 -8 32 272
use FILL  FILL_0__971_
timestamp 1701859473
transform -1 0 4530 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__972_
timestamp 1701859473
transform 1 0 4890 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__973_
timestamp 1701859473
transform -1 0 4470 0 1 270
box -12 -8 32 272
use FILL  FILL_0__974_
timestamp 1701859473
transform -1 0 4590 0 1 270
box -12 -8 32 272
use FILL  FILL_0__975_
timestamp 1701859473
transform -1 0 5150 0 1 270
box -12 -8 32 272
use FILL  FILL_0__976_
timestamp 1701859473
transform -1 0 5030 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__977_
timestamp 1701859473
transform -1 0 4990 0 1 270
box -12 -8 32 272
use FILL  FILL_0__978_
timestamp 1701859473
transform 1 0 3730 0 1 270
box -12 -8 32 272
use FILL  FILL_0__979_
timestamp 1701859473
transform -1 0 3370 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__980_
timestamp 1701859473
transform -1 0 3510 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__981_
timestamp 1701859473
transform -1 0 5290 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__982_
timestamp 1701859473
transform -1 0 4350 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__983_
timestamp 1701859473
transform -1 0 5150 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__984_
timestamp 1701859473
transform -1 0 5330 0 1 790
box -12 -8 32 272
use FILL  FILL_0__985_
timestamp 1701859473
transform -1 0 3210 0 1 790
box -12 -8 32 272
use FILL  FILL_0__986_
timestamp 1701859473
transform 1 0 5190 0 1 790
box -12 -8 32 272
use FILL  FILL_0__987_
timestamp 1701859473
transform 1 0 4490 0 1 790
box -12 -8 32 272
use FILL  FILL_0__988_
timestamp 1701859473
transform -1 0 3630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__989_
timestamp 1701859473
transform -1 0 3770 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__990_
timestamp 1701859473
transform 1 0 3670 0 1 790
box -12 -8 32 272
use FILL  FILL_0__991_
timestamp 1701859473
transform -1 0 4670 0 1 790
box -12 -8 32 272
use FILL  FILL_0__992_
timestamp 1701859473
transform -1 0 5510 0 1 790
box -12 -8 32 272
use FILL  FILL_0__993_
timestamp 1701859473
transform -1 0 5750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__994_
timestamp 1701859473
transform -1 0 5770 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__995_
timestamp 1701859473
transform -1 0 5150 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__996_
timestamp 1701859473
transform -1 0 5170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__997_
timestamp 1701859473
transform 1 0 5630 0 1 270
box -12 -8 32 272
use FILL  FILL_0__998_
timestamp 1701859473
transform -1 0 5790 0 1 270
box -12 -8 32 272
use FILL  FILL_0__999_
timestamp 1701859473
transform 1 0 6290 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1000_
timestamp 1701859473
transform -1 0 6110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1001_
timestamp 1701859473
transform -1 0 6250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1002_
timestamp 1701859473
transform 1 0 6270 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1003_
timestamp 1701859473
transform 1 0 6090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1004_
timestamp 1701859473
transform -1 0 6230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1005_
timestamp 1701859473
transform 1 0 5150 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1006_
timestamp 1701859473
transform -1 0 5470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1007_
timestamp 1701859473
transform 1 0 5250 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1008_
timestamp 1701859473
transform 1 0 5930 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1009_
timestamp 1701859473
transform 1 0 6190 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1010_
timestamp 1701859473
transform -1 0 6230 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1011_
timestamp 1701859473
transform 1 0 3290 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1012_
timestamp 1701859473
transform -1 0 2650 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1013_
timestamp 1701859473
transform 1 0 1710 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1014_
timestamp 1701859473
transform 1 0 3450 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1015_
timestamp 1701859473
transform 1 0 2690 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1016_
timestamp 1701859473
transform -1 0 3370 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1017_
timestamp 1701859473
transform -1 0 3250 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1018_
timestamp 1701859473
transform -1 0 3390 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1019_
timestamp 1701859473
transform 1 0 3130 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1020_
timestamp 1701859473
transform -1 0 3010 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1021_
timestamp 1701859473
transform -1 0 2950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1022_
timestamp 1701859473
transform 1 0 2630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1023_
timestamp 1701859473
transform 1 0 3050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1024_
timestamp 1701859473
transform 1 0 3190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1025_
timestamp 1701859473
transform 1 0 3310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1026_
timestamp 1701859473
transform 1 0 3410 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1027_
timestamp 1701859473
transform 1 0 3570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1028_
timestamp 1701859473
transform -1 0 3510 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1029_
timestamp 1701859473
transform -1 0 3650 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1030_
timestamp 1701859473
transform -1 0 3790 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1031_
timestamp 1701859473
transform 1 0 4350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1032_
timestamp 1701859473
transform 1 0 3950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1033_
timestamp 1701859473
transform 1 0 3370 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1034_
timestamp 1701859473
transform -1 0 2790 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1035_
timestamp 1701859473
transform 1 0 930 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1036_
timestamp 1701859473
transform 1 0 2770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1037_
timestamp 1701859473
transform -1 0 3030 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1038_
timestamp 1701859473
transform 1 0 2510 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1039_
timestamp 1701859473
transform 1 0 3110 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1040_
timestamp 1701859473
transform 1 0 2330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1041_
timestamp 1701859473
transform 1 0 2170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1042_
timestamp 1701859473
transform 1 0 2130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1043_
timestamp 1701859473
transform -1 0 2290 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1044_
timestamp 1701859473
transform -1 0 2710 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1045_
timestamp 1701859473
transform -1 0 2070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1046_
timestamp 1701859473
transform 1 0 2150 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1047_
timestamp 1701859473
transform 1 0 2410 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1048_
timestamp 1701859473
transform -1 0 2870 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1049_
timestamp 1701859473
transform -1 0 2570 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1050_
timestamp 1701859473
transform -1 0 2250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1051_
timestamp 1701859473
transform -1 0 2390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1052_
timestamp 1701859473
transform 1 0 2790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1053_
timestamp 1701859473
transform 1 0 2470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1054_
timestamp 1701859473
transform 1 0 2030 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1055_
timestamp 1701859473
transform 1 0 2690 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1056_
timestamp 1701859473
transform 1 0 2790 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1057_
timestamp 1701859473
transform 1 0 2630 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1058_
timestamp 1701859473
transform 1 0 2470 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1059_
timestamp 1701859473
transform -1 0 2970 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1060_
timestamp 1701859473
transform 1 0 3090 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1061_
timestamp 1701859473
transform 1 0 4870 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1062_
timestamp 1701859473
transform -1 0 2550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1063_
timestamp 1701859473
transform 1 0 2530 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1064_
timestamp 1701859473
transform -1 0 1470 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1065_
timestamp 1701859473
transform -1 0 2230 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1066_
timestamp 1701859473
transform -1 0 1890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1067_
timestamp 1701859473
transform 1 0 2090 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1068_
timestamp 1701859473
transform -1 0 1990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1069_
timestamp 1701859473
transform -1 0 1450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1070_
timestamp 1701859473
transform 1 0 1870 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1071_
timestamp 1701859473
transform 1 0 2030 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1072_
timestamp 1701859473
transform -1 0 1750 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1073_
timestamp 1701859473
transform -1 0 1830 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1074_
timestamp 1701859473
transform -1 0 1730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1075_
timestamp 1701859473
transform -1 0 1610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1076_
timestamp 1701859473
transform 1 0 1470 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1077_
timestamp 1701859473
transform -1 0 1970 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1078_
timestamp 1701859473
transform -1 0 1550 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1079_
timestamp 1701859473
transform -1 0 1830 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1080_
timestamp 1701859473
transform 1 0 1650 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1081_
timestamp 1701859473
transform -1 0 1730 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1082_
timestamp 1701859473
transform 1 0 1930 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1083_
timestamp 1701859473
transform 1 0 1630 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1084_
timestamp 1701859473
transform 1 0 1710 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1085_
timestamp 1701859473
transform -1 0 1730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1086_
timestamp 1701859473
transform -1 0 2550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1087_
timestamp 1701859473
transform 1 0 1570 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1088_
timestamp 1701859473
transform -1 0 1570 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1089_
timestamp 1701859473
transform 1 0 1790 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1090_
timestamp 1701859473
transform 1 0 1830 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1091_
timestamp 1701859473
transform -1 0 2270 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1092_
timestamp 1701859473
transform -1 0 2410 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1093_
timestamp 1701859473
transform -1 0 2370 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1094_
timestamp 1701859473
transform 1 0 2750 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1095_
timestamp 1701859473
transform -1 0 2530 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1096_
timestamp 1701859473
transform 1 0 2890 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1097_
timestamp 1701859473
transform -1 0 3010 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1098_
timestamp 1701859473
transform 1 0 4470 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1099_
timestamp 1701859473
transform 1 0 3230 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1100_
timestamp 1701859473
transform -1 0 590 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1101_
timestamp 1701859473
transform -1 0 1590 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1102_
timestamp 1701859473
transform 1 0 1430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1103_
timestamp 1701859473
transform -1 0 770 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1104_
timestamp 1701859473
transform -1 0 1610 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1105_
timestamp 1701859473
transform 1 0 1190 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1106_
timestamp 1701859473
transform -1 0 1470 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1107_
timestamp 1701859473
transform 1 0 1310 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1108_
timestamp 1701859473
transform -1 0 1290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1109_
timestamp 1701859473
transform -1 0 770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1110_
timestamp 1701859473
transform 1 0 990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1111_
timestamp 1701859473
transform -1 0 630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1112_
timestamp 1701859473
transform -1 0 470 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1113_
timestamp 1701859473
transform -1 0 1130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1114_
timestamp 1701859473
transform 1 0 850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1115_
timestamp 1701859473
transform -1 0 890 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1116_
timestamp 1701859473
transform -1 0 1950 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1117_
timestamp 1701859473
transform 1 0 1530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1118_
timestamp 1701859473
transform -1 0 2370 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1119_
timestamp 1701859473
transform -1 0 1970 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1120_
timestamp 1701859473
transform -1 0 1830 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1121_
timestamp 1701859473
transform -1 0 2870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1122_
timestamp 1701859473
transform -1 0 2110 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1123_
timestamp 1701859473
transform -1 0 1590 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1124_
timestamp 1701859473
transform -1 0 1670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1125_
timestamp 1701859473
transform -1 0 3710 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1126_
timestamp 1701859473
transform -1 0 1830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1127_
timestamp 1701859473
transform -1 0 1390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1128_
timestamp 1701859473
transform -1 0 1210 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1129_
timestamp 1701859473
transform 1 0 610 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1130_
timestamp 1701859473
transform 1 0 1030 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1131_
timestamp 1701859473
transform 1 0 610 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1132_
timestamp 1701859473
transform -1 0 1350 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1133_
timestamp 1701859473
transform -1 0 950 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1134_
timestamp 1701859473
transform -1 0 790 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1135_
timestamp 1701859473
transform -1 0 1270 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1136_
timestamp 1701859473
transform -1 0 1250 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1137_
timestamp 1701859473
transform 1 0 1070 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1138_
timestamp 1701859473
transform -1 0 1110 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1139_
timestamp 1701859473
transform -1 0 710 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1140_
timestamp 1701859473
transform -1 0 1430 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1141_
timestamp 1701859473
transform -1 0 970 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1142_
timestamp 1701859473
transform -1 0 810 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1143_
timestamp 1701859473
transform 1 0 850 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1144_
timestamp 1701859473
transform 1 0 1250 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1145_
timestamp 1701859473
transform -1 0 2150 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1146_
timestamp 1701859473
transform -1 0 1150 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1147_
timestamp 1701859473
transform -1 0 2010 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1148_
timestamp 1701859473
transform 1 0 2370 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1149_
timestamp 1701859473
transform -1 0 2230 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1150_
timestamp 1701859473
transform -1 0 2730 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1151_
timestamp 1701859473
transform 1 0 2850 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1152_
timestamp 1701859473
transform 1 0 4050 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1153_
timestamp 1701859473
transform -1 0 1750 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1154_
timestamp 1701859473
transform -1 0 430 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1155_
timestamp 1701859473
transform 1 0 2870 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1156_
timestamp 1701859473
transform -1 0 2290 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1157_
timestamp 1701859473
transform 1 0 850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1158_
timestamp 1701859473
transform -1 0 1490 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1159_
timestamp 1701859473
transform -1 0 1330 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1160_
timestamp 1701859473
transform -1 0 990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1161_
timestamp 1701859473
transform -1 0 310 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1162_
timestamp 1701859473
transform -1 0 1670 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1163_
timestamp 1701859473
transform 1 0 1790 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1164_
timestamp 1701859473
transform 1 0 1190 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1165_
timestamp 1701859473
transform 1 0 1430 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1166_
timestamp 1701859473
transform -1 0 1510 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1167_
timestamp 1701859473
transform -1 0 1050 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1168_
timestamp 1701859473
transform -1 0 790 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1169_
timestamp 1701859473
transform -1 0 1370 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1170_
timestamp 1701859473
transform -1 0 1110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1171_
timestamp 1701859473
transform 1 0 870 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1172_
timestamp 1701859473
transform 1 0 790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1173_
timestamp 1701859473
transform -1 0 1070 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1174_
timestamp 1701859473
transform -1 0 950 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1175_
timestamp 1701859473
transform 1 0 1330 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1176_
timestamp 1701859473
transform 1 0 1290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1177_
timestamp 1701859473
transform -1 0 1190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1178_
timestamp 1701859473
transform 1 0 1150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1179_
timestamp 1701859473
transform -1 0 1030 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1180_
timestamp 1701859473
transform -1 0 930 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1181_
timestamp 1701859473
transform -1 0 910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1182_
timestamp 1701859473
transform -1 0 610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1183_
timestamp 1701859473
transform -1 0 470 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1184_
timestamp 1701859473
transform 1 0 730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1185_
timestamp 1701859473
transform -1 0 1630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1186_
timestamp 1701859473
transform -1 0 1470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1187_
timestamp 1701859473
transform -1 0 1730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1188_
timestamp 1701859473
transform -1 0 1190 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1189_
timestamp 1701859473
transform 1 0 770 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1190_
timestamp 1701859473
transform -1 0 330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1191_
timestamp 1701859473
transform -1 0 650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1192_
timestamp 1701859473
transform -1 0 330 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1193_
timestamp 1701859473
transform -1 0 630 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1194_
timestamp 1701859473
transform -1 0 30 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1195_
timestamp 1701859473
transform 1 0 150 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1196_
timestamp 1701859473
transform 1 0 1370 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1197_
timestamp 1701859473
transform 1 0 170 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1198_
timestamp 1701859473
transform -1 0 470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1199_
timestamp 1701859473
transform 1 0 450 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1200_
timestamp 1701859473
transform 1 0 130 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1201_
timestamp 1701859473
transform -1 0 30 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1202_
timestamp 1701859473
transform -1 0 30 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1203_
timestamp 1701859473
transform -1 0 310 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1204_
timestamp 1701859473
transform 1 0 10 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1205_
timestamp 1701859473
transform 1 0 270 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1206_
timestamp 1701859473
transform -1 0 650 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1207_
timestamp 1701859473
transform 1 0 170 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1208_
timestamp 1701859473
transform 1 0 310 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1209_
timestamp 1701859473
transform 1 0 470 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1210_
timestamp 1701859473
transform 1 0 1590 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1211_
timestamp 1701859473
transform 1 0 1830 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1212_
timestamp 1701859473
transform 1 0 990 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1213_
timestamp 1701859473
transform 1 0 1410 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1214_
timestamp 1701859473
transform -1 0 1970 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1215_
timestamp 1701859473
transform 1 0 2510 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1216_
timestamp 1701859473
transform 1 0 3650 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1217_
timestamp 1701859473
transform 1 0 2070 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1218_
timestamp 1701859473
transform -1 0 810 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1219_
timestamp 1701859473
transform 1 0 1190 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1220_
timestamp 1701859473
transform 1 0 10 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1221_
timestamp 1701859473
transform -1 0 150 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1222_
timestamp 1701859473
transform 1 0 2410 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1223_
timestamp 1701859473
transform 1 0 1870 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1224_
timestamp 1701859473
transform -1 0 1450 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1225_
timestamp 1701859473
transform -1 0 870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1226_
timestamp 1701859473
transform -1 0 650 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1227_
timestamp 1701859473
transform 1 0 1250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1228_
timestamp 1701859473
transform -1 0 950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1229_
timestamp 1701859473
transform -1 0 30 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1230_
timestamp 1701859473
transform -1 0 190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1231_
timestamp 1701859473
transform 1 0 10 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1232_
timestamp 1701859473
transform -1 0 1610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1233_
timestamp 1701859473
transform -1 0 1310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1234_
timestamp 1701859473
transform 1 0 1010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1235_
timestamp 1701859473
transform -1 0 1150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1236_
timestamp 1701859473
transform -1 0 870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1237_
timestamp 1701859473
transform 1 0 910 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1238_
timestamp 1701859473
transform 1 0 1550 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1239_
timestamp 1701859473
transform -1 0 1330 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1240_
timestamp 1701859473
transform -1 0 1450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1241_
timestamp 1701859473
transform -1 0 790 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1242_
timestamp 1701859473
transform 1 0 710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1243_
timestamp 1701859473
transform -1 0 1030 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1244_
timestamp 1701859473
transform 1 0 870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1245_
timestamp 1701859473
transform -1 0 1590 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1246_
timestamp 1701859473
transform -1 0 1510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1247_
timestamp 1701859473
transform 1 0 1010 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1248_
timestamp 1701859473
transform -1 0 1650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1249_
timestamp 1701859473
transform 1 0 1130 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1250_
timestamp 1701859473
transform -1 0 1390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1251_
timestamp 1701859473
transform -1 0 1290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1252_
timestamp 1701859473
transform -1 0 990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1253_
timestamp 1701859473
transform -1 0 870 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1254_
timestamp 1701859473
transform -1 0 1150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1255_
timestamp 1701859473
transform -1 0 2350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1256_
timestamp 1701859473
transform -1 0 2210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1257_
timestamp 1701859473
transform -1 0 2710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1258_
timestamp 1701859473
transform -1 0 2050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1259_
timestamp 1701859473
transform -1 0 590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1260_
timestamp 1701859473
transform -1 0 330 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1261_
timestamp 1701859473
transform -1 0 590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1262_
timestamp 1701859473
transform 1 0 690 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1263_
timestamp 1701859473
transform 1 0 710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1264_
timestamp 1701859473
transform -1 0 290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1265_
timestamp 1701859473
transform -1 0 30 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1266_
timestamp 1701859473
transform -1 0 470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1267_
timestamp 1701859473
transform -1 0 310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1268_
timestamp 1701859473
transform 1 0 410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1269_
timestamp 1701859473
transform -1 0 490 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1270_
timestamp 1701859473
transform -1 0 330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1271_
timestamp 1701859473
transform 1 0 170 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1272_
timestamp 1701859473
transform 1 0 190 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1273_
timestamp 1701859473
transform 1 0 170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1274_
timestamp 1701859473
transform 1 0 470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1275_
timestamp 1701859473
transform 1 0 470 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1276_
timestamp 1701859473
transform -1 0 190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1277_
timestamp 1701859473
transform 1 0 10 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1278_
timestamp 1701859473
transform -1 0 190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1279_
timestamp 1701859473
transform -1 0 330 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1280_
timestamp 1701859473
transform -1 0 30 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1281_
timestamp 1701859473
transform 1 0 10 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1282_
timestamp 1701859473
transform 1 0 150 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1283_
timestamp 1701859473
transform -1 0 770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1284_
timestamp 1701859473
transform 1 0 310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1285_
timestamp 1701859473
transform 1 0 10 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1286_
timestamp 1701859473
transform 1 0 610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1287_
timestamp 1701859473
transform -1 0 650 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1288_
timestamp 1701859473
transform 1 0 470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1289_
timestamp 1701859473
transform 1 0 310 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1290_
timestamp 1701859473
transform 1 0 470 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1291_
timestamp 1701859473
transform 1 0 2330 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1292_
timestamp 1701859473
transform 1 0 2170 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1293_
timestamp 1701859473
transform -1 0 2910 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1294_
timestamp 1701859473
transform -1 0 3030 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1295_
timestamp 1701859473
transform 1 0 2670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1296_
timestamp 1701859473
transform -1 0 2930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1297_
timestamp 1701859473
transform -1 0 1090 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1298_
timestamp 1701859473
transform 1 0 770 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1299_
timestamp 1701859473
transform 1 0 10 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1300_
timestamp 1701859473
transform 1 0 10 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1301_
timestamp 1701859473
transform -1 0 150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1302_
timestamp 1701859473
transform 1 0 2890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1303_
timestamp 1701859473
transform -1 0 2370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1304_
timestamp 1701859473
transform -1 0 2590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1305_
timestamp 1701859473
transform 1 0 2030 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1306_
timestamp 1701859473
transform 1 0 1910 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1307_
timestamp 1701859473
transform -1 0 2210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1308_
timestamp 1701859473
transform -1 0 1910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1309_
timestamp 1701859473
transform 1 0 3110 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1310_
timestamp 1701859473
transform -1 0 2590 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1311_
timestamp 1701859473
transform -1 0 1730 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1312_
timestamp 1701859473
transform -1 0 1610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1313_
timestamp 1701859473
transform 1 0 1170 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1314_
timestamp 1701859473
transform -1 0 1450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1315_
timestamp 1701859473
transform -1 0 1770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1316_
timestamp 1701859473
transform -1 0 2050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1317_
timestamp 1701859473
transform 1 0 1010 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1318_
timestamp 1701859473
transform -1 0 1150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1319_
timestamp 1701859473
transform -1 0 990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1320_
timestamp 1701859473
transform -1 0 1210 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1321_
timestamp 1701859473
transform -1 0 1290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1322_
timestamp 1701859473
transform 1 0 770 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1323_
timestamp 1701859473
transform 1 0 610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1324_
timestamp 1701859473
transform -1 0 310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1325_
timestamp 1701859473
transform -1 0 170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1326_
timestamp 1701859473
transform 1 0 1470 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1327_
timestamp 1701859473
transform -1 0 1350 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1328_
timestamp 1701859473
transform 1 0 1010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1329_
timestamp 1701859473
transform 1 0 1050 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1330_
timestamp 1701859473
transform 1 0 1310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1331_
timestamp 1701859473
transform 1 0 1150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1332_
timestamp 1701859473
transform 1 0 1730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1333_
timestamp 1701859473
transform 1 0 2690 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1334_
timestamp 1701859473
transform 1 0 1970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1335_
timestamp 1701859473
transform -1 0 1630 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1336_
timestamp 1701859473
transform -1 0 1690 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1337_
timestamp 1701859473
transform 1 0 1310 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1338_
timestamp 1701859473
transform 1 0 1270 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1339_
timestamp 1701859473
transform -1 0 750 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1340_
timestamp 1701859473
transform 1 0 1430 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1341_
timestamp 1701859473
transform 1 0 1550 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1342_
timestamp 1701859473
transform -1 0 1650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1343_
timestamp 1701859473
transform -1 0 1790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1344_
timestamp 1701859473
transform 1 0 1490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1345_
timestamp 1701859473
transform -1 0 1470 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1346_
timestamp 1701859473
transform 1 0 1890 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1347_
timestamp 1701859473
transform -1 0 2090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1348_
timestamp 1701859473
transform -1 0 1610 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1349_
timestamp 1701859473
transform -1 0 1650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1350_
timestamp 1701859473
transform -1 0 870 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1351_
timestamp 1701859473
transform 1 0 1730 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1352_
timestamp 1701859473
transform -1 0 1370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1353_
timestamp 1701859473
transform -1 0 1210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1354_
timestamp 1701859473
transform -1 0 910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1355_
timestamp 1701859473
transform -1 0 1190 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1356_
timestamp 1701859473
transform -1 0 1010 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1357_
timestamp 1701859473
transform -1 0 1070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1358_
timestamp 1701859473
transform -1 0 630 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1359_
timestamp 1701859473
transform -1 0 330 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1360_
timestamp 1701859473
transform -1 0 570 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1361_
timestamp 1701859473
transform -1 0 430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1362_
timestamp 1701859473
transform -1 0 790 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1363_
timestamp 1701859473
transform -1 0 750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1364_
timestamp 1701859473
transform -1 0 490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1365_
timestamp 1701859473
transform 1 0 150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1366_
timestamp 1701859473
transform -1 0 870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1367_
timestamp 1701859473
transform -1 0 490 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1368_
timestamp 1701859473
transform -1 0 330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1369_
timestamp 1701859473
transform 1 0 170 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1370_
timestamp 1701859473
transform -1 0 170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1371_
timestamp 1701859473
transform -1 0 170 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1372_
timestamp 1701859473
transform 1 0 10 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1373_
timestamp 1701859473
transform -1 0 30 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1374_
timestamp 1701859473
transform 1 0 10 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1375_
timestamp 1701859473
transform 1 0 10 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1376_
timestamp 1701859473
transform 1 0 170 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1377_
timestamp 1701859473
transform 1 0 470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1378_
timestamp 1701859473
transform 1 0 310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1379_
timestamp 1701859473
transform 1 0 10 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1380_
timestamp 1701859473
transform 1 0 470 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1381_
timestamp 1701859473
transform 1 0 610 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1382_
timestamp 1701859473
transform 1 0 630 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1383_
timestamp 1701859473
transform 1 0 910 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1384_
timestamp 1701859473
transform -1 0 350 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1385_
timestamp 1701859473
transform 1 0 10 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1386_
timestamp 1701859473
transform -1 0 410 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1387_
timestamp 1701859473
transform 1 0 2150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1388_
timestamp 1701859473
transform 1 0 3130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1389_
timestamp 1701859473
transform -1 0 3030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1390_
timestamp 1701859473
transform 1 0 3230 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1391_
timestamp 1701859473
transform 1 0 3290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1392_
timestamp 1701859473
transform -1 0 3450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1393_
timestamp 1701859473
transform -1 0 4530 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1394_
timestamp 1701859473
transform -1 0 2290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1395_
timestamp 1701859473
transform 1 0 1990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1396_
timestamp 1701859473
transform 1 0 2370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1397_
timestamp 1701859473
transform 1 0 170 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1398_
timestamp 1701859473
transform 1 0 330 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1399_
timestamp 1701859473
transform -1 0 750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1400_
timestamp 1701859473
transform 1 0 10 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1401_
timestamp 1701859473
transform 1 0 10 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1402_
timestamp 1701859473
transform 1 0 110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1403_
timestamp 1701859473
transform 1 0 1750 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1404_
timestamp 1701859473
transform 1 0 2770 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1405_
timestamp 1701859473
transform 1 0 2510 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1406_
timestamp 1701859473
transform -1 0 2990 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1407_
timestamp 1701859473
transform -1 0 3590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1408_
timestamp 1701859473
transform 1 0 3030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1409_
timestamp 1701859473
transform -1 0 3350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1410_
timestamp 1701859473
transform 1 0 3170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1411_
timestamp 1701859473
transform -1 0 2430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1412_
timestamp 1701859473
transform 1 0 2730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1413_
timestamp 1701859473
transform 1 0 2710 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1414_
timestamp 1701859473
transform -1 0 2230 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1415_
timestamp 1701859473
transform 1 0 1430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1416_
timestamp 1701859473
transform 1 0 1830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1417_
timestamp 1701859473
transform -1 0 2130 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1418_
timestamp 1701859473
transform 1 0 2350 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1419_
timestamp 1701859473
transform 1 0 2550 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1420_
timestamp 1701859473
transform -1 0 1610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1421_
timestamp 1701859473
transform 1 0 1830 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1422_
timestamp 1701859473
transform -1 0 2430 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1423_
timestamp 1701859473
transform 1 0 1970 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1424_
timestamp 1701859473
transform -1 0 2470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1425_
timestamp 1701859473
transform -1 0 2070 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1426_
timestamp 1701859473
transform -1 0 2290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1427_
timestamp 1701859473
transform -1 0 2270 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1428_
timestamp 1701859473
transform 1 0 2110 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1429_
timestamp 1701859473
transform -1 0 1510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1430_
timestamp 1701859473
transform -1 0 1070 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1431_
timestamp 1701859473
transform -1 0 930 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1432_
timestamp 1701859473
transform 1 0 3030 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1433_
timestamp 1701859473
transform 1 0 3290 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1434_
timestamp 1701859473
transform -1 0 3030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1435_
timestamp 1701859473
transform 1 0 3410 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1436_
timestamp 1701859473
transform -1 0 2910 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1437_
timestamp 1701859473
transform -1 0 2870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1438_
timestamp 1701859473
transform -1 0 3050 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1439_
timestamp 1701859473
transform 1 0 3730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1440_
timestamp 1701859473
transform 1 0 3470 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1441_
timestamp 1701859473
transform -1 0 3350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1442_
timestamp 1701859473
transform -1 0 2890 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1443_
timestamp 1701859473
transform 1 0 2650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1444_
timestamp 1701859473
transform 1 0 2490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1445_
timestamp 1701859473
transform 1 0 2330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1446_
timestamp 1701859473
transform -1 0 4250 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1447_
timestamp 1701859473
transform 1 0 2550 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1448_
timestamp 1701859473
transform 1 0 1930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1449_
timestamp 1701859473
transform 1 0 1910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1450_
timestamp 1701859473
transform 1 0 2010 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1451_
timestamp 1701859473
transform -1 0 2410 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1452_
timestamp 1701859473
transform -1 0 2090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1453_
timestamp 1701859473
transform -1 0 2710 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1454_
timestamp 1701859473
transform -1 0 2290 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1455_
timestamp 1701859473
transform 1 0 2150 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1456_
timestamp 1701859473
transform 1 0 1630 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1457_
timestamp 1701859473
transform -1 0 1370 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1458_
timestamp 1701859473
transform -1 0 1230 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1459_
timestamp 1701859473
transform -1 0 750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1460_
timestamp 1701859473
transform -1 0 1330 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1461_
timestamp 1701859473
transform -1 0 1170 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1462_
timestamp 1701859473
transform -1 0 2390 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1463_
timestamp 1701859473
transform 1 0 1770 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1464_
timestamp 1701859473
transform -1 0 1490 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1465_
timestamp 1701859473
transform 1 0 2230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1466_
timestamp 1701859473
transform -1 0 670 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1467_
timestamp 1701859473
transform -1 0 350 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1468_
timestamp 1701859473
transform -1 0 1370 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1469_
timestamp 1701859473
transform 1 0 890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1470_
timestamp 1701859473
transform -1 0 830 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1471_
timestamp 1701859473
transform -1 0 510 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1472_
timestamp 1701859473
transform 1 0 170 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1473_
timestamp 1701859473
transform -1 0 450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1474_
timestamp 1701859473
transform -1 0 290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1475_
timestamp 1701859473
transform -1 0 490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1476_
timestamp 1701859473
transform -1 0 330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1477_
timestamp 1701859473
transform -1 0 30 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1478_
timestamp 1701859473
transform 1 0 130 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1479_
timestamp 1701859473
transform -1 0 30 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1480_
timestamp 1701859473
transform 1 0 170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1481_
timestamp 1701859473
transform -1 0 590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1482_
timestamp 1701859473
transform 1 0 490 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1483_
timestamp 1701859473
transform -1 0 750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1484_
timestamp 1701859473
transform 1 0 570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1485_
timestamp 1701859473
transform -1 0 450 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1486_
timestamp 1701859473
transform 1 0 270 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1487_
timestamp 1701859473
transform 1 0 630 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1488_
timestamp 1701859473
transform -1 0 3110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1489_
timestamp 1701859473
transform -1 0 3830 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1490_
timestamp 1701859473
transform 1 0 4370 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1491_
timestamp 1701859473
transform 1 0 3230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1492_
timestamp 1701859473
transform 1 0 3350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1493_
timestamp 1701859473
transform -1 0 630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1494_
timestamp 1701859473
transform 1 0 570 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1495_
timestamp 1701859473
transform -1 0 2230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1496_
timestamp 1701859473
transform 1 0 2810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1497_
timestamp 1701859473
transform -1 0 1130 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1498_
timestamp 1701859473
transform 1 0 950 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1499_
timestamp 1701859473
transform 1 0 2710 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1500_
timestamp 1701859473
transform -1 0 3470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1501_
timestamp 1701859473
transform -1 0 3810 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1502_
timestamp 1701859473
transform 1 0 3670 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1503_
timestamp 1701859473
transform -1 0 3950 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1504_
timestamp 1701859473
transform -1 0 3630 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1505_
timestamp 1701859473
transform -1 0 3490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1506_
timestamp 1701859473
transform -1 0 4870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1507_
timestamp 1701859473
transform 1 0 3890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1508_
timestamp 1701859473
transform -1 0 3870 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1509_
timestamp 1701859473
transform -1 0 3550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1510_
timestamp 1701859473
transform -1 0 3190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1511_
timestamp 1701859473
transform 1 0 3130 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1512_
timestamp 1701859473
transform -1 0 3250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1513_
timestamp 1701859473
transform 1 0 3670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1514_
timestamp 1701859473
transform -1 0 3590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1515_
timestamp 1701859473
transform -1 0 3310 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1516_
timestamp 1701859473
transform -1 0 2930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1517_
timestamp 1701859473
transform 1 0 2770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1518_
timestamp 1701859473
transform -1 0 2650 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1519_
timestamp 1701859473
transform 1 0 2570 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1520_
timestamp 1701859473
transform 1 0 3070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1521_
timestamp 1701859473
transform -1 0 3390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1522_
timestamp 1701859473
transform 1 0 3470 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1523_
timestamp 1701859473
transform 1 0 3210 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1524_
timestamp 1701859473
transform 1 0 1790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1525_
timestamp 1701859473
transform 1 0 1910 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1526_
timestamp 1701859473
transform 1 0 4110 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1527_
timestamp 1701859473
transform -1 0 4370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1528_
timestamp 1701859473
transform 1 0 4190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1529_
timestamp 1701859473
transform 1 0 3890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1530_
timestamp 1701859473
transform -1 0 4050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1531_
timestamp 1701859473
transform 1 0 4270 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1532_
timestamp 1701859473
transform -1 0 4710 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1533_
timestamp 1701859473
transform 1 0 3710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1534_
timestamp 1701859473
transform -1 0 4150 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1535_
timestamp 1701859473
transform -1 0 3990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1536_
timestamp 1701859473
transform -1 0 4130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1537_
timestamp 1701859473
transform -1 0 4150 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1538_
timestamp 1701859473
transform -1 0 4010 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1539_
timestamp 1701859473
transform -1 0 3850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1540_
timestamp 1701859473
transform -1 0 3770 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1541_
timestamp 1701859473
transform 1 0 3630 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1542_
timestamp 1701859473
transform 1 0 2510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1543_
timestamp 1701859473
transform 1 0 2650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1544_
timestamp 1701859473
transform 1 0 4330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1545_
timestamp 1701859473
transform -1 0 4190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1546_
timestamp 1701859473
transform 1 0 3890 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1547_
timestamp 1701859473
transform 1 0 4470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1548_
timestamp 1701859473
transform -1 0 3370 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1549_
timestamp 1701859473
transform -1 0 4050 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1550_
timestamp 1701859473
transform -1 0 3250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1551_
timestamp 1701859473
transform 1 0 1050 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1552_
timestamp 1701859473
transform -1 0 1210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1553_
timestamp 1701859473
transform 1 0 3850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1554_
timestamp 1701859473
transform -1 0 3510 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1555_
timestamp 1701859473
transform 1 0 2210 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1556_
timestamp 1701859473
transform -1 0 3090 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1557_
timestamp 1701859473
transform 1 0 2910 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1558_
timestamp 1701859473
transform 1 0 3070 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1559_
timestamp 1701859473
transform 1 0 3390 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1560_
timestamp 1701859473
transform 1 0 2610 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1561_
timestamp 1701859473
transform -1 0 3350 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1562_
timestamp 1701859473
transform -1 0 3190 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1563_
timestamp 1701859473
transform -1 0 3030 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1564_
timestamp 1701859473
transform -1 0 2950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1565_
timestamp 1701859473
transform -1 0 2850 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1566_
timestamp 1701859473
transform -1 0 3190 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1567_
timestamp 1701859473
transform 1 0 3490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1568_
timestamp 1701859473
transform 1 0 4090 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1569_
timestamp 1701859473
transform -1 0 3910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1570_
timestamp 1701859473
transform -1 0 4570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1571_
timestamp 1701859473
transform -1 0 3230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1572_
timestamp 1701859473
transform 1 0 3690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1573_
timestamp 1701859473
transform 1 0 4690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1574_
timestamp 1701859473
transform -1 0 3710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1575_
timestamp 1701859473
transform -1 0 3550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1576_
timestamp 1701859473
transform 1 0 3870 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1577_
timestamp 1701859473
transform 1 0 4170 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1578_
timestamp 1701859473
transform 1 0 4030 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1579_
timestamp 1701859473
transform 1 0 3970 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1580_
timestamp 1701859473
transform 1 0 4890 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1581_
timestamp 1701859473
transform -1 0 4270 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1582_
timestamp 1701859473
transform -1 0 4810 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1583_
timestamp 1701859473
transform 1 0 4970 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1584_
timestamp 1701859473
transform 1 0 4650 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1585_
timestamp 1701859473
transform 1 0 4930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1586_
timestamp 1701859473
transform 1 0 5710 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1587_
timestamp 1701859473
transform 1 0 5310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1588_
timestamp 1701859473
transform -1 0 5310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1589_
timestamp 1701859473
transform 1 0 5010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1590_
timestamp 1701859473
transform 1 0 5550 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1591_
timestamp 1701859473
transform -1 0 4830 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1592_
timestamp 1701859473
transform 1 0 4930 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1593_
timestamp 1701859473
transform -1 0 5110 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1594_
timestamp 1701859473
transform -1 0 5410 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1595_
timestamp 1701859473
transform -1 0 4790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1596_
timestamp 1701859473
transform -1 0 4570 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1597_
timestamp 1701859473
transform 1 0 4390 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1598_
timestamp 1701859473
transform -1 0 5050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1599_
timestamp 1701859473
transform 1 0 5010 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1600_
timestamp 1701859473
transform -1 0 4910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1601_
timestamp 1701859473
transform -1 0 5250 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1602_
timestamp 1701859473
transform 1 0 4730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1603_
timestamp 1701859473
transform 1 0 5650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1604_
timestamp 1701859473
transform 1 0 4170 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1605_
timestamp 1701859473
transform 1 0 4310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1606_
timestamp 1701859473
transform 1 0 4250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1607_
timestamp 1701859473
transform 1 0 4290 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1608_
timestamp 1701859473
transform 1 0 4370 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1609_
timestamp 1701859473
transform -1 0 4690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1610_
timestamp 1701859473
transform -1 0 4530 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1611_
timestamp 1701859473
transform -1 0 4530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1612_
timestamp 1701859473
transform 1 0 4370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1613_
timestamp 1701859473
transform 1 0 4630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1614_
timestamp 1701859473
transform -1 0 4610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1615_
timestamp 1701859473
transform 1 0 4330 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1616_
timestamp 1701859473
transform 1 0 4490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1617_
timestamp 1701859473
transform 1 0 4450 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1618_
timestamp 1701859473
transform 1 0 5870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1619_
timestamp 1701859473
transform 1 0 6090 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1620_
timestamp 1701859473
transform 1 0 4610 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1621_
timestamp 1701859473
transform -1 0 4470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1622_
timestamp 1701859473
transform 1 0 4750 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1623_
timestamp 1701859473
transform -1 0 5530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1624_
timestamp 1701859473
transform -1 0 5390 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1625_
timestamp 1701859473
transform 1 0 4630 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1626_
timestamp 1701859473
transform -1 0 5090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1627_
timestamp 1701859473
transform 1 0 5950 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1628_
timestamp 1701859473
transform -1 0 4930 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1629_
timestamp 1701859473
transform 1 0 4750 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1630_
timestamp 1701859473
transform -1 0 5550 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1631_
timestamp 1701859473
transform 1 0 5050 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1632_
timestamp 1701859473
transform -1 0 4950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1633_
timestamp 1701859473
transform -1 0 4790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1634_
timestamp 1701859473
transform -1 0 2390 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1635_
timestamp 1701859473
transform 1 0 2770 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1636_
timestamp 1701859473
transform -1 0 4470 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1637_
timestamp 1701859473
transform -1 0 4630 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1638_
timestamp 1701859473
transform -1 0 4310 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1639_
timestamp 1701859473
transform -1 0 4890 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1640_
timestamp 1701859473
transform -1 0 4790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1641_
timestamp 1701859473
transform -1 0 4850 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1642_
timestamp 1701859473
transform -1 0 4710 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1643_
timestamp 1701859473
transform 1 0 5390 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1644_
timestamp 1701859473
transform 1 0 4970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1645_
timestamp 1701859473
transform -1 0 5690 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1646_
timestamp 1701859473
transform 1 0 5210 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1647_
timestamp 1701859473
transform 1 0 5170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1648_
timestamp 1701859473
transform 1 0 5590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1649_
timestamp 1701859473
transform 1 0 5170 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1650_
timestamp 1701859473
transform 1 0 5770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1651_
timestamp 1701859473
transform 1 0 5630 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1652_
timestamp 1701859473
transform 1 0 5170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1653_
timestamp 1701859473
transform 1 0 5250 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1654_
timestamp 1701859473
transform -1 0 5830 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1655_
timestamp 1701859473
transform 1 0 5090 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1656_
timestamp 1701859473
transform 1 0 5390 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1657_
timestamp 1701859473
transform 1 0 4450 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1658_
timestamp 1701859473
transform 1 0 5150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1659_
timestamp 1701859473
transform 1 0 5670 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1660_
timestamp 1701859473
transform -1 0 5170 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1661_
timestamp 1701859473
transform -1 0 5310 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1662_
timestamp 1701859473
transform 1 0 5770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1663_
timestamp 1701859473
transform 1 0 6090 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1664_
timestamp 1701859473
transform -1 0 5750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1665_
timestamp 1701859473
transform -1 0 5550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1666_
timestamp 1701859473
transform 1 0 5510 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1667_
timestamp 1701859473
transform 1 0 5590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1668_
timestamp 1701859473
transform -1 0 6230 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1669_
timestamp 1701859473
transform 1 0 5810 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1670_
timestamp 1701859473
transform -1 0 5450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1671_
timestamp 1701859473
transform -1 0 5950 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1672_
timestamp 1701859473
transform 1 0 5910 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1673_
timestamp 1701859473
transform 1 0 3970 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1674_
timestamp 1701859473
transform -1 0 4150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1675_
timestamp 1701859473
transform 1 0 5910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1676_
timestamp 1701859473
transform 1 0 6190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1677_
timestamp 1701859473
transform -1 0 6090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1678_
timestamp 1701859473
transform -1 0 6070 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1679_
timestamp 1701859473
transform 1 0 5830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1680_
timestamp 1701859473
transform 1 0 6230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1681_
timestamp 1701859473
transform 1 0 6110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1682_
timestamp 1701859473
transform 1 0 5970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1683_
timestamp 1701859473
transform -1 0 5730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1684_
timestamp 1701859473
transform 1 0 5870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1685_
timestamp 1701859473
transform 1 0 5790 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1686_
timestamp 1701859473
transform -1 0 5450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1687_
timestamp 1701859473
transform -1 0 6010 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1688_
timestamp 1701859473
transform 1 0 5990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1689_
timestamp 1701859473
transform -1 0 6270 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1690_
timestamp 1701859473
transform 1 0 6090 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1691_
timestamp 1701859473
transform -1 0 5310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1692_
timestamp 1701859473
transform -1 0 5410 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1693_
timestamp 1701859473
transform 1 0 5230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1694_
timestamp 1701859473
transform -1 0 5970 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1695_
timestamp 1701859473
transform -1 0 5490 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1696_
timestamp 1701859473
transform -1 0 5350 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1697_
timestamp 1701859473
transform 1 0 5310 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1698_
timestamp 1701859473
transform 1 0 5690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1699_
timestamp 1701859473
transform 1 0 5570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1700_
timestamp 1701859473
transform -1 0 5270 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1701_
timestamp 1701859473
transform 1 0 5250 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1702_
timestamp 1701859473
transform 1 0 5970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1703_
timestamp 1701859473
transform -1 0 5150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1704_
timestamp 1701859473
transform 1 0 4830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1705_
timestamp 1701859473
transform -1 0 5290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1706_
timestamp 1701859473
transform -1 0 5430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1707_
timestamp 1701859473
transform 1 0 5410 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1708_
timestamp 1701859473
transform 1 0 6150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1709_
timestamp 1701859473
transform 1 0 6250 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1710_
timestamp 1701859473
transform 1 0 5590 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1711_
timestamp 1701859473
transform 1 0 5390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1712_
timestamp 1701859473
transform -1 0 5030 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1713_
timestamp 1701859473
transform 1 0 4710 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1714_
timestamp 1701859473
transform 1 0 4590 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1715_
timestamp 1701859473
transform -1 0 4490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1716_
timestamp 1701859473
transform 1 0 4610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1717_
timestamp 1701859473
transform -1 0 4930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1718_
timestamp 1701859473
transform 1 0 5050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1719_
timestamp 1701859473
transform 1 0 5230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1720_
timestamp 1701859473
transform -1 0 5450 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1721_
timestamp 1701859473
transform 1 0 5770 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1722_
timestamp 1701859473
transform 1 0 4650 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1723_
timestamp 1701859473
transform 1 0 4090 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1724_
timestamp 1701859473
transform 1 0 4770 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1725_
timestamp 1701859473
transform 1 0 4910 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1726_
timestamp 1701859473
transform 1 0 5070 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1727_
timestamp 1701859473
transform -1 0 5690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1728_
timestamp 1701859473
transform 1 0 5370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1729_
timestamp 1701859473
transform 1 0 5190 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1730_
timestamp 1701859473
transform 1 0 5510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1731_
timestamp 1701859473
transform 1 0 5970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1732_
timestamp 1701859473
transform 1 0 5830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1733_
timestamp 1701859473
transform 1 0 5750 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1734_
timestamp 1701859473
transform -1 0 6270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1735_
timestamp 1701859473
transform -1 0 6270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1736_
timestamp 1701859473
transform -1 0 6030 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1737_
timestamp 1701859473
transform 1 0 5890 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1738_
timestamp 1701859473
transform 1 0 6110 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1739_
timestamp 1701859473
transform -1 0 6130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1740_
timestamp 1701859473
transform 1 0 6150 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1741_
timestamp 1701859473
transform 1 0 6270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1742_
timestamp 1701859473
transform 1 0 6270 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1743_
timestamp 1701859473
transform 1 0 5870 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1744_
timestamp 1701859473
transform 1 0 5590 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1745_
timestamp 1701859473
transform 1 0 5570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1746_
timestamp 1701859473
transform 1 0 6230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1747_
timestamp 1701859473
transform 1 0 6070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1748_
timestamp 1701859473
transform -1 0 6270 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1749_
timestamp 1701859473
transform 1 0 4730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1750_
timestamp 1701859473
transform -1 0 4050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1751_
timestamp 1701859473
transform 1 0 4310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1752_
timestamp 1701859473
transform 1 0 3890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1753_
timestamp 1701859473
transform 1 0 4210 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1754_
timestamp 1701859473
transform 1 0 4330 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1755_
timestamp 1701859473
transform 1 0 4670 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1756_
timestamp 1701859473
transform -1 0 4190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1757_
timestamp 1701859473
transform 1 0 5450 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1758_
timestamp 1701859473
transform 1 0 6010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1759_
timestamp 1701859473
transform 1 0 5610 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1760_
timestamp 1701859473
transform 1 0 6110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1761_
timestamp 1701859473
transform 1 0 5870 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1762_
timestamp 1701859473
transform 1 0 5990 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1763_
timestamp 1701859473
transform 1 0 6130 0 -1 5990
box -12 -8 32 272
use FILL  FILL_0__1764_
timestamp 1701859473
transform -1 0 6190 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1765_
timestamp 1701859473
transform 1 0 5990 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1766_
timestamp 1701859473
transform -1 0 6110 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1767_
timestamp 1701859473
transform -1 0 6270 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1768_
timestamp 1701859473
transform -1 0 6310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1769_
timestamp 1701859473
transform -1 0 6130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1770_
timestamp 1701859473
transform 1 0 5310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1771_
timestamp 1701859473
transform -1 0 5730 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1772_
timestamp 1701859473
transform 1 0 5550 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1773_
timestamp 1701859473
transform -1 0 6250 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1774_
timestamp 1701859473
transform -1 0 6030 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1775_
timestamp 1701859473
transform -1 0 5970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1776_
timestamp 1701859473
transform -1 0 5870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1777_
timestamp 1701859473
transform -1 0 4870 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1778_
timestamp 1701859473
transform 1 0 3450 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1779_
timestamp 1701859473
transform 1 0 4490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1780_
timestamp 1701859473
transform 1 0 4370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1781_
timestamp 1701859473
transform 1 0 4610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1782_
timestamp 1701859473
transform -1 0 4510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1783_
timestamp 1701859473
transform 1 0 4910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1784_
timestamp 1701859473
transform -1 0 4990 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1785_
timestamp 1701859473
transform 1 0 5110 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1786_
timestamp 1701859473
transform 1 0 5210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1787_
timestamp 1701859473
transform -1 0 5530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1788_
timestamp 1701859473
transform 1 0 5630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1789_
timestamp 1701859473
transform -1 0 5810 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1790_
timestamp 1701859473
transform -1 0 5450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1791_
timestamp 1701859473
transform -1 0 5810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1792_
timestamp 1701859473
transform 1 0 5370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1793_
timestamp 1701859473
transform -1 0 5070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1794_
timestamp 1701859473
transform -1 0 4510 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1795_
timestamp 1701859473
transform -1 0 4530 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1796_
timestamp 1701859473
transform -1 0 5010 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1797_
timestamp 1701859473
transform 1 0 5350 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1798_
timestamp 1701859473
transform -1 0 5470 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1799_
timestamp 1701859473
transform -1 0 5210 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1800_
timestamp 1701859473
transform 1 0 5170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1801_
timestamp 1701859473
transform -1 0 5530 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1802_
timestamp 1701859473
transform -1 0 3450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1803_
timestamp 1701859473
transform -1 0 4470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1804_
timestamp 1701859473
transform -1 0 4310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1805_
timestamp 1701859473
transform -1 0 4070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1806_
timestamp 1701859473
transform 1 0 3890 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1807_
timestamp 1701859473
transform -1 0 3350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1808_
timestamp 1701859473
transform 1 0 4170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1809_
timestamp 1701859473
transform 1 0 4030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1810_
timestamp 1701859473
transform -1 0 3590 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1811_
timestamp 1701859473
transform -1 0 4310 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1812_
timestamp 1701859473
transform 1 0 4150 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1813_
timestamp 1701859473
transform 1 0 3870 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1814_
timestamp 1701859473
transform -1 0 4170 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1815_
timestamp 1701859473
transform 1 0 3990 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1816_
timestamp 1701859473
transform -1 0 4250 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1817_
timestamp 1701859473
transform 1 0 3850 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1818_
timestamp 1701859473
transform 1 0 3830 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1819_
timestamp 1701859473
transform 1 0 3530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1820_
timestamp 1701859473
transform -1 0 3750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1821_
timestamp 1701859473
transform 1 0 3590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1822_
timestamp 1701859473
transform -1 0 4050 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1823_
timestamp 1701859473
transform 1 0 4010 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1824_
timestamp 1701859473
transform 1 0 3990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1825_
timestamp 1701859473
transform 1 0 3110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1826_
timestamp 1701859473
transform 1 0 2830 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1827_
timestamp 1701859473
transform -1 0 2670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1828_
timestamp 1701859473
transform 1 0 2790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1829_
timestamp 1701859473
transform -1 0 3210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1830_
timestamp 1701859473
transform -1 0 2770 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1831_
timestamp 1701859473
transform -1 0 2690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1832_
timestamp 1701859473
transform 1 0 3190 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1833_
timestamp 1701859473
transform -1 0 3250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1834_
timestamp 1701859473
transform -1 0 3990 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1835_
timestamp 1701859473
transform 1 0 3570 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1836_
timestamp 1701859473
transform -1 0 3250 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1837_
timestamp 1701859473
transform -1 0 3390 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1838_
timestamp 1701859473
transform -1 0 2990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1839_
timestamp 1701859473
transform 1 0 2830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1840_
timestamp 1701859473
transform 1 0 2310 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1841_
timestamp 1701859473
transform 1 0 2050 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1842_
timestamp 1701859473
transform -1 0 2010 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1843_
timestamp 1701859473
transform -1 0 2150 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1844_
timestamp 1701859473
transform -1 0 2490 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1845_
timestamp 1701859473
transform -1 0 2610 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1846_
timestamp 1701859473
transform -1 0 2310 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1847_
timestamp 1701859473
transform -1 0 2430 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1848_
timestamp 1701859473
transform 1 0 2770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1849_
timestamp 1701859473
transform 1 0 2630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1911_
timestamp 1701859473
transform 1 0 6230 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1912_
timestamp 1701859473
transform 1 0 2150 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1913_
timestamp 1701859473
transform 1 0 2070 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1914_
timestamp 1701859473
transform 1 0 3610 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1915_
timestamp 1701859473
transform 1 0 3750 0 1 5470
box -12 -8 32 272
use FILL  FILL_0__1916_
timestamp 1701859473
transform 1 0 6250 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1917_
timestamp 1701859473
transform 1 0 6110 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1918_
timestamp 1701859473
transform 1 0 5810 0 1 5990
box -12 -8 32 272
use FILL  FILL_0__1919_
timestamp 1701859473
transform -1 0 5670 0 1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert0
timestamp 1701859473
transform 1 0 4730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert1
timestamp 1701859473
transform -1 0 4350 0 1 270
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert2
timestamp 1701859473
transform -1 0 4210 0 -1 270
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert3
timestamp 1701859473
transform 1 0 5330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert4
timestamp 1701859473
transform 1 0 5490 0 1 270
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert12
timestamp 1701859473
transform 1 0 2050 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert13
timestamp 1701859473
transform 1 0 2190 0 1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert14
timestamp 1701859473
transform 1 0 1290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert15
timestamp 1701859473
transform -1 0 1870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert16
timestamp 1701859473
transform -1 0 3530 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert17
timestamp 1701859473
transform 1 0 3050 0 1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert18
timestamp 1701859473
transform -1 0 3350 0 1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert19
timestamp 1701859473
transform -1 0 2970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert20
timestamp 1701859473
transform 1 0 3890 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert21
timestamp 1701859473
transform -1 0 4050 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert22
timestamp 1701859473
transform -1 0 5610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert23
timestamp 1701859473
transform -1 0 3570 0 1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert24
timestamp 1701859473
transform 1 0 4050 0 1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert25
timestamp 1701859473
transform 1 0 4870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert5
timestamp 1701859473
transform 1 0 4890 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert6
timestamp 1701859473
transform 1 0 4890 0 1 1830
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert7
timestamp 1701859473
transform -1 0 4090 0 1 270
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert8
timestamp 1701859473
transform -1 0 3650 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert9
timestamp 1701859473
transform -1 0 3410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert10
timestamp 1701859473
transform 1 0 4630 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert11
timestamp 1701859473
transform -1 0 4670 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__922_
timestamp 1701859473
transform -1 0 4090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__923_
timestamp 1701859473
transform 1 0 4190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__924_
timestamp 1701859473
transform -1 0 5730 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__925_
timestamp 1701859473
transform -1 0 5830 0 1 790
box -12 -8 32 272
use FILL  FILL_1__926_
timestamp 1701859473
transform -1 0 6130 0 1 790
box -12 -8 32 272
use FILL  FILL_1__927_
timestamp 1701859473
transform -1 0 3750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__928_
timestamp 1701859473
transform -1 0 2950 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__929_
timestamp 1701859473
transform -1 0 4230 0 1 790
box -12 -8 32 272
use FILL  FILL_1__930_
timestamp 1701859473
transform -1 0 5970 0 1 790
box -12 -8 32 272
use FILL  FILL_1__931_
timestamp 1701859473
transform 1 0 5670 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__932_
timestamp 1701859473
transform -1 0 5950 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__933_
timestamp 1701859473
transform -1 0 5970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__934_
timestamp 1701859473
transform 1 0 5310 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__935_
timestamp 1701859473
transform -1 0 5990 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__936_
timestamp 1701859473
transform 1 0 5070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__937_
timestamp 1701859473
transform 1 0 5330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__938_
timestamp 1701859473
transform 1 0 5190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__939_
timestamp 1701859473
transform -1 0 5070 0 1 790
box -12 -8 32 272
use FILL  FILL_1__940_
timestamp 1701859473
transform 1 0 5030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__941_
timestamp 1701859473
transform 1 0 5870 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__942_
timestamp 1701859473
transform -1 0 5950 0 1 270
box -12 -8 32 272
use FILL  FILL_1__943_
timestamp 1701859473
transform -1 0 6090 0 1 270
box -12 -8 32 272
use FILL  FILL_1__944_
timestamp 1701859473
transform -1 0 5170 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__945_
timestamp 1701859473
transform -1 0 5830 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__946_
timestamp 1701859473
transform 1 0 1730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__947_
timestamp 1701859473
transform 1 0 1990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__948_
timestamp 1701859473
transform -1 0 1850 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__949_
timestamp 1701859473
transform -1 0 2290 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__950_
timestamp 1701859473
transform 1 0 2270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__951_
timestamp 1701859473
transform 1 0 2130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__952_
timestamp 1701859473
transform 1 0 4390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__953_
timestamp 1701859473
transform 1 0 3250 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__954_
timestamp 1701859473
transform 1 0 3390 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__955_
timestamp 1701859473
transform 1 0 3570 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__956_
timestamp 1701859473
transform 1 0 3530 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__957_
timestamp 1701859473
transform 1 0 3650 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__958_
timestamp 1701859473
transform 1 0 1730 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__959_
timestamp 1701859473
transform -1 0 1890 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__960_
timestamp 1701859473
transform 1 0 2350 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__961_
timestamp 1701859473
transform 1 0 2210 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__962_
timestamp 1701859473
transform 1 0 2830 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__963_
timestamp 1701859473
transform -1 0 2990 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__964_
timestamp 1701859473
transform 1 0 2930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__965_
timestamp 1701859473
transform -1 0 3090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__966_
timestamp 1701859473
transform -1 0 4450 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__967_
timestamp 1701859473
transform 1 0 3910 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__968_
timestamp 1701859473
transform -1 0 4310 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__969_
timestamp 1701859473
transform -1 0 5050 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__970_
timestamp 1701859473
transform -1 0 4390 0 1 790
box -12 -8 32 272
use FILL  FILL_1__971_
timestamp 1701859473
transform -1 0 4550 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__972_
timestamp 1701859473
transform 1 0 4910 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__973_
timestamp 1701859473
transform -1 0 4490 0 1 270
box -12 -8 32 272
use FILL  FILL_1__974_
timestamp 1701859473
transform -1 0 4610 0 1 270
box -12 -8 32 272
use FILL  FILL_1__975_
timestamp 1701859473
transform -1 0 5170 0 1 270
box -12 -8 32 272
use FILL  FILL_1__976_
timestamp 1701859473
transform -1 0 5050 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__977_
timestamp 1701859473
transform -1 0 5010 0 1 270
box -12 -8 32 272
use FILL  FILL_1__978_
timestamp 1701859473
transform 1 0 3750 0 1 270
box -12 -8 32 272
use FILL  FILL_1__979_
timestamp 1701859473
transform -1 0 3390 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__980_
timestamp 1701859473
transform -1 0 3530 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__981_
timestamp 1701859473
transform -1 0 5310 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__982_
timestamp 1701859473
transform -1 0 4370 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__983_
timestamp 1701859473
transform -1 0 5170 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__984_
timestamp 1701859473
transform -1 0 5350 0 1 790
box -12 -8 32 272
use FILL  FILL_1__985_
timestamp 1701859473
transform -1 0 3230 0 1 790
box -12 -8 32 272
use FILL  FILL_1__986_
timestamp 1701859473
transform 1 0 5210 0 1 790
box -12 -8 32 272
use FILL  FILL_1__987_
timestamp 1701859473
transform 1 0 4510 0 1 790
box -12 -8 32 272
use FILL  FILL_1__988_
timestamp 1701859473
transform -1 0 3650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__989_
timestamp 1701859473
transform -1 0 3790 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__990_
timestamp 1701859473
transform 1 0 3690 0 1 790
box -12 -8 32 272
use FILL  FILL_1__991_
timestamp 1701859473
transform -1 0 4690 0 1 790
box -12 -8 32 272
use FILL  FILL_1__992_
timestamp 1701859473
transform -1 0 5530 0 1 790
box -12 -8 32 272
use FILL  FILL_1__993_
timestamp 1701859473
transform -1 0 5770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__994_
timestamp 1701859473
transform -1 0 5790 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__995_
timestamp 1701859473
transform -1 0 5170 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__996_
timestamp 1701859473
transform -1 0 5190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__997_
timestamp 1701859473
transform 1 0 5650 0 1 270
box -12 -8 32 272
use FILL  FILL_1__998_
timestamp 1701859473
transform -1 0 5810 0 1 270
box -12 -8 32 272
use FILL  FILL_1__999_
timestamp 1701859473
transform 1 0 6310 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1000_
timestamp 1701859473
transform -1 0 6130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1001_
timestamp 1701859473
transform -1 0 6270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1002_
timestamp 1701859473
transform 1 0 6290 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1003_
timestamp 1701859473
transform 1 0 6110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1004_
timestamp 1701859473
transform -1 0 6250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1005_
timestamp 1701859473
transform 1 0 5170 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1006_
timestamp 1701859473
transform -1 0 5490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1007_
timestamp 1701859473
transform 1 0 5270 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1008_
timestamp 1701859473
transform 1 0 5950 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1009_
timestamp 1701859473
transform 1 0 6210 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1010_
timestamp 1701859473
transform -1 0 6250 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1011_
timestamp 1701859473
transform 1 0 3310 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1012_
timestamp 1701859473
transform -1 0 2670 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1013_
timestamp 1701859473
transform 1 0 1730 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1014_
timestamp 1701859473
transform 1 0 3470 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1015_
timestamp 1701859473
transform 1 0 2710 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1016_
timestamp 1701859473
transform -1 0 3390 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1017_
timestamp 1701859473
transform -1 0 3270 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1018_
timestamp 1701859473
transform -1 0 3410 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1019_
timestamp 1701859473
transform 1 0 3150 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1020_
timestamp 1701859473
transform -1 0 3030 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1021_
timestamp 1701859473
transform -1 0 2970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1022_
timestamp 1701859473
transform 1 0 2650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1023_
timestamp 1701859473
transform 1 0 3070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1024_
timestamp 1701859473
transform 1 0 3210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1025_
timestamp 1701859473
transform 1 0 3330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1026_
timestamp 1701859473
transform 1 0 3430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1027_
timestamp 1701859473
transform 1 0 3590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1028_
timestamp 1701859473
transform -1 0 3530 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1029_
timestamp 1701859473
transform -1 0 3670 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1030_
timestamp 1701859473
transform -1 0 3810 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1031_
timestamp 1701859473
transform 1 0 4370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1032_
timestamp 1701859473
transform 1 0 3970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1033_
timestamp 1701859473
transform 1 0 3390 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1034_
timestamp 1701859473
transform -1 0 2810 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1035_
timestamp 1701859473
transform 1 0 950 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1036_
timestamp 1701859473
transform 1 0 2790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1037_
timestamp 1701859473
transform -1 0 3050 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1038_
timestamp 1701859473
transform 1 0 2530 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1039_
timestamp 1701859473
transform 1 0 3130 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1040_
timestamp 1701859473
transform 1 0 2350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1041_
timestamp 1701859473
transform 1 0 2190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1042_
timestamp 1701859473
transform 1 0 2150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1043_
timestamp 1701859473
transform -1 0 2310 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1044_
timestamp 1701859473
transform -1 0 2730 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1045_
timestamp 1701859473
transform -1 0 2090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1046_
timestamp 1701859473
transform 1 0 2170 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1047_
timestamp 1701859473
transform 1 0 2430 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1048_
timestamp 1701859473
transform -1 0 2890 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1049_
timestamp 1701859473
transform -1 0 2590 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1050_
timestamp 1701859473
transform -1 0 2270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1051_
timestamp 1701859473
transform -1 0 2410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1052_
timestamp 1701859473
transform 1 0 2810 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1053_
timestamp 1701859473
transform 1 0 2490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1054_
timestamp 1701859473
transform 1 0 2050 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1055_
timestamp 1701859473
transform 1 0 2710 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1056_
timestamp 1701859473
transform 1 0 2810 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1057_
timestamp 1701859473
transform 1 0 2650 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1058_
timestamp 1701859473
transform 1 0 2490 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1059_
timestamp 1701859473
transform -1 0 2990 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1060_
timestamp 1701859473
transform 1 0 3110 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1061_
timestamp 1701859473
transform 1 0 4890 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1062_
timestamp 1701859473
transform -1 0 2570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1063_
timestamp 1701859473
transform 1 0 2550 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1064_
timestamp 1701859473
transform -1 0 1490 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1065_
timestamp 1701859473
transform -1 0 2250 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1066_
timestamp 1701859473
transform -1 0 1910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1067_
timestamp 1701859473
transform 1 0 2110 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1068_
timestamp 1701859473
transform -1 0 2010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1069_
timestamp 1701859473
transform -1 0 1470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1070_
timestamp 1701859473
transform 1 0 1890 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1071_
timestamp 1701859473
transform 1 0 2050 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1072_
timestamp 1701859473
transform -1 0 1770 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1073_
timestamp 1701859473
transform -1 0 1850 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1074_
timestamp 1701859473
transform -1 0 1750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1075_
timestamp 1701859473
transform -1 0 1630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1076_
timestamp 1701859473
transform 1 0 1490 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1077_
timestamp 1701859473
transform -1 0 1990 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1078_
timestamp 1701859473
transform -1 0 1570 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1079_
timestamp 1701859473
transform -1 0 1850 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1080_
timestamp 1701859473
transform 1 0 1670 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1081_
timestamp 1701859473
transform -1 0 1750 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1082_
timestamp 1701859473
transform 1 0 1950 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1083_
timestamp 1701859473
transform 1 0 1650 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1084_
timestamp 1701859473
transform 1 0 1730 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1085_
timestamp 1701859473
transform -1 0 1750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1086_
timestamp 1701859473
transform -1 0 2570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1087_
timestamp 1701859473
transform 1 0 1590 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1088_
timestamp 1701859473
transform -1 0 1590 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1089_
timestamp 1701859473
transform 1 0 1810 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1090_
timestamp 1701859473
transform 1 0 1850 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1091_
timestamp 1701859473
transform -1 0 2290 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1092_
timestamp 1701859473
transform -1 0 2430 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1093_
timestamp 1701859473
transform -1 0 2390 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1094_
timestamp 1701859473
transform 1 0 2770 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1095_
timestamp 1701859473
transform -1 0 2550 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1096_
timestamp 1701859473
transform 1 0 2910 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1097_
timestamp 1701859473
transform -1 0 3030 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1098_
timestamp 1701859473
transform 1 0 4490 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1099_
timestamp 1701859473
transform 1 0 3250 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1100_
timestamp 1701859473
transform -1 0 610 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1101_
timestamp 1701859473
transform -1 0 1610 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1102_
timestamp 1701859473
transform 1 0 1450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1103_
timestamp 1701859473
transform -1 0 790 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1104_
timestamp 1701859473
transform -1 0 1630 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1105_
timestamp 1701859473
transform 1 0 1210 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1106_
timestamp 1701859473
transform -1 0 1490 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1107_
timestamp 1701859473
transform 1 0 1330 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1108_
timestamp 1701859473
transform -1 0 1310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1109_
timestamp 1701859473
transform -1 0 790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1110_
timestamp 1701859473
transform 1 0 1010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1111_
timestamp 1701859473
transform -1 0 650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1112_
timestamp 1701859473
transform -1 0 490 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1113_
timestamp 1701859473
transform -1 0 1150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1114_
timestamp 1701859473
transform 1 0 870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1115_
timestamp 1701859473
transform -1 0 910 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1116_
timestamp 1701859473
transform -1 0 1970 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1117_
timestamp 1701859473
transform 1 0 1550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1118_
timestamp 1701859473
transform -1 0 2390 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1119_
timestamp 1701859473
transform -1 0 1990 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1120_
timestamp 1701859473
transform -1 0 1850 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1121_
timestamp 1701859473
transform -1 0 2890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1122_
timestamp 1701859473
transform -1 0 2130 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1123_
timestamp 1701859473
transform -1 0 1610 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1124_
timestamp 1701859473
transform -1 0 1690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1125_
timestamp 1701859473
transform -1 0 3730 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1126_
timestamp 1701859473
transform -1 0 1850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1127_
timestamp 1701859473
transform -1 0 1410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1128_
timestamp 1701859473
transform -1 0 1230 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1129_
timestamp 1701859473
transform 1 0 630 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1130_
timestamp 1701859473
transform 1 0 1050 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1131_
timestamp 1701859473
transform 1 0 630 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1132_
timestamp 1701859473
transform -1 0 1370 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1133_
timestamp 1701859473
transform -1 0 970 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1134_
timestamp 1701859473
transform -1 0 810 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1135_
timestamp 1701859473
transform -1 0 1290 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1136_
timestamp 1701859473
transform -1 0 1270 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1137_
timestamp 1701859473
transform 1 0 1090 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1138_
timestamp 1701859473
transform -1 0 1130 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1139_
timestamp 1701859473
transform -1 0 730 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1140_
timestamp 1701859473
transform -1 0 1450 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1141_
timestamp 1701859473
transform -1 0 990 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1142_
timestamp 1701859473
transform -1 0 830 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1143_
timestamp 1701859473
transform 1 0 870 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1144_
timestamp 1701859473
transform 1 0 1270 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1145_
timestamp 1701859473
transform -1 0 2170 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1146_
timestamp 1701859473
transform -1 0 1170 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1147_
timestamp 1701859473
transform -1 0 2030 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1148_
timestamp 1701859473
transform 1 0 2390 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1149_
timestamp 1701859473
transform -1 0 2250 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1150_
timestamp 1701859473
transform -1 0 2750 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1151_
timestamp 1701859473
transform 1 0 2870 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1152_
timestamp 1701859473
transform 1 0 4070 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1153_
timestamp 1701859473
transform -1 0 1770 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1154_
timestamp 1701859473
transform -1 0 450 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1155_
timestamp 1701859473
transform 1 0 2890 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1156_
timestamp 1701859473
transform -1 0 2310 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1157_
timestamp 1701859473
transform 1 0 870 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1158_
timestamp 1701859473
transform -1 0 1510 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1159_
timestamp 1701859473
transform -1 0 1350 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1160_
timestamp 1701859473
transform -1 0 1010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1161_
timestamp 1701859473
transform -1 0 330 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1162_
timestamp 1701859473
transform -1 0 1690 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1163_
timestamp 1701859473
transform 1 0 1810 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1164_
timestamp 1701859473
transform 1 0 1210 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1165_
timestamp 1701859473
transform 1 0 1450 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1166_
timestamp 1701859473
transform -1 0 1530 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1167_
timestamp 1701859473
transform -1 0 1070 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1168_
timestamp 1701859473
transform -1 0 810 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1169_
timestamp 1701859473
transform -1 0 1390 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1170_
timestamp 1701859473
transform -1 0 1130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1171_
timestamp 1701859473
transform 1 0 890 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1172_
timestamp 1701859473
transform 1 0 810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1173_
timestamp 1701859473
transform -1 0 1090 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1174_
timestamp 1701859473
transform -1 0 970 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1175_
timestamp 1701859473
transform 1 0 1350 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1176_
timestamp 1701859473
transform 1 0 1310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1177_
timestamp 1701859473
transform -1 0 1210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1178_
timestamp 1701859473
transform 1 0 1170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1179_
timestamp 1701859473
transform -1 0 1050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1180_
timestamp 1701859473
transform -1 0 950 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1181_
timestamp 1701859473
transform -1 0 930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1182_
timestamp 1701859473
transform -1 0 630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1183_
timestamp 1701859473
transform -1 0 490 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1184_
timestamp 1701859473
transform 1 0 750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1185_
timestamp 1701859473
transform -1 0 1650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1186_
timestamp 1701859473
transform -1 0 1490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1187_
timestamp 1701859473
transform -1 0 1750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1188_
timestamp 1701859473
transform -1 0 1210 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1189_
timestamp 1701859473
transform 1 0 790 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1190_
timestamp 1701859473
transform -1 0 350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1191_
timestamp 1701859473
transform -1 0 670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1192_
timestamp 1701859473
transform -1 0 350 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1193_
timestamp 1701859473
transform -1 0 650 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1194_
timestamp 1701859473
transform -1 0 50 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1195_
timestamp 1701859473
transform 1 0 170 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1196_
timestamp 1701859473
transform 1 0 1390 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1197_
timestamp 1701859473
transform 1 0 190 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1198_
timestamp 1701859473
transform -1 0 490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1199_
timestamp 1701859473
transform 1 0 470 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1200_
timestamp 1701859473
transform 1 0 150 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1201_
timestamp 1701859473
transform -1 0 50 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1202_
timestamp 1701859473
transform -1 0 50 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1203_
timestamp 1701859473
transform -1 0 330 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1204_
timestamp 1701859473
transform 1 0 30 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1205_
timestamp 1701859473
transform 1 0 290 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1206_
timestamp 1701859473
transform -1 0 670 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1207_
timestamp 1701859473
transform 1 0 190 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1208_
timestamp 1701859473
transform 1 0 330 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1209_
timestamp 1701859473
transform 1 0 490 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1210_
timestamp 1701859473
transform 1 0 1610 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1211_
timestamp 1701859473
transform 1 0 1850 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1212_
timestamp 1701859473
transform 1 0 1010 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1213_
timestamp 1701859473
transform 1 0 1430 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1214_
timestamp 1701859473
transform -1 0 1990 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1215_
timestamp 1701859473
transform 1 0 2530 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1216_
timestamp 1701859473
transform 1 0 3670 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1217_
timestamp 1701859473
transform 1 0 2090 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1218_
timestamp 1701859473
transform -1 0 830 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1219_
timestamp 1701859473
transform 1 0 1210 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1220_
timestamp 1701859473
transform 1 0 30 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1221_
timestamp 1701859473
transform -1 0 170 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1222_
timestamp 1701859473
transform 1 0 2430 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1223_
timestamp 1701859473
transform 1 0 1890 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1224_
timestamp 1701859473
transform -1 0 1470 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1225_
timestamp 1701859473
transform -1 0 890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1226_
timestamp 1701859473
transform -1 0 670 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1227_
timestamp 1701859473
transform 1 0 1270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1228_
timestamp 1701859473
transform -1 0 970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1229_
timestamp 1701859473
transform -1 0 50 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1230_
timestamp 1701859473
transform -1 0 210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1231_
timestamp 1701859473
transform 1 0 30 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1232_
timestamp 1701859473
transform -1 0 1630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1233_
timestamp 1701859473
transform -1 0 1330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1234_
timestamp 1701859473
transform 1 0 1030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1235_
timestamp 1701859473
transform -1 0 1170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1236_
timestamp 1701859473
transform -1 0 890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1237_
timestamp 1701859473
transform 1 0 930 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1238_
timestamp 1701859473
transform 1 0 1570 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1239_
timestamp 1701859473
transform -1 0 1350 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1240_
timestamp 1701859473
transform -1 0 1470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1241_
timestamp 1701859473
transform -1 0 810 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1242_
timestamp 1701859473
transform 1 0 730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1243_
timestamp 1701859473
transform -1 0 1050 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1244_
timestamp 1701859473
transform 1 0 890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1245_
timestamp 1701859473
transform -1 0 1610 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1246_
timestamp 1701859473
transform -1 0 1530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1247_
timestamp 1701859473
transform 1 0 1030 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1248_
timestamp 1701859473
transform -1 0 1670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1249_
timestamp 1701859473
transform 1 0 1150 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1250_
timestamp 1701859473
transform -1 0 1410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1251_
timestamp 1701859473
transform -1 0 1310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1252_
timestamp 1701859473
transform -1 0 1010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1253_
timestamp 1701859473
transform -1 0 890 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1254_
timestamp 1701859473
transform -1 0 1170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1255_
timestamp 1701859473
transform -1 0 2370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1256_
timestamp 1701859473
transform -1 0 2230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1257_
timestamp 1701859473
transform -1 0 2730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1258_
timestamp 1701859473
transform -1 0 2070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1259_
timestamp 1701859473
transform -1 0 610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1260_
timestamp 1701859473
transform -1 0 350 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1261_
timestamp 1701859473
transform -1 0 610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1262_
timestamp 1701859473
transform 1 0 710 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1263_
timestamp 1701859473
transform 1 0 730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1264_
timestamp 1701859473
transform -1 0 310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1265_
timestamp 1701859473
transform -1 0 50 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1266_
timestamp 1701859473
transform -1 0 490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1267_
timestamp 1701859473
transform -1 0 330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1268_
timestamp 1701859473
transform 1 0 430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1269_
timestamp 1701859473
transform -1 0 510 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1270_
timestamp 1701859473
transform -1 0 350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1271_
timestamp 1701859473
transform 1 0 190 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1272_
timestamp 1701859473
transform 1 0 210 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1273_
timestamp 1701859473
transform 1 0 190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1274_
timestamp 1701859473
transform 1 0 490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1275_
timestamp 1701859473
transform 1 0 490 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1276_
timestamp 1701859473
transform -1 0 210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1277_
timestamp 1701859473
transform 1 0 30 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1278_
timestamp 1701859473
transform -1 0 210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1279_
timestamp 1701859473
transform -1 0 350 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1280_
timestamp 1701859473
transform -1 0 50 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1281_
timestamp 1701859473
transform 1 0 30 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1282_
timestamp 1701859473
transform 1 0 170 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1283_
timestamp 1701859473
transform -1 0 790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1284_
timestamp 1701859473
transform 1 0 330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1285_
timestamp 1701859473
transform 1 0 30 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1286_
timestamp 1701859473
transform 1 0 630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1287_
timestamp 1701859473
transform -1 0 670 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1288_
timestamp 1701859473
transform 1 0 490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1289_
timestamp 1701859473
transform 1 0 330 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1290_
timestamp 1701859473
transform 1 0 490 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1291_
timestamp 1701859473
transform 1 0 2350 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1292_
timestamp 1701859473
transform 1 0 2190 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1293_
timestamp 1701859473
transform -1 0 2930 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1294_
timestamp 1701859473
transform -1 0 3050 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1295_
timestamp 1701859473
transform 1 0 2690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1296_
timestamp 1701859473
transform -1 0 2950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1297_
timestamp 1701859473
transform -1 0 1110 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1298_
timestamp 1701859473
transform 1 0 790 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1299_
timestamp 1701859473
transform 1 0 30 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1300_
timestamp 1701859473
transform 1 0 30 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1301_
timestamp 1701859473
transform -1 0 170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1302_
timestamp 1701859473
transform 1 0 2910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1303_
timestamp 1701859473
transform -1 0 2390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1304_
timestamp 1701859473
transform -1 0 2610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1305_
timestamp 1701859473
transform 1 0 2050 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1306_
timestamp 1701859473
transform 1 0 1930 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1307_
timestamp 1701859473
transform -1 0 2230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1308_
timestamp 1701859473
transform -1 0 1930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1309_
timestamp 1701859473
transform 1 0 3130 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1310_
timestamp 1701859473
transform -1 0 2610 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1311_
timestamp 1701859473
transform -1 0 1750 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1312_
timestamp 1701859473
transform -1 0 1630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1313_
timestamp 1701859473
transform 1 0 1190 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1314_
timestamp 1701859473
transform -1 0 1470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1315_
timestamp 1701859473
transform -1 0 1790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1316_
timestamp 1701859473
transform -1 0 2070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1317_
timestamp 1701859473
transform 1 0 1030 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1318_
timestamp 1701859473
transform -1 0 1170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1319_
timestamp 1701859473
transform -1 0 1010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1320_
timestamp 1701859473
transform -1 0 1230 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1321_
timestamp 1701859473
transform -1 0 1310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1322_
timestamp 1701859473
transform 1 0 790 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1323_
timestamp 1701859473
transform 1 0 630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1324_
timestamp 1701859473
transform -1 0 330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1325_
timestamp 1701859473
transform -1 0 190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1326_
timestamp 1701859473
transform 1 0 1490 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1327_
timestamp 1701859473
transform -1 0 1370 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1328_
timestamp 1701859473
transform 1 0 1030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1329_
timestamp 1701859473
transform 1 0 1070 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1330_
timestamp 1701859473
transform 1 0 1330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1331_
timestamp 1701859473
transform 1 0 1170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1332_
timestamp 1701859473
transform 1 0 1750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1333_
timestamp 1701859473
transform 1 0 2710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1334_
timestamp 1701859473
transform 1 0 1990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1335_
timestamp 1701859473
transform -1 0 1650 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1336_
timestamp 1701859473
transform -1 0 1710 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1337_
timestamp 1701859473
transform 1 0 1330 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1338_
timestamp 1701859473
transform 1 0 1290 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1339_
timestamp 1701859473
transform -1 0 770 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1340_
timestamp 1701859473
transform 1 0 1450 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1341_
timestamp 1701859473
transform 1 0 1570 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1342_
timestamp 1701859473
transform -1 0 1670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1343_
timestamp 1701859473
transform -1 0 1810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1344_
timestamp 1701859473
transform 1 0 1510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1345_
timestamp 1701859473
transform -1 0 1490 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1346_
timestamp 1701859473
transform 1 0 1910 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1347_
timestamp 1701859473
transform -1 0 2110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1348_
timestamp 1701859473
transform -1 0 1630 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1349_
timestamp 1701859473
transform -1 0 1670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1350_
timestamp 1701859473
transform -1 0 890 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1351_
timestamp 1701859473
transform 1 0 1750 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1352_
timestamp 1701859473
transform -1 0 1390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1353_
timestamp 1701859473
transform -1 0 1230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1354_
timestamp 1701859473
transform -1 0 930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1355_
timestamp 1701859473
transform -1 0 1210 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1356_
timestamp 1701859473
transform -1 0 1030 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1357_
timestamp 1701859473
transform -1 0 1090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1358_
timestamp 1701859473
transform -1 0 650 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1359_
timestamp 1701859473
transform -1 0 350 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1360_
timestamp 1701859473
transform -1 0 590 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1361_
timestamp 1701859473
transform -1 0 450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1362_
timestamp 1701859473
transform -1 0 810 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1363_
timestamp 1701859473
transform -1 0 770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1364_
timestamp 1701859473
transform -1 0 510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1365_
timestamp 1701859473
transform 1 0 170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1366_
timestamp 1701859473
transform -1 0 890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1367_
timestamp 1701859473
transform -1 0 510 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1368_
timestamp 1701859473
transform -1 0 350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1369_
timestamp 1701859473
transform 1 0 190 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1370_
timestamp 1701859473
transform -1 0 190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1371_
timestamp 1701859473
transform -1 0 190 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1372_
timestamp 1701859473
transform 1 0 30 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1373_
timestamp 1701859473
transform -1 0 50 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1374_
timestamp 1701859473
transform 1 0 30 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1375_
timestamp 1701859473
transform 1 0 30 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1376_
timestamp 1701859473
transform 1 0 190 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1377_
timestamp 1701859473
transform 1 0 490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1378_
timestamp 1701859473
transform 1 0 330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1379_
timestamp 1701859473
transform 1 0 30 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1380_
timestamp 1701859473
transform 1 0 490 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1381_
timestamp 1701859473
transform 1 0 630 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1382_
timestamp 1701859473
transform 1 0 650 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1383_
timestamp 1701859473
transform 1 0 930 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1384_
timestamp 1701859473
transform -1 0 370 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1385_
timestamp 1701859473
transform 1 0 30 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1386_
timestamp 1701859473
transform -1 0 430 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1387_
timestamp 1701859473
transform 1 0 2170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1388_
timestamp 1701859473
transform 1 0 3150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1389_
timestamp 1701859473
transform -1 0 3050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1390_
timestamp 1701859473
transform 1 0 3250 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1391_
timestamp 1701859473
transform 1 0 3310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1392_
timestamp 1701859473
transform -1 0 3470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1393_
timestamp 1701859473
transform -1 0 4550 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1394_
timestamp 1701859473
transform -1 0 2310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1395_
timestamp 1701859473
transform 1 0 2010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1396_
timestamp 1701859473
transform 1 0 2390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1397_
timestamp 1701859473
transform 1 0 190 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1398_
timestamp 1701859473
transform 1 0 350 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1399_
timestamp 1701859473
transform -1 0 770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1400_
timestamp 1701859473
transform 1 0 30 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1401_
timestamp 1701859473
transform 1 0 30 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1402_
timestamp 1701859473
transform 1 0 130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1403_
timestamp 1701859473
transform 1 0 1770 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1404_
timestamp 1701859473
transform 1 0 2790 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1405_
timestamp 1701859473
transform 1 0 2530 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1406_
timestamp 1701859473
transform -1 0 3010 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1407_
timestamp 1701859473
transform -1 0 3610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1408_
timestamp 1701859473
transform 1 0 3050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1409_
timestamp 1701859473
transform -1 0 3370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1410_
timestamp 1701859473
transform 1 0 3190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1411_
timestamp 1701859473
transform -1 0 2450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1412_
timestamp 1701859473
transform 1 0 2750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1413_
timestamp 1701859473
transform 1 0 2730 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1414_
timestamp 1701859473
transform -1 0 2250 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1415_
timestamp 1701859473
transform 1 0 1450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1416_
timestamp 1701859473
transform 1 0 1850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1417_
timestamp 1701859473
transform -1 0 2150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1418_
timestamp 1701859473
transform 1 0 2370 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1419_
timestamp 1701859473
transform 1 0 2570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1420_
timestamp 1701859473
transform -1 0 1630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1421_
timestamp 1701859473
transform 1 0 1850 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1422_
timestamp 1701859473
transform -1 0 2450 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1423_
timestamp 1701859473
transform 1 0 1990 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1424_
timestamp 1701859473
transform -1 0 2490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1425_
timestamp 1701859473
transform -1 0 2090 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1426_
timestamp 1701859473
transform -1 0 2310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1427_
timestamp 1701859473
transform -1 0 2290 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1428_
timestamp 1701859473
transform 1 0 2130 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1429_
timestamp 1701859473
transform -1 0 1530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1430_
timestamp 1701859473
transform -1 0 1090 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1431_
timestamp 1701859473
transform -1 0 950 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1432_
timestamp 1701859473
transform 1 0 3050 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1433_
timestamp 1701859473
transform 1 0 3310 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1434_
timestamp 1701859473
transform -1 0 3050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1435_
timestamp 1701859473
transform 1 0 3430 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1436_
timestamp 1701859473
transform -1 0 2930 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1437_
timestamp 1701859473
transform -1 0 2890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1438_
timestamp 1701859473
transform -1 0 3070 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1439_
timestamp 1701859473
transform 1 0 3750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1440_
timestamp 1701859473
transform 1 0 3490 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1441_
timestamp 1701859473
transform -1 0 3370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1442_
timestamp 1701859473
transform -1 0 2910 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1443_
timestamp 1701859473
transform 1 0 2670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1444_
timestamp 1701859473
transform 1 0 2510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1445_
timestamp 1701859473
transform 1 0 2350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1446_
timestamp 1701859473
transform -1 0 4270 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1447_
timestamp 1701859473
transform 1 0 2570 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1448_
timestamp 1701859473
transform 1 0 1950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1449_
timestamp 1701859473
transform 1 0 1930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1450_
timestamp 1701859473
transform 1 0 2030 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1451_
timestamp 1701859473
transform -1 0 2430 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1452_
timestamp 1701859473
transform -1 0 2110 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1453_
timestamp 1701859473
transform -1 0 2730 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1454_
timestamp 1701859473
transform -1 0 2310 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1455_
timestamp 1701859473
transform 1 0 2170 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1456_
timestamp 1701859473
transform 1 0 1650 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1457_
timestamp 1701859473
transform -1 0 1390 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1458_
timestamp 1701859473
transform -1 0 1250 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1459_
timestamp 1701859473
transform -1 0 770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1460_
timestamp 1701859473
transform -1 0 1350 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1461_
timestamp 1701859473
transform -1 0 1190 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1462_
timestamp 1701859473
transform -1 0 2410 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1463_
timestamp 1701859473
transform 1 0 1790 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1464_
timestamp 1701859473
transform -1 0 1510 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1465_
timestamp 1701859473
transform 1 0 2250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1466_
timestamp 1701859473
transform -1 0 690 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1467_
timestamp 1701859473
transform -1 0 370 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1468_
timestamp 1701859473
transform -1 0 1390 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1469_
timestamp 1701859473
transform 1 0 910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1470_
timestamp 1701859473
transform -1 0 850 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1471_
timestamp 1701859473
transform -1 0 530 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1472_
timestamp 1701859473
transform 1 0 190 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1473_
timestamp 1701859473
transform -1 0 470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1474_
timestamp 1701859473
transform -1 0 310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1475_
timestamp 1701859473
transform -1 0 510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1476_
timestamp 1701859473
transform -1 0 350 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1477_
timestamp 1701859473
transform -1 0 50 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1478_
timestamp 1701859473
transform 1 0 150 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1479_
timestamp 1701859473
transform -1 0 50 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1480_
timestamp 1701859473
transform 1 0 190 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1481_
timestamp 1701859473
transform -1 0 610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1482_
timestamp 1701859473
transform 1 0 510 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1483_
timestamp 1701859473
transform -1 0 770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1484_
timestamp 1701859473
transform 1 0 590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1485_
timestamp 1701859473
transform -1 0 470 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1486_
timestamp 1701859473
transform 1 0 290 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1487_
timestamp 1701859473
transform 1 0 650 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1488_
timestamp 1701859473
transform -1 0 3130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1489_
timestamp 1701859473
transform -1 0 3850 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1490_
timestamp 1701859473
transform 1 0 4390 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1491_
timestamp 1701859473
transform 1 0 3250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1492_
timestamp 1701859473
transform 1 0 3370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1493_
timestamp 1701859473
transform -1 0 650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1494_
timestamp 1701859473
transform 1 0 590 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1495_
timestamp 1701859473
transform -1 0 2250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1496_
timestamp 1701859473
transform 1 0 2830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1497_
timestamp 1701859473
transform -1 0 1150 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1498_
timestamp 1701859473
transform 1 0 970 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1499_
timestamp 1701859473
transform 1 0 2730 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1500_
timestamp 1701859473
transform -1 0 3490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1501_
timestamp 1701859473
transform -1 0 3830 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1502_
timestamp 1701859473
transform 1 0 3690 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1503_
timestamp 1701859473
transform -1 0 3970 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1504_
timestamp 1701859473
transform -1 0 3650 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1505_
timestamp 1701859473
transform -1 0 3510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1506_
timestamp 1701859473
transform -1 0 4890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1507_
timestamp 1701859473
transform 1 0 3910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1508_
timestamp 1701859473
transform -1 0 3890 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1509_
timestamp 1701859473
transform -1 0 3570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1510_
timestamp 1701859473
transform -1 0 3210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1511_
timestamp 1701859473
transform 1 0 3150 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1512_
timestamp 1701859473
transform -1 0 3270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1513_
timestamp 1701859473
transform 1 0 3690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1514_
timestamp 1701859473
transform -1 0 3610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1515_
timestamp 1701859473
transform -1 0 3330 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1516_
timestamp 1701859473
transform -1 0 2950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1517_
timestamp 1701859473
transform 1 0 2790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1518_
timestamp 1701859473
transform -1 0 2670 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1519_
timestamp 1701859473
transform 1 0 2590 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1520_
timestamp 1701859473
transform 1 0 3090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1521_
timestamp 1701859473
transform -1 0 3410 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1522_
timestamp 1701859473
transform 1 0 3490 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1523_
timestamp 1701859473
transform 1 0 3230 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1524_
timestamp 1701859473
transform 1 0 1810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1525_
timestamp 1701859473
transform 1 0 1930 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1526_
timestamp 1701859473
transform 1 0 4130 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1527_
timestamp 1701859473
transform -1 0 4390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1528_
timestamp 1701859473
transform 1 0 4210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1529_
timestamp 1701859473
transform 1 0 3910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1530_
timestamp 1701859473
transform -1 0 4070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1531_
timestamp 1701859473
transform 1 0 4290 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1532_
timestamp 1701859473
transform -1 0 4730 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1533_
timestamp 1701859473
transform 1 0 3730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1534_
timestamp 1701859473
transform -1 0 4170 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1535_
timestamp 1701859473
transform -1 0 4010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1536_
timestamp 1701859473
transform -1 0 4150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1537_
timestamp 1701859473
transform -1 0 4170 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1538_
timestamp 1701859473
transform -1 0 4030 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1539_
timestamp 1701859473
transform -1 0 3870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1540_
timestamp 1701859473
transform -1 0 3790 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1541_
timestamp 1701859473
transform 1 0 3650 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1542_
timestamp 1701859473
transform 1 0 2530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1543_
timestamp 1701859473
transform 1 0 2670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1544_
timestamp 1701859473
transform 1 0 4350 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1545_
timestamp 1701859473
transform -1 0 4210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1546_
timestamp 1701859473
transform 1 0 3910 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1547_
timestamp 1701859473
transform 1 0 4490 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1548_
timestamp 1701859473
transform -1 0 3390 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1549_
timestamp 1701859473
transform -1 0 4070 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1550_
timestamp 1701859473
transform -1 0 3270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1551_
timestamp 1701859473
transform 1 0 1070 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1552_
timestamp 1701859473
transform -1 0 1230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1553_
timestamp 1701859473
transform 1 0 3870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1554_
timestamp 1701859473
transform -1 0 3530 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1555_
timestamp 1701859473
transform 1 0 2230 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1556_
timestamp 1701859473
transform -1 0 3110 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1557_
timestamp 1701859473
transform 1 0 2930 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1558_
timestamp 1701859473
transform 1 0 3090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1559_
timestamp 1701859473
transform 1 0 3410 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1560_
timestamp 1701859473
transform 1 0 2630 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1561_
timestamp 1701859473
transform -1 0 3370 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1562_
timestamp 1701859473
transform -1 0 3210 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1563_
timestamp 1701859473
transform -1 0 3050 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1564_
timestamp 1701859473
transform -1 0 2970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1565_
timestamp 1701859473
transform -1 0 2870 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1566_
timestamp 1701859473
transform -1 0 3210 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1567_
timestamp 1701859473
transform 1 0 3510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1568_
timestamp 1701859473
transform 1 0 4110 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1569_
timestamp 1701859473
transform -1 0 3930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1570_
timestamp 1701859473
transform -1 0 4590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1571_
timestamp 1701859473
transform -1 0 3250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1572_
timestamp 1701859473
transform 1 0 3710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1573_
timestamp 1701859473
transform 1 0 4710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1574_
timestamp 1701859473
transform -1 0 3730 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1575_
timestamp 1701859473
transform -1 0 3570 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1576_
timestamp 1701859473
transform 1 0 3890 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1577_
timestamp 1701859473
transform 1 0 4190 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1578_
timestamp 1701859473
transform 1 0 4050 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1579_
timestamp 1701859473
transform 1 0 3990 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1580_
timestamp 1701859473
transform 1 0 4910 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1581_
timestamp 1701859473
transform -1 0 4290 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1582_
timestamp 1701859473
transform -1 0 4830 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1583_
timestamp 1701859473
transform 1 0 4990 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1584_
timestamp 1701859473
transform 1 0 4670 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1585_
timestamp 1701859473
transform 1 0 4950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1586_
timestamp 1701859473
transform 1 0 5730 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1587_
timestamp 1701859473
transform 1 0 5330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1588_
timestamp 1701859473
transform -1 0 5330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1589_
timestamp 1701859473
transform 1 0 5030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1590_
timestamp 1701859473
transform 1 0 5570 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1591_
timestamp 1701859473
transform -1 0 4850 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1592_
timestamp 1701859473
transform 1 0 4950 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1593_
timestamp 1701859473
transform -1 0 5130 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1594_
timestamp 1701859473
transform -1 0 5430 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1595_
timestamp 1701859473
transform -1 0 4810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1596_
timestamp 1701859473
transform -1 0 4590 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1597_
timestamp 1701859473
transform 1 0 4410 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1598_
timestamp 1701859473
transform -1 0 5070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1599_
timestamp 1701859473
transform 1 0 5030 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1600_
timestamp 1701859473
transform -1 0 4930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1601_
timestamp 1701859473
transform -1 0 5270 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1602_
timestamp 1701859473
transform 1 0 4750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1603_
timestamp 1701859473
transform 1 0 5670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1604_
timestamp 1701859473
transform 1 0 4190 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1605_
timestamp 1701859473
transform 1 0 4330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1606_
timestamp 1701859473
transform 1 0 4270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1607_
timestamp 1701859473
transform 1 0 4310 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1608_
timestamp 1701859473
transform 1 0 4390 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1609_
timestamp 1701859473
transform -1 0 4710 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1610_
timestamp 1701859473
transform -1 0 4550 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1611_
timestamp 1701859473
transform -1 0 4550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1612_
timestamp 1701859473
transform 1 0 4390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1613_
timestamp 1701859473
transform 1 0 4650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1614_
timestamp 1701859473
transform -1 0 4630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1615_
timestamp 1701859473
transform 1 0 4350 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1616_
timestamp 1701859473
transform 1 0 4510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1617_
timestamp 1701859473
transform 1 0 4470 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1618_
timestamp 1701859473
transform 1 0 5890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1619_
timestamp 1701859473
transform 1 0 6110 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1620_
timestamp 1701859473
transform 1 0 4630 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1621_
timestamp 1701859473
transform -1 0 4490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1622_
timestamp 1701859473
transform 1 0 4770 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1623_
timestamp 1701859473
transform -1 0 5550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1624_
timestamp 1701859473
transform -1 0 5410 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1625_
timestamp 1701859473
transform 1 0 4650 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1626_
timestamp 1701859473
transform -1 0 5110 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1627_
timestamp 1701859473
transform 1 0 5970 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1628_
timestamp 1701859473
transform -1 0 4950 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1629_
timestamp 1701859473
transform 1 0 4770 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1630_
timestamp 1701859473
transform -1 0 5570 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1631_
timestamp 1701859473
transform 1 0 5070 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1632_
timestamp 1701859473
transform -1 0 4970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1633_
timestamp 1701859473
transform -1 0 4810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1634_
timestamp 1701859473
transform -1 0 2410 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1635_
timestamp 1701859473
transform 1 0 2790 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1636_
timestamp 1701859473
transform -1 0 4490 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1637_
timestamp 1701859473
transform -1 0 4650 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1638_
timestamp 1701859473
transform -1 0 4330 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1639_
timestamp 1701859473
transform -1 0 4910 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1640_
timestamp 1701859473
transform -1 0 4810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1641_
timestamp 1701859473
transform -1 0 4870 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1642_
timestamp 1701859473
transform -1 0 4730 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1643_
timestamp 1701859473
transform 1 0 5410 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1644_
timestamp 1701859473
transform 1 0 4990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1645_
timestamp 1701859473
transform -1 0 5710 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1646_
timestamp 1701859473
transform 1 0 5230 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1647_
timestamp 1701859473
transform 1 0 5190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1648_
timestamp 1701859473
transform 1 0 5610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1649_
timestamp 1701859473
transform 1 0 5190 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1650_
timestamp 1701859473
transform 1 0 5790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1651_
timestamp 1701859473
transform 1 0 5650 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1652_
timestamp 1701859473
transform 1 0 5190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1653_
timestamp 1701859473
transform 1 0 5270 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1654_
timestamp 1701859473
transform -1 0 5850 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1655_
timestamp 1701859473
transform 1 0 5110 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1656_
timestamp 1701859473
transform 1 0 5410 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1657_
timestamp 1701859473
transform 1 0 4470 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1658_
timestamp 1701859473
transform 1 0 5170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1659_
timestamp 1701859473
transform 1 0 5690 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1660_
timestamp 1701859473
transform -1 0 5190 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1661_
timestamp 1701859473
transform -1 0 5330 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1662_
timestamp 1701859473
transform 1 0 5790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1663_
timestamp 1701859473
transform 1 0 6110 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1664_
timestamp 1701859473
transform -1 0 5770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1665_
timestamp 1701859473
transform -1 0 5570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1666_
timestamp 1701859473
transform 1 0 5530 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1667_
timestamp 1701859473
transform 1 0 5610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1668_
timestamp 1701859473
transform -1 0 6250 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1669_
timestamp 1701859473
transform 1 0 5830 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1670_
timestamp 1701859473
transform -1 0 5470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1671_
timestamp 1701859473
transform -1 0 5970 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1672_
timestamp 1701859473
transform 1 0 5930 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1673_
timestamp 1701859473
transform 1 0 3990 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1674_
timestamp 1701859473
transform -1 0 4170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1675_
timestamp 1701859473
transform 1 0 5930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1676_
timestamp 1701859473
transform 1 0 6210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1677_
timestamp 1701859473
transform -1 0 6110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1678_
timestamp 1701859473
transform -1 0 6090 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1679_
timestamp 1701859473
transform 1 0 5850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1680_
timestamp 1701859473
transform 1 0 6250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1681_
timestamp 1701859473
transform 1 0 6130 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1682_
timestamp 1701859473
transform 1 0 5990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1683_
timestamp 1701859473
transform -1 0 5750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1684_
timestamp 1701859473
transform 1 0 5890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1685_
timestamp 1701859473
transform 1 0 5810 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1686_
timestamp 1701859473
transform -1 0 5470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1687_
timestamp 1701859473
transform -1 0 6030 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1688_
timestamp 1701859473
transform 1 0 6010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1689_
timestamp 1701859473
transform -1 0 6290 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1690_
timestamp 1701859473
transform 1 0 6110 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1691_
timestamp 1701859473
transform -1 0 5330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1692_
timestamp 1701859473
transform -1 0 5430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1693_
timestamp 1701859473
transform 1 0 5250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1694_
timestamp 1701859473
transform -1 0 5990 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1695_
timestamp 1701859473
transform -1 0 5510 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1696_
timestamp 1701859473
transform -1 0 5370 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1697_
timestamp 1701859473
transform 1 0 5330 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1698_
timestamp 1701859473
transform 1 0 5710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1699_
timestamp 1701859473
transform 1 0 5590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1700_
timestamp 1701859473
transform -1 0 5290 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1701_
timestamp 1701859473
transform 1 0 5270 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1702_
timestamp 1701859473
transform 1 0 5990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1703_
timestamp 1701859473
transform -1 0 5170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1704_
timestamp 1701859473
transform 1 0 4850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1705_
timestamp 1701859473
transform -1 0 5310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1706_
timestamp 1701859473
transform -1 0 5450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1707_
timestamp 1701859473
transform 1 0 5430 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1708_
timestamp 1701859473
transform 1 0 6170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1709_
timestamp 1701859473
transform 1 0 6270 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1710_
timestamp 1701859473
transform 1 0 5610 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1711_
timestamp 1701859473
transform 1 0 5410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1712_
timestamp 1701859473
transform -1 0 5050 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1713_
timestamp 1701859473
transform 1 0 4730 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1714_
timestamp 1701859473
transform 1 0 4610 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1715_
timestamp 1701859473
transform -1 0 4510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1716_
timestamp 1701859473
transform 1 0 4630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1717_
timestamp 1701859473
transform -1 0 4950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1718_
timestamp 1701859473
transform 1 0 5070 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1719_
timestamp 1701859473
transform 1 0 5250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1720_
timestamp 1701859473
transform -1 0 5470 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1721_
timestamp 1701859473
transform 1 0 5790 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1722_
timestamp 1701859473
transform 1 0 4670 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1723_
timestamp 1701859473
transform 1 0 4110 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1724_
timestamp 1701859473
transform 1 0 4790 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1725_
timestamp 1701859473
transform 1 0 4930 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1726_
timestamp 1701859473
transform 1 0 5090 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1727_
timestamp 1701859473
transform -1 0 5710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1728_
timestamp 1701859473
transform 1 0 5390 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1729_
timestamp 1701859473
transform 1 0 5210 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1730_
timestamp 1701859473
transform 1 0 5530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1731_
timestamp 1701859473
transform 1 0 5990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1732_
timestamp 1701859473
transform 1 0 5850 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1733_
timestamp 1701859473
transform 1 0 5770 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1734_
timestamp 1701859473
transform -1 0 6290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1735_
timestamp 1701859473
transform -1 0 6290 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1736_
timestamp 1701859473
transform -1 0 6050 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1737_
timestamp 1701859473
transform 1 0 5910 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1738_
timestamp 1701859473
transform 1 0 6130 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1739_
timestamp 1701859473
transform -1 0 6150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1740_
timestamp 1701859473
transform 1 0 6170 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1741_
timestamp 1701859473
transform 1 0 6290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1742_
timestamp 1701859473
transform 1 0 6290 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1743_
timestamp 1701859473
transform 1 0 5890 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1744_
timestamp 1701859473
transform 1 0 5610 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1745_
timestamp 1701859473
transform 1 0 5590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1746_
timestamp 1701859473
transform 1 0 6250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1747_
timestamp 1701859473
transform 1 0 6090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1748_
timestamp 1701859473
transform -1 0 6290 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1749_
timestamp 1701859473
transform 1 0 4750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1750_
timestamp 1701859473
transform -1 0 4070 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1751_
timestamp 1701859473
transform 1 0 4330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1752_
timestamp 1701859473
transform 1 0 3910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1753_
timestamp 1701859473
transform 1 0 4230 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1754_
timestamp 1701859473
transform 1 0 4350 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1755_
timestamp 1701859473
transform 1 0 4690 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1756_
timestamp 1701859473
transform -1 0 4210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1757_
timestamp 1701859473
transform 1 0 5470 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1758_
timestamp 1701859473
transform 1 0 6030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1759_
timestamp 1701859473
transform 1 0 5630 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1760_
timestamp 1701859473
transform 1 0 6130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1761_
timestamp 1701859473
transform 1 0 5890 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1762_
timestamp 1701859473
transform 1 0 6010 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1763_
timestamp 1701859473
transform 1 0 6150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_1__1764_
timestamp 1701859473
transform -1 0 6210 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1765_
timestamp 1701859473
transform 1 0 6010 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1766_
timestamp 1701859473
transform -1 0 6130 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1767_
timestamp 1701859473
transform -1 0 6290 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1768_
timestamp 1701859473
transform -1 0 6330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1769_
timestamp 1701859473
transform -1 0 6150 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1770_
timestamp 1701859473
transform 1 0 5330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1771_
timestamp 1701859473
transform -1 0 5750 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1772_
timestamp 1701859473
transform 1 0 5570 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1773_
timestamp 1701859473
transform -1 0 6270 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1774_
timestamp 1701859473
transform -1 0 6050 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1775_
timestamp 1701859473
transform -1 0 5990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1776_
timestamp 1701859473
transform -1 0 5890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1777_
timestamp 1701859473
transform -1 0 4890 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1778_
timestamp 1701859473
transform 1 0 3470 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1779_
timestamp 1701859473
transform 1 0 4510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1780_
timestamp 1701859473
transform 1 0 4390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1781_
timestamp 1701859473
transform 1 0 4630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1782_
timestamp 1701859473
transform -1 0 4530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1783_
timestamp 1701859473
transform 1 0 4930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1784_
timestamp 1701859473
transform -1 0 5010 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1785_
timestamp 1701859473
transform 1 0 5130 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1786_
timestamp 1701859473
transform 1 0 5230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1787_
timestamp 1701859473
transform -1 0 5550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1788_
timestamp 1701859473
transform 1 0 5650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1789_
timestamp 1701859473
transform -1 0 5830 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1790_
timestamp 1701859473
transform -1 0 5470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1791_
timestamp 1701859473
transform -1 0 5830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1792_
timestamp 1701859473
transform 1 0 5390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1793_
timestamp 1701859473
transform -1 0 5090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1794_
timestamp 1701859473
transform -1 0 4530 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1795_
timestamp 1701859473
transform -1 0 4550 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1796_
timestamp 1701859473
transform -1 0 5030 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1797_
timestamp 1701859473
transform 1 0 5370 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1798_
timestamp 1701859473
transform -1 0 5490 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1799_
timestamp 1701859473
transform -1 0 5230 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1800_
timestamp 1701859473
transform 1 0 5190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1801_
timestamp 1701859473
transform -1 0 5550 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1802_
timestamp 1701859473
transform -1 0 3470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1803_
timestamp 1701859473
transform -1 0 4490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1804_
timestamp 1701859473
transform -1 0 4330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1805_
timestamp 1701859473
transform -1 0 4090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1806_
timestamp 1701859473
transform 1 0 3910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1807_
timestamp 1701859473
transform -1 0 3370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1808_
timestamp 1701859473
transform 1 0 4190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1809_
timestamp 1701859473
transform 1 0 4050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1810_
timestamp 1701859473
transform -1 0 3610 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1811_
timestamp 1701859473
transform -1 0 4330 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1812_
timestamp 1701859473
transform 1 0 4170 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1813_
timestamp 1701859473
transform 1 0 3890 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1814_
timestamp 1701859473
transform -1 0 4190 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1815_
timestamp 1701859473
transform 1 0 4010 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1816_
timestamp 1701859473
transform -1 0 4270 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1817_
timestamp 1701859473
transform 1 0 3870 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1818_
timestamp 1701859473
transform 1 0 3850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1819_
timestamp 1701859473
transform 1 0 3550 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1820_
timestamp 1701859473
transform -1 0 3770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1821_
timestamp 1701859473
transform 1 0 3610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1822_
timestamp 1701859473
transform -1 0 4070 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1823_
timestamp 1701859473
transform 1 0 4030 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1824_
timestamp 1701859473
transform 1 0 4010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1825_
timestamp 1701859473
transform 1 0 3130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1826_
timestamp 1701859473
transform 1 0 2850 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1827_
timestamp 1701859473
transform -1 0 2690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1828_
timestamp 1701859473
transform 1 0 2810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1829_
timestamp 1701859473
transform -1 0 3230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1830_
timestamp 1701859473
transform -1 0 2790 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1831_
timestamp 1701859473
transform -1 0 2710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1832_
timestamp 1701859473
transform 1 0 3210 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1833_
timestamp 1701859473
transform -1 0 3270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1834_
timestamp 1701859473
transform -1 0 4010 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1835_
timestamp 1701859473
transform 1 0 3590 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1836_
timestamp 1701859473
transform -1 0 3270 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1837_
timestamp 1701859473
transform -1 0 3410 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1838_
timestamp 1701859473
transform -1 0 3010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1839_
timestamp 1701859473
transform 1 0 2850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1840_
timestamp 1701859473
transform 1 0 2330 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1841_
timestamp 1701859473
transform 1 0 2070 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1842_
timestamp 1701859473
transform -1 0 2030 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1843_
timestamp 1701859473
transform -1 0 2170 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1844_
timestamp 1701859473
transform -1 0 2510 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1845_
timestamp 1701859473
transform -1 0 2630 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1846_
timestamp 1701859473
transform -1 0 2330 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1847_
timestamp 1701859473
transform -1 0 2450 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1848_
timestamp 1701859473
transform 1 0 2790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1849_
timestamp 1701859473
transform 1 0 2650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1911_
timestamp 1701859473
transform 1 0 6250 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1912_
timestamp 1701859473
transform 1 0 2170 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1913_
timestamp 1701859473
transform 1 0 2090 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1914_
timestamp 1701859473
transform 1 0 3630 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1915_
timestamp 1701859473
transform 1 0 3770 0 1 5470
box -12 -8 32 272
use FILL  FILL_1__1916_
timestamp 1701859473
transform 1 0 6270 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1917_
timestamp 1701859473
transform 1 0 6130 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1918_
timestamp 1701859473
transform 1 0 5830 0 1 5990
box -12 -8 32 272
use FILL  FILL_1__1919_
timestamp 1701859473
transform -1 0 5690 0 1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert0
timestamp 1701859473
transform 1 0 4750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert1
timestamp 1701859473
transform -1 0 4370 0 1 270
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert2
timestamp 1701859473
transform -1 0 4230 0 -1 270
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert3
timestamp 1701859473
transform 1 0 5350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert4
timestamp 1701859473
transform 1 0 5510 0 1 270
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert12
timestamp 1701859473
transform 1 0 2070 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert13
timestamp 1701859473
transform 1 0 2210 0 1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert14
timestamp 1701859473
transform 1 0 1310 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert15
timestamp 1701859473
transform -1 0 1890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert16
timestamp 1701859473
transform -1 0 3550 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert17
timestamp 1701859473
transform 1 0 3070 0 1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert18
timestamp 1701859473
transform -1 0 3370 0 1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert19
timestamp 1701859473
transform -1 0 2990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert20
timestamp 1701859473
transform 1 0 3910 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert21
timestamp 1701859473
transform -1 0 4070 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert22
timestamp 1701859473
transform -1 0 5630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert23
timestamp 1701859473
transform -1 0 3590 0 1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert24
timestamp 1701859473
transform 1 0 4070 0 1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert25
timestamp 1701859473
transform 1 0 4890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert5
timestamp 1701859473
transform 1 0 4910 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert6
timestamp 1701859473
transform 1 0 4910 0 1 1830
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert7
timestamp 1701859473
transform -1 0 4110 0 1 270
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert8
timestamp 1701859473
transform -1 0 3670 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert9
timestamp 1701859473
transform -1 0 3430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert10
timestamp 1701859473
transform 1 0 4650 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert11
timestamp 1701859473
transform -1 0 4690 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__922_
timestamp 1701859473
transform -1 0 4110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__923_
timestamp 1701859473
transform 1 0 4210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__924_
timestamp 1701859473
transform -1 0 5750 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__925_
timestamp 1701859473
transform -1 0 5850 0 1 790
box -12 -8 32 272
use FILL  FILL_2__926_
timestamp 1701859473
transform -1 0 6150 0 1 790
box -12 -8 32 272
use FILL  FILL_2__927_
timestamp 1701859473
transform -1 0 3770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__928_
timestamp 1701859473
transform -1 0 2970 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__929_
timestamp 1701859473
transform -1 0 4250 0 1 790
box -12 -8 32 272
use FILL  FILL_2__930_
timestamp 1701859473
transform -1 0 5990 0 1 790
box -12 -8 32 272
use FILL  FILL_2__931_
timestamp 1701859473
transform 1 0 5690 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__932_
timestamp 1701859473
transform -1 0 5970 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__933_
timestamp 1701859473
transform -1 0 5990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__934_
timestamp 1701859473
transform 1 0 5330 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__935_
timestamp 1701859473
transform -1 0 6010 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__936_
timestamp 1701859473
transform 1 0 5090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__937_
timestamp 1701859473
transform 1 0 5350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__938_
timestamp 1701859473
transform 1 0 5210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__939_
timestamp 1701859473
transform -1 0 5090 0 1 790
box -12 -8 32 272
use FILL  FILL_2__940_
timestamp 1701859473
transform 1 0 5050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__941_
timestamp 1701859473
transform 1 0 5890 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__942_
timestamp 1701859473
transform -1 0 5970 0 1 270
box -12 -8 32 272
use FILL  FILL_2__943_
timestamp 1701859473
transform -1 0 6110 0 1 270
box -12 -8 32 272
use FILL  FILL_2__944_
timestamp 1701859473
transform -1 0 5190 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__945_
timestamp 1701859473
transform -1 0 5850 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__946_
timestamp 1701859473
transform 1 0 1750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__947_
timestamp 1701859473
transform 1 0 2010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__948_
timestamp 1701859473
transform -1 0 1870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__949_
timestamp 1701859473
transform -1 0 2310 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__950_
timestamp 1701859473
transform 1 0 2290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__951_
timestamp 1701859473
transform 1 0 2150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__952_
timestamp 1701859473
transform 1 0 4410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__953_
timestamp 1701859473
transform 1 0 3270 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__954_
timestamp 1701859473
transform 1 0 3410 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__955_
timestamp 1701859473
transform 1 0 3590 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__956_
timestamp 1701859473
transform 1 0 3550 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__957_
timestamp 1701859473
transform 1 0 3670 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__958_
timestamp 1701859473
transform 1 0 1750 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__959_
timestamp 1701859473
transform -1 0 1910 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__960_
timestamp 1701859473
transform 1 0 2370 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__961_
timestamp 1701859473
transform 1 0 2230 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__962_
timestamp 1701859473
transform 1 0 2850 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__963_
timestamp 1701859473
transform -1 0 3010 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__964_
timestamp 1701859473
transform 1 0 2950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__965_
timestamp 1701859473
transform -1 0 3110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__966_
timestamp 1701859473
transform -1 0 4470 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__967_
timestamp 1701859473
transform 1 0 3930 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__968_
timestamp 1701859473
transform -1 0 4330 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__969_
timestamp 1701859473
transform -1 0 5070 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__970_
timestamp 1701859473
transform -1 0 4410 0 1 790
box -12 -8 32 272
use FILL  FILL_2__971_
timestamp 1701859473
transform -1 0 4570 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__972_
timestamp 1701859473
transform 1 0 4930 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__973_
timestamp 1701859473
transform -1 0 4510 0 1 270
box -12 -8 32 272
use FILL  FILL_2__974_
timestamp 1701859473
transform -1 0 4630 0 1 270
box -12 -8 32 272
use FILL  FILL_2__975_
timestamp 1701859473
transform -1 0 5190 0 1 270
box -12 -8 32 272
use FILL  FILL_2__976_
timestamp 1701859473
transform -1 0 5070 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__977_
timestamp 1701859473
transform -1 0 5030 0 1 270
box -12 -8 32 272
use FILL  FILL_2__978_
timestamp 1701859473
transform 1 0 3770 0 1 270
box -12 -8 32 272
use FILL  FILL_2__979_
timestamp 1701859473
transform -1 0 3410 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__980_
timestamp 1701859473
transform -1 0 3550 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__981_
timestamp 1701859473
transform -1 0 5330 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__982_
timestamp 1701859473
transform -1 0 4390 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__983_
timestamp 1701859473
transform -1 0 5190 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__984_
timestamp 1701859473
transform -1 0 5370 0 1 790
box -12 -8 32 272
use FILL  FILL_2__985_
timestamp 1701859473
transform -1 0 3250 0 1 790
box -12 -8 32 272
use FILL  FILL_2__986_
timestamp 1701859473
transform 1 0 5230 0 1 790
box -12 -8 32 272
use FILL  FILL_2__987_
timestamp 1701859473
transform 1 0 4530 0 1 790
box -12 -8 32 272
use FILL  FILL_2__988_
timestamp 1701859473
transform -1 0 3670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__989_
timestamp 1701859473
transform -1 0 3810 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__990_
timestamp 1701859473
transform 1 0 3710 0 1 790
box -12 -8 32 272
use FILL  FILL_2__991_
timestamp 1701859473
transform -1 0 4710 0 1 790
box -12 -8 32 272
use FILL  FILL_2__992_
timestamp 1701859473
transform -1 0 5550 0 1 790
box -12 -8 32 272
use FILL  FILL_2__993_
timestamp 1701859473
transform -1 0 5790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__994_
timestamp 1701859473
transform -1 0 5810 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__995_
timestamp 1701859473
transform -1 0 5190 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__996_
timestamp 1701859473
transform -1 0 5210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__997_
timestamp 1701859473
transform 1 0 5670 0 1 270
box -12 -8 32 272
use FILL  FILL_2__998_
timestamp 1701859473
transform -1 0 5830 0 1 270
box -12 -8 32 272
use FILL  FILL_2__999_
timestamp 1701859473
transform 1 0 6330 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1000_
timestamp 1701859473
transform -1 0 6150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1001_
timestamp 1701859473
transform -1 0 6290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1002_
timestamp 1701859473
transform 1 0 6310 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1003_
timestamp 1701859473
transform 1 0 6130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1004_
timestamp 1701859473
transform -1 0 6270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1005_
timestamp 1701859473
transform 1 0 5190 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1006_
timestamp 1701859473
transform -1 0 5510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1007_
timestamp 1701859473
transform 1 0 5290 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1008_
timestamp 1701859473
transform 1 0 5970 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1009_
timestamp 1701859473
transform 1 0 6230 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1010_
timestamp 1701859473
transform -1 0 6270 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1011_
timestamp 1701859473
transform 1 0 3330 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1012_
timestamp 1701859473
transform -1 0 2690 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1013_
timestamp 1701859473
transform 1 0 1750 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1014_
timestamp 1701859473
transform 1 0 3490 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1015_
timestamp 1701859473
transform 1 0 2730 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1016_
timestamp 1701859473
transform -1 0 3410 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1017_
timestamp 1701859473
transform -1 0 3290 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1018_
timestamp 1701859473
transform -1 0 3430 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1019_
timestamp 1701859473
transform 1 0 3170 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1020_
timestamp 1701859473
transform -1 0 3050 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1021_
timestamp 1701859473
transform -1 0 2990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1022_
timestamp 1701859473
transform 1 0 2670 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1023_
timestamp 1701859473
transform 1 0 3090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1024_
timestamp 1701859473
transform 1 0 3230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1025_
timestamp 1701859473
transform 1 0 3350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1026_
timestamp 1701859473
transform 1 0 3450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1027_
timestamp 1701859473
transform 1 0 3610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1028_
timestamp 1701859473
transform -1 0 3550 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1029_
timestamp 1701859473
transform -1 0 3690 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1030_
timestamp 1701859473
transform -1 0 3830 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1031_
timestamp 1701859473
transform 1 0 4390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1032_
timestamp 1701859473
transform 1 0 3990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1033_
timestamp 1701859473
transform 1 0 3410 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1034_
timestamp 1701859473
transform -1 0 2830 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1035_
timestamp 1701859473
transform 1 0 970 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1036_
timestamp 1701859473
transform 1 0 2810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1037_
timestamp 1701859473
transform -1 0 3070 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1038_
timestamp 1701859473
transform 1 0 2550 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1039_
timestamp 1701859473
transform 1 0 3150 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1040_
timestamp 1701859473
transform 1 0 2370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1041_
timestamp 1701859473
transform 1 0 2210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1042_
timestamp 1701859473
transform 1 0 2170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1043_
timestamp 1701859473
transform -1 0 2330 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1044_
timestamp 1701859473
transform -1 0 2750 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1045_
timestamp 1701859473
transform -1 0 2110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1046_
timestamp 1701859473
transform 1 0 2190 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1047_
timestamp 1701859473
transform 1 0 2450 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1048_
timestamp 1701859473
transform -1 0 2910 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1049_
timestamp 1701859473
transform -1 0 2610 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1050_
timestamp 1701859473
transform -1 0 2290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1051_
timestamp 1701859473
transform -1 0 2430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1052_
timestamp 1701859473
transform 1 0 2830 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1053_
timestamp 1701859473
transform 1 0 2510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1054_
timestamp 1701859473
transform 1 0 2070 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1055_
timestamp 1701859473
transform 1 0 2730 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1056_
timestamp 1701859473
transform 1 0 2830 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1057_
timestamp 1701859473
transform 1 0 2670 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1058_
timestamp 1701859473
transform 1 0 2510 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1059_
timestamp 1701859473
transform -1 0 3010 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1060_
timestamp 1701859473
transform 1 0 3130 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1061_
timestamp 1701859473
transform 1 0 4910 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1062_
timestamp 1701859473
transform -1 0 2590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1063_
timestamp 1701859473
transform 1 0 2570 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1064_
timestamp 1701859473
transform -1 0 1510 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1065_
timestamp 1701859473
transform -1 0 2270 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1066_
timestamp 1701859473
transform -1 0 1930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1067_
timestamp 1701859473
transform 1 0 2130 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1068_
timestamp 1701859473
transform -1 0 2030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1069_
timestamp 1701859473
transform -1 0 1490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1070_
timestamp 1701859473
transform 1 0 1910 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1071_
timestamp 1701859473
transform 1 0 2070 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1072_
timestamp 1701859473
transform -1 0 1790 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1073_
timestamp 1701859473
transform -1 0 1870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1074_
timestamp 1701859473
transform -1 0 1770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1075_
timestamp 1701859473
transform -1 0 1650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1076_
timestamp 1701859473
transform 1 0 1510 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1077_
timestamp 1701859473
transform -1 0 2010 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1078_
timestamp 1701859473
transform -1 0 1590 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1079_
timestamp 1701859473
transform -1 0 1870 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1080_
timestamp 1701859473
transform 1 0 1690 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1081_
timestamp 1701859473
transform -1 0 1770 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1082_
timestamp 1701859473
transform 1 0 1970 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1083_
timestamp 1701859473
transform 1 0 1670 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1084_
timestamp 1701859473
transform 1 0 1750 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1085_
timestamp 1701859473
transform -1 0 1770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1086_
timestamp 1701859473
transform -1 0 2590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1087_
timestamp 1701859473
transform 1 0 1610 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1088_
timestamp 1701859473
transform -1 0 1610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1089_
timestamp 1701859473
transform 1 0 1830 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1090_
timestamp 1701859473
transform 1 0 1870 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1091_
timestamp 1701859473
transform -1 0 2310 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1092_
timestamp 1701859473
transform -1 0 2450 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1093_
timestamp 1701859473
transform -1 0 2410 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1094_
timestamp 1701859473
transform 1 0 2790 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1095_
timestamp 1701859473
transform -1 0 2570 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1096_
timestamp 1701859473
transform 1 0 2930 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1097_
timestamp 1701859473
transform -1 0 3050 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1098_
timestamp 1701859473
transform 1 0 4510 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1099_
timestamp 1701859473
transform 1 0 3270 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1100_
timestamp 1701859473
transform -1 0 630 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1101_
timestamp 1701859473
transform -1 0 1630 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1102_
timestamp 1701859473
transform 1 0 1470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1103_
timestamp 1701859473
transform -1 0 810 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1104_
timestamp 1701859473
transform -1 0 1650 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1105_
timestamp 1701859473
transform 1 0 1230 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1106_
timestamp 1701859473
transform -1 0 1510 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1107_
timestamp 1701859473
transform 1 0 1350 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1108_
timestamp 1701859473
transform -1 0 1330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1109_
timestamp 1701859473
transform -1 0 810 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1110_
timestamp 1701859473
transform 1 0 1030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1111_
timestamp 1701859473
transform -1 0 670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1112_
timestamp 1701859473
transform -1 0 510 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1113_
timestamp 1701859473
transform -1 0 1170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1114_
timestamp 1701859473
transform 1 0 890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1115_
timestamp 1701859473
transform -1 0 930 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1116_
timestamp 1701859473
transform -1 0 1990 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1117_
timestamp 1701859473
transform 1 0 1570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1118_
timestamp 1701859473
transform -1 0 2410 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1119_
timestamp 1701859473
transform -1 0 2010 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1120_
timestamp 1701859473
transform -1 0 1870 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1121_
timestamp 1701859473
transform -1 0 2910 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1122_
timestamp 1701859473
transform -1 0 2150 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1123_
timestamp 1701859473
transform -1 0 1630 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1124_
timestamp 1701859473
transform -1 0 1710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1125_
timestamp 1701859473
transform -1 0 3750 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1126_
timestamp 1701859473
transform -1 0 1870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1127_
timestamp 1701859473
transform -1 0 1430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1128_
timestamp 1701859473
transform -1 0 1250 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1129_
timestamp 1701859473
transform 1 0 650 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1130_
timestamp 1701859473
transform 1 0 1070 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1131_
timestamp 1701859473
transform 1 0 650 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1132_
timestamp 1701859473
transform -1 0 1390 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1133_
timestamp 1701859473
transform -1 0 990 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1134_
timestamp 1701859473
transform -1 0 830 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1135_
timestamp 1701859473
transform -1 0 1310 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1136_
timestamp 1701859473
transform -1 0 1290 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1137_
timestamp 1701859473
transform 1 0 1110 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1138_
timestamp 1701859473
transform -1 0 1150 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1139_
timestamp 1701859473
transform -1 0 750 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1140_
timestamp 1701859473
transform -1 0 1470 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1141_
timestamp 1701859473
transform -1 0 1010 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1142_
timestamp 1701859473
transform -1 0 850 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1143_
timestamp 1701859473
transform 1 0 890 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1144_
timestamp 1701859473
transform 1 0 1290 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1145_
timestamp 1701859473
transform -1 0 2190 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1146_
timestamp 1701859473
transform -1 0 1190 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1147_
timestamp 1701859473
transform -1 0 2050 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1148_
timestamp 1701859473
transform 1 0 2410 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1149_
timestamp 1701859473
transform -1 0 2270 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1150_
timestamp 1701859473
transform -1 0 2770 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1151_
timestamp 1701859473
transform 1 0 2890 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1152_
timestamp 1701859473
transform 1 0 4090 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1153_
timestamp 1701859473
transform -1 0 1790 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1154_
timestamp 1701859473
transform -1 0 470 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1155_
timestamp 1701859473
transform 1 0 2910 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1156_
timestamp 1701859473
transform -1 0 2330 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1157_
timestamp 1701859473
transform 1 0 890 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1158_
timestamp 1701859473
transform -1 0 1530 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1159_
timestamp 1701859473
transform -1 0 1370 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1160_
timestamp 1701859473
transform -1 0 1030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1161_
timestamp 1701859473
transform -1 0 350 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1162_
timestamp 1701859473
transform -1 0 1710 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1163_
timestamp 1701859473
transform 1 0 1830 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1164_
timestamp 1701859473
transform 1 0 1230 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1165_
timestamp 1701859473
transform 1 0 1470 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1166_
timestamp 1701859473
transform -1 0 1550 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1167_
timestamp 1701859473
transform -1 0 1090 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1168_
timestamp 1701859473
transform -1 0 830 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1169_
timestamp 1701859473
transform -1 0 1410 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1170_
timestamp 1701859473
transform -1 0 1150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1171_
timestamp 1701859473
transform 1 0 910 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1172_
timestamp 1701859473
transform 1 0 830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1173_
timestamp 1701859473
transform -1 0 1110 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1174_
timestamp 1701859473
transform -1 0 990 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1175_
timestamp 1701859473
transform 1 0 1370 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1176_
timestamp 1701859473
transform 1 0 1330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1177_
timestamp 1701859473
transform -1 0 1230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1178_
timestamp 1701859473
transform 1 0 1190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1179_
timestamp 1701859473
transform -1 0 1070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1180_
timestamp 1701859473
transform -1 0 970 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1181_
timestamp 1701859473
transform -1 0 950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1182_
timestamp 1701859473
transform -1 0 650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1183_
timestamp 1701859473
transform -1 0 510 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1184_
timestamp 1701859473
transform 1 0 770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1185_
timestamp 1701859473
transform -1 0 1670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1186_
timestamp 1701859473
transform -1 0 1510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1187_
timestamp 1701859473
transform -1 0 1770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1188_
timestamp 1701859473
transform -1 0 1230 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1189_
timestamp 1701859473
transform 1 0 810 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1190_
timestamp 1701859473
transform -1 0 370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1191_
timestamp 1701859473
transform -1 0 690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1192_
timestamp 1701859473
transform -1 0 370 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1193_
timestamp 1701859473
transform -1 0 670 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1194_
timestamp 1701859473
transform -1 0 70 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1195_
timestamp 1701859473
transform 1 0 190 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1196_
timestamp 1701859473
transform 1 0 1410 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1197_
timestamp 1701859473
transform 1 0 210 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1198_
timestamp 1701859473
transform -1 0 510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1199_
timestamp 1701859473
transform 1 0 490 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1200_
timestamp 1701859473
transform 1 0 170 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1201_
timestamp 1701859473
transform -1 0 70 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1202_
timestamp 1701859473
transform -1 0 70 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1203_
timestamp 1701859473
transform -1 0 350 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1204_
timestamp 1701859473
transform 1 0 50 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1205_
timestamp 1701859473
transform 1 0 310 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1206_
timestamp 1701859473
transform -1 0 690 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1207_
timestamp 1701859473
transform 1 0 210 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1208_
timestamp 1701859473
transform 1 0 350 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1209_
timestamp 1701859473
transform 1 0 510 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1210_
timestamp 1701859473
transform 1 0 1630 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1211_
timestamp 1701859473
transform 1 0 1870 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1212_
timestamp 1701859473
transform 1 0 1030 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1213_
timestamp 1701859473
transform 1 0 1450 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1214_
timestamp 1701859473
transform -1 0 2010 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1215_
timestamp 1701859473
transform 1 0 2550 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1216_
timestamp 1701859473
transform 1 0 3690 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1217_
timestamp 1701859473
transform 1 0 2110 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1218_
timestamp 1701859473
transform -1 0 850 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1219_
timestamp 1701859473
transform 1 0 1230 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1220_
timestamp 1701859473
transform 1 0 50 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1221_
timestamp 1701859473
transform -1 0 190 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1222_
timestamp 1701859473
transform 1 0 2450 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1223_
timestamp 1701859473
transform 1 0 1910 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1224_
timestamp 1701859473
transform -1 0 1490 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1225_
timestamp 1701859473
transform -1 0 910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1226_
timestamp 1701859473
transform -1 0 690 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1227_
timestamp 1701859473
transform 1 0 1290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1228_
timestamp 1701859473
transform -1 0 990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1229_
timestamp 1701859473
transform -1 0 70 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1230_
timestamp 1701859473
transform -1 0 230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1231_
timestamp 1701859473
transform 1 0 50 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1232_
timestamp 1701859473
transform -1 0 1650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1233_
timestamp 1701859473
transform -1 0 1350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1234_
timestamp 1701859473
transform 1 0 1050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1235_
timestamp 1701859473
transform -1 0 1190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1236_
timestamp 1701859473
transform -1 0 910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1237_
timestamp 1701859473
transform 1 0 950 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1238_
timestamp 1701859473
transform 1 0 1590 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1239_
timestamp 1701859473
transform -1 0 1370 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1240_
timestamp 1701859473
transform -1 0 1490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1241_
timestamp 1701859473
transform -1 0 830 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1242_
timestamp 1701859473
transform 1 0 750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1243_
timestamp 1701859473
transform -1 0 1070 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1244_
timestamp 1701859473
transform 1 0 910 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1245_
timestamp 1701859473
transform -1 0 1630 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1246_
timestamp 1701859473
transform -1 0 1550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1247_
timestamp 1701859473
transform 1 0 1050 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1248_
timestamp 1701859473
transform -1 0 1690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1249_
timestamp 1701859473
transform 1 0 1170 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1250_
timestamp 1701859473
transform -1 0 1430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1251_
timestamp 1701859473
transform -1 0 1330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1252_
timestamp 1701859473
transform -1 0 1030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1253_
timestamp 1701859473
transform -1 0 910 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1254_
timestamp 1701859473
transform -1 0 1190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1255_
timestamp 1701859473
transform -1 0 2390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1256_
timestamp 1701859473
transform -1 0 2250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1257_
timestamp 1701859473
transform -1 0 2750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1258_
timestamp 1701859473
transform -1 0 2090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1259_
timestamp 1701859473
transform -1 0 630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1260_
timestamp 1701859473
transform -1 0 370 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1261_
timestamp 1701859473
transform -1 0 630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1262_
timestamp 1701859473
transform 1 0 730 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1263_
timestamp 1701859473
transform 1 0 750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1264_
timestamp 1701859473
transform -1 0 330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1265_
timestamp 1701859473
transform -1 0 70 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1266_
timestamp 1701859473
transform -1 0 510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1267_
timestamp 1701859473
transform -1 0 350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1268_
timestamp 1701859473
transform 1 0 450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1269_
timestamp 1701859473
transform -1 0 530 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1270_
timestamp 1701859473
transform -1 0 370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1271_
timestamp 1701859473
transform 1 0 210 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1272_
timestamp 1701859473
transform 1 0 230 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1273_
timestamp 1701859473
transform 1 0 210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1274_
timestamp 1701859473
transform 1 0 510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1275_
timestamp 1701859473
transform 1 0 510 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1276_
timestamp 1701859473
transform -1 0 230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1277_
timestamp 1701859473
transform 1 0 50 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1278_
timestamp 1701859473
transform -1 0 230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1279_
timestamp 1701859473
transform -1 0 370 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1280_
timestamp 1701859473
transform -1 0 70 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1281_
timestamp 1701859473
transform 1 0 50 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1282_
timestamp 1701859473
transform 1 0 190 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1283_
timestamp 1701859473
transform -1 0 810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1284_
timestamp 1701859473
transform 1 0 350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1285_
timestamp 1701859473
transform 1 0 50 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1286_
timestamp 1701859473
transform 1 0 650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1287_
timestamp 1701859473
transform -1 0 690 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1288_
timestamp 1701859473
transform 1 0 510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1289_
timestamp 1701859473
transform 1 0 350 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1290_
timestamp 1701859473
transform 1 0 510 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1291_
timestamp 1701859473
transform 1 0 2370 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1292_
timestamp 1701859473
transform 1 0 2210 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1293_
timestamp 1701859473
transform -1 0 2950 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1294_
timestamp 1701859473
transform -1 0 3070 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1295_
timestamp 1701859473
transform 1 0 2710 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1296_
timestamp 1701859473
transform -1 0 2970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1297_
timestamp 1701859473
transform -1 0 1130 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1298_
timestamp 1701859473
transform 1 0 810 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1299_
timestamp 1701859473
transform 1 0 50 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1300_
timestamp 1701859473
transform 1 0 50 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1301_
timestamp 1701859473
transform -1 0 190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1302_
timestamp 1701859473
transform 1 0 2930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1303_
timestamp 1701859473
transform -1 0 2410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1304_
timestamp 1701859473
transform -1 0 2630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1305_
timestamp 1701859473
transform 1 0 2070 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1306_
timestamp 1701859473
transform 1 0 1950 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1307_
timestamp 1701859473
transform -1 0 2250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1308_
timestamp 1701859473
transform -1 0 1950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1309_
timestamp 1701859473
transform 1 0 3150 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1310_
timestamp 1701859473
transform -1 0 2630 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1311_
timestamp 1701859473
transform -1 0 1770 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1312_
timestamp 1701859473
transform -1 0 1650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1313_
timestamp 1701859473
transform 1 0 1210 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1314_
timestamp 1701859473
transform -1 0 1490 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1315_
timestamp 1701859473
transform -1 0 1810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1316_
timestamp 1701859473
transform -1 0 2090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1317_
timestamp 1701859473
transform 1 0 1050 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1318_
timestamp 1701859473
transform -1 0 1190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1319_
timestamp 1701859473
transform -1 0 1030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1320_
timestamp 1701859473
transform -1 0 1250 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1321_
timestamp 1701859473
transform -1 0 1330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1322_
timestamp 1701859473
transform 1 0 810 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1323_
timestamp 1701859473
transform 1 0 650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1324_
timestamp 1701859473
transform -1 0 350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1325_
timestamp 1701859473
transform -1 0 210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1326_
timestamp 1701859473
transform 1 0 1510 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1327_
timestamp 1701859473
transform -1 0 1390 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1328_
timestamp 1701859473
transform 1 0 1050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1329_
timestamp 1701859473
transform 1 0 1090 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1330_
timestamp 1701859473
transform 1 0 1350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1331_
timestamp 1701859473
transform 1 0 1190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1332_
timestamp 1701859473
transform 1 0 1770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1333_
timestamp 1701859473
transform 1 0 2730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1334_
timestamp 1701859473
transform 1 0 2010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1335_
timestamp 1701859473
transform -1 0 1670 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1336_
timestamp 1701859473
transform -1 0 1730 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1337_
timestamp 1701859473
transform 1 0 1350 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1338_
timestamp 1701859473
transform 1 0 1310 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1339_
timestamp 1701859473
transform -1 0 790 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1340_
timestamp 1701859473
transform 1 0 1470 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1341_
timestamp 1701859473
transform 1 0 1590 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1342_
timestamp 1701859473
transform -1 0 1690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1343_
timestamp 1701859473
transform -1 0 1830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1344_
timestamp 1701859473
transform 1 0 1530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1345_
timestamp 1701859473
transform -1 0 1510 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1346_
timestamp 1701859473
transform 1 0 1930 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1347_
timestamp 1701859473
transform -1 0 2130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1348_
timestamp 1701859473
transform -1 0 1650 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1349_
timestamp 1701859473
transform -1 0 1690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1350_
timestamp 1701859473
transform -1 0 910 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1351_
timestamp 1701859473
transform 1 0 1770 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1352_
timestamp 1701859473
transform -1 0 1410 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1353_
timestamp 1701859473
transform -1 0 1250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1354_
timestamp 1701859473
transform -1 0 950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1355_
timestamp 1701859473
transform -1 0 1230 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1356_
timestamp 1701859473
transform -1 0 1050 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1357_
timestamp 1701859473
transform -1 0 1110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1358_
timestamp 1701859473
transform -1 0 670 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1359_
timestamp 1701859473
transform -1 0 370 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1360_
timestamp 1701859473
transform -1 0 610 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1361_
timestamp 1701859473
transform -1 0 470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1362_
timestamp 1701859473
transform -1 0 830 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1363_
timestamp 1701859473
transform -1 0 790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1364_
timestamp 1701859473
transform -1 0 530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1365_
timestamp 1701859473
transform 1 0 190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1366_
timestamp 1701859473
transform -1 0 910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1367_
timestamp 1701859473
transform -1 0 530 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1368_
timestamp 1701859473
transform -1 0 370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1369_
timestamp 1701859473
transform 1 0 210 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1370_
timestamp 1701859473
transform -1 0 210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1371_
timestamp 1701859473
transform -1 0 210 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1372_
timestamp 1701859473
transform 1 0 50 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1373_
timestamp 1701859473
transform -1 0 70 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1374_
timestamp 1701859473
transform 1 0 50 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1375_
timestamp 1701859473
transform 1 0 50 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1376_
timestamp 1701859473
transform 1 0 210 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1377_
timestamp 1701859473
transform 1 0 510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1378_
timestamp 1701859473
transform 1 0 350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1379_
timestamp 1701859473
transform 1 0 50 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1380_
timestamp 1701859473
transform 1 0 510 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1381_
timestamp 1701859473
transform 1 0 650 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1382_
timestamp 1701859473
transform 1 0 670 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1383_
timestamp 1701859473
transform 1 0 950 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1384_
timestamp 1701859473
transform -1 0 390 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1385_
timestamp 1701859473
transform 1 0 50 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1386_
timestamp 1701859473
transform -1 0 450 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1387_
timestamp 1701859473
transform 1 0 2190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1388_
timestamp 1701859473
transform 1 0 3170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1389_
timestamp 1701859473
transform -1 0 3070 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1390_
timestamp 1701859473
transform 1 0 3270 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1391_
timestamp 1701859473
transform 1 0 3330 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1392_
timestamp 1701859473
transform -1 0 3490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1393_
timestamp 1701859473
transform -1 0 4570 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1394_
timestamp 1701859473
transform -1 0 2330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1395_
timestamp 1701859473
transform 1 0 2030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1396_
timestamp 1701859473
transform 1 0 2410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1397_
timestamp 1701859473
transform 1 0 210 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1398_
timestamp 1701859473
transform 1 0 370 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1399_
timestamp 1701859473
transform -1 0 790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1400_
timestamp 1701859473
transform 1 0 50 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1401_
timestamp 1701859473
transform 1 0 50 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1402_
timestamp 1701859473
transform 1 0 150 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1403_
timestamp 1701859473
transform 1 0 1790 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1404_
timestamp 1701859473
transform 1 0 2810 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1405_
timestamp 1701859473
transform 1 0 2550 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1406_
timestamp 1701859473
transform -1 0 3030 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1407_
timestamp 1701859473
transform -1 0 3630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1408_
timestamp 1701859473
transform 1 0 3070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1409_
timestamp 1701859473
transform -1 0 3390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1410_
timestamp 1701859473
transform 1 0 3210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1411_
timestamp 1701859473
transform -1 0 2470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1412_
timestamp 1701859473
transform 1 0 2770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1413_
timestamp 1701859473
transform 1 0 2750 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1414_
timestamp 1701859473
transform -1 0 2270 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1415_
timestamp 1701859473
transform 1 0 1470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1416_
timestamp 1701859473
transform 1 0 1870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1417_
timestamp 1701859473
transform -1 0 2170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1418_
timestamp 1701859473
transform 1 0 2390 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1419_
timestamp 1701859473
transform 1 0 2590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1420_
timestamp 1701859473
transform -1 0 1650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1421_
timestamp 1701859473
transform 1 0 1870 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1422_
timestamp 1701859473
transform -1 0 2470 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1423_
timestamp 1701859473
transform 1 0 2010 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1424_
timestamp 1701859473
transform -1 0 2510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1425_
timestamp 1701859473
transform -1 0 2110 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1426_
timestamp 1701859473
transform -1 0 2330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1427_
timestamp 1701859473
transform -1 0 2310 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1428_
timestamp 1701859473
transform 1 0 2150 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1429_
timestamp 1701859473
transform -1 0 1550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1430_
timestamp 1701859473
transform -1 0 1110 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1431_
timestamp 1701859473
transform -1 0 970 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1432_
timestamp 1701859473
transform 1 0 3070 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1433_
timestamp 1701859473
transform 1 0 3330 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1434_
timestamp 1701859473
transform -1 0 3070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1435_
timestamp 1701859473
transform 1 0 3450 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1436_
timestamp 1701859473
transform -1 0 2950 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1437_
timestamp 1701859473
transform -1 0 2910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1438_
timestamp 1701859473
transform -1 0 3090 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1439_
timestamp 1701859473
transform 1 0 3770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1440_
timestamp 1701859473
transform 1 0 3510 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1441_
timestamp 1701859473
transform -1 0 3390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1442_
timestamp 1701859473
transform -1 0 2930 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1443_
timestamp 1701859473
transform 1 0 2690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1444_
timestamp 1701859473
transform 1 0 2530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1445_
timestamp 1701859473
transform 1 0 2370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1446_
timestamp 1701859473
transform -1 0 4290 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1447_
timestamp 1701859473
transform 1 0 2590 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1448_
timestamp 1701859473
transform 1 0 1970 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1449_
timestamp 1701859473
transform 1 0 1950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1450_
timestamp 1701859473
transform 1 0 2050 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1451_
timestamp 1701859473
transform -1 0 2450 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1452_
timestamp 1701859473
transform -1 0 2130 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1453_
timestamp 1701859473
transform -1 0 2750 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1454_
timestamp 1701859473
transform -1 0 2330 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1455_
timestamp 1701859473
transform 1 0 2190 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1456_
timestamp 1701859473
transform 1 0 1670 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1457_
timestamp 1701859473
transform -1 0 1410 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1458_
timestamp 1701859473
transform -1 0 1270 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1459_
timestamp 1701859473
transform -1 0 790 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1460_
timestamp 1701859473
transform -1 0 1370 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1461_
timestamp 1701859473
transform -1 0 1210 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1462_
timestamp 1701859473
transform -1 0 2430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1463_
timestamp 1701859473
transform 1 0 1810 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1464_
timestamp 1701859473
transform -1 0 1530 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1465_
timestamp 1701859473
transform 1 0 2270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1466_
timestamp 1701859473
transform -1 0 710 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1467_
timestamp 1701859473
transform -1 0 390 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1468_
timestamp 1701859473
transform -1 0 1410 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1469_
timestamp 1701859473
transform 1 0 930 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1470_
timestamp 1701859473
transform -1 0 870 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1471_
timestamp 1701859473
transform -1 0 550 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1472_
timestamp 1701859473
transform 1 0 210 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1473_
timestamp 1701859473
transform -1 0 490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1474_
timestamp 1701859473
transform -1 0 330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1475_
timestamp 1701859473
transform -1 0 530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1476_
timestamp 1701859473
transform -1 0 370 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1477_
timestamp 1701859473
transform -1 0 70 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1478_
timestamp 1701859473
transform 1 0 170 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1479_
timestamp 1701859473
transform -1 0 70 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1480_
timestamp 1701859473
transform 1 0 210 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1481_
timestamp 1701859473
transform -1 0 630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1482_
timestamp 1701859473
transform 1 0 530 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1483_
timestamp 1701859473
transform -1 0 790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1484_
timestamp 1701859473
transform 1 0 610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1485_
timestamp 1701859473
transform -1 0 490 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1486_
timestamp 1701859473
transform 1 0 310 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1487_
timestamp 1701859473
transform 1 0 670 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1488_
timestamp 1701859473
transform -1 0 3150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1489_
timestamp 1701859473
transform -1 0 3870 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1490_
timestamp 1701859473
transform 1 0 4410 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1491_
timestamp 1701859473
transform 1 0 3270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1492_
timestamp 1701859473
transform 1 0 3390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1493_
timestamp 1701859473
transform -1 0 670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1494_
timestamp 1701859473
transform 1 0 610 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1495_
timestamp 1701859473
transform -1 0 2270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1496_
timestamp 1701859473
transform 1 0 2850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1497_
timestamp 1701859473
transform -1 0 1170 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1498_
timestamp 1701859473
transform 1 0 990 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1499_
timestamp 1701859473
transform 1 0 2750 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1500_
timestamp 1701859473
transform -1 0 3510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1501_
timestamp 1701859473
transform -1 0 3850 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1502_
timestamp 1701859473
transform 1 0 3710 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1503_
timestamp 1701859473
transform -1 0 3990 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1504_
timestamp 1701859473
transform -1 0 3670 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1505_
timestamp 1701859473
transform -1 0 3530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1506_
timestamp 1701859473
transform -1 0 4910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1507_
timestamp 1701859473
transform 1 0 3930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1508_
timestamp 1701859473
transform -1 0 3910 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1509_
timestamp 1701859473
transform -1 0 3590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1510_
timestamp 1701859473
transform -1 0 3230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1511_
timestamp 1701859473
transform 1 0 3170 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1512_
timestamp 1701859473
transform -1 0 3290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1513_
timestamp 1701859473
transform 1 0 3710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1514_
timestamp 1701859473
transform -1 0 3630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1515_
timestamp 1701859473
transform -1 0 3350 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1516_
timestamp 1701859473
transform -1 0 2970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1517_
timestamp 1701859473
transform 1 0 2810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1518_
timestamp 1701859473
transform -1 0 2690 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1519_
timestamp 1701859473
transform 1 0 2610 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1520_
timestamp 1701859473
transform 1 0 3110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1521_
timestamp 1701859473
transform -1 0 3430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1522_
timestamp 1701859473
transform 1 0 3510 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1523_
timestamp 1701859473
transform 1 0 3250 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1524_
timestamp 1701859473
transform 1 0 1830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1525_
timestamp 1701859473
transform 1 0 1950 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1526_
timestamp 1701859473
transform 1 0 4150 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1527_
timestamp 1701859473
transform -1 0 4410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1528_
timestamp 1701859473
transform 1 0 4230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1529_
timestamp 1701859473
transform 1 0 3930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1530_
timestamp 1701859473
transform -1 0 4090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1531_
timestamp 1701859473
transform 1 0 4310 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1532_
timestamp 1701859473
transform -1 0 4750 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1533_
timestamp 1701859473
transform 1 0 3750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1534_
timestamp 1701859473
transform -1 0 4190 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1535_
timestamp 1701859473
transform -1 0 4030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1536_
timestamp 1701859473
transform -1 0 4170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1537_
timestamp 1701859473
transform -1 0 4190 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1538_
timestamp 1701859473
transform -1 0 4050 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1539_
timestamp 1701859473
transform -1 0 3890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1540_
timestamp 1701859473
transform -1 0 3810 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1541_
timestamp 1701859473
transform 1 0 3670 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1542_
timestamp 1701859473
transform 1 0 2550 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1543_
timestamp 1701859473
transform 1 0 2690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1544_
timestamp 1701859473
transform 1 0 4370 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1545_
timestamp 1701859473
transform -1 0 4230 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1546_
timestamp 1701859473
transform 1 0 3930 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1547_
timestamp 1701859473
transform 1 0 4510 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1548_
timestamp 1701859473
transform -1 0 3410 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1549_
timestamp 1701859473
transform -1 0 4090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1550_
timestamp 1701859473
transform -1 0 3290 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1551_
timestamp 1701859473
transform 1 0 1090 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1552_
timestamp 1701859473
transform -1 0 1250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1553_
timestamp 1701859473
transform 1 0 3890 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1554_
timestamp 1701859473
transform -1 0 3550 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1555_
timestamp 1701859473
transform 1 0 2250 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1556_
timestamp 1701859473
transform -1 0 3130 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1557_
timestamp 1701859473
transform 1 0 2950 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1558_
timestamp 1701859473
transform 1 0 3110 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1559_
timestamp 1701859473
transform 1 0 3430 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1560_
timestamp 1701859473
transform 1 0 2650 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1561_
timestamp 1701859473
transform -1 0 3390 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1562_
timestamp 1701859473
transform -1 0 3230 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1563_
timestamp 1701859473
transform -1 0 3070 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1564_
timestamp 1701859473
transform -1 0 2990 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1565_
timestamp 1701859473
transform -1 0 2890 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1566_
timestamp 1701859473
transform -1 0 3230 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1567_
timestamp 1701859473
transform 1 0 3530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1568_
timestamp 1701859473
transform 1 0 4130 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1569_
timestamp 1701859473
transform -1 0 3950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1570_
timestamp 1701859473
transform -1 0 4610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1571_
timestamp 1701859473
transform -1 0 3270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1572_
timestamp 1701859473
transform 1 0 3730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1573_
timestamp 1701859473
transform 1 0 4730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1574_
timestamp 1701859473
transform -1 0 3750 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1575_
timestamp 1701859473
transform -1 0 3590 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1576_
timestamp 1701859473
transform 1 0 3910 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1577_
timestamp 1701859473
transform 1 0 4210 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1578_
timestamp 1701859473
transform 1 0 4070 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1579_
timestamp 1701859473
transform 1 0 4010 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1580_
timestamp 1701859473
transform 1 0 4930 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1581_
timestamp 1701859473
transform -1 0 4310 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1582_
timestamp 1701859473
transform -1 0 4850 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1583_
timestamp 1701859473
transform 1 0 5010 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1584_
timestamp 1701859473
transform 1 0 4690 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1585_
timestamp 1701859473
transform 1 0 4970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1586_
timestamp 1701859473
transform 1 0 5750 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1587_
timestamp 1701859473
transform 1 0 5350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1588_
timestamp 1701859473
transform -1 0 5350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1589_
timestamp 1701859473
transform 1 0 5050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1590_
timestamp 1701859473
transform 1 0 5590 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1591_
timestamp 1701859473
transform -1 0 4870 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1592_
timestamp 1701859473
transform 1 0 4970 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1593_
timestamp 1701859473
transform -1 0 5150 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1594_
timestamp 1701859473
transform -1 0 5450 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1595_
timestamp 1701859473
transform -1 0 4830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1596_
timestamp 1701859473
transform -1 0 4610 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1597_
timestamp 1701859473
transform 1 0 4430 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1598_
timestamp 1701859473
transform -1 0 5090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1599_
timestamp 1701859473
transform 1 0 5050 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1600_
timestamp 1701859473
transform -1 0 4950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1601_
timestamp 1701859473
transform -1 0 5290 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1602_
timestamp 1701859473
transform 1 0 4770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1603_
timestamp 1701859473
transform 1 0 5690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1604_
timestamp 1701859473
transform 1 0 4210 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1605_
timestamp 1701859473
transform 1 0 4350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1606_
timestamp 1701859473
transform 1 0 4290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1607_
timestamp 1701859473
transform 1 0 4330 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1608_
timestamp 1701859473
transform 1 0 4410 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1609_
timestamp 1701859473
transform -1 0 4730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1610_
timestamp 1701859473
transform -1 0 4570 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1611_
timestamp 1701859473
transform -1 0 4570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1612_
timestamp 1701859473
transform 1 0 4410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1613_
timestamp 1701859473
transform 1 0 4670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1614_
timestamp 1701859473
transform -1 0 4650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1615_
timestamp 1701859473
transform 1 0 4370 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1616_
timestamp 1701859473
transform 1 0 4530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1617_
timestamp 1701859473
transform 1 0 4490 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1618_
timestamp 1701859473
transform 1 0 5910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1619_
timestamp 1701859473
transform 1 0 6130 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1620_
timestamp 1701859473
transform 1 0 4650 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1621_
timestamp 1701859473
transform -1 0 4510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1622_
timestamp 1701859473
transform 1 0 4790 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1623_
timestamp 1701859473
transform -1 0 5570 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1624_
timestamp 1701859473
transform -1 0 5430 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1625_
timestamp 1701859473
transform 1 0 4670 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1626_
timestamp 1701859473
transform -1 0 5130 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1627_
timestamp 1701859473
transform 1 0 5990 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1628_
timestamp 1701859473
transform -1 0 4970 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1629_
timestamp 1701859473
transform 1 0 4790 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1630_
timestamp 1701859473
transform -1 0 5590 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1631_
timestamp 1701859473
transform 1 0 5090 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1632_
timestamp 1701859473
transform -1 0 4990 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1633_
timestamp 1701859473
transform -1 0 4830 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1634_
timestamp 1701859473
transform -1 0 2430 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1635_
timestamp 1701859473
transform 1 0 2810 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1636_
timestamp 1701859473
transform -1 0 4510 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1637_
timestamp 1701859473
transform -1 0 4670 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1638_
timestamp 1701859473
transform -1 0 4350 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1639_
timestamp 1701859473
transform -1 0 4930 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1640_
timestamp 1701859473
transform -1 0 4830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1641_
timestamp 1701859473
transform -1 0 4890 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1642_
timestamp 1701859473
transform -1 0 4750 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1643_
timestamp 1701859473
transform 1 0 5430 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1644_
timestamp 1701859473
transform 1 0 5010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1645_
timestamp 1701859473
transform -1 0 5730 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1646_
timestamp 1701859473
transform 1 0 5250 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1647_
timestamp 1701859473
transform 1 0 5210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1648_
timestamp 1701859473
transform 1 0 5630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1649_
timestamp 1701859473
transform 1 0 5210 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1650_
timestamp 1701859473
transform 1 0 5810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1651_
timestamp 1701859473
transform 1 0 5670 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1652_
timestamp 1701859473
transform 1 0 5210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1653_
timestamp 1701859473
transform 1 0 5290 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1654_
timestamp 1701859473
transform -1 0 5870 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1655_
timestamp 1701859473
transform 1 0 5130 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1656_
timestamp 1701859473
transform 1 0 5430 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1657_
timestamp 1701859473
transform 1 0 4490 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1658_
timestamp 1701859473
transform 1 0 5190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1659_
timestamp 1701859473
transform 1 0 5710 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1660_
timestamp 1701859473
transform -1 0 5210 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1661_
timestamp 1701859473
transform -1 0 5350 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1662_
timestamp 1701859473
transform 1 0 5810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1663_
timestamp 1701859473
transform 1 0 6130 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1664_
timestamp 1701859473
transform -1 0 5790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1665_
timestamp 1701859473
transform -1 0 5590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1666_
timestamp 1701859473
transform 1 0 5550 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1667_
timestamp 1701859473
transform 1 0 5630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1668_
timestamp 1701859473
transform -1 0 6270 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1669_
timestamp 1701859473
transform 1 0 5850 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1670_
timestamp 1701859473
transform -1 0 5490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1671_
timestamp 1701859473
transform -1 0 5990 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1672_
timestamp 1701859473
transform 1 0 5950 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1673_
timestamp 1701859473
transform 1 0 4010 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1674_
timestamp 1701859473
transform -1 0 4190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1675_
timestamp 1701859473
transform 1 0 5950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1676_
timestamp 1701859473
transform 1 0 6230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1677_
timestamp 1701859473
transform -1 0 6130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1678_
timestamp 1701859473
transform -1 0 6110 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1679_
timestamp 1701859473
transform 1 0 5870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1680_
timestamp 1701859473
transform 1 0 6270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1681_
timestamp 1701859473
transform 1 0 6150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1682_
timestamp 1701859473
transform 1 0 6010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1683_
timestamp 1701859473
transform -1 0 5770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1684_
timestamp 1701859473
transform 1 0 5910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1685_
timestamp 1701859473
transform 1 0 5830 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1686_
timestamp 1701859473
transform -1 0 5490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1687_
timestamp 1701859473
transform -1 0 6050 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1688_
timestamp 1701859473
transform 1 0 6030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1689_
timestamp 1701859473
transform -1 0 6310 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1690_
timestamp 1701859473
transform 1 0 6130 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1691_
timestamp 1701859473
transform -1 0 5350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1692_
timestamp 1701859473
transform -1 0 5450 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1693_
timestamp 1701859473
transform 1 0 5270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1694_
timestamp 1701859473
transform -1 0 6010 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1695_
timestamp 1701859473
transform -1 0 5530 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1696_
timestamp 1701859473
transform -1 0 5390 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1697_
timestamp 1701859473
transform 1 0 5350 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1698_
timestamp 1701859473
transform 1 0 5730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1699_
timestamp 1701859473
transform 1 0 5610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1700_
timestamp 1701859473
transform -1 0 5310 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1701_
timestamp 1701859473
transform 1 0 5290 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1702_
timestamp 1701859473
transform 1 0 6010 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1703_
timestamp 1701859473
transform -1 0 5190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1704_
timestamp 1701859473
transform 1 0 4870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1705_
timestamp 1701859473
transform -1 0 5330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1706_
timestamp 1701859473
transform -1 0 5470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1707_
timestamp 1701859473
transform 1 0 5450 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1708_
timestamp 1701859473
transform 1 0 6190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1709_
timestamp 1701859473
transform 1 0 6290 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1710_
timestamp 1701859473
transform 1 0 5630 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1711_
timestamp 1701859473
transform 1 0 5430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1712_
timestamp 1701859473
transform -1 0 5070 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1713_
timestamp 1701859473
transform 1 0 4750 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1714_
timestamp 1701859473
transform 1 0 4630 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1715_
timestamp 1701859473
transform -1 0 4530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1716_
timestamp 1701859473
transform 1 0 4650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1717_
timestamp 1701859473
transform -1 0 4970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1718_
timestamp 1701859473
transform 1 0 5090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1719_
timestamp 1701859473
transform 1 0 5270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1720_
timestamp 1701859473
transform -1 0 5490 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1721_
timestamp 1701859473
transform 1 0 5810 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1722_
timestamp 1701859473
transform 1 0 4690 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1723_
timestamp 1701859473
transform 1 0 4130 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1724_
timestamp 1701859473
transform 1 0 4810 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1725_
timestamp 1701859473
transform 1 0 4950 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1726_
timestamp 1701859473
transform 1 0 5110 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1727_
timestamp 1701859473
transform -1 0 5730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1728_
timestamp 1701859473
transform 1 0 5410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1729_
timestamp 1701859473
transform 1 0 5230 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1730_
timestamp 1701859473
transform 1 0 5550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1731_
timestamp 1701859473
transform 1 0 6010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1732_
timestamp 1701859473
transform 1 0 5870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1733_
timestamp 1701859473
transform 1 0 5790 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1734_
timestamp 1701859473
transform -1 0 6310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1735_
timestamp 1701859473
transform -1 0 6310 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1736_
timestamp 1701859473
transform -1 0 6070 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1737_
timestamp 1701859473
transform 1 0 5930 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1738_
timestamp 1701859473
transform 1 0 6150 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1739_
timestamp 1701859473
transform -1 0 6170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1740_
timestamp 1701859473
transform 1 0 6190 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1741_
timestamp 1701859473
transform 1 0 6310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1742_
timestamp 1701859473
transform 1 0 6310 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1743_
timestamp 1701859473
transform 1 0 5910 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1744_
timestamp 1701859473
transform 1 0 5630 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1745_
timestamp 1701859473
transform 1 0 5610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1746_
timestamp 1701859473
transform 1 0 6270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1747_
timestamp 1701859473
transform 1 0 6110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1748_
timestamp 1701859473
transform -1 0 6310 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1749_
timestamp 1701859473
transform 1 0 4770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1750_
timestamp 1701859473
transform -1 0 4090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1751_
timestamp 1701859473
transform 1 0 4350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1752_
timestamp 1701859473
transform 1 0 3930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1753_
timestamp 1701859473
transform 1 0 4250 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1754_
timestamp 1701859473
transform 1 0 4370 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1755_
timestamp 1701859473
transform 1 0 4710 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1756_
timestamp 1701859473
transform -1 0 4230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1757_
timestamp 1701859473
transform 1 0 5490 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1758_
timestamp 1701859473
transform 1 0 6050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1759_
timestamp 1701859473
transform 1 0 5650 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1760_
timestamp 1701859473
transform 1 0 6150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1761_
timestamp 1701859473
transform 1 0 5910 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1762_
timestamp 1701859473
transform 1 0 6030 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1763_
timestamp 1701859473
transform 1 0 6170 0 -1 5990
box -12 -8 32 272
use FILL  FILL_2__1764_
timestamp 1701859473
transform -1 0 6230 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1765_
timestamp 1701859473
transform 1 0 6030 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1766_
timestamp 1701859473
transform -1 0 6150 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1767_
timestamp 1701859473
transform -1 0 6310 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1768_
timestamp 1701859473
transform -1 0 6350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1769_
timestamp 1701859473
transform -1 0 6170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1770_
timestamp 1701859473
transform 1 0 5350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1771_
timestamp 1701859473
transform -1 0 5770 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1772_
timestamp 1701859473
transform 1 0 5590 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1773_
timestamp 1701859473
transform -1 0 6290 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1774_
timestamp 1701859473
transform -1 0 6070 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1775_
timestamp 1701859473
transform -1 0 6010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1776_
timestamp 1701859473
transform -1 0 5910 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1777_
timestamp 1701859473
transform -1 0 4910 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1778_
timestamp 1701859473
transform 1 0 3490 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1779_
timestamp 1701859473
transform 1 0 4530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1780_
timestamp 1701859473
transform 1 0 4410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1781_
timestamp 1701859473
transform 1 0 4650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1782_
timestamp 1701859473
transform -1 0 4550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1783_
timestamp 1701859473
transform 1 0 4950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1784_
timestamp 1701859473
transform -1 0 5030 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1785_
timestamp 1701859473
transform 1 0 5150 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1786_
timestamp 1701859473
transform 1 0 5250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1787_
timestamp 1701859473
transform -1 0 5570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1788_
timestamp 1701859473
transform 1 0 5670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1789_
timestamp 1701859473
transform -1 0 5850 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1790_
timestamp 1701859473
transform -1 0 5490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1791_
timestamp 1701859473
transform -1 0 5850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1792_
timestamp 1701859473
transform 1 0 5410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1793_
timestamp 1701859473
transform -1 0 5110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1794_
timestamp 1701859473
transform -1 0 4550 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1795_
timestamp 1701859473
transform -1 0 4570 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1796_
timestamp 1701859473
transform -1 0 5050 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1797_
timestamp 1701859473
transform 1 0 5390 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1798_
timestamp 1701859473
transform -1 0 5510 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1799_
timestamp 1701859473
transform -1 0 5250 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1800_
timestamp 1701859473
transform 1 0 5210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1801_
timestamp 1701859473
transform -1 0 5570 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1802_
timestamp 1701859473
transform -1 0 3490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1803_
timestamp 1701859473
transform -1 0 4510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1804_
timestamp 1701859473
transform -1 0 4350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1805_
timestamp 1701859473
transform -1 0 4110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1806_
timestamp 1701859473
transform 1 0 3930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1807_
timestamp 1701859473
transform -1 0 3390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1808_
timestamp 1701859473
transform 1 0 4210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1809_
timestamp 1701859473
transform 1 0 4070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1810_
timestamp 1701859473
transform -1 0 3630 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1811_
timestamp 1701859473
transform -1 0 4350 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1812_
timestamp 1701859473
transform 1 0 4190 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1813_
timestamp 1701859473
transform 1 0 3910 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1814_
timestamp 1701859473
transform -1 0 4210 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1815_
timestamp 1701859473
transform 1 0 4030 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1816_
timestamp 1701859473
transform -1 0 4290 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1817_
timestamp 1701859473
transform 1 0 3890 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1818_
timestamp 1701859473
transform 1 0 3870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1819_
timestamp 1701859473
transform 1 0 3570 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1820_
timestamp 1701859473
transform -1 0 3790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1821_
timestamp 1701859473
transform 1 0 3630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1822_
timestamp 1701859473
transform -1 0 4090 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1823_
timestamp 1701859473
transform 1 0 4050 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1824_
timestamp 1701859473
transform 1 0 4030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1825_
timestamp 1701859473
transform 1 0 3150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1826_
timestamp 1701859473
transform 1 0 2870 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1827_
timestamp 1701859473
transform -1 0 2710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1828_
timestamp 1701859473
transform 1 0 2830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1829_
timestamp 1701859473
transform -1 0 3250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1830_
timestamp 1701859473
transform -1 0 2810 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1831_
timestamp 1701859473
transform -1 0 2730 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1832_
timestamp 1701859473
transform 1 0 3230 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1833_
timestamp 1701859473
transform -1 0 3290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1834_
timestamp 1701859473
transform -1 0 4030 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1835_
timestamp 1701859473
transform 1 0 3610 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1836_
timestamp 1701859473
transform -1 0 3290 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1837_
timestamp 1701859473
transform -1 0 3430 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1838_
timestamp 1701859473
transform -1 0 3030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1839_
timestamp 1701859473
transform 1 0 2870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1840_
timestamp 1701859473
transform 1 0 2350 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1841_
timestamp 1701859473
transform 1 0 2090 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1842_
timestamp 1701859473
transform -1 0 2050 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1843_
timestamp 1701859473
transform -1 0 2190 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1844_
timestamp 1701859473
transform -1 0 2530 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1845_
timestamp 1701859473
transform -1 0 2650 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1846_
timestamp 1701859473
transform -1 0 2350 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1847_
timestamp 1701859473
transform -1 0 2470 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1848_
timestamp 1701859473
transform 1 0 2810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1849_
timestamp 1701859473
transform 1 0 2670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1911_
timestamp 1701859473
transform 1 0 6270 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1912_
timestamp 1701859473
transform 1 0 2190 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1913_
timestamp 1701859473
transform 1 0 2110 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1914_
timestamp 1701859473
transform 1 0 3650 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1915_
timestamp 1701859473
transform 1 0 3790 0 1 5470
box -12 -8 32 272
use FILL  FILL_2__1916_
timestamp 1701859473
transform 1 0 6290 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1917_
timestamp 1701859473
transform 1 0 6150 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1918_
timestamp 1701859473
transform 1 0 5850 0 1 5990
box -12 -8 32 272
use FILL  FILL_2__1919_
timestamp 1701859473
transform -1 0 5710 0 1 790
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert0
timestamp 1701859473
transform 1 0 4770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert1
timestamp 1701859473
transform -1 0 4390 0 1 270
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert2
timestamp 1701859473
transform -1 0 4250 0 -1 270
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert3
timestamp 1701859473
transform 1 0 5370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert4
timestamp 1701859473
transform 1 0 5530 0 1 270
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert12
timestamp 1701859473
transform 1 0 2090 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert13
timestamp 1701859473
transform 1 0 2230 0 1 1830
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert14
timestamp 1701859473
transform 1 0 1330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert15
timestamp 1701859473
transform -1 0 1910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert16
timestamp 1701859473
transform -1 0 3570 0 1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert17
timestamp 1701859473
transform 1 0 3090 0 1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert18
timestamp 1701859473
transform -1 0 3390 0 1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert19
timestamp 1701859473
transform -1 0 3010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert20
timestamp 1701859473
transform 1 0 3930 0 1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert21
timestamp 1701859473
transform -1 0 4090 0 1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert22
timestamp 1701859473
transform -1 0 5650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert23
timestamp 1701859473
transform -1 0 3610 0 1 790
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert24
timestamp 1701859473
transform 1 0 4090 0 1 790
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert25
timestamp 1701859473
transform 1 0 4910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert5
timestamp 1701859473
transform 1 0 4930 0 1 1310
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert6
timestamp 1701859473
transform 1 0 4930 0 1 1830
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert7
timestamp 1701859473
transform -1 0 4130 0 1 270
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert8
timestamp 1701859473
transform -1 0 3690 0 1 2350
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert9
timestamp 1701859473
transform -1 0 3450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert10
timestamp 1701859473
transform 1 0 4670 0 1 1310
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert11
timestamp 1701859473
transform -1 0 4710 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__923_
timestamp 1701859473
transform 1 0 4230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__925_
timestamp 1701859473
transform -1 0 5870 0 1 790
box -12 -8 32 272
use FILL  FILL_3__926_
timestamp 1701859473
transform -1 0 6170 0 1 790
box -12 -8 32 272
use FILL  FILL_3__928_
timestamp 1701859473
transform -1 0 2990 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__930_
timestamp 1701859473
transform -1 0 6010 0 1 790
box -12 -8 32 272
use FILL  FILL_3__932_
timestamp 1701859473
transform -1 0 5990 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__933_
timestamp 1701859473
transform -1 0 6010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__935_
timestamp 1701859473
transform -1 0 6030 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__937_
timestamp 1701859473
transform 1 0 5370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__938_
timestamp 1701859473
transform 1 0 5230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__940_
timestamp 1701859473
transform 1 0 5070 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__942_
timestamp 1701859473
transform -1 0 5990 0 1 270
box -12 -8 32 272
use FILL  FILL_3__943_
timestamp 1701859473
transform -1 0 6130 0 1 270
box -12 -8 32 272
use FILL  FILL_3__945_
timestamp 1701859473
transform -1 0 5870 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__947_
timestamp 1701859473
transform 1 0 2030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__948_
timestamp 1701859473
transform -1 0 1890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__950_
timestamp 1701859473
transform 1 0 2310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__952_
timestamp 1701859473
transform 1 0 4430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__953_
timestamp 1701859473
transform 1 0 3290 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__955_
timestamp 1701859473
transform 1 0 3610 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__957_
timestamp 1701859473
transform 1 0 3690 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__958_
timestamp 1701859473
transform 1 0 1770 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__960_
timestamp 1701859473
transform 1 0 2390 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__962_
timestamp 1701859473
transform 1 0 2870 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__964_
timestamp 1701859473
transform 1 0 2970 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__965_
timestamp 1701859473
transform -1 0 3130 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__967_
timestamp 1701859473
transform 1 0 3950 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__969_
timestamp 1701859473
transform -1 0 5090 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__970_
timestamp 1701859473
transform -1 0 4430 0 1 790
box -12 -8 32 272
use FILL  FILL_3__972_
timestamp 1701859473
transform 1 0 4950 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__974_
timestamp 1701859473
transform -1 0 4650 0 1 270
box -12 -8 32 272
use FILL  FILL_3__975_
timestamp 1701859473
transform -1 0 5210 0 1 270
box -12 -8 32 272
use FILL  FILL_3__977_
timestamp 1701859473
transform -1 0 5050 0 1 270
box -12 -8 32 272
use FILL  FILL_3__979_
timestamp 1701859473
transform -1 0 3430 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__980_
timestamp 1701859473
transform -1 0 3570 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__982_
timestamp 1701859473
transform -1 0 4410 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__984_
timestamp 1701859473
transform -1 0 5390 0 1 790
box -12 -8 32 272
use FILL  FILL_3__985_
timestamp 1701859473
transform -1 0 3270 0 1 790
box -12 -8 32 272
use FILL  FILL_3__987_
timestamp 1701859473
transform 1 0 4550 0 1 790
box -12 -8 32 272
use FILL  FILL_3__989_
timestamp 1701859473
transform -1 0 3830 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__991_
timestamp 1701859473
transform -1 0 4730 0 1 790
box -12 -8 32 272
use FILL  FILL_3__992_
timestamp 1701859473
transform -1 0 5570 0 1 790
box -12 -8 32 272
use FILL  FILL_3__994_
timestamp 1701859473
transform -1 0 5830 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__996_
timestamp 1701859473
transform -1 0 5230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__997_
timestamp 1701859473
transform 1 0 5690 0 1 270
box -12 -8 32 272
use FILL  FILL_3__999_
timestamp 1701859473
transform 1 0 6350 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1000_
timestamp 1701859473
transform -1 0 6170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1002_
timestamp 1701859473
transform 1 0 6330 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1004_
timestamp 1701859473
transform -1 0 6290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1006_
timestamp 1701859473
transform -1 0 5530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1007_
timestamp 1701859473
transform 1 0 5310 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1009_
timestamp 1701859473
transform 1 0 6250 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1011_
timestamp 1701859473
transform 1 0 3350 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1012_
timestamp 1701859473
transform -1 0 2710 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1014_
timestamp 1701859473
transform 1 0 3510 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1016_
timestamp 1701859473
transform -1 0 3430 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1017_
timestamp 1701859473
transform -1 0 3310 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1019_
timestamp 1701859473
transform 1 0 3190 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1021_
timestamp 1701859473
transform -1 0 3010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1022_
timestamp 1701859473
transform 1 0 2690 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1024_
timestamp 1701859473
transform 1 0 3250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1026_
timestamp 1701859473
transform 1 0 3470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1027_
timestamp 1701859473
transform 1 0 3630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1029_
timestamp 1701859473
transform -1 0 3710 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1031_
timestamp 1701859473
transform 1 0 4410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1032_
timestamp 1701859473
transform 1 0 4010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1034_
timestamp 1701859473
transform -1 0 2850 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1036_
timestamp 1701859473
transform 1 0 2830 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1038_
timestamp 1701859473
transform 1 0 2570 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1039_
timestamp 1701859473
transform 1 0 3170 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1041_
timestamp 1701859473
transform 1 0 2230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1043_
timestamp 1701859473
transform -1 0 2350 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1044_
timestamp 1701859473
transform -1 0 2770 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1046_
timestamp 1701859473
transform 1 0 2210 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1048_
timestamp 1701859473
transform -1 0 2930 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1049_
timestamp 1701859473
transform -1 0 2630 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1051_
timestamp 1701859473
transform -1 0 2450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1053_
timestamp 1701859473
transform 1 0 2530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1054_
timestamp 1701859473
transform 1 0 2090 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1056_
timestamp 1701859473
transform 1 0 2850 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1058_
timestamp 1701859473
transform 1 0 2530 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1059_
timestamp 1701859473
transform -1 0 3030 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1061_
timestamp 1701859473
transform 1 0 4930 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1063_
timestamp 1701859473
transform 1 0 2590 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1065_
timestamp 1701859473
transform -1 0 2290 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1066_
timestamp 1701859473
transform -1 0 1950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1068_
timestamp 1701859473
transform -1 0 2050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1070_
timestamp 1701859473
transform 1 0 1930 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1071_
timestamp 1701859473
transform 1 0 2090 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1073_
timestamp 1701859473
transform -1 0 1890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1075_
timestamp 1701859473
transform -1 0 1670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1076_
timestamp 1701859473
transform 1 0 1530 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1078_
timestamp 1701859473
transform -1 0 1610 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1080_
timestamp 1701859473
transform 1 0 1710 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1081_
timestamp 1701859473
transform -1 0 1790 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1083_
timestamp 1701859473
transform 1 0 1690 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1085_
timestamp 1701859473
transform -1 0 1790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1086_
timestamp 1701859473
transform -1 0 2610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1088_
timestamp 1701859473
transform -1 0 1630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1090_
timestamp 1701859473
transform 1 0 1890 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1091_
timestamp 1701859473
transform -1 0 2330 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1093_
timestamp 1701859473
transform -1 0 2430 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1095_
timestamp 1701859473
transform -1 0 2590 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1097_
timestamp 1701859473
transform -1 0 3070 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1098_
timestamp 1701859473
transform 1 0 4530 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1100_
timestamp 1701859473
transform -1 0 650 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1102_
timestamp 1701859473
transform 1 0 1490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1103_
timestamp 1701859473
transform -1 0 830 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1105_
timestamp 1701859473
transform 1 0 1250 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1107_
timestamp 1701859473
transform 1 0 1370 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1108_
timestamp 1701859473
transform -1 0 1350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1110_
timestamp 1701859473
transform 1 0 1050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1112_
timestamp 1701859473
transform -1 0 530 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1113_
timestamp 1701859473
transform -1 0 1190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1115_
timestamp 1701859473
transform -1 0 950 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1117_
timestamp 1701859473
transform 1 0 1590 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1118_
timestamp 1701859473
transform -1 0 2430 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1120_
timestamp 1701859473
transform -1 0 1890 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1122_
timestamp 1701859473
transform -1 0 2170 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1124_
timestamp 1701859473
transform -1 0 1730 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1125_
timestamp 1701859473
transform -1 0 3770 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1127_
timestamp 1701859473
transform -1 0 1450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1129_
timestamp 1701859473
transform 1 0 670 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1130_
timestamp 1701859473
transform 1 0 1090 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1132_
timestamp 1701859473
transform -1 0 1410 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1134_
timestamp 1701859473
transform -1 0 850 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1135_
timestamp 1701859473
transform -1 0 1330 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1137_
timestamp 1701859473
transform 1 0 1130 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1139_
timestamp 1701859473
transform -1 0 770 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1140_
timestamp 1701859473
transform -1 0 1490 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1142_
timestamp 1701859473
transform -1 0 870 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1144_
timestamp 1701859473
transform 1 0 1310 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1145_
timestamp 1701859473
transform -1 0 2210 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1147_
timestamp 1701859473
transform -1 0 2070 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1149_
timestamp 1701859473
transform -1 0 2290 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1150_
timestamp 1701859473
transform -1 0 2790 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1152_
timestamp 1701859473
transform 1 0 4110 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1154_
timestamp 1701859473
transform -1 0 490 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1156_
timestamp 1701859473
transform -1 0 2350 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1157_
timestamp 1701859473
transform 1 0 910 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1159_
timestamp 1701859473
transform -1 0 1390 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1161_
timestamp 1701859473
transform -1 0 370 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1162_
timestamp 1701859473
transform -1 0 1730 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1164_
timestamp 1701859473
transform 1 0 1250 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1166_
timestamp 1701859473
transform -1 0 1570 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1167_
timestamp 1701859473
transform -1 0 1110 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1169_
timestamp 1701859473
transform -1 0 1430 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1171_
timestamp 1701859473
transform 1 0 930 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1172_
timestamp 1701859473
transform 1 0 850 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1174_
timestamp 1701859473
transform -1 0 1010 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1176_
timestamp 1701859473
transform 1 0 1350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1177_
timestamp 1701859473
transform -1 0 1250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1179_
timestamp 1701859473
transform -1 0 1090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1181_
timestamp 1701859473
transform -1 0 970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1183_
timestamp 1701859473
transform -1 0 530 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1184_
timestamp 1701859473
transform 1 0 790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1186_
timestamp 1701859473
transform -1 0 1530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1188_
timestamp 1701859473
transform -1 0 1250 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1189_
timestamp 1701859473
transform 1 0 830 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1191_
timestamp 1701859473
transform -1 0 710 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1193_
timestamp 1701859473
transform -1 0 690 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1194_
timestamp 1701859473
transform -1 0 90 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1196_
timestamp 1701859473
transform 1 0 1430 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1198_
timestamp 1701859473
transform -1 0 530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1199_
timestamp 1701859473
transform 1 0 510 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1201_
timestamp 1701859473
transform -1 0 90 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1203_
timestamp 1701859473
transform -1 0 370 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1204_
timestamp 1701859473
transform 1 0 70 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1206_
timestamp 1701859473
transform -1 0 710 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1208_
timestamp 1701859473
transform 1 0 370 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1209_
timestamp 1701859473
transform 1 0 530 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1211_
timestamp 1701859473
transform 1 0 1890 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1213_
timestamp 1701859473
transform 1 0 1470 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1215_
timestamp 1701859473
transform 1 0 2570 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1216_
timestamp 1701859473
transform 1 0 3710 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1218_
timestamp 1701859473
transform -1 0 870 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1220_
timestamp 1701859473
transform 1 0 70 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1221_
timestamp 1701859473
transform -1 0 210 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1223_
timestamp 1701859473
transform 1 0 1930 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1225_
timestamp 1701859473
transform -1 0 930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1226_
timestamp 1701859473
transform -1 0 710 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1228_
timestamp 1701859473
transform -1 0 1010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1230_
timestamp 1701859473
transform -1 0 250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1231_
timestamp 1701859473
transform 1 0 70 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1233_
timestamp 1701859473
transform -1 0 1370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1235_
timestamp 1701859473
transform -1 0 1210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1236_
timestamp 1701859473
transform -1 0 930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1238_
timestamp 1701859473
transform 1 0 1610 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1240_
timestamp 1701859473
transform -1 0 1510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1242_
timestamp 1701859473
transform 1 0 770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1243_
timestamp 1701859473
transform -1 0 1090 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1245_
timestamp 1701859473
transform -1 0 1650 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1247_
timestamp 1701859473
transform 1 0 1070 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1248_
timestamp 1701859473
transform -1 0 1710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1250_
timestamp 1701859473
transform -1 0 1450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1252_
timestamp 1701859473
transform -1 0 1050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1253_
timestamp 1701859473
transform -1 0 930 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1255_
timestamp 1701859473
transform -1 0 2410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1257_
timestamp 1701859473
transform -1 0 2770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1258_
timestamp 1701859473
transform -1 0 2110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1260_
timestamp 1701859473
transform -1 0 390 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1262_
timestamp 1701859473
transform 1 0 750 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1263_
timestamp 1701859473
transform 1 0 770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1265_
timestamp 1701859473
transform -1 0 90 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1267_
timestamp 1701859473
transform -1 0 370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1268_
timestamp 1701859473
transform 1 0 470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1270_
timestamp 1701859473
transform -1 0 390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1272_
timestamp 1701859473
transform 1 0 250 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1274_
timestamp 1701859473
transform 1 0 530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1275_
timestamp 1701859473
transform 1 0 530 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1277_
timestamp 1701859473
transform 1 0 70 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1279_
timestamp 1701859473
transform -1 0 390 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1280_
timestamp 1701859473
transform -1 0 90 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1282_
timestamp 1701859473
transform 1 0 210 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1284_
timestamp 1701859473
transform 1 0 370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1285_
timestamp 1701859473
transform 1 0 70 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1287_
timestamp 1701859473
transform -1 0 710 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1289_
timestamp 1701859473
transform 1 0 370 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1290_
timestamp 1701859473
transform 1 0 530 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1292_
timestamp 1701859473
transform 1 0 2230 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1294_
timestamp 1701859473
transform -1 0 3090 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1295_
timestamp 1701859473
transform 1 0 2730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1297_
timestamp 1701859473
transform -1 0 1150 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1299_
timestamp 1701859473
transform 1 0 70 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1300_
timestamp 1701859473
transform 1 0 70 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1302_
timestamp 1701859473
transform 1 0 2950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1304_
timestamp 1701859473
transform -1 0 2650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1306_
timestamp 1701859473
transform 1 0 1970 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1307_
timestamp 1701859473
transform -1 0 2270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1309_
timestamp 1701859473
transform 1 0 3170 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1311_
timestamp 1701859473
transform -1 0 1790 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1312_
timestamp 1701859473
transform -1 0 1670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1314_
timestamp 1701859473
transform -1 0 1510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1316_
timestamp 1701859473
transform -1 0 2110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1317_
timestamp 1701859473
transform 1 0 1070 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1319_
timestamp 1701859473
transform -1 0 1050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1321_
timestamp 1701859473
transform -1 0 1350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1322_
timestamp 1701859473
transform 1 0 830 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1324_
timestamp 1701859473
transform -1 0 370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1326_
timestamp 1701859473
transform 1 0 1530 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1327_
timestamp 1701859473
transform -1 0 1410 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1329_
timestamp 1701859473
transform 1 0 1110 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1331_
timestamp 1701859473
transform 1 0 1210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1333_
timestamp 1701859473
transform 1 0 2750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1334_
timestamp 1701859473
transform 1 0 2030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1336_
timestamp 1701859473
transform -1 0 1750 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1338_
timestamp 1701859473
transform 1 0 1330 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1339_
timestamp 1701859473
transform -1 0 810 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1341_
timestamp 1701859473
transform 1 0 1610 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1343_
timestamp 1701859473
transform -1 0 1850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1344_
timestamp 1701859473
transform 1 0 1550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1346_
timestamp 1701859473
transform 1 0 1950 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1348_
timestamp 1701859473
transform -1 0 1670 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1349_
timestamp 1701859473
transform -1 0 1710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1351_
timestamp 1701859473
transform 1 0 1790 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1353_
timestamp 1701859473
transform -1 0 1270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1354_
timestamp 1701859473
transform -1 0 970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1356_
timestamp 1701859473
transform -1 0 1070 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1358_
timestamp 1701859473
transform -1 0 690 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1359_
timestamp 1701859473
transform -1 0 390 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1361_
timestamp 1701859473
transform -1 0 490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1363_
timestamp 1701859473
transform -1 0 810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1365_
timestamp 1701859473
transform 1 0 210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1366_
timestamp 1701859473
transform -1 0 930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1368_
timestamp 1701859473
transform -1 0 390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1370_
timestamp 1701859473
transform -1 0 230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1371_
timestamp 1701859473
transform -1 0 230 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1373_
timestamp 1701859473
transform -1 0 90 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1375_
timestamp 1701859473
transform 1 0 70 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1376_
timestamp 1701859473
transform 1 0 230 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1378_
timestamp 1701859473
transform 1 0 370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1380_
timestamp 1701859473
transform 1 0 530 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1381_
timestamp 1701859473
transform 1 0 670 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1383_
timestamp 1701859473
transform 1 0 970 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1385_
timestamp 1701859473
transform 1 0 70 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1386_
timestamp 1701859473
transform -1 0 470 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1388_
timestamp 1701859473
transform 1 0 3190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1390_
timestamp 1701859473
transform 1 0 3290 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1392_
timestamp 1701859473
transform -1 0 3510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1393_
timestamp 1701859473
transform -1 0 4590 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1395_
timestamp 1701859473
transform 1 0 2050 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1397_
timestamp 1701859473
transform 1 0 230 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1398_
timestamp 1701859473
transform 1 0 390 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1400_
timestamp 1701859473
transform 1 0 70 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1402_
timestamp 1701859473
transform 1 0 170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1403_
timestamp 1701859473
transform 1 0 1810 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1405_
timestamp 1701859473
transform 1 0 2570 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1407_
timestamp 1701859473
transform -1 0 3650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1408_
timestamp 1701859473
transform 1 0 3090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1410_
timestamp 1701859473
transform 1 0 3230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1412_
timestamp 1701859473
transform 1 0 2790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1413_
timestamp 1701859473
transform 1 0 2770 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1415_
timestamp 1701859473
transform 1 0 1490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1417_
timestamp 1701859473
transform -1 0 2190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1418_
timestamp 1701859473
transform 1 0 2410 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1420_
timestamp 1701859473
transform -1 0 1670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1422_
timestamp 1701859473
transform -1 0 2490 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1424_
timestamp 1701859473
transform -1 0 2530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1425_
timestamp 1701859473
transform -1 0 2130 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1427_
timestamp 1701859473
transform -1 0 2330 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1429_
timestamp 1701859473
transform -1 0 1570 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1430_
timestamp 1701859473
transform -1 0 1130 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1432_
timestamp 1701859473
transform 1 0 3090 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1434_
timestamp 1701859473
transform -1 0 3090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1435_
timestamp 1701859473
transform 1 0 3470 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1437_
timestamp 1701859473
transform -1 0 2930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1439_
timestamp 1701859473
transform 1 0 3790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1440_
timestamp 1701859473
transform 1 0 3530 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1442_
timestamp 1701859473
transform -1 0 2950 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1444_
timestamp 1701859473
transform 1 0 2550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1445_
timestamp 1701859473
transform 1 0 2390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1447_
timestamp 1701859473
transform 1 0 2610 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1449_
timestamp 1701859473
transform 1 0 1970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1451_
timestamp 1701859473
transform -1 0 2470 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1452_
timestamp 1701859473
transform -1 0 2150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1454_
timestamp 1701859473
transform -1 0 2350 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1456_
timestamp 1701859473
transform 1 0 1690 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1457_
timestamp 1701859473
transform -1 0 1430 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1459_
timestamp 1701859473
transform -1 0 810 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1461_
timestamp 1701859473
transform -1 0 1230 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1462_
timestamp 1701859473
transform -1 0 2450 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1464_
timestamp 1701859473
transform -1 0 1550 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1466_
timestamp 1701859473
transform -1 0 730 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1467_
timestamp 1701859473
transform -1 0 410 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1469_
timestamp 1701859473
transform 1 0 950 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1471_
timestamp 1701859473
transform -1 0 570 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1472_
timestamp 1701859473
transform 1 0 230 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1474_
timestamp 1701859473
transform -1 0 350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1476_
timestamp 1701859473
transform -1 0 390 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1477_
timestamp 1701859473
transform -1 0 90 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1479_
timestamp 1701859473
transform -1 0 90 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1481_
timestamp 1701859473
transform -1 0 650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1483_
timestamp 1701859473
transform -1 0 810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1484_
timestamp 1701859473
transform 1 0 630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1486_
timestamp 1701859473
transform 1 0 330 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1488_
timestamp 1701859473
transform -1 0 3170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1489_
timestamp 1701859473
transform -1 0 3890 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1491_
timestamp 1701859473
transform 1 0 3290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1493_
timestamp 1701859473
transform -1 0 690 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1494_
timestamp 1701859473
transform 1 0 630 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1496_
timestamp 1701859473
transform 1 0 2870 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1498_
timestamp 1701859473
transform 1 0 1010 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1499_
timestamp 1701859473
transform 1 0 2770 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1501_
timestamp 1701859473
transform -1 0 3870 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1503_
timestamp 1701859473
transform -1 0 4010 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1504_
timestamp 1701859473
transform -1 0 3690 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1506_
timestamp 1701859473
transform -1 0 4930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1508_
timestamp 1701859473
transform -1 0 3930 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1510_
timestamp 1701859473
transform -1 0 3250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1511_
timestamp 1701859473
transform 1 0 3190 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1513_
timestamp 1701859473
transform 1 0 3730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1515_
timestamp 1701859473
transform -1 0 3370 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1516_
timestamp 1701859473
transform -1 0 2990 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1518_
timestamp 1701859473
transform -1 0 2710 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1520_
timestamp 1701859473
transform 1 0 3130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1521_
timestamp 1701859473
transform -1 0 3450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1523_
timestamp 1701859473
transform 1 0 3270 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1525_
timestamp 1701859473
transform 1 0 1970 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1526_
timestamp 1701859473
transform 1 0 4170 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1528_
timestamp 1701859473
transform 1 0 4250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1530_
timestamp 1701859473
transform -1 0 4110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1531_
timestamp 1701859473
transform 1 0 4330 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1533_
timestamp 1701859473
transform 1 0 3770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1535_
timestamp 1701859473
transform -1 0 4050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1536_
timestamp 1701859473
transform -1 0 4190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1538_
timestamp 1701859473
transform -1 0 4070 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1540_
timestamp 1701859473
transform -1 0 3830 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1542_
timestamp 1701859473
transform 1 0 2570 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1543_
timestamp 1701859473
transform 1 0 2710 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1545_
timestamp 1701859473
transform -1 0 4250 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1547_
timestamp 1701859473
transform 1 0 4530 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1548_
timestamp 1701859473
transform -1 0 3430 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1550_
timestamp 1701859473
transform -1 0 3310 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1552_
timestamp 1701859473
transform -1 0 1270 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1553_
timestamp 1701859473
transform 1 0 3910 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1555_
timestamp 1701859473
transform 1 0 2270 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1557_
timestamp 1701859473
transform 1 0 2970 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1558_
timestamp 1701859473
transform 1 0 3130 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1560_
timestamp 1701859473
transform 1 0 2670 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1562_
timestamp 1701859473
transform -1 0 3250 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1563_
timestamp 1701859473
transform -1 0 3090 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1565_
timestamp 1701859473
transform -1 0 2910 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1567_
timestamp 1701859473
transform 1 0 3550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1568_
timestamp 1701859473
transform 1 0 4150 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1570_
timestamp 1701859473
transform -1 0 4630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1572_
timestamp 1701859473
transform 1 0 3750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1574_
timestamp 1701859473
transform -1 0 3770 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1575_
timestamp 1701859473
transform -1 0 3610 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1577_
timestamp 1701859473
transform 1 0 4230 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1579_
timestamp 1701859473
transform 1 0 4030 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1580_
timestamp 1701859473
transform 1 0 4950 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1582_
timestamp 1701859473
transform -1 0 4870 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1584_
timestamp 1701859473
transform 1 0 4710 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1585_
timestamp 1701859473
transform 1 0 4990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1587_
timestamp 1701859473
transform 1 0 5370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1589_
timestamp 1701859473
transform 1 0 5070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1590_
timestamp 1701859473
transform 1 0 5610 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1592_
timestamp 1701859473
transform 1 0 4990 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1594_
timestamp 1701859473
transform -1 0 5470 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1595_
timestamp 1701859473
transform -1 0 4850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1597_
timestamp 1701859473
transform 1 0 4450 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1599_
timestamp 1701859473
transform 1 0 5070 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1601_
timestamp 1701859473
transform -1 0 5310 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1602_
timestamp 1701859473
transform 1 0 4790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1604_
timestamp 1701859473
transform 1 0 4230 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1606_
timestamp 1701859473
transform 1 0 4310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1607_
timestamp 1701859473
transform 1 0 4350 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1609_
timestamp 1701859473
transform -1 0 4750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1611_
timestamp 1701859473
transform -1 0 4590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1612_
timestamp 1701859473
transform 1 0 4430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1614_
timestamp 1701859473
transform -1 0 4670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1616_
timestamp 1701859473
transform 1 0 4550 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1617_
timestamp 1701859473
transform 1 0 4510 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1619_
timestamp 1701859473
transform 1 0 6150 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1621_
timestamp 1701859473
transform -1 0 4530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1622_
timestamp 1701859473
transform 1 0 4810 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1624_
timestamp 1701859473
transform -1 0 5450 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1626_
timestamp 1701859473
transform -1 0 5150 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1627_
timestamp 1701859473
transform 1 0 6010 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1629_
timestamp 1701859473
transform 1 0 4810 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1631_
timestamp 1701859473
transform 1 0 5110 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1633_
timestamp 1701859473
transform -1 0 4850 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1634_
timestamp 1701859473
transform -1 0 2450 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1636_
timestamp 1701859473
transform -1 0 4530 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1638_
timestamp 1701859473
transform -1 0 4370 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1639_
timestamp 1701859473
transform -1 0 4950 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1641_
timestamp 1701859473
transform -1 0 4910 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1643_
timestamp 1701859473
transform 1 0 5450 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1644_
timestamp 1701859473
transform 1 0 5030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1646_
timestamp 1701859473
transform 1 0 5270 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1648_
timestamp 1701859473
transform 1 0 5650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1649_
timestamp 1701859473
transform 1 0 5230 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1651_
timestamp 1701859473
transform 1 0 5690 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1653_
timestamp 1701859473
transform 1 0 5310 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1654_
timestamp 1701859473
transform -1 0 5890 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1656_
timestamp 1701859473
transform 1 0 5450 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1658_
timestamp 1701859473
transform 1 0 5210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1660_
timestamp 1701859473
transform -1 0 5230 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1661_
timestamp 1701859473
transform -1 0 5370 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1663_
timestamp 1701859473
transform 1 0 6150 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1665_
timestamp 1701859473
transform -1 0 5610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1666_
timestamp 1701859473
transform 1 0 5570 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1668_
timestamp 1701859473
transform -1 0 6290 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1670_
timestamp 1701859473
transform -1 0 5510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1671_
timestamp 1701859473
transform -1 0 6010 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1673_
timestamp 1701859473
transform 1 0 4030 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1675_
timestamp 1701859473
transform 1 0 5970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1676_
timestamp 1701859473
transform 1 0 6250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1678_
timestamp 1701859473
transform -1 0 6130 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1680_
timestamp 1701859473
transform 1 0 6290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1681_
timestamp 1701859473
transform 1 0 6170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1683_
timestamp 1701859473
transform -1 0 5790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1685_
timestamp 1701859473
transform 1 0 5850 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1686_
timestamp 1701859473
transform -1 0 5510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1688_
timestamp 1701859473
transform 1 0 6050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1690_
timestamp 1701859473
transform 1 0 6150 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1692_
timestamp 1701859473
transform -1 0 5470 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1693_
timestamp 1701859473
transform 1 0 5290 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1695_
timestamp 1701859473
transform -1 0 5550 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1697_
timestamp 1701859473
transform 1 0 5370 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1698_
timestamp 1701859473
transform 1 0 5750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1700_
timestamp 1701859473
transform -1 0 5330 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1702_
timestamp 1701859473
transform 1 0 6030 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1703_
timestamp 1701859473
transform -1 0 5210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1705_
timestamp 1701859473
transform -1 0 5350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1707_
timestamp 1701859473
transform 1 0 5470 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1708_
timestamp 1701859473
transform 1 0 6210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1710_
timestamp 1701859473
transform 1 0 5650 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1712_
timestamp 1701859473
transform -1 0 5090 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1713_
timestamp 1701859473
transform 1 0 4770 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1715_
timestamp 1701859473
transform -1 0 4550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1717_
timestamp 1701859473
transform -1 0 4990 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1719_
timestamp 1701859473
transform 1 0 5290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1720_
timestamp 1701859473
transform -1 0 5510 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1722_
timestamp 1701859473
transform 1 0 4710 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1724_
timestamp 1701859473
transform 1 0 4830 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1725_
timestamp 1701859473
transform 1 0 4970 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1727_
timestamp 1701859473
transform -1 0 5750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1729_
timestamp 1701859473
transform 1 0 5250 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1730_
timestamp 1701859473
transform 1 0 5570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1732_
timestamp 1701859473
transform 1 0 5890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1734_
timestamp 1701859473
transform -1 0 6330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1735_
timestamp 1701859473
transform -1 0 6330 0 -1 5990
box -12 -8 32 272
use FILL  FILL_3__1737_
timestamp 1701859473
transform 1 0 5950 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1739_
timestamp 1701859473
transform -1 0 6190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1740_
timestamp 1701859473
transform 1 0 6210 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1742_
timestamp 1701859473
transform 1 0 6330 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1744_
timestamp 1701859473
transform 1 0 5650 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1745_
timestamp 1701859473
transform 1 0 5630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1747_
timestamp 1701859473
transform 1 0 6130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1749_
timestamp 1701859473
transform 1 0 4790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1751_
timestamp 1701859473
transform 1 0 4370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1752_
timestamp 1701859473
transform 1 0 3950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1754_
timestamp 1701859473
transform 1 0 4390 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1756_
timestamp 1701859473
transform -1 0 4250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1757_
timestamp 1701859473
transform 1 0 5510 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1759_
timestamp 1701859473
transform 1 0 5670 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1761_
timestamp 1701859473
transform 1 0 5930 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1762_
timestamp 1701859473
transform 1 0 6050 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1764_
timestamp 1701859473
transform -1 0 6250 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1766_
timestamp 1701859473
transform -1 0 6170 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1767_
timestamp 1701859473
transform -1 0 6330 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1769_
timestamp 1701859473
transform -1 0 6190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1771_
timestamp 1701859473
transform -1 0 5790 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1772_
timestamp 1701859473
transform 1 0 5610 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1774_
timestamp 1701859473
transform -1 0 6090 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1776_
timestamp 1701859473
transform -1 0 5930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1778_
timestamp 1701859473
transform 1 0 3510 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1779_
timestamp 1701859473
transform 1 0 4550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1781_
timestamp 1701859473
transform 1 0 4670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1783_
timestamp 1701859473
transform 1 0 4970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1784_
timestamp 1701859473
transform -1 0 5050 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1786_
timestamp 1701859473
transform 1 0 5270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1788_
timestamp 1701859473
transform 1 0 5690 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1789_
timestamp 1701859473
transform -1 0 5870 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1791_
timestamp 1701859473
transform -1 0 5870 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1793_
timestamp 1701859473
transform -1 0 5130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1794_
timestamp 1701859473
transform -1 0 4570 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1796_
timestamp 1701859473
transform -1 0 5070 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1798_
timestamp 1701859473
transform -1 0 5530 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1799_
timestamp 1701859473
transform -1 0 5270 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1801_
timestamp 1701859473
transform -1 0 5590 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1803_
timestamp 1701859473
transform -1 0 4530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1804_
timestamp 1701859473
transform -1 0 4370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1806_
timestamp 1701859473
transform 1 0 3950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1808_
timestamp 1701859473
transform 1 0 4230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1810_
timestamp 1701859473
transform -1 0 3650 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1811_
timestamp 1701859473
transform -1 0 4370 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1813_
timestamp 1701859473
transform 1 0 3930 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1815_
timestamp 1701859473
transform 1 0 4050 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1816_
timestamp 1701859473
transform -1 0 4310 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1818_
timestamp 1701859473
transform 1 0 3890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1820_
timestamp 1701859473
transform -1 0 3810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1821_
timestamp 1701859473
transform 1 0 3650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1823_
timestamp 1701859473
transform 1 0 4070 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1825_
timestamp 1701859473
transform 1 0 3170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1826_
timestamp 1701859473
transform 1 0 2890 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1828_
timestamp 1701859473
transform 1 0 2850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1830_
timestamp 1701859473
transform -1 0 2830 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1831_
timestamp 1701859473
transform -1 0 2750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1833_
timestamp 1701859473
transform -1 0 3310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1835_
timestamp 1701859473
transform 1 0 3630 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1836_
timestamp 1701859473
transform -1 0 3310 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1838_
timestamp 1701859473
transform -1 0 3050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1840_
timestamp 1701859473
transform 1 0 2370 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1842_
timestamp 1701859473
transform -1 0 2070 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1843_
timestamp 1701859473
transform -1 0 2210 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1845_
timestamp 1701859473
transform -1 0 2670 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1847_
timestamp 1701859473
transform -1 0 2490 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1848_
timestamp 1701859473
transform 1 0 2830 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1911_
timestamp 1701859473
transform 1 0 6290 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1913_
timestamp 1701859473
transform 1 0 2130 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1914_
timestamp 1701859473
transform 1 0 3670 0 1 5470
box -12 -8 32 272
use FILL  FILL_3__1916_
timestamp 1701859473
transform 1 0 6310 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1918_
timestamp 1701859473
transform 1 0 5870 0 1 5990
box -12 -8 32 272
use FILL  FILL_3__1919_
timestamp 1701859473
transform -1 0 5730 0 1 790
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert0
timestamp 1701859473
transform 1 0 4790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert2
timestamp 1701859473
transform -1 0 4270 0 -1 270
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert4
timestamp 1701859473
transform 1 0 5550 0 1 270
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert12
timestamp 1701859473
transform 1 0 2110 0 1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert14
timestamp 1701859473
transform 1 0 1350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert15
timestamp 1701859473
transform -1 0 1930 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert17
timestamp 1701859473
transform 1 0 3110 0 1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert19
timestamp 1701859473
transform -1 0 3030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert20
timestamp 1701859473
transform 1 0 3950 0 1 1310
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert22
timestamp 1701859473
transform -1 0 5670 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert24
timestamp 1701859473
transform 1 0 4110 0 1 790
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert25
timestamp 1701859473
transform 1 0 4930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert5
timestamp 1701859473
transform 1 0 4950 0 1 1310
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert7
timestamp 1701859473
transform -1 0 4150 0 1 270
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert9
timestamp 1701859473
transform -1 0 3470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert10
timestamp 1701859473
transform 1 0 4690 0 1 1310
box -12 -8 32 272
<< labels >>
flabel metal1 s 6443 2 6503 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal3 s 6476 4596 6484 4604 3 FreeSans 16 0 0 0 Cin[7]
port 2 nsew
flabel metal3 s 6476 4556 6484 4564 3 FreeSans 16 0 0 0 Cin[6]
port 3 nsew
flabel metal3 s 6476 4516 6484 4524 3 FreeSans 16 0 0 0 Cin[5]
port 4 nsew
flabel metal3 s 6476 4376 6484 4384 3 FreeSans 16 0 0 0 Cin[4]
port 5 nsew
flabel metal3 s 6476 4336 6484 4344 3 FreeSans 16 0 0 0 Cin[3]
port 6 nsew
flabel metal2 s 3217 -23 3223 -17 7 FreeSans 16 270 0 0 Cin[2]
port 7 nsew
flabel metal2 s 3177 -23 3183 -17 7 FreeSans 16 270 0 0 Cin[1]
port 8 nsew
flabel metal2 s 1397 -23 1403 -17 7 FreeSans 16 270 0 0 Cin[0]
port 9 nsew
flabel metal2 s 4057 -23 4063 -17 7 FreeSans 16 270 0 0 Rdy
port 10 nsew
flabel metal3 s 6476 656 6484 664 3 FreeSans 16 0 0 0 Vld
port 11 nsew
flabel metal3 s -24 3936 -16 3944 7 FreeSans 16 0 0 0 Xin[3]
port 12 nsew
flabel metal3 s -24 3896 -16 3904 7 FreeSans 16 0 0 0 Xin[2]
port 13 nsew
flabel metal3 s -24 3856 -16 3864 7 FreeSans 16 0 0 0 Xin[1]
port 14 nsew
flabel metal3 s -24 3816 -16 3824 7 FreeSans 16 0 0 0 Xin[0]
port 15 nsew
flabel metal2 s 3837 6297 3843 6303 3 FreeSans 16 90 0 0 Xout[3]
port 16 nsew
flabel metal2 s 3717 6297 3723 6303 3 FreeSans 16 90 0 0 Xout[2]
port 17 nsew
flabel metal2 s 2177 6297 2183 6303 3 FreeSans 16 90 0 0 Xout[1]
port 18 nsew
flabel metal2 s 2137 6297 2143 6303 3 FreeSans 16 90 0 0 Xout[0]
port 19 nsew
flabel metal3 s -24 1956 -16 1964 7 FreeSans 16 0 0 0 Yin[3]
port 20 nsew
flabel metal3 s -24 3776 -16 3784 7 FreeSans 16 0 0 0 Yin[2]
port 21 nsew
flabel metal2 s 3557 -23 3563 -17 7 FreeSans 16 270 0 0 Yin[1]
port 22 nsew
flabel metal2 s 4017 -23 4023 -17 7 FreeSans 16 270 0 0 Yin[0]
port 23 nsew
flabel metal2 s 5757 6297 5763 6303 3 FreeSans 16 90 0 0 Yout[3]
port 24 nsew
flabel metal2 s 5917 6297 5923 6303 3 FreeSans 16 90 0 0 Yout[2]
port 25 nsew
flabel metal3 s 6476 696 6484 704 3 FreeSans 16 0 0 0 Yout[1]
port 26 nsew
flabel metal3 s 6476 916 6484 924 3 FreeSans 16 0 0 0 Yout[0]
port 27 nsew
flabel metal2 s 4137 -23 4143 -17 7 FreeSans 16 270 0 0 clk
port 28 nsew
<< properties >>
string FIXED_BBOX -40 -40 6480 6300
<< end >>
