magic
tech scmos
magscale 1 3
timestamp 1725338204
<< checkpaint >>
rect 10 480 480 505
rect 10 474 505 480
rect -14 16 505 474
rect 10 10 505 16
rect 10 -15 480 10
<< nwell >>
rect 110 110 380 380
<< psubstratepdiff >>
rect 45 425 445 445
rect 45 65 65 425
rect 195 195 295 295
rect 425 65 445 425
rect 45 45 445 65
<< nsubstratendiff >>
rect 130 340 360 360
rect 130 150 150 340
rect 340 150 360 340
rect 130 130 360 150
<< genericcontact >>
rect 70 425 420 445
rect 45 70 65 420
rect 150 340 340 360
rect 130 150 150 340
rect 195 195 295 295
rect 340 150 360 340
rect 150 130 340 150
rect 425 70 445 420
rect 70 45 420 65
<< metal1 >>
rect 45 425 445 445
rect 45 65 65 425
rect 130 340 360 360
rect 130 150 150 340
rect 195 195 295 295
rect 340 150 360 340
rect 130 130 360 150
rect 425 65 445 425
rect 45 45 445 65
<< end >>
