magic
tech scmos
magscale 1 2
timestamp 1728387359
<< nwell >>
rect -12 174 492 252
<< ntransistor >>
rect 24 14 28 54
rect 36 14 40 54
rect 60 14 64 54
rect 72 14 76 54
rect 122 14 126 34
rect 142 14 146 34
rect 162 14 166 34
rect 212 14 216 34
rect 232 14 236 34
rect 277 14 281 34
rect 297 14 301 34
rect 350 14 354 54
rect 362 14 366 54
rect 387 14 391 54
rect 399 14 403 54
rect 447 14 451 34
<< ptransistor >>
rect 22 186 26 226
rect 42 186 46 226
rect 62 186 66 226
rect 82 186 86 226
rect 127 206 131 226
rect 147 206 151 226
rect 167 186 171 226
rect 212 186 216 226
rect 232 186 236 226
rect 277 206 281 226
rect 297 206 301 226
rect 342 186 346 226
rect 362 186 366 226
rect 382 186 386 226
rect 402 186 406 226
rect 447 186 451 226
<< ndiffusion >>
rect 20 14 24 54
rect 28 14 36 54
rect 40 14 44 54
rect 56 14 60 54
rect 64 14 72 54
rect 76 14 80 54
rect 120 14 122 34
rect 126 14 128 34
rect 140 14 142 34
rect 146 14 148 34
rect 160 14 162 34
rect 166 14 168 34
rect 210 14 212 34
rect 216 14 218 34
rect 230 14 232 34
rect 236 14 238 34
rect 275 14 277 34
rect 281 14 283 34
rect 295 14 297 34
rect 301 14 303 34
rect 346 14 350 54
rect 354 14 362 54
rect 366 14 371 54
rect 383 14 387 54
rect 391 14 399 54
rect 403 14 407 54
rect 445 14 447 34
rect 451 14 453 34
<< pdiffusion >>
rect 20 186 22 226
rect 26 186 28 226
rect 40 186 42 226
rect 46 186 48 226
rect 60 186 62 226
rect 66 186 68 226
rect 80 186 82 226
rect 86 203 88 226
rect 125 206 127 226
rect 131 206 133 226
rect 145 206 147 226
rect 151 206 153 226
rect 165 206 167 226
rect 86 186 100 203
rect 155 186 167 206
rect 171 186 173 226
rect 210 186 212 226
rect 216 186 218 226
rect 230 186 232 226
rect 236 186 238 226
rect 275 206 277 226
rect 281 206 283 226
rect 295 206 297 226
rect 301 206 303 226
rect 340 186 342 226
rect 346 186 348 226
rect 360 186 362 226
rect 366 186 368 226
rect 380 186 382 226
rect 386 186 388 226
rect 400 186 402 226
rect 406 186 408 226
rect 445 186 447 226
rect 451 186 453 226
<< ndcontact >>
rect 8 14 20 54
rect 44 14 56 54
rect 80 14 92 54
rect 108 14 120 34
rect 128 14 140 34
rect 148 14 160 34
rect 168 14 180 34
rect 198 14 210 34
rect 218 14 230 34
rect 238 14 250 34
rect 263 14 275 34
rect 283 14 295 34
rect 303 14 315 34
rect 334 14 346 54
rect 371 14 383 54
rect 407 14 419 54
rect 433 14 445 34
rect 453 14 465 34
<< pdcontact >>
rect 8 186 20 226
rect 28 186 40 226
rect 48 186 60 226
rect 68 186 80 226
rect 88 203 100 226
rect 113 206 125 226
rect 133 206 145 226
rect 153 206 165 226
rect 173 186 185 226
rect 198 186 210 226
rect 218 186 230 226
rect 238 186 250 226
rect 263 206 275 226
rect 283 206 295 226
rect 303 206 315 226
rect 328 186 340 226
rect 348 186 360 226
rect 368 186 380 226
rect 388 186 400 226
rect 408 186 420 226
rect 433 186 445 226
rect 453 186 465 226
<< psubstratepcontact >>
rect -6 -6 486 6
<< nsubstratencontact >>
rect -6 234 486 246
<< polysilicon >>
rect 22 226 26 230
rect 42 226 46 230
rect 62 226 66 230
rect 82 226 86 230
rect 127 226 131 230
rect 147 226 151 230
rect 167 226 171 230
rect 212 226 216 230
rect 232 226 236 230
rect 277 226 281 230
rect 297 226 301 230
rect 342 226 346 230
rect 362 226 366 230
rect 382 226 386 230
rect 402 226 406 230
rect 447 226 451 230
rect 22 109 26 186
rect 42 168 46 186
rect 22 97 24 109
rect 24 54 28 97
rect 44 72 48 156
rect 62 151 66 186
rect 36 54 40 60
rect 60 54 64 139
rect 82 131 86 186
rect 82 84 86 119
rect 127 95 131 206
rect 147 121 151 206
rect 146 87 150 109
rect 167 91 171 186
rect 212 105 216 186
rect 232 128 236 186
rect 277 178 281 206
rect 256 166 281 178
rect 232 122 244 128
rect 212 93 219 105
rect 72 80 86 84
rect 122 83 150 87
rect 72 54 76 80
rect 122 34 126 83
rect 162 79 171 91
rect 142 34 146 63
rect 162 34 166 79
rect 212 54 216 93
rect 240 72 244 122
rect 275 88 280 166
rect 297 117 301 206
rect 342 180 346 186
rect 341 168 346 180
rect 300 105 314 117
rect 275 82 301 88
rect 236 66 244 72
rect 192 42 216 54
rect 212 34 216 42
rect 232 34 236 60
rect 277 34 281 60
rect 297 34 301 82
rect 309 72 314 105
rect 330 62 335 168
rect 362 166 366 186
rect 382 180 386 186
rect 350 160 366 166
rect 350 122 356 160
rect 381 150 385 168
rect 370 144 385 150
rect 402 147 406 186
rect 344 70 350 110
rect 370 90 374 144
rect 405 135 406 147
rect 402 104 406 135
rect 372 78 374 90
rect 344 66 366 70
rect 330 58 354 62
rect 350 54 354 58
rect 362 54 366 66
rect 370 62 374 78
rect 380 98 406 104
rect 380 70 384 98
rect 447 90 451 186
rect 404 78 451 90
rect 380 66 403 70
rect 370 58 391 62
rect 387 54 391 58
rect 399 54 403 66
rect 447 34 451 78
rect 24 10 28 14
rect 36 10 40 14
rect 60 10 64 14
rect 72 10 76 14
rect 122 10 126 14
rect 142 10 146 14
rect 162 10 166 14
rect 212 10 216 14
rect 232 10 236 14
rect 277 10 281 14
rect 297 10 301 14
rect 350 10 354 14
rect 362 10 366 14
rect 387 10 391 14
rect 399 10 403 14
rect 447 10 451 14
<< polycontact >>
rect 38 156 50 168
rect 24 97 36 109
rect 36 60 48 72
rect 60 139 72 151
rect 77 119 89 131
rect 115 95 127 107
rect 146 109 158 121
rect 244 166 256 178
rect 219 93 231 105
rect 171 79 183 91
rect 137 63 149 75
rect 329 168 341 180
rect 288 105 300 117
rect 224 60 236 72
rect 276 60 288 72
rect 180 42 192 54
rect 309 60 321 72
rect 374 168 386 180
rect 344 110 356 122
rect 393 135 405 147
rect 360 78 372 90
rect 392 78 404 90
<< metal1 >>
rect -6 246 486 248
rect -6 232 486 234
rect 8 226 20 232
rect 48 226 60 232
rect 88 226 100 232
rect 173 226 185 232
rect 218 226 230 232
rect 328 226 340 232
rect 368 226 380 232
rect 408 226 420 232
rect 453 226 465 232
rect 109 206 113 226
rect 131 206 133 226
rect 152 206 153 226
rect 109 197 117 206
rect 131 197 137 206
rect 152 197 160 206
rect 28 180 35 186
rect 8 174 35 180
rect 8 84 16 174
rect 68 168 80 186
rect 157 186 160 197
rect 201 180 210 186
rect 238 180 250 186
rect 201 169 203 180
rect 50 161 156 168
rect 244 178 250 180
rect 72 143 123 151
rect 143 154 156 161
rect 264 159 273 206
rect 283 183 295 206
rect 304 198 314 206
rect 348 180 360 186
rect 297 169 329 177
rect 348 172 374 180
rect 392 159 400 186
rect 143 145 263 154
rect 317 153 419 159
rect 323 139 393 147
rect 143 133 330 139
rect 65 131 330 133
rect 89 127 156 131
rect 95 113 140 119
rect 95 97 103 113
rect 24 90 103 97
rect 133 103 140 113
rect 158 113 203 121
rect 217 117 300 125
rect 133 97 213 103
rect 8 78 110 84
rect 8 54 16 78
rect 48 60 92 68
rect 82 54 92 60
rect 103 57 110 78
rect 120 72 127 95
rect 206 87 213 97
rect 309 110 344 122
rect 309 99 315 110
rect 363 104 377 117
rect 251 92 315 99
rect 322 97 377 104
rect 251 87 257 92
rect 206 78 257 87
rect 322 85 329 97
rect 263 78 329 85
rect 352 78 360 90
rect 372 78 392 90
rect 120 64 137 72
rect 263 72 270 78
rect 149 63 171 69
rect 165 54 171 63
rect 236 60 270 72
rect 288 60 309 72
rect 352 54 362 78
rect 411 54 419 153
rect 165 45 180 54
rect 108 34 117 43
rect 128 34 137 43
rect 148 34 157 43
rect 198 40 203 52
rect 245 40 250 52
rect 198 34 210 40
rect 238 34 250 40
rect 263 34 275 40
rect 283 34 295 40
rect 303 34 315 40
rect 346 46 362 54
rect 433 34 443 186
rect 44 8 56 14
rect 168 8 180 14
rect 218 8 230 14
rect 371 8 383 14
rect 453 8 465 14
rect -6 6 486 8
rect -6 -8 486 -6
<< m2contact >>
rect 103 183 117 197
rect 123 183 137 197
rect 143 183 157 197
rect 203 166 217 180
rect 230 166 244 180
rect 123 141 137 155
rect 304 184 318 198
rect 283 169 297 183
rect 263 145 277 159
rect 303 145 317 159
rect 23 109 37 123
rect 63 117 77 131
rect 203 111 217 125
rect 183 77 197 91
rect 231 93 245 107
rect 363 117 377 131
rect 103 43 117 57
rect 123 43 137 57
rect 143 43 157 57
rect 203 40 217 54
rect 231 40 245 54
rect 263 40 277 54
rect 283 40 297 54
rect 303 40 317 54
rect 443 89 457 103
<< metal2 >>
rect 23 123 37 137
rect 63 103 77 117
rect 107 57 115 183
rect 127 155 135 183
rect 127 57 135 141
rect 147 57 155 183
rect 205 125 213 166
rect 183 63 197 77
rect 205 54 213 111
rect 233 107 241 166
rect 233 54 241 93
rect 266 54 274 145
rect 287 54 295 169
rect 305 159 313 184
rect 305 54 313 145
rect 363 103 377 117
rect 443 103 457 117
<< m1p >>
rect -6 232 486 248
rect -6 -8 486 8
<< m2p >>
rect 23 123 37 137
rect 63 103 77 117
rect 363 103 377 117
rect 443 103 457 117
rect 183 63 197 77
<< labels >>
rlabel metal1 -6 -8 486 8 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal1 -6 232 486 248 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal2 63 103 77 117 0 S
port 1 nsew signal input
rlabel metal2 183 63 197 77 0 D
port 2 nsew signal input
rlabel metal2 363 103 377 117 0 CLK
port 3 nsew signal input
rlabel metal2 23 123 37 137 0 R
port 0 nsew signal input
rlabel metal2 443 103 457 117 0 Q
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 480 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
