magic
tech scmos
magscale 1 2
timestamp 1727572430
<< nwell >>
rect -12 154 112 272
<< ntransistor >>
rect 20 14 24 54
rect 30 14 34 54
rect 52 14 56 34
<< ptransistor >>
rect 20 206 24 246
rect 40 206 44 246
rect 60 206 64 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 14 30 54
rect 34 14 36 54
rect 48 14 52 34
rect 56 14 58 34
<< pdiffusion >>
rect 18 206 20 246
rect 24 206 26 246
rect 38 206 40 246
rect 44 206 46 246
rect 58 206 60 246
rect 64 206 66 246
<< ndcontact >>
rect 6 14 18 54
rect 36 14 48 54
rect 58 14 70 34
<< pdcontact >>
rect 6 206 18 246
rect 26 206 38 246
rect 46 206 58 246
rect 66 206 78 246
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 254 106 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 20 103 24 206
rect 40 129 44 206
rect 60 202 64 206
rect 60 198 68 202
rect 16 91 24 103
rect 20 54 24 91
rect 30 117 44 129
rect 30 54 34 117
rect 64 72 68 198
rect 56 66 68 72
rect 52 34 56 60
rect 20 10 24 14
rect 30 10 34 14
rect 52 10 56 14
<< polycontact >>
rect 4 91 16 103
rect 44 117 56 129
rect 44 60 56 72
<< metal1 >>
rect -6 266 106 268
rect -6 252 106 254
rect 6 246 18 252
rect 46 246 58 252
rect 27 72 34 206
rect 66 137 74 206
rect 6 64 44 72
rect 6 54 18 64
rect 63 39 70 123
rect 58 34 70 39
rect 36 8 48 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m2contact >>
rect 3 103 17 117
rect 63 123 77 137
rect 43 103 57 117
<< metal2 >>
rect 63 137 77 157
rect 3 117 17 137
rect 43 83 57 103
<< m2p >>
rect 63 143 77 157
rect 3 123 17 137
rect 43 83 57 97
<< labels >>
rlabel metal2 3 123 17 137 0 A
port 0 nsew signal input
rlabel metal2 43 83 57 97 0 B
port 1 nsew signal input
rlabel metal2 63 143 77 157 0 Y
port 2 nsew signal output
rlabel metal1 -6 252 106 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -6 -8 106 8 0 gnd
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
