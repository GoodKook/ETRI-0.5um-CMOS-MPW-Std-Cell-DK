magic
tech scmos
magscale 1 6
timestamp 1569139307
<< checkpaint >>
rect -120 -120 2520 5180
<< metal1 >>
rect 207 3660 429 3700
rect 459 3660 2340 3720
rect 120 1400 284 1440
rect 393 1400 2340 1460
<< metal2 >>
rect 112 4644 152 5060
rect 112 4606 298 4644
rect 472 4200 540 4312
rect 100 4160 540 4200
rect 0 2260 80 3820
rect 12 1560 80 2160
rect 0 0 80 1560
rect 100 1440 120 4160
rect 302 3660 374 4160
rect 100 1400 195 1440
rect 264 140 372 3640
rect 516 140 624 3640
rect 768 140 876 3640
rect 1020 140 1128 3640
rect 1272 140 1380 3640
rect 1524 140 1632 3640
rect 1776 140 1884 3640
rect 2028 140 2136 3640
rect 2300 2260 2400 3820
rect 2300 1660 2388 2260
rect 264 0 2136 140
rect 2300 0 2400 1560
use VIA1  VIA1_0
timestamp 1569139307
transform 1 0 354 0 1 3680
box -8 -8 8 8
use VIA1  VIA1_1
timestamp 1569139307
transform 1 0 322 0 1 3680
box -8 -8 8 8
use VIA1  VIA1_2
array 0 1 32 0 0 0
timestamp 1569139307
transform 1 0 140 0 1 1420
box -8 -8 8 8
use VIA1  VIA1_3
array 0 1 36 0 4 36
timestamp 1569139307
transform 1 0 2325 0 1 1691
box -8 -8 8 8
use VIA1  VIA1_4
array 0 0 0 0 4 32
timestamp 1569139307
transform 1 0 45 0 1 1998
box -8 -8 8 8
<< end >>
