magic
tech scmos
magscale 1 3
timestamp 1569140870
<< checkpaint >>
rect -58 -58 202 182
<< polysilicon >>
rect 2 2 142 122
<< pseudo_rpoly2 >>
rect 12 12 112 112
use poly1cont_CDNS_723012252915  poly1cont_CDNS_723012252915_0
timestamp 1569140870
transform 1 0 120 0 1 16
box 0 0 18 92
use poly2cont_CDNS_723012252916  poly2cont_CDNS_723012252916_0
timestamp 1569140870
transform 1 0 16 0 1 16
box 0 0 92 92
<< end >>
