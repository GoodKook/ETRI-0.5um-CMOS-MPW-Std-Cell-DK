magic
tech scmos
timestamp 1700315010
<< checkpaint >>
rect -23 107 33 153
rect -23 -23 33 23
<< nwell >>
rect -6 77 16 136
<< psubstratepcontact >>
rect -3 -3 13 3
<< nsubstratencontact >>
rect -3 127 13 133
<< metal1 >>
rect -3 133 13 134
rect -3 126 13 127
rect -3 3 13 4
rect -3 -4 13 -3
<< m1p >>
rect -3 126 13 134
rect -3 -4 13 4
<< labels >>
rlabel metal1 -3 -4 13 4 0 gnd
port 2 nsew ground bidirectional abutment
rlabel nsubstratencontact 3 129 3 129 0 vdd
port 3 nsew power bidirectional abutment
rlabel psubstratepcontact 4 0 4 0 0 gnd
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 10 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
