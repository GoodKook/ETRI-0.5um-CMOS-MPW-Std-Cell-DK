* NGSPICE file created from ALU8_Mult.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL vdd gnd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A Y vdd gnd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 D CLK Q vdd gnd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S Y vdd gnd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A Y vdd gnd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A Y vdd gnd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR R S D CLK Q vdd gnd
.ends

.subckt ALU8_Mult gnd vdd ABCmd_i[7] ABCmd_i[6] ABCmd_i[5] ABCmd_i[4] ABCmd_i[3] ABCmd_i[2]
+ ABCmd_i[1] ABCmd_i[0] ACC_o[7] ACC_o[6] ACC_o[5] ACC_o[4] ACC_o[3] ACC_o[2] ACC_o[1]
+ ACC_o[0] Flag_i LoadA_i LoadB_i LoadCmd_i MulH_i MulL_i clk reset
XFILL_0__1828_ vdd gnd FILL
XFILL_0__1759_ vdd gnd FILL
XFILL_2__992_ vdd gnd FILL
XFILL_1__1104_ vdd gnd FILL
XFILL86250x68550 vdd gnd FILL
XFILL_1__1035_ vdd gnd FILL
XFILL_1__1868_ vdd gnd FILL
XFILL_1__1799_ vdd gnd FILL
XFILL_2__1213_ vdd gnd FILL
XFILL_0__1613_ vdd gnd FILL
XFILL_0__1544_ vdd gnd FILL
X_1270_ _1358_/A _1270_/B _1278_/B vdd gnd NAND2X1
XFILL_0__1475_ vdd gnd FILL
X_1606_ _1686_/A _1608_/B vdd gnd INVX1
X_1399_ _1439_/B _1462_/A vdd gnd INVX1
X_1468_ _1468_/A _1468_/B _1468_/C _1469_/B vdd gnd AOI21X1
X_1537_ _1567_/A _1537_/B _1539_/B vdd gnd NAND2X1
XFILL_1__1722_ vdd gnd FILL
XFILL_1__1584_ vdd gnd FILL
X_981_ _981_/A _982_/C _992_/A vdd gnd NOR2X1
XFILL_1__1018_ vdd gnd FILL
XFILL_0__1260_ vdd gnd FILL
XFILL_0__1191_ vdd gnd FILL
X_1322_ _1322_/A _1322_/B _1322_/C _1409_/A vdd gnd NAND3X1
XFILL_1__993_ vdd gnd FILL
X_1253_ _1253_/A _1253_/B _1352_/C _1257_/C vdd gnd OAI21X1
XFILL_0__1527_ vdd gnd FILL
X_1184_ _1530_/A _1530_/C _1530_/B _1529_/A vdd gnd NOR3X1
XFILL_0__1458_ vdd gnd FILL
XFILL_0__1389_ vdd gnd FILL
XFILL_1__1636_ vdd gnd FILL
XFILL_1__1705_ vdd gnd FILL
XFILL_1__1498_ vdd gnd FILL
XFILL_1__1567_ vdd gnd FILL
X_964_ _980_/A _964_/B _964_/C _973_/B vdd gnd NAND3X1
XFILL_0__1312_ vdd gnd FILL
XFILL_0__1174_ vdd gnd FILL
X_1871_ _1871_/A _1871_/B _1871_/C _1873_/B vdd gnd AOI21X1
XFILL_0__1243_ vdd gnd FILL
X_1305_ _923_/A _958_/C _977_/A _1319_/A vdd gnd NAND3X1
X_1236_ _1236_/A _1236_/B _1236_/C _1340_/C vdd gnd OAI21X1
XFILL_1__976_ vdd gnd FILL
XFILL_1__1421_ vdd gnd FILL
X_1167_ _1265_/B _1265_/A _1190_/C vdd gnd AND2X2
X_1098_ _1113_/C _1113_/A _1113_/B _1246_/C vdd gnd AOI21X1
XFILL_1__1352_ vdd gnd FILL
XFILL_1__1283_ vdd gnd FILL
XFILL_2__1461_ vdd gnd FILL
XFILL_1__1619_ vdd gnd FILL
XFILL_0__994_ vdd gnd FILL
X_947_ _971_/A _971_/B _957_/C _955_/A vdd gnd NAND3X1
XFILL_0__1861_ vdd gnd FILL
XFILL_2__1728_ vdd gnd FILL
XFILL_0__1792_ vdd gnd FILL
X_1021_ _1101_/B _1022_/B vdd gnd INVX1
XFILL_0__1157_ vdd gnd FILL
X_1854_ _1854_/A _1854_/B _1871_/B _1858_/B vdd gnd OAI21X1
X_1785_ _958_/C _1787_/B _1786_/C vdd gnd NAND2X1
XFILL_0__1226_ vdd gnd FILL
XFILL_0__1088_ vdd gnd FILL
XFILL_1__1404_ vdd gnd FILL
XFILL_1__959_ vdd gnd FILL
X_1219_ _1297_/A _1297_/B _1294_/C _1237_/B vdd gnd NAND3X1
XFILL_1__1335_ vdd gnd FILL
XFILL_1__1266_ vdd gnd FILL
XFILL_1__1197_ vdd gnd FILL
XFILL_0__977_ vdd gnd FILL
XFILL_0__1011_ vdd gnd FILL
X_1570_ _1833_/Y _1594_/A _1571_/C vdd gnd NAND2X1
XFILL_0__1844_ vdd gnd FILL
XFILL_0__1775_ vdd gnd FILL
X_1004_ _1062_/A _964_/B _958_/C _1070_/A vdd gnd NAND3X1
XFILL_1__1120_ vdd gnd FILL
XFILL_0__1209_ vdd gnd FILL
X_1768_ _1809_/A _980_/B _1842_/C _1769_/C vdd gnd OAI21X1
X_1837_ _1837_/A _1843_/B _1840_/B vdd gnd AND2X2
XFILL_1__1051_ vdd gnd FILL
XFILL_1__1884_ vdd gnd FILL
X_1699_ _1744_/A _1729_/B _1863_/A _1732_/B vdd gnd OAI21X1
XFILL_1__1318_ vdd gnd FILL
XFILL_1__1249_ vdd gnd FILL
XFILL_0__1560_ vdd gnd FILL
XFILL_0__1491_ vdd gnd FILL
X_1622_ ABCmd_i[1] LoadA_i _1623_/C vdd gnd NAND2X1
XFILL_1_CLKBUF1_insert0 vdd gnd FILL
X_1553_ _1554_/A _1553_/B _1556_/B vdd gnd NAND2X1
XFILL_2_BUFX2_insert14 vdd gnd FILL
X_1484_ Flag_i _1776_/Y _1592_/C _1485_/C vdd gnd OAI21X1
XFILL_0__1758_ vdd gnd FILL
XFILL_0__1689_ vdd gnd FILL
XFILL_0__1827_ vdd gnd FILL
XFILL_1__1034_ vdd gnd FILL
XFILL_1__1103_ vdd gnd FILL
XFILL_1__1867_ vdd gnd FILL
XFILL_1__1798_ vdd gnd FILL
XFILL_0__1543_ vdd gnd FILL
XFILL_0__1612_ vdd gnd FILL
XFILL_0__1474_ vdd gnd FILL
X_1605_ LoadCmd_i _1605_/B _1605_/C _1655_/D vdd gnd OAI21X1
X_1536_ _920_/Y _1536_/B _1536_/C _1665_/D vdd gnd OAI21X1
X_1398_ _1408_/A _1410_/C _1409_/A _1439_/B vdd gnd NAND3X1
X_1467_ _1519_/A _1519_/B _1525_/A vdd gnd NAND2X1
XFILL_1__1652_ vdd gnd FILL
XFILL_1__1583_ vdd gnd FILL
XFILL_1__1721_ vdd gnd FILL
XFILL_1__1017_ vdd gnd FILL
X_980_ _980_/A _980_/B _980_/C _982_/C vdd gnd NAND3X1
XFILL_2__1761_ vdd gnd FILL
XFILL85650x46950 vdd gnd FILL
XFILL_0__1190_ vdd gnd FILL
X_1321_ _1321_/A _1410_/A _1322_/B vdd gnd NOR2X1
XFILL_1__992_ vdd gnd FILL
X_1252_ _1352_/A _1352_/B _1285_/A _1257_/B vdd gnd NAND3X1
XFILL_0__1457_ vdd gnd FILL
X_1183_ _1183_/A _1183_/B _1183_/C _1530_/A vdd gnd AOI21X1
XFILL_0__1526_ vdd gnd FILL
XFILL_0__1388_ vdd gnd FILL
X_1519_ _1519_/A _1519_/B _1519_/C _1525_/B vdd gnd OAI21X1
XFILL_1__1635_ vdd gnd FILL
XFILL_1__1704_ vdd gnd FILL
XFILL_1__1566_ vdd gnd FILL
XFILL_1__1497_ vdd gnd FILL
X_963_ _963_/A _963_/B _967_/A _999_/A vdd gnd OAI21X1
XFILL_2__1813_ vdd gnd FILL
XFILL_0__1311_ vdd gnd FILL
X_1870_ _1870_/A _1870_/B _1870_/C _1888_/A vdd gnd OAI21X1
XFILL_2__1109_ vdd gnd FILL
XFILL_0__1242_ vdd gnd FILL
XFILL_0__1173_ vdd gnd FILL
X_1304_ _1332_/B _1332_/A _1405_/A vdd gnd NAND2X1
XFILL_1__1420_ vdd gnd FILL
X_1166_ _1166_/A _1166_/B _1166_/C _1265_/B vdd gnd NAND3X1
X_1235_ _1340_/A _1340_/B _1289_/C _1248_/A vdd gnd NAND3X1
XFILL_1__975_ vdd gnd FILL
XFILL_0__1509_ vdd gnd FILL
XFILL_1__1351_ vdd gnd FILL
X_1097_ _1209_/A _1236_/C _1236_/A _1113_/A vdd gnd NAND3X1
XFILL_1__1282_ vdd gnd FILL
XFILL_1__1618_ vdd gnd FILL
XFILL_1__1549_ vdd gnd FILL
XFILL_0__993_ vdd gnd FILL
XFILL_0__1860_ vdd gnd FILL
X_946_ _946_/A _946_/B _946_/C _971_/B vdd gnd OAI21X1
XFILL_0__1791_ vdd gnd FILL
X_1020_ _935_/A _982_/B _1080_/A _1101_/B vdd gnd OAI21X1
XFILL_0__1156_ vdd gnd FILL
X_1853_ _1874_/B _1874_/A _1854_/B vdd gnd NOR2X1
XFILL_0__1087_ vdd gnd FILL
X_1784_ _1837_/A _979_/B _1787_/B vdd gnd AND2X2
XFILL_0__1225_ vdd gnd FILL
XFILL_1__1403_ vdd gnd FILL
XFILL_1__958_ vdd gnd FILL
X_1218_ _1643_/B _963_/B _1218_/C _1297_/B vdd gnd OAI21X1
X_1149_ _964_/B _977_/B _1172_/B vdd gnd NAND2X1
XFILL_1__1196_ vdd gnd FILL
XFILL_1__1334_ vdd gnd FILL
XFILL_1__1265_ vdd gnd FILL
XFILL_0__1010_ vdd gnd FILL
XFILL_0__976_ vdd gnd FILL
XFILL_0__1843_ vdd gnd FILL
X_929_ _980_/A _958_/B _980_/C _930_/B vdd gnd NAND3X1
XFILL_0__1774_ vdd gnd FILL
X_1003_ _1007_/A _1008_/C _1070_/B vdd gnd AND2X2
XFILL_1__1050_ vdd gnd FILL
XFILL_0__1139_ vdd gnd FILL
X_1836_ _1836_/A _1836_/B _1841_/C vdd gnd NAND2X1
X_1767_ _1767_/A _1767_/B _1767_/C _1771_/A vdd gnd OAI21X1
X_1698_ _975_/B _1863_/A vdd gnd INVX1
XFILL_0__1208_ vdd gnd FILL
XFILL_1__1883_ vdd gnd FILL
XFILL86850x75750 vdd gnd FILL
XFILL_1__1317_ vdd gnd FILL
XFILL_1__1248_ vdd gnd FILL
XFILL_1__1179_ vdd gnd FILL
XFILL_0__1490_ vdd gnd FILL
XFILL_2__1357_ vdd gnd FILL
XFILL_1_CLKBUF1_insert1 vdd gnd FILL
X_1552_ _1555_/B _1555_/C _1553_/B vdd gnd NAND2X1
XFILL_0__959_ vdd gnd FILL
X_1621_ LoadA_i _953_/A _1621_/C _1669_/D vdd gnd OAI21X1
X_1483_ _1889_/Y _1485_/B vdd gnd INVX1
XFILL_0__1826_ vdd gnd FILL
XFILL_0__1757_ vdd gnd FILL
XFILL_0__1688_ vdd gnd FILL
XFILL_1__1033_ vdd gnd FILL
XFILL_1__1102_ vdd gnd FILL
XFILL86850x50550 vdd gnd FILL
X_1819_ _1881_/B _1824_/B vdd gnd INVX1
XFILL_1__1866_ vdd gnd FILL
XFILL_1__1797_ vdd gnd FILL
XFILL_2__1409_ vdd gnd FILL
XFILL_0__1473_ vdd gnd FILL
XFILL_0__1611_ vdd gnd FILL
XFILL_0__1542_ vdd gnd FILL
X_1604_ LoadCmd_i ABCmd_i[2] _1605_/C vdd gnd NAND2X1
XFILL_1__1720_ vdd gnd FILL
X_1535_ _920_/Y _1535_/B _1536_/C vdd gnd NAND2X1
X_1466_ _1488_/C _1470_/A _1519_/B vdd gnd NAND2X1
X_1397_ _1409_/A _1408_/A _1410_/C _1460_/A vdd gnd AOI21X1
XFILL_1__1651_ vdd gnd FILL
XFILL_1__1582_ vdd gnd FILL
XFILL_0__1809_ vdd gnd FILL
XFILL_1__1016_ vdd gnd FILL
XFILL_1__1849_ vdd gnd FILL
XFILL_2__1056_ vdd gnd FILL
X_1320_ _1378_/A _1378_/B _1320_/C _1322_/C vdd gnd NAND3X1
XFILL_1__991_ vdd gnd FILL
X_1182_ _1428_/B _1480_/A _1480_/B _1530_/C vdd gnd NAND3X1
X_1251_ _1286_/A _1353_/A vdd gnd INVX1
XFILL_0__1456_ vdd gnd FILL
XFILL_0__1525_ vdd gnd FILL
XFILL_0__1387_ vdd gnd FILL
X_1518_ _1519_/A _1519_/B _1518_/C _1584_/A vdd gnd OAI21X1
X_1449_ _977_/A _1577_/A _1495_/A vdd gnd NAND2X1
XFILL_1__1703_ vdd gnd FILL
XFILL_1__1634_ vdd gnd FILL
XFILL_1__1496_ vdd gnd FILL
XFILL_1__1565_ vdd gnd FILL
X_962_ _962_/A _962_/B _963_/B vdd gnd NAND2X1
XFILL_0__1310_ vdd gnd FILL
XFILL_0__1241_ vdd gnd FILL
XFILL_0__1172_ vdd gnd FILL
XFILL_1__974_ vdd gnd FILL
X_1303_ _1303_/A _1367_/B _1367_/A _1332_/A vdd gnd OAI21X1
XFILL_1__1350_ vdd gnd FILL
X_1096_ _1209_/C _1236_/B _1209_/B _1113_/C vdd gnd OAI21X1
X_1165_ _997_/Y _1166_/C vdd gnd INVX1
X_1234_ _1329_/C _1336_/B _1336_/A _1340_/B vdd gnd NAND3X1
XFILL_0__1508_ vdd gnd FILL
XFILL_0__1439_ vdd gnd FILL
XFILL_1__1281_ vdd gnd FILL
XFILL_1__1617_ vdd gnd FILL
XFILL_1__1548_ vdd gnd FILL
XFILL_1__1479_ vdd gnd FILL
XFILL_0__992_ vdd gnd FILL
X_945_ _962_/A _964_/C _946_/B vdd gnd NAND2X1
XFILL_0__1790_ vdd gnd FILL
XFILL_0__1224_ vdd gnd FILL
X_1852_ _1852_/A _1852_/B _1856_/B vdd gnd NOR2X1
XFILL_0__1155_ vdd gnd FILL
XFILL_0__1086_ vdd gnd FILL
X_1783_ _1836_/A _962_/B _1788_/C vdd gnd NAND2X1
XFILL_1__957_ vdd gnd FILL
XFILL_1__1402_ vdd gnd FILL
X_1148_ _1148_/A _1148_/B _1171_/B vdd gnd NAND2X1
X_1079_ _1645_/B _946_/B _1079_/C _1201_/C vdd gnd OAI21X1
X_1217_ _980_/B _1643_/B vdd gnd INVX1
XFILL_1__1333_ vdd gnd FILL
XFILL_1__1264_ vdd gnd FILL
XFILL_1__1195_ vdd gnd FILL
XFILL_2__1442_ vdd gnd FILL
XFILL_0__975_ vdd gnd FILL
X_928_ _962_/A _961_/A _964_/C _935_/C vdd gnd NAND3X1
XFILL_0__1773_ vdd gnd FILL
XFILL_2__1709_ vdd gnd FILL
XFILL_0__1842_ vdd gnd FILL
X_1002_ _1007_/A _1008_/C _1057_/C vdd gnd NOR2X1
X_1835_ _1866_/A _1866_/B _1861_/B _1854_/A vdd gnd AOI21X1
XFILL_0__1207_ vdd gnd FILL
XFILL_0__1138_ vdd gnd FILL
XFILL_0__1069_ vdd gnd FILL
XFILL_1__1882_ vdd gnd FILL
X_1766_ _964_/C _1766_/B _1863_/B _1767_/A vdd gnd OAI21X1
X_1697_ _961_/A _1729_/B vdd gnd INVX1
XFILL_1__1316_ vdd gnd FILL
XFILL_1__1247_ vdd gnd FILL
XFILL_1__1178_ vdd gnd FILL
XFILL_0__958_ vdd gnd FILL
XFILL_1_CLKBUF1_insert2 vdd gnd FILL
X_1551_ _1551_/A _1551_/B _1576_/B _1555_/B vdd gnd OAI21X1
X_1620_ ABCmd_i[0] LoadA_i _1621_/C vdd gnd NAND2X1
X_1482_ _1482_/A _1482_/B _1482_/C _1486_/B vdd gnd AOI21X1
XFILL_0__1756_ vdd gnd FILL
XFILL_0__1825_ vdd gnd FILL
XFILL_1__1101_ vdd gnd FILL
XFILL_0__1687_ vdd gnd FILL
X_1818_ _1818_/A _1818_/B _1866_/B _1874_/A vdd gnd OAI21X1
XFILL_1__1032_ vdd gnd FILL
XFILL_1__1865_ vdd gnd FILL
X_1749_ _1750_/A _964_/B _1842_/C _1750_/C vdd gnd OAI21X1
XFILL_1__1796_ vdd gnd FILL
XFILL_2__1141_ vdd gnd FILL
XFILL_0__1610_ vdd gnd FILL
XFILL_0__1472_ vdd gnd FILL
XFILL_0__1541_ vdd gnd FILL
X_1465_ _1465_/A _1465_/B _1465_/C _1488_/C vdd gnd NAND3X1
X_1534_ _1534_/A _1534_/B _1534_/C _1535_/B vdd gnd OAI21X1
X_1603_ _1843_/A _1605_/B vdd gnd INVX1
XFILL_1__1650_ vdd gnd FILL
X_1396_ _1396_/A _1396_/B _1410_/C vdd gnd NAND2X1
XFILL_1__1581_ vdd gnd FILL
XFILL_0__1739_ vdd gnd FILL
XFILL_0__1808_ vdd gnd FILL
XFILL_2__972_ vdd gnd FILL
XFILL_1__1015_ vdd gnd FILL
XFILL_1__1779_ vdd gnd FILL
XFILL_1__1848_ vdd gnd FILL
XFILL_1__990_ vdd gnd FILL
XFILL_0__1524_ vdd gnd FILL
X_1181_ _1181_/A _1181_/B _1181_/C _1480_/B vdd gnd OAI21X1
X_1250_ _1353_/C _1286_/B _1286_/A _1255_/B vdd gnd AOI21X1
XFILL_0__1455_ vdd gnd FILL
XFILL_0__1386_ vdd gnd FILL
XFILL_1__1633_ vdd gnd FILL
X_1448_ _1491_/C _1490_/A _1448_/C _1455_/A vdd gnd AOI21X1
X_1517_ _1525_/A _1517_/B _1518_/C vdd gnd NAND2X1
XFILL_1__1702_ vdd gnd FILL
X_1379_ _1629_/B _1548_/D _1382_/A _1380_/B vdd gnd OAI21X1
XFILL_1__1495_ vdd gnd FILL
XFILL_1__1564_ vdd gnd FILL
X_961_ _961_/A _963_/A vdd gnd INVX1
XFILL_0__1240_ vdd gnd FILL
XFILL_0__1171_ vdd gnd FILL
XFILL_1__973_ vdd gnd FILL
X_1302_ _1302_/A _1302_/B _1367_/B vdd gnd AND2X2
X_1233_ _1410_/A _1233_/B _1233_/C _1336_/B vdd gnd OAI21X1
XFILL_0__1507_ vdd gnd FILL
X_1164_ _1567_/A _1265_/C vdd gnd INVX1
X_1095_ _1095_/A _1095_/B _1095_/C _1113_/B vdd gnd AOI21X1
XFILL_1__1280_ vdd gnd FILL
XFILL_0__1438_ vdd gnd FILL
XFILL_0__1369_ vdd gnd FILL
XFILL_1__1616_ vdd gnd FILL
XFILL_0__991_ vdd gnd FILL
XFILL_1__1547_ vdd gnd FILL
XFILL_1__1478_ vdd gnd FILL
XFILL85950x50550 vdd gnd FILL
X_944_ _958_/B _946_/A vdd gnd INVX1
XFILL_0__1154_ vdd gnd FILL
X_1851_ _1851_/A _1851_/B _1852_/A vdd gnd NAND2X1
XFILL_0__1223_ vdd gnd FILL
X_1782_ _1782_/A _1782_/B _1782_/C _1797_/C vdd gnd AOI21X1
XFILL_0__1085_ vdd gnd FILL
XFILL_1__956_ vdd gnd FILL
X_1216_ _1218_/C _1216_/B _1294_/C vdd gnd OR2X2
XFILL_1__1401_ vdd gnd FILL
X_1147_ _1147_/A _1148_/B vdd gnd INVX1
X_1078_ _962_/A _980_/B _958_/C _1079_/C vdd gnd NAND3X1
XFILL_1__1332_ vdd gnd FILL
XFILL_1__1263_ vdd gnd FILL
XFILL_1__1194_ vdd gnd FILL
XFILL_0__974_ vdd gnd FILL
X_927_ _953_/C _927_/B _997_/A vdd gnd OR2X2
XFILL_0__1772_ vdd gnd FILL
XFILL_0__1841_ vdd gnd FILL
X_1001_ _1062_/A _961_/A _1823_/A _1008_/C vdd gnd NAND3X1
XFILL_0__1137_ vdd gnd FILL
X_1834_ _1859_/A _1874_/C vdd gnd INVX1
X_1765_ _1839_/A _980_/B _1765_/C _1839_/D _1767_/B vdd gnd AOI22X1
XFILL_0__1206_ vdd gnd FILL
XFILL_0__1068_ vdd gnd FILL
XFILL_1__1881_ vdd gnd FILL
XFILL86850x10950 vdd gnd FILL
X_1696_ _1836_/A _1863_/B vdd gnd INVX2
XFILL_1__939_ vdd gnd FILL
XFILL_1__1315_ vdd gnd FILL
XFILL_1__1246_ vdd gnd FILL
XFILL_1__1177_ vdd gnd FILL
XFILL_1_CLKBUF1_insert3 vdd gnd FILL
XFILL_0__957_ vdd gnd FILL
X_1550_ _1576_/A _1576_/B _1555_/C vdd gnd OR2X2
X_1481_ _1482_/A _1482_/B MulL_i _1482_/C vdd gnd OAI21X1
XFILL_0__1686_ vdd gnd FILL
XFILL_0__1755_ vdd gnd FILL
XFILL_0__1824_ vdd gnd FILL
XFILL_1__1100_ vdd gnd FILL
XFILL_1__1031_ vdd gnd FILL
X_1817_ _1871_/B _1817_/Y vdd gnd INVX1
X_1748_ _1748_/A _1748_/B _1748_/C _1756_/A vdd gnd OAI21X1
X_1679_ _1679_/D _1679_/CLK _964_/B vdd gnd DFFPOSX1
XFILL_1__1795_ vdd gnd FILL
XFILL_1__1864_ vdd gnd FILL
XFILL_1__1229_ vdd gnd FILL
XFILL_0__1540_ vdd gnd FILL
XFILL_0__1471_ vdd gnd FILL
X_1602_ LoadCmd_i _1602_/B _1602_/C _1654_/D vdd gnd OAI21X1
X_1464_ _1488_/B _1488_/A _1465_/C vdd gnd NAND2X1
X_1395_ _1444_/C _1442_/B _1442_/A _1396_/A vdd gnd OAI21X1
X_1533_ _1888_/A _1533_/B _1592_/C _1534_/B vdd gnd OAI21X1
XFILL_1__1580_ vdd gnd FILL
XFILL_0__1738_ vdd gnd FILL
XFILL_0__1807_ vdd gnd FILL
XFILL_1__1014_ vdd gnd FILL
XFILL86550x32550 vdd gnd FILL
XFILL_1__1778_ vdd gnd FILL
XFILL_1__1847_ vdd gnd FILL
X_1180_ _1180_/A _1181_/B vdd gnd INVX1
XFILL_0__1523_ vdd gnd FILL
XFILL_0__1454_ vdd gnd FILL
XFILL_0__1385_ vdd gnd FILL
X_1516_ _1583_/B _1522_/A vdd gnd INVX1
X_1447_ _1457_/A _1454_/B vdd gnd INVX1
XFILL_1__1632_ vdd gnd FILL
X_1378_ _1378_/A _1378_/B _1378_/C _1382_/A vdd gnd AOI21X1
XFILL_1__1701_ vdd gnd FILL
XFILL_1__1563_ vdd gnd FILL
XFILL_1__1494_ vdd gnd FILL
X_960_ _967_/A _967_/B _973_/C vdd gnd OR2X2
XFILL_2__1741_ vdd gnd FILL
XFILL_0__1170_ vdd gnd FILL
XFILL_2__1037_ vdd gnd FILL
XFILL_1__972_ vdd gnd FILL
X_1301_ _1302_/B _1302_/A _1303_/A vdd gnd NOR2X1
X_1232_ _1333_/B _1333_/A _1329_/C vdd gnd NAND2X1
XFILL_0__1506_ vdd gnd FILL
X_1163_ _1163_/A _1530_/B _1163_/C _1567_/A vdd gnd NAND3X1
XFILL_0__1437_ vdd gnd FILL
X_1094_ _1114_/A _1114_/B _1114_/C _1195_/B vdd gnd AOI21X1
XFILL_0__1368_ vdd gnd FILL
XFILL_0__1299_ vdd gnd FILL
XFILL_1__1615_ vdd gnd FILL
XFILL_1__1546_ vdd gnd FILL
XFILL_0__990_ vdd gnd FILL
XFILL_1__1477_ vdd gnd FILL
X_943_ _971_/C _957_/C vdd gnd INVX1
XFILL_0__1153_ vdd gnd FILL
XFILL_0__1222_ vdd gnd FILL
X_1781_ _1781_/A _1782_/C vdd gnd INVX1
X_1850_ _1850_/A _1850_/B _1851_/B vdd gnd NOR2X1
XFILL_0__1084_ vdd gnd FILL
XFILL_1__1400_ vdd gnd FILL
XFILL_1__955_ vdd gnd FILL
X_1146_ _952_/A _958_/B _979_/C _1147_/A vdd gnd NAND3X1
X_1215_ _1294_/A _1297_/A vdd gnd INVX1
X_1077_ _979_/B _1645_/B vdd gnd INVX1
XFILL_1__1331_ vdd gnd FILL
XFILL_1__1193_ vdd gnd FILL
XFILL_1__1262_ vdd gnd FILL
XFILL_1__1529_ vdd gnd FILL
XFILL_0__973_ vdd gnd FILL
XFILL_0__1840_ vdd gnd FILL
X_926_ _980_/B _926_/B _953_/C vdd gnd NAND2X1
XFILL_2__1638_ vdd gnd FILL
X_1000_ _1062_/A _958_/B _962_/B _1007_/A vdd gnd NAND3X1
XFILL_0__1771_ vdd gnd FILL
XFILL_0__1136_ vdd gnd FILL
X_1833_ _1871_/A _1833_/Y vdd gnd INVX1
XFILL_0__1067_ vdd gnd FILL
X_1764_ _964_/C _1766_/B _1765_/C vdd gnd NAND2X1
XFILL_0__1205_ vdd gnd FILL
XFILL_1__1880_ vdd gnd FILL
X_1695_ _961_/A _1695_/B _1839_/D _1695_/D _1702_/A vdd gnd AOI22X1
XFILL_1__938_ vdd gnd FILL
X_1129_ _937_/A _1143_/A vdd gnd INVX1
XFILL_1__1314_ vdd gnd FILL
XFILL_1__1176_ vdd gnd FILL
XFILL_1__1245_ vdd gnd FILL
XFILL_2__1285_ vdd gnd FILL
XFILL_0__956_ vdd gnd FILL
XFILL_1_CLKBUF1_insert4 vdd gnd FILL
X_1480_ _1480_/A _1480_/B _1482_/B vdd gnd NAND2X1
XFILL_0__1823_ vdd gnd FILL
XFILL_0__1754_ vdd gnd FILL
XFILL_0__1685_ vdd gnd FILL
XFILL_1__1030_ vdd gnd FILL
X_1678_ _1678_/D _1681_/CLK _958_/B vdd gnd DFFPOSX1
X_1816_ _1866_/A _1816_/B _1871_/B vdd gnd NAND2X1
XFILL_0__1119_ vdd gnd FILL
X_1747_ _980_/C _1747_/B _1863_/B _1748_/A vdd gnd OAI21X1
XFILL_1__1794_ vdd gnd FILL
XFILL_1__1863_ vdd gnd FILL
XFILL_1__1159_ vdd gnd FILL
XFILL_1__1228_ vdd gnd FILL
XFILL_0__1470_ vdd gnd FILL
XFILL_2__1337_ vdd gnd FILL
X_1601_ LoadCmd_i ABCmd_i[1] _1602_/C vdd gnd NAND2X1
XFILL_0__939_ vdd gnd FILL
X_1532_ Flag_i _1852_/B _1534_/A vdd gnd NOR2X1
X_1463_ _1463_/A _1510_/A _1463_/C _1465_/B vdd gnd NAND3X1
X_1394_ _1394_/A _1394_/B _1442_/B vdd gnd AND2X2
XFILL_0__1806_ vdd gnd FILL
XFILL_0__1599_ vdd gnd FILL
XFILL_0__1737_ vdd gnd FILL
XFILL_1__1013_ vdd gnd FILL
XFILL_1__1846_ vdd gnd FILL
XFILL_1__1777_ vdd gnd FILL
XFILL_2__1122_ vdd gnd FILL
XFILL_0__1453_ vdd gnd FILL
XFILL_0__1522_ vdd gnd FILL
XFILL_0__1384_ vdd gnd FILL
X_1515_ _1575_/A _1573_/A _1583_/B vdd gnd NAND2X1
XFILL_1__1700_ vdd gnd FILL
XFILL_1__1631_ vdd gnd FILL
X_1446_ _1448_/C _1490_/A _1491_/C _1457_/A vdd gnd NAND3X1
X_1377_ _1378_/C _1377_/B _1377_/C _1437_/C vdd gnd OAI21X1
XFILL_1__1562_ vdd gnd FILL
XFILL_2__953_ vdd gnd FILL
XFILL_1__1493_ vdd gnd FILL
XFILL_1__1829_ vdd gnd FILL
XFILL85950x10950 vdd gnd FILL
X_1162_ _997_/B _1185_/B _997_/A _1163_/C vdd gnd OAI21X1
XFILL_1__971_ vdd gnd FILL
X_1300_ _1826_/B _1370_/B _1302_/B vdd gnd NAND2X1
X_1231_ _1237_/B _1237_/A _1336_/A vdd gnd AND2X2
XFILL_0__1436_ vdd gnd FILL
XFILL_0__1505_ vdd gnd FILL
X_1093_ _1209_/C _1236_/B _1236_/A _1114_/B vdd gnd OAI21X1
XBUFX2_insert5 _1660_/Q _975_/A vdd gnd BUFX2
XFILL_0__1298_ vdd gnd FILL
XFILL_0__1367_ vdd gnd FILL
X_1429_ _1429_/A _1429_/B _1429_/C _1432_/C vdd gnd OAI21X1
XFILL_1__1614_ vdd gnd FILL
XFILL_1__1545_ vdd gnd FILL
XFILL_1__1476_ vdd gnd FILL
XFILL_2__1585_ vdd gnd FILL
X_942_ _946_/C _942_/B _971_/C vdd gnd NOR2X1
XFILL_0__1221_ vdd gnd FILL
XFILL_0__1152_ vdd gnd FILL
X_1780_ _1780_/A _1780_/B _1782_/A vdd gnd NAND2X1
XFILL_0__1083_ vdd gnd FILL
XFILL_1__954_ vdd gnd FILL
X_1145_ _1150_/C _1148_/A vdd gnd INVX1
XFILL_1__1330_ vdd gnd FILL
X_1214_ _1297_/C _1294_/B _1294_/A _1237_/A vdd gnd OAI21X1
XFILL_0__1419_ vdd gnd FILL
XFILL_1__1192_ vdd gnd FILL
X_1076_ _975_/A _958_/C _979_/B _1218_/C vdd gnd NAND3X1
XFILL_1__1261_ vdd gnd FILL
XFILL_1__1459_ vdd gnd FILL
XFILL_2__1370_ vdd gnd FILL
XFILL_1__1528_ vdd gnd FILL
XFILL_0__972_ vdd gnd FILL
X_925_ _925_/A _982_/A _926_/B vdd gnd NOR2X1
XFILL_0__1770_ vdd gnd FILL
X_1832_ _1832_/A _1848_/C _1871_/A vdd gnd NAND2X1
XFILL_0__1204_ vdd gnd FILL
XFILL_0__1135_ vdd gnd FILL
XFILL_0__1066_ vdd gnd FILL
X_1763_ _1837_/A _980_/B _1766_/B vdd gnd AND2X2
X_1694_ _975_/B _1729_/A _1695_/B vdd gnd NAND2X1
XFILL_1__937_ vdd gnd FILL
X_1128_ _927_/B _953_/C _1185_/C vdd gnd NOR2X1
XFILL_1__1313_ vdd gnd FILL
X_1059_ _975_/A _961_/A _1881_/B _1067_/C vdd gnd NAND3X1
XFILL_1__1244_ vdd gnd FILL
XFILL_1__1175_ vdd gnd FILL
XFILL_2__1422_ vdd gnd FILL
XFILL_0__955_ vdd gnd FILL
XFILL_0__1753_ vdd gnd FILL
XFILL_0__1822_ vdd gnd FILL
X_1815_ _1818_/A _1818_/B _1816_/B vdd gnd NAND2X1
X_1677_ _1677_/D _1684_/CLK _961_/A vdd gnd DFFPOSX1
XFILL_1__1862_ vdd gnd FILL
XFILL_0__1049_ vdd gnd FILL
XFILL_0__1118_ vdd gnd FILL
X_1746_ _1839_/A _964_/B _1746_/C _1839_/D _1748_/B vdd gnd AOI22X1
XFILL_1__1793_ vdd gnd FILL
XFILL_1_BUFX2_insert5 vdd gnd FILL
XFILL_1__1158_ vdd gnd FILL
XFILL_1__1089_ vdd gnd FILL
XFILL_1__1227_ vdd gnd FILL
XFILL_0__938_ vdd gnd FILL
X_1462_ _1462_/A _1462_/B _1462_/C _1463_/C vdd gnd OAI21X1
X_1531_ MulL_i _1531_/B _1539_/A _1534_/C vdd gnd NAND3X1
X_1600_ _1729_/A _1602_/B vdd gnd INVX1
X_1393_ _1394_/A _1394_/B _1444_/C vdd gnd NOR2X1
XFILL_0__1736_ vdd gnd FILL
XFILL_0__1805_ vdd gnd FILL
XFILL_0__1598_ vdd gnd FILL
XFILL_1__1012_ vdd gnd FILL
XFILL86250x39750 vdd gnd FILL
XFILL_1__1845_ vdd gnd FILL
X_1729_ _1729_/A _1729_/B _1744_/A _1731_/B vdd gnd MUX2X1
XFILL86250x82950 vdd gnd FILL
XFILL_1__1776_ vdd gnd FILL
XFILL_2__1885_ vdd gnd FILL
XFILL_0__1383_ vdd gnd FILL
XFILL_0__1452_ vdd gnd FILL
XFILL_0__1521_ vdd gnd FILL
X_1445_ _1631_/B _1548_/D _1445_/C _1490_/A vdd gnd OAI21X1
X_1514_ _1514_/A _1514_/B _1514_/C _1575_/A vdd gnd NAND3X1
XFILL_1__1630_ vdd gnd FILL
XFILL_1__1492_ vdd gnd FILL
X_1376_ _1382_/B _1377_/C vdd gnd INVX1
XFILL_1__1561_ vdd gnd FILL
XFILL86850x18150 vdd gnd FILL
XFILL_0__1719_ vdd gnd FILL
XFILL_1__1828_ vdd gnd FILL
XFILL_1__1759_ vdd gnd FILL
XFILL_1__970_ vdd gnd FILL
X_1161_ _1161_/A _1161_/B _1161_/C _1185_/B vdd gnd AOI21X1
XBUFX2_insert6 _1660_/Q _980_/A vdd gnd BUFX2
X_1092_ _1092_/A _1092_/B _1236_/A vdd gnd NAND2X1
X_1230_ _1238_/B _1329_/A _1238_/A _1340_/A vdd gnd NAND3X1
XFILL_0__1435_ vdd gnd FILL
XFILL_0__1504_ vdd gnd FILL
XFILL_0__1366_ vdd gnd FILL
XFILL_0__1297_ vdd gnd FILL
XFILL_1__1613_ vdd gnd FILL
XFILL_1_BUFX2_insert10 vdd gnd FILL
X_1428_ _1592_/C _1428_/B _1429_/C vdd gnd NOR2X1
XFILL_1__1544_ vdd gnd FILL
XFILL_1__1475_ vdd gnd FILL
X_1359_ _1474_/A _1521_/B _1523_/A _1361_/B vdd gnd OAI21X1
X_941_ _980_/A _958_/B _964_/C _942_/B vdd gnd NAND3X1
XFILL_2__1722_ vdd gnd FILL
XFILL_0__1220_ vdd gnd FILL
XFILL_0__1151_ vdd gnd FILL
XFILL_0__1082_ vdd gnd FILL
XFILL_1__953_ vdd gnd FILL
X_1213_ _1218_/C _1216_/B _1294_/B vdd gnd AND2X2
X_1144_ _952_/A _961_/A _980_/C _1150_/C vdd gnd NAND3X1
X_1075_ _1084_/A _1201_/D vdd gnd INVX1
XFILL_1__1260_ vdd gnd FILL
XFILL_0__1418_ vdd gnd FILL
XFILL_0__1349_ vdd gnd FILL
XFILL_1__1191_ vdd gnd FILL
XFILL_1__1458_ vdd gnd FILL
XFILL_1__1389_ vdd gnd FILL
XFILL_0__971_ vdd gnd FILL
XFILL_1__1527_ vdd gnd FILL
X_924_ _979_/C _982_/A vdd gnd INVX2
XFILL_0__1134_ vdd gnd FILL
X_1831_ _1866_/B _1861_/B _1866_/A _1832_/A vdd gnd NAND3X1
XFILL_0__1203_ vdd gnd FILL
XFILL_0__1065_ vdd gnd FILL
X_1693_ _961_/A _1837_/A _1695_/D vdd gnd NAND2X1
X_1762_ _1836_/A _958_/C _1767_/C vdd gnd NAND2X1
XFILL_1__936_ vdd gnd FILL
XFILL_1__1312_ vdd gnd FILL
X_1058_ _975_/A _958_/B _1823_/A _1065_/A vdd gnd NAND3X1
XFILL_1__1243_ vdd gnd FILL
X_1127_ _1127_/A _1127_/B _1127_/C _1591_/A vdd gnd AOI21X1
XFILL_1__1174_ vdd gnd FILL
XFILL_0__954_ vdd gnd FILL
XFILL_0__1752_ vdd gnd FILL
XFILL_0__1821_ vdd gnd FILL
X_1814_ _1814_/A _1814_/B _1814_/C _1818_/B vdd gnd AOI21X1
XFILL_0__1117_ vdd gnd FILL
X_1745_ _980_/C _1747_/B _1746_/C vdd gnd NAND2X1
X_1676_ _1676_/D _1683_/CLK _1881_/B vdd gnd DFFPOSX1
XFILL_0__1048_ vdd gnd FILL
XFILL_1__1861_ vdd gnd FILL
XFILL_1__1792_ vdd gnd FILL
XFILL_1_BUFX2_insert6 vdd gnd FILL
XFILL_1__1226_ vdd gnd FILL
XFILL_1__1157_ vdd gnd FILL
XFILL_1__1088_ vdd gnd FILL
XFILL_0__937_ vdd gnd FILL
X_1461_ _1461_/A _1461_/B _1461_/C _1470_/A vdd gnd NAND3X1
X_1392_ _1444_/A _1444_/B _1442_/C _1396_/B vdd gnd NAND3X1
X_1530_ _1530_/A _1530_/B _1530_/C _1531_/B vdd gnd OAI21X1
XFILL_0__1735_ vdd gnd FILL
XFILL_0__1804_ vdd gnd FILL
XFILL_0__1597_ vdd gnd FILL
XFILL_1__1011_ vdd gnd FILL
X_1728_ _1752_/A _1842_/C _1733_/B _1734_/B vdd gnd OAI21X1
X_1659_ _1659_/D _1684_/CLK _1858_/A vdd gnd DFFPOSX1
XFILL_1__1844_ vdd gnd FILL
XFILL_1__1775_ vdd gnd FILL
XFILL_1__1209_ vdd gnd FILL
XFILL_0__1520_ vdd gnd FILL
XFILL_0__1382_ vdd gnd FILL
XFILL_2__1318_ vdd gnd FILL
XFILL_0__1451_ vdd gnd FILL
X_1513_ _1513_/A _1513_/B _1573_/A vdd gnd NAND2X1
X_1444_ _1444_/A _1444_/B _1444_/C _1445_/C vdd gnd AOI21X1
X_1375_ _1826_/B _1440_/B _1382_/B vdd gnd NAND2X1
XFILL_1__1491_ vdd gnd FILL
XFILL_0__1649_ vdd gnd FILL
XFILL_1__1560_ vdd gnd FILL
XFILL_0__1718_ vdd gnd FILL
XFILL_1__1758_ vdd gnd FILL
XFILL_1__1827_ vdd gnd FILL
XFILL_1__1689_ vdd gnd FILL
X_1160_ _1187_/A _1530_/B vdd gnd INVX1
XBUFX2_insert7 _1660_/Q _923_/A vdd gnd BUFX2
XFILL_0__1503_ vdd gnd FILL
X_1091_ _935_/A _1501_/A _1091_/C _1092_/B vdd gnd OAI21X1
XFILL_0__1365_ vdd gnd FILL
XFILL_0__1296_ vdd gnd FILL
XFILL_0__1434_ vdd gnd FILL
XFILL_1__1612_ vdd gnd FILL
XFILL_1_BUFX2_insert11 vdd gnd FILL
X_1427_ _1427_/A _1427_/B _1429_/B vdd gnd AND2X2
X_1358_ _1358_/A _1523_/A _1523_/B _1362_/A vdd gnd AOI21X1
XFILL_1__1543_ vdd gnd FILL
XFILL_1__1474_ vdd gnd FILL
X_1289_ _1289_/A _1344_/B _1289_/C _1290_/C vdd gnd NOR3X1
X_940_ _952_/A _961_/A _958_/C _946_/C vdd gnd NAND3X1
XFILL_0__1150_ vdd gnd FILL
XFILL_0__1081_ vdd gnd FILL
XFILL_2__1017_ vdd gnd FILL
XFILL_1__952_ vdd gnd FILL
X_1212_ _1218_/C _1216_/B _1297_/C vdd gnd NOR2X1
XFILL_0__1417_ vdd gnd FILL
X_1143_ _1143_/A _936_/A _937_/C _1156_/A vdd gnd NAND3X1
X_1074_ _975_/A _977_/A _980_/C _1084_/A vdd gnd NAND3X1
XFILL_0__1348_ vdd gnd FILL
XFILL_1__1190_ vdd gnd FILL
XFILL_0__1279_ vdd gnd FILL
XFILL_1__1526_ vdd gnd FILL
XFILL_1__1457_ vdd gnd FILL
XFILL_1__1388_ vdd gnd FILL
XFILL_0__970_ vdd gnd FILL
X_923_ _923_/A _925_/A vdd gnd INVX1
XFILL_2__1566_ vdd gnd FILL
XFILL_0__1133_ vdd gnd FILL
X_1830_ _1874_/B _1874_/A _1848_/C vdd gnd NAND2X1
X_1761_ _1794_/B _1794_/A _1795_/B vdd gnd AND2X2
XFILL_0__1202_ vdd gnd FILL
XFILL_0__1064_ vdd gnd FILL
X_1692_ _1744_/A _1837_/A vdd gnd INVX2
XFILL_1__935_ vdd gnd FILL
XFILL_0__1897_ vdd gnd FILL
X_1126_ _1127_/C _1127_/B _1127_/A _1262_/A vdd gnd NAND3X1
XFILL_1__1311_ vdd gnd FILL
X_1057_ _1057_/A _1057_/B _1057_/C _1088_/C vdd gnd AOI21X1
XFILL_1__1242_ vdd gnd FILL
XFILL_1__1173_ vdd gnd FILL
XFILL_1__1509_ vdd gnd FILL
XFILL85950x18150 vdd gnd FILL
XFILL_0__953_ vdd gnd FILL
XFILL_0__1820_ vdd gnd FILL
XFILL_2__1618_ vdd gnd FILL
XFILL_0__1751_ vdd gnd FILL
X_1813_ _1814_/C _1813_/B _1813_/C _1866_/A vdd gnd OAI21X1
XFILL_0__1047_ vdd gnd FILL
XFILL_0__1116_ vdd gnd FILL
X_1744_ _1744_/A _1744_/B _1747_/B vdd gnd NOR2X1
X_1675_ _1675_/D _1683_/CLK _1823_/A vdd gnd DFFPOSX1
XFILL_1__1860_ vdd gnd FILL
XFILL_1__1791_ vdd gnd FILL
XFILL_1_BUFX2_insert7 vdd gnd FILL
XFILL86850x46950 vdd gnd FILL
X_1109_ _982_/A _1548_/D _1109_/C _1110_/B vdd gnd OAI21X1
XFILL_1__1156_ vdd gnd FILL
XFILL_1__1225_ vdd gnd FILL
XFILL_1__1087_ vdd gnd FILL
XFILL_2__1265_ vdd gnd FILL
XFILL_0__936_ vdd gnd FILL
X_1460_ _1460_/A _1460_/B _1488_/B _1461_/B vdd gnd OAI21X1
X_1391_ _1633_/B _982_/B _1394_/B _1444_/B vdd gnd OAI21X1
XFILL_0__1803_ vdd gnd FILL
XFILL_0__1734_ vdd gnd FILL
XFILL_0__1596_ vdd gnd FILL
XFILL_1__1010_ vdd gnd FILL
X_1727_ _1727_/A _1733_/B vdd gnd INVX1
X_1658_ _1658_/D _1684_/CLK _1836_/A vdd gnd DFFPOSX1
XFILL86850x21750 vdd gnd FILL
X_1589_ _1589_/A _1589_/B _1589_/C _1590_/B vdd gnd OAI21X1
XFILL_1__1774_ vdd gnd FILL
XFILL_1__1843_ vdd gnd FILL
XFILL_1__1139_ vdd gnd FILL
XFILL_2__1050_ vdd gnd FILL
XFILL_1__1208_ vdd gnd FILL
XFILL_0__1450_ vdd gnd FILL
XFILL_0__1381_ vdd gnd FILL
X_1512_ _1514_/B _1514_/C _1513_/B vdd gnd NAND2X1
X_1443_ _962_/B _1577_/B _1443_/C _1491_/C vdd gnd NAND3X1
X_1374_ _925_/A _1629_/B _1440_/B vdd gnd NOR2X1
XFILL_0__1648_ vdd gnd FILL
XFILL_1__1490_ vdd gnd FILL
XFILL_0__1579_ vdd gnd FILL
XFILL_0__1717_ vdd gnd FILL
XFILL86550x68550 vdd gnd FILL
XFILL_1__1757_ vdd gnd FILL
XFILL_1__1688_ vdd gnd FILL
XFILL_1__1826_ vdd gnd FILL
XFILL_2__1102_ vdd gnd FILL
XFILL_2__1866_ vdd gnd FILL
XFILL_0__1502_ vdd gnd FILL
X_1090_ _952_/A _977_/A _1501_/A vdd gnd NAND2X1
XBUFX2_insert8 _1660_/Q _962_/A vdd gnd BUFX2
XFILL_0__1433_ vdd gnd FILL
XFILL_0__1295_ vdd gnd FILL
XFILL_0__1364_ vdd gnd FILL
X_1426_ _1472_/C _1426_/B _1434_/B vdd gnd NAND2X1
XFILL_1__1611_ vdd gnd FILL
X_1288_ _1354_/A _1420_/A vdd gnd INVX1
X_1357_ _1523_/C _1520_/D _1523_/B vdd gnd NAND2X1
XFILL_1_BUFX2_insert12 vdd gnd FILL
XFILL_1__1542_ vdd gnd FILL
XFILL_1__1473_ vdd gnd FILL
XFILL86550x43350 vdd gnd FILL
XFILL_2__933_ vdd gnd FILL
XFILL_2__1651_ vdd gnd FILL
XFILL_1__1809_ vdd gnd FILL
XFILL_0__1080_ vdd gnd FILL
X_1142_ _956_/C _1142_/B _1142_/C _1183_/B vdd gnd NAND3X1
XFILL_1__951_ vdd gnd FILL
X_999_ _999_/A _999_/B _999_/C _999_/Y vdd gnd AOI21X1
X_1211_ _975_/A _962_/B _980_/B _1216_/B vdd gnd NAND3X1
XFILL_0__1416_ vdd gnd FILL
X_1073_ _1087_/B _1087_/C _1087_/A _1236_/C vdd gnd NAND3X1
XFILL_0__1347_ vdd gnd FILL
XFILL_0__1278_ vdd gnd FILL
X_1409_ _1409_/A _1410_/B vdd gnd INVX1
XFILL_1__1525_ vdd gnd FILL
XFILL_1__1456_ vdd gnd FILL
XFILL_1__1387_ vdd gnd FILL
X_922_ _975_/B _922_/B _927_/B vdd gnd NAND2X1
XFILL_0__1201_ vdd gnd FILL
XFILL_2_CLKBUF1_insert1 vdd gnd FILL
XFILL_0__1132_ vdd gnd FILL
X_1760_ _1780_/A _1773_/A vdd gnd INVX1
XFILL_0__1063_ vdd gnd FILL
X_1691_ _1744_/A _1839_/A _1839_/D vdd gnd NAND2X1
XCLKBUF1_insert0 clk _1668_/CLK vdd gnd CLKBUF1
XFILL_1__934_ vdd gnd FILL
XFILL_1__1310_ vdd gnd FILL
XFILL_0__1896_ vdd gnd FILL
X_1125_ _1256_/B _1192_/C _1256_/A _1127_/A vdd gnd OAI21X1
XFILL_1__1172_ vdd gnd FILL
X_1056_ _1056_/A _1056_/B _1056_/C _1114_/C vdd gnd OAI21X1
XFILL_1__1241_ vdd gnd FILL
X_1889_ _1889_/A _1889_/B _1889_/Y vdd gnd AND2X2
XFILL_1__1508_ vdd gnd FILL
XFILL_1__1439_ vdd gnd FILL
XFILL_2__1350_ vdd gnd FILL
XFILL_0__952_ vdd gnd FILL
XFILL_0__1750_ vdd gnd FILL
X_1674_ _1674_/D _1683_/CLK _962_/B vdd gnd DFFPOSX1
X_1812_ _1818_/A _1813_/C vdd gnd INVX1
XFILL_0__1046_ vdd gnd FILL
XFILL_0__1115_ vdd gnd FILL
X_1743_ _964_/B _1744_/B vdd gnd INVX1
XFILL_1_BUFX2_insert8 vdd gnd FILL
XFILL_1__1790_ vdd gnd FILL
X_1039_ _991_/C _991_/A _992_/A _1044_/C vdd gnd AOI21X1
XFILL_0__1879_ vdd gnd FILL
X_1108_ _1193_/A _1193_/B _1194_/C vdd gnd NAND2X1
XFILL_1__1155_ vdd gnd FILL
XFILL_1__1224_ vdd gnd FILL
XFILL_1__1086_ vdd gnd FILL
XFILL_2__1402_ vdd gnd FILL
XFILL_0__935_ vdd gnd FILL
X_1390_ _1823_/A _1633_/B vdd gnd INVX1
XFILL_0__1733_ vdd gnd FILL
XFILL_0__1802_ vdd gnd FILL
XFILL_0__1595_ vdd gnd FILL
X_1657_ _1657_/D _1679_/CLK _1836_/B vdd gnd DFFPOSX1
X_1726_ _1726_/A _1726_/B _1757_/C vdd gnd NAND2X1
XFILL_0__1029_ vdd gnd FILL
XFILL_1__1842_ vdd gnd FILL
X_1588_ _1588_/A _1588_/B _1667_/D vdd gnd NAND2X1
XFILL_1__1773_ vdd gnd FILL
XFILL_1__1138_ vdd gnd FILL
XFILL_1__1069_ vdd gnd FILL
XFILL_1__1207_ vdd gnd FILL
XFILL_0__1380_ vdd gnd FILL
X_1511_ _1543_/A _1543_/B _1511_/C _1514_/C vdd gnd NAND3X1
X_1442_ _1442_/A _1442_/B _1442_/C _1443_/C vdd gnd OAI21X1
X_1373_ _958_/C _1629_/B vdd gnd INVX1
XFILL_0__1716_ vdd gnd FILL
XFILL_0__1647_ vdd gnd FILL
XFILL_0__1578_ vdd gnd FILL
X_1709_ _1836_/A _1709_/B _1709_/C _1710_/A vdd gnd OAI21X1
XFILL_1__1825_ vdd gnd FILL
XFILL_1__1756_ vdd gnd FILL
XFILL_1__1687_ vdd gnd FILL
XFILL_0__1501_ vdd gnd FILL
XFILL_0__1363_ vdd gnd FILL
XFILL_0__1432_ vdd gnd FILL
XBUFX2_insert9 _1660_/Q _1062_/A vdd gnd BUFX2
XFILL_0__1294_ vdd gnd FILL
X_1425_ _1425_/A _1425_/B _1426_/B vdd gnd OR2X2
XFILL_1_BUFX2_insert13 vdd gnd FILL
XFILL_1__1472_ vdd gnd FILL
XFILL_1__1610_ vdd gnd FILL
X_1356_ _1418_/B _1356_/B _1356_/C _1523_/C vdd gnd NAND3X1
XFILL_1__1541_ vdd gnd FILL
X_1287_ _1287_/A _1287_/B _1287_/C _1354_/A vdd gnd OAI21X1
XFILL_1__1808_ vdd gnd FILL
XFILL85950x46950 vdd gnd FILL
XFILL_1__1739_ vdd gnd FILL
XFILL_1__950_ vdd gnd FILL
X_1141_ _1185_/C _997_/C _1186_/C _1163_/A vdd gnd NAND3X1
X_998_ _998_/A _998_/B _998_/C _998_/Y vdd gnd OAI21X1
X_1210_ _962_/A _964_/C _977_/A _1294_/A vdd gnd NAND3X1
X_1072_ _1221_/C _1228_/A _1228_/B _1087_/B vdd gnd OAI21X1
XFILL_0__1415_ vdd gnd FILL
XFILL_0__1346_ vdd gnd FILL
XFILL_0__1277_ vdd gnd FILL
X_1408_ _1408_/A _1409_/A _1408_/C _1411_/A vdd gnd NAND3X1
XFILL_1__1455_ vdd gnd FILL
XFILL_1__1524_ vdd gnd FILL
X_1339_ _1419_/A _1419_/B _1349_/C _1355_/C vdd gnd NAND3X1
XFILL_1__1386_ vdd gnd FILL
X_921_ _923_/A _979_/B _922_/B vdd gnd AND2X2
XFILL_2__1702_ vdd gnd FILL
XFILL_0__1200_ vdd gnd FILL
XFILL_0__1131_ vdd gnd FILL
XFILL_0__1062_ vdd gnd FILL
XCLKBUF1_insert1 clk _1679_/CLK vdd gnd CLKBUF1
X_1690_ _1729_/A _1839_/A vdd gnd INVX2
XFILL_0__1895_ vdd gnd FILL
XFILL_1__933_ vdd gnd FILL
X_1055_ _1055_/A _1055_/B _1055_/C _1124_/C vdd gnd AOI21X1
X_1124_ _1124_/A _1124_/B _1124_/C _1192_/C vdd gnd AOI21X1
XFILL_1__1171_ vdd gnd FILL
XFILL_0__1329_ vdd gnd FILL
XFILL_1__1240_ vdd gnd FILL
X_1888_ _1888_/A _1888_/B _1889_/B vdd gnd NAND2X1
XFILL_1__1507_ vdd gnd FILL
XFILL_1__1438_ vdd gnd FILL
XFILL_0__951_ vdd gnd FILL
XFILL_1__1369_ vdd gnd FILL
X_1811_ _1811_/A _1811_/B _1866_/B _1818_/A vdd gnd OAI21X1
XFILL_0__1114_ vdd gnd FILL
X_1673_ _1673_/D _1684_/CLK _958_/C vdd gnd DFFPOSX1
X_1742_ _1836_/A _964_/C _1748_/C vdd gnd NAND2X1
XFILL_0__1045_ vdd gnd FILL
XFILL_0__1878_ vdd gnd FILL
XFILL_1_BUFX2_insert9 vdd gnd FILL
X_1107_ _1107_/A _1107_/B _1107_/C _1115_/A vdd gnd NAND3X1
X_1038_ _1826_/B _977_/B _1040_/B vdd gnd NAND2X1
XFILL_1__1223_ vdd gnd FILL
XFILL_1__1154_ vdd gnd FILL
XFILL_1__1085_ vdd gnd FILL
XFILL_0__934_ vdd gnd FILL
XFILL_0__1801_ vdd gnd FILL
XFILL_0__1732_ vdd gnd FILL
XFILL_0__1594_ vdd gnd FILL
X_1725_ _1725_/A _1725_/B _1740_/B _1726_/A vdd gnd MUX2X1
X_1656_ _1656_/D _1679_/CLK _1686_/A vdd gnd DFFPOSX1
XFILL_0__1028_ vdd gnd FILL
XFILL_1__1772_ vdd gnd FILL
XFILL_1__1841_ vdd gnd FILL
X_1587_ MulH_i _1587_/B _1595_/C _1588_/B vdd gnd NAND3X1
XFILL_1__1206_ vdd gnd FILL
XFILL_1__1137_ vdd gnd FILL
XFILL_1__1068_ vdd gnd FILL
XFILL_2__1246_ vdd gnd FILL
X_1441_ _1491_/A _1448_/C vdd gnd INVX1
X_1510_ _1510_/A _1510_/B _1543_/B vdd gnd NAND2X1
XFILL_0__1646_ vdd gnd FILL
X_1372_ _1372_/A _1372_/B _1378_/C vdd gnd NOR2X1
XFILL_0__1715_ vdd gnd FILL
XFILL_0__1577_ vdd gnd FILL
X_1708_ _1709_/C _1713_/A _1710_/B vdd gnd OR2X2
X_1639_ LoadB_i _946_/A _1639_/C _1678_/D vdd gnd OAI21X1
XFILL_1__1755_ vdd gnd FILL
XFILL_1__1824_ vdd gnd FILL
XFILL_1__1686_ vdd gnd FILL
XFILL_0__1500_ vdd gnd FILL
XFILL_0__1293_ vdd gnd FILL
XFILL_0__1431_ vdd gnd FILL
XFILL_0__1362_ vdd gnd FILL
X_1424_ _1425_/B _1425_/A _1472_/C vdd gnd NAND2X1
X_1355_ _1420_/A _1355_/B _1355_/C _1356_/B vdd gnd NAND3X1
XFILL_1_BUFX2_insert14 vdd gnd FILL
XFILL_0__1629_ vdd gnd FILL
XFILL_1__1471_ vdd gnd FILL
X_1286_ _1286_/A _1286_/B _1286_/C _1351_/C vdd gnd AOI21X1
XFILL_1__1540_ vdd gnd FILL
XFILL_1__1738_ vdd gnd FILL
XFILL_1__1807_ vdd gnd FILL
X_997_ _997_/A _997_/B _997_/C _997_/Y vdd gnd OAI21X1
X_1140_ _1161_/B _1161_/A _1161_/C _1186_/C vdd gnd NAND3X1
X_1071_ _1221_/A _1221_/B _1228_/C _1087_/A vdd gnd NAND3X1
XFILL_0__1414_ vdd gnd FILL
XFILL_0__1345_ vdd gnd FILL
XFILL_0__1276_ vdd gnd FILL
X_1407_ _1410_/C _1408_/C vdd gnd INVX1
X_1338_ _1369_/B _1369_/A _1405_/C _1419_/B vdd gnd NAND3X1
XFILL_1__1454_ vdd gnd FILL
XFILL_1__1385_ vdd gnd FILL
XFILL_1__1523_ vdd gnd FILL
X_1269_ _1474_/A _1521_/B _1270_/B vdd gnd NAND2X1
XFILL86250x25350 vdd gnd FILL
X_920_ MulH_i _920_/Y vdd gnd INVX2
XFILL_2__1494_ vdd gnd FILL
XFILL_0__1130_ vdd gnd FILL
XCLKBUF1_insert2 clk _1684_/CLK vdd gnd CLKBUF1
XFILL_0__1061_ vdd gnd FILL
XFILL_1__932_ vdd gnd FILL
XFILL_0__1894_ vdd gnd FILL
X_1123_ _1123_/A _1123_/B _1123_/C _1256_/B vdd gnd AOI21X1
X_1054_ _1256_/A _1192_/B vdd gnd INVX1
XFILL_1__1170_ vdd gnd FILL
XFILL_0__1328_ vdd gnd FILL
X_1887_ _1887_/A _1887_/B _1888_/B vdd gnd NAND2X1
XFILL_0__1259_ vdd gnd FILL
XFILL_1__1506_ vdd gnd FILL
XFILL_1__1437_ vdd gnd FILL
XFILL_1__1368_ vdd gnd FILL
XFILL_0__950_ vdd gnd FILL
XFILL_1__1299_ vdd gnd FILL
XFILL_2__1546_ vdd gnd FILL
X_1741_ _1741_/A _1741_/B _1757_/A _1794_/B vdd gnd OAI21X1
X_1810_ _1878_/A _1811_/B _1811_/A _1866_/B vdd gnd OAI21X1
XFILL_0__1113_ vdd gnd FILL
X_1672_ _1672_/D _1681_/CLK _964_/C vdd gnd DFFPOSX1
XFILL_0__1044_ vdd gnd FILL
XFILL_0__1877_ vdd gnd FILL
X_1106_ _1109_/C _1193_/A _1107_/B vdd gnd NAND2X1
XFILL_1__1153_ vdd gnd FILL
XFILL_1__1222_ vdd gnd FILL
X_1037_ _1048_/B _1048_/A _1048_/C _1055_/C vdd gnd AOI21X1
XFILL_1__1084_ vdd gnd FILL
XFILL_2__1331_ vdd gnd FILL
XFILL_2__1193_ vdd gnd FILL
XFILL_0__933_ vdd gnd FILL
XFILL_0__1731_ vdd gnd FILL
XFILL_0__1800_ vdd gnd FILL
XFILL_0__1593_ vdd gnd FILL
X_1724_ _1752_/A _1842_/C _1725_/B _1725_/A vdd gnd OAI21X1
XFILL_0__1027_ vdd gnd FILL
X_1586_ _1586_/A _1586_/B _1586_/C _1587_/B vdd gnd NAND3X1
XFILL_1__1771_ vdd gnd FILL
XFILL_1__1840_ vdd gnd FILL
X_1655_ _1655_/D _1679_/CLK _1655_/Q vdd gnd DFFPOSX1
XFILL_1__1136_ vdd gnd FILL
XFILL_1__1205_ vdd gnd FILL
XFILL_1__1067_ vdd gnd FILL
X_1440_ _1843_/B _1440_/B _1491_/A vdd gnd NAND2X1
X_1371_ _1437_/A _1380_/A vdd gnd INVX1
XFILL_0__1645_ vdd gnd FILL
XFILL_0__1714_ vdd gnd FILL
XFILL_0__1576_ vdd gnd FILL
X_1638_ ABCmd_i[1] LoadB_i _1639_/C vdd gnd NAND2X1
X_1707_ _1734_/A _1727_/A _1713_/C _1709_/C vdd gnd OAI21X1
X_1569_ _1569_/A _1569_/B MulL_i _1571_/A vdd gnd OAI21X1
XFILL_1__1754_ vdd gnd FILL
XFILL_1__1685_ vdd gnd FILL
XFILL_1__1823_ vdd gnd FILL
XFILL_2__1030_ vdd gnd FILL
XFILL_1__1119_ vdd gnd FILL
XFILL_2__1794_ vdd gnd FILL
XFILL_0__1430_ vdd gnd FILL
XFILL_0__1292_ vdd gnd FILL
XFILL_0__1361_ vdd gnd FILL
X_1423_ _1524_/B _1425_/B vdd gnd INVX1
X_1354_ _1354_/A _1420_/C _1354_/C _1418_/B vdd gnd NAND3X1
X_1285_ _1285_/A _1285_/B _1286_/C vdd gnd NOR2X1
XFILL_1__1470_ vdd gnd FILL
XFILL_0__1628_ vdd gnd FILL
XFILL_0__1559_ vdd gnd FILL
XFILL_1__1737_ vdd gnd FILL
XFILL_1__1806_ vdd gnd FILL
XFILL_1__1599_ vdd gnd FILL
X_996_ _996_/A _996_/B _996_/C _997_/B vdd gnd AOI21X1
XFILL_2__1846_ vdd gnd FILL
XFILL_0__1413_ vdd gnd FILL
X_1070_ _1070_/A _1070_/B _1070_/C _1087_/C vdd gnd OAI21X1
XFILL_0__1344_ vdd gnd FILL
XFILL_0__1275_ vdd gnd FILL
X_1406_ _1406_/A _1406_/B _1462_/C _1439_/B _1435_/A vdd gnd AOI22X1
XFILL_1__1522_ vdd gnd FILL
X_1337_ _1344_/C _1343_/A _1369_/B vdd gnd NAND2X1
X_1268_ _1523_/A _1268_/B _1474_/A vdd gnd NAND2X1
XFILL_1__1384_ vdd gnd FILL
XFILL_1__1453_ vdd gnd FILL
X_1199_ _1287_/A _1204_/A vdd gnd INVX1
XFILL_2__1631_ vdd gnd FILL
XFILL_0__1060_ vdd gnd FILL
XCLKBUF1_insert3 clk _1683_/CLK vdd gnd CLKBUF1
X_979_ _980_/A _979_/B _979_/C _981_/A vdd gnd NAND3X1
XFILL_1__931_ vdd gnd FILL
XFILL_0__1893_ vdd gnd FILL
X_1122_ _1192_/B _1256_/C _1192_/A _1127_/B vdd gnd NAND3X1
X_1053_ _1265_/A _1127_/C vdd gnd INVX1
XFILL_0__1327_ vdd gnd FILL
XFILL_0__1189_ vdd gnd FILL
X_1886_ _1887_/B _1887_/A _1886_/C _1889_/A vdd gnd NAND3X1
XFILL_0__1258_ vdd gnd FILL
XFILL_1__1505_ vdd gnd FILL
XFILL_1__1436_ vdd gnd FILL
XFILL_1__1298_ vdd gnd FILL
XFILL_1__1367_ vdd gnd FILL
X_1671_ _1671_/D _1679_/CLK _980_/C vdd gnd DFFPOSX1
X_1740_ _1740_/A _1740_/B _1741_/A vdd gnd NOR2X1
XFILL_0__1112_ vdd gnd FILL
XFILL_0__1043_ vdd gnd FILL
XFILL_0__1876_ vdd gnd FILL
X_1105_ _1105_/A _1193_/A vdd gnd INVX1
XFILL_1__1152_ vdd gnd FILL
XFILL_1__1221_ vdd gnd FILL
X_1036_ _1095_/B _1056_/C _1056_/B _1048_/A vdd gnd NAND3X1
X_1869_ _1872_/B _1872_/A _1870_/C vdd gnd AND2X2
XFILL_1__1083_ vdd gnd FILL
XFILL_1__1419_ vdd gnd FILL
XFILL_0__932_ vdd gnd FILL
XFILL_0__1730_ vdd gnd FILL
XFILL_0__1592_ vdd gnd FILL
X_1654_ _1654_/D _1684_/CLK _1729_/A vdd gnd DFFPOSX1
X_1723_ _1740_/A _1725_/B vdd gnd INVX1
XFILL_0__1026_ vdd gnd FILL
X_1585_ _1585_/A _1586_/A vdd gnd INVX1
XFILL_1__1770_ vdd gnd FILL
XFILL_0__1859_ vdd gnd FILL
X_1019_ _1023_/A _1080_/A _1101_/C vdd gnd NOR2X1
XFILL_1__1135_ vdd gnd FILL
XFILL_1__1066_ vdd gnd FILL
XFILL_1__1204_ vdd gnd FILL
X_1370_ _1843_/B _1370_/B _1437_/A vdd gnd NAND2X1
XFILL_0__1713_ vdd gnd FILL
XFILL_0__1575_ vdd gnd FILL
XFILL_0__1644_ vdd gnd FILL
X_1637_ LoadB_i _963_/A _1637_/C _1677_/D vdd gnd OAI21X1
XFILL_0__1009_ vdd gnd FILL
X_1706_ _1878_/A _1727_/A _1734_/A _1713_/C vdd gnd OAI21X1
XFILL_1__1822_ vdd gnd FILL
XFILL86850x57750 vdd gnd FILL
X_1499_ _1504_/A _1504_/C _1551_/B vdd gnd NAND2X1
X_1568_ _1568_/A _1568_/B _1568_/C _1571_/B vdd gnd AOI21X1
XFILL_1__1753_ vdd gnd FILL
XFILL_1__1049_ vdd gnd FILL
XFILL_1__1118_ vdd gnd FILL
XFILL_0__1291_ vdd gnd FILL
XFILL_0__1360_ vdd gnd FILL
X_1422_ _1519_/C _1517_/B _1524_/B vdd gnd NAND2X1
XFILL85950x7350 vdd gnd FILL
XFILL_2__1089_ vdd gnd FILL
X_1284_ _1352_/A _1352_/B _1285_/B vdd gnd NAND2X1
X_1353_ _1353_/A _1353_/B _1353_/C _1356_/C vdd gnd OAI21X1
XFILL_0__1489_ vdd gnd FILL
XFILL_0__1558_ vdd gnd FILL
XFILL_0__1627_ vdd gnd FILL
XFILL86850x32550 vdd gnd FILL
XFILL_1__1805_ vdd gnd FILL
XFILL_1__1598_ vdd gnd FILL
XFILL_1__1736_ vdd gnd FILL
X_995_ _996_/B _996_/A _996_/C _997_/C vdd gnd NAND3X1
XFILL_0__1412_ vdd gnd FILL
XFILL_0__1343_ vdd gnd FILL
XFILL_0__1274_ vdd gnd FILL
X_1405_ _1405_/A _1405_/B _1405_/C _1468_/C vdd gnd OAI21X1
XFILL_1__1452_ vdd gnd FILL
XFILL_1__1521_ vdd gnd FILL
X_1336_ _1336_/A _1336_/B _1344_/A _1343_/A vdd gnd AOI21X1
X_1267_ _1267_/A _1593_/B _1591_/B _1521_/B vdd gnd AOI21X1
X_1198_ _979_/C _1547_/B _1287_/A vdd gnd NAND2X1
XFILL_1__1383_ vdd gnd FILL
XFILL_1__1719_ vdd gnd FILL
XFILL_1__930_ vdd gnd FILL
XCLKBUF1_insert4 clk _1681_/CLK vdd gnd CLKBUF1
XFILL_0__1892_ vdd gnd FILL
X_978_ _992_/C _991_/C vdd gnd INVX1
X_1121_ _1123_/B _1123_/C _1123_/A _1256_/C vdd gnd NAND3X1
X_1052_ _997_/Y _1052_/B _1265_/A vdd gnd NAND2X1
XFILL_0__1326_ vdd gnd FILL
XFILL_0__1188_ vdd gnd FILL
X_1885_ _1885_/A _1885_/B _1885_/C _1887_/A vdd gnd NAND3X1
XFILL_0__1257_ vdd gnd FILL
XFILL_1__1435_ vdd gnd FILL
X_1319_ _1319_/A _1319_/B _1319_/C _1322_/A vdd gnd NAND3X1
XFILL86550x54150 vdd gnd FILL
XFILL_1__1504_ vdd gnd FILL
XFILL_1__1366_ vdd gnd FILL
XFILL_1__1297_ vdd gnd FILL
XFILL_0__1042_ vdd gnd FILL
X_1670_ _1670_/D _1681_/CLK _979_/C vdd gnd DFFPOSX1
XFILL_0__1111_ vdd gnd FILL
XFILL_0__1875_ vdd gnd FILL
X_1035_ _1095_/C _1056_/A _1095_/A _1048_/B vdd gnd OAI21X1
X_1104_ _979_/C _1577_/B _1105_/A vdd gnd NAND2X1
XFILL_0__1309_ vdd gnd FILL
XFILL_1__1151_ vdd gnd FILL
XFILL_1__1220_ vdd gnd FILL
XFILL_1__1082_ vdd gnd FILL
X_1868_ _1868_/A _1868_/B _1868_/C _1872_/B vdd gnd OAI21X1
X_1799_ _1814_/B _1814_/A _1800_/B vdd gnd NOR2X1
XFILL_0__931_ vdd gnd FILL
XFILL_1__1418_ vdd gnd FILL
XFILL_1__1349_ vdd gnd FILL
XFILL_2__1527_ vdd gnd FILL
XFILL_0__1591_ vdd gnd FILL
XFILL_2__1389_ vdd gnd FILL
X_1584_ _1584_/A _1584_/B _1584_/C _1586_/C vdd gnd NAND3X1
X_1653_ _1653_/D _1679_/CLK _1744_/A vdd gnd DFFPOSX1
X_1722_ _1752_/A _958_/B _1722_/C _1740_/A vdd gnd AOI21X1
XFILL_0__1025_ vdd gnd FILL
XFILL_0__1858_ vdd gnd FILL
XFILL_0__1789_ vdd gnd FILL
X_1018_ _1062_/A _980_/B _964_/C _1080_/A vdd gnd NAND3X1
XFILL_1__1203_ vdd gnd FILL
XFILL_1__1134_ vdd gnd FILL
XFILL_1__1065_ vdd gnd FILL
XFILL_2__1174_ vdd gnd FILL
XFILL_0__1712_ vdd gnd FILL
XFILL_0__1574_ vdd gnd FILL
XFILL_0__1643_ vdd gnd FILL
X_1705_ _1809_/A _1842_/C _1878_/A vdd gnd NOR2X1
X_1636_ ABCmd_i[0] LoadB_i _1637_/C vdd gnd NAND2X1
X_1567_ _1567_/A _1569_/B _1568_/A vdd gnd NAND2X1
XFILL_0__1008_ vdd gnd FILL
XFILL_1__1821_ vdd gnd FILL
X_1498_ _1652_/B _963_/B _1498_/C _1504_/A vdd gnd OAI21X1
XFILL_1__1752_ vdd gnd FILL
XFILL_1__1048_ vdd gnd FILL
XFILL_1__1117_ vdd gnd FILL
XFILL_0__1290_ vdd gnd FILL
XFILL_2__1226_ vdd gnd FILL
X_1421_ _1421_/A _1421_/B _1421_/C _1519_/C vdd gnd NAND3X1
XFILL_0__1626_ vdd gnd FILL
X_1352_ _1352_/A _1352_/B _1352_/C _1353_/B vdd gnd AOI21X1
X_1283_ _1283_/A _1283_/B _1362_/C vdd gnd NAND2X1
XFILL_0__1488_ vdd gnd FILL
XFILL_0__1557_ vdd gnd FILL
X_1619_ LoadCmd_i _925_/A _1619_/C _1660_/D vdd gnd OAI21X1
XFILL_1__1735_ vdd gnd FILL
XFILL_1__1804_ vdd gnd FILL
XFILL_1__1597_ vdd gnd FILL
XFILL_2__1011_ vdd gnd FILL
XFILL86850x3750 vdd gnd FILL
XFILL86550x7350 vdd gnd FILL
X_994_ _994_/A _998_/B _998_/A _996_/A vdd gnd OAI21X1
XFILL_0__1411_ vdd gnd FILL
XFILL_0__1342_ vdd gnd FILL
XFILL_0__1273_ vdd gnd FILL
X_1404_ _1468_/A _1468_/B _1435_/C _1413_/C vdd gnd NAND3X1
X_1335_ _1344_/A _1344_/B _1343_/B _1405_/C vdd gnd OAI21X1
XFILL_1__1382_ vdd gnd FILL
XFILL_1__1451_ vdd gnd FILL
X_1197_ _925_/A _1652_/B _1547_/B vdd gnd NOR2X1
XFILL_1__1520_ vdd gnd FILL
XFILL_0__1609_ vdd gnd FILL
X_1266_ _1569_/A _1569_/B _1568_/B _1593_/B vdd gnd OAI21X1
XFILL_1__1718_ vdd gnd FILL
XFILL_1__1649_ vdd gnd FILL
X_977_ _977_/A _977_/B _992_/C vdd gnd NAND2X1
XFILL_0__1891_ vdd gnd FILL
XFILL_2__1689_ vdd gnd FILL
X_1120_ _1246_/C _1195_/B _1195_/A _1123_/A vdd gnd OAI21X1
X_1051_ _1166_/B _1166_/A _1052_/B vdd gnd NAND2X1
XFILL_0__1325_ vdd gnd FILL
X_1884_ _1884_/A _1884_/B _1884_/C _1887_/B vdd gnd OAI21X1
XFILL_0__1256_ vdd gnd FILL
XFILL_0__1187_ vdd gnd FILL
X_1318_ _1410_/A _1321_/A _1377_/B _1318_/D _1334_/A vdd gnd OAI22X1
XFILL_1__989_ vdd gnd FILL
XFILL_1__1503_ vdd gnd FILL
XFILL_1__1365_ vdd gnd FILL
X_1249_ _1253_/A _1253_/B _1285_/A _1286_/B vdd gnd OAI21X1
XFILL_1__1434_ vdd gnd FILL
XFILL_1__1296_ vdd gnd FILL
XFILL_2__1474_ vdd gnd FILL
XFILL_0__1110_ vdd gnd FILL
XFILL_0__1041_ vdd gnd FILL
XFILL_0__1874_ vdd gnd FILL
X_1034_ _988_/C _988_/A _994_/A _1048_/C vdd gnd AOI21X1
X_1103_ _982_/A _1548_/D _1193_/B _1107_/C vdd gnd OAI21X1
XFILL_0__1308_ vdd gnd FILL
XFILL_1__1150_ vdd gnd FILL
X_1867_ _1867_/A _1868_/C vdd gnd INVX1
XFILL_1__1081_ vdd gnd FILL
XFILL_0__1239_ vdd gnd FILL
X_1798_ _1798_/A _1814_/B vdd gnd INVX1
XFILL_1__1417_ vdd gnd FILL
XFILL_0__930_ vdd gnd FILL
XFILL_1__1348_ vdd gnd FILL
XFILL_1__1279_ vdd gnd FILL
XFILL_0__1590_ vdd gnd FILL
X_1721_ _1752_/A _958_/B _1842_/C _1722_/C vdd gnd OAI21X1
X_1652_ LoadB_i _1652_/B _1652_/C _1684_/D vdd gnd OAI21X1
X_1583_ _1583_/A _1583_/B _1584_/B vdd gnd NOR2X1
XFILL_0__1024_ vdd gnd FILL
XFILL_0__1857_ vdd gnd FILL
XFILL_0__1788_ vdd gnd FILL
X_1017_ _1062_/A _979_/B _980_/C _1023_/A vdd gnd NAND3X1
XFILL_1__1202_ vdd gnd FILL
XFILL_1__1133_ vdd gnd FILL
XFILL_1__1064_ vdd gnd FILL
XFILL_1__1897_ vdd gnd FILL
XFILL_2__1311_ vdd gnd FILL
XFILL_0__1642_ vdd gnd FILL
XFILL_0__1711_ vdd gnd FILL
XFILL_0__1573_ vdd gnd FILL
XFILL_0__1007_ vdd gnd FILL
X_1704_ _961_/A _1750_/A _1704_/C _1727_/A vdd gnd AOI21X1
X_1635_ LoadA_i _1635_/B _1635_/C _1676_/D vdd gnd OAI21X1
X_1497_ _1498_/C _1544_/A _1504_/C vdd gnd OR2X2
XFILL_1__1751_ vdd gnd FILL
XFILL_1__1820_ vdd gnd FILL
X_1566_ _1566_/A _1566_/B _1666_/D vdd gnd NAND2X1
XFILL_1__1116_ vdd gnd FILL
XFILL_1__1047_ vdd gnd FILL
X_1420_ _1420_/A _1420_/B _1420_/C _1421_/C vdd gnd OAI21X1
X_1351_ _1351_/A _1351_/B _1351_/C _1520_/D vdd gnd OAI21X1
XFILL_0__1625_ vdd gnd FILL
X_1282_ _1282_/A _1592_/C MulH_i _1283_/A vdd gnd AOI21X1
XFILL_0__1556_ vdd gnd FILL
XFILL_0__1487_ vdd gnd FILL
X_1618_ LoadCmd_i ABCmd_i[7] _1619_/C vdd gnd NAND2X1
X_1549_ _1589_/A _1589_/B _1549_/C _1576_/B vdd gnd OAI21X1
XFILL86550x39750 vdd gnd FILL
XFILL_1__1734_ vdd gnd FILL
XFILL_1__1803_ vdd gnd FILL
XFILL86550x82950 vdd gnd FILL
XFILL_1__1596_ vdd gnd FILL
XBUFX2_insert10 _1660_/Q _952_/A vdd gnd BUFX2
X_993_ _993_/A _993_/B _998_/A vdd gnd NAND2X1
XFILL_2__1774_ vdd gnd FILL
XFILL_0__1410_ vdd gnd FILL
XFILL_0__1272_ vdd gnd FILL
XFILL_0__1341_ vdd gnd FILL
X_1403_ _1462_/C _1439_/B _1439_/A _1468_/B vdd gnd NAND3X1
X_1334_ _1334_/A _1409_/A _1343_/B vdd gnd AND2X2
X_1265_ _1265_/A _1265_/B _1265_/C _1568_/B vdd gnd NAND3X1
XFILL_1__1381_ vdd gnd FILL
XFILL_1__1450_ vdd gnd FILL
X_1196_ _1843_/B _1652_/B vdd gnd INVX1
XFILL_0__1539_ vdd gnd FILL
XFILL_0__1608_ vdd gnd FILL
XFILL_1__1648_ vdd gnd FILL
XFILL_1__1717_ vdd gnd FILL
XFILL_1__1579_ vdd gnd FILL
XFILL_2__1826_ vdd gnd FILL
XFILL_0__1890_ vdd gnd FILL
X_976_ _976_/A _977_/B vdd gnd INVX2
X_1050_ _1118_/A _1118_/C _1055_/B _1166_/B vdd gnd NAND3X1
XFILL_0__1186_ vdd gnd FILL
XFILL_0__1324_ vdd gnd FILL
X_1883_ _1885_/A _1884_/C vdd gnd INVX1
XFILL_0__1255_ vdd gnd FILL
XFILL_1__988_ vdd gnd FILL
X_1317_ _952_/A _1881_/B _964_/B _1321_/A vdd gnd NAND3X1
XFILL_1__1502_ vdd gnd FILL
X_1248_ _1248_/A _1248_/B _1341_/A _1253_/B vdd gnd AOI21X1
XFILL_1__1295_ vdd gnd FILL
XFILL_1__1364_ vdd gnd FILL
XFILL_1__1433_ vdd gnd FILL
X_1179_ _1482_/A _1428_/B vdd gnd INVX1
XFILL_2__1611_ vdd gnd FILL
XFILL_0__1040_ vdd gnd FILL
X_959_ _962_/A _961_/A _962_/B _967_/B vdd gnd NAND3X1
XFILL_0__1873_ vdd gnd FILL
X_1102_ _1109_/C _1193_/B vdd gnd INVX1
X_1033_ _1049_/A _1049_/B _998_/Y _1118_/B vdd gnd AOI21X1
XFILL_0__1307_ vdd gnd FILL
XFILL_0__1169_ vdd gnd FILL
X_1866_ _1866_/A _1866_/B _1866_/C _1868_/B vdd gnd AOI21X1
X_1797_ _1851_/A _1797_/B _1797_/C _1814_/A vdd gnd OAI21X1
XFILL_1__1080_ vdd gnd FILL
XFILL_0__1238_ vdd gnd FILL
XFILL_1__1416_ vdd gnd FILL
XFILL_1__1347_ vdd gnd FILL
XFILL_1__1278_ vdd gnd FILL
X_1651_ ABCmd_i[7] LoadB_i _1652_/C vdd gnd NAND2X1
XFILL_0__989_ vdd gnd FILL
XFILL_0__1023_ vdd gnd FILL
X_1720_ _1720_/A _1720_/B _1720_/C _1740_/B vdd gnd OAI21X1
X_1582_ _1585_/A _1582_/B _1582_/C _1595_/C vdd gnd OAI21X1
XFILL_0__1856_ vdd gnd FILL
XFILL_0__1787_ vdd gnd FILL
XFILL_1__1132_ vdd gnd FILL
X_1016_ _1026_/A _1101_/A vdd gnd INVX1
XFILL_1__1201_ vdd gnd FILL
X_1849_ _1885_/C _1885_/B _1873_/A vdd gnd AND2X2
XFILL_1__1063_ vdd gnd FILL
XFILL_1__1896_ vdd gnd FILL
XFILL_0__1641_ vdd gnd FILL
XFILL_0__1710_ vdd gnd FILL
XFILL_0__1572_ vdd gnd FILL
X_1634_ ABCmd_i[7] LoadA_i _1635_/C vdd gnd NAND2X1
XFILL_0__1006_ vdd gnd FILL
X_1703_ _961_/A _1750_/A _1842_/C _1704_/C vdd gnd OAI21X1
X_1496_ _1548_/D _1545_/B _1546_/B _1498_/C vdd gnd OAI21X1
X_1565_ MulH_i _1565_/B _1565_/C _1566_/B vdd gnd NAND3X1
XFILL_1__1750_ vdd gnd FILL
XFILL_0__1839_ vdd gnd FILL
XFILL_1__1046_ vdd gnd FILL
XFILL_1__1115_ vdd gnd FILL
XFILL_1__1879_ vdd gnd FILL
X_1350_ _1354_/C _1420_/C _1354_/A _1351_/B vdd gnd AOI21X1
X_1281_ _1873_/A _1739_/Y Flag_i _1282_/A vdd gnd MUX2X1
XFILL_0__1555_ vdd gnd FILL
XFILL_0__1624_ vdd gnd FILL
XFILL_0__1486_ vdd gnd FILL
X_1617_ LoadCmd_i _1617_/B _1617_/C _1659_/D vdd gnd OAI21X1
XFILL_1__1802_ vdd gnd FILL
X_1548_ _1652_/B _1548_/B _1635_/B _1548_/D _1549_/C vdd gnd OAI22X1
X_1479_ _1479_/A _1479_/B _1487_/B vdd gnd NAND2X1
XFILL_1__1733_ vdd gnd FILL
XFILL_1__1595_ vdd gnd FILL
XFILL_2__986_ vdd gnd FILL
XFILL_1__1029_ vdd gnd FILL
XBUFX2_insert11 _1655_/Q _1809_/A vdd gnd BUFX2
X_992_ _992_/A _992_/B _992_/C _993_/A vdd gnd OAI21X1
XFILL_0__1271_ vdd gnd FILL
XFILL_0__1340_ vdd gnd FILL
XFILL_2__1207_ vdd gnd FILL
X_1402_ _1460_/A _1462_/C vdd gnd INVX1
XFILL_2__1069_ vdd gnd FILL
X_1264_ _1265_/A _1265_/B _1569_/B vdd gnd NAND2X1
X_1333_ _1333_/A _1333_/B _1344_/A vdd gnd AND2X2
XFILL_0__1469_ vdd gnd FILL
XFILL_1__1380_ vdd gnd FILL
XFILL_0__1607_ vdd gnd FILL
XFILL_0__1538_ vdd gnd FILL
X_1195_ _1195_/A _1195_/B _1195_/C _1352_/C vdd gnd OAI21X1
XFILL_1__1647_ vdd gnd FILL
XFILL_1__1578_ vdd gnd FILL
XFILL_1__1716_ vdd gnd FILL
X_975_ _975_/A _975_/B _976_/A vdd gnd NAND2X1
XFILL_0__1323_ vdd gnd FILL
XFILL_0__1185_ vdd gnd FILL
X_1882_ _1882_/A _1882_/B _1885_/A vdd gnd NAND2X1
XFILL_0__1254_ vdd gnd FILL
XFILL_1__987_ vdd gnd FILL
X_1316_ _1319_/B _1319_/C _1319_/A _1377_/B vdd gnd AOI21X1
XFILL_1__1501_ vdd gnd FILL
XFILL_1__1432_ vdd gnd FILL
X_1247_ _1341_/C _1290_/B _1290_/A _1253_/A vdd gnd AOI21X1
X_1178_ _1429_/A _1427_/B _1427_/A _1482_/A vdd gnd NAND3X1
XFILL_1__1363_ vdd gnd FILL
XFILL_1__1294_ vdd gnd FILL
X_958_ _980_/A _958_/B _958_/C _967_/A vdd gnd NAND3X1
XFILL_0__1872_ vdd gnd FILL
X_1032_ _1095_/C _1056_/A _1056_/B _1049_/B vdd gnd OAI21X1
X_1101_ _1101_/A _1101_/B _1101_/C _1109_/C vdd gnd AOI21X1
XFILL_0__1306_ vdd gnd FILL
XFILL_0__1168_ vdd gnd FILL
XFILL_0__1237_ vdd gnd FILL
X_1865_ _1865_/A _1866_/C vdd gnd INVX1
X_1796_ _1858_/A _1850_/B _1797_/B vdd gnd NAND2X1
XFILL_0__1099_ vdd gnd FILL
XFILL_1__1415_ vdd gnd FILL
XFILL_0_BUFX2_insert10 vdd gnd FILL
XFILL_1__1346_ vdd gnd FILL
XFILL_1__1277_ vdd gnd FILL
XFILL85650x39750 vdd gnd FILL
XFILL85650x82950 vdd gnd FILL
XFILL_2__1455_ vdd gnd FILL
X_1650_ LoadB_i _1650_/B _1650_/C _1683_/D vdd gnd OAI21X1
XFILL_0__988_ vdd gnd FILL
X_1581_ _1586_/B _1582_/C vdd gnd INVX1
XFILL_0__1022_ vdd gnd FILL
XFILL_0__1855_ vdd gnd FILL
X_1015_ _1062_/A _977_/A _979_/C _1026_/A vdd gnd NAND3X1
XFILL_0__1786_ vdd gnd FILL
XFILL_1__1131_ vdd gnd FILL
XFILL_1__1062_ vdd gnd FILL
XFILL_1__1200_ vdd gnd FILL
X_1779_ _1779_/A _1779_/B _1779_/C _1793_/A vdd gnd NAND3X1
X_1848_ _1859_/A _1876_/B _1848_/C _1885_/B vdd gnd NAND3X1
XFILL_1__1895_ vdd gnd FILL
XFILL_1__1329_ vdd gnd FILL
XFILL_2__1507_ vdd gnd FILL
XFILL_0__1640_ vdd gnd FILL
XFILL_0__1571_ vdd gnd FILL
X_1633_ LoadA_i _1633_/B _1633_/C _1675_/D vdd gnd OAI21X1
X_1564_ _1564_/A _1564_/B _1573_/C _1565_/C vdd gnd OAI21X1
XFILL_0__1005_ vdd gnd FILL
X_1702_ _1702_/A _1702_/B _1733_/A _1734_/A vdd gnd OAI21X1
X_1495_ _1495_/A _1495_/B _1589_/A _1546_/B vdd gnd OAI21X1
XFILL_0__1838_ vdd gnd FILL
XFILL_0__1769_ vdd gnd FILL
XFILL_1__1114_ vdd gnd FILL
XFILL_1__1045_ vdd gnd FILL
XFILL_1__1878_ vdd gnd FILL
XFILL_2__1154_ vdd gnd FILL
X_1280_ _1429_/A _1280_/B MulL_i _1283_/B vdd gnd OAI21X1
XFILL_0__1554_ vdd gnd FILL
XFILL_0__1623_ vdd gnd FILL
XFILL_0__1485_ vdd gnd FILL
X_1616_ LoadCmd_i ABCmd_i[6] _1617_/C vdd gnd NAND2X1
X_1547_ _1881_/B _1547_/B _1589_/B vdd gnd NAND2X1
XFILL_1__1801_ vdd gnd FILL
X_1478_ _1478_/A _1478_/B _1478_/C _1479_/B vdd gnd OAI21X1
XFILL_1__1732_ vdd gnd FILL
XFILL_1__1594_ vdd gnd FILL
XFILL_1__1028_ vdd gnd FILL
XBUFX2_insert12 _1655_/Q _1843_/A vdd gnd BUFX2
X_991_ _991_/A _991_/B _991_/C _993_/B vdd gnd NAND3X1
XFILL_0__1270_ vdd gnd FILL
X_1401_ _1406_/B _1406_/A _1439_/A vdd gnd AND2X2
X_1332_ _1332_/A _1332_/B _1369_/A vdd gnd AND2X2
XFILL_0__1606_ vdd gnd FILL
X_1194_ _1194_/A _1194_/B _1194_/C _1286_/A vdd gnd OAI21X1
X_1263_ _1591_/A _1267_/A vdd gnd INVX1
XFILL_0__1468_ vdd gnd FILL
XFILL_0__1537_ vdd gnd FILL
XFILL_0__1399_ vdd gnd FILL
XFILL86850x68550 vdd gnd FILL
XFILL_1__1715_ vdd gnd FILL
XFILL_1__1646_ vdd gnd FILL
XFILL86250x64950 vdd gnd FILL
XFILL_1__1577_ vdd gnd FILL
X_974_ _989_/C _989_/B _989_/A _988_/A vdd gnd NAND3X1
XFILL_2__1755_ vdd gnd FILL
XFILL_0__1322_ vdd gnd FILL
XFILL_0__1184_ vdd gnd FILL
X_1881_ _1881_/A _1881_/B _1882_/B vdd gnd OR2X2
XFILL_0__1253_ vdd gnd FILL
X_1315_ _980_/B _1372_/A _1577_/A _1319_/C vdd gnd NAND3X1
XFILL_1__986_ vdd gnd FILL
XFILL_1__1500_ vdd gnd FILL
X_1246_ _1246_/A _1246_/B _1246_/C _1285_/A vdd gnd AOI21X1
XFILL_1__1431_ vdd gnd FILL
XFILL_1__1362_ vdd gnd FILL
X_1177_ _1641_/B _976_/A _1177_/C _1427_/B vdd gnd OAI21X1
XFILL_1__1293_ vdd gnd FILL
XFILL86850x43350 vdd gnd FILL
XFILL_2__1540_ vdd gnd FILL
XFILL_1__1629_ vdd gnd FILL
X_957_ _957_/A _957_/B _957_/C _990_/C vdd gnd OAI21X1
XFILL_0__1871_ vdd gnd FILL
XFILL_2__1807_ vdd gnd FILL
X_1031_ _1031_/A _1031_/B _1056_/B vdd gnd AND2X2
X_1100_ _1194_/A _1107_/A vdd gnd INVX1
XFILL_0__1305_ vdd gnd FILL
XFILL_0__1236_ vdd gnd FILL
XFILL_0__1167_ vdd gnd FILL
X_1795_ _1795_/A _1795_/B _1795_/C _1850_/B vdd gnd OAI21X1
X_1864_ _1864_/A _1867_/A _1864_/C _1872_/A vdd gnd NAND3X1
XFILL_0__1098_ vdd gnd FILL
XFILL_1__969_ vdd gnd FILL
XFILL_0_BUFX2_insert11 vdd gnd FILL
XFILL_1__1414_ vdd gnd FILL
XFILL_1__1345_ vdd gnd FILL
X_1229_ _1410_/A _1233_/B _1333_/B _1238_/A vdd gnd OAI21X1
XFILL_1__1276_ vdd gnd FILL
XFILL_0__987_ vdd gnd FILL
X_1580_ _1589_/C _1580_/B _1586_/B vdd gnd NAND2X1
XFILL_0__1021_ vdd gnd FILL
XFILL_0__1854_ vdd gnd FILL
XFILL_0__1785_ vdd gnd FILL
X_1014_ _1029_/A _1029_/B _1029_/C _1056_/C vdd gnd NAND3X1
XFILL_1__1130_ vdd gnd FILL
XFILL_0__1219_ vdd gnd FILL
X_1847_ _1874_/C _1854_/A _1847_/C _1885_/C vdd gnd OAI21X1
XFILL_1__1061_ vdd gnd FILL
X_1778_ _1778_/A _1795_/C _1871_/C _1779_/C vdd gnd AOI21X1
XFILL_1__1894_ vdd gnd FILL
XFILL_1__1328_ vdd gnd FILL
XFILL_1__1259_ vdd gnd FILL
XFILL_0__1570_ vdd gnd FILL
X_1701_ _979_/C _1836_/A _1733_/A vdd gnd NAND2X1
X_1632_ ABCmd_i[6] LoadA_i _1633_/C vdd gnd NAND2X1
X_1563_ _1575_/C _1563_/B _1573_/C vdd gnd AND2X2
X_1494_ _1826_/B _1577_/A _1589_/A vdd gnd NAND2X1
XFILL_0__1004_ vdd gnd FILL
XFILL_0__1768_ vdd gnd FILL
XFILL_0__1837_ vdd gnd FILL
XFILL_0__1699_ vdd gnd FILL
XFILL_1__1113_ vdd gnd FILL
XFILL_1__1044_ vdd gnd FILL
XFILL_1__1877_ vdd gnd FILL
XFILL_0__1622_ vdd gnd FILL
XFILL_0__1553_ vdd gnd FILL
XFILL_0__1484_ vdd gnd FILL
X_1615_ _1858_/A _1617_/B vdd gnd INVX1
X_1546_ _1546_/A _1546_/B _1546_/C _1554_/A vdd gnd AOI21X1
X_1477_ _1524_/A _1478_/C vdd gnd INVX1
XFILL_1__1731_ vdd gnd FILL
XFILL_1__1800_ vdd gnd FILL
XFILL_1__1593_ vdd gnd FILL
XBUFX2_insert13 _1655_/Q _1750_/A vdd gnd BUFX2
X_990_ _990_/A _990_/B _990_/C _998_/B vdd gnd AOI21X1
XFILL_1__1027_ vdd gnd FILL
X_1400_ _1460_/A _1462_/A _1462_/B _1468_/A vdd gnd OAI21X1
X_1331_ _1369_/C _1405_/B _1405_/A _1419_/A vdd gnd OAI21X1
XFILL_0__1605_ vdd gnd FILL
X_1193_ _1193_/A _1193_/B _1194_/B vdd gnd NOR2X1
X_1262_ _1262_/A _1591_/B vdd gnd INVX1
XFILL_0__1398_ vdd gnd FILL
XFILL_0__1467_ vdd gnd FILL
XFILL_0__1536_ vdd gnd FILL
XFILL_1__1645_ vdd gnd FILL
X_1529_ _1529_/A _1539_/A vdd gnd INVX1
XFILL_1__1714_ vdd gnd FILL
XFILL_1__1576_ vdd gnd FILL
X_973_ _999_/A _973_/B _973_/C _989_/B vdd gnd NAND3X1
XFILL_0__1321_ vdd gnd FILL
X_1880_ _1881_/B _1881_/A _1882_/A vdd gnd NAND2X1
XFILL_0__1252_ vdd gnd FILL
XFILL_0__1183_ vdd gnd FILL
X_1314_ _923_/A _1823_/A _1577_/A vdd gnd AND2X2
XFILL_1__985_ vdd gnd FILL
XFILL_0__1519_ vdd gnd FILL
XFILL_1__1361_ vdd gnd FILL
X_1176_ _964_/B _1641_/B vdd gnd INVX1
X_1245_ _1352_/A _1352_/B _1352_/C _1353_/C vdd gnd NAND3X1
XFILL_1__1430_ vdd gnd FILL
XFILL_1__1292_ vdd gnd FILL
XFILL_1__1628_ vdd gnd FILL
XFILL_1__1559_ vdd gnd FILL
X_956_ _956_/A _956_/B _956_/C _996_/C vdd gnd OAI21X1
XFILL_0__1870_ vdd gnd FILL
X_1030_ _1030_/A _1030_/B _999_/Y _1095_/C vdd gnd AOI21X1
XFILL_0__1304_ vdd gnd FILL
X_1863_ _1863_/A _1863_/B _1867_/A vdd gnd NOR2X1
XFILL_0__1166_ vdd gnd FILL
XFILL_0__1235_ vdd gnd FILL
X_1794_ _1794_/A _1794_/B _1795_/A vdd gnd NOR2X1
XFILL_0__1097_ vdd gnd FILL
XFILL_1__968_ vdd gnd FILL
X_1228_ _1228_/A _1228_/B _1228_/C _1333_/B vdd gnd OAI21X1
XFILL_0_BUFX2_insert12 vdd gnd FILL
XFILL_1__1413_ vdd gnd FILL
X_1159_ _1183_/B _1183_/C _1183_/A _1187_/A vdd gnd NAND3X1
XFILL_1__1344_ vdd gnd FILL
XFILL_1__1275_ vdd gnd FILL
XFILL_0__986_ vdd gnd FILL
XFILL_0__1020_ vdd gnd FILL
X_939_ _957_/A _971_/A vdd gnd INVX1
XFILL_0__1853_ vdd gnd FILL
XFILL_0__1784_ vdd gnd FILL
X_1013_ _1057_/C _1070_/B _1070_/A _1029_/B vdd gnd OAI21X1
XFILL_0__1218_ vdd gnd FILL
XFILL_0__1149_ vdd gnd FILL
XFILL_1__1060_ vdd gnd FILL
X_1846_ _1876_/B _1847_/C vdd gnd INVX1
X_1777_ _1858_/A _1871_/C vdd gnd INVX1
XFILL_1__1893_ vdd gnd FILL
XFILL_1__1327_ vdd gnd FILL
XFILL_1__1258_ vdd gnd FILL
XFILL_1__1189_ vdd gnd FILL
X_1631_ LoadA_i _1631_/B _1631_/C _1674_/D vdd gnd OAI21X1
XFILL_0__969_ vdd gnd FILL
XFILL_2__1298_ vdd gnd FILL
XFILL_0__1003_ vdd gnd FILL
X_1700_ _1863_/B _1732_/B _1702_/B vdd gnd NAND2X1
X_1562_ _1574_/A _1574_/B _1583_/B _1564_/B vdd gnd AOI21X1
X_1493_ _962_/B _1547_/B _1544_/A vdd gnd NAND2X1
XFILL_0__1836_ vdd gnd FILL
XFILL_0__1767_ vdd gnd FILL
XFILL_0__1698_ vdd gnd FILL
XFILL_1__1112_ vdd gnd FILL
X_1829_ _1861_/B _1874_/B vdd gnd INVX1
XFILL_1__1043_ vdd gnd FILL
XFILL_1__1876_ vdd gnd FILL
XFILL_0__1552_ vdd gnd FILL
XFILL_0__1621_ vdd gnd FILL
XFILL_0__1483_ vdd gnd FILL
X_1614_ LoadCmd_i _1614_/B _1614_/C _1658_/D vdd gnd OAI21X1
X_1545_ _1548_/D _1545_/B _1546_/C vdd gnd NOR2X1
X_1476_ _1476_/A _1476_/B _1524_/B _1478_/B vdd gnd AOI21X1
XFILL_1__1730_ vdd gnd FILL
XFILL_0__1819_ vdd gnd FILL
XFILL86850x28950 vdd gnd FILL
XFILL_1__1592_ vdd gnd FILL
XBUFX2_insert14 _1655_/Q _1752_/A vdd gnd BUFX2
XFILL_1__1026_ vdd gnd FILL
XFILL_1__1859_ vdd gnd FILL
XFILL_2__1135_ vdd gnd FILL
X_1330_ _1334_/A _1409_/A _1330_/C _1405_/B vdd gnd AOI21X1
X_1261_ _1363_/A _1526_/A _1358_/A vdd gnd NAND2X1
XFILL_0__1604_ vdd gnd FILL
XFILL_0__1535_ vdd gnd FILL
X_1192_ _1192_/A _1192_/B _1192_/C _1255_/C vdd gnd AOI21X1
XFILL_0__1466_ vdd gnd FILL
XFILL_0__1397_ vdd gnd FILL
X_1459_ _1463_/A _1510_/A _1488_/B vdd gnd NAND2X1
X_1528_ _1528_/A _1560_/C _1536_/B vdd gnd NAND2X1
XFILL_1__1644_ vdd gnd FILL
XFILL_1__1713_ vdd gnd FILL
XFILL_1__1575_ vdd gnd FILL
XFILL_2__966_ vdd gnd FILL
XFILL_1__1009_ vdd gnd FILL
X_972_ _999_/C _972_/B _999_/B _989_/A vdd gnd OAI21X1
XFILL_0__1320_ vdd gnd FILL
XFILL_0__1182_ vdd gnd FILL
XFILL_0__1251_ vdd gnd FILL
XFILL_1__984_ vdd gnd FILL
X_1313_ _962_/B _1372_/B _922_/B _1319_/B vdd gnd NAND3X1
X_1244_ _1290_/A _1290_/B _1341_/C _1352_/B vdd gnd NAND3X1
XFILL_0__1518_ vdd gnd FILL
XFILL_1__1291_ vdd gnd FILL
XFILL_1__1360_ vdd gnd FILL
X_1175_ _1279_/B _1279_/A _1429_/A vdd gnd NOR2X1
XFILL_0__1449_ vdd gnd FILL
XFILL_1__1558_ vdd gnd FILL
XFILL_1__1627_ vdd gnd FILL
XFILL_1__1489_ vdd gnd FILL
X_955_ _955_/A _955_/B _955_/C _956_/B vdd gnd AOI21X1
XFILL_0__1303_ vdd gnd FILL
XFILL_2__1598_ vdd gnd FILL
X_1793_ _1793_/A _1797_/C _1798_/A _1813_/B vdd gnd AOI21X1
X_1862_ _1865_/A _1874_/A _1864_/C vdd gnd NAND2X1
XFILL_0__1165_ vdd gnd FILL
XFILL_0__1234_ vdd gnd FILL
XFILL_0__1096_ vdd gnd FILL
X_1158_ _1158_/A _956_/B _956_/A _1183_/A vdd gnd OAI21X1
XFILL_1__1412_ vdd gnd FILL
XFILL_1__967_ vdd gnd FILL
XFILL_0_BUFX2_insert13 vdd gnd FILL
X_1227_ _1233_/C _1333_/A _1238_/B vdd gnd NAND2X1
XFILL_1__1343_ vdd gnd FILL
X_1089_ _1201_/D _1201_/C _1089_/C _1092_/A vdd gnd NAND3X1
XFILL_1__1274_ vdd gnd FILL
XFILL86550x25350 vdd gnd FILL
XFILL_2__1383_ vdd gnd FILL
XFILL_0__985_ vdd gnd FILL
X_938_ _980_/A _964_/B _980_/C _957_/A vdd gnd NAND3X1
X_1012_ _1057_/A _1057_/B _1070_/C _1029_/A vdd gnd NAND3X1
XFILL_0__1852_ vdd gnd FILL
XFILL_0__1783_ vdd gnd FILL
XFILL_0__1148_ vdd gnd FILL
XFILL_0__1079_ vdd gnd FILL
XFILL_0__1217_ vdd gnd FILL
X_1845_ _1878_/B _1877_/A _1859_/C _1876_/B vdd gnd OAI21X1
X_1776_ _1851_/A _1776_/Y vdd gnd INVX1
XFILL_1__1892_ vdd gnd FILL
XFILL_1__1326_ vdd gnd FILL
XFILL_1__1188_ vdd gnd FILL
XFILL_1__1257_ vdd gnd FILL
XFILL_2__1435_ vdd gnd FILL
XFILL_0_BUFX2_insert5 vdd gnd FILL
X_1630_ ABCmd_i[5] LoadA_i _1631_/C vdd gnd NAND2X1
XFILL_0__968_ vdd gnd FILL
XFILL_0__1002_ vdd gnd FILL
X_1492_ _1543_/A _1508_/C vdd gnd INVX1
X_1561_ _1575_/A _1564_/A vdd gnd INVX1
XFILL_0__1835_ vdd gnd FILL
XFILL_0__1766_ vdd gnd FILL
XFILL_0__1697_ vdd gnd FILL
XFILL_1__1042_ vdd gnd FILL
XFILL_1__1111_ vdd gnd FILL
X_1828_ _1828_/A _1828_/B _1859_/A _1861_/B vdd gnd OAI21X1
X_1759_ _1778_/A _1759_/Y vdd gnd INVX1
XFILL_1__1875_ vdd gnd FILL
XFILL_2__1220_ vdd gnd FILL
XFILL_1__1309_ vdd gnd FILL
XFILL_2__1082_ vdd gnd FILL
XFILL_0__1551_ vdd gnd FILL
XFILL_0__1620_ vdd gnd FILL
XFILL_0__1482_ vdd gnd FILL
X_1613_ LoadCmd_i ABCmd_i[5] _1614_/C vdd gnd NAND2X1
X_1544_ _1544_/A _1546_/A vdd gnd INVX1
X_1475_ _1526_/A _1526_/C _1476_/A vdd gnd NAND2X1
XFILL_0__1818_ vdd gnd FILL
XFILL_1__1591_ vdd gnd FILL
XFILL_0__1749_ vdd gnd FILL
XFILL_1__1025_ vdd gnd FILL
XFILL_1__1858_ vdd gnd FILL
XFILL_1__1789_ vdd gnd FILL
X_1191_ _1591_/A _1191_/B _1262_/A _1526_/A vdd gnd OAI21X1
X_1260_ _1268_/B _1523_/A _1363_/A vdd gnd AND2X2
XFILL_0__1465_ vdd gnd FILL
XFILL_0__1534_ vdd gnd FILL
XFILL_0__1603_ vdd gnd FILL
XFILL_0__1396_ vdd gnd FILL
X_1527_ _1583_/B _1574_/B _1574_/A _1528_/A vdd gnd NAND3X1
X_1458_ _1463_/A _1510_/A _1488_/A _1461_/C vdd gnd NAND3X1
X_1389_ _1394_/A _1394_/B _1442_/C vdd gnd OR2X2
XFILL_1__1574_ vdd gnd FILL
XFILL_1__1643_ vdd gnd FILL
XFILL_1__1712_ vdd gnd FILL
XFILL_1__1008_ vdd gnd FILL
X_971_ _971_/A _971_/B _971_/C _989_/C vdd gnd AOI21X1
XFILL_0__1181_ vdd gnd FILL
XFILL_0__1250_ vdd gnd FILL
X_1312_ _1320_/C _1378_/B _1378_/A _1318_/D vdd gnd AOI21X1
XFILL_1__983_ vdd gnd FILL
X_1174_ _961_/A _926_/B _1279_/A vdd gnd NAND2X1
X_1243_ _1289_/A _1344_/B _1289_/C _1290_/B vdd gnd OAI21X1
XFILL_0__1448_ vdd gnd FILL
XFILL_0__1517_ vdd gnd FILL
XFILL_1__1290_ vdd gnd FILL
XFILL_0__1379_ vdd gnd FILL
XFILL_1__1557_ vdd gnd FILL
XFILL_1__1626_ vdd gnd FILL
XFILL_1__1488_ vdd gnd FILL
X_954_ _954_/A _997_/A _956_/A vdd gnd NAND2X1
XFILL_2__1735_ vdd gnd FILL
XFILL_0__1302_ vdd gnd FILL
XFILL_0__1164_ vdd gnd FILL
XFILL_0__1095_ vdd gnd FILL
X_1861_ _1876_/B _1861_/B _1865_/A vdd gnd NOR2X1
X_1792_ _1792_/A _1792_/B _1801_/A _1798_/A vdd gnd OAI21X1
XFILL_0__1233_ vdd gnd FILL
XFILL_1__966_ vdd gnd FILL
XFILL_1__1411_ vdd gnd FILL
X_1157_ _1181_/C _1181_/A _1180_/A _1183_/C vdd gnd OAI21X1
XFILL_1__1342_ vdd gnd FILL
XFILL_0_BUFX2_insert14 vdd gnd FILL
X_1226_ _1410_/A _1233_/B _1333_/A vdd gnd NOR2X1
X_1088_ _1088_/A _1088_/B _1088_/C _1209_/C vdd gnd AOI21X1
XFILL_1__1273_ vdd gnd FILL
XFILL_2__1520_ vdd gnd FILL
XFILL_1__1609_ vdd gnd FILL
XFILL_0__984_ vdd gnd FILL
XFILL_0__1851_ vdd gnd FILL
X_937_ _937_/A _937_/B _937_/C _955_/C vdd gnd OAI21X1
X_1011_ _973_/B _972_/B _973_/C _1029_/C vdd gnd OAI21X1
XFILL_0__1782_ vdd gnd FILL
XFILL_0__1216_ vdd gnd FILL
XFILL_0__1147_ vdd gnd FILL
XFILL_0__1078_ vdd gnd FILL
X_1844_ _1878_/A _1877_/A _1878_/B _1859_/C vdd gnd OAI21X1
X_1775_ _1779_/B _1779_/A _1851_/A vdd gnd NAND2X1
XFILL_1__949_ vdd gnd FILL
XFILL_1__1891_ vdd gnd FILL
XFILL_1__1325_ vdd gnd FILL
X_1209_ _1209_/A _1209_/B _1209_/C _1289_/C vdd gnd AOI21X1
XFILL_1__1187_ vdd gnd FILL
XFILL_1__1256_ vdd gnd FILL
XFILL_0_BUFX2_insert6 vdd gnd FILL
X_1560_ _1575_/A _1583_/A _1560_/C _1565_/B vdd gnd NAND3X1
XFILL_0__967_ vdd gnd FILL
XFILL_0__1001_ vdd gnd FILL
X_1491_ _1491_/A _1491_/B _1491_/C _1543_/A vdd gnd OAI21X1
XFILL_0__1834_ vdd gnd FILL
XFILL_0__1765_ vdd gnd FILL
XFILL_0__1696_ vdd gnd FILL
XFILL_1__1041_ vdd gnd FILL
X_1827_ _1878_/A _1828_/B _1828_/A _1859_/A vdd gnd OAI21X1
XFILL_1__1110_ vdd gnd FILL
X_1758_ _1780_/B _1758_/B _1778_/A vdd gnd NAND2X1
XFILL_1__1874_ vdd gnd FILL
X_1689_ _1734_/D _1713_/A vdd gnd INVX1
XFILL_1__1308_ vdd gnd FILL
XFILL_1__1239_ vdd gnd FILL
XFILL_0__1550_ vdd gnd FILL
XFILL_0__1481_ vdd gnd FILL
X_1543_ _1543_/A _1543_/B _1543_/C _1558_/B vdd gnd AOI21X1
X_1474_ _1474_/A _1523_/B _1526_/C vdd gnd NOR2X1
X_1612_ _1836_/A _1614_/B vdd gnd INVX1
XFILL_0__1817_ vdd gnd FILL
XFILL_0__1748_ vdd gnd FILL
XFILL_1__1590_ vdd gnd FILL
XFILL_1__1024_ vdd gnd FILL
XFILL_1__1857_ vdd gnd FILL
XFILL_1__1788_ vdd gnd FILL
XFILL_0__1602_ vdd gnd FILL
X_1190_ _1265_/C _1568_/C _1190_/C _1191_/B vdd gnd OAI21X1
XFILL_0__1464_ vdd gnd FILL
XFILL_0__1395_ vdd gnd FILL
XFILL_0__1533_ vdd gnd FILL
X_1457_ _1457_/A _1457_/B _1457_/C _1510_/A vdd gnd NAND3X1
X_1526_ _1526_/A _1526_/B _1526_/C _1574_/B vdd gnd NAND3X1
XFILL_1__1711_ vdd gnd FILL
X_1388_ _923_/A _1881_/B _980_/B _1394_/B vdd gnd NAND3X1
XFILL_1__1573_ vdd gnd FILL
XFILL_1__1642_ vdd gnd FILL
X_970_ _990_/A _990_/B _990_/C _998_/C vdd gnd NAND3X1
XFILL_1__1007_ vdd gnd FILL
XFILL_2__1820_ vdd gnd FILL
XFILL_0__1180_ vdd gnd FILL
X_1311_ _1631_/B _982_/B _1372_/B _1378_/B vdd gnd OAI21X1
XFILL_1__982_ vdd gnd FILL
X_1242_ _1340_/A _1340_/B _1340_/C _1341_/C vdd gnd NAND3X1
X_1173_ _958_/B _977_/B _1279_/B vdd gnd NAND2X1
XFILL_0__1447_ vdd gnd FILL
XFILL_0__1378_ vdd gnd FILL
XFILL_0__1516_ vdd gnd FILL
X_1509_ _1510_/B _1510_/A _1511_/C vdd gnd OR2X2
XFILL_1__1556_ vdd gnd FILL
XFILL_1__1625_ vdd gnd FILL
XFILL_1__1487_ vdd gnd FILL
X_953_ _953_/A _982_/B _953_/C _954_/A vdd gnd OAI21X1
XFILL_0__1301_ vdd gnd FILL
X_1860_ _1868_/A _1864_/A vdd gnd INVX1
XFILL_0__1232_ vdd gnd FILL
XFILL_0__1163_ vdd gnd FILL
XFILL_0__1094_ vdd gnd FILL
X_1791_ _1878_/A _1792_/B _1792_/A _1801_/A vdd gnd OAI21X1
XFILL_1__965_ vdd gnd FILL
XFILL_1__1410_ vdd gnd FILL
X_1156_ _1156_/A _1156_/B _1156_/C _1181_/A vdd gnd AOI21X1
X_1087_ _1087_/A _1087_/B _1087_/C _1236_/B vdd gnd AOI21X1
XFILL_1__1341_ vdd gnd FILL
X_1225_ _1327_/C _1325_/B _1233_/B vdd gnd AND2X2
XFILL_1__1272_ vdd gnd FILL
XFILL86850x79350 vdd gnd FILL
XFILL_1__1608_ vdd gnd FILL
XFILL_0__983_ vdd gnd FILL
XFILL_1__1539_ vdd gnd FILL
X_936_ _936_/A _937_/B vdd gnd INVX1
XFILL_0__1781_ vdd gnd FILL
XFILL_0__1850_ vdd gnd FILL
XFILL_2__1579_ vdd gnd FILL
X_1010_ _999_/Y _1030_/B _1030_/A _1095_/B vdd gnd NAND3X1
XFILL_0__1215_ vdd gnd FILL
X_1843_ _1843_/A _1843_/B _1843_/C _1877_/A vdd gnd AOI21X1
XFILL_0__1077_ vdd gnd FILL
XFILL_0__1146_ vdd gnd FILL
X_1774_ _1780_/A _1774_/B _1780_/B _1779_/B vdd gnd NAND3X1
XFILL_1__1890_ vdd gnd FILL
XFILL_1__948_ vdd gnd FILL
X_1208_ _1241_/B _1241_/A _1341_/A vdd gnd NAND2X1
X_1139_ _988_/A _998_/C _998_/A _1161_/B vdd gnd NAND3X1
XFILL86850x54150 vdd gnd FILL
XFILL86250x50550 vdd gnd FILL
XFILL_1__1324_ vdd gnd FILL
XFILL_1__1255_ vdd gnd FILL
XFILL_1__1186_ vdd gnd FILL
XFILL_0_BUFX2_insert7 vdd gnd FILL
XFILL_0__966_ vdd gnd FILL
XFILL_0__1000_ vdd gnd FILL
X_1490_ _1490_/A _1491_/C _1491_/B vdd gnd NAND2X1
XFILL_0__1833_ vdd gnd FILL
XFILL_0__1764_ vdd gnd FILL
XFILL_0__1695_ vdd gnd FILL
XFILL_0__1129_ vdd gnd FILL
X_1826_ _1843_/A _1826_/B _1826_/C _1828_/B vdd gnd AOI21X1
XFILL_1__1040_ vdd gnd FILL
X_1757_ _1757_/A _1757_/B _1757_/C _1758_/B vdd gnd NAND3X1
XFILL_1__1873_ vdd gnd FILL
X_1688_ _1836_/A _1709_/B _1734_/D vdd gnd NOR2X1
XFILL_1__1307_ vdd gnd FILL
XFILL_1__1238_ vdd gnd FILL
XFILL_1__1169_ vdd gnd FILL
XFILL_2__1416_ vdd gnd FILL
XFILL_0__1480_ vdd gnd FILL
XFILL_0__949_ vdd gnd FILL
X_1611_ LoadCmd_i _1611_/B _1611_/C _1657_/D vdd gnd OAI21X1
XFILL_2__1278_ vdd gnd FILL
X_1473_ _1519_/C _1478_/A vdd gnd INVX1
X_1542_ _1542_/A _1542_/B _920_/Y _1566_/A vdd gnd OAI21X1
XFILL_0__1816_ vdd gnd FILL
XFILL_0__1747_ vdd gnd FILL
XFILL_1__1023_ vdd gnd FILL
X_1809_ _1809_/A _977_/A _1809_/C _1811_/B vdd gnd AOI21X1
XFILL_1__1856_ vdd gnd FILL
XFILL_1__1787_ vdd gnd FILL
XFILL_2__1063_ vdd gnd FILL
XFILL_0__1601_ vdd gnd FILL
XFILL_0__1532_ vdd gnd FILL
XFILL_0__1463_ vdd gnd FILL
XFILL_0__1394_ vdd gnd FILL
X_1456_ _1456_/A _1457_/B vdd gnd INVX1
X_1387_ _923_/A _1823_/A _979_/B _1394_/A vdd gnd NAND3X1
X_1525_ _1525_/A _1525_/B _1526_/B _1525_/D _1574_/A vdd gnd AOI22X1
XFILL_1__1641_ vdd gnd FILL
XFILL_1__1710_ vdd gnd FILL
XFILL_1__1572_ vdd gnd FILL
XFILL_1__1006_ vdd gnd FILL
XFILL_1__1839_ vdd gnd FILL
XFILL_2__1115_ vdd gnd FILL
X_1310_ _962_/B _1631_/B vdd gnd INVX1
XFILL_1__981_ vdd gnd FILL
XFILL_2__1879_ vdd gnd FILL
X_1241_ _1241_/A _1241_/B _1290_/A vdd gnd AND2X2
XFILL_0__1515_ vdd gnd FILL
X_1172_ _1177_/C _1172_/B _1427_/A vdd gnd OR2X2
XFILL_0__1446_ vdd gnd FILL
XFILL_0__1377_ vdd gnd FILL
X_1508_ _1543_/C _1508_/B _1508_/C _1514_/B vdd gnd OAI21X1
X_1439_ _1439_/A _1439_/B _1460_/A _1488_/A vdd gnd AOI21X1
XFILL_1__1624_ vdd gnd FILL
XFILL_1__1555_ vdd gnd FILL
XFILL_1__1486_ vdd gnd FILL
XFILL_2__946_ vdd gnd FILL
X_952_ _952_/A _979_/B _982_/B vdd gnd NAND2X1
XFILL_0__1162_ vdd gnd FILL
XFILL_0__1300_ vdd gnd FILL
XFILL_0__1231_ vdd gnd FILL
X_1790_ _1843_/A _979_/B _1790_/C _1792_/B vdd gnd AOI21X1
XFILL_0__1093_ vdd gnd FILL
XFILL_1__964_ vdd gnd FILL
X_1224_ _1327_/C _1325_/B _1410_/A vdd gnd NOR2X1
X_1155_ _980_/B _977_/B _1181_/C vdd gnd NAND2X1
X_1086_ _1209_/A _1209_/B _1236_/C _1114_/A vdd gnd NAND3X1
XFILL_1__1271_ vdd gnd FILL
XFILL_1__1340_ vdd gnd FILL
XFILL_0__1429_ vdd gnd FILL
XFILL_1__1607_ vdd gnd FILL
XFILL_1__1538_ vdd gnd FILL
XFILL_1__1469_ vdd gnd FILL
XFILL_0__982_ vdd gnd FILL
X_935_ _935_/A _935_/B _935_/C _936_/A vdd gnd OAI21X1
XFILL_0__1780_ vdd gnd FILL
XFILL_0__1145_ vdd gnd FILL
XFILL_0__1214_ vdd gnd FILL
X_1773_ _1773_/A _1795_/B _1782_/B _1779_/A vdd gnd OAI21X1
X_1842_ _1843_/A _1843_/B _1842_/C _1843_/C vdd gnd OAI21X1
XFILL_0__1076_ vdd gnd FILL
XFILL_1__947_ vdd gnd FILL
X_1207_ _1207_/A _1287_/B _1287_/A _1241_/B vdd gnd OAI21X1
X_1138_ _994_/A _998_/B _988_/C _1161_/A vdd gnd OAI21X1
XFILL_1__1323_ vdd gnd FILL
X_1069_ _1088_/C _1088_/B _1088_/A _1209_/A vdd gnd NAND3X1
XFILL_1__1254_ vdd gnd FILL
XFILL_1__1185_ vdd gnd FILL
XFILL_0_BUFX2_insert8 vdd gnd FILL
XFILL_2__1363_ vdd gnd FILL
XFILL_0__965_ vdd gnd FILL
XFILL_0__1832_ vdd gnd FILL
XFILL_0__1763_ vdd gnd FILL
XFILL_0__1694_ vdd gnd FILL
XFILL_0__1128_ vdd gnd FILL
X_1756_ _1756_/A _1756_/B _1780_/A _1757_/B vdd gnd OAI21X1
XFILL_0__1059_ vdd gnd FILL
X_1825_ _1843_/A _1826_/B _1842_/C _1826_/C vdd gnd OAI21X1
XFILL_1__1872_ vdd gnd FILL
X_1687_ _1687_/A _1842_/C _1836_/B _1709_/B vdd gnd OAI21X1
XFILL_1__1306_ vdd gnd FILL
XFILL_1__1168_ vdd gnd FILL
XFILL_1__1237_ vdd gnd FILL
XFILL_1__1099_ vdd gnd FILL
XFILL_0__948_ vdd gnd FILL
X_1610_ LoadCmd_i ABCmd_i[4] _1611_/C vdd gnd NAND2X1
X_1472_ _1519_/C _1524_/A _1472_/C _1479_/A vdd gnd NAND3X1
XFILL_0__1815_ vdd gnd FILL
X_1541_ _1594_/A _1817_/Y _1542_/A vdd gnd AND2X2
XFILL_0__1746_ vdd gnd FILL
XFILL_1__1022_ vdd gnd FILL
X_1739_ _1795_/C _1739_/Y vdd gnd INVX1
X_1808_ _1809_/A _977_/A _1842_/C _1809_/C vdd gnd OAI21X1
XFILL_1__1855_ vdd gnd FILL
XFILL_1__1786_ vdd gnd FILL
XFILL_2__1200_ vdd gnd FILL
XFILL_0__1462_ vdd gnd FILL
XFILL_0__1531_ vdd gnd FILL
XFILL_0__1600_ vdd gnd FILL
XFILL_0__1393_ vdd gnd FILL
X_1524_ _1524_/A _1524_/B _1526_/B vdd gnd NOR2X1
X_1455_ _1455_/A _1457_/C vdd gnd INVX1
X_1386_ _1442_/A _1444_/A vdd gnd INVX1
XFILL_1__1640_ vdd gnd FILL
XFILL_1__1571_ vdd gnd FILL
XFILL_0__1729_ vdd gnd FILL
XFILL_1__1005_ vdd gnd FILL
XFILL_1__1769_ vdd gnd FILL
XFILL_1__1838_ vdd gnd FILL
XFILL_1__980_ vdd gnd FILL
X_1171_ _1171_/A _1171_/B _1177_/C vdd gnd NAND2X1
X_1240_ _1341_/A _1248_/B _1248_/A _1352_/A vdd gnd NAND3X1
XFILL_0__1445_ vdd gnd FILL
XFILL_0__1514_ vdd gnd FILL
XFILL_0__1376_ vdd gnd FILL
X_1507_ _1510_/B _1510_/A _1508_/B vdd gnd AND2X2
XFILL_1__1554_ vdd gnd FILL
X_1438_ _1465_/A _1461_/A vdd gnd INVX1
X_1369_ _1369_/A _1369_/B _1369_/C _1435_/C vdd gnd AOI21X1
XFILL_1__1623_ vdd gnd FILL
XFILL86850x39750 vdd gnd FILL
XFILL86850x82950 vdd gnd FILL
XFILL_1__1485_ vdd gnd FILL
X_951_ _975_/B _953_/A vdd gnd INVX1
XFILL_0__1161_ vdd gnd FILL
XFILL_0__1092_ vdd gnd FILL
XFILL_0__1230_ vdd gnd FILL
X_1154_ _1156_/C _1156_/B _1156_/A _1180_/A vdd gnd NAND3X1
XFILL_1__963_ vdd gnd FILL
X_1223_ _975_/A _1881_/B _958_/B _1325_/B vdd gnd NAND3X1
X_1085_ _1085_/A _1085_/B _1209_/B vdd gnd NAND2X1
XFILL_0__1428_ vdd gnd FILL
XFILL_1__1270_ vdd gnd FILL
XFILL_0__1359_ vdd gnd FILL
XFILL86250x10950 vdd gnd FILL
XFILL86850x14550 vdd gnd FILL
XFILL_1__1537_ vdd gnd FILL
XFILL_1__1606_ vdd gnd FILL
XFILL_1__1399_ vdd gnd FILL
XFILL_1__1468_ vdd gnd FILL
XFILL_0__981_ vdd gnd FILL
X_934_ _962_/A _958_/B _935_/B vdd gnd NAND2X1
XFILL_2__1715_ vdd gnd FILL
XFILL_0__1144_ vdd gnd FILL
XFILL_0__1213_ vdd gnd FILL
X_1772_ _1774_/B _1782_/B vdd gnd INVX1
XFILL_0__1075_ vdd gnd FILL
X_1841_ _1841_/A _1841_/B _1841_/C _1878_/B vdd gnd OAI21X1
X_1137_ _1142_/C _1142_/B _1158_/A _1161_/C vdd gnd AOI21X1
XFILL_1__946_ vdd gnd FILL
X_1206_ _1206_/A _1206_/B _1287_/B vdd gnd AND2X2
XFILL_1__1322_ vdd gnd FILL
XFILL_1__1184_ vdd gnd FILL
X_1068_ _1221_/A _1228_/B _1228_/C _1088_/A vdd gnd NAND3X1
XFILL_1__1253_ vdd gnd FILL
XFILL_2__1500_ vdd gnd FILL
XFILL_0_BUFX2_insert9 vdd gnd FILL
XFILL_0__964_ vdd gnd FILL
XFILL_0__1831_ vdd gnd FILL
XFILL_0__1693_ vdd gnd FILL
XFILL_0__1762_ vdd gnd FILL
X_1686_ _1686_/A _1842_/C vdd gnd INVX4
X_1755_ _1878_/A _1756_/B _1756_/A _1780_/A vdd gnd OAI21X1
XFILL_0__1058_ vdd gnd FILL
X_1824_ _1863_/B _1824_/B _1824_/C _1824_/D _1828_/A vdd gnd OAI22X1
XFILL_0__1127_ vdd gnd FILL
XFILL_1__929_ vdd gnd FILL
XFILL_1__1871_ vdd gnd FILL
XFILL_1__1305_ vdd gnd FILL
XFILL86550x36150 vdd gnd FILL
XFILL_1__1167_ vdd gnd FILL
XFILL_1__1098_ vdd gnd FILL
XFILL_1__1236_ vdd gnd FILL
XFILL_0__947_ vdd gnd FILL
X_1540_ Flag_i MulL_i _1594_/A vdd gnd NOR2X1
X_1471_ _1471_/A _1525_/A _1524_/A vdd gnd NAND2X1
XFILL_0__1814_ vdd gnd FILL
XFILL_0__1745_ vdd gnd FILL
XFILL_1__1021_ vdd gnd FILL
X_1807_ _1807_/A _1807_/B _1807_/C _1811_/A vdd gnd OAI21X1
X_1669_ _1669_/D _1681_/CLK _975_/B vdd gnd DFFPOSX1
XFILL_1__1854_ vdd gnd FILL
X_1738_ _1738_/A _1757_/C _1795_/C vdd gnd NAND2X1
XFILL_1__1785_ vdd gnd FILL
XFILL_1__1219_ vdd gnd FILL
XFILL_0__1461_ vdd gnd FILL
XFILL_0__1530_ vdd gnd FILL
XFILL_0__1392_ vdd gnd FILL
XFILL_2__1259_ vdd gnd FILL
X_1454_ _1455_/A _1454_/B _1456_/A _1463_/A vdd gnd OAI21X1
X_1523_ _1523_/A _1523_/B _1523_/C _1525_/D vdd gnd OAI21X1
X_1385_ _923_/A _962_/B _977_/A _1442_/A vdd gnd NAND3X1
XFILL_0__1728_ vdd gnd FILL
XFILL_1__1570_ vdd gnd FILL
XFILL_1__1004_ vdd gnd FILL
XFILL_1__1837_ vdd gnd FILL
XFILL_1__1768_ vdd gnd FILL
XFILL_1__1699_ vdd gnd FILL
X_1170_ _1180_/A _1170_/B _1170_/C _1480_/A vdd gnd NAND3X1
XFILL_0__1513_ vdd gnd FILL
XFILL_0__1444_ vdd gnd FILL
XFILL_0__1375_ vdd gnd FILL
X_1506_ _1510_/A _1510_/B _1543_/C vdd gnd NOR2X1
X_1437_ _1437_/A _1437_/B _1437_/C _1465_/A vdd gnd OAI21X1
X_1368_ _1436_/A _1469_/A vdd gnd INVX1
XFILL_1__1553_ vdd gnd FILL
X_1299_ _1299_/A _1299_/B _1367_/C _1332_/B vdd gnd NAND3X1
XFILL_1__1622_ vdd gnd FILL
XFILL_1__1484_ vdd gnd FILL
X_950_ _955_/B _955_/C _955_/A _956_/C vdd gnd NAND3X1
XFILL_2__1800_ vdd gnd FILL
XFILL_0__1160_ vdd gnd FILL
XFILL_0__1091_ vdd gnd FILL
XFILL_1__962_ vdd gnd FILL
X_1153_ _931_/A _937_/B _937_/A _1156_/B vdd gnd OAI21X1
X_1222_ _962_/A _1823_/A _964_/B _1327_/C vdd gnd NAND3X1
X_1084_ _1084_/A _1201_/C _1089_/C _1085_/A vdd gnd NAND3X1
XFILL_0__1427_ vdd gnd FILL
XFILL_0__1358_ vdd gnd FILL
XFILL_0__1289_ vdd gnd FILL
XFILL_1__1467_ vdd gnd FILL
XFILL_1__1605_ vdd gnd FILL
XFILL_1__1536_ vdd gnd FILL
XFILL_2__927_ vdd gnd FILL
XFILL_1__1398_ vdd gnd FILL
XFILL_0__980_ vdd gnd FILL
X_933_ _980_/C _935_/A vdd gnd INVX2
XFILL_0__1212_ vdd gnd FILL
X_1840_ _1881_/B _1840_/B _1863_/B _1841_/A vdd gnd OAI21X1
XFILL_0__1143_ vdd gnd FILL
X_1771_ _1771_/A _1771_/B _1781_/A _1774_/B vdd gnd OAI21X1
XFILL_0__1074_ vdd gnd FILL
XFILL_1__945_ vdd gnd FILL
X_1136_ _1136_/A _1136_/B _1136_/C _1142_/B vdd gnd NAND3X1
XFILL_1__1321_ vdd gnd FILL
X_1067_ _946_/A _1548_/B _1067_/C _1221_/A vdd gnd OAI21X1
X_1205_ _1206_/B _1206_/A _1207_/A vdd gnd NOR2X1
XFILL_1__1183_ vdd gnd FILL
XFILL_1__1252_ vdd gnd FILL
XFILL_1__1519_ vdd gnd FILL
XFILL_0__963_ vdd gnd FILL
XFILL_0__1830_ vdd gnd FILL
XFILL_0__1761_ vdd gnd FILL
XFILL_2__1559_ vdd gnd FILL
XFILL_0__1692_ vdd gnd FILL
X_1823_ _1823_/A _1823_/B _1863_/B _1824_/C vdd gnd OAI21X1
X_1754_ _1794_/A _1794_/B _1780_/B vdd gnd NAND2X1
XFILL_1__1870_ vdd gnd FILL
XFILL_0__1057_ vdd gnd FILL
X_1685_ _1750_/A _1687_/A vdd gnd INVX1
XFILL_0__1126_ vdd gnd FILL
XFILL_1__928_ vdd gnd FILL
XFILL_1__1304_ vdd gnd FILL
X_1119_ _1246_/A _1246_/B _1195_/C _1123_/B vdd gnd NAND3X1
XFILL_1__1235_ vdd gnd FILL
XFILL_1__1097_ vdd gnd FILL
XFILL_1__1166_ vdd gnd FILL
XFILL_2__1344_ vdd gnd FILL
XFILL85950x39750 vdd gnd FILL
XFILL85950x82950 vdd gnd FILL
XFILL_0__946_ vdd gnd FILL
X_1470_ _1470_/A _1488_/C _1470_/C _1471_/A vdd gnd NAND3X1
XFILL_0__1813_ vdd gnd FILL
XFILL_0__1744_ vdd gnd FILL
XFILL_0__1109_ vdd gnd FILL
XFILL_1__1020_ vdd gnd FILL
X_1806_ _962_/B _1806_/B _1863_/B _1807_/A vdd gnd OAI21X1
X_1599_ LoadCmd_i _1599_/B _1599_/C _1653_/D vdd gnd OAI21X1
XFILL_1__1853_ vdd gnd FILL
X_1737_ _1741_/B _1737_/B _1738_/A vdd gnd NAND2X1
X_1668_ _1668_/R vdd _1668_/D _1668_/CLK _1897_/A vdd gnd DFFSR
XFILL_1__1784_ vdd gnd FILL
XFILL_1__1218_ vdd gnd FILL
XFILL_1__1149_ vdd gnd FILL
XFILL_0__1460_ vdd gnd FILL
XFILL_0__1391_ vdd gnd FILL
XFILL_0__929_ vdd gnd FILL
X_1453_ _1453_/A _1545_/B _1456_/A vdd gnd NAND2X1
X_1522_ _1522_/A _1584_/A _1584_/C _1560_/C vdd gnd NAND3X1
XFILL_0__1727_ vdd gnd FILL
X_1384_ _1406_/A _1406_/B _1462_/B vdd gnd NAND2X1
XFILL_0__1589_ vdd gnd FILL
XFILL_1__1003_ vdd gnd FILL
XFILL_1__1836_ vdd gnd FILL
XFILL_1__1767_ vdd gnd FILL
XFILL_1__1698_ vdd gnd FILL
XFILL_2__1043_ vdd gnd FILL
XFILL_0__1512_ vdd gnd FILL
XFILL_0__1443_ vdd gnd FILL
XFILL_0__1374_ vdd gnd FILL
X_1436_ _1436_/A _1436_/B _1436_/C _1519_/A vdd gnd AOI21X1
X_1505_ _1576_/A _1505_/B _1510_/B vdd gnd NAND2X1
X_1367_ _1367_/A _1367_/B _1367_/C _1436_/A vdd gnd OAI21X1
XFILL_1__1621_ vdd gnd FILL
XFILL_1__1552_ vdd gnd FILL
X_1298_ _1627_/B _1548_/D _1302_/A _1299_/B vdd gnd OAI21X1
XFILL_1__1483_ vdd gnd FILL
XFILL_1__1819_ vdd gnd FILL
XFILL_2__1592_ vdd gnd FILL
XFILL_0__1090_ vdd gnd FILL
XFILL_1__961_ vdd gnd FILL
X_1221_ _1221_/A _1221_/B _1221_/C _1233_/C vdd gnd AOI21X1
XFILL_2__1859_ vdd gnd FILL
X_1152_ _1172_/B _1152_/B _1171_/B _1156_/C vdd gnd OAI21X1
X_1083_ _1201_/A _1201_/B _1089_/C vdd gnd NAND2X1
XFILL_0__1426_ vdd gnd FILL
XFILL_0__1288_ vdd gnd FILL
XFILL_0__1357_ vdd gnd FILL
X_1419_ _1419_/A _1419_/B _1419_/C _1420_/B vdd gnd AOI21X1
XFILL_1__1604_ vdd gnd FILL
XFILL_1__1466_ vdd gnd FILL
XFILL_1__1397_ vdd gnd FILL
XFILL86550x64950 vdd gnd FILL
XFILL_1__1535_ vdd gnd FILL
X_932_ _980_/A _964_/B _979_/C _937_/A vdd gnd NAND3X1
XFILL_2__1644_ vdd gnd FILL
XFILL_0__1142_ vdd gnd FILL
XFILL_0__1211_ vdd gnd FILL
X_1770_ _1878_/A _1771_/B _1771_/A _1781_/A vdd gnd OAI21X1
XFILL_0__1073_ vdd gnd FILL
XFILL_1__944_ vdd gnd FILL
X_1204_ _1204_/A _1204_/B _1287_/C _1241_/A vdd gnd NAND3X1
X_1135_ _1185_/C _1135_/B _1142_/C vdd gnd NOR2X1
XFILL_1__1320_ vdd gnd FILL
XFILL_1__1251_ vdd gnd FILL
X_1066_ _975_/A _1823_/A _1548_/B vdd gnd NAND2X1
XFILL_0__1409_ vdd gnd FILL
XFILL_1__1182_ vdd gnd FILL
XFILL_1__1518_ vdd gnd FILL
XFILL_1__1449_ vdd gnd FILL
XFILL_2__1291_ vdd gnd FILL
XFILL_0__962_ vdd gnd FILL
XFILL_0__1760_ vdd gnd FILL
XFILL_0__1691_ vdd gnd FILL
X_1753_ _1753_/A _1753_/B _1756_/A _1794_/A vdd gnd MUX2X1
X_1822_ _1839_/A _1826_/B _1822_/C _1839_/D _1824_/D vdd gnd AOI22X1
XFILL_0__1125_ vdd gnd FILL
X_1684_ _1684_/D _1684_/CLK _1843_/B vdd gnd DFFPOSX1
XFILL_0__1056_ vdd gnd FILL
XFILL_1__927_ vdd gnd FILL
XFILL_0__1889_ vdd gnd FILL
XFILL_1__1303_ vdd gnd FILL
X_1049_ _1049_/A _1049_/B _998_/Y _1118_/C vdd gnd NAND3X1
X_1118_ _1118_/A _1118_/B _1118_/C _1123_/C vdd gnd OAI21X1
XFILL_1__1234_ vdd gnd FILL
XFILL_1__1096_ vdd gnd FILL
XFILL_1__1165_ vdd gnd FILL
XFILL_0__945_ vdd gnd FILL
XFILL_0__1812_ vdd gnd FILL
XFILL_0__1743_ vdd gnd FILL
XFILL_0__1039_ vdd gnd FILL
X_1736_ _1740_/B _1740_/A _1757_/A _1737_/B vdd gnd OAI21X1
XFILL_0__1108_ vdd gnd FILL
X_1805_ _1839_/A _977_/A _1805_/C _1839_/D _1807_/B vdd gnd AOI22X1
X_1598_ ABCmd_i[0] LoadCmd_i _1599_/C vdd gnd NAND2X1
XFILL_1__1852_ vdd gnd FILL
XFILL86250x18150 vdd gnd FILL
XFILL_1__1783_ vdd gnd FILL
X_1667_ _1668_/R vdd _1667_/D _1668_/CLK _1896_/A vdd gnd DFFSR
XFILL_1__1148_ vdd gnd FILL
XFILL_1__1217_ vdd gnd FILL
XFILL_1__1079_ vdd gnd FILL
XFILL_2__1892_ vdd gnd FILL
XFILL_0__1390_ vdd gnd FILL
XFILL_0__928_ vdd gnd FILL
X_1383_ _1383_/A _1437_/B _1437_/A _1406_/B vdd gnd OAI21X1
X_1452_ _1635_/B _982_/B _1495_/A _1453_/A vdd gnd OAI21X1
X_1521_ _1521_/A _1521_/B _1521_/C _1584_/C vdd gnd OAI21X1
XFILL_0__1726_ vdd gnd FILL
XFILL_1__1002_ vdd gnd FILL
XFILL_0__1588_ vdd gnd FILL
X_1719_ _979_/C _1719_/B _1863_/B _1720_/B vdd gnd OAI21X1
XFILL_1__1835_ vdd gnd FILL
XFILL_1__1766_ vdd gnd FILL
XFILL_1__1697_ vdd gnd FILL
XFILL_0__1511_ vdd gnd FILL
XFILL_0__1442_ vdd gnd FILL
XFILL_0__1373_ vdd gnd FILL
X_1504_ _1504_/A _1504_/B _1504_/C _1576_/A vdd gnd NAND3X1
X_1435_ _1435_/A _1460_/B _1435_/C _1436_/C vdd gnd NOR3X1
XFILL_1__1551_ vdd gnd FILL
X_1366_ _1521_/A _1521_/B _1476_/B _1425_/A vdd gnd OAI21X1
XFILL_1__1620_ vdd gnd FILL
X_1297_ _1297_/A _1297_/B _1297_/C _1302_/A vdd gnd AOI21X1
XFILL_0__1709_ vdd gnd FILL
XFILL_1__1482_ vdd gnd FILL
XFILL_1__1818_ vdd gnd FILL
XFILL_1__1749_ vdd gnd FILL
XFILL_1__960_ vdd gnd FILL
X_1151_ _1171_/A _1152_/B vdd gnd INVX1
X_1220_ _1237_/A _1237_/B _1329_/A vdd gnd NAND2X1
XFILL_0__1425_ vdd gnd FILL
X_1082_ _1218_/C _1201_/B vdd gnd INVX1
XFILL_0__1356_ vdd gnd FILL
XFILL_0__1287_ vdd gnd FILL
X_1418_ _1420_/C _1418_/B _1418_/C _1517_/B vdd gnd NAND3X1
X_1349_ _1349_/A _1349_/B _1349_/C _1354_/C vdd gnd OAI21X1
XFILL_1__1534_ vdd gnd FILL
XFILL_1__1603_ vdd gnd FILL
XFILL_1__1465_ vdd gnd FILL
XFILL_1__1396_ vdd gnd FILL
X_931_ _931_/A _937_/C vdd gnd INVX1
XFILL_0__1141_ vdd gnd FILL
XFILL_0__1210_ vdd gnd FILL
XFILL_0__1072_ vdd gnd FILL
X_1134_ _953_/C _927_/B _1135_/B vdd gnd AND2X2
XFILL_1__943_ vdd gnd FILL
X_1203_ _935_/A _1548_/D _1206_/A _1204_/B vdd gnd OAI21X1
XFILL_0__1408_ vdd gnd FILL
XFILL_1__1181_ vdd gnd FILL
X_1065_ _1065_/A _1067_/C _1228_/C vdd gnd OR2X2
XFILL_1__1250_ vdd gnd FILL
XFILL_0__1339_ vdd gnd FILL
XFILL_1__1517_ vdd gnd FILL
XFILL_1__1448_ vdd gnd FILL
XFILL_1__1379_ vdd gnd FILL
XFILL_0__961_ vdd gnd FILL
XFILL_0__1690_ vdd gnd FILL
X_1683_ _1683_/D _1683_/CLK _1826_/B vdd gnd DFFPOSX1
X_1752_ _1752_/A _1842_/C _1753_/B _1753_/A vdd gnd OAI21X1
XFILL_0__1055_ vdd gnd FILL
XFILL_0__1124_ vdd gnd FILL
X_1821_ _1823_/A _1823_/B _1822_/C vdd gnd NAND2X1
XFILL_1__926_ vdd gnd FILL
XFILL_0__1888_ vdd gnd FILL
X_1117_ _1124_/B _1124_/A _1124_/C _1192_/A vdd gnd NAND3X1
XFILL_1__1302_ vdd gnd FILL
XFILL_1__1164_ vdd gnd FILL
X_1048_ _1048_/A _1048_/B _1048_/C _1055_/B vdd gnd NAND3X1
XFILL_1__1233_ vdd gnd FILL
XFILL_1__1095_ vdd gnd FILL
XFILL_0__944_ vdd gnd FILL
XFILL_0__1811_ vdd gnd FILL
XFILL_0__1742_ vdd gnd FILL
X_1735_ _1878_/A _1740_/A _1740_/B _1757_/A vdd gnd OAI21X1
XFILL_0__1107_ vdd gnd FILL
X_1804_ _962_/B _1806_/B _1805_/C vdd gnd NAND2X1
XFILL_0__1038_ vdd gnd FILL
X_1666_ _1668_/R vdd _1666_/D _1679_/CLK _1895_/A vdd gnd DFFSR
XFILL_1__1782_ vdd gnd FILL
XFILL_1__1851_ vdd gnd FILL
X_1597_ _1744_/A _1599_/B vdd gnd INVX1
XFILL_1__1147_ vdd gnd FILL
XFILL_1__1216_ vdd gnd FILL
XFILL_1__1078_ vdd gnd FILL
XFILL_2__1187_ vdd gnd FILL
XFILL_0__927_ vdd gnd FILL
X_1520_ _1525_/A _1525_/B _1520_/C _1520_/D _1521_/C vdd gnd AOI22X1
X_1382_ _1382_/A _1382_/B _1437_/B vdd gnd AND2X2
X_1451_ _1495_/A _1495_/B _1545_/B vdd gnd OR2X2
XFILL_0__1725_ vdd gnd FILL
XFILL_0__1587_ vdd gnd FILL
XFILL_1__1001_ vdd gnd FILL
X_1649_ ABCmd_i[6] LoadB_i _1650_/C vdd gnd NAND2X1
XFILL_1__1834_ vdd gnd FILL
X_1718_ _1744_/A _1718_/B _1719_/B vdd gnd NOR2X1
XFILL_1__1696_ vdd gnd FILL
XFILL_1__1765_ vdd gnd FILL
XFILL_0__1441_ vdd gnd FILL
XFILL_0__1510_ vdd gnd FILL
XFILL_0__1372_ vdd gnd FILL
XFILL_2__1239_ vdd gnd FILL
X_1503_ _1551_/A _1504_/B vdd gnd INVX1
XFILL_1__1550_ vdd gnd FILL
X_1365_ _1520_/D _1520_/C _1476_/B vdd gnd NAND2X1
X_1296_ _964_/C _1627_/B vdd gnd INVX1
XFILL_0__1708_ vdd gnd FILL
X_1434_ _920_/Y _1434_/B _1434_/C _1663_/D vdd gnd OAI21X1
XFILL_0__1639_ vdd gnd FILL
XFILL_1__1481_ vdd gnd FILL
XFILL_1__1817_ vdd gnd FILL
XFILL_1__1748_ vdd gnd FILL
XFILL_2__1024_ vdd gnd FILL
X_1150_ _982_/A _935_/B _1150_/C _1171_/A vdd gnd OAI21X1
XFILL_0__1424_ vdd gnd FILL
XFILL_0__1355_ vdd gnd FILL
X_1081_ _1201_/D _1091_/C _1085_/B vdd gnd NAND2X1
XFILL_0__1286_ vdd gnd FILL
X_1417_ _1421_/A _1421_/B _1418_/C vdd gnd NAND2X1
XFILL_1__1464_ vdd gnd FILL
XFILL_1__1602_ vdd gnd FILL
X_1348_ _1419_/B _1419_/A _1419_/C _1420_/C vdd gnd NAND3X1
XFILL_1__1533_ vdd gnd FILL
X_1279_ _1279_/A _1279_/B _1280_/B vdd gnd AND2X2
XFILL_1__1395_ vdd gnd FILL
X_930_ _935_/C _930_/B _931_/A vdd gnd NOR2X1
XFILL_0__1140_ vdd gnd FILL
XFILL_0__1071_ vdd gnd FILL
XFILL_1__942_ vdd gnd FILL
X_1133_ _1136_/C _1136_/B _1136_/A _1158_/A vdd gnd AOI21X1
X_1064_ _1221_/C _1228_/A _1221_/B _1088_/B vdd gnd OAI21X1
XFILL86850x150 vdd gnd FILL
X_1202_ _1206_/A _1206_/B _1287_/C vdd gnd OR2X2
XFILL_0__1407_ vdd gnd FILL
XFILL_1__1180_ vdd gnd FILL
XFILL_0__1338_ vdd gnd FILL
XFILL_0__1269_ vdd gnd FILL
X_1897_ _1897_/A ACC_o[7] vdd gnd BUFX2
XFILL86250x46950 vdd gnd FILL
XFILL_1__1447_ vdd gnd FILL
XFILL_1__1516_ vdd gnd FILL
XFILL_1__1378_ vdd gnd FILL
XFILL_0__960_ vdd gnd FILL
XFILL_2__1625_ vdd gnd FILL
X_1820_ _1837_/A _1826_/B _1823_/B vdd gnd AND2X2
XFILL_2__1487_ vdd gnd FILL
X_1682_ _1682_/D _1683_/CLK _977_/A vdd gnd DFFPOSX1
X_1751_ _1756_/B _1753_/B vdd gnd INVX1
XFILL_0__1123_ vdd gnd FILL
XFILL_0__1054_ vdd gnd FILL
XFILL_1__925_ vdd gnd FILL
XFILL_0__1887_ vdd gnd FILL
XFILL_1__1301_ vdd gnd FILL
X_1047_ _1055_/C _1118_/B _1055_/A _1166_/A vdd gnd OAI21X1
X_1116_ _1246_/B _1195_/C _1195_/A _1124_/B vdd gnd NAND3X1
XFILL_1__1163_ vdd gnd FILL
XFILL_1__1094_ vdd gnd FILL
XFILL86850x25350 vdd gnd FILL
XFILL_1__1232_ vdd gnd FILL
XFILL_2__1272_ vdd gnd FILL
XFILL_0__943_ vdd gnd FILL
XFILL_0__1741_ vdd gnd FILL
XFILL_0__1810_ vdd gnd FILL
X_1803_ _1837_/A _977_/A _1806_/B vdd gnd AND2X2
XFILL_0__1037_ vdd gnd FILL
X_1734_ _1734_/A _1734_/B _1734_/C _1734_/D _1741_/B vdd gnd AOI22X1
XFILL_1__1850_ vdd gnd FILL
XFILL_0__1106_ vdd gnd FILL
X_1665_ _1668_/R vdd _1665_/D _1668_/CLK _1894_/A vdd gnd DFFSR
X_1596_ reset _1668_/R vdd gnd INVX4
XFILL_1__1781_ vdd gnd FILL
XFILL_1__1215_ vdd gnd FILL
XFILL_1__1077_ vdd gnd FILL
XFILL_1__1146_ vdd gnd FILL
XFILL_2__1324_ vdd gnd FILL
XFILL_0__926_ vdd gnd FILL
X_1450_ _1881_/B _922_/B _1495_/B vdd gnd NAND2X1
XFILL_0__1724_ vdd gnd FILL
X_1381_ _1382_/B _1382_/A _1383_/A vdd gnd NOR2X1
XFILL_0__1586_ vdd gnd FILL
XFILL_1__1000_ vdd gnd FILL
X_1648_ LoadB_i _1648_/B _1648_/C _1682_/D vdd gnd OAI21X1
X_1579_ _1579_/A _1579_/B _1589_/C vdd gnd NAND2X1
XFILL_1__1833_ vdd gnd FILL
X_1717_ _958_/B _1718_/B vdd gnd INVX1
XFILL_1__1695_ vdd gnd FILL
XFILL_1__1764_ vdd gnd FILL
XFILL_1__1129_ vdd gnd FILL
XFILL_0__1440_ vdd gnd FILL
XFILL_0__1371_ vdd gnd FILL
X_1502_ _1881_/B _1502_/B _1551_/A vdd gnd NAND2X1
X_1433_ _920_/Y _1433_/B _1434_/C vdd gnd NAND2X1
X_1295_ _1370_/B _1577_/B _1295_/C _1367_/C vdd gnd NAND3X1
XFILL_1__1480_ vdd gnd FILL
X_1364_ _1523_/C _1523_/A _1520_/C vdd gnd NAND2X1
XFILL_0__1707_ vdd gnd FILL
XFILL_2__940_ vdd gnd FILL
XFILL_0__1638_ vdd gnd FILL
XFILL_0__1569_ vdd gnd FILL
XFILL_1__1816_ vdd gnd FILL
XFILL_1__1747_ vdd gnd FILL
X_1080_ _1080_/A _1218_/C _1201_/C _1091_/C vdd gnd OAI21X1
XFILL_2__1787_ vdd gnd FILL
XFILL_0__1423_ vdd gnd FILL
XFILL_0__1354_ vdd gnd FILL
XFILL_0__1285_ vdd gnd FILL
XFILL_1__1601_ vdd gnd FILL
X_1416_ _1436_/A _1469_/C _1436_/B _1421_/B vdd gnd NAND3X1
X_1347_ _1355_/C _1355_/B _1420_/A _1351_/A vdd gnd AOI21X1
XFILL_1__1463_ vdd gnd FILL
XFILL_1__1394_ vdd gnd FILL
XFILL_1__1532_ vdd gnd FILL
X_1278_ _920_/Y _1278_/B _1278_/C _1661_/D vdd gnd OAI21X1
XFILL_2__1572_ vdd gnd FILL
XFILL_0__1070_ vdd gnd FILL
XFILL_1__941_ vdd gnd FILL
X_1201_ _1201_/A _1201_/B _1201_/C _1201_/D _1206_/A vdd gnd AOI22X1
XFILL_2__1839_ vdd gnd FILL
X_1132_ _957_/A _971_/B _957_/C _1136_/C vdd gnd NAND3X1
X_989_ _989_/A _989_/B _989_/C _994_/A vdd gnd AOI21X1
X_1063_ _1228_/B _1221_/B vdd gnd INVX1
XFILL_0__1406_ vdd gnd FILL
XFILL_0__1337_ vdd gnd FILL
XFILL_0__1268_ vdd gnd FILL
X_1896_ _1896_/A ACC_o[6] vdd gnd BUFX2
XFILL_0__1199_ vdd gnd FILL
XFILL_1__1446_ vdd gnd FILL
XFILL_1__1377_ vdd gnd FILL
XFILL_1__1515_ vdd gnd FILL
X_1750_ _1750_/A _964_/B _1750_/C _1756_/B vdd gnd AOI21X1
XFILL_0__1122_ vdd gnd FILL
X_1681_ _1681_/D _1681_/CLK _979_/B vdd gnd DFFPOSX1
XFILL_0__1053_ vdd gnd FILL
XFILL_0__1886_ vdd gnd FILL
XFILL_1__924_ vdd gnd FILL
XFILL_1__1300_ vdd gnd FILL
XFILL_1__1231_ vdd gnd FILL
X_1046_ _1118_/A _1055_/A vdd gnd INVX1
X_1115_ _1115_/A _1115_/B _1195_/A vdd gnd AND2X2
XFILL_1__1162_ vdd gnd FILL
XFILL_1__1093_ vdd gnd FILL
X_1879_ _1879_/A _1879_/B _1881_/A vdd gnd NAND2X1
XFILL_0__942_ vdd gnd FILL
XFILL_1__1429_ vdd gnd FILL
XFILL_0__1740_ vdd gnd FILL
X_1733_ _1733_/A _1733_/B _1733_/C _1734_/C vdd gnd NAND3X1
X_1802_ _1836_/A _1823_/A _1807_/C vdd gnd NAND2X1
XFILL_0__1105_ vdd gnd FILL
XFILL_1__1780_ vdd gnd FILL
XFILL_0__1036_ vdd gnd FILL
X_1664_ _1668_/R vdd _1664_/D _1668_/CLK _1893_/A vdd gnd DFFSR
X_1595_ _1595_/A _1595_/B _1595_/C _1595_/D _1668_/D vdd gnd AOI22X1
XFILL_0__1869_ vdd gnd FILL
XFILL_1__1214_ vdd gnd FILL
X_1029_ _1029_/A _1029_/B _1029_/C _1056_/A vdd gnd AOI21X1
XFILL_1__1145_ vdd gnd FILL
XFILL_1__1076_ vdd gnd FILL
XFILL_0__925_ vdd gnd FILL
X_1380_ _1380_/A _1380_/B _1437_/C _1406_/A vdd gnd NAND3X1
XFILL_0__1723_ vdd gnd FILL
XFILL_0__1585_ vdd gnd FILL
X_1716_ _1839_/A _958_/B _1716_/C _1839_/D _1720_/A vdd gnd AOI22X1
X_1647_ ABCmd_i[5] LoadB_i _1648_/C vdd gnd NAND2X1
X_1578_ _1579_/B _1579_/A _1580_/B vdd gnd OR2X2
XFILL_1__1832_ vdd gnd FILL
XFILL_0__1019_ vdd gnd FILL
XFILL_1__1763_ vdd gnd FILL
XFILL_1__1694_ vdd gnd FILL
XFILL_1__1128_ vdd gnd FILL
XFILL_2__1872_ vdd gnd FILL
XFILL_1__1059_ vdd gnd FILL
XFILL_0__1370_ vdd gnd FILL
X_1501_ _1501_/A _1502_/B vdd gnd INVX1
X_1363_ _1363_/A _1363_/B _1521_/A vdd gnd NAND2X1
X_1432_ _1432_/A _1432_/B _1432_/C _1433_/B vdd gnd OAI21X1
XFILL_0__1637_ vdd gnd FILL
X_1294_ _1294_/A _1294_/B _1294_/C _1295_/C vdd gnd OAI21X1
XFILL_0__1706_ vdd gnd FILL
XFILL_0__1499_ vdd gnd FILL
XFILL_0__1568_ vdd gnd FILL
XFILL_1__1815_ vdd gnd FILL
XFILL_1__1746_ vdd gnd FILL
XFILL_2__999_ vdd gnd FILL
XFILL85950x25350 vdd gnd FILL
XFILL_0__1422_ vdd gnd FILL
XFILL_0__1284_ vdd gnd FILL
XFILL_0__1353_ vdd gnd FILL
X_1415_ _1435_/A _1460_/B _1435_/C _1436_/B vdd gnd OAI21X1
XFILL_1__1531_ vdd gnd FILL
X_1346_ _1349_/B _1349_/A _1419_/C _1355_/B vdd gnd OAI21X1
XFILL_1__1600_ vdd gnd FILL
XFILL_1__1462_ vdd gnd FILL
XFILL_1__1393_ vdd gnd FILL
X_1277_ _920_/Y _1277_/B _1278_/C vdd gnd NAND2X1
XFILL_1__1729_ vdd gnd FILL
X_988_ _988_/A _998_/C _988_/C _996_/B vdd gnd NAND3X1
XFILL_1__940_ vdd gnd FILL
X_1200_ _980_/C _1577_/B _1206_/B vdd gnd NAND2X1
X_1131_ _971_/C _957_/B _971_/A _1136_/B vdd gnd OAI21X1
XFILL_0__1405_ vdd gnd FILL
X_1062_ _1062_/A _964_/B _962_/B _1228_/B vdd gnd NAND3X1
XFILL_0__1336_ vdd gnd FILL
X_1895_ _1895_/A ACC_o[5] vdd gnd BUFX2
XFILL_0__1267_ vdd gnd FILL
XFILL_0__1198_ vdd gnd FILL
XFILL_1__1514_ vdd gnd FILL
X_1329_ _1329_/A _1329_/B _1329_/C _1330_/C vdd gnd OAI21X1
XFILL_1__1445_ vdd gnd FILL
XFILL_1__1376_ vdd gnd FILL
XFILL_0__1121_ vdd gnd FILL
XFILL_0__1052_ vdd gnd FILL
X_1680_ _1680_/D _1681_/CLK _980_/B vdd gnd DFFPOSX1
XFILL_1__923_ vdd gnd FILL
XFILL_0__1885_ vdd gnd FILL
X_1114_ _1114_/A _1114_/B _1114_/C _1195_/C vdd gnd NAND3X1
XFILL_1__1161_ vdd gnd FILL
X_1045_ _1045_/A _1256_/A _1118_/A vdd gnd NAND2X1
XFILL_1__1230_ vdd gnd FILL
XFILL_0__1319_ vdd gnd FILL
X_1878_ _1878_/A _1878_/B _1879_/B vdd gnd NAND2X1
XFILL_1__1092_ vdd gnd FILL
XFILL86550x75750 vdd gnd FILL
XFILL_0__941_ vdd gnd FILL
XFILL_1__1359_ vdd gnd FILL
XFILL_1__1428_ vdd gnd FILL
XFILL_2__1468_ vdd gnd FILL
XFILL_0__1035_ vdd gnd FILL
X_1801_ _1801_/A _1814_/C vdd gnd INVX1
X_1732_ _1863_/B _1732_/B _1732_/C _1733_/C vdd gnd NAND3X1
XFILL_0__1104_ vdd gnd FILL
X_1663_ _1668_/R vdd _1663_/D _1668_/CLK _1892_/A vdd gnd DFFSR
X_1594_ _1594_/A _1873_/A MulH_i _1595_/B vdd gnd AOI21X1
XFILL_0__1868_ vdd gnd FILL
XFILL_0__1799_ vdd gnd FILL
XFILL_1__1144_ vdd gnd FILL
XFILL_1__1213_ vdd gnd FILL
X_1028_ _1095_/B _1095_/A _1056_/C _1049_/A vdd gnd NAND3X1
XFILL86550x50550 vdd gnd FILL
XFILL_1__1075_ vdd gnd FILL
XFILL_0__924_ vdd gnd FILL
XFILL_0__1584_ vdd gnd FILL
XFILL_0__1722_ vdd gnd FILL
X_1646_ _977_/A _1648_/B vdd gnd INVX1
X_1715_ _979_/C _958_/B _1837_/A _1716_/C vdd gnd NAND3X1
XFILL_0__1018_ vdd gnd FILL
X_1577_ _1577_/A _1577_/B _1589_/B _1579_/A vdd gnd AOI21X1
XFILL_1__1831_ vdd gnd FILL
XFILL_1__1693_ vdd gnd FILL
XFILL_1__1762_ vdd gnd FILL
XFILL_1__1127_ vdd gnd FILL
XFILL_1__1058_ vdd gnd FILL
XFILL_2__1305_ vdd gnd FILL
XFILL_2__1167_ vdd gnd FILL
X_1500_ _1635_/B _1501_/A _1551_/B _1505_/B vdd gnd OAI21X1
X_1293_ _946_/B _1370_/B vdd gnd INVX1
X_1431_ _1856_/Y _1533_/B _1592_/C _1432_/B vdd gnd OAI21X1
X_1362_ _1362_/A _1362_/B _1362_/C _1662_/D vdd gnd OAI21X1
XFILL_0__1636_ vdd gnd FILL
XFILL_0__1567_ vdd gnd FILL
XFILL_0__1705_ vdd gnd FILL
XFILL_0__1498_ vdd gnd FILL
X_1629_ LoadA_i _1629_/B _1629_/C _1673_/D vdd gnd OAI21X1
XFILL_1__1814_ vdd gnd FILL
XFILL_1__1745_ vdd gnd FILL
XFILL_0__1421_ vdd gnd FILL
XFILL_0__1352_ vdd gnd FILL
XFILL_0__1283_ vdd gnd FILL
XFILL_0_CLKBUF1_insert0 vdd gnd FILL
X_1414_ _1468_/A _1468_/B _1468_/C _1469_/C vdd gnd NAND3X1
XFILL_1__1530_ vdd gnd FILL
X_1345_ _1345_/A _1345_/B _1405_/A _1349_/B vdd gnd AOI21X1
X_1276_ _1276_/A _1276_/B _1276_/C _1277_/B vdd gnd OAI21X1
XFILL_1__1461_ vdd gnd FILL
XFILL_0__1619_ vdd gnd FILL
XFILL_1__1392_ vdd gnd FILL
XFILL_1__1728_ vdd gnd FILL
XFILL_2__1004_ vdd gnd FILL
X_987_ _987_/A _987_/B _988_/C vdd gnd NAND2X1
X_1130_ _1143_/A _936_/A _931_/A _1136_/A vdd gnd AOI21X1
XFILL_2__1768_ vdd gnd FILL
XFILL_0__1404_ vdd gnd FILL
XFILL_0__1335_ vdd gnd FILL
X_1061_ _1065_/A _1067_/C _1228_/A vdd gnd AND2X2
XFILL_0__1197_ vdd gnd FILL
XFILL_0__1266_ vdd gnd FILL
X_1894_ _1894_/A ACC_o[4] vdd gnd BUFX2
XFILL_1__1513_ vdd gnd FILL
XFILL_1__1444_ vdd gnd FILL
XFILL_1__999_ vdd gnd FILL
X_1328_ _1408_/A _1328_/B _1333_/B _1329_/B vdd gnd AOI21X1
X_1259_ _1259_/A _1259_/B _1259_/C _1523_/A vdd gnd NAND3X1
XFILL_1__1375_ vdd gnd FILL
XFILL86250x7350 vdd gnd FILL
XFILL_2__1553_ vdd gnd FILL
XFILL_0__1120_ vdd gnd FILL
XFILL_0__1051_ vdd gnd FILL
XFILL_1__922_ vdd gnd FILL
XFILL_0__1884_ vdd gnd FILL
X_1113_ _1113_/A _1113_/B _1113_/C _1246_/B vdd gnd NAND3X1
X_1044_ _953_/A _1548_/D _1044_/C _1045_/A vdd gnd OAI21X1
XFILL_1__1160_ vdd gnd FILL
XFILL_0__1318_ vdd gnd FILL
XFILL_1__1091_ vdd gnd FILL
X_1877_ _1877_/A _1879_/A vdd gnd INVX1
XFILL_0__1249_ vdd gnd FILL
XFILL_1__1427_ vdd gnd FILL
XFILL_0__940_ vdd gnd FILL
XFILL_1__1289_ vdd gnd FILL
XFILL_1__1358_ vdd gnd FILL
XFILL_2__1605_ vdd gnd FILL
X_1800_ _1813_/B _1800_/B _1852_/B vdd gnd NOR2X1
XFILL_0__1034_ vdd gnd FILL
X_1731_ _1731_/A _1731_/B _1732_/C vdd gnd NAND2X1
XFILL_0__1103_ vdd gnd FILL
X_1662_ _1668_/R vdd _1662_/D _1668_/CLK _1891_/A vdd gnd DFFSR
XFILL_0__1867_ vdd gnd FILL
X_1593_ _1593_/A _1593_/B _1593_/C _1595_/A vdd gnd OAI21X1
X_1027_ _1031_/B _1031_/A _1095_/A vdd gnd NAND2X1
XFILL_0__1798_ vdd gnd FILL
XFILL_1__1143_ vdd gnd FILL
XFILL_1__1212_ vdd gnd FILL
XFILL_1__1074_ vdd gnd FILL
XFILL_2__1252_ vdd gnd FILL
XFILL_0__923_ vdd gnd FILL
XFILL_0__1721_ vdd gnd FILL
XFILL_0__1652_ vdd gnd FILL
XFILL_0__1583_ vdd gnd FILL
X_1576_ _1576_/A _1576_/B _1576_/C _1579_/B vdd gnd OAI21X1
X_1645_ LoadB_i _1645_/B _1645_/C _1681_/D vdd gnd OAI21X1
XFILL_1__1830_ vdd gnd FILL
XFILL_0__1017_ vdd gnd FILL
X_1714_ _1836_/A _980_/C _1720_/C vdd gnd NAND2X1
XFILL_1__1761_ vdd gnd FILL
XFILL_1__1692_ vdd gnd FILL
XFILL_1__1057_ vdd gnd FILL
XFILL_1__1126_ vdd gnd FILL
X_1430_ Flag_i _1759_/Y _1432_/A vdd gnd NOR2X1
X_1292_ _1367_/A _1299_/A vdd gnd INVX1
X_1361_ _1363_/B _1361_/B MulH_i _1362_/B vdd gnd OAI21X1
XFILL_0__1704_ vdd gnd FILL
XFILL_0__1635_ vdd gnd FILL
XFILL_0__1497_ vdd gnd FILL
XFILL_0__1566_ vdd gnd FILL
X_1628_ ABCmd_i[4] LoadA_i _1629_/C vdd gnd NAND2X1
X_1559_ _1563_/B _1575_/C _1583_/A vdd gnd NAND2X1
XFILL_1__1813_ vdd gnd FILL
XFILL_1__1744_ vdd gnd FILL
XFILL_1__1109_ vdd gnd FILL
XFILL_0__1420_ vdd gnd FILL
XFILL_0__1351_ vdd gnd FILL
XFILL_0__1282_ vdd gnd FILL
X_1413_ _1469_/A _1413_/B _1413_/C _1421_/A vdd gnd NAND3X1
XFILL86550x150 vdd gnd FILL
XFILL_0_CLKBUF1_insert1 vdd gnd FILL
XFILL_1__1460_ vdd gnd FILL
X_1344_ _1344_/A _1344_/B _1344_/C _1345_/B vdd gnd OAI21X1
X_1275_ _961_/A MulL_i _977_/B _1276_/C vdd gnd NAND3X1
XFILL_0__1618_ vdd gnd FILL
XFILL_1__1391_ vdd gnd FILL
XFILL_0__1549_ vdd gnd FILL
XFILL_2__920_ vdd gnd FILL
XFILL_1__1727_ vdd gnd FILL
XFILL_1__1589_ vdd gnd FILL
X_986_ _992_/C _991_/A _991_/B _987_/A vdd gnd NAND3X1
X_1060_ _1065_/A _1067_/C _1221_/C vdd gnd NOR2X1
XFILL_0__1403_ vdd gnd FILL
XFILL_0__1334_ vdd gnd FILL
XFILL_0__1196_ vdd gnd FILL
XFILL_0__1265_ vdd gnd FILL
X_1893_ _1893_/A ACC_o[3] vdd gnd BUFX2
XFILL_1__1512_ vdd gnd FILL
XFILL_1__1443_ vdd gnd FILL
XFILL_1__998_ vdd gnd FILL
X_1327_ _1635_/B _935_/B _1327_/C _1328_/B vdd gnd OAI21X1
X_1189_ _1569_/A _1568_/C vdd gnd INVX1
X_1258_ _1286_/A _1286_/B _1353_/C _1259_/B vdd gnd NAND3X1
XFILL_1__1374_ vdd gnd FILL
XFILL_0__1050_ vdd gnd FILL
XFILL_1__921_ vdd gnd FILL
XFILL_0__1883_ vdd gnd FILL
X_969_ _999_/C _972_/B _973_/B _990_/B vdd gnd OAI21X1
X_1112_ _1246_/C _1195_/B _1246_/A _1124_/A vdd gnd OAI21X1
X_1043_ _1577_/B _1548_/D vdd gnd INVX4
XFILL_0__1317_ vdd gnd FILL
XFILL_1__1090_ vdd gnd FILL
XFILL_0__1248_ vdd gnd FILL
X_1876_ _1876_/A _1876_/B _1884_/B vdd gnd AND2X2
XFILL86550x10950 vdd gnd FILL
XFILL_0__1179_ vdd gnd FILL
XFILL_1__1426_ vdd gnd FILL
XFILL_1__1357_ vdd gnd FILL
XFILL_1__1288_ vdd gnd FILL
XFILL_0__1102_ vdd gnd FILL
XFILL_0__999_ vdd gnd FILL
XFILL_0__1033_ vdd gnd FILL
X_1661_ _1668_/R vdd _1661_/D _1668_/CLK _1890_/A vdd gnd DFFSR
X_1730_ _1863_/A _1839_/A _961_/A _1731_/A vdd gnd OAI21X1
X_1592_ _1593_/A _1593_/B _1592_/C _1593_/C vdd gnd AOI21X1
XFILL_0__1866_ vdd gnd FILL
XFILL_1__1211_ vdd gnd FILL
X_1026_ _1026_/A _1101_/B _1026_/C _1031_/B vdd gnd NAND3X1
XFILL_0__1797_ vdd gnd FILL
XFILL_1__1142_ vdd gnd FILL
X_1859_ _1859_/A _1876_/B _1859_/C _1868_/A vdd gnd OAI21X1
XFILL_1__1073_ vdd gnd FILL
XFILL_1__1409_ vdd gnd FILL
XFILL_0__922_ vdd gnd FILL
XFILL_0__1651_ vdd gnd FILL
XFILL_2_BUFX2_insert8 vdd gnd FILL
XFILL_0__1720_ vdd gnd FILL
XFILL_0__1582_ vdd gnd FILL
X_1713_ _1713_/A _1713_/B _1713_/C _1726_/B vdd gnd OAI21X1
X_1575_ _1575_/A _1583_/A _1575_/C _1585_/A vdd gnd OAI21X1
X_1644_ ABCmd_i[4] LoadB_i _1645_/C vdd gnd NAND2X1
XFILL_1__1760_ vdd gnd FILL
XFILL_0__1016_ vdd gnd FILL
XFILL_0__1849_ vdd gnd FILL
XFILL_1__1691_ vdd gnd FILL
X_1009_ _1057_/A _1070_/A _1070_/C _1030_/A vdd gnd NAND3X1
XFILL86250x32550 vdd gnd FILL
XFILL86850x36150 vdd gnd FILL
XFILL_1__1056_ vdd gnd FILL
XFILL_1__1125_ vdd gnd FILL
XFILL_1__1889_ vdd gnd FILL
XFILL_2__1096_ vdd gnd FILL
X_1360_ _1520_/D _1523_/C _1363_/B vdd gnd AND2X2
XFILL_0__1634_ vdd gnd FILL
X_1291_ _980_/C _1547_/B _1367_/A vdd gnd NAND2X1
XFILL_0__1703_ vdd gnd FILL
XFILL_0__1496_ vdd gnd FILL
XFILL_0__1565_ vdd gnd FILL
X_1489_ _1514_/A _1513_/A vdd gnd INVX1
X_1558_ _1558_/A _1558_/B _1575_/C vdd gnd OR2X2
X_1627_ LoadA_i _1627_/B _1627_/C _1672_/D vdd gnd OAI21X1
XFILL_1__1812_ vdd gnd FILL
XFILL_1__1743_ vdd gnd FILL
XFILL_1__1108_ vdd gnd FILL
XFILL_1__1039_ vdd gnd FILL
XFILL_2__1852_ vdd gnd FILL
XFILL_0__1350_ vdd gnd FILL
XFILL_0__1281_ vdd gnd FILL
XFILL_0_CLKBUF1_insert2 vdd gnd FILL
XFILL_2__1148_ vdd gnd FILL
X_1412_ _1435_/A _1460_/B _1468_/C _1413_/B vdd gnd OAI21X1
X_1343_ _1343_/A _1343_/B _1345_/A vdd gnd NAND2X1
XFILL_1__1390_ vdd gnd FILL
XFILL_0__1617_ vdd gnd FILL
X_1274_ _1814_/A _1533_/B _1592_/C _1276_/B vdd gnd OAI21X1
XFILL_0__1548_ vdd gnd FILL
XFILL_0__1479_ vdd gnd FILL
XFILL_1__1726_ vdd gnd FILL
XFILL_1__1588_ vdd gnd FILL
XFILL_2__979_ vdd gnd FILL
X_985_ _992_/A _991_/B vdd gnd INVX1
XFILL_0__1402_ vdd gnd FILL
XFILL_0__1264_ vdd gnd FILL
X_1892_ _1892_/A ACC_o[2] vdd gnd BUFX2
XFILL_0__1333_ vdd gnd FILL
XFILL_0__1195_ vdd gnd FILL
XFILL_1__1511_ vdd gnd FILL
XFILL_1__997_ vdd gnd FILL
X_1326_ _1881_/B _1635_/B vdd gnd INVX2
XFILL_1__1442_ vdd gnd FILL
XFILL_1__1373_ vdd gnd FILL
X_1188_ _1529_/A _1567_/A _1537_/B _1569_/A vdd gnd NAND3X1
X_1257_ _1353_/A _1257_/B _1257_/C _1259_/A vdd gnd NAND3X1
XFILL_1__1709_ vdd gnd FILL
X_968_ _999_/A _972_/B vdd gnd INVX1
XFILL_0__1882_ vdd gnd FILL
XFILL_1__920_ vdd gnd FILL
X_1042_ _925_/A _1650_/B _1577_/B vdd gnd NOR2X1
X_1111_ _1115_/B _1115_/A _1246_/A vdd gnd NAND2X1
XFILL_0__1316_ vdd gnd FILL
X_1875_ _1876_/B _1876_/A _1884_/A vdd gnd NOR2X1
XFILL_0__1247_ vdd gnd FILL
XFILL_0__1178_ vdd gnd FILL
X_1309_ _1372_/A _1372_/B _1320_/C vdd gnd OR2X2
XFILL_1__1425_ vdd gnd FILL
XFILL_1__1356_ vdd gnd FILL
XFILL_1__1287_ vdd gnd FILL
XFILL_2__1396_ vdd gnd FILL
XFILL_0__998_ vdd gnd FILL
XFILL_0__1032_ vdd gnd FILL
XFILL_0__1101_ vdd gnd FILL
X_1660_ _1660_/D _1683_/CLK _1660_/Q vdd gnd DFFPOSX1
X_1591_ _1591_/A _1591_/B _1593_/A vdd gnd NOR2X1
XFILL_0__1865_ vdd gnd FILL
XFILL_0__1796_ vdd gnd FILL
XFILL_1__1141_ vdd gnd FILL
XFILL_1__1210_ vdd gnd FILL
X_1025_ _1025_/A _1201_/A _1026_/C vdd gnd NAND2X1
XFILL_1__1072_ vdd gnd FILL
X_1858_ _1858_/A _1858_/B _1870_/B vdd gnd NAND2X1
X_1789_ _1809_/A _979_/B _1842_/C _1790_/C vdd gnd OAI21X1
XFILL_1__1408_ vdd gnd FILL
XFILL_0__921_ vdd gnd FILL
XFILL_1__1339_ vdd gnd FILL
XFILL_0__1650_ vdd gnd FILL
XFILL_2__1448_ vdd gnd FILL
XFILL_0__1581_ vdd gnd FILL
X_1643_ LoadB_i _1643_/B _1643_/C _1680_/D vdd gnd OAI21X1
X_1712_ _1727_/A _1734_/A _1713_/B vdd gnd NOR2X1
XFILL_0__1015_ vdd gnd FILL
X_1574_ _1574_/A _1574_/B _1574_/C _1582_/B vdd gnd AOI21X1
XFILL_0__1779_ vdd gnd FILL
XFILL_0__1848_ vdd gnd FILL
XFILL_1__1690_ vdd gnd FILL
X_1008_ _946_/A _963_/B _1008_/C _1057_/A vdd gnd OAI21X1
XFILL_1__1124_ vdd gnd FILL
XFILL_1__1055_ vdd gnd FILL
XFILL_1__1888_ vdd gnd FILL
XFILL86850x7350 vdd gnd FILL
XFILL_2__1233_ vdd gnd FILL
XFILL_0__1633_ vdd gnd FILL
XFILL_0__1564_ vdd gnd FILL
XFILL_0__1702_ vdd gnd FILL
X_1290_ _1290_/A _1290_/B _1290_/C _1349_/C vdd gnd AOI21X1
XFILL_0__1495_ vdd gnd FILL
X_1626_ ABCmd_i[3] LoadA_i _1627_/C vdd gnd NAND2X1
X_1488_ _1488_/A _1488_/B _1488_/C _1514_/A vdd gnd OAI21X1
X_1557_ _1558_/B _1558_/A _1563_/B vdd gnd NAND2X1
XFILL_1__1811_ vdd gnd FILL
XFILL_1__1742_ vdd gnd FILL
XFILL_1__1107_ vdd gnd FILL
XFILL_1__1038_ vdd gnd FILL
XFILL_0__1280_ vdd gnd FILL
XFILL_0_CLKBUF1_insert3 vdd gnd FILL
X_1411_ _1411_/A _1411_/B _1462_/B _1460_/B vdd gnd AOI21X1
X_1342_ _1405_/C _1369_/B _1369_/A _1349_/A vdd gnd AOI21X1
X_1273_ MulL_i _1592_/C vdd gnd INVX2
XFILL_0__1616_ vdd gnd FILL
XFILL_0__1547_ vdd gnd FILL
XFILL_0__1478_ vdd gnd FILL
X_1609_ _1836_/B _1611_/B vdd gnd INVX1
XFILL_1__1725_ vdd gnd FILL
XFILL_1__1587_ vdd gnd FILL
X_984_ _992_/A _992_/B _991_/C _987_/B vdd gnd OAI21X1
XFILL_0__1401_ vdd gnd FILL
XFILL_2__1696_ vdd gnd FILL
XFILL_0__1332_ vdd gnd FILL
XFILL_0__1194_ vdd gnd FILL
X_1891_ _1891_/A ACC_o[1] vdd gnd BUFX2
XFILL_0__1263_ vdd gnd FILL
XFILL_1__1510_ vdd gnd FILL
XFILL_1__996_ vdd gnd FILL
X_1325_ _1327_/C _1325_/B _1408_/A vdd gnd OR2X2
X_1256_ _1256_/A _1256_/B _1256_/C _1259_/C vdd gnd OAI21X1
XFILL_1__1441_ vdd gnd FILL
X_1187_ _1187_/A _1187_/B _1187_/C _1537_/B vdd gnd NAND3X1
XFILL_1__1372_ vdd gnd FILL
XFILL_1__1639_ vdd gnd FILL
XFILL_1__1708_ vdd gnd FILL
XFILL_2__1481_ vdd gnd FILL
X_967_ _967_/A _967_/B _999_/C vdd gnd NOR2X1
XFILL_0__1881_ vdd gnd FILL
X_1110_ _1194_/A _1110_/B _1194_/C _1115_/B vdd gnd NAND3X1
XFILL_2__1748_ vdd gnd FILL
X_1041_ _1826_/B _1650_/B vdd gnd INVX1
XFILL_0__1315_ vdd gnd FILL
X_1874_ _1874_/A _1874_/B _1874_/C _1876_/A vdd gnd AOI21X1
XFILL_0__1246_ vdd gnd FILL
XFILL_0__1177_ vdd gnd FILL
XFILL_1__979_ vdd gnd FILL
X_1308_ _952_/A _1823_/A _980_/B _1372_/B vdd gnd NAND3X1
XFILL_1__1424_ vdd gnd FILL
X_1239_ _1289_/A _1344_/B _1340_/C _1248_/B vdd gnd OAI21X1
XFILL86850x64950 vdd gnd FILL
XFILL_1__1355_ vdd gnd FILL
XFILL_1__1286_ vdd gnd FILL
XFILL_2__1533_ vdd gnd FILL
XFILL_0__997_ vdd gnd FILL
XFILL_0__1031_ vdd gnd FILL
XFILL_0__1100_ vdd gnd FILL
X_1590_ _920_/Y _1590_/B _1595_/D vdd gnd NOR2X1
XFILL_0__1795_ vdd gnd FILL
XFILL_0__1864_ vdd gnd FILL
X_1024_ _1080_/A _1201_/A vdd gnd INVX1
XFILL_1__1140_ vdd gnd FILL
X_1857_ _1885_/B _1885_/C _1870_/A vdd gnd NAND2X1
XFILL_1__1071_ vdd gnd FILL
X_1788_ _1788_/A _1788_/B _1788_/C _1792_/A vdd gnd OAI21X1
XFILL_0__1229_ vdd gnd FILL
XFILL_1__1407_ vdd gnd FILL
XFILL_2__1180_ vdd gnd FILL
XFILL_1__1338_ vdd gnd FILL
XFILL_1__1269_ vdd gnd FILL
XFILL_0__920_ vdd gnd FILL
XFILL_0__1580_ vdd gnd FILL
X_1642_ ABCmd_i[3] LoadB_i _1643_/C vdd gnd NAND2X1
XFILL_0__1014_ vdd gnd FILL
X_1711_ _1711_/A _1850_/A vdd gnd INVX1
X_1573_ _1573_/A _1575_/A _1573_/C _1574_/C vdd gnd NAND3X1
XFILL_0__1847_ vdd gnd FILL
XFILL_0__1778_ vdd gnd FILL
X_1007_ _1007_/A _1008_/C _1070_/C vdd gnd OR2X2
XFILL_1__1123_ vdd gnd FILL
XFILL_1__1054_ vdd gnd FILL
XFILL_1__1887_ vdd gnd FILL
XFILL_0__1701_ vdd gnd FILL
XFILL_0__1632_ vdd gnd FILL
XFILL_0__1563_ vdd gnd FILL
XFILL_0__1494_ vdd gnd FILL
X_1556_ _1576_/C _1556_/B _1558_/A vdd gnd NAND2X1
X_1625_ LoadA_i _935_/A _1625_/C _1671_/D vdd gnd OAI21X1
XFILL_1__1810_ vdd gnd FILL
XFILL_1__1741_ vdd gnd FILL
XFILL86550x18150 vdd gnd FILL
X_1487_ _920_/Y _1487_/B _1487_/C _1664_/D vdd gnd OAI21X1
XFILL_1__1037_ vdd gnd FILL
XFILL_1__1106_ vdd gnd FILL
XFILL_2__1781_ vdd gnd FILL
X_1410_ _1410_/A _1410_/B _1410_/C _1411_/B vdd gnd OAI21X1
XFILL_0_CLKBUF1_insert4 vdd gnd FILL
X_1272_ Flag_i _1533_/B vdd gnd INVX1
X_1341_ _1341_/A _1341_/B _1341_/C _1419_/C vdd gnd OAI21X1
XFILL_0__1615_ vdd gnd FILL
XFILL_0__1546_ vdd gnd FILL
XFILL_0__1477_ vdd gnd FILL
X_1539_ _1539_/A _1539_/B _1539_/C _1542_/B vdd gnd AOI21X1
X_1608_ LoadCmd_i _1608_/B _1608_/C _1656_/D vdd gnd OAI21X1
XFILL_1__1724_ vdd gnd FILL
XFILL_1__1586_ vdd gnd FILL
X_983_ _991_/A _992_/B vdd gnd INVX1
XFILL_2__1833_ vdd gnd FILL
XFILL_0__1400_ vdd gnd FILL
XFILL_0__1331_ vdd gnd FILL
XFILL_0__1193_ vdd gnd FILL
X_1890_ _1890_/A ACC_o[0] vdd gnd BUFX2
XFILL_0__1262_ vdd gnd FILL
X_1186_ _997_/A _997_/C _1186_/C _1187_/B vdd gnd NAND3X1
XFILL_1__1440_ vdd gnd FILL
XFILL_1__995_ vdd gnd FILL
X_1324_ _1340_/B _1329_/C _1344_/C _1369_/C vdd gnd AOI21X1
X_1255_ _1255_/A _1255_/B _1255_/C _1268_/B vdd gnd OAI21X1
XFILL_1__1371_ vdd gnd FILL
XFILL_0__1529_ vdd gnd FILL
XFILL_1__1638_ vdd gnd FILL
XFILL_1__1569_ vdd gnd FILL
XFILL_1__1707_ vdd gnd FILL
XFILL_0__1880_ vdd gnd FILL
X_966_ _999_/A _999_/B _973_/C _990_/A vdd gnd NAND3X1
X_1040_ _1044_/C _1040_/B _1256_/A vdd gnd OR2X2
XFILL_0__1314_ vdd gnd FILL
XFILL_0__1176_ vdd gnd FILL
X_1873_ _1873_/A _1873_/B _1873_/C _1886_/C vdd gnd AOI21X1
XFILL_0__1245_ vdd gnd FILL
X_1307_ _923_/A _962_/B _979_/B _1372_/A vdd gnd NAND3X1
XFILL_1__978_ vdd gnd FILL
X_1169_ _1181_/A _1170_/C vdd gnd INVX1
XFILL_1__1423_ vdd gnd FILL
X_1238_ _1238_/A _1238_/B _1329_/A _1344_/B vdd gnd AOI21X1
XFILL_1__1354_ vdd gnd FILL
XFILL_1__1285_ vdd gnd FILL
XFILL_0__996_ vdd gnd FILL
XFILL_0__1030_ vdd gnd FILL
XFILL_0__1863_ vdd gnd FILL
X_949_ _971_/C _957_/B _957_/A _955_/B vdd gnd OAI21X1
XFILL_0__1794_ vdd gnd FILL
X_1023_ _1023_/A _1025_/A vdd gnd INVX1
XFILL_1__1070_ vdd gnd FILL
XFILL_0__1228_ vdd gnd FILL
XFILL_0__1159_ vdd gnd FILL
X_1856_ _1856_/A _1856_/B _1856_/Y vdd gnd AND2X2
X_1787_ _958_/C _1787_/B _1863_/B _1788_/A vdd gnd OAI21X1
XFILL_1__1406_ vdd gnd FILL
XFILL_1__1337_ vdd gnd FILL
XFILL_1__1199_ vdd gnd FILL
XFILL_1__1268_ vdd gnd FILL
XFILL_0__979_ vdd gnd FILL
X_1641_ LoadB_i _1641_/B _1641_/C _1679_/D vdd gnd OAI21X1
XFILL_0__1013_ vdd gnd FILL
X_1710_ _1710_/A _1710_/B _1711_/A vdd gnd NAND2X1
X_1572_ _920_/Y _1572_/B _1588_/A vdd gnd NAND2X1
XFILL_0__1846_ vdd gnd FILL
X_1006_ _1057_/C _1070_/B _1057_/B _1030_/B vdd gnd OAI21X1
XFILL_0__1777_ vdd gnd FILL
X_1839_ _1839_/A _1843_/B _1839_/C _1839_/D _1841_/B vdd gnd AOI22X1
XFILL_1__1122_ vdd gnd FILL
XFILL_1__1053_ vdd gnd FILL
XFILL_1__1886_ vdd gnd FILL
XFILL_0__1700_ vdd gnd FILL
XFILL_0__1631_ vdd gnd FILL
XFILL_0__1562_ vdd gnd FILL
XFILL_0__1493_ vdd gnd FILL
XFILL_2__1429_ vdd gnd FILL
XFILL86250x150 vdd gnd FILL
X_1555_ _1555_/A _1555_/B _1555_/C _1576_/C vdd gnd NAND3X1
X_1624_ ABCmd_i[2] LoadA_i _1625_/C vdd gnd NAND2X1
XFILL_1__1740_ vdd gnd FILL
XFILL_0__1829_ vdd gnd FILL
X_1486_ _1486_/A _1486_/B _920_/Y _1487_/C vdd gnd OAI21X1
XFILL_1__1036_ vdd gnd FILL
XFILL_1__1105_ vdd gnd FILL
XFILL_1__1869_ vdd gnd FILL
XFILL85950x64950 vdd gnd FILL
XFILL_2__1076_ vdd gnd FILL
X_1340_ _1340_/A _1340_/B _1340_/C _1341_/B vdd gnd AOI21X1
XFILL_0__1614_ vdd gnd FILL
X_1271_ _1850_/A Flag_i _1276_/A vdd gnd NOR2X1
XFILL_0__1545_ vdd gnd FILL
XFILL_0__1476_ vdd gnd FILL
X_1469_ _1469_/A _1469_/B _1469_/C _1470_/C vdd gnd OAI21X1
X_1607_ LoadCmd_i ABCmd_i[3] _1608_/C vdd gnd NAND2X1
X_1538_ _1539_/A _1539_/B MulL_i _1539_/C vdd gnd OAI21X1
XFILL_1__1723_ vdd gnd FILL
XFILL_1__1585_ vdd gnd FILL
XFILL_1__1019_ vdd gnd FILL
X_982_ _982_/A _982_/B _982_/C _991_/A vdd gnd OAI21X1
XFILL_0__1330_ vdd gnd FILL
XFILL_0__1261_ vdd gnd FILL
XFILL_2__1128_ vdd gnd FILL
XFILL_0__1192_ vdd gnd FILL
XFILL_1__994_ vdd gnd FILL
X_1323_ _1409_/A _1334_/A _1344_/C vdd gnd NAND2X1
X_1185_ _997_/B _1185_/B _1185_/C _1187_/C vdd gnd OAI21X1
XFILL_1__1370_ vdd gnd FILL
X_1254_ _1257_/C _1257_/B _1353_/A _1255_/A vdd gnd AOI21X1
XFILL_0__1459_ vdd gnd FILL
XFILL_0__1528_ vdd gnd FILL
XFILL_1__1706_ vdd gnd FILL
XFILL_1__1637_ vdd gnd FILL
XFILL_1__1499_ vdd gnd FILL
XFILL_1__1568_ vdd gnd FILL
XFILL_2__959_ vdd gnd FILL
X_965_ _973_/B _999_/B vdd gnd INVX1
XFILL_0__1313_ vdd gnd FILL
X_1872_ _1872_/A _1872_/B _1873_/C vdd gnd NAND2X1
XFILL_0__1244_ vdd gnd FILL
XFILL_0__1175_ vdd gnd FILL
X_1306_ _1319_/A _1378_/A vdd gnd INVX1
XFILL_1__977_ vdd gnd FILL
XFILL_1__1422_ vdd gnd FILL
X_1168_ _1181_/C _1170_/B vdd gnd INVX1
X_1237_ _1237_/A _1237_/B _1329_/C _1336_/B _1289_/A vdd gnd AOI22X1
XFILL_1__1353_ vdd gnd FILL
X_1099_ _1843_/B _977_/B _1194_/A vdd gnd NAND2X1
XFILL_1__1284_ vdd gnd FILL
XFILL_0__995_ vdd gnd FILL
X_948_ _971_/B _957_/B vdd gnd INVX1
XFILL_0__1793_ vdd gnd FILL
XFILL_0__1862_ vdd gnd FILL
X_1022_ _1101_/C _1022_/B _1101_/A _1031_/A vdd gnd OAI21X1
X_1855_ _1858_/B _1873_/A _1856_/A vdd gnd NOR2X1
XFILL_0__1227_ vdd gnd FILL
XFILL_0__1158_ vdd gnd FILL
XFILL_0__1089_ vdd gnd FILL
X_1786_ _1839_/A _979_/B _1786_/C _1839_/D _1788_/B vdd gnd AOI22X1
XFILL86550x46950 vdd gnd FILL
XFILL_1__1405_ vdd gnd FILL
XFILL_1__1336_ vdd gnd FILL
XFILL_1__1267_ vdd gnd FILL
XFILL_1__1198_ vdd gnd FILL
XFILL_2__1514_ vdd gnd FILL
XFILL_2__1376_ vdd gnd FILL
XFILL_0__978_ vdd gnd FILL
X_1640_ ABCmd_i[2] LoadB_i _1641_/C vdd gnd NAND2X1
XFILL_0__1012_ vdd gnd FILL
X_1571_ _1571_/A _1571_/B _1571_/C _1572_/B vdd gnd OAI21X1
XFILL_0__1845_ vdd gnd FILL
XFILL_0__1776_ vdd gnd FILL
X_1005_ _1070_/A _1057_/B vdd gnd INVX1
XFILL_1__1121_ vdd gnd FILL
X_1838_ _1881_/B _1840_/B _1839_/C vdd gnd NAND2X1
XFILL_1__1052_ vdd gnd FILL
XFILL_1__1885_ vdd gnd FILL
X_1769_ _1809_/A _980_/B _1769_/C _1771_/B vdd gnd AOI21X1
XFILL_2__1161_ vdd gnd FILL
XFILL_1__1319_ vdd gnd FILL
XFILL_0__1630_ vdd gnd FILL
XFILL_0__1492_ vdd gnd FILL
XFILL_0__1561_ vdd gnd FILL
X_1554_ _1554_/A _1555_/A vdd gnd INVX1
X_1623_ LoadA_i _982_/A _1623_/C _1670_/D vdd gnd OAI21X1
X_1485_ Flag_i _1485_/B _1485_/C _1486_/A vdd gnd AOI21X1
.ends

