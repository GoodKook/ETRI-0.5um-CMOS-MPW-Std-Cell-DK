magic
tech scmos
magscale 1 2
timestamp 1701862152
<< checkpaint >>
rect -14 142 74 159
rect -34 61 114 142
<< nwell >>
rect -13 154 93 272
<< ntransistor >>
rect 18 14 22 34
rect 38 14 42 34
rect 58 14 62 34
<< ptransistor >>
rect 18 166 22 246
rect 28 166 32 246
rect 52 206 56 246
<< ndiffusion >>
rect 16 14 18 34
rect 22 14 24 34
rect 36 14 38 34
rect 42 14 44 34
rect 56 14 58 34
rect 62 14 64 34
<< pdiffusion >>
rect 16 166 18 246
rect 22 166 28 246
rect 32 166 34 246
rect 46 206 52 246
rect 56 206 58 246
<< ndcontact >>
rect 4 14 16 34
rect 24 14 36 34
rect 44 14 56 34
rect 64 14 76 34
<< pdcontact >>
rect 4 166 16 246
rect 34 166 46 246
rect 58 206 70 246
<< psubstratepcontact >>
rect -7 -6 87 6
<< nsubstratencontact >>
rect -7 254 87 266
<< polysilicon >>
rect 18 246 22 250
rect 28 246 32 250
rect 52 246 56 250
rect 52 204 56 206
rect 52 200 62 204
rect 18 34 22 166
rect 28 142 32 166
rect 58 160 62 200
rect 28 138 42 142
rect 38 103 42 138
rect 38 34 42 91
rect 58 34 62 44
rect 18 10 22 14
rect 38 10 42 14
rect 58 10 62 14
<< polycontact >>
rect 6 117 18 129
rect 50 148 62 160
rect 30 91 42 103
rect 50 44 62 56
<< metal1 >>
rect -7 266 87 268
rect -7 252 87 254
rect 34 246 46 252
rect 60 200 74 206
rect 4 160 16 166
rect 4 154 50 160
rect 50 56 56 148
rect 68 117 74 200
rect 26 44 50 50
rect 26 34 32 44
rect 68 34 74 103
rect 4 8 16 14
rect 44 8 56 14
rect -7 6 87 8
rect -7 -8 87 -6
<< m2contact >>
rect 4 103 18 117
rect 28 103 42 117
rect 62 103 76 117
<< metal2 >>
rect 26 117 34 134
rect 26 103 28 117
rect 6 86 14 103
rect 66 86 74 103
<< m1p >>
rect -7 252 87 268
rect -7 -8 87 8
<< m2p >>
rect 26 119 34 134
rect 6 86 14 101
rect 66 86 74 101
<< labels >>
rlabel metal2 10 90 10 90 1 A
port 1 n signal input
rlabel metal2 30 131 30 131 1 B
port 2 n signal input
rlabel metal2 70 89 70 89 5 Y
port 3 n signal output
rlabel metal1 -7 252 87 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -7 -8 87 8 0 gnd
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
