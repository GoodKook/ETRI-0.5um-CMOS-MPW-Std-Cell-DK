magic
tech scmos
magscale 1 2
timestamp 1702305602
<< checkpaint >>
rect 8 177 95 180
rect -37 83 97 177
rect -35 77 95 83
rect 6 66 95 77
rect 8 65 95 66
<< nwell >>
rect -13 154 73 272
<< ntransistor >>
rect 18 14 22 34
rect 38 14 42 54
<< ptransistor >>
rect 18 206 22 246
rect 38 166 42 246
<< ndiffusion >>
rect 16 14 18 34
rect 22 14 24 34
rect 36 14 38 54
rect 42 14 44 54
<< pdiffusion >>
rect 16 206 18 246
rect 22 206 24 246
rect 36 178 38 246
rect 24 166 38 178
rect 42 167 44 246
rect 42 166 56 167
<< ndcontact >>
rect 4 14 16 34
rect 24 14 36 54
rect 44 14 56 54
<< pdcontact >>
rect 4 206 16 246
rect 24 178 36 246
rect 44 167 56 246
<< psubstratepcontact >>
rect -6 -6 66 6
<< nsubstratencontact >>
rect -6 254 66 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 18 117 22 206
rect 38 161 42 166
rect 17 105 22 117
rect 18 34 22 105
rect 38 54 42 60
rect 18 10 22 14
rect 38 10 42 14
<< polycontact >>
rect 30 149 42 161
rect 5 105 17 117
rect 30 60 42 72
<< metal1 >>
rect -6 266 66 268
rect -6 252 66 254
rect 24 246 36 252
rect 4 161 12 206
rect 4 154 30 161
rect 3 123 17 137
rect 5 117 17 123
rect 30 72 37 149
rect 48 137 56 167
rect 43 123 57 137
rect 4 60 30 68
rect 4 34 12 60
rect 48 54 56 123
rect 24 8 36 14
rect -6 6 66 8
rect -6 -8 66 -6
<< m1p >>
rect -6 252 66 268
rect 3 123 17 137
rect 43 123 57 137
rect -6 -8 66 8
<< labels >>
rlabel nsubstratencontact 29 260 29 260 0 vdd
port 3 nsew power bidirectional abutment
rlabel psubstratepcontact 31 0 31 0 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 10 127 10 127 0 A
port 1 nsew signal input
rlabel metal1 50 127 50 127 0 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 60 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
