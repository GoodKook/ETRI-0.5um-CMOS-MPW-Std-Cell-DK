magic
tech scmos
magscale 1 2
timestamp 1701862152
<< checkpaint >>
rect -14 142 74 159
rect -34 78 74 142
rect -34 61 54 78
<< nwell >>
rect -12 154 52 272
<< ntransistor >>
rect 18 14 22 34
<< ptransistor >>
rect 18 206 22 246
<< ndiffusion >>
rect 16 14 18 34
rect 22 14 24 34
<< pdiffusion >>
rect 16 206 18 246
rect 22 206 24 246
<< ndcontact >>
rect 4 14 16 34
rect 24 14 36 34
<< pdcontact >>
rect 4 206 16 246
rect 24 206 36 246
<< psubstratepcontact >>
rect -6 -6 46 6
<< nsubstratencontact >>
rect -6 254 46 266
<< polysilicon >>
rect 18 246 22 250
rect 18 129 22 206
rect 16 117 22 129
rect 18 34 22 117
rect 18 10 22 14
<< polycontact >>
rect 4 117 16 129
<< metal1 >>
rect -6 266 46 268
rect -6 252 46 254
rect 4 246 16 252
rect 24 117 32 206
rect 24 34 32 103
rect 4 8 16 14
rect -6 6 46 8
rect -6 -8 46 -6
<< m2contact >>
rect 3 103 17 117
rect 23 103 37 117
<< metal2 >>
rect 26 117 34 134
rect 6 86 14 103
<< m1p >>
rect -6 252 46 268
rect -6 -8 46 8
<< m2p >>
rect 26 119 34 134
rect 6 86 14 101
<< labels >>
rlabel metal2 10 90 10 90 1 A
port 1 n signal input
rlabel metal2 28 128 28 128 1 Y
port 2 n signal output
rlabel metal1 -6 252 46 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -6 -8 46 8 0 gnd
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 40 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
