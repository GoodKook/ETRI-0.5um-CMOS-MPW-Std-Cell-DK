magic
tech scmos
magscale 1 3
timestamp 1569140870
<< checkpaint >>
rect -56 -56 84 84
<< diffusion >>
rect 5 5 23 23
<< genericcontact >>
rect 11 11 17 17
<< metal1 >>
rect 4 4 24 24
<< end >>
