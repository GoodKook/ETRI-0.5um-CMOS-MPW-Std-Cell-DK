magic
tech scmos
magscale 1 30
timestamp 1726627926
<< checkpaint >>
rect -229 25660 2111 25670
rect 2250 25660 5865 26265
rect -600 23455 5865 25660
rect -660 20400 5865 23455
rect -600 19795 5865 20400
rect -660 11805 5865 19795
rect -735 10515 5865 11805
rect -600 -590 5865 10515
rect -570 -600 5865 -590
rect -229 -604 3786 -600
rect -175 -606 3786 -604
rect 1516 -615 3786 -606
<< nwell >>
rect -60 21000 2940 22855
rect -60 11205 2940 19195
<< psubstratepdiff >>
rect 30 23400 2850 25060
rect 30 0 2850 7800
<< nsubstratendiff >>
rect 30 21100 2850 22760
rect 30 11290 2850 19100
<< metal1 >>
rect 30 23400 2850 25060
rect 30 21100 2850 22760
rect 30 11290 2850 19100
rect 30 0 2850 7800
<< metal2 >>
rect 30 23400 2850 25060
rect 30 21100 2850 22760
rect 30 11290 2850 19100
rect 30 0 2850 7800
<< metal3 >>
rect 30 23400 2850 25060
rect 30 21100 2850 22760
rect 30 11290 2850 19100
rect 30 0 2850 7800
use IOFILLER10  IOFILLER10_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1537935238
transform 1 0 415 0 1 0
box -35 0 1035 25060
use IOFILLER10  IOFILLER10_1
timestamp 1537935238
transform 1 0 1495 0 1 0
box -35 0 1035 25060
<< end >>
