magic
tech scmos
magscale 2 1
timestamp 1756365015
<< checkpaint >>
rect -39 402 403 450
rect -39 41 451 402
rect -40 -40 451 41
<< metal1 >>
rect 1 143 407 362
rect 1 142 204 143
rect 224 142 407 143
rect 1 141 196 142
rect 240 141 407 142
rect 1 140 192 141
rect 249 140 407 141
rect 1 139 187 140
rect 258 139 407 140
rect 1 138 184 139
rect 265 138 407 139
rect 1 137 180 138
rect 185 137 188 138
rect 206 137 223 138
rect 272 137 407 138
rect 1 136 177 137
rect 182 136 188 137
rect 201 136 232 137
rect 279 136 407 137
rect 1 135 175 136
rect 179 135 187 136
rect 197 135 239 136
rect 284 135 407 136
rect 1 134 171 135
rect 176 134 185 135
rect 194 134 245 135
rect 290 134 407 135
rect 1 133 169 134
rect 174 133 183 134
rect 191 133 250 134
rect 295 133 407 134
rect 1 132 166 133
rect 171 132 181 133
rect 188 132 254 133
rect 301 132 407 133
rect 1 131 164 132
rect 169 131 179 132
rect 186 131 258 132
rect 306 131 407 132
rect 1 130 162 131
rect 166 130 177 131
rect 183 130 262 131
rect 310 130 407 131
rect 1 129 159 130
rect 163 129 175 130
rect 181 129 264 130
rect 315 129 407 130
rect 1 128 157 129
rect 161 128 174 129
rect 179 128 267 129
rect 319 128 407 129
rect 1 127 155 128
rect 158 127 172 128
rect 177 127 268 128
rect 324 127 407 128
rect 1 126 153 127
rect 156 126 170 127
rect 175 126 269 127
rect 328 126 407 127
rect 1 125 151 126
rect 153 125 168 126
rect 173 125 270 126
rect 333 125 407 126
rect 1 124 149 125
rect 151 124 166 125
rect 171 124 268 125
rect 337 124 407 125
rect 1 123 147 124
rect 148 123 165 124
rect 170 123 265 124
rect 341 123 407 124
rect 1 122 163 123
rect 168 122 260 123
rect 287 122 300 123
rect 345 122 407 123
rect 1 121 161 122
rect 166 121 256 122
rect 275 121 282 122
rect 287 121 318 122
rect 349 121 407 122
rect 1 120 159 121
rect 165 120 250 121
rect 268 120 281 121
rect 287 120 333 121
rect 353 120 407 121
rect 1 119 157 120
rect 163 119 244 120
rect 262 119 280 120
rect 286 119 344 120
rect 356 119 407 120
rect 1 118 155 119
rect 161 118 237 119
rect 256 118 279 119
rect 285 118 356 119
rect 359 118 407 119
rect 1 117 154 118
rect 160 117 229 118
rect 251 117 278 118
rect 285 117 407 118
rect 1 116 152 117
rect 158 116 220 117
rect 245 116 277 117
rect 284 116 407 117
rect 1 115 150 116
rect 157 115 206 116
rect 240 115 276 116
rect 282 115 407 116
rect 1 114 108 115
rect 234 114 275 115
rect 281 114 407 115
rect 1 113 101 114
rect 227 113 274 114
rect 279 113 407 114
rect 1 112 97 113
rect 220 112 273 113
rect 277 112 407 113
rect 1 111 93 112
rect 209 111 272 112
rect 274 111 407 112
rect 1 110 90 111
rect 197 110 407 111
rect 1 109 87 110
rect 106 109 300 110
rect 310 109 407 110
rect 1 108 84 109
rect 101 108 296 109
rect 314 108 407 109
rect 1 107 81 108
rect 96 107 108 108
rect 119 107 294 108
rect 316 107 407 108
rect 1 106 78 107
rect 92 106 104 107
rect 123 106 292 107
rect 297 106 313 107
rect 319 106 407 107
rect 1 105 76 106
rect 89 105 102 106
rect 112 105 115 106
rect 125 105 290 106
rect 295 105 316 106
rect 320 105 407 106
rect 1 104 73 105
rect 85 104 100 105
rect 106 104 122 105
rect 127 104 289 105
rect 292 104 318 105
rect 321 104 407 105
rect 1 103 71 104
rect 82 103 99 104
rect 103 103 125 104
rect 129 103 288 104
rect 290 103 320 104
rect 323 103 407 104
rect 1 102 69 103
rect 78 102 97 103
rect 101 102 127 103
rect 130 102 287 103
rect 289 102 322 103
rect 324 102 407 103
rect 1 101 66 102
rect 75 101 96 102
rect 99 101 129 102
rect 131 101 286 102
rect 287 101 323 102
rect 325 101 407 102
rect 1 100 64 101
rect 73 100 95 101
rect 97 100 130 101
rect 132 100 285 101
rect 286 100 324 101
rect 326 100 407 101
rect 1 99 61 100
rect 69 99 94 100
rect 96 99 132 100
rect 133 99 284 100
rect 285 99 325 100
rect 1 98 59 99
rect 67 98 93 99
rect 95 98 133 99
rect 134 98 283 99
rect 284 98 326 99
rect 327 98 407 100
rect 1 97 57 98
rect 64 97 92 98
rect 1 96 55 97
rect 61 96 92 97
rect 93 97 134 98
rect 135 97 327 98
rect 328 97 407 98
rect 93 96 135 97
rect 136 96 328 97
rect 329 96 407 97
rect 1 95 53 96
rect 58 95 91 96
rect 92 95 407 96
rect 1 94 51 95
rect 55 94 407 95
rect 1 93 49 94
rect 53 93 407 94
rect 1 92 47 93
rect 50 92 407 93
rect 1 91 45 92
rect 48 91 407 92
rect 1 90 43 91
rect 45 90 407 91
rect 1 89 41 90
rect 42 89 407 90
rect 1 74 407 89
rect 1 73 193 74
rect 199 73 371 74
rect 374 73 407 74
rect 1 72 52 73
rect 66 72 190 73
rect 200 72 209 73
rect 213 72 224 73
rect 228 72 244 73
rect 260 72 295 73
rect 302 72 370 73
rect 1 71 44 72
rect 67 71 82 72
rect 85 71 145 72
rect 149 71 187 72
rect 202 71 208 72
rect 215 71 223 72
rect 229 71 236 72
rect 263 71 290 72
rect 304 71 314 72
rect 1 70 42 71
rect 68 70 81 71
rect 85 70 143 71
rect 149 70 185 71
rect 202 70 207 71
rect 215 70 221 71
rect 230 70 234 71
rect 264 70 286 71
rect 305 70 312 71
rect 318 70 369 72
rect 376 70 407 73
rect 1 68 40 70
rect 69 69 79 70
rect 85 69 142 70
rect 148 69 183 70
rect 202 69 206 70
rect 216 69 220 70
rect 230 69 233 70
rect 265 69 284 70
rect 305 69 310 70
rect 69 68 78 69
rect 85 68 140 69
rect 148 68 181 69
rect 202 68 205 69
rect 215 68 219 69
rect 1 65 39 68
rect 69 67 77 68
rect 85 67 139 68
rect 147 67 181 68
rect 195 67 196 68
rect 202 67 204 68
rect 215 67 218 68
rect 230 67 232 69
rect 265 68 282 69
rect 305 68 308 69
rect 318 68 368 70
rect 375 68 407 70
rect 265 67 281 68
rect 304 67 307 68
rect 317 67 367 68
rect 69 66 76 67
rect 84 66 138 67
rect 146 66 180 67
rect 193 66 196 67
rect 56 65 63 66
rect 69 65 75 66
rect 83 65 137 66
rect 145 65 180 66
rect 191 65 196 66
rect 201 66 203 67
rect 215 66 217 67
rect 229 66 231 67
rect 249 66 259 67
rect 201 65 202 66
rect 214 65 216 66
rect 228 65 231 66
rect 243 65 260 66
rect 1 62 38 65
rect 50 64 63 65
rect 68 64 74 65
rect 82 64 136 65
rect 144 64 180 65
rect 189 64 195 65
rect 206 64 207 65
rect 213 64 215 65
rect 47 63 62 64
rect 67 63 73 64
rect 82 63 135 64
rect 143 63 180 64
rect 49 62 61 63
rect 66 62 72 63
rect 81 62 134 63
rect 142 62 180 63
rect 190 63 195 64
rect 205 63 206 64
rect 213 63 214 64
rect 227 63 230 65
rect 240 64 244 65
rect 248 64 259 65
rect 265 64 280 67
rect 295 66 298 67
rect 303 66 305 67
rect 316 66 367 67
rect 374 66 407 68
rect 292 64 297 66
rect 311 65 312 66
rect 315 65 367 66
rect 373 65 407 66
rect 309 64 323 65
rect 190 62 194 63
rect 204 62 206 63
rect 212 62 213 63
rect 226 62 230 63
rect 241 63 243 64
rect 247 63 258 64
rect 265 63 279 64
rect 292 63 296 64
rect 307 63 322 64
rect 327 63 366 65
rect 372 63 407 65
rect 241 62 242 63
rect 1 61 39 62
rect 49 61 60 62
rect 65 61 71 62
rect 80 61 133 62
rect 141 61 157 62
rect 160 61 180 62
rect 187 61 193 62
rect 203 61 205 62
rect 211 61 212 62
rect 225 61 242 62
rect 246 62 257 63
rect 264 62 279 63
rect 289 62 295 63
rect 305 62 321 63
rect 246 61 254 62
rect 263 61 280 62
rect 285 61 294 62
rect 303 61 321 62
rect 327 61 365 63
rect 371 61 407 63
rect 1 59 59 61
rect 64 59 70 61
rect 79 60 132 61
rect 140 60 155 61
rect 161 60 193 61
rect 202 60 204 61
rect 78 59 95 60
rect 103 59 122 60
rect 125 59 132 60
rect 139 59 142 60
rect 1 58 58 59
rect 63 58 69 59
rect 77 58 93 59
rect 104 58 113 59
rect 117 58 120 59
rect 126 58 131 59
rect 138 58 140 59
rect 147 58 154 60
rect 1 57 57 58
rect 1 56 56 57
rect 62 56 68 58
rect 76 57 79 58
rect 82 57 91 58
rect 104 57 111 58
rect 118 57 119 58
rect 75 56 77 57
rect 84 56 89 57
rect 1 54 55 56
rect 61 55 67 56
rect 60 54 67 55
rect 74 55 76 56
rect 84 55 88 56
rect 104 55 110 57
rect 117 56 118 57
rect 126 56 130 58
rect 137 57 139 58
rect 148 57 154 58
rect 161 59 192 60
rect 201 59 204 60
rect 215 60 217 61
rect 224 60 241 61
rect 245 60 251 61
rect 262 60 293 61
rect 301 60 321 61
rect 326 60 364 61
rect 215 59 216 60
rect 223 59 240 60
rect 245 59 248 60
rect 261 59 291 60
rect 299 59 321 60
rect 325 59 341 60
rect 346 59 351 60
rect 353 59 364 60
rect 370 59 407 61
rect 161 58 191 59
rect 200 58 203 59
rect 214 58 215 59
rect 223 58 239 59
rect 259 58 289 59
rect 161 57 190 58
rect 199 57 202 58
rect 213 57 215 58
rect 222 57 238 58
rect 256 57 289 58
rect 297 58 319 59
rect 322 58 331 59
rect 336 58 340 59
rect 346 58 350 59
rect 354 58 364 59
rect 297 57 317 58
rect 323 57 330 58
rect 336 57 339 58
rect 346 57 348 58
rect 136 56 137 57
rect 148 56 153 57
rect 161 56 189 57
rect 198 56 202 57
rect 212 56 214 57
rect 221 56 235 57
rect 253 56 288 57
rect 297 56 316 57
rect 323 56 329 57
rect 336 56 337 57
rect 346 56 347 57
rect 116 55 117 56
rect 126 55 129 56
rect 135 55 136 56
rect 141 55 142 56
rect 148 55 152 56
rect 74 54 75 55
rect 83 54 87 55
rect 96 54 97 55
rect 104 54 109 55
rect 115 54 116 55
rect 125 54 128 55
rect 134 54 135 55
rect 140 54 142 55
rect 147 54 151 55
rect 155 54 156 55
rect 1 53 54 54
rect 60 53 66 54
rect 73 53 74 54
rect 83 53 86 54
rect 94 53 96 54
rect 1 52 53 53
rect 1 50 52 52
rect 59 51 66 53
rect 72 52 73 53
rect 82 52 85 53
rect 92 52 95 53
rect 103 52 108 54
rect 114 53 115 54
rect 113 52 114 53
rect 124 52 128 54
rect 133 53 134 54
rect 139 53 141 54
rect 146 53 150 54
rect 154 53 156 54
rect 161 54 188 56
rect 197 55 201 56
rect 211 55 213 56
rect 196 54 200 55
rect 210 54 213 55
rect 220 54 233 56
rect 248 55 288 56
rect 299 55 315 56
rect 242 54 288 55
rect 300 54 315 55
rect 322 54 328 56
rect 335 55 336 56
rect 345 55 346 56
rect 334 54 335 55
rect 355 54 363 58
rect 369 54 407 59
rect 161 53 187 54
rect 196 53 199 54
rect 209 53 212 54
rect 219 53 232 54
rect 246 53 288 54
rect 302 53 314 54
rect 321 53 327 54
rect 333 53 334 54
rect 354 53 363 54
rect 368 53 407 54
rect 132 52 133 53
rect 138 52 140 53
rect 146 52 149 53
rect 153 52 155 53
rect 71 51 72 52
rect 81 51 85 52
rect 91 51 94 52
rect 102 51 106 52
rect 123 51 126 52
rect 137 51 139 52
rect 145 51 147 52
rect 152 51 155 52
rect 161 52 186 53
rect 195 52 198 53
rect 208 52 211 53
rect 161 51 164 52
rect 165 51 185 52
rect 194 51 198 52
rect 207 51 211 52
rect 218 52 231 53
rect 249 52 287 53
rect 303 52 313 53
rect 320 52 327 53
rect 353 52 363 53
rect 367 52 407 53
rect 218 51 227 52
rect 229 51 232 52
rect 253 51 286 52
rect 292 51 293 52
rect 305 51 313 52
rect 319 51 326 52
rect 352 51 356 52
rect 358 51 364 52
rect 59 50 65 51
rect 70 50 71 51
rect 81 50 84 51
rect 90 50 93 51
rect 101 50 105 51
rect 122 50 125 51
rect 143 50 146 51
rect 151 50 155 51
rect 160 50 162 51
rect 165 50 184 51
rect 193 50 197 51
rect 1 49 51 50
rect 1 47 50 49
rect 1 42 49 47
rect 58 46 65 50
rect 80 49 82 50
rect 89 49 92 50
rect 101 49 103 50
rect 121 49 123 50
rect 142 49 145 50
rect 151 49 154 50
rect 159 49 161 50
rect 165 49 183 50
rect 89 48 91 49
rect 100 48 101 49
rect 140 48 144 49
rect 158 48 159 49
rect 164 48 182 49
rect 192 48 196 50
rect 206 49 210 51
rect 218 50 225 51
rect 229 50 234 51
rect 255 50 285 51
rect 291 50 295 51
rect 307 50 313 51
rect 205 48 210 49
rect 217 49 223 50
rect 229 49 233 50
rect 257 49 267 50
rect 272 49 284 50
rect 290 49 296 50
rect 308 49 313 50
rect 318 50 324 51
rect 336 50 337 51
rect 351 50 354 51
rect 358 50 361 51
rect 365 50 407 52
rect 318 49 323 50
rect 335 49 336 50
rect 351 49 353 50
rect 358 49 360 50
rect 217 48 222 49
rect 227 48 232 49
rect 73 47 74 48
rect 114 47 115 48
rect 126 47 127 48
rect 141 47 142 48
rect 163 47 183 48
rect 191 47 195 48
rect 204 47 210 48
rect 218 47 219 48
rect 226 47 232 48
rect 238 48 241 49
rect 259 48 266 49
rect 273 48 283 49
rect 290 48 298 49
rect 310 48 313 49
rect 317 48 321 49
rect 334 48 336 49
rect 350 48 351 49
rect 357 48 360 49
rect 238 47 244 48
rect 72 46 73 47
rect 83 46 84 47
rect 105 46 106 47
rect 113 46 115 47
rect 125 46 127 47
rect 133 46 134 47
rect 146 46 147 47
rect 162 46 183 47
rect 58 45 66 46
rect 71 45 73 46
rect 82 45 85 46
rect 93 45 94 46
rect 103 45 107 46
rect 112 45 115 46
rect 123 45 127 46
rect 132 45 135 46
rect 145 45 148 46
rect 160 45 183 46
rect 190 45 195 47
rect 203 45 210 47
rect 225 46 231 47
rect 238 46 247 47
rect 260 46 265 48
rect 273 47 282 48
rect 224 45 230 46
rect 238 45 249 46
rect 261 45 265 46
rect 272 46 282 47
rect 289 47 299 48
rect 311 47 313 48
rect 318 47 319 48
rect 334 47 335 48
rect 343 47 344 48
rect 356 47 360 48
rect 289 46 301 47
rect 272 45 281 46
rect 289 45 302 46
rect 56 44 66 45
rect 70 44 73 45
rect 80 44 86 45
rect 91 44 94 45
rect 102 44 107 45
rect 111 44 116 45
rect 121 44 128 45
rect 131 44 136 45
rect 144 44 150 45
rect 159 44 184 45
rect 189 44 196 45
rect 202 44 210 45
rect 222 44 230 45
rect 237 44 252 45
rect 261 44 266 45
rect 271 44 281 45
rect 287 44 304 45
rect 312 44 313 47
rect 324 46 325 47
rect 333 46 335 47
rect 342 46 344 47
rect 355 46 360 47
rect 323 45 326 46
rect 332 45 334 46
rect 341 45 344 46
rect 353 45 360 46
rect 366 45 407 50
rect 322 44 327 45
rect 331 44 334 45
rect 340 44 344 45
rect 352 44 361 45
rect 365 44 407 45
rect 55 43 74 44
rect 78 43 95 44
rect 100 43 137 44
rect 142 43 185 44
rect 187 43 196 44
rect 201 43 211 44
rect 221 43 230 44
rect 236 43 254 44
rect 261 43 306 44
rect 312 43 314 44
rect 320 43 335 44
rect 339 43 344 44
rect 350 43 407 44
rect 53 42 197 43
rect 200 42 213 43
rect 219 42 230 43
rect 235 42 256 43
rect 260 42 308 43
rect 312 42 407 43
rect 1 41 231 42
rect 232 41 407 42
rect 1 4 407 41
<< metal2 >>
rect 3 141 409 360
rect 3 140 206 141
rect 226 140 409 141
rect 3 139 198 140
rect 242 139 409 140
rect 3 138 194 139
rect 251 138 409 139
rect 3 137 189 138
rect 260 137 409 138
rect 3 136 186 137
rect 267 136 409 137
rect 3 135 182 136
rect 187 135 190 136
rect 208 135 225 136
rect 274 135 409 136
rect 3 134 179 135
rect 184 134 190 135
rect 203 134 234 135
rect 281 134 409 135
rect 3 133 177 134
rect 181 133 189 134
rect 199 133 241 134
rect 286 133 409 134
rect 3 132 173 133
rect 178 132 187 133
rect 196 132 247 133
rect 292 132 409 133
rect 3 131 171 132
rect 176 131 185 132
rect 193 131 252 132
rect 297 131 409 132
rect 3 130 168 131
rect 173 130 183 131
rect 190 130 256 131
rect 303 130 409 131
rect 3 129 166 130
rect 171 129 181 130
rect 188 129 260 130
rect 308 129 409 130
rect 3 128 164 129
rect 168 128 179 129
rect 185 128 264 129
rect 312 128 409 129
rect 3 127 161 128
rect 165 127 177 128
rect 183 127 266 128
rect 317 127 409 128
rect 3 126 159 127
rect 163 126 176 127
rect 181 126 269 127
rect 321 126 409 127
rect 3 125 157 126
rect 160 125 174 126
rect 179 125 270 126
rect 326 125 409 126
rect 3 124 155 125
rect 158 124 172 125
rect 177 124 271 125
rect 330 124 409 125
rect 3 123 153 124
rect 155 123 170 124
rect 175 123 272 124
rect 335 123 409 124
rect 3 122 151 123
rect 153 122 168 123
rect 173 122 270 123
rect 339 122 409 123
rect 3 121 149 122
rect 150 121 167 122
rect 172 121 267 122
rect 343 121 409 122
rect 3 120 165 121
rect 170 120 262 121
rect 289 120 302 121
rect 347 120 409 121
rect 3 119 163 120
rect 168 119 258 120
rect 277 119 284 120
rect 289 119 320 120
rect 351 119 409 120
rect 3 118 161 119
rect 167 118 252 119
rect 270 118 283 119
rect 289 118 335 119
rect 355 118 409 119
rect 3 117 159 118
rect 165 117 246 118
rect 264 117 282 118
rect 288 117 346 118
rect 358 117 409 118
rect 3 116 157 117
rect 163 116 239 117
rect 258 116 281 117
rect 287 116 358 117
rect 361 116 409 117
rect 3 115 156 116
rect 162 115 231 116
rect 253 115 280 116
rect 287 115 409 116
rect 3 114 154 115
rect 160 114 222 115
rect 247 114 279 115
rect 286 114 409 115
rect 3 113 152 114
rect 159 113 208 114
rect 242 113 278 114
rect 284 113 409 114
rect 3 112 110 113
rect 236 112 277 113
rect 283 112 409 113
rect 3 111 103 112
rect 229 111 276 112
rect 281 111 409 112
rect 3 110 99 111
rect 222 110 275 111
rect 279 110 409 111
rect 3 109 95 110
rect 211 109 274 110
rect 276 109 409 110
rect 3 108 92 109
rect 199 108 409 109
rect 3 107 89 108
rect 108 107 302 108
rect 312 107 409 108
rect 3 106 86 107
rect 103 106 298 107
rect 316 106 409 107
rect 3 105 83 106
rect 98 105 110 106
rect 121 105 296 106
rect 318 105 409 106
rect 3 104 80 105
rect 94 104 106 105
rect 125 104 294 105
rect 299 104 315 105
rect 321 104 409 105
rect 3 103 78 104
rect 91 103 104 104
rect 114 103 117 104
rect 127 103 292 104
rect 297 103 318 104
rect 322 103 409 104
rect 3 102 75 103
rect 87 102 102 103
rect 108 102 124 103
rect 129 102 291 103
rect 294 102 320 103
rect 323 102 409 103
rect 3 101 73 102
rect 84 101 101 102
rect 105 101 127 102
rect 131 101 290 102
rect 292 101 322 102
rect 325 101 409 102
rect 3 100 71 101
rect 80 100 99 101
rect 103 100 129 101
rect 132 100 289 101
rect 291 100 324 101
rect 326 100 409 101
rect 3 99 68 100
rect 77 99 98 100
rect 101 99 131 100
rect 133 99 288 100
rect 289 99 325 100
rect 327 99 409 100
rect 3 98 66 99
rect 75 98 97 99
rect 99 98 132 99
rect 134 98 287 99
rect 288 98 326 99
rect 328 98 409 99
rect 3 97 63 98
rect 71 97 96 98
rect 98 97 134 98
rect 135 97 286 98
rect 287 97 327 98
rect 3 96 61 97
rect 69 96 95 97
rect 97 96 135 97
rect 136 96 285 97
rect 286 96 328 97
rect 329 96 409 98
rect 3 95 59 96
rect 66 95 94 96
rect 3 94 57 95
rect 63 94 94 95
rect 95 95 136 96
rect 137 95 329 96
rect 330 95 409 96
rect 95 94 137 95
rect 138 94 330 95
rect 331 94 409 95
rect 3 93 55 94
rect 60 93 93 94
rect 94 93 409 94
rect 3 92 53 93
rect 57 92 409 93
rect 3 91 51 92
rect 55 91 409 92
rect 3 90 49 91
rect 52 90 409 91
rect 3 89 47 90
rect 50 89 409 90
rect 3 88 45 89
rect 47 88 409 89
rect 3 87 43 88
rect 44 87 409 88
rect 3 72 409 87
rect 3 71 195 72
rect 201 71 373 72
rect 376 71 409 72
rect 3 70 54 71
rect 68 70 192 71
rect 202 70 211 71
rect 215 70 226 71
rect 230 70 246 71
rect 262 70 297 71
rect 304 70 372 71
rect 3 69 46 70
rect 69 69 84 70
rect 87 69 147 70
rect 151 69 189 70
rect 204 69 210 70
rect 217 69 225 70
rect 231 69 238 70
rect 265 69 292 70
rect 306 69 316 70
rect 3 68 44 69
rect 70 68 83 69
rect 87 68 145 69
rect 151 68 187 69
rect 204 68 209 69
rect 217 68 223 69
rect 232 68 236 69
rect 266 68 288 69
rect 307 68 314 69
rect 320 68 371 70
rect 378 68 409 71
rect 3 66 42 68
rect 71 67 81 68
rect 87 67 144 68
rect 150 67 185 68
rect 204 67 208 68
rect 218 67 222 68
rect 232 67 235 68
rect 267 67 286 68
rect 307 67 312 68
rect 71 66 80 67
rect 87 66 142 67
rect 150 66 183 67
rect 204 66 207 67
rect 217 66 221 67
rect 3 63 41 66
rect 71 65 79 66
rect 87 65 141 66
rect 149 65 183 66
rect 197 65 198 66
rect 204 65 206 66
rect 217 65 220 66
rect 232 65 234 67
rect 267 66 284 67
rect 307 66 310 67
rect 320 66 370 68
rect 377 66 409 68
rect 267 65 283 66
rect 306 65 309 66
rect 319 65 369 66
rect 71 64 78 65
rect 86 64 140 65
rect 148 64 182 65
rect 195 64 198 65
rect 58 63 65 64
rect 71 63 77 64
rect 85 63 139 64
rect 147 63 182 64
rect 193 63 198 64
rect 203 64 205 65
rect 217 64 219 65
rect 231 64 233 65
rect 251 64 261 65
rect 203 63 204 64
rect 216 63 218 64
rect 230 63 233 64
rect 245 63 262 64
rect 3 60 40 63
rect 52 62 65 63
rect 70 62 76 63
rect 84 62 138 63
rect 146 62 182 63
rect 191 62 197 63
rect 208 62 209 63
rect 215 62 217 63
rect 49 61 64 62
rect 69 61 75 62
rect 84 61 137 62
rect 145 61 182 62
rect 51 60 63 61
rect 68 60 74 61
rect 83 60 136 61
rect 144 60 182 61
rect 192 61 197 62
rect 207 61 208 62
rect 215 61 216 62
rect 229 61 232 63
rect 242 62 246 63
rect 250 62 261 63
rect 267 62 282 65
rect 297 64 300 65
rect 305 64 307 65
rect 318 64 369 65
rect 376 64 409 66
rect 294 62 299 64
rect 313 63 314 64
rect 317 63 369 64
rect 375 63 409 64
rect 311 62 325 63
rect 192 60 196 61
rect 206 60 208 61
rect 214 60 215 61
rect 228 60 232 61
rect 243 61 245 62
rect 249 61 260 62
rect 267 61 281 62
rect 294 61 298 62
rect 309 61 324 62
rect 329 61 368 63
rect 374 61 409 63
rect 243 60 244 61
rect 3 59 41 60
rect 51 59 62 60
rect 67 59 73 60
rect 82 59 135 60
rect 143 59 159 60
rect 162 59 182 60
rect 189 59 195 60
rect 205 59 207 60
rect 213 59 214 60
rect 227 59 244 60
rect 248 60 259 61
rect 266 60 281 61
rect 291 60 297 61
rect 307 60 323 61
rect 248 59 256 60
rect 265 59 282 60
rect 287 59 296 60
rect 305 59 323 60
rect 329 59 367 61
rect 373 59 409 61
rect 3 57 61 59
rect 66 57 72 59
rect 81 58 134 59
rect 142 58 157 59
rect 163 58 195 59
rect 204 58 206 59
rect 80 57 97 58
rect 105 57 124 58
rect 127 57 134 58
rect 141 57 144 58
rect 3 56 60 57
rect 65 56 71 57
rect 79 56 95 57
rect 106 56 115 57
rect 119 56 122 57
rect 128 56 133 57
rect 140 56 142 57
rect 149 56 156 58
rect 3 55 59 56
rect 3 54 58 55
rect 64 54 70 56
rect 78 55 81 56
rect 84 55 93 56
rect 106 55 113 56
rect 120 55 121 56
rect 77 54 79 55
rect 86 54 91 55
rect 3 52 57 54
rect 63 53 69 54
rect 62 52 69 53
rect 76 53 78 54
rect 86 53 90 54
rect 106 53 112 55
rect 119 54 120 55
rect 128 54 132 56
rect 139 55 141 56
rect 150 55 156 56
rect 163 57 194 58
rect 203 57 206 58
rect 217 58 219 59
rect 226 58 243 59
rect 247 58 253 59
rect 264 58 295 59
rect 303 58 323 59
rect 328 58 366 59
rect 217 57 218 58
rect 225 57 242 58
rect 247 57 250 58
rect 263 57 293 58
rect 301 57 323 58
rect 327 57 343 58
rect 348 57 353 58
rect 355 57 366 58
rect 372 57 409 59
rect 163 56 193 57
rect 202 56 205 57
rect 216 56 217 57
rect 225 56 241 57
rect 261 56 291 57
rect 163 55 192 56
rect 201 55 204 56
rect 215 55 217 56
rect 224 55 240 56
rect 258 55 291 56
rect 299 56 321 57
rect 324 56 333 57
rect 338 56 342 57
rect 348 56 352 57
rect 356 56 366 57
rect 299 55 319 56
rect 325 55 332 56
rect 338 55 341 56
rect 348 55 350 56
rect 138 54 139 55
rect 150 54 155 55
rect 163 54 191 55
rect 200 54 204 55
rect 214 54 216 55
rect 223 54 237 55
rect 255 54 290 55
rect 299 54 318 55
rect 325 54 331 55
rect 338 54 339 55
rect 348 54 349 55
rect 118 53 119 54
rect 128 53 131 54
rect 137 53 138 54
rect 143 53 144 54
rect 150 53 154 54
rect 76 52 77 53
rect 85 52 89 53
rect 98 52 99 53
rect 106 52 111 53
rect 117 52 118 53
rect 127 52 130 53
rect 136 52 137 53
rect 142 52 144 53
rect 149 52 153 53
rect 157 52 158 53
rect 3 51 56 52
rect 62 51 68 52
rect 75 51 76 52
rect 85 51 88 52
rect 96 51 98 52
rect 3 50 55 51
rect 3 48 54 50
rect 61 49 68 51
rect 74 50 75 51
rect 84 50 87 51
rect 94 50 97 51
rect 105 50 110 52
rect 116 51 117 52
rect 115 50 116 51
rect 126 50 130 52
rect 135 51 136 52
rect 141 51 143 52
rect 148 51 152 52
rect 156 51 158 52
rect 163 52 190 54
rect 199 53 203 54
rect 213 53 215 54
rect 198 52 202 53
rect 212 52 215 53
rect 222 52 235 54
rect 250 53 290 54
rect 301 53 317 54
rect 244 52 290 53
rect 302 52 317 53
rect 324 52 330 54
rect 337 53 338 54
rect 347 53 348 54
rect 336 52 337 53
rect 357 52 365 56
rect 371 52 409 57
rect 163 51 189 52
rect 198 51 201 52
rect 211 51 214 52
rect 221 51 234 52
rect 248 51 290 52
rect 304 51 316 52
rect 323 51 329 52
rect 335 51 336 52
rect 356 51 365 52
rect 370 51 409 52
rect 134 50 135 51
rect 140 50 142 51
rect 148 50 151 51
rect 155 50 157 51
rect 73 49 74 50
rect 83 49 87 50
rect 93 49 96 50
rect 104 49 108 50
rect 125 49 128 50
rect 139 49 141 50
rect 147 49 149 50
rect 154 49 157 50
rect 163 50 188 51
rect 197 50 200 51
rect 210 50 213 51
rect 163 49 166 50
rect 167 49 187 50
rect 196 49 200 50
rect 209 49 213 50
rect 220 50 233 51
rect 251 50 289 51
rect 305 50 315 51
rect 322 50 329 51
rect 355 50 365 51
rect 369 50 409 51
rect 220 49 229 50
rect 231 49 234 50
rect 255 49 288 50
rect 294 49 295 50
rect 307 49 315 50
rect 321 49 328 50
rect 354 49 358 50
rect 360 49 366 50
rect 61 48 67 49
rect 72 48 73 49
rect 83 48 86 49
rect 92 48 95 49
rect 103 48 107 49
rect 124 48 127 49
rect 145 48 148 49
rect 153 48 157 49
rect 162 48 164 49
rect 167 48 186 49
rect 195 48 199 49
rect 3 47 53 48
rect 3 45 52 47
rect 3 40 51 45
rect 60 44 67 48
rect 82 47 84 48
rect 91 47 94 48
rect 103 47 105 48
rect 123 47 125 48
rect 144 47 147 48
rect 153 47 156 48
rect 161 47 163 48
rect 167 47 185 48
rect 91 46 93 47
rect 102 46 103 47
rect 142 46 146 47
rect 160 46 161 47
rect 166 46 184 47
rect 194 46 198 48
rect 208 47 212 49
rect 220 48 227 49
rect 231 48 236 49
rect 257 48 287 49
rect 293 48 297 49
rect 309 48 315 49
rect 207 46 212 47
rect 219 47 225 48
rect 231 47 235 48
rect 259 47 269 48
rect 274 47 286 48
rect 292 47 298 48
rect 310 47 315 48
rect 320 48 326 49
rect 338 48 339 49
rect 353 48 356 49
rect 360 48 363 49
rect 367 48 409 50
rect 320 47 325 48
rect 337 47 338 48
rect 353 47 355 48
rect 360 47 362 48
rect 219 46 224 47
rect 229 46 234 47
rect 75 45 76 46
rect 116 45 117 46
rect 128 45 129 46
rect 143 45 144 46
rect 165 45 185 46
rect 193 45 197 46
rect 206 45 212 46
rect 220 45 221 46
rect 228 45 234 46
rect 240 46 243 47
rect 261 46 268 47
rect 275 46 285 47
rect 292 46 300 47
rect 312 46 315 47
rect 319 46 323 47
rect 336 46 338 47
rect 352 46 353 47
rect 359 46 362 47
rect 240 45 246 46
rect 74 44 75 45
rect 85 44 86 45
rect 107 44 108 45
rect 115 44 117 45
rect 127 44 129 45
rect 135 44 136 45
rect 148 44 149 45
rect 164 44 185 45
rect 60 43 68 44
rect 73 43 75 44
rect 84 43 87 44
rect 95 43 96 44
rect 105 43 109 44
rect 114 43 117 44
rect 125 43 129 44
rect 134 43 137 44
rect 147 43 150 44
rect 162 43 185 44
rect 192 43 197 45
rect 205 43 212 45
rect 227 44 233 45
rect 240 44 249 45
rect 262 44 267 46
rect 275 45 284 46
rect 226 43 232 44
rect 240 43 251 44
rect 263 43 267 44
rect 274 44 284 45
rect 291 45 301 46
rect 313 45 315 46
rect 320 45 321 46
rect 336 45 337 46
rect 345 45 346 46
rect 358 45 362 46
rect 291 44 303 45
rect 274 43 283 44
rect 291 43 304 44
rect 58 42 68 43
rect 72 42 75 43
rect 82 42 88 43
rect 93 42 96 43
rect 104 42 109 43
rect 113 42 118 43
rect 123 42 130 43
rect 133 42 138 43
rect 146 42 152 43
rect 161 42 186 43
rect 191 42 198 43
rect 204 42 212 43
rect 224 42 232 43
rect 239 42 254 43
rect 263 42 268 43
rect 273 42 283 43
rect 289 42 306 43
rect 314 42 315 45
rect 326 44 327 45
rect 335 44 337 45
rect 344 44 346 45
rect 357 44 362 45
rect 325 43 328 44
rect 334 43 336 44
rect 343 43 346 44
rect 355 43 362 44
rect 368 43 409 48
rect 324 42 329 43
rect 333 42 336 43
rect 342 42 346 43
rect 354 42 363 43
rect 367 42 409 43
rect 57 41 76 42
rect 80 41 97 42
rect 102 41 139 42
rect 144 41 187 42
rect 189 41 198 42
rect 203 41 213 42
rect 223 41 232 42
rect 238 41 256 42
rect 263 41 308 42
rect 314 41 316 42
rect 322 41 337 42
rect 341 41 346 42
rect 352 41 409 42
rect 55 40 199 41
rect 202 40 215 41
rect 221 40 232 41
rect 237 40 258 41
rect 262 40 310 41
rect 314 40 409 41
rect 3 39 233 40
rect 234 39 409 40
rect 3 2 409 39
<< metal3 >>
rect 5 139 411 358
rect 5 138 208 139
rect 228 138 411 139
rect 5 137 200 138
rect 244 137 411 138
rect 5 136 196 137
rect 253 136 411 137
rect 5 135 191 136
rect 262 135 411 136
rect 5 134 188 135
rect 269 134 411 135
rect 5 133 184 134
rect 189 133 192 134
rect 210 133 227 134
rect 276 133 411 134
rect 5 132 181 133
rect 186 132 192 133
rect 205 132 236 133
rect 283 132 411 133
rect 5 131 179 132
rect 183 131 191 132
rect 201 131 243 132
rect 288 131 411 132
rect 5 130 175 131
rect 180 130 189 131
rect 198 130 249 131
rect 294 130 411 131
rect 5 129 173 130
rect 178 129 187 130
rect 195 129 254 130
rect 299 129 411 130
rect 5 128 170 129
rect 175 128 185 129
rect 192 128 258 129
rect 305 128 411 129
rect 5 127 168 128
rect 173 127 183 128
rect 190 127 262 128
rect 310 127 411 128
rect 5 126 166 127
rect 170 126 181 127
rect 187 126 266 127
rect 314 126 411 127
rect 5 125 163 126
rect 167 125 179 126
rect 185 125 268 126
rect 319 125 411 126
rect 5 124 161 125
rect 165 124 178 125
rect 183 124 271 125
rect 323 124 411 125
rect 5 123 159 124
rect 162 123 176 124
rect 181 123 272 124
rect 328 123 411 124
rect 5 122 157 123
rect 160 122 174 123
rect 179 122 273 123
rect 332 122 411 123
rect 5 121 155 122
rect 157 121 172 122
rect 177 121 274 122
rect 337 121 411 122
rect 5 120 153 121
rect 155 120 170 121
rect 175 120 272 121
rect 341 120 411 121
rect 5 119 151 120
rect 152 119 169 120
rect 174 119 269 120
rect 345 119 411 120
rect 5 118 167 119
rect 172 118 264 119
rect 291 118 304 119
rect 349 118 411 119
rect 5 117 165 118
rect 170 117 260 118
rect 279 117 286 118
rect 291 117 322 118
rect 353 117 411 118
rect 5 116 163 117
rect 169 116 254 117
rect 272 116 285 117
rect 291 116 337 117
rect 357 116 411 117
rect 5 115 161 116
rect 167 115 248 116
rect 266 115 284 116
rect 290 115 348 116
rect 360 115 411 116
rect 5 114 159 115
rect 165 114 241 115
rect 260 114 283 115
rect 289 114 360 115
rect 363 114 411 115
rect 5 113 158 114
rect 164 113 233 114
rect 255 113 282 114
rect 289 113 411 114
rect 5 112 156 113
rect 162 112 224 113
rect 249 112 281 113
rect 288 112 411 113
rect 5 111 154 112
rect 161 111 210 112
rect 244 111 280 112
rect 286 111 411 112
rect 5 110 112 111
rect 238 110 279 111
rect 285 110 411 111
rect 5 109 105 110
rect 231 109 278 110
rect 283 109 411 110
rect 5 108 101 109
rect 224 108 277 109
rect 281 108 411 109
rect 5 107 97 108
rect 213 107 276 108
rect 278 107 411 108
rect 5 106 94 107
rect 201 106 411 107
rect 5 105 91 106
rect 110 105 304 106
rect 314 105 411 106
rect 5 104 88 105
rect 105 104 300 105
rect 318 104 411 105
rect 5 103 85 104
rect 100 103 112 104
rect 123 103 298 104
rect 320 103 411 104
rect 5 102 82 103
rect 96 102 108 103
rect 127 102 296 103
rect 301 102 317 103
rect 323 102 411 103
rect 5 101 80 102
rect 93 101 106 102
rect 116 101 119 102
rect 129 101 294 102
rect 299 101 320 102
rect 324 101 411 102
rect 5 100 77 101
rect 89 100 104 101
rect 110 100 126 101
rect 131 100 293 101
rect 296 100 322 101
rect 325 100 411 101
rect 5 99 75 100
rect 86 99 103 100
rect 107 99 129 100
rect 133 99 292 100
rect 294 99 324 100
rect 327 99 411 100
rect 5 98 73 99
rect 82 98 101 99
rect 105 98 131 99
rect 134 98 291 99
rect 293 98 326 99
rect 328 98 411 99
rect 5 97 70 98
rect 79 97 100 98
rect 103 97 133 98
rect 135 97 290 98
rect 291 97 327 98
rect 329 97 411 98
rect 5 96 68 97
rect 77 96 99 97
rect 101 96 134 97
rect 136 96 289 97
rect 290 96 328 97
rect 330 96 411 97
rect 5 95 65 96
rect 73 95 98 96
rect 100 95 136 96
rect 137 95 288 96
rect 289 95 329 96
rect 5 94 63 95
rect 71 94 97 95
rect 99 94 137 95
rect 138 94 287 95
rect 288 94 330 95
rect 331 94 411 96
rect 5 93 61 94
rect 68 93 96 94
rect 5 92 59 93
rect 65 92 96 93
rect 97 93 138 94
rect 139 93 331 94
rect 332 93 411 94
rect 97 92 139 93
rect 140 92 332 93
rect 333 92 411 93
rect 5 91 57 92
rect 62 91 95 92
rect 96 91 411 92
rect 5 90 55 91
rect 59 90 411 91
rect 5 89 53 90
rect 57 89 411 90
rect 5 88 51 89
rect 54 88 411 89
rect 5 87 49 88
rect 52 87 411 88
rect 5 86 47 87
rect 49 86 411 87
rect 5 85 45 86
rect 46 85 411 86
rect 5 70 411 85
rect 5 69 197 70
rect 203 69 375 70
rect 378 69 411 70
rect 5 68 56 69
rect 70 68 194 69
rect 204 68 213 69
rect 217 68 228 69
rect 232 68 248 69
rect 264 68 299 69
rect 306 68 374 69
rect 5 67 48 68
rect 71 67 86 68
rect 89 67 149 68
rect 153 67 191 68
rect 206 67 212 68
rect 219 67 227 68
rect 233 67 240 68
rect 267 67 294 68
rect 308 67 318 68
rect 5 66 46 67
rect 72 66 85 67
rect 89 66 147 67
rect 153 66 189 67
rect 206 66 211 67
rect 219 66 225 67
rect 234 66 238 67
rect 268 66 290 67
rect 309 66 316 67
rect 322 66 373 68
rect 380 66 411 69
rect 5 64 44 66
rect 73 65 83 66
rect 89 65 146 66
rect 152 65 187 66
rect 206 65 210 66
rect 220 65 224 66
rect 234 65 237 66
rect 269 65 288 66
rect 309 65 314 66
rect 73 64 82 65
rect 89 64 144 65
rect 152 64 185 65
rect 206 64 209 65
rect 219 64 223 65
rect 5 61 43 64
rect 73 63 81 64
rect 89 63 143 64
rect 151 63 185 64
rect 199 63 200 64
rect 206 63 208 64
rect 219 63 222 64
rect 234 63 236 65
rect 269 64 286 65
rect 309 64 312 65
rect 322 64 372 66
rect 379 64 411 66
rect 269 63 285 64
rect 308 63 311 64
rect 321 63 371 64
rect 73 62 80 63
rect 88 62 142 63
rect 150 62 184 63
rect 197 62 200 63
rect 60 61 67 62
rect 73 61 79 62
rect 87 61 141 62
rect 149 61 184 62
rect 195 61 200 62
rect 205 62 207 63
rect 219 62 221 63
rect 233 62 235 63
rect 253 62 263 63
rect 205 61 206 62
rect 218 61 220 62
rect 232 61 235 62
rect 247 61 264 62
rect 5 58 42 61
rect 54 60 67 61
rect 72 60 78 61
rect 86 60 140 61
rect 148 60 184 61
rect 193 60 199 61
rect 210 60 211 61
rect 217 60 219 61
rect 51 59 66 60
rect 71 59 77 60
rect 86 59 139 60
rect 147 59 184 60
rect 53 58 65 59
rect 70 58 76 59
rect 85 58 138 59
rect 146 58 184 59
rect 194 59 199 60
rect 209 59 210 60
rect 217 59 218 60
rect 231 59 234 61
rect 244 60 248 61
rect 252 60 263 61
rect 269 60 284 63
rect 299 62 302 63
rect 307 62 309 63
rect 320 62 371 63
rect 378 62 411 64
rect 296 60 301 62
rect 315 61 316 62
rect 319 61 371 62
rect 377 61 411 62
rect 313 60 327 61
rect 194 58 198 59
rect 208 58 210 59
rect 216 58 217 59
rect 230 58 234 59
rect 245 59 247 60
rect 251 59 262 60
rect 269 59 283 60
rect 296 59 300 60
rect 311 59 326 60
rect 331 59 370 61
rect 376 59 411 61
rect 245 58 246 59
rect 5 57 43 58
rect 53 57 64 58
rect 69 57 75 58
rect 84 57 137 58
rect 145 57 161 58
rect 164 57 184 58
rect 191 57 197 58
rect 207 57 209 58
rect 215 57 216 58
rect 229 57 246 58
rect 250 58 261 59
rect 268 58 283 59
rect 293 58 299 59
rect 309 58 325 59
rect 250 57 258 58
rect 267 57 284 58
rect 289 57 298 58
rect 307 57 325 58
rect 331 57 369 59
rect 375 57 411 59
rect 5 55 63 57
rect 68 55 74 57
rect 83 56 136 57
rect 144 56 159 57
rect 165 56 197 57
rect 206 56 208 57
rect 82 55 99 56
rect 107 55 126 56
rect 129 55 136 56
rect 143 55 146 56
rect 5 54 62 55
rect 67 54 73 55
rect 81 54 97 55
rect 108 54 117 55
rect 121 54 124 55
rect 130 54 135 55
rect 142 54 144 55
rect 151 54 158 56
rect 5 53 61 54
rect 5 52 60 53
rect 66 52 72 54
rect 80 53 83 54
rect 86 53 95 54
rect 108 53 115 54
rect 122 53 123 54
rect 79 52 81 53
rect 88 52 93 53
rect 5 50 59 52
rect 65 51 71 52
rect 64 50 71 51
rect 78 51 80 52
rect 88 51 92 52
rect 108 51 114 53
rect 121 52 122 53
rect 130 52 134 54
rect 141 53 143 54
rect 152 53 158 54
rect 165 55 196 56
rect 205 55 208 56
rect 219 56 221 57
rect 228 56 245 57
rect 249 56 255 57
rect 266 56 297 57
rect 305 56 325 57
rect 330 56 368 57
rect 219 55 220 56
rect 227 55 244 56
rect 249 55 252 56
rect 265 55 295 56
rect 303 55 325 56
rect 329 55 345 56
rect 350 55 355 56
rect 357 55 368 56
rect 374 55 411 57
rect 165 54 195 55
rect 204 54 207 55
rect 218 54 219 55
rect 227 54 243 55
rect 263 54 293 55
rect 165 53 194 54
rect 203 53 206 54
rect 217 53 219 54
rect 226 53 242 54
rect 260 53 293 54
rect 301 54 323 55
rect 326 54 335 55
rect 340 54 344 55
rect 350 54 354 55
rect 358 54 368 55
rect 301 53 321 54
rect 327 53 334 54
rect 340 53 343 54
rect 350 53 352 54
rect 140 52 141 53
rect 152 52 157 53
rect 165 52 193 53
rect 202 52 206 53
rect 216 52 218 53
rect 225 52 239 53
rect 257 52 292 53
rect 301 52 320 53
rect 327 52 333 53
rect 340 52 341 53
rect 350 52 351 53
rect 120 51 121 52
rect 130 51 133 52
rect 139 51 140 52
rect 145 51 146 52
rect 152 51 156 52
rect 78 50 79 51
rect 87 50 91 51
rect 100 50 101 51
rect 108 50 113 51
rect 119 50 120 51
rect 129 50 132 51
rect 138 50 139 51
rect 144 50 146 51
rect 151 50 155 51
rect 159 50 160 51
rect 5 49 58 50
rect 64 49 70 50
rect 77 49 78 50
rect 87 49 90 50
rect 98 49 100 50
rect 5 48 57 49
rect 5 46 56 48
rect 63 47 70 49
rect 76 48 77 49
rect 86 48 89 49
rect 96 48 99 49
rect 107 48 112 50
rect 118 49 119 50
rect 117 48 118 49
rect 128 48 132 50
rect 137 49 138 50
rect 143 49 145 50
rect 150 49 154 50
rect 158 49 160 50
rect 165 50 192 52
rect 201 51 205 52
rect 215 51 217 52
rect 200 50 204 51
rect 214 50 217 51
rect 224 50 237 52
rect 252 51 292 52
rect 303 51 319 52
rect 246 50 292 51
rect 304 50 319 51
rect 326 50 332 52
rect 339 51 340 52
rect 349 51 350 52
rect 338 50 339 51
rect 359 50 367 54
rect 373 50 411 55
rect 165 49 191 50
rect 200 49 203 50
rect 213 49 216 50
rect 223 49 236 50
rect 250 49 292 50
rect 306 49 318 50
rect 325 49 331 50
rect 337 49 338 50
rect 358 49 367 50
rect 372 49 411 50
rect 136 48 137 49
rect 142 48 144 49
rect 150 48 153 49
rect 157 48 159 49
rect 75 47 76 48
rect 85 47 89 48
rect 95 47 98 48
rect 106 47 110 48
rect 127 47 130 48
rect 141 47 143 48
rect 149 47 151 48
rect 156 47 159 48
rect 165 48 190 49
rect 199 48 202 49
rect 212 48 215 49
rect 165 47 168 48
rect 169 47 189 48
rect 198 47 202 48
rect 211 47 215 48
rect 222 48 235 49
rect 253 48 291 49
rect 307 48 317 49
rect 324 48 331 49
rect 357 48 367 49
rect 371 48 411 49
rect 222 47 231 48
rect 233 47 236 48
rect 257 47 290 48
rect 296 47 297 48
rect 309 47 317 48
rect 323 47 330 48
rect 356 47 360 48
rect 362 47 368 48
rect 63 46 69 47
rect 74 46 75 47
rect 85 46 88 47
rect 94 46 97 47
rect 105 46 109 47
rect 126 46 129 47
rect 147 46 150 47
rect 155 46 159 47
rect 164 46 166 47
rect 169 46 188 47
rect 197 46 201 47
rect 5 45 55 46
rect 5 43 54 45
rect 5 38 53 43
rect 62 42 69 46
rect 84 45 86 46
rect 93 45 96 46
rect 105 45 107 46
rect 125 45 127 46
rect 146 45 149 46
rect 155 45 158 46
rect 163 45 165 46
rect 169 45 187 46
rect 93 44 95 45
rect 104 44 105 45
rect 144 44 148 45
rect 162 44 163 45
rect 168 44 186 45
rect 196 44 200 46
rect 210 45 214 47
rect 222 46 229 47
rect 233 46 238 47
rect 259 46 289 47
rect 295 46 299 47
rect 311 46 317 47
rect 209 44 214 45
rect 221 45 227 46
rect 233 45 237 46
rect 261 45 271 46
rect 276 45 288 46
rect 294 45 300 46
rect 312 45 317 46
rect 322 46 328 47
rect 340 46 341 47
rect 355 46 358 47
rect 362 46 365 47
rect 369 46 411 48
rect 322 45 327 46
rect 339 45 340 46
rect 355 45 357 46
rect 362 45 364 46
rect 221 44 226 45
rect 231 44 236 45
rect 77 43 78 44
rect 118 43 119 44
rect 130 43 131 44
rect 145 43 146 44
rect 167 43 187 44
rect 195 43 199 44
rect 208 43 214 44
rect 222 43 223 44
rect 230 43 236 44
rect 242 44 245 45
rect 263 44 270 45
rect 277 44 287 45
rect 294 44 302 45
rect 314 44 317 45
rect 321 44 325 45
rect 338 44 340 45
rect 354 44 355 45
rect 361 44 364 45
rect 242 43 248 44
rect 76 42 77 43
rect 87 42 88 43
rect 109 42 110 43
rect 117 42 119 43
rect 129 42 131 43
rect 137 42 138 43
rect 150 42 151 43
rect 166 42 187 43
rect 62 41 70 42
rect 75 41 77 42
rect 86 41 89 42
rect 97 41 98 42
rect 107 41 111 42
rect 116 41 119 42
rect 127 41 131 42
rect 136 41 139 42
rect 149 41 152 42
rect 164 41 187 42
rect 194 41 199 43
rect 207 41 214 43
rect 229 42 235 43
rect 242 42 251 43
rect 264 42 269 44
rect 277 43 286 44
rect 228 41 234 42
rect 242 41 253 42
rect 265 41 269 42
rect 276 42 286 43
rect 293 43 303 44
rect 315 43 317 44
rect 322 43 323 44
rect 338 43 339 44
rect 347 43 348 44
rect 360 43 364 44
rect 293 42 305 43
rect 276 41 285 42
rect 293 41 306 42
rect 60 40 70 41
rect 74 40 77 41
rect 84 40 90 41
rect 95 40 98 41
rect 106 40 111 41
rect 115 40 120 41
rect 125 40 132 41
rect 135 40 140 41
rect 148 40 154 41
rect 163 40 188 41
rect 193 40 200 41
rect 206 40 214 41
rect 226 40 234 41
rect 241 40 256 41
rect 265 40 270 41
rect 275 40 285 41
rect 291 40 308 41
rect 316 40 317 43
rect 328 42 329 43
rect 337 42 339 43
rect 346 42 348 43
rect 359 42 364 43
rect 327 41 330 42
rect 336 41 338 42
rect 345 41 348 42
rect 357 41 364 42
rect 370 41 411 46
rect 326 40 331 41
rect 335 40 338 41
rect 344 40 348 41
rect 356 40 365 41
rect 369 40 411 41
rect 59 39 78 40
rect 82 39 99 40
rect 104 39 141 40
rect 146 39 189 40
rect 191 39 200 40
rect 205 39 215 40
rect 225 39 234 40
rect 240 39 258 40
rect 265 39 310 40
rect 316 39 318 40
rect 324 39 339 40
rect 343 39 348 40
rect 354 39 411 40
rect 57 38 201 39
rect 204 38 217 39
rect 223 38 234 39
rect 239 38 260 39
rect 264 38 312 39
rect 316 38 411 39
rect 5 37 235 38
rect 236 37 411 38
rect 5 0 411 37
<< end >>
