magic
tech scmos
magscale 1 30
timestamp 1725930584
<< checkpaint >>
rect -229 25660 2111 25670
rect -600 25645 2400 25660
rect -600 23455 3786 25645
rect -660 20400 3786 23455
rect -600 19795 3786 20400
rect -660 11805 3786 19795
rect -735 10515 3786 11805
rect -600 -590 3786 10515
rect -570 -600 3786 -590
rect -229 -604 3786 -600
rect -175 -606 3786 -604
rect 1516 -615 3786 -606
<< nwell >>
rect -60 21000 1860 22855
rect -60 11205 1860 19195
<< psubstratepdiff >>
rect 30 23400 1770 25060
rect 30 0 1770 7800
<< nsubstratendiff >>
rect 30 21100 1770 22760
rect 30 11290 1770 19100
<< metal1 >>
rect 30 23400 1770 25060
rect 30 21100 1770 22760
rect 30 11290 1770 19100
rect 30 0 1770 7800
<< metal2 >>
rect 30 23400 1770 25060
rect 30 21100 1770 22760
rect 30 11290 1770 19100
rect 30 0 1770 7800
<< metal3 >>
rect 30 23400 1770 25060
rect 30 21100 1770 22760
rect 30 11290 1770 19100
rect 30 0 1770 7800
use IOFILLER10  IOFILLER10_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1537935238
transform 1 0 460 0 1 0
box -35 0 1035 25060
<< end >>
