magic
tech scmos
magscale 1 3
timestamp 1537935238
<< checkpaint >>
rect -60 -975 1260 2590
<< metal2 >>
rect 126 2516 1074 2530
use METAL_RING  METAL_RING_0
timestamp 1537935238
transform 1 0 0 0 1 0
box 0 0 1200 2506
use NDRV1  NDRV1_0
timestamp 1537935238
transform 1 0 126 0 1 1560
box 0 0 948 780
use NDRV1  NDRV1_1
timestamp 1537935238
transform 1 0 126 0 1 780
box 0 0 948 780
use NDRV1  NDRV1_2
timestamp 1537935238
transform 1 0 126 0 1 0
box 0 0 948 780
use PAD_80  PAD_80_0
timestamp 1537935238
transform 1 0 600 0 1 -490
box -425 -425 425 490
use PAD_METAL_PVSS  PAD_METAL_PVSS_0
timestamp 1537935238
transform 1 0 0 0 1 0
box 126 -1 1074 2530
<< labels >>
flabel space 600 -490 600 -490 0 FreeSans 500 0 0 0 VSS
flabel m3p s 0 2195 0 2195 0 FreeSans 500 0 0 0 VDD
flabel m3p s 0 1463 0 1463 0 FreeSans 500 0 0 0 VDD
flabel m3p s 0 2400 0 2400 0 FreeSans 500 0 0 0 VSS
flabel m3p s 0 350 0 350 0 FreeSans 500 0 0 0 VSS
flabel m2p s 575 2530 575 2530 0 FreeSans 500 0 0 0 VSS
<< end >>
