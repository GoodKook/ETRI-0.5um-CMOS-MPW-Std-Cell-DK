magic
tech scmos
magscale 1 30
timestamp 1725924400
<< checkpaint >>
rect -25900 -9750 114735 26213
use IOFILLER1  IOFILLER1_0
timestamp 1537935238
transform 1 0 114000 0 1 0
box -35 0 135 25060
use IOFILLER10  IOFILLER10_0
timestamp 1537935238
transform 1 0 113000 0 1 0
box -35 0 1035 25060
use IOFILLER50  IOFILLER50_0
timestamp 1537935238
transform 1 0 108000 0 1 0
box -35 0 5035 25060
use PANA  PANA_0
timestamp 1537935238
transform 1 0 96000 0 1 0
box -100 -9150 12095 25300
use PBCT4  PBCT4_0
timestamp 1537935238
transform 1 0 24000 0 1 0
box -100 -9150 12100 25351
use PBCT8  PBCT8_0
timestamp 1537935238
transform 1 0 72000 0 1 0
box -100 -9150 12100 25351
use PCORNER  PCORNER_0
timestamp 1537935238
transform 1 0 -25300 0 1 0
box 0 0 25300 25300
use PIC  PIC_0
timestamp 1537935238
transform 1 0 84000 0 1 0
box -100 -9150 12100 25300
use POB4  POB4_0
timestamp 1537935238
transform 1 0 12000 0 1 0
box -100 -9150 12100 25300
use POB8  POB8_0
timestamp 1537935238
transform 1 0 60000 0 1 0
box -100 -9150 12100 25300
use POB24  POB24_0
timestamp 1537935238
transform 1 0 0 0 1 0
box -100 -9150 12100 25300
use PVDD  PVDD_0
timestamp 1537935238
transform 1 0 36000 0 1 0
box 0 -9150 12000 25300
use PVSS  PVSS_0
timestamp 1537935238
transform 1 0 48000 0 1 0
box 0 -9150 12000 25300
<< labels >>
flabel space 102000 -4900 102000 -4900 0 FreeSans 10000 0 0 0 PAD6
flabel space 90000 -4900 90000 -4900 0 FreeSans 10000 0 0 0 PAD5
flabel space 78000 -4900 78000 -4900 0 FreeSans 10000 0 0 0 PAD4
flabel space 66000 -4900 66000 -4900 0 FreeSans 10000 0 0 0 PAD3
flabel space 54000 -4900 54000 -4900 0 FreeSans 10000 0 0 0 VSS
flabel space 42000 -4900 42000 -4900 0 FreeSans 10000 0 0 0 VDD
flabel space 30000 -4900 30000 -4900 0 FreeSans 10000 0 0 0 PAD2
flabel space 18000 -4900 18000 -4900 0 FreeSans 10000 0 0 0 PAD1
flabel space 6000 -4900 6000 -4900 0 FreeSans 10000 0 0 0 PAD0
<< end >>
